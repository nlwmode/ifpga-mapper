module top (\CarrierSense_Tx2_reg/NET0131 , \Collision_Tx1_reg/NET0131 , \Collision_Tx2_reg/NET0131 , \RstTxPauseRq_reg/NET0131 , \RxAbortRst_reg/NET0131 , \RxAbort_latch_reg/NET0131 , \RxAbort_wb_reg/NET0131 , \RxEnSync_reg/NET0131 , \TPauseRq_reg/NET0131 , \TxPauseRq_sync2_reg/NET0131 , \TxPauseRq_sync3_reg/NET0131 , \WillSendControlFrame_sync2_reg/NET0131 , \WillSendControlFrame_sync3_reg/NET0131 , \WillTransmit_q2_reg/P0001 , \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 , \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 , \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 , \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 , \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[0]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[1]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[2]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[3]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[4]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[5]/NET0131 , \ethreg1_IPGT_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 , \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 , \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 , \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 , \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131 , \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 , \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 , \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 , \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131 , \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 , \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 , \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 , \ethreg1_MODER_0_DataOut_reg[0]/NET0131 , \ethreg1_MODER_0_DataOut_reg[1]/NET0131 , \ethreg1_MODER_0_DataOut_reg[2]/NET0131 , \ethreg1_MODER_0_DataOut_reg[3]/NET0131 , \ethreg1_MODER_0_DataOut_reg[4]/NET0131 , \ethreg1_MODER_0_DataOut_reg[5]/NET0131 , \ethreg1_MODER_0_DataOut_reg[6]/NET0131 , \ethreg1_MODER_0_DataOut_reg[7]/NET0131 , \ethreg1_MODER_1_DataOut_reg[0]/NET0131 , \ethreg1_MODER_1_DataOut_reg[1]/NET0131 , \ethreg1_MODER_1_DataOut_reg[2]/NET0131 , \ethreg1_MODER_1_DataOut_reg[3]/NET0131 , \ethreg1_MODER_1_DataOut_reg[4]/NET0131 , \ethreg1_MODER_1_DataOut_reg[5]/NET0131 , \ethreg1_MODER_1_DataOut_reg[6]/NET0131 , \ethreg1_MODER_1_DataOut_reg[7]/NET0131 , \ethreg1_MODER_2_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 , \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 , \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 , \ethreg1_ResetRxCIrq_sync2_reg/NET0131 , \ethreg1_ResetRxCIrq_sync3_reg/NET0131 , \ethreg1_ResetTxCIrq_sync2_reg/NET0131 , \ethreg1_SetRxCIrq_reg/NET0131 , \ethreg1_SetRxCIrq_rxclk_reg/NET0131 , \ethreg1_SetRxCIrq_sync2_reg/NET0131 , \ethreg1_SetRxCIrq_sync3_reg/NET0131 , \ethreg1_SetTxCIrq_reg/NET0131 , \ethreg1_SetTxCIrq_sync2_reg/NET0131 , \ethreg1_SetTxCIrq_sync3_reg/NET0131 , \ethreg1_SetTxCIrq_txclk_reg/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 , \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 , \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 , \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 , \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 , \ethreg1_irq_busy_reg/NET0131 , \ethreg1_irq_rxb_reg/NET0131 , \ethreg1_irq_rxc_reg/NET0131 , \ethreg1_irq_rxe_reg/NET0131 , \ethreg1_irq_txb_reg/NET0131 , \ethreg1_irq_txc_reg/NET0131 , \ethreg1_irq_txe_reg/NET0131 , m_wb_ack_i_pad, \m_wb_adr_o[10]_pad , \m_wb_adr_o[11]_pad , \m_wb_adr_o[12]_pad , \m_wb_adr_o[13]_pad , \m_wb_adr_o[14]_pad , \m_wb_adr_o[15]_pad , \m_wb_adr_o[16]_pad , \m_wb_adr_o[17]_pad , \m_wb_adr_o[18]_pad , \m_wb_adr_o[19]_pad , \m_wb_adr_o[20]_pad , \m_wb_adr_o[21]_pad , \m_wb_adr_o[22]_pad , \m_wb_adr_o[23]_pad , \m_wb_adr_o[24]_pad , \m_wb_adr_o[25]_pad , \m_wb_adr_o[26]_pad , \m_wb_adr_o[27]_pad , \m_wb_adr_o[28]_pad , \m_wb_adr_o[29]_pad , \m_wb_adr_o[2]_pad , \m_wb_adr_o[30]_pad , \m_wb_adr_o[31]_pad , \m_wb_adr_o[3]_pad , \m_wb_adr_o[4]_pad , \m_wb_adr_o[5]_pad , \m_wb_adr_o[6]_pad , \m_wb_adr_o[7]_pad , \m_wb_adr_o[8]_pad , \m_wb_adr_o[9]_pad , \m_wb_dat_i[10]_pad , \m_wb_dat_i[11]_pad , \m_wb_dat_i[12]_pad , \m_wb_dat_i[13]_pad , \m_wb_dat_i[14]_pad , \m_wb_dat_i[15]_pad , \m_wb_dat_i[16]_pad , \m_wb_dat_i[17]_pad , \m_wb_dat_i[18]_pad , \m_wb_dat_i[19]_pad , \m_wb_dat_i[1]_pad , \m_wb_dat_i[20]_pad , \m_wb_dat_i[22]_pad , \m_wb_dat_i[23]_pad , \m_wb_dat_i[24]_pad , \m_wb_dat_i[25]_pad , \m_wb_dat_i[26]_pad , \m_wb_dat_i[27]_pad , \m_wb_dat_i[28]_pad , \m_wb_dat_i[29]_pad , \m_wb_dat_i[2]_pad , \m_wb_dat_i[30]_pad , \m_wb_dat_i[31]_pad , \m_wb_dat_i[3]_pad , \m_wb_dat_i[4]_pad , \m_wb_dat_i[5]_pad , \m_wb_dat_i[6]_pad , \m_wb_dat_i[7]_pad , \m_wb_dat_i[8]_pad , m_wb_err_i_pad, \m_wb_sel_o[0]_pad , \m_wb_sel_o[1]_pad , \m_wb_sel_o[2]_pad , \m_wb_sel_o[3]_pad , m_wb_stb_o_pad, m_wb_we_o_pad, \maccontrol1_MuxedAbort_reg/NET0131 , \maccontrol1_MuxedDone_reg/NET0131 , \maccontrol1_TxAbortInLatched_reg/NET0131 , \maccontrol1_TxDoneInLatched_reg/NET0131 , \maccontrol1_TxUsedDataOutDetected_reg/NET0131 , \maccontrol1_receivecontrol1_AddressOK_reg/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 , \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 , \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 , \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 , \maccontrol1_receivecontrol1_Divider2_reg/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 , \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 , \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 , \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 , \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 , \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 , \maccontrol1_receivecontrol1_Pause_reg/NET0131 , \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 , \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 , \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 , \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 , \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 , \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131 , \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131 , \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001 , \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 , \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 , \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001 , \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 , \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131 , \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 , \macstatus1_CarrierSenseLost_reg/NET0131 , \macstatus1_DeferLatched_reg/NET0131 , \macstatus1_DribbleNibble_reg/NET0131 , \macstatus1_InvalidSymbol_reg/NET0131 , \macstatus1_LatchedCrcError_reg/NET0131 , \macstatus1_LatchedMRxErr_reg/NET0131 , \macstatus1_LateCollLatched_reg/P0002 , \macstatus1_LoadRxStatus_reg/NET0131 , \macstatus1_ReceiveEnd_reg/NET0131 , \macstatus1_ReceivedPacketTooBig_reg/NET0131 , \macstatus1_RetryCntLatched_reg[0]/P0002 , \macstatus1_RetryCntLatched_reg[1]/P0002 , \macstatus1_RetryCntLatched_reg[2]/P0002 , \macstatus1_RetryCntLatched_reg[3]/P0002 , \macstatus1_RetryLimit_reg/P0002 , \macstatus1_RxColWindow_reg/NET0131 , \macstatus1_RxLateCollision_reg/NET0131 , \macstatus1_ShortFrame_reg/NET0131 , mcoll_pad_i_pad, md_pad_i_pad, mdc_pad_o_pad, \miim1_BitCounter_reg[0]/NET0131 , \miim1_BitCounter_reg[1]/NET0131 , \miim1_BitCounter_reg[2]/NET0131 , \miim1_BitCounter_reg[3]/NET0131 , \miim1_BitCounter_reg[4]/NET0131 , \miim1_BitCounter_reg[5]/NET0131 , \miim1_BitCounter_reg[6]/NET0131 , \miim1_EndBusy_reg/NET0131 , \miim1_InProgress_q1_reg/NET0131 , \miim1_InProgress_q2_reg/NET0131 , \miim1_InProgress_q3_reg/NET0131 , \miim1_InProgress_reg/NET0131 , \miim1_LatchByte0_d_reg/NET0131 , \miim1_LatchByte1_d_reg/NET0131 , \miim1_LatchByte_reg[0]/NET0131 , \miim1_LatchByte_reg[1]/NET0131 , \miim1_Nvalid_reg/NET0131 , \miim1_RStatStart_q1_reg/NET0131 , \miim1_RStatStart_q2_reg/NET0131 , \miim1_RStatStart_reg/NET0131 , \miim1_RStat_q2_reg/NET0131 , \miim1_RStat_q3_reg/NET0131 , \miim1_ScanStat_q2_reg/NET0131 , \miim1_SyncStatMdcEn_reg/NET0131 , \miim1_WCtrlDataStart_q1_reg/NET0131 , \miim1_WCtrlDataStart_q2_reg/NET0131 , \miim1_WCtrlDataStart_q_reg/NET0131 , \miim1_WCtrlDataStart_reg/NET0131 , \miim1_WCtrlData_q2_reg/NET0131 , \miim1_WCtrlData_q3_reg/NET0131 , \miim1_WriteOp_reg/NET0131 , \miim1_clkgen_Counter_reg[0]/NET0131 , \miim1_clkgen_Counter_reg[1]/NET0131 , \miim1_clkgen_Counter_reg[2]/NET0131 , \miim1_clkgen_Counter_reg[3]/NET0131 , \miim1_clkgen_Counter_reg[4]/NET0131 , \miim1_clkgen_Counter_reg[5]/NET0131 , \miim1_clkgen_Counter_reg[6]/NET0131 , \miim1_outctrl_Mdo_2d_reg/NET0131 , \miim1_shftrg_LinkFail_reg/NET0131 , \miim1_shftrg_ShiftReg_reg[0]/NET0131 , \miim1_shftrg_ShiftReg_reg[1]/NET0131 , \miim1_shftrg_ShiftReg_reg[2]/NET0131 , \miim1_shftrg_ShiftReg_reg[3]/NET0131 , \miim1_shftrg_ShiftReg_reg[4]/NET0131 , \miim1_shftrg_ShiftReg_reg[5]/NET0131 , \miim1_shftrg_ShiftReg_reg[6]/NET0131 , \miim1_shftrg_ShiftReg_reg[7]/NET0131 , \mrxd_pad_i[0]_pad , \mrxd_pad_i[1]_pad , \mrxd_pad_i[2]_pad , \mrxd_pad_i[3]_pad , mrxdv_pad_i_pad, mrxerr_pad_i_pad, \mtxd_pad_o[0]_pad , \mtxd_pad_o[1]_pad , \mtxd_pad_o[2]_pad , \mtxd_pad_o[3]_pad , mtxen_pad_o_pad, mtxerr_pad_o_pad, \rxethmac1_Broadcast_reg/NET0131 , \rxethmac1_CrcHashGood_reg/P0001 , \rxethmac1_CrcHash_reg[0]/P0001 , \rxethmac1_CrcHash_reg[1]/P0001 , \rxethmac1_CrcHash_reg[2]/P0001 , \rxethmac1_CrcHash_reg[3]/P0001 , \rxethmac1_CrcHash_reg[4]/P0001 , \rxethmac1_CrcHash_reg[5]/P0001 , \rxethmac1_DelayData_reg/NET0131 , \rxethmac1_LatchedByte_reg[0]/NET0131 , \rxethmac1_LatchedByte_reg[1]/NET0131 , \rxethmac1_LatchedByte_reg[2]/NET0131 , \rxethmac1_LatchedByte_reg[3]/NET0131 , \rxethmac1_LatchedByte_reg[4]/NET0131 , \rxethmac1_LatchedByte_reg[5]/NET0131 , \rxethmac1_LatchedByte_reg[6]/NET0131 , \rxethmac1_LatchedByte_reg[7]/NET0131 , \rxethmac1_Multicast_reg/NET0131 , \rxethmac1_RxData_d_reg[0]/NET0131 , \rxethmac1_RxData_d_reg[1]/NET0131 , \rxethmac1_RxData_d_reg[2]/NET0131 , \rxethmac1_RxData_d_reg[3]/NET0131 , \rxethmac1_RxData_d_reg[4]/NET0131 , \rxethmac1_RxData_d_reg[5]/NET0131 , \rxethmac1_RxData_d_reg[6]/NET0131 , \rxethmac1_RxData_d_reg[7]/NET0131 , \rxethmac1_RxData_reg[0]/NET0131 , \rxethmac1_RxData_reg[1]/NET0131 , \rxethmac1_RxData_reg[2]/NET0131 , \rxethmac1_RxData_reg[3]/NET0131 , \rxethmac1_RxData_reg[4]/NET0131 , \rxethmac1_RxData_reg[5]/NET0131 , \rxethmac1_RxData_reg[6]/NET0131 , \rxethmac1_RxData_reg[7]/NET0131 , \rxethmac1_RxEndFrm_d_reg/NET0131 , \rxethmac1_RxEndFrm_reg/NET0131 , \rxethmac1_RxStartFrm_reg/NET0131 , \rxethmac1_RxValid_reg/NET0131 , \rxethmac1_crcrx_Crc_reg[0]/NET0131 , \rxethmac1_crcrx_Crc_reg[10]/NET0131 , \rxethmac1_crcrx_Crc_reg[11]/NET0131 , \rxethmac1_crcrx_Crc_reg[12]/NET0131 , \rxethmac1_crcrx_Crc_reg[13]/NET0131 , \rxethmac1_crcrx_Crc_reg[14]/NET0131 , \rxethmac1_crcrx_Crc_reg[15]/NET0131 , \rxethmac1_crcrx_Crc_reg[16]/NET0131 , \rxethmac1_crcrx_Crc_reg[17]/NET0131 , \rxethmac1_crcrx_Crc_reg[18]/NET0131 , \rxethmac1_crcrx_Crc_reg[19]/NET0131 , \rxethmac1_crcrx_Crc_reg[1]/NET0131 , \rxethmac1_crcrx_Crc_reg[20]/NET0131 , \rxethmac1_crcrx_Crc_reg[21]/NET0131 , \rxethmac1_crcrx_Crc_reg[22]/NET0131 , \rxethmac1_crcrx_Crc_reg[23]/NET0131 , \rxethmac1_crcrx_Crc_reg[24]/NET0131 , \rxethmac1_crcrx_Crc_reg[25]/NET0131 , \rxethmac1_crcrx_Crc_reg[26]/NET0131 , \rxethmac1_crcrx_Crc_reg[27]/NET0131 , \rxethmac1_crcrx_Crc_reg[28]/NET0131 , \rxethmac1_crcrx_Crc_reg[29]/NET0131 , \rxethmac1_crcrx_Crc_reg[2]/NET0131 , \rxethmac1_crcrx_Crc_reg[30]/NET0131 , \rxethmac1_crcrx_Crc_reg[31]/NET0131 , \rxethmac1_crcrx_Crc_reg[3]/NET0131 , \rxethmac1_crcrx_Crc_reg[4]/NET0131 , \rxethmac1_crcrx_Crc_reg[5]/NET0131 , \rxethmac1_crcrx_Crc_reg[6]/NET0131 , \rxethmac1_crcrx_Crc_reg[7]/NET0131 , \rxethmac1_crcrx_Crc_reg[8]/NET0131 , \rxethmac1_crcrx_Crc_reg[9]/NET0131 , \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131 , \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 , \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 , \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 , \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 , \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 , \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 , \rxethmac1_rxstatem1_StateData0_reg/NET0131 , \rxethmac1_rxstatem1_StateData1_reg/NET0131 , \rxethmac1_rxstatem1_StateDrop_reg/NET0131 , \rxethmac1_rxstatem1_StateIdle_reg/NET0131 , \rxethmac1_rxstatem1_StatePreamble_reg/NET0131 , \rxethmac1_rxstatem1_StateSFD_reg/NET0131 , \txethmac1_ColWindow_reg/NET0131 , \txethmac1_PacketFinished_q_reg/NET0131 , \txethmac1_RetryCnt_reg[0]/NET0131 , \txethmac1_RetryCnt_reg[1]/NET0131 , \txethmac1_RetryCnt_reg[2]/NET0131 , \txethmac1_RetryCnt_reg[3]/NET0131 , \txethmac1_StatusLatch_reg/NET0131 , \txethmac1_StopExcessiveDeferOccured_reg/NET0131 , \txethmac1_TxAbort_reg/NET0131 , \txethmac1_TxDone_reg/NET0131 , \txethmac1_TxRetry_reg/NET0131 , \txethmac1_TxUsedData_reg/NET0131 , \txethmac1_random1_RandomLatched_reg[0]/NET0131 , \txethmac1_random1_RandomLatched_reg[1]/NET0131 , \txethmac1_random1_RandomLatched_reg[2]/NET0131 , \txethmac1_random1_RandomLatched_reg[3]/NET0131 , \txethmac1_random1_RandomLatched_reg[4]/NET0131 , \txethmac1_random1_RandomLatched_reg[5]/NET0131 , \txethmac1_random1_RandomLatched_reg[6]/NET0131 , \txethmac1_random1_RandomLatched_reg[7]/NET0131 , \txethmac1_random1_RandomLatched_reg[8]/NET0131 , \txethmac1_random1_RandomLatched_reg[9]/NET0131 , \txethmac1_random1_x_reg[1]/NET0131 , \txethmac1_random1_x_reg[2]/NET0131 , \txethmac1_random1_x_reg[3]/NET0131 , \txethmac1_random1_x_reg[4]/NET0131 , \txethmac1_random1_x_reg[5]/NET0131 , \txethmac1_random1_x_reg[6]/NET0131 , \txethmac1_random1_x_reg[7]/NET0131 , \txethmac1_random1_x_reg[8]/NET0131 , \txethmac1_random1_x_reg[9]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 , \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 , \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[0]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[10]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[11]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[12]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[13]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[14]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[15]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[1]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[2]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[3]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[4]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[5]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[6]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[7]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[8]/NET0131 , \txethmac1_txcounters1_NibCnt_reg[9]/NET0131 , \txethmac1_txcrc_Crc_reg[0]/NET0131 , \txethmac1_txcrc_Crc_reg[10]/NET0131 , \txethmac1_txcrc_Crc_reg[11]/NET0131 , \txethmac1_txcrc_Crc_reg[12]/NET0131 , \txethmac1_txcrc_Crc_reg[13]/NET0131 , \txethmac1_txcrc_Crc_reg[14]/NET0131 , \txethmac1_txcrc_Crc_reg[15]/NET0131 , \txethmac1_txcrc_Crc_reg[16]/NET0131 , \txethmac1_txcrc_Crc_reg[17]/NET0131 , \txethmac1_txcrc_Crc_reg[18]/NET0131 , \txethmac1_txcrc_Crc_reg[19]/NET0131 , \txethmac1_txcrc_Crc_reg[1]/NET0131 , \txethmac1_txcrc_Crc_reg[20]/NET0131 , \txethmac1_txcrc_Crc_reg[21]/NET0131 , \txethmac1_txcrc_Crc_reg[22]/NET0131 , \txethmac1_txcrc_Crc_reg[23]/NET0131 , \txethmac1_txcrc_Crc_reg[24]/NET0131 , \txethmac1_txcrc_Crc_reg[25]/NET0131 , \txethmac1_txcrc_Crc_reg[26]/NET0131 , \txethmac1_txcrc_Crc_reg[27]/NET0131 , \txethmac1_txcrc_Crc_reg[28]/NET0131 , \txethmac1_txcrc_Crc_reg[29]/NET0131 , \txethmac1_txcrc_Crc_reg[2]/NET0131 , \txethmac1_txcrc_Crc_reg[30]/NET0131 , \txethmac1_txcrc_Crc_reg[31]/NET0131 , \txethmac1_txcrc_Crc_reg[3]/NET0131 , \txethmac1_txcrc_Crc_reg[4]/NET0131 , \txethmac1_txcrc_Crc_reg[5]/NET0131 , \txethmac1_txcrc_Crc_reg[6]/NET0131 , \txethmac1_txcrc_Crc_reg[7]/NET0131 , \txethmac1_txcrc_Crc_reg[8]/NET0131 , \txethmac1_txcrc_Crc_reg[9]/NET0131 , \txethmac1_txstatem1_Rule1_reg/NET0131 , \txethmac1_txstatem1_StateBackOff_reg/NET0131 , \txethmac1_txstatem1_StateData_reg[0]/NET0131 , \txethmac1_txstatem1_StateData_reg[1]/NET0131 , \txethmac1_txstatem1_StateDefer_reg/NET0131 , \txethmac1_txstatem1_StateFCS_reg/NET0131 , \txethmac1_txstatem1_StateIPG_reg/NET0131 , \txethmac1_txstatem1_StateIdle_reg/NET0131 , \txethmac1_txstatem1_StateJam_q_reg/NET0131 , \txethmac1_txstatem1_StateJam_reg/NET0131 , \txethmac1_txstatem1_StatePAD_reg/NET0131 , \txethmac1_txstatem1_StatePreamble_reg/NET0131 , wb_ack_o_pad, \wb_adr_i[10]_pad , \wb_adr_i[11]_pad , \wb_adr_i[2]_pad , \wb_adr_i[3]_pad , \wb_adr_i[4]_pad , \wb_adr_i[5]_pad , \wb_adr_i[6]_pad , \wb_adr_i[7]_pad , \wb_adr_i[8]_pad , \wb_adr_i[9]_pad , wb_cyc_i_pad, \wb_dat_i[0]_pad , \wb_dat_i[10]_pad , \wb_dat_i[11]_pad , \wb_dat_i[12]_pad , \wb_dat_i[13]_pad , \wb_dat_i[14]_pad , \wb_dat_i[15]_pad , \wb_dat_i[16]_pad , \wb_dat_i[17]_pad , \wb_dat_i[18]_pad , \wb_dat_i[19]_pad , \wb_dat_i[1]_pad , \wb_dat_i[20]_pad , \wb_dat_i[21]_pad , \wb_dat_i[22]_pad , \wb_dat_i[23]_pad , \wb_dat_i[24]_pad , \wb_dat_i[25]_pad , \wb_dat_i[26]_pad , \wb_dat_i[27]_pad , \wb_dat_i[28]_pad , \wb_dat_i[29]_pad , \wb_dat_i[2]_pad , \wb_dat_i[30]_pad , \wb_dat_i[31]_pad , \wb_dat_i[3]_pad , \wb_dat_i[4]_pad , \wb_dat_i[5]_pad , \wb_dat_i[6]_pad , \wb_dat_i[7]_pad , \wb_dat_i[8]_pad , \wb_dat_i[9]_pad , wb_err_o_pad, wb_rst_i_pad, \wb_sel_i[0]_pad , \wb_sel_i[1]_pad , \wb_sel_i[2]_pad , \wb_sel_i[3]_pad , wb_stb_i_pad, wb_we_i_pad, \wishbone_BDRead_reg/NET0131 , \wishbone_BDWrite_reg[0]/NET0131 , \wishbone_BDWrite_reg[1]/NET0131 , \wishbone_BDWrite_reg[2]/NET0131 , \wishbone_BDWrite_reg[3]/NET0131 , \wishbone_BlockReadTxDataFromMemory_reg/NET0131 , \wishbone_BlockingIncrementTxPointer_reg/NET0131 , \wishbone_BlockingTxBDRead_reg/NET0131 , \wishbone_BlockingTxStatusWrite_reg/NET0131 , \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 , \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131 , \wishbone_Busy_IRQ_rck_reg/NET0131 , \wishbone_Busy_IRQ_sync2_reg/P0001 , \wishbone_Busy_IRQ_sync3_reg/P0001 , \wishbone_Busy_IRQ_syncb2_reg/P0001 , \wishbone_Flop_reg/NET0131 , \wishbone_IncrTxPointer_reg/NET0131 , \wishbone_LastByteIn_reg/NET0131 , \wishbone_LastWord_reg/NET0131 , \wishbone_LatchValidBytes_q_reg/NET0131 , \wishbone_LatchValidBytes_reg/NET0131 , \wishbone_LatchedRxLength_reg[0]/NET0131 , \wishbone_LatchedRxLength_reg[10]/NET0131 , \wishbone_LatchedRxLength_reg[11]/NET0131 , \wishbone_LatchedRxLength_reg[12]/NET0131 , \wishbone_LatchedRxLength_reg[13]/NET0131 , \wishbone_LatchedRxLength_reg[14]/NET0131 , \wishbone_LatchedRxLength_reg[15]/NET0131 , \wishbone_LatchedRxLength_reg[1]/NET0131 , \wishbone_LatchedRxLength_reg[2]/NET0131 , \wishbone_LatchedRxLength_reg[3]/NET0131 , \wishbone_LatchedRxLength_reg[4]/NET0131 , \wishbone_LatchedRxLength_reg[5]/NET0131 , \wishbone_LatchedRxLength_reg[6]/NET0131 , \wishbone_LatchedRxLength_reg[7]/NET0131 , \wishbone_LatchedRxLength_reg[8]/NET0131 , \wishbone_LatchedRxLength_reg[9]/NET0131 , \wishbone_LatchedRxStartFrm_reg/NET0131 , \wishbone_LatchedTxLength_reg[0]/NET0131 , \wishbone_LatchedTxLength_reg[10]/NET0131 , \wishbone_LatchedTxLength_reg[11]/NET0131 , \wishbone_LatchedTxLength_reg[12]/NET0131 , \wishbone_LatchedTxLength_reg[13]/NET0131 , \wishbone_LatchedTxLength_reg[14]/NET0131 , \wishbone_LatchedTxLength_reg[15]/NET0131 , \wishbone_LatchedTxLength_reg[1]/NET0131 , \wishbone_LatchedTxLength_reg[2]/NET0131 , \wishbone_LatchedTxLength_reg[3]/NET0131 , \wishbone_LatchedTxLength_reg[4]/NET0131 , \wishbone_LatchedTxLength_reg[5]/NET0131 , \wishbone_LatchedTxLength_reg[6]/NET0131 , \wishbone_LatchedTxLength_reg[7]/NET0131 , \wishbone_LatchedTxLength_reg[8]/NET0131 , \wishbone_LatchedTxLength_reg[9]/NET0131 , \wishbone_MasterWbRX_reg/NET0131 , \wishbone_MasterWbTX_reg/NET0131 , \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 , \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 , \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131 , \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131 , \wishbone_ReadTxDataFromFifo_tck_reg/NET0131 , \wishbone_ReadTxDataFromMemory_reg/NET0131 , \wishbone_RxAbortLatched_reg/NET0131 , \wishbone_RxAbortSync2_reg/NET0131 , \wishbone_RxAbortSync3_reg/NET0131 , \wishbone_RxAbortSync4_reg/NET0131 , \wishbone_RxAbortSyncb2_reg/NET0131 , \wishbone_RxBDAddress_reg[1]/NET0131 , \wishbone_RxBDAddress_reg[2]/NET0131 , \wishbone_RxBDAddress_reg[3]/NET0131 , \wishbone_RxBDAddress_reg[4]/NET0131 , \wishbone_RxBDAddress_reg[5]/NET0131 , \wishbone_RxBDAddress_reg[6]/NET0131 , \wishbone_RxBDAddress_reg[7]/NET0131 , \wishbone_RxBDRead_reg/NET0131 , \wishbone_RxBDReady_reg/NET0131 , \wishbone_RxB_IRQ_reg/NET0131 , \wishbone_RxByteCnt_reg[0]/NET0131 , \wishbone_RxByteCnt_reg[1]/NET0131 , \wishbone_RxDataLatched1_reg[10]/NET0131 , \wishbone_RxDataLatched1_reg[11]/NET0131 , \wishbone_RxDataLatched1_reg[12]/NET0131 , \wishbone_RxDataLatched1_reg[13]/NET0131 , \wishbone_RxDataLatched1_reg[14]/NET0131 , \wishbone_RxDataLatched1_reg[15]/NET0131 , \wishbone_RxDataLatched1_reg[16]/NET0131 , \wishbone_RxDataLatched1_reg[17]/NET0131 , \wishbone_RxDataLatched1_reg[18]/NET0131 , \wishbone_RxDataLatched1_reg[19]/NET0131 , \wishbone_RxDataLatched1_reg[20]/NET0131 , \wishbone_RxDataLatched1_reg[21]/NET0131 , \wishbone_RxDataLatched1_reg[22]/NET0131 , \wishbone_RxDataLatched1_reg[23]/NET0131 , \wishbone_RxDataLatched1_reg[24]/NET0131 , \wishbone_RxDataLatched1_reg[25]/NET0131 , \wishbone_RxDataLatched1_reg[26]/NET0131 , \wishbone_RxDataLatched1_reg[27]/NET0131 , \wishbone_RxDataLatched1_reg[28]/NET0131 , \wishbone_RxDataLatched1_reg[29]/NET0131 , \wishbone_RxDataLatched1_reg[30]/NET0131 , \wishbone_RxDataLatched1_reg[31]/NET0131 , \wishbone_RxDataLatched1_reg[8]/NET0131 , \wishbone_RxDataLatched1_reg[9]/NET0131 , \wishbone_RxDataLatched2_reg[0]/NET0131 , \wishbone_RxDataLatched2_reg[10]/NET0131 , \wishbone_RxDataLatched2_reg[11]/NET0131 , \wishbone_RxDataLatched2_reg[12]/NET0131 , \wishbone_RxDataLatched2_reg[13]/NET0131 , \wishbone_RxDataLatched2_reg[14]/NET0131 , \wishbone_RxDataLatched2_reg[15]/NET0131 , \wishbone_RxDataLatched2_reg[16]/NET0131 , \wishbone_RxDataLatched2_reg[17]/NET0131 , \wishbone_RxDataLatched2_reg[18]/NET0131 , \wishbone_RxDataLatched2_reg[19]/NET0131 , \wishbone_RxDataLatched2_reg[1]/NET0131 , \wishbone_RxDataLatched2_reg[20]/NET0131 , \wishbone_RxDataLatched2_reg[21]/NET0131 , \wishbone_RxDataLatched2_reg[22]/NET0131 , \wishbone_RxDataLatched2_reg[23]/NET0131 , \wishbone_RxDataLatched2_reg[24]/NET0131 , \wishbone_RxDataLatched2_reg[25]/NET0131 , \wishbone_RxDataLatched2_reg[26]/NET0131 , \wishbone_RxDataLatched2_reg[27]/NET0131 , \wishbone_RxDataLatched2_reg[28]/NET0131 , \wishbone_RxDataLatched2_reg[29]/NET0131 , \wishbone_RxDataLatched2_reg[2]/NET0131 , \wishbone_RxDataLatched2_reg[30]/NET0131 , \wishbone_RxDataLatched2_reg[31]/NET0131 , \wishbone_RxDataLatched2_reg[3]/NET0131 , \wishbone_RxDataLatched2_reg[4]/NET0131 , \wishbone_RxDataLatched2_reg[5]/NET0131 , \wishbone_RxDataLatched2_reg[6]/NET0131 , \wishbone_RxDataLatched2_reg[7]/NET0131 , \wishbone_RxDataLatched2_reg[8]/NET0131 , \wishbone_RxDataLatched2_reg[9]/NET0131 , \wishbone_RxE_IRQ_reg/NET0131 , \wishbone_RxEn_needed_reg/NET0131 , \wishbone_RxEn_q_reg/NET0131 , \wishbone_RxEn_reg/NET0131 , \wishbone_RxEnableWindow_reg/NET0131 , \wishbone_RxOverrun_reg/NET0131 , \wishbone_RxPointerLSB_rst_reg[0]/NET0131 , \wishbone_RxPointerLSB_rst_reg[1]/NET0131 , \wishbone_RxPointerMSB_reg[10]/NET0131 , \wishbone_RxPointerMSB_reg[11]/NET0131 , \wishbone_RxPointerMSB_reg[12]/NET0131 , \wishbone_RxPointerMSB_reg[13]/NET0131 , \wishbone_RxPointerMSB_reg[14]/NET0131 , \wishbone_RxPointerMSB_reg[15]/NET0131 , \wishbone_RxPointerMSB_reg[16]/NET0131 , \wishbone_RxPointerMSB_reg[17]/NET0131 , \wishbone_RxPointerMSB_reg[18]/NET0131 , \wishbone_RxPointerMSB_reg[19]/NET0131 , \wishbone_RxPointerMSB_reg[20]/NET0131 , \wishbone_RxPointerMSB_reg[21]/NET0131 , \wishbone_RxPointerMSB_reg[22]/NET0131 , \wishbone_RxPointerMSB_reg[23]/NET0131 , \wishbone_RxPointerMSB_reg[24]/NET0131 , \wishbone_RxPointerMSB_reg[25]/NET0131 , \wishbone_RxPointerMSB_reg[26]/NET0131 , \wishbone_RxPointerMSB_reg[27]/NET0131 , \wishbone_RxPointerMSB_reg[28]/NET0131 , \wishbone_RxPointerMSB_reg[29]/NET0131 , \wishbone_RxPointerMSB_reg[2]/NET0131 , \wishbone_RxPointerMSB_reg[30]/NET0131 , \wishbone_RxPointerMSB_reg[31]/NET0131 , \wishbone_RxPointerMSB_reg[3]/NET0131 , \wishbone_RxPointerMSB_reg[4]/NET0131 , \wishbone_RxPointerMSB_reg[5]/NET0131 , \wishbone_RxPointerMSB_reg[6]/NET0131 , \wishbone_RxPointerMSB_reg[7]/NET0131 , \wishbone_RxPointerMSB_reg[8]/NET0131 , \wishbone_RxPointerMSB_reg[9]/NET0131 , \wishbone_RxPointerRead_reg/NET0131 , \wishbone_RxReady_reg/NET0131 , \wishbone_RxStatusInLatched_reg[0]/NET0131 , \wishbone_RxStatusInLatched_reg[1]/NET0131 , \wishbone_RxStatusInLatched_reg[2]/NET0131 , \wishbone_RxStatusInLatched_reg[3]/NET0131 , \wishbone_RxStatusInLatched_reg[4]/NET0131 , \wishbone_RxStatusInLatched_reg[5]/NET0131 , \wishbone_RxStatusInLatched_reg[6]/NET0131 , \wishbone_RxStatusInLatched_reg[7]/NET0131 , \wishbone_RxStatusInLatched_reg[8]/NET0131 , \wishbone_RxStatusWriteLatched_reg/NET0131 , \wishbone_RxStatusWriteLatched_sync2_reg/NET0131 , \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131 , \wishbone_RxStatus_reg[13]/NET0131 , \wishbone_RxStatus_reg[14]/NET0131 , \wishbone_RxValidBytes_reg[0]/NET0131 , \wishbone_RxValidBytes_reg[1]/NET0131 , \wishbone_ShiftEndedSync1_reg/NET0131 , \wishbone_ShiftEndedSync2_reg/NET0131 , \wishbone_ShiftEndedSync3_reg/NET0131 , \wishbone_ShiftEndedSync_c1_reg/NET0131 , \wishbone_ShiftEndedSync_c2_reg/NET0131 , \wishbone_ShiftEnded_rck_reg/NET0131 , \wishbone_ShiftEnded_reg/NET0131 , \wishbone_ShiftWillEnd_reg/NET0131 , \wishbone_StartOccured_reg/NET0131 , \wishbone_SyncRxStartFrm_q2_reg/NET0131 , \wishbone_SyncRxStartFrm_q_reg/NET0131 , \wishbone_TxAbortPacketBlocked_reg/NET0131 , \wishbone_TxAbortPacket_NotCleared_reg/NET0131 , \wishbone_TxAbortPacket_reg/NET0131 , \wishbone_TxAbort_q_reg/NET0131 , \wishbone_TxAbort_wb_q_reg/NET0131 , \wishbone_TxAbort_wb_reg/NET0131 , \wishbone_TxBDAddress_reg[1]/NET0131 , \wishbone_TxBDAddress_reg[2]/NET0131 , \wishbone_TxBDAddress_reg[3]/NET0131 , \wishbone_TxBDAddress_reg[4]/NET0131 , \wishbone_TxBDAddress_reg[5]/NET0131 , \wishbone_TxBDAddress_reg[6]/NET0131 , \wishbone_TxBDAddress_reg[7]/NET0131 , \wishbone_TxBDRead_reg/NET0131 , \wishbone_TxBDReady_reg/NET0131 , \wishbone_TxB_IRQ_reg/NET0131 , \wishbone_TxByteCnt_reg[0]/NET0131 , \wishbone_TxByteCnt_reg[1]/NET0131 , \wishbone_TxDataLatched_reg[0]/NET0131 , \wishbone_TxDataLatched_reg[10]/NET0131 , \wishbone_TxDataLatched_reg[11]/NET0131 , \wishbone_TxDataLatched_reg[12]/NET0131 , \wishbone_TxDataLatched_reg[13]/NET0131 , \wishbone_TxDataLatched_reg[14]/NET0131 , \wishbone_TxDataLatched_reg[15]/NET0131 , \wishbone_TxDataLatched_reg[16]/NET0131 , \wishbone_TxDataLatched_reg[17]/NET0131 , \wishbone_TxDataLatched_reg[18]/NET0131 , \wishbone_TxDataLatched_reg[19]/NET0131 , \wishbone_TxDataLatched_reg[1]/NET0131 , \wishbone_TxDataLatched_reg[20]/NET0131 , \wishbone_TxDataLatched_reg[21]/NET0131 , \wishbone_TxDataLatched_reg[22]/NET0131 , \wishbone_TxDataLatched_reg[23]/NET0131 , \wishbone_TxDataLatched_reg[24]/NET0131 , \wishbone_TxDataLatched_reg[25]/NET0131 , \wishbone_TxDataLatched_reg[26]/NET0131 , \wishbone_TxDataLatched_reg[27]/NET0131 , \wishbone_TxDataLatched_reg[28]/NET0131 , \wishbone_TxDataLatched_reg[29]/NET0131 , \wishbone_TxDataLatched_reg[2]/NET0131 , \wishbone_TxDataLatched_reg[30]/NET0131 , \wishbone_TxDataLatched_reg[31]/NET0131 , \wishbone_TxDataLatched_reg[3]/NET0131 , \wishbone_TxDataLatched_reg[4]/NET0131 , \wishbone_TxDataLatched_reg[5]/NET0131 , \wishbone_TxDataLatched_reg[6]/NET0131 , \wishbone_TxDataLatched_reg[7]/NET0131 , \wishbone_TxDataLatched_reg[8]/NET0131 , \wishbone_TxDataLatched_reg[9]/NET0131 , \wishbone_TxData_reg[0]/NET0131 , \wishbone_TxData_reg[1]/NET0131 , \wishbone_TxData_reg[2]/NET0131 , \wishbone_TxData_reg[3]/NET0131 , \wishbone_TxData_reg[4]/NET0131 , \wishbone_TxData_reg[5]/NET0131 , \wishbone_TxData_reg[6]/NET0131 , \wishbone_TxData_reg[7]/NET0131 , \wishbone_TxDonePacketBlocked_reg/NET0131 , \wishbone_TxDonePacket_NotCleared_reg/NET0131 , \wishbone_TxDonePacket_reg/NET0131 , \wishbone_TxDone_wb_q_reg/NET0131 , \wishbone_TxDone_wb_reg/NET0131 , \wishbone_TxE_IRQ_reg/NET0131 , \wishbone_TxEn_needed_reg/NET0131 , \wishbone_TxEn_q_reg/NET0131 , \wishbone_TxEn_reg/NET0131 , \wishbone_TxEndFrm_reg/NET0131 , \wishbone_TxEndFrm_wb_reg/NET0131 , \wishbone_TxLength_reg[0]/NET0131 , \wishbone_TxLength_reg[10]/NET0131 , \wishbone_TxLength_reg[11]/NET0131 , \wishbone_TxLength_reg[12]/NET0131 , \wishbone_TxLength_reg[13]/NET0131 , \wishbone_TxLength_reg[14]/NET0131 , \wishbone_TxLength_reg[15]/NET0131 , \wishbone_TxLength_reg[1]/NET0131 , \wishbone_TxLength_reg[2]/NET0131 , \wishbone_TxLength_reg[3]/NET0131 , \wishbone_TxLength_reg[4]/NET0131 , \wishbone_TxLength_reg[5]/NET0131 , \wishbone_TxLength_reg[6]/NET0131 , \wishbone_TxLength_reg[7]/NET0131 , \wishbone_TxLength_reg[8]/NET0131 , \wishbone_TxLength_reg[9]/NET0131 , \wishbone_TxPointerLSB_reg[0]/NET0131 , \wishbone_TxPointerLSB_reg[1]/NET0131 , \wishbone_TxPointerLSB_rst_reg[0]/NET0131 , \wishbone_TxPointerLSB_rst_reg[1]/NET0131 , \wishbone_TxPointerMSB_reg[10]/NET0131 , \wishbone_TxPointerMSB_reg[11]/NET0131 , \wishbone_TxPointerMSB_reg[12]/NET0131 , \wishbone_TxPointerMSB_reg[13]/NET0131 , \wishbone_TxPointerMSB_reg[14]/NET0131 , \wishbone_TxPointerMSB_reg[15]/NET0131 , \wishbone_TxPointerMSB_reg[16]/NET0131 , \wishbone_TxPointerMSB_reg[17]/NET0131 , \wishbone_TxPointerMSB_reg[18]/NET0131 , \wishbone_TxPointerMSB_reg[19]/NET0131 , \wishbone_TxPointerMSB_reg[20]/NET0131 , \wishbone_TxPointerMSB_reg[21]/NET0131 , \wishbone_TxPointerMSB_reg[22]/NET0131 , \wishbone_TxPointerMSB_reg[23]/NET0131 , \wishbone_TxPointerMSB_reg[24]/NET0131 , \wishbone_TxPointerMSB_reg[25]/NET0131 , \wishbone_TxPointerMSB_reg[26]/NET0131 , \wishbone_TxPointerMSB_reg[27]/NET0131 , \wishbone_TxPointerMSB_reg[28]/NET0131 , \wishbone_TxPointerMSB_reg[29]/NET0131 , \wishbone_TxPointerMSB_reg[2]/NET0131 , \wishbone_TxPointerMSB_reg[30]/NET0131 , \wishbone_TxPointerMSB_reg[31]/NET0131 , \wishbone_TxPointerMSB_reg[3]/NET0131 , \wishbone_TxPointerMSB_reg[4]/NET0131 , \wishbone_TxPointerMSB_reg[5]/NET0131 , \wishbone_TxPointerMSB_reg[6]/NET0131 , \wishbone_TxPointerMSB_reg[7]/NET0131 , \wishbone_TxPointerMSB_reg[8]/NET0131 , \wishbone_TxPointerMSB_reg[9]/NET0131 , \wishbone_TxPointerRead_reg/NET0131 , \wishbone_TxRetryPacketBlocked_reg/NET0131 , \wishbone_TxRetryPacket_NotCleared_reg/NET0131 , \wishbone_TxRetryPacket_reg/NET0131 , \wishbone_TxRetry_q_reg/NET0131 , \wishbone_TxRetry_wb_q_reg/NET0131 , \wishbone_TxRetry_wb_reg/NET0131 , \wishbone_TxStartFrm_reg/NET0131 , \wishbone_TxStartFrm_sync2_reg/NET0131 , \wishbone_TxStartFrm_syncb2_reg/NET0131 , \wishbone_TxStartFrm_wb_reg/NET0131 , \wishbone_TxStatus_reg[11]/NET0131 , \wishbone_TxStatus_reg[12]/NET0131 , \wishbone_TxStatus_reg[13]/NET0131 , \wishbone_TxStatus_reg[14]/NET0131 , \wishbone_TxUnderRun_reg/NET0131 , \wishbone_TxUnderRun_sync1_reg/NET0131 , \wishbone_TxUnderRun_wb_reg/NET0131 , \wishbone_TxUsedData_q_reg/NET0131 , \wishbone_TxValidBytesLatched_reg[0]/NET0131 , \wishbone_TxValidBytesLatched_reg[1]/NET0131 , \wishbone_WB_ACK_O_reg/P0001 , \wishbone_WbEn_q_reg/NET0131 , \wishbone_WbEn_reg/NET0131 , \wishbone_WriteRxDataToFifoSync2_reg/NET0131 , \wishbone_WriteRxDataToFifoSync3_reg/NET0131 , \wishbone_WriteRxDataToFifo_reg/NET0131 , \wishbone_bd_ram_mem0_reg[0][0]/P0001 , \wishbone_bd_ram_mem0_reg[0][1]/P0001 , \wishbone_bd_ram_mem0_reg[0][2]/P0001 , \wishbone_bd_ram_mem0_reg[0][3]/P0001 , \wishbone_bd_ram_mem0_reg[0][4]/P0001 , \wishbone_bd_ram_mem0_reg[0][5]/P0001 , \wishbone_bd_ram_mem0_reg[0][6]/P0001 , \wishbone_bd_ram_mem0_reg[0][7]/P0001 , \wishbone_bd_ram_mem0_reg[100][0]/P0001 , \wishbone_bd_ram_mem0_reg[100][1]/P0001 , \wishbone_bd_ram_mem0_reg[100][2]/P0001 , \wishbone_bd_ram_mem0_reg[100][3]/P0001 , \wishbone_bd_ram_mem0_reg[100][4]/P0001 , \wishbone_bd_ram_mem0_reg[100][5]/P0001 , \wishbone_bd_ram_mem0_reg[100][6]/P0001 , \wishbone_bd_ram_mem0_reg[100][7]/P0001 , \wishbone_bd_ram_mem0_reg[101][0]/P0001 , \wishbone_bd_ram_mem0_reg[101][1]/P0001 , \wishbone_bd_ram_mem0_reg[101][2]/P0001 , \wishbone_bd_ram_mem0_reg[101][3]/P0001 , \wishbone_bd_ram_mem0_reg[101][4]/P0001 , \wishbone_bd_ram_mem0_reg[101][5]/P0001 , \wishbone_bd_ram_mem0_reg[101][6]/P0001 , \wishbone_bd_ram_mem0_reg[101][7]/P0001 , \wishbone_bd_ram_mem0_reg[102][0]/P0001 , \wishbone_bd_ram_mem0_reg[102][1]/P0001 , \wishbone_bd_ram_mem0_reg[102][2]/P0001 , \wishbone_bd_ram_mem0_reg[102][3]/P0001 , \wishbone_bd_ram_mem0_reg[102][4]/P0001 , \wishbone_bd_ram_mem0_reg[102][5]/P0001 , \wishbone_bd_ram_mem0_reg[102][6]/P0001 , \wishbone_bd_ram_mem0_reg[102][7]/P0001 , \wishbone_bd_ram_mem0_reg[103][0]/P0001 , \wishbone_bd_ram_mem0_reg[103][1]/P0001 , \wishbone_bd_ram_mem0_reg[103][2]/P0001 , \wishbone_bd_ram_mem0_reg[103][3]/P0001 , \wishbone_bd_ram_mem0_reg[103][4]/P0001 , \wishbone_bd_ram_mem0_reg[103][5]/P0001 , \wishbone_bd_ram_mem0_reg[103][6]/P0001 , \wishbone_bd_ram_mem0_reg[103][7]/P0001 , \wishbone_bd_ram_mem0_reg[104][0]/P0001 , \wishbone_bd_ram_mem0_reg[104][1]/P0001 , \wishbone_bd_ram_mem0_reg[104][2]/P0001 , \wishbone_bd_ram_mem0_reg[104][3]/P0001 , \wishbone_bd_ram_mem0_reg[104][4]/P0001 , \wishbone_bd_ram_mem0_reg[104][5]/P0001 , \wishbone_bd_ram_mem0_reg[104][6]/P0001 , \wishbone_bd_ram_mem0_reg[104][7]/P0001 , \wishbone_bd_ram_mem0_reg[105][0]/P0001 , \wishbone_bd_ram_mem0_reg[105][1]/P0001 , \wishbone_bd_ram_mem0_reg[105][2]/P0001 , \wishbone_bd_ram_mem0_reg[105][3]/P0001 , \wishbone_bd_ram_mem0_reg[105][4]/P0001 , \wishbone_bd_ram_mem0_reg[105][5]/P0001 , \wishbone_bd_ram_mem0_reg[105][6]/P0001 , \wishbone_bd_ram_mem0_reg[105][7]/P0001 , \wishbone_bd_ram_mem0_reg[106][0]/P0001 , \wishbone_bd_ram_mem0_reg[106][1]/P0001 , \wishbone_bd_ram_mem0_reg[106][2]/P0001 , \wishbone_bd_ram_mem0_reg[106][3]/P0001 , \wishbone_bd_ram_mem0_reg[106][4]/P0001 , \wishbone_bd_ram_mem0_reg[106][5]/P0001 , \wishbone_bd_ram_mem0_reg[106][6]/P0001 , \wishbone_bd_ram_mem0_reg[106][7]/P0001 , \wishbone_bd_ram_mem0_reg[107][0]/P0001 , \wishbone_bd_ram_mem0_reg[107][1]/P0001 , \wishbone_bd_ram_mem0_reg[107][2]/P0001 , \wishbone_bd_ram_mem0_reg[107][3]/P0001 , \wishbone_bd_ram_mem0_reg[107][4]/P0001 , \wishbone_bd_ram_mem0_reg[107][5]/P0001 , \wishbone_bd_ram_mem0_reg[107][6]/P0001 , \wishbone_bd_ram_mem0_reg[107][7]/P0001 , \wishbone_bd_ram_mem0_reg[108][0]/P0001 , \wishbone_bd_ram_mem0_reg[108][1]/P0001 , \wishbone_bd_ram_mem0_reg[108][2]/P0001 , \wishbone_bd_ram_mem0_reg[108][3]/P0001 , \wishbone_bd_ram_mem0_reg[108][4]/P0001 , \wishbone_bd_ram_mem0_reg[108][5]/P0001 , \wishbone_bd_ram_mem0_reg[108][6]/P0001 , \wishbone_bd_ram_mem0_reg[108][7]/P0001 , \wishbone_bd_ram_mem0_reg[109][0]/P0001 , \wishbone_bd_ram_mem0_reg[109][1]/P0001 , \wishbone_bd_ram_mem0_reg[109][2]/P0001 , \wishbone_bd_ram_mem0_reg[109][3]/P0001 , \wishbone_bd_ram_mem0_reg[109][4]/P0001 , \wishbone_bd_ram_mem0_reg[109][5]/P0001 , \wishbone_bd_ram_mem0_reg[109][6]/P0001 , \wishbone_bd_ram_mem0_reg[109][7]/P0001 , \wishbone_bd_ram_mem0_reg[10][0]/P0001 , \wishbone_bd_ram_mem0_reg[10][1]/P0001 , \wishbone_bd_ram_mem0_reg[10][2]/P0001 , \wishbone_bd_ram_mem0_reg[10][3]/P0001 , \wishbone_bd_ram_mem0_reg[10][4]/P0001 , \wishbone_bd_ram_mem0_reg[10][5]/P0001 , \wishbone_bd_ram_mem0_reg[10][6]/P0001 , \wishbone_bd_ram_mem0_reg[10][7]/P0001 , \wishbone_bd_ram_mem0_reg[110][0]/P0001 , \wishbone_bd_ram_mem0_reg[110][1]/P0001 , \wishbone_bd_ram_mem0_reg[110][2]/P0001 , \wishbone_bd_ram_mem0_reg[110][3]/P0001 , \wishbone_bd_ram_mem0_reg[110][4]/P0001 , \wishbone_bd_ram_mem0_reg[110][5]/P0001 , \wishbone_bd_ram_mem0_reg[110][6]/P0001 , \wishbone_bd_ram_mem0_reg[110][7]/P0001 , \wishbone_bd_ram_mem0_reg[111][0]/P0001 , \wishbone_bd_ram_mem0_reg[111][1]/P0001 , \wishbone_bd_ram_mem0_reg[111][2]/P0001 , \wishbone_bd_ram_mem0_reg[111][3]/P0001 , \wishbone_bd_ram_mem0_reg[111][4]/P0001 , \wishbone_bd_ram_mem0_reg[111][5]/P0001 , \wishbone_bd_ram_mem0_reg[111][6]/P0001 , \wishbone_bd_ram_mem0_reg[111][7]/P0001 , \wishbone_bd_ram_mem0_reg[112][0]/P0001 , \wishbone_bd_ram_mem0_reg[112][1]/P0001 , \wishbone_bd_ram_mem0_reg[112][2]/P0001 , \wishbone_bd_ram_mem0_reg[112][3]/P0001 , \wishbone_bd_ram_mem0_reg[112][4]/P0001 , \wishbone_bd_ram_mem0_reg[112][5]/P0001 , \wishbone_bd_ram_mem0_reg[112][6]/P0001 , \wishbone_bd_ram_mem0_reg[112][7]/P0001 , \wishbone_bd_ram_mem0_reg[113][0]/P0001 , \wishbone_bd_ram_mem0_reg[113][1]/P0001 , \wishbone_bd_ram_mem0_reg[113][2]/P0001 , \wishbone_bd_ram_mem0_reg[113][3]/P0001 , \wishbone_bd_ram_mem0_reg[113][4]/P0001 , \wishbone_bd_ram_mem0_reg[113][5]/P0001 , \wishbone_bd_ram_mem0_reg[113][6]/P0001 , \wishbone_bd_ram_mem0_reg[113][7]/P0001 , \wishbone_bd_ram_mem0_reg[114][0]/P0001 , \wishbone_bd_ram_mem0_reg[114][1]/P0001 , \wishbone_bd_ram_mem0_reg[114][2]/P0001 , \wishbone_bd_ram_mem0_reg[114][3]/P0001 , \wishbone_bd_ram_mem0_reg[114][4]/P0001 , \wishbone_bd_ram_mem0_reg[114][5]/P0001 , \wishbone_bd_ram_mem0_reg[114][6]/P0001 , \wishbone_bd_ram_mem0_reg[114][7]/P0001 , \wishbone_bd_ram_mem0_reg[115][0]/P0001 , \wishbone_bd_ram_mem0_reg[115][1]/P0001 , \wishbone_bd_ram_mem0_reg[115][2]/P0001 , \wishbone_bd_ram_mem0_reg[115][3]/P0001 , \wishbone_bd_ram_mem0_reg[115][4]/P0001 , \wishbone_bd_ram_mem0_reg[115][5]/P0001 , \wishbone_bd_ram_mem0_reg[115][6]/P0001 , \wishbone_bd_ram_mem0_reg[115][7]/P0001 , \wishbone_bd_ram_mem0_reg[116][0]/P0001 , \wishbone_bd_ram_mem0_reg[116][1]/P0001 , \wishbone_bd_ram_mem0_reg[116][2]/P0001 , \wishbone_bd_ram_mem0_reg[116][3]/P0001 , \wishbone_bd_ram_mem0_reg[116][4]/P0001 , \wishbone_bd_ram_mem0_reg[116][5]/P0001 , \wishbone_bd_ram_mem0_reg[116][6]/P0001 , \wishbone_bd_ram_mem0_reg[116][7]/P0001 , \wishbone_bd_ram_mem0_reg[117][0]/P0001 , \wishbone_bd_ram_mem0_reg[117][1]/P0001 , \wishbone_bd_ram_mem0_reg[117][2]/P0001 , \wishbone_bd_ram_mem0_reg[117][3]/P0001 , \wishbone_bd_ram_mem0_reg[117][4]/P0001 , \wishbone_bd_ram_mem0_reg[117][5]/P0001 , \wishbone_bd_ram_mem0_reg[117][6]/P0001 , \wishbone_bd_ram_mem0_reg[117][7]/P0001 , \wishbone_bd_ram_mem0_reg[118][0]/P0001 , \wishbone_bd_ram_mem0_reg[118][1]/P0001 , \wishbone_bd_ram_mem0_reg[118][2]/P0001 , \wishbone_bd_ram_mem0_reg[118][3]/P0001 , \wishbone_bd_ram_mem0_reg[118][4]/P0001 , \wishbone_bd_ram_mem0_reg[118][5]/P0001 , \wishbone_bd_ram_mem0_reg[118][6]/P0001 , \wishbone_bd_ram_mem0_reg[118][7]/P0001 , \wishbone_bd_ram_mem0_reg[119][0]/P0001 , \wishbone_bd_ram_mem0_reg[119][1]/P0001 , \wishbone_bd_ram_mem0_reg[119][2]/P0001 , \wishbone_bd_ram_mem0_reg[119][3]/P0001 , \wishbone_bd_ram_mem0_reg[119][4]/P0001 , \wishbone_bd_ram_mem0_reg[119][5]/P0001 , \wishbone_bd_ram_mem0_reg[119][6]/P0001 , \wishbone_bd_ram_mem0_reg[119][7]/P0001 , \wishbone_bd_ram_mem0_reg[11][0]/P0001 , \wishbone_bd_ram_mem0_reg[11][1]/P0001 , \wishbone_bd_ram_mem0_reg[11][2]/P0001 , \wishbone_bd_ram_mem0_reg[11][3]/P0001 , \wishbone_bd_ram_mem0_reg[11][4]/P0001 , \wishbone_bd_ram_mem0_reg[11][5]/P0001 , \wishbone_bd_ram_mem0_reg[11][6]/P0001 , \wishbone_bd_ram_mem0_reg[11][7]/P0001 , \wishbone_bd_ram_mem0_reg[120][0]/P0001 , \wishbone_bd_ram_mem0_reg[120][1]/P0001 , \wishbone_bd_ram_mem0_reg[120][2]/P0001 , \wishbone_bd_ram_mem0_reg[120][3]/P0001 , \wishbone_bd_ram_mem0_reg[120][4]/P0001 , \wishbone_bd_ram_mem0_reg[120][5]/P0001 , \wishbone_bd_ram_mem0_reg[120][6]/P0001 , \wishbone_bd_ram_mem0_reg[120][7]/P0001 , \wishbone_bd_ram_mem0_reg[121][0]/P0001 , \wishbone_bd_ram_mem0_reg[121][1]/P0001 , \wishbone_bd_ram_mem0_reg[121][2]/P0001 , \wishbone_bd_ram_mem0_reg[121][3]/P0001 , \wishbone_bd_ram_mem0_reg[121][4]/P0001 , \wishbone_bd_ram_mem0_reg[121][5]/P0001 , \wishbone_bd_ram_mem0_reg[121][6]/P0001 , \wishbone_bd_ram_mem0_reg[121][7]/P0001 , \wishbone_bd_ram_mem0_reg[122][0]/P0001 , \wishbone_bd_ram_mem0_reg[122][1]/P0001 , \wishbone_bd_ram_mem0_reg[122][2]/P0001 , \wishbone_bd_ram_mem0_reg[122][3]/P0001 , \wishbone_bd_ram_mem0_reg[122][4]/P0001 , \wishbone_bd_ram_mem0_reg[122][5]/P0001 , \wishbone_bd_ram_mem0_reg[122][6]/P0001 , \wishbone_bd_ram_mem0_reg[122][7]/P0001 , \wishbone_bd_ram_mem0_reg[123][0]/P0001 , \wishbone_bd_ram_mem0_reg[123][1]/P0001 , \wishbone_bd_ram_mem0_reg[123][2]/P0001 , \wishbone_bd_ram_mem0_reg[123][3]/P0001 , \wishbone_bd_ram_mem0_reg[123][4]/P0001 , \wishbone_bd_ram_mem0_reg[123][5]/P0001 , \wishbone_bd_ram_mem0_reg[123][6]/P0001 , \wishbone_bd_ram_mem0_reg[123][7]/P0001 , \wishbone_bd_ram_mem0_reg[124][0]/P0001 , \wishbone_bd_ram_mem0_reg[124][1]/P0001 , \wishbone_bd_ram_mem0_reg[124][2]/P0001 , \wishbone_bd_ram_mem0_reg[124][3]/P0001 , \wishbone_bd_ram_mem0_reg[124][4]/P0001 , \wishbone_bd_ram_mem0_reg[124][5]/P0001 , \wishbone_bd_ram_mem0_reg[124][6]/P0001 , \wishbone_bd_ram_mem0_reg[124][7]/P0001 , \wishbone_bd_ram_mem0_reg[125][0]/P0001 , \wishbone_bd_ram_mem0_reg[125][1]/P0001 , \wishbone_bd_ram_mem0_reg[125][2]/P0001 , \wishbone_bd_ram_mem0_reg[125][3]/P0001 , \wishbone_bd_ram_mem0_reg[125][4]/P0001 , \wishbone_bd_ram_mem0_reg[125][5]/P0001 , \wishbone_bd_ram_mem0_reg[125][6]/P0001 , \wishbone_bd_ram_mem0_reg[125][7]/P0001 , \wishbone_bd_ram_mem0_reg[126][0]/P0001 , \wishbone_bd_ram_mem0_reg[126][1]/P0001 , \wishbone_bd_ram_mem0_reg[126][2]/P0001 , \wishbone_bd_ram_mem0_reg[126][3]/P0001 , \wishbone_bd_ram_mem0_reg[126][4]/P0001 , \wishbone_bd_ram_mem0_reg[126][5]/P0001 , \wishbone_bd_ram_mem0_reg[126][6]/P0001 , \wishbone_bd_ram_mem0_reg[126][7]/P0001 , \wishbone_bd_ram_mem0_reg[127][0]/P0001 , \wishbone_bd_ram_mem0_reg[127][1]/P0001 , \wishbone_bd_ram_mem0_reg[127][2]/P0001 , \wishbone_bd_ram_mem0_reg[127][3]/P0001 , \wishbone_bd_ram_mem0_reg[127][4]/P0001 , \wishbone_bd_ram_mem0_reg[127][5]/P0001 , \wishbone_bd_ram_mem0_reg[127][6]/P0001 , \wishbone_bd_ram_mem0_reg[127][7]/P0001 , \wishbone_bd_ram_mem0_reg[128][0]/P0001 , \wishbone_bd_ram_mem0_reg[128][1]/P0001 , \wishbone_bd_ram_mem0_reg[128][2]/P0001 , \wishbone_bd_ram_mem0_reg[128][3]/P0001 , \wishbone_bd_ram_mem0_reg[128][4]/P0001 , \wishbone_bd_ram_mem0_reg[128][5]/P0001 , \wishbone_bd_ram_mem0_reg[128][6]/P0001 , \wishbone_bd_ram_mem0_reg[128][7]/P0001 , \wishbone_bd_ram_mem0_reg[129][0]/P0001 , \wishbone_bd_ram_mem0_reg[129][1]/P0001 , \wishbone_bd_ram_mem0_reg[129][2]/P0001 , \wishbone_bd_ram_mem0_reg[129][3]/P0001 , \wishbone_bd_ram_mem0_reg[129][4]/P0001 , \wishbone_bd_ram_mem0_reg[129][5]/P0001 , \wishbone_bd_ram_mem0_reg[129][6]/P0001 , \wishbone_bd_ram_mem0_reg[129][7]/P0001 , \wishbone_bd_ram_mem0_reg[12][0]/P0001 , \wishbone_bd_ram_mem0_reg[12][1]/P0001 , \wishbone_bd_ram_mem0_reg[12][2]/P0001 , \wishbone_bd_ram_mem0_reg[12][3]/P0001 , \wishbone_bd_ram_mem0_reg[12][4]/P0001 , \wishbone_bd_ram_mem0_reg[12][5]/P0001 , \wishbone_bd_ram_mem0_reg[12][6]/P0001 , \wishbone_bd_ram_mem0_reg[12][7]/P0001 , \wishbone_bd_ram_mem0_reg[130][0]/P0001 , \wishbone_bd_ram_mem0_reg[130][1]/P0001 , \wishbone_bd_ram_mem0_reg[130][2]/P0001 , \wishbone_bd_ram_mem0_reg[130][3]/P0001 , \wishbone_bd_ram_mem0_reg[130][4]/P0001 , \wishbone_bd_ram_mem0_reg[130][5]/P0001 , \wishbone_bd_ram_mem0_reg[130][6]/P0001 , \wishbone_bd_ram_mem0_reg[130][7]/P0001 , \wishbone_bd_ram_mem0_reg[131][0]/P0001 , \wishbone_bd_ram_mem0_reg[131][1]/P0001 , \wishbone_bd_ram_mem0_reg[131][2]/P0001 , \wishbone_bd_ram_mem0_reg[131][3]/P0001 , \wishbone_bd_ram_mem0_reg[131][4]/P0001 , \wishbone_bd_ram_mem0_reg[131][5]/P0001 , \wishbone_bd_ram_mem0_reg[131][6]/P0001 , \wishbone_bd_ram_mem0_reg[131][7]/P0001 , \wishbone_bd_ram_mem0_reg[132][0]/P0001 , \wishbone_bd_ram_mem0_reg[132][1]/P0001 , \wishbone_bd_ram_mem0_reg[132][2]/P0001 , \wishbone_bd_ram_mem0_reg[132][3]/P0001 , \wishbone_bd_ram_mem0_reg[132][4]/P0001 , \wishbone_bd_ram_mem0_reg[132][5]/P0001 , \wishbone_bd_ram_mem0_reg[132][6]/P0001 , \wishbone_bd_ram_mem0_reg[132][7]/P0001 , \wishbone_bd_ram_mem0_reg[133][0]/P0001 , \wishbone_bd_ram_mem0_reg[133][1]/P0001 , \wishbone_bd_ram_mem0_reg[133][2]/P0001 , \wishbone_bd_ram_mem0_reg[133][3]/P0001 , \wishbone_bd_ram_mem0_reg[133][4]/P0001 , \wishbone_bd_ram_mem0_reg[133][5]/P0001 , \wishbone_bd_ram_mem0_reg[133][6]/P0001 , \wishbone_bd_ram_mem0_reg[133][7]/P0001 , \wishbone_bd_ram_mem0_reg[134][0]/P0001 , \wishbone_bd_ram_mem0_reg[134][1]/P0001 , \wishbone_bd_ram_mem0_reg[134][2]/P0001 , \wishbone_bd_ram_mem0_reg[134][3]/P0001 , \wishbone_bd_ram_mem0_reg[134][4]/P0001 , \wishbone_bd_ram_mem0_reg[134][5]/P0001 , \wishbone_bd_ram_mem0_reg[134][6]/P0001 , \wishbone_bd_ram_mem0_reg[134][7]/P0001 , \wishbone_bd_ram_mem0_reg[135][0]/P0001 , \wishbone_bd_ram_mem0_reg[135][1]/P0001 , \wishbone_bd_ram_mem0_reg[135][2]/P0001 , \wishbone_bd_ram_mem0_reg[135][3]/P0001 , \wishbone_bd_ram_mem0_reg[135][4]/P0001 , \wishbone_bd_ram_mem0_reg[135][5]/P0001 , \wishbone_bd_ram_mem0_reg[135][6]/P0001 , \wishbone_bd_ram_mem0_reg[135][7]/P0001 , \wishbone_bd_ram_mem0_reg[136][0]/P0001 , \wishbone_bd_ram_mem0_reg[136][1]/P0001 , \wishbone_bd_ram_mem0_reg[136][2]/P0001 , \wishbone_bd_ram_mem0_reg[136][3]/P0001 , \wishbone_bd_ram_mem0_reg[136][4]/P0001 , \wishbone_bd_ram_mem0_reg[136][5]/P0001 , \wishbone_bd_ram_mem0_reg[136][6]/P0001 , \wishbone_bd_ram_mem0_reg[136][7]/P0001 , \wishbone_bd_ram_mem0_reg[137][0]/P0001 , \wishbone_bd_ram_mem0_reg[137][1]/P0001 , \wishbone_bd_ram_mem0_reg[137][2]/P0001 , \wishbone_bd_ram_mem0_reg[137][3]/P0001 , \wishbone_bd_ram_mem0_reg[137][4]/P0001 , \wishbone_bd_ram_mem0_reg[137][5]/P0001 , \wishbone_bd_ram_mem0_reg[137][6]/P0001 , \wishbone_bd_ram_mem0_reg[137][7]/P0001 , \wishbone_bd_ram_mem0_reg[138][0]/P0001 , \wishbone_bd_ram_mem0_reg[138][1]/P0001 , \wishbone_bd_ram_mem0_reg[138][2]/P0001 , \wishbone_bd_ram_mem0_reg[138][3]/P0001 , \wishbone_bd_ram_mem0_reg[138][4]/P0001 , \wishbone_bd_ram_mem0_reg[138][5]/P0001 , \wishbone_bd_ram_mem0_reg[138][6]/P0001 , \wishbone_bd_ram_mem0_reg[138][7]/P0001 , \wishbone_bd_ram_mem0_reg[139][0]/P0001 , \wishbone_bd_ram_mem0_reg[139][1]/P0001 , \wishbone_bd_ram_mem0_reg[139][2]/P0001 , \wishbone_bd_ram_mem0_reg[139][3]/P0001 , \wishbone_bd_ram_mem0_reg[139][4]/P0001 , \wishbone_bd_ram_mem0_reg[139][5]/P0001 , \wishbone_bd_ram_mem0_reg[139][6]/P0001 , \wishbone_bd_ram_mem0_reg[139][7]/P0001 , \wishbone_bd_ram_mem0_reg[13][0]/P0001 , \wishbone_bd_ram_mem0_reg[13][1]/P0001 , \wishbone_bd_ram_mem0_reg[13][2]/P0001 , \wishbone_bd_ram_mem0_reg[13][3]/P0001 , \wishbone_bd_ram_mem0_reg[13][4]/P0001 , \wishbone_bd_ram_mem0_reg[13][5]/P0001 , \wishbone_bd_ram_mem0_reg[13][6]/P0001 , \wishbone_bd_ram_mem0_reg[13][7]/P0001 , \wishbone_bd_ram_mem0_reg[140][0]/P0001 , \wishbone_bd_ram_mem0_reg[140][1]/P0001 , \wishbone_bd_ram_mem0_reg[140][2]/P0001 , \wishbone_bd_ram_mem0_reg[140][3]/P0001 , \wishbone_bd_ram_mem0_reg[140][4]/P0001 , \wishbone_bd_ram_mem0_reg[140][5]/P0001 , \wishbone_bd_ram_mem0_reg[140][6]/P0001 , \wishbone_bd_ram_mem0_reg[140][7]/P0001 , \wishbone_bd_ram_mem0_reg[141][0]/P0001 , \wishbone_bd_ram_mem0_reg[141][1]/P0001 , \wishbone_bd_ram_mem0_reg[141][2]/P0001 , \wishbone_bd_ram_mem0_reg[141][3]/P0001 , \wishbone_bd_ram_mem0_reg[141][4]/P0001 , \wishbone_bd_ram_mem0_reg[141][5]/P0001 , \wishbone_bd_ram_mem0_reg[141][6]/P0001 , \wishbone_bd_ram_mem0_reg[141][7]/P0001 , \wishbone_bd_ram_mem0_reg[142][0]/P0001 , \wishbone_bd_ram_mem0_reg[142][1]/P0001 , \wishbone_bd_ram_mem0_reg[142][2]/P0001 , \wishbone_bd_ram_mem0_reg[142][3]/P0001 , \wishbone_bd_ram_mem0_reg[142][4]/P0001 , \wishbone_bd_ram_mem0_reg[142][5]/P0001 , \wishbone_bd_ram_mem0_reg[142][6]/P0001 , \wishbone_bd_ram_mem0_reg[142][7]/P0001 , \wishbone_bd_ram_mem0_reg[143][0]/P0001 , \wishbone_bd_ram_mem0_reg[143][1]/P0001 , \wishbone_bd_ram_mem0_reg[143][2]/P0001 , \wishbone_bd_ram_mem0_reg[143][3]/P0001 , \wishbone_bd_ram_mem0_reg[143][4]/P0001 , \wishbone_bd_ram_mem0_reg[143][5]/P0001 , \wishbone_bd_ram_mem0_reg[143][6]/P0001 , \wishbone_bd_ram_mem0_reg[143][7]/P0001 , \wishbone_bd_ram_mem0_reg[144][0]/P0001 , \wishbone_bd_ram_mem0_reg[144][1]/P0001 , \wishbone_bd_ram_mem0_reg[144][2]/P0001 , \wishbone_bd_ram_mem0_reg[144][3]/P0001 , \wishbone_bd_ram_mem0_reg[144][4]/P0001 , \wishbone_bd_ram_mem0_reg[144][5]/P0001 , \wishbone_bd_ram_mem0_reg[144][6]/P0001 , \wishbone_bd_ram_mem0_reg[144][7]/P0001 , \wishbone_bd_ram_mem0_reg[145][0]/P0001 , \wishbone_bd_ram_mem0_reg[145][1]/P0001 , \wishbone_bd_ram_mem0_reg[145][2]/P0001 , \wishbone_bd_ram_mem0_reg[145][3]/P0001 , \wishbone_bd_ram_mem0_reg[145][4]/P0001 , \wishbone_bd_ram_mem0_reg[145][5]/P0001 , \wishbone_bd_ram_mem0_reg[145][6]/P0001 , \wishbone_bd_ram_mem0_reg[145][7]/P0001 , \wishbone_bd_ram_mem0_reg[146][0]/P0001 , \wishbone_bd_ram_mem0_reg[146][1]/P0001 , \wishbone_bd_ram_mem0_reg[146][2]/P0001 , \wishbone_bd_ram_mem0_reg[146][3]/P0001 , \wishbone_bd_ram_mem0_reg[146][4]/P0001 , \wishbone_bd_ram_mem0_reg[146][5]/P0001 , \wishbone_bd_ram_mem0_reg[146][6]/P0001 , \wishbone_bd_ram_mem0_reg[146][7]/P0001 , \wishbone_bd_ram_mem0_reg[147][0]/P0001 , \wishbone_bd_ram_mem0_reg[147][1]/P0001 , \wishbone_bd_ram_mem0_reg[147][2]/P0001 , \wishbone_bd_ram_mem0_reg[147][3]/P0001 , \wishbone_bd_ram_mem0_reg[147][4]/P0001 , \wishbone_bd_ram_mem0_reg[147][5]/P0001 , \wishbone_bd_ram_mem0_reg[147][6]/P0001 , \wishbone_bd_ram_mem0_reg[147][7]/P0001 , \wishbone_bd_ram_mem0_reg[148][0]/P0001 , \wishbone_bd_ram_mem0_reg[148][1]/P0001 , \wishbone_bd_ram_mem0_reg[148][2]/P0001 , \wishbone_bd_ram_mem0_reg[148][3]/P0001 , \wishbone_bd_ram_mem0_reg[148][4]/P0001 , \wishbone_bd_ram_mem0_reg[148][5]/P0001 , \wishbone_bd_ram_mem0_reg[148][6]/P0001 , \wishbone_bd_ram_mem0_reg[148][7]/P0001 , \wishbone_bd_ram_mem0_reg[149][0]/P0001 , \wishbone_bd_ram_mem0_reg[149][1]/P0001 , \wishbone_bd_ram_mem0_reg[149][2]/P0001 , \wishbone_bd_ram_mem0_reg[149][3]/P0001 , \wishbone_bd_ram_mem0_reg[149][4]/P0001 , \wishbone_bd_ram_mem0_reg[149][5]/P0001 , \wishbone_bd_ram_mem0_reg[149][6]/P0001 , \wishbone_bd_ram_mem0_reg[149][7]/P0001 , \wishbone_bd_ram_mem0_reg[14][0]/P0001 , \wishbone_bd_ram_mem0_reg[14][1]/P0001 , \wishbone_bd_ram_mem0_reg[14][2]/P0001 , \wishbone_bd_ram_mem0_reg[14][3]/P0001 , \wishbone_bd_ram_mem0_reg[14][4]/P0001 , \wishbone_bd_ram_mem0_reg[14][5]/P0001 , \wishbone_bd_ram_mem0_reg[14][6]/P0001 , \wishbone_bd_ram_mem0_reg[14][7]/P0001 , \wishbone_bd_ram_mem0_reg[150][0]/P0001 , \wishbone_bd_ram_mem0_reg[150][1]/P0001 , \wishbone_bd_ram_mem0_reg[150][2]/P0001 , \wishbone_bd_ram_mem0_reg[150][3]/P0001 , \wishbone_bd_ram_mem0_reg[150][4]/P0001 , \wishbone_bd_ram_mem0_reg[150][5]/P0001 , \wishbone_bd_ram_mem0_reg[150][6]/P0001 , \wishbone_bd_ram_mem0_reg[150][7]/P0001 , \wishbone_bd_ram_mem0_reg[151][0]/P0001 , \wishbone_bd_ram_mem0_reg[151][1]/P0001 , \wishbone_bd_ram_mem0_reg[151][2]/P0001 , \wishbone_bd_ram_mem0_reg[151][3]/P0001 , \wishbone_bd_ram_mem0_reg[151][4]/P0001 , \wishbone_bd_ram_mem0_reg[151][5]/P0001 , \wishbone_bd_ram_mem0_reg[151][6]/P0001 , \wishbone_bd_ram_mem0_reg[151][7]/P0001 , \wishbone_bd_ram_mem0_reg[152][0]/P0001 , \wishbone_bd_ram_mem0_reg[152][1]/P0001 , \wishbone_bd_ram_mem0_reg[152][2]/P0001 , \wishbone_bd_ram_mem0_reg[152][3]/P0001 , \wishbone_bd_ram_mem0_reg[152][4]/P0001 , \wishbone_bd_ram_mem0_reg[152][5]/P0001 , \wishbone_bd_ram_mem0_reg[152][6]/P0001 , \wishbone_bd_ram_mem0_reg[152][7]/P0001 , \wishbone_bd_ram_mem0_reg[153][0]/P0001 , \wishbone_bd_ram_mem0_reg[153][1]/P0001 , \wishbone_bd_ram_mem0_reg[153][2]/P0001 , \wishbone_bd_ram_mem0_reg[153][3]/P0001 , \wishbone_bd_ram_mem0_reg[153][4]/P0001 , \wishbone_bd_ram_mem0_reg[153][5]/P0001 , \wishbone_bd_ram_mem0_reg[153][6]/P0001 , \wishbone_bd_ram_mem0_reg[153][7]/P0001 , \wishbone_bd_ram_mem0_reg[154][0]/P0001 , \wishbone_bd_ram_mem0_reg[154][1]/P0001 , \wishbone_bd_ram_mem0_reg[154][2]/P0001 , \wishbone_bd_ram_mem0_reg[154][3]/P0001 , \wishbone_bd_ram_mem0_reg[154][4]/P0001 , \wishbone_bd_ram_mem0_reg[154][5]/P0001 , \wishbone_bd_ram_mem0_reg[154][6]/P0001 , \wishbone_bd_ram_mem0_reg[154][7]/P0001 , \wishbone_bd_ram_mem0_reg[155][0]/P0001 , \wishbone_bd_ram_mem0_reg[155][1]/P0001 , \wishbone_bd_ram_mem0_reg[155][2]/P0001 , \wishbone_bd_ram_mem0_reg[155][3]/P0001 , \wishbone_bd_ram_mem0_reg[155][4]/P0001 , \wishbone_bd_ram_mem0_reg[155][5]/P0001 , \wishbone_bd_ram_mem0_reg[155][6]/P0001 , \wishbone_bd_ram_mem0_reg[155][7]/P0001 , \wishbone_bd_ram_mem0_reg[156][0]/P0001 , \wishbone_bd_ram_mem0_reg[156][1]/P0001 , \wishbone_bd_ram_mem0_reg[156][2]/P0001 , \wishbone_bd_ram_mem0_reg[156][3]/P0001 , \wishbone_bd_ram_mem0_reg[156][4]/P0001 , \wishbone_bd_ram_mem0_reg[156][5]/P0001 , \wishbone_bd_ram_mem0_reg[156][6]/P0001 , \wishbone_bd_ram_mem0_reg[156][7]/P0001 , \wishbone_bd_ram_mem0_reg[157][0]/P0001 , \wishbone_bd_ram_mem0_reg[157][1]/P0001 , \wishbone_bd_ram_mem0_reg[157][2]/P0001 , \wishbone_bd_ram_mem0_reg[157][3]/P0001 , \wishbone_bd_ram_mem0_reg[157][4]/P0001 , \wishbone_bd_ram_mem0_reg[157][5]/P0001 , \wishbone_bd_ram_mem0_reg[157][6]/P0001 , \wishbone_bd_ram_mem0_reg[157][7]/P0001 , \wishbone_bd_ram_mem0_reg[158][0]/P0001 , \wishbone_bd_ram_mem0_reg[158][1]/P0001 , \wishbone_bd_ram_mem0_reg[158][2]/P0001 , \wishbone_bd_ram_mem0_reg[158][3]/P0001 , \wishbone_bd_ram_mem0_reg[158][4]/P0001 , \wishbone_bd_ram_mem0_reg[158][5]/P0001 , \wishbone_bd_ram_mem0_reg[158][6]/P0001 , \wishbone_bd_ram_mem0_reg[158][7]/P0001 , \wishbone_bd_ram_mem0_reg[159][0]/P0001 , \wishbone_bd_ram_mem0_reg[159][1]/P0001 , \wishbone_bd_ram_mem0_reg[159][2]/P0001 , \wishbone_bd_ram_mem0_reg[159][3]/P0001 , \wishbone_bd_ram_mem0_reg[159][4]/P0001 , \wishbone_bd_ram_mem0_reg[159][5]/P0001 , \wishbone_bd_ram_mem0_reg[159][6]/P0001 , \wishbone_bd_ram_mem0_reg[159][7]/P0001 , \wishbone_bd_ram_mem0_reg[15][0]/P0001 , \wishbone_bd_ram_mem0_reg[15][1]/P0001 , \wishbone_bd_ram_mem0_reg[15][2]/P0001 , \wishbone_bd_ram_mem0_reg[15][3]/P0001 , \wishbone_bd_ram_mem0_reg[15][4]/P0001 , \wishbone_bd_ram_mem0_reg[15][5]/P0001 , \wishbone_bd_ram_mem0_reg[15][6]/P0001 , \wishbone_bd_ram_mem0_reg[15][7]/P0001 , \wishbone_bd_ram_mem0_reg[160][0]/P0001 , \wishbone_bd_ram_mem0_reg[160][1]/P0001 , \wishbone_bd_ram_mem0_reg[160][2]/P0001 , \wishbone_bd_ram_mem0_reg[160][3]/P0001 , \wishbone_bd_ram_mem0_reg[160][4]/P0001 , \wishbone_bd_ram_mem0_reg[160][5]/P0001 , \wishbone_bd_ram_mem0_reg[160][6]/P0001 , \wishbone_bd_ram_mem0_reg[160][7]/P0001 , \wishbone_bd_ram_mem0_reg[161][0]/P0001 , \wishbone_bd_ram_mem0_reg[161][1]/P0001 , \wishbone_bd_ram_mem0_reg[161][2]/P0001 , \wishbone_bd_ram_mem0_reg[161][3]/P0001 , \wishbone_bd_ram_mem0_reg[161][4]/P0001 , \wishbone_bd_ram_mem0_reg[161][5]/P0001 , \wishbone_bd_ram_mem0_reg[161][6]/P0001 , \wishbone_bd_ram_mem0_reg[161][7]/P0001 , \wishbone_bd_ram_mem0_reg[162][0]/P0001 , \wishbone_bd_ram_mem0_reg[162][1]/P0001 , \wishbone_bd_ram_mem0_reg[162][2]/P0001 , \wishbone_bd_ram_mem0_reg[162][3]/P0001 , \wishbone_bd_ram_mem0_reg[162][4]/P0001 , \wishbone_bd_ram_mem0_reg[162][5]/P0001 , \wishbone_bd_ram_mem0_reg[162][6]/P0001 , \wishbone_bd_ram_mem0_reg[162][7]/P0001 , \wishbone_bd_ram_mem0_reg[163][0]/P0001 , \wishbone_bd_ram_mem0_reg[163][1]/P0001 , \wishbone_bd_ram_mem0_reg[163][2]/P0001 , \wishbone_bd_ram_mem0_reg[163][3]/P0001 , \wishbone_bd_ram_mem0_reg[163][4]/P0001 , \wishbone_bd_ram_mem0_reg[163][5]/P0001 , \wishbone_bd_ram_mem0_reg[163][6]/P0001 , \wishbone_bd_ram_mem0_reg[163][7]/P0001 , \wishbone_bd_ram_mem0_reg[164][0]/P0001 , \wishbone_bd_ram_mem0_reg[164][1]/P0001 , \wishbone_bd_ram_mem0_reg[164][2]/P0001 , \wishbone_bd_ram_mem0_reg[164][3]/P0001 , \wishbone_bd_ram_mem0_reg[164][4]/P0001 , \wishbone_bd_ram_mem0_reg[164][5]/P0001 , \wishbone_bd_ram_mem0_reg[164][6]/P0001 , \wishbone_bd_ram_mem0_reg[164][7]/P0001 , \wishbone_bd_ram_mem0_reg[165][0]/P0001 , \wishbone_bd_ram_mem0_reg[165][1]/P0001 , \wishbone_bd_ram_mem0_reg[165][2]/P0001 , \wishbone_bd_ram_mem0_reg[165][3]/P0001 , \wishbone_bd_ram_mem0_reg[165][4]/P0001 , \wishbone_bd_ram_mem0_reg[165][5]/P0001 , \wishbone_bd_ram_mem0_reg[165][6]/P0001 , \wishbone_bd_ram_mem0_reg[165][7]/P0001 , \wishbone_bd_ram_mem0_reg[166][0]/P0001 , \wishbone_bd_ram_mem0_reg[166][1]/P0001 , \wishbone_bd_ram_mem0_reg[166][2]/P0001 , \wishbone_bd_ram_mem0_reg[166][3]/P0001 , \wishbone_bd_ram_mem0_reg[166][4]/P0001 , \wishbone_bd_ram_mem0_reg[166][5]/P0001 , \wishbone_bd_ram_mem0_reg[166][6]/P0001 , \wishbone_bd_ram_mem0_reg[166][7]/P0001 , \wishbone_bd_ram_mem0_reg[167][0]/P0001 , \wishbone_bd_ram_mem0_reg[167][1]/P0001 , \wishbone_bd_ram_mem0_reg[167][2]/P0001 , \wishbone_bd_ram_mem0_reg[167][3]/P0001 , \wishbone_bd_ram_mem0_reg[167][4]/P0001 , \wishbone_bd_ram_mem0_reg[167][5]/P0001 , \wishbone_bd_ram_mem0_reg[167][6]/P0001 , \wishbone_bd_ram_mem0_reg[167][7]/P0001 , \wishbone_bd_ram_mem0_reg[168][0]/P0001 , \wishbone_bd_ram_mem0_reg[168][1]/P0001 , \wishbone_bd_ram_mem0_reg[168][2]/P0001 , \wishbone_bd_ram_mem0_reg[168][3]/P0001 , \wishbone_bd_ram_mem0_reg[168][4]/P0001 , \wishbone_bd_ram_mem0_reg[168][5]/P0001 , \wishbone_bd_ram_mem0_reg[168][6]/P0001 , \wishbone_bd_ram_mem0_reg[168][7]/P0001 , \wishbone_bd_ram_mem0_reg[169][0]/P0001 , \wishbone_bd_ram_mem0_reg[169][1]/P0001 , \wishbone_bd_ram_mem0_reg[169][2]/P0001 , \wishbone_bd_ram_mem0_reg[169][3]/P0001 , \wishbone_bd_ram_mem0_reg[169][4]/P0001 , \wishbone_bd_ram_mem0_reg[169][5]/P0001 , \wishbone_bd_ram_mem0_reg[169][6]/P0001 , \wishbone_bd_ram_mem0_reg[169][7]/P0001 , \wishbone_bd_ram_mem0_reg[16][0]/P0001 , \wishbone_bd_ram_mem0_reg[16][1]/P0001 , \wishbone_bd_ram_mem0_reg[16][2]/P0001 , \wishbone_bd_ram_mem0_reg[16][3]/P0001 , \wishbone_bd_ram_mem0_reg[16][4]/P0001 , \wishbone_bd_ram_mem0_reg[16][5]/P0001 , \wishbone_bd_ram_mem0_reg[16][6]/P0001 , \wishbone_bd_ram_mem0_reg[16][7]/P0001 , \wishbone_bd_ram_mem0_reg[170][0]/P0001 , \wishbone_bd_ram_mem0_reg[170][1]/P0001 , \wishbone_bd_ram_mem0_reg[170][2]/P0001 , \wishbone_bd_ram_mem0_reg[170][3]/P0001 , \wishbone_bd_ram_mem0_reg[170][4]/P0001 , \wishbone_bd_ram_mem0_reg[170][5]/P0001 , \wishbone_bd_ram_mem0_reg[170][6]/P0001 , \wishbone_bd_ram_mem0_reg[170][7]/P0001 , \wishbone_bd_ram_mem0_reg[171][0]/P0001 , \wishbone_bd_ram_mem0_reg[171][1]/P0001 , \wishbone_bd_ram_mem0_reg[171][2]/P0001 , \wishbone_bd_ram_mem0_reg[171][3]/P0001 , \wishbone_bd_ram_mem0_reg[171][4]/P0001 , \wishbone_bd_ram_mem0_reg[171][5]/P0001 , \wishbone_bd_ram_mem0_reg[171][6]/P0001 , \wishbone_bd_ram_mem0_reg[171][7]/P0001 , \wishbone_bd_ram_mem0_reg[172][0]/P0001 , \wishbone_bd_ram_mem0_reg[172][1]/P0001 , \wishbone_bd_ram_mem0_reg[172][2]/P0001 , \wishbone_bd_ram_mem0_reg[172][3]/P0001 , \wishbone_bd_ram_mem0_reg[172][4]/P0001 , \wishbone_bd_ram_mem0_reg[172][5]/P0001 , \wishbone_bd_ram_mem0_reg[172][6]/P0001 , \wishbone_bd_ram_mem0_reg[172][7]/P0001 , \wishbone_bd_ram_mem0_reg[173][0]/P0001 , \wishbone_bd_ram_mem0_reg[173][1]/P0001 , \wishbone_bd_ram_mem0_reg[173][2]/P0001 , \wishbone_bd_ram_mem0_reg[173][3]/P0001 , \wishbone_bd_ram_mem0_reg[173][4]/P0001 , \wishbone_bd_ram_mem0_reg[173][5]/P0001 , \wishbone_bd_ram_mem0_reg[173][6]/P0001 , \wishbone_bd_ram_mem0_reg[173][7]/P0001 , \wishbone_bd_ram_mem0_reg[174][0]/P0001 , \wishbone_bd_ram_mem0_reg[174][1]/P0001 , \wishbone_bd_ram_mem0_reg[174][2]/P0001 , \wishbone_bd_ram_mem0_reg[174][3]/P0001 , \wishbone_bd_ram_mem0_reg[174][4]/P0001 , \wishbone_bd_ram_mem0_reg[174][5]/P0001 , \wishbone_bd_ram_mem0_reg[174][6]/P0001 , \wishbone_bd_ram_mem0_reg[174][7]/P0001 , \wishbone_bd_ram_mem0_reg[175][0]/P0001 , \wishbone_bd_ram_mem0_reg[175][1]/P0001 , \wishbone_bd_ram_mem0_reg[175][2]/P0001 , \wishbone_bd_ram_mem0_reg[175][3]/P0001 , \wishbone_bd_ram_mem0_reg[175][4]/P0001 , \wishbone_bd_ram_mem0_reg[175][5]/P0001 , \wishbone_bd_ram_mem0_reg[175][6]/P0001 , \wishbone_bd_ram_mem0_reg[175][7]/P0001 , \wishbone_bd_ram_mem0_reg[176][0]/P0001 , \wishbone_bd_ram_mem0_reg[176][1]/P0001 , \wishbone_bd_ram_mem0_reg[176][2]/P0001 , \wishbone_bd_ram_mem0_reg[176][3]/P0001 , \wishbone_bd_ram_mem0_reg[176][4]/P0001 , \wishbone_bd_ram_mem0_reg[176][5]/P0001 , \wishbone_bd_ram_mem0_reg[176][6]/P0001 , \wishbone_bd_ram_mem0_reg[176][7]/P0001 , \wishbone_bd_ram_mem0_reg[177][0]/P0001 , \wishbone_bd_ram_mem0_reg[177][1]/P0001 , \wishbone_bd_ram_mem0_reg[177][2]/P0001 , \wishbone_bd_ram_mem0_reg[177][3]/P0001 , \wishbone_bd_ram_mem0_reg[177][4]/P0001 , \wishbone_bd_ram_mem0_reg[177][5]/P0001 , \wishbone_bd_ram_mem0_reg[177][6]/P0001 , \wishbone_bd_ram_mem0_reg[177][7]/P0001 , \wishbone_bd_ram_mem0_reg[178][0]/P0001 , \wishbone_bd_ram_mem0_reg[178][1]/P0001 , \wishbone_bd_ram_mem0_reg[178][2]/P0001 , \wishbone_bd_ram_mem0_reg[178][3]/P0001 , \wishbone_bd_ram_mem0_reg[178][4]/P0001 , \wishbone_bd_ram_mem0_reg[178][5]/P0001 , \wishbone_bd_ram_mem0_reg[178][6]/P0001 , \wishbone_bd_ram_mem0_reg[178][7]/P0001 , \wishbone_bd_ram_mem0_reg[179][0]/P0001 , \wishbone_bd_ram_mem0_reg[179][1]/P0001 , \wishbone_bd_ram_mem0_reg[179][2]/P0001 , \wishbone_bd_ram_mem0_reg[179][3]/P0001 , \wishbone_bd_ram_mem0_reg[179][4]/P0001 , \wishbone_bd_ram_mem0_reg[179][5]/P0001 , \wishbone_bd_ram_mem0_reg[179][6]/P0001 , \wishbone_bd_ram_mem0_reg[179][7]/P0001 , \wishbone_bd_ram_mem0_reg[17][0]/P0001 , \wishbone_bd_ram_mem0_reg[17][1]/P0001 , \wishbone_bd_ram_mem0_reg[17][2]/P0001 , \wishbone_bd_ram_mem0_reg[17][3]/P0001 , \wishbone_bd_ram_mem0_reg[17][4]/P0001 , \wishbone_bd_ram_mem0_reg[17][5]/P0001 , \wishbone_bd_ram_mem0_reg[17][6]/P0001 , \wishbone_bd_ram_mem0_reg[17][7]/P0001 , \wishbone_bd_ram_mem0_reg[180][0]/P0001 , \wishbone_bd_ram_mem0_reg[180][1]/P0001 , \wishbone_bd_ram_mem0_reg[180][2]/P0001 , \wishbone_bd_ram_mem0_reg[180][3]/P0001 , \wishbone_bd_ram_mem0_reg[180][4]/P0001 , \wishbone_bd_ram_mem0_reg[180][5]/P0001 , \wishbone_bd_ram_mem0_reg[180][6]/P0001 , \wishbone_bd_ram_mem0_reg[180][7]/P0001 , \wishbone_bd_ram_mem0_reg[181][0]/P0001 , \wishbone_bd_ram_mem0_reg[181][1]/P0001 , \wishbone_bd_ram_mem0_reg[181][2]/P0001 , \wishbone_bd_ram_mem0_reg[181][3]/P0001 , \wishbone_bd_ram_mem0_reg[181][4]/P0001 , \wishbone_bd_ram_mem0_reg[181][5]/P0001 , \wishbone_bd_ram_mem0_reg[181][6]/P0001 , \wishbone_bd_ram_mem0_reg[181][7]/P0001 , \wishbone_bd_ram_mem0_reg[182][0]/P0001 , \wishbone_bd_ram_mem0_reg[182][1]/P0001 , \wishbone_bd_ram_mem0_reg[182][2]/P0001 , \wishbone_bd_ram_mem0_reg[182][3]/P0001 , \wishbone_bd_ram_mem0_reg[182][4]/P0001 , \wishbone_bd_ram_mem0_reg[182][5]/P0001 , \wishbone_bd_ram_mem0_reg[182][6]/P0001 , \wishbone_bd_ram_mem0_reg[182][7]/P0001 , \wishbone_bd_ram_mem0_reg[183][0]/P0001 , \wishbone_bd_ram_mem0_reg[183][1]/P0001 , \wishbone_bd_ram_mem0_reg[183][2]/P0001 , \wishbone_bd_ram_mem0_reg[183][3]/P0001 , \wishbone_bd_ram_mem0_reg[183][4]/P0001 , \wishbone_bd_ram_mem0_reg[183][5]/P0001 , \wishbone_bd_ram_mem0_reg[183][6]/P0001 , \wishbone_bd_ram_mem0_reg[183][7]/P0001 , \wishbone_bd_ram_mem0_reg[184][0]/P0001 , \wishbone_bd_ram_mem0_reg[184][1]/P0001 , \wishbone_bd_ram_mem0_reg[184][2]/P0001 , \wishbone_bd_ram_mem0_reg[184][3]/P0001 , \wishbone_bd_ram_mem0_reg[184][4]/P0001 , \wishbone_bd_ram_mem0_reg[184][5]/P0001 , \wishbone_bd_ram_mem0_reg[184][6]/P0001 , \wishbone_bd_ram_mem0_reg[184][7]/P0001 , \wishbone_bd_ram_mem0_reg[185][0]/P0001 , \wishbone_bd_ram_mem0_reg[185][1]/P0001 , \wishbone_bd_ram_mem0_reg[185][2]/P0001 , \wishbone_bd_ram_mem0_reg[185][3]/P0001 , \wishbone_bd_ram_mem0_reg[185][4]/P0001 , \wishbone_bd_ram_mem0_reg[185][5]/P0001 , \wishbone_bd_ram_mem0_reg[185][6]/P0001 , \wishbone_bd_ram_mem0_reg[185][7]/P0001 , \wishbone_bd_ram_mem0_reg[186][0]/P0001 , \wishbone_bd_ram_mem0_reg[186][1]/P0001 , \wishbone_bd_ram_mem0_reg[186][2]/P0001 , \wishbone_bd_ram_mem0_reg[186][3]/P0001 , \wishbone_bd_ram_mem0_reg[186][4]/P0001 , \wishbone_bd_ram_mem0_reg[186][5]/P0001 , \wishbone_bd_ram_mem0_reg[186][6]/P0001 , \wishbone_bd_ram_mem0_reg[186][7]/P0001 , \wishbone_bd_ram_mem0_reg[187][0]/P0001 , \wishbone_bd_ram_mem0_reg[187][1]/P0001 , \wishbone_bd_ram_mem0_reg[187][2]/P0001 , \wishbone_bd_ram_mem0_reg[187][3]/P0001 , \wishbone_bd_ram_mem0_reg[187][4]/P0001 , \wishbone_bd_ram_mem0_reg[187][5]/P0001 , \wishbone_bd_ram_mem0_reg[187][6]/P0001 , \wishbone_bd_ram_mem0_reg[187][7]/P0001 , \wishbone_bd_ram_mem0_reg[188][0]/P0001 , \wishbone_bd_ram_mem0_reg[188][1]/P0001 , \wishbone_bd_ram_mem0_reg[188][2]/P0001 , \wishbone_bd_ram_mem0_reg[188][3]/P0001 , \wishbone_bd_ram_mem0_reg[188][4]/P0001 , \wishbone_bd_ram_mem0_reg[188][5]/P0001 , \wishbone_bd_ram_mem0_reg[188][6]/P0001 , \wishbone_bd_ram_mem0_reg[188][7]/P0001 , \wishbone_bd_ram_mem0_reg[189][0]/P0001 , \wishbone_bd_ram_mem0_reg[189][1]/P0001 , \wishbone_bd_ram_mem0_reg[189][2]/P0001 , \wishbone_bd_ram_mem0_reg[189][3]/P0001 , \wishbone_bd_ram_mem0_reg[189][4]/P0001 , \wishbone_bd_ram_mem0_reg[189][5]/P0001 , \wishbone_bd_ram_mem0_reg[189][6]/P0001 , \wishbone_bd_ram_mem0_reg[189][7]/P0001 , \wishbone_bd_ram_mem0_reg[18][0]/P0001 , \wishbone_bd_ram_mem0_reg[18][1]/P0001 , \wishbone_bd_ram_mem0_reg[18][2]/P0001 , \wishbone_bd_ram_mem0_reg[18][3]/P0001 , \wishbone_bd_ram_mem0_reg[18][4]/P0001 , \wishbone_bd_ram_mem0_reg[18][5]/P0001 , \wishbone_bd_ram_mem0_reg[18][6]/P0001 , \wishbone_bd_ram_mem0_reg[18][7]/P0001 , \wishbone_bd_ram_mem0_reg[190][0]/P0001 , \wishbone_bd_ram_mem0_reg[190][1]/P0001 , \wishbone_bd_ram_mem0_reg[190][2]/P0001 , \wishbone_bd_ram_mem0_reg[190][3]/P0001 , \wishbone_bd_ram_mem0_reg[190][4]/P0001 , \wishbone_bd_ram_mem0_reg[190][5]/P0001 , \wishbone_bd_ram_mem0_reg[190][6]/P0001 , \wishbone_bd_ram_mem0_reg[190][7]/P0001 , \wishbone_bd_ram_mem0_reg[191][0]/P0001 , \wishbone_bd_ram_mem0_reg[191][1]/P0001 , \wishbone_bd_ram_mem0_reg[191][2]/P0001 , \wishbone_bd_ram_mem0_reg[191][3]/P0001 , \wishbone_bd_ram_mem0_reg[191][4]/P0001 , \wishbone_bd_ram_mem0_reg[191][5]/P0001 , \wishbone_bd_ram_mem0_reg[191][6]/P0001 , \wishbone_bd_ram_mem0_reg[191][7]/P0001 , \wishbone_bd_ram_mem0_reg[192][0]/P0001 , \wishbone_bd_ram_mem0_reg[192][1]/P0001 , \wishbone_bd_ram_mem0_reg[192][2]/P0001 , \wishbone_bd_ram_mem0_reg[192][3]/P0001 , \wishbone_bd_ram_mem0_reg[192][4]/P0001 , \wishbone_bd_ram_mem0_reg[192][5]/P0001 , \wishbone_bd_ram_mem0_reg[192][6]/P0001 , \wishbone_bd_ram_mem0_reg[192][7]/P0001 , \wishbone_bd_ram_mem0_reg[193][0]/P0001 , \wishbone_bd_ram_mem0_reg[193][1]/P0001 , \wishbone_bd_ram_mem0_reg[193][2]/P0001 , \wishbone_bd_ram_mem0_reg[193][3]/P0001 , \wishbone_bd_ram_mem0_reg[193][4]/P0001 , \wishbone_bd_ram_mem0_reg[193][5]/P0001 , \wishbone_bd_ram_mem0_reg[193][6]/P0001 , \wishbone_bd_ram_mem0_reg[193][7]/P0001 , \wishbone_bd_ram_mem0_reg[194][0]/P0001 , \wishbone_bd_ram_mem0_reg[194][1]/P0001 , \wishbone_bd_ram_mem0_reg[194][2]/P0001 , \wishbone_bd_ram_mem0_reg[194][3]/P0001 , \wishbone_bd_ram_mem0_reg[194][4]/P0001 , \wishbone_bd_ram_mem0_reg[194][5]/P0001 , \wishbone_bd_ram_mem0_reg[194][6]/P0001 , \wishbone_bd_ram_mem0_reg[194][7]/P0001 , \wishbone_bd_ram_mem0_reg[195][0]/P0001 , \wishbone_bd_ram_mem0_reg[195][1]/P0001 , \wishbone_bd_ram_mem0_reg[195][2]/P0001 , \wishbone_bd_ram_mem0_reg[195][3]/P0001 , \wishbone_bd_ram_mem0_reg[195][4]/P0001 , \wishbone_bd_ram_mem0_reg[195][5]/P0001 , \wishbone_bd_ram_mem0_reg[195][6]/P0001 , \wishbone_bd_ram_mem0_reg[195][7]/P0001 , \wishbone_bd_ram_mem0_reg[196][0]/P0001 , \wishbone_bd_ram_mem0_reg[196][1]/P0001 , \wishbone_bd_ram_mem0_reg[196][2]/P0001 , \wishbone_bd_ram_mem0_reg[196][3]/P0001 , \wishbone_bd_ram_mem0_reg[196][4]/P0001 , \wishbone_bd_ram_mem0_reg[196][5]/P0001 , \wishbone_bd_ram_mem0_reg[196][6]/P0001 , \wishbone_bd_ram_mem0_reg[196][7]/P0001 , \wishbone_bd_ram_mem0_reg[197][0]/P0001 , \wishbone_bd_ram_mem0_reg[197][1]/P0001 , \wishbone_bd_ram_mem0_reg[197][2]/P0001 , \wishbone_bd_ram_mem0_reg[197][3]/P0001 , \wishbone_bd_ram_mem0_reg[197][4]/P0001 , \wishbone_bd_ram_mem0_reg[197][5]/P0001 , \wishbone_bd_ram_mem0_reg[197][6]/P0001 , \wishbone_bd_ram_mem0_reg[197][7]/P0001 , \wishbone_bd_ram_mem0_reg[198][0]/P0001 , \wishbone_bd_ram_mem0_reg[198][1]/P0001 , \wishbone_bd_ram_mem0_reg[198][2]/P0001 , \wishbone_bd_ram_mem0_reg[198][3]/P0001 , \wishbone_bd_ram_mem0_reg[198][4]/P0001 , \wishbone_bd_ram_mem0_reg[198][5]/P0001 , \wishbone_bd_ram_mem0_reg[198][6]/P0001 , \wishbone_bd_ram_mem0_reg[198][7]/P0001 , \wishbone_bd_ram_mem0_reg[199][0]/P0001 , \wishbone_bd_ram_mem0_reg[199][1]/P0001 , \wishbone_bd_ram_mem0_reg[199][2]/P0001 , \wishbone_bd_ram_mem0_reg[199][3]/P0001 , \wishbone_bd_ram_mem0_reg[199][4]/P0001 , \wishbone_bd_ram_mem0_reg[199][5]/P0001 , \wishbone_bd_ram_mem0_reg[199][6]/P0001 , \wishbone_bd_ram_mem0_reg[199][7]/P0001 , \wishbone_bd_ram_mem0_reg[19][0]/P0001 , \wishbone_bd_ram_mem0_reg[19][1]/P0001 , \wishbone_bd_ram_mem0_reg[19][2]/P0001 , \wishbone_bd_ram_mem0_reg[19][3]/P0001 , \wishbone_bd_ram_mem0_reg[19][4]/P0001 , \wishbone_bd_ram_mem0_reg[19][5]/P0001 , \wishbone_bd_ram_mem0_reg[19][6]/P0001 , \wishbone_bd_ram_mem0_reg[19][7]/P0001 , \wishbone_bd_ram_mem0_reg[1][0]/P0001 , \wishbone_bd_ram_mem0_reg[1][1]/P0001 , \wishbone_bd_ram_mem0_reg[1][2]/P0001 , \wishbone_bd_ram_mem0_reg[1][3]/P0001 , \wishbone_bd_ram_mem0_reg[1][4]/P0001 , \wishbone_bd_ram_mem0_reg[1][5]/P0001 , \wishbone_bd_ram_mem0_reg[1][6]/P0001 , \wishbone_bd_ram_mem0_reg[1][7]/P0001 , \wishbone_bd_ram_mem0_reg[200][0]/P0001 , \wishbone_bd_ram_mem0_reg[200][1]/P0001 , \wishbone_bd_ram_mem0_reg[200][2]/P0001 , \wishbone_bd_ram_mem0_reg[200][3]/P0001 , \wishbone_bd_ram_mem0_reg[200][4]/P0001 , \wishbone_bd_ram_mem0_reg[200][5]/P0001 , \wishbone_bd_ram_mem0_reg[200][6]/P0001 , \wishbone_bd_ram_mem0_reg[200][7]/P0001 , \wishbone_bd_ram_mem0_reg[201][0]/P0001 , \wishbone_bd_ram_mem0_reg[201][1]/P0001 , \wishbone_bd_ram_mem0_reg[201][2]/P0001 , \wishbone_bd_ram_mem0_reg[201][3]/P0001 , \wishbone_bd_ram_mem0_reg[201][4]/P0001 , \wishbone_bd_ram_mem0_reg[201][5]/P0001 , \wishbone_bd_ram_mem0_reg[201][6]/P0001 , \wishbone_bd_ram_mem0_reg[201][7]/P0001 , \wishbone_bd_ram_mem0_reg[202][0]/P0001 , \wishbone_bd_ram_mem0_reg[202][1]/P0001 , \wishbone_bd_ram_mem0_reg[202][2]/P0001 , \wishbone_bd_ram_mem0_reg[202][3]/P0001 , \wishbone_bd_ram_mem0_reg[202][4]/P0001 , \wishbone_bd_ram_mem0_reg[202][5]/P0001 , \wishbone_bd_ram_mem0_reg[202][6]/P0001 , \wishbone_bd_ram_mem0_reg[202][7]/P0001 , \wishbone_bd_ram_mem0_reg[203][0]/P0001 , \wishbone_bd_ram_mem0_reg[203][1]/P0001 , \wishbone_bd_ram_mem0_reg[203][2]/P0001 , \wishbone_bd_ram_mem0_reg[203][3]/P0001 , \wishbone_bd_ram_mem0_reg[203][4]/P0001 , \wishbone_bd_ram_mem0_reg[203][5]/P0001 , \wishbone_bd_ram_mem0_reg[203][6]/P0001 , \wishbone_bd_ram_mem0_reg[203][7]/P0001 , \wishbone_bd_ram_mem0_reg[204][0]/P0001 , \wishbone_bd_ram_mem0_reg[204][1]/P0001 , \wishbone_bd_ram_mem0_reg[204][2]/P0001 , \wishbone_bd_ram_mem0_reg[204][3]/P0001 , \wishbone_bd_ram_mem0_reg[204][4]/P0001 , \wishbone_bd_ram_mem0_reg[204][5]/P0001 , \wishbone_bd_ram_mem0_reg[204][6]/P0001 , \wishbone_bd_ram_mem0_reg[204][7]/P0001 , \wishbone_bd_ram_mem0_reg[205][0]/P0001 , \wishbone_bd_ram_mem0_reg[205][1]/P0001 , \wishbone_bd_ram_mem0_reg[205][2]/P0001 , \wishbone_bd_ram_mem0_reg[205][3]/P0001 , \wishbone_bd_ram_mem0_reg[205][4]/P0001 , \wishbone_bd_ram_mem0_reg[205][5]/P0001 , \wishbone_bd_ram_mem0_reg[205][6]/P0001 , \wishbone_bd_ram_mem0_reg[205][7]/P0001 , \wishbone_bd_ram_mem0_reg[206][0]/P0001 , \wishbone_bd_ram_mem0_reg[206][1]/P0001 , \wishbone_bd_ram_mem0_reg[206][2]/P0001 , \wishbone_bd_ram_mem0_reg[206][3]/P0001 , \wishbone_bd_ram_mem0_reg[206][4]/P0001 , \wishbone_bd_ram_mem0_reg[206][5]/P0001 , \wishbone_bd_ram_mem0_reg[206][6]/P0001 , \wishbone_bd_ram_mem0_reg[206][7]/P0001 , \wishbone_bd_ram_mem0_reg[207][0]/P0001 , \wishbone_bd_ram_mem0_reg[207][1]/P0001 , \wishbone_bd_ram_mem0_reg[207][2]/P0001 , \wishbone_bd_ram_mem0_reg[207][3]/P0001 , \wishbone_bd_ram_mem0_reg[207][4]/P0001 , \wishbone_bd_ram_mem0_reg[207][5]/P0001 , \wishbone_bd_ram_mem0_reg[207][6]/P0001 , \wishbone_bd_ram_mem0_reg[207][7]/P0001 , \wishbone_bd_ram_mem0_reg[208][0]/P0001 , \wishbone_bd_ram_mem0_reg[208][1]/P0001 , \wishbone_bd_ram_mem0_reg[208][2]/P0001 , \wishbone_bd_ram_mem0_reg[208][3]/P0001 , \wishbone_bd_ram_mem0_reg[208][4]/P0001 , \wishbone_bd_ram_mem0_reg[208][5]/P0001 , \wishbone_bd_ram_mem0_reg[208][6]/P0001 , \wishbone_bd_ram_mem0_reg[208][7]/P0001 , \wishbone_bd_ram_mem0_reg[209][0]/P0001 , \wishbone_bd_ram_mem0_reg[209][1]/P0001 , \wishbone_bd_ram_mem0_reg[209][2]/P0001 , \wishbone_bd_ram_mem0_reg[209][3]/P0001 , \wishbone_bd_ram_mem0_reg[209][4]/P0001 , \wishbone_bd_ram_mem0_reg[209][5]/P0001 , \wishbone_bd_ram_mem0_reg[209][6]/P0001 , \wishbone_bd_ram_mem0_reg[209][7]/P0001 , \wishbone_bd_ram_mem0_reg[20][0]/P0001 , \wishbone_bd_ram_mem0_reg[20][1]/P0001 , \wishbone_bd_ram_mem0_reg[20][2]/P0001 , \wishbone_bd_ram_mem0_reg[20][3]/P0001 , \wishbone_bd_ram_mem0_reg[20][4]/P0001 , \wishbone_bd_ram_mem0_reg[20][5]/P0001 , \wishbone_bd_ram_mem0_reg[20][6]/P0001 , \wishbone_bd_ram_mem0_reg[20][7]/P0001 , \wishbone_bd_ram_mem0_reg[210][0]/P0001 , \wishbone_bd_ram_mem0_reg[210][1]/P0001 , \wishbone_bd_ram_mem0_reg[210][2]/P0001 , \wishbone_bd_ram_mem0_reg[210][3]/P0001 , \wishbone_bd_ram_mem0_reg[210][4]/P0001 , \wishbone_bd_ram_mem0_reg[210][5]/P0001 , \wishbone_bd_ram_mem0_reg[210][6]/P0001 , \wishbone_bd_ram_mem0_reg[210][7]/P0001 , \wishbone_bd_ram_mem0_reg[211][0]/P0001 , \wishbone_bd_ram_mem0_reg[211][1]/P0001 , \wishbone_bd_ram_mem0_reg[211][2]/P0001 , \wishbone_bd_ram_mem0_reg[211][3]/P0001 , \wishbone_bd_ram_mem0_reg[211][4]/P0001 , \wishbone_bd_ram_mem0_reg[211][5]/P0001 , \wishbone_bd_ram_mem0_reg[211][6]/P0001 , \wishbone_bd_ram_mem0_reg[211][7]/P0001 , \wishbone_bd_ram_mem0_reg[212][0]/P0001 , \wishbone_bd_ram_mem0_reg[212][1]/P0001 , \wishbone_bd_ram_mem0_reg[212][2]/P0001 , \wishbone_bd_ram_mem0_reg[212][3]/P0001 , \wishbone_bd_ram_mem0_reg[212][4]/P0001 , \wishbone_bd_ram_mem0_reg[212][5]/P0001 , \wishbone_bd_ram_mem0_reg[212][6]/P0001 , \wishbone_bd_ram_mem0_reg[212][7]/P0001 , \wishbone_bd_ram_mem0_reg[213][0]/P0001 , \wishbone_bd_ram_mem0_reg[213][1]/P0001 , \wishbone_bd_ram_mem0_reg[213][2]/P0001 , \wishbone_bd_ram_mem0_reg[213][3]/P0001 , \wishbone_bd_ram_mem0_reg[213][4]/P0001 , \wishbone_bd_ram_mem0_reg[213][5]/P0001 , \wishbone_bd_ram_mem0_reg[213][6]/P0001 , \wishbone_bd_ram_mem0_reg[213][7]/P0001 , \wishbone_bd_ram_mem0_reg[214][0]/P0001 , \wishbone_bd_ram_mem0_reg[214][1]/P0001 , \wishbone_bd_ram_mem0_reg[214][2]/P0001 , \wishbone_bd_ram_mem0_reg[214][3]/P0001 , \wishbone_bd_ram_mem0_reg[214][4]/P0001 , \wishbone_bd_ram_mem0_reg[214][5]/P0001 , \wishbone_bd_ram_mem0_reg[214][6]/P0001 , \wishbone_bd_ram_mem0_reg[214][7]/P0001 , \wishbone_bd_ram_mem0_reg[215][0]/P0001 , \wishbone_bd_ram_mem0_reg[215][1]/P0001 , \wishbone_bd_ram_mem0_reg[215][2]/P0001 , \wishbone_bd_ram_mem0_reg[215][3]/P0001 , \wishbone_bd_ram_mem0_reg[215][4]/P0001 , \wishbone_bd_ram_mem0_reg[215][5]/P0001 , \wishbone_bd_ram_mem0_reg[215][6]/P0001 , \wishbone_bd_ram_mem0_reg[215][7]/P0001 , \wishbone_bd_ram_mem0_reg[216][0]/P0001 , \wishbone_bd_ram_mem0_reg[216][1]/P0001 , \wishbone_bd_ram_mem0_reg[216][2]/P0001 , \wishbone_bd_ram_mem0_reg[216][3]/P0001 , \wishbone_bd_ram_mem0_reg[216][4]/P0001 , \wishbone_bd_ram_mem0_reg[216][5]/P0001 , \wishbone_bd_ram_mem0_reg[216][6]/P0001 , \wishbone_bd_ram_mem0_reg[216][7]/P0001 , \wishbone_bd_ram_mem0_reg[217][0]/P0001 , \wishbone_bd_ram_mem0_reg[217][1]/P0001 , \wishbone_bd_ram_mem0_reg[217][2]/P0001 , \wishbone_bd_ram_mem0_reg[217][3]/P0001 , \wishbone_bd_ram_mem0_reg[217][4]/P0001 , \wishbone_bd_ram_mem0_reg[217][5]/P0001 , \wishbone_bd_ram_mem0_reg[217][6]/P0001 , \wishbone_bd_ram_mem0_reg[217][7]/P0001 , \wishbone_bd_ram_mem0_reg[218][0]/P0001 , \wishbone_bd_ram_mem0_reg[218][1]/P0001 , \wishbone_bd_ram_mem0_reg[218][2]/P0001 , \wishbone_bd_ram_mem0_reg[218][3]/P0001 , \wishbone_bd_ram_mem0_reg[218][4]/P0001 , \wishbone_bd_ram_mem0_reg[218][5]/P0001 , \wishbone_bd_ram_mem0_reg[218][6]/P0001 , \wishbone_bd_ram_mem0_reg[218][7]/P0001 , \wishbone_bd_ram_mem0_reg[219][0]/P0001 , \wishbone_bd_ram_mem0_reg[219][1]/P0001 , \wishbone_bd_ram_mem0_reg[219][2]/P0001 , \wishbone_bd_ram_mem0_reg[219][3]/P0001 , \wishbone_bd_ram_mem0_reg[219][4]/P0001 , \wishbone_bd_ram_mem0_reg[219][5]/P0001 , \wishbone_bd_ram_mem0_reg[219][6]/P0001 , \wishbone_bd_ram_mem0_reg[219][7]/P0001 , \wishbone_bd_ram_mem0_reg[21][0]/P0001 , \wishbone_bd_ram_mem0_reg[21][1]/P0001 , \wishbone_bd_ram_mem0_reg[21][2]/P0001 , \wishbone_bd_ram_mem0_reg[21][3]/P0001 , \wishbone_bd_ram_mem0_reg[21][4]/P0001 , \wishbone_bd_ram_mem0_reg[21][5]/P0001 , \wishbone_bd_ram_mem0_reg[21][6]/P0001 , \wishbone_bd_ram_mem0_reg[21][7]/P0001 , \wishbone_bd_ram_mem0_reg[220][0]/P0001 , \wishbone_bd_ram_mem0_reg[220][1]/P0001 , \wishbone_bd_ram_mem0_reg[220][2]/P0001 , \wishbone_bd_ram_mem0_reg[220][3]/P0001 , \wishbone_bd_ram_mem0_reg[220][4]/P0001 , \wishbone_bd_ram_mem0_reg[220][5]/P0001 , \wishbone_bd_ram_mem0_reg[220][6]/P0001 , \wishbone_bd_ram_mem0_reg[220][7]/P0001 , \wishbone_bd_ram_mem0_reg[221][0]/P0001 , \wishbone_bd_ram_mem0_reg[221][1]/P0001 , \wishbone_bd_ram_mem0_reg[221][2]/P0001 , \wishbone_bd_ram_mem0_reg[221][3]/P0001 , \wishbone_bd_ram_mem0_reg[221][4]/P0001 , \wishbone_bd_ram_mem0_reg[221][5]/P0001 , \wishbone_bd_ram_mem0_reg[221][6]/P0001 , \wishbone_bd_ram_mem0_reg[221][7]/P0001 , \wishbone_bd_ram_mem0_reg[222][0]/P0001 , \wishbone_bd_ram_mem0_reg[222][1]/P0001 , \wishbone_bd_ram_mem0_reg[222][2]/P0001 , \wishbone_bd_ram_mem0_reg[222][3]/P0001 , \wishbone_bd_ram_mem0_reg[222][4]/P0001 , \wishbone_bd_ram_mem0_reg[222][5]/P0001 , \wishbone_bd_ram_mem0_reg[222][6]/P0001 , \wishbone_bd_ram_mem0_reg[222][7]/P0001 , \wishbone_bd_ram_mem0_reg[223][0]/P0001 , \wishbone_bd_ram_mem0_reg[223][1]/P0001 , \wishbone_bd_ram_mem0_reg[223][2]/P0001 , \wishbone_bd_ram_mem0_reg[223][3]/P0001 , \wishbone_bd_ram_mem0_reg[223][4]/P0001 , \wishbone_bd_ram_mem0_reg[223][5]/P0001 , \wishbone_bd_ram_mem0_reg[223][6]/P0001 , \wishbone_bd_ram_mem0_reg[223][7]/P0001 , \wishbone_bd_ram_mem0_reg[224][0]/P0001 , \wishbone_bd_ram_mem0_reg[224][1]/P0001 , \wishbone_bd_ram_mem0_reg[224][2]/P0001 , \wishbone_bd_ram_mem0_reg[224][3]/P0001 , \wishbone_bd_ram_mem0_reg[224][4]/P0001 , \wishbone_bd_ram_mem0_reg[224][5]/P0001 , \wishbone_bd_ram_mem0_reg[224][6]/P0001 , \wishbone_bd_ram_mem0_reg[224][7]/P0001 , \wishbone_bd_ram_mem0_reg[225][0]/P0001 , \wishbone_bd_ram_mem0_reg[225][1]/P0001 , \wishbone_bd_ram_mem0_reg[225][2]/P0001 , \wishbone_bd_ram_mem0_reg[225][3]/P0001 , \wishbone_bd_ram_mem0_reg[225][4]/P0001 , \wishbone_bd_ram_mem0_reg[225][5]/P0001 , \wishbone_bd_ram_mem0_reg[225][6]/P0001 , \wishbone_bd_ram_mem0_reg[225][7]/P0001 , \wishbone_bd_ram_mem0_reg[226][0]/P0001 , \wishbone_bd_ram_mem0_reg[226][1]/P0001 , \wishbone_bd_ram_mem0_reg[226][2]/P0001 , \wishbone_bd_ram_mem0_reg[226][3]/P0001 , \wishbone_bd_ram_mem0_reg[226][4]/P0001 , \wishbone_bd_ram_mem0_reg[226][5]/P0001 , \wishbone_bd_ram_mem0_reg[226][6]/P0001 , \wishbone_bd_ram_mem0_reg[226][7]/P0001 , \wishbone_bd_ram_mem0_reg[227][0]/P0001 , \wishbone_bd_ram_mem0_reg[227][1]/P0001 , \wishbone_bd_ram_mem0_reg[227][2]/P0001 , \wishbone_bd_ram_mem0_reg[227][3]/P0001 , \wishbone_bd_ram_mem0_reg[227][4]/P0001 , \wishbone_bd_ram_mem0_reg[227][5]/P0001 , \wishbone_bd_ram_mem0_reg[227][6]/P0001 , \wishbone_bd_ram_mem0_reg[227][7]/P0001 , \wishbone_bd_ram_mem0_reg[228][0]/P0001 , \wishbone_bd_ram_mem0_reg[228][1]/P0001 , \wishbone_bd_ram_mem0_reg[228][2]/P0001 , \wishbone_bd_ram_mem0_reg[228][3]/P0001 , \wishbone_bd_ram_mem0_reg[228][4]/P0001 , \wishbone_bd_ram_mem0_reg[228][5]/P0001 , \wishbone_bd_ram_mem0_reg[228][6]/P0001 , \wishbone_bd_ram_mem0_reg[228][7]/P0001 , \wishbone_bd_ram_mem0_reg[229][0]/P0001 , \wishbone_bd_ram_mem0_reg[229][1]/P0001 , \wishbone_bd_ram_mem0_reg[229][2]/P0001 , \wishbone_bd_ram_mem0_reg[229][3]/P0001 , \wishbone_bd_ram_mem0_reg[229][4]/P0001 , \wishbone_bd_ram_mem0_reg[229][5]/P0001 , \wishbone_bd_ram_mem0_reg[229][6]/P0001 , \wishbone_bd_ram_mem0_reg[229][7]/P0001 , \wishbone_bd_ram_mem0_reg[22][0]/P0001 , \wishbone_bd_ram_mem0_reg[22][1]/P0001 , \wishbone_bd_ram_mem0_reg[22][2]/P0001 , \wishbone_bd_ram_mem0_reg[22][3]/P0001 , \wishbone_bd_ram_mem0_reg[22][4]/P0001 , \wishbone_bd_ram_mem0_reg[22][5]/P0001 , \wishbone_bd_ram_mem0_reg[22][6]/P0001 , \wishbone_bd_ram_mem0_reg[22][7]/P0001 , \wishbone_bd_ram_mem0_reg[230][0]/P0001 , \wishbone_bd_ram_mem0_reg[230][1]/P0001 , \wishbone_bd_ram_mem0_reg[230][2]/P0001 , \wishbone_bd_ram_mem0_reg[230][3]/P0001 , \wishbone_bd_ram_mem0_reg[230][4]/P0001 , \wishbone_bd_ram_mem0_reg[230][5]/P0001 , \wishbone_bd_ram_mem0_reg[230][6]/P0001 , \wishbone_bd_ram_mem0_reg[230][7]/P0001 , \wishbone_bd_ram_mem0_reg[231][0]/P0001 , \wishbone_bd_ram_mem0_reg[231][1]/P0001 , \wishbone_bd_ram_mem0_reg[231][2]/P0001 , \wishbone_bd_ram_mem0_reg[231][3]/P0001 , \wishbone_bd_ram_mem0_reg[231][4]/P0001 , \wishbone_bd_ram_mem0_reg[231][5]/P0001 , \wishbone_bd_ram_mem0_reg[231][6]/P0001 , \wishbone_bd_ram_mem0_reg[231][7]/P0001 , \wishbone_bd_ram_mem0_reg[232][0]/P0001 , \wishbone_bd_ram_mem0_reg[232][1]/P0001 , \wishbone_bd_ram_mem0_reg[232][2]/P0001 , \wishbone_bd_ram_mem0_reg[232][3]/P0001 , \wishbone_bd_ram_mem0_reg[232][4]/P0001 , \wishbone_bd_ram_mem0_reg[232][5]/P0001 , \wishbone_bd_ram_mem0_reg[232][6]/P0001 , \wishbone_bd_ram_mem0_reg[232][7]/P0001 , \wishbone_bd_ram_mem0_reg[233][0]/P0001 , \wishbone_bd_ram_mem0_reg[233][1]/P0001 , \wishbone_bd_ram_mem0_reg[233][2]/P0001 , \wishbone_bd_ram_mem0_reg[233][3]/P0001 , \wishbone_bd_ram_mem0_reg[233][4]/P0001 , \wishbone_bd_ram_mem0_reg[233][5]/P0001 , \wishbone_bd_ram_mem0_reg[233][6]/P0001 , \wishbone_bd_ram_mem0_reg[233][7]/P0001 , \wishbone_bd_ram_mem0_reg[234][0]/P0001 , \wishbone_bd_ram_mem0_reg[234][1]/P0001 , \wishbone_bd_ram_mem0_reg[234][2]/P0001 , \wishbone_bd_ram_mem0_reg[234][3]/P0001 , \wishbone_bd_ram_mem0_reg[234][4]/P0001 , \wishbone_bd_ram_mem0_reg[234][5]/P0001 , \wishbone_bd_ram_mem0_reg[234][6]/P0001 , \wishbone_bd_ram_mem0_reg[234][7]/P0001 , \wishbone_bd_ram_mem0_reg[235][0]/P0001 , \wishbone_bd_ram_mem0_reg[235][1]/P0001 , \wishbone_bd_ram_mem0_reg[235][2]/P0001 , \wishbone_bd_ram_mem0_reg[235][3]/P0001 , \wishbone_bd_ram_mem0_reg[235][4]/P0001 , \wishbone_bd_ram_mem0_reg[235][5]/P0001 , \wishbone_bd_ram_mem0_reg[235][6]/P0001 , \wishbone_bd_ram_mem0_reg[235][7]/P0001 , \wishbone_bd_ram_mem0_reg[236][0]/P0001 , \wishbone_bd_ram_mem0_reg[236][1]/P0001 , \wishbone_bd_ram_mem0_reg[236][2]/P0001 , \wishbone_bd_ram_mem0_reg[236][3]/P0001 , \wishbone_bd_ram_mem0_reg[236][4]/P0001 , \wishbone_bd_ram_mem0_reg[236][5]/P0001 , \wishbone_bd_ram_mem0_reg[236][6]/P0001 , \wishbone_bd_ram_mem0_reg[236][7]/P0001 , \wishbone_bd_ram_mem0_reg[237][0]/P0001 , \wishbone_bd_ram_mem0_reg[237][1]/P0001 , \wishbone_bd_ram_mem0_reg[237][2]/P0001 , \wishbone_bd_ram_mem0_reg[237][3]/P0001 , \wishbone_bd_ram_mem0_reg[237][4]/P0001 , \wishbone_bd_ram_mem0_reg[237][5]/P0001 , \wishbone_bd_ram_mem0_reg[237][6]/P0001 , \wishbone_bd_ram_mem0_reg[237][7]/P0001 , \wishbone_bd_ram_mem0_reg[238][0]/P0001 , \wishbone_bd_ram_mem0_reg[238][1]/P0001 , \wishbone_bd_ram_mem0_reg[238][2]/P0001 , \wishbone_bd_ram_mem0_reg[238][3]/P0001 , \wishbone_bd_ram_mem0_reg[238][4]/P0001 , \wishbone_bd_ram_mem0_reg[238][5]/P0001 , \wishbone_bd_ram_mem0_reg[238][6]/P0001 , \wishbone_bd_ram_mem0_reg[238][7]/P0001 , \wishbone_bd_ram_mem0_reg[239][0]/P0001 , \wishbone_bd_ram_mem0_reg[239][1]/P0001 , \wishbone_bd_ram_mem0_reg[239][2]/P0001 , \wishbone_bd_ram_mem0_reg[239][3]/P0001 , \wishbone_bd_ram_mem0_reg[239][4]/P0001 , \wishbone_bd_ram_mem0_reg[239][5]/P0001 , \wishbone_bd_ram_mem0_reg[239][6]/P0001 , \wishbone_bd_ram_mem0_reg[239][7]/P0001 , \wishbone_bd_ram_mem0_reg[23][0]/P0001 , \wishbone_bd_ram_mem0_reg[23][1]/P0001 , \wishbone_bd_ram_mem0_reg[23][2]/P0001 , \wishbone_bd_ram_mem0_reg[23][3]/P0001 , \wishbone_bd_ram_mem0_reg[23][4]/P0001 , \wishbone_bd_ram_mem0_reg[23][5]/P0001 , \wishbone_bd_ram_mem0_reg[23][6]/P0001 , \wishbone_bd_ram_mem0_reg[23][7]/P0001 , \wishbone_bd_ram_mem0_reg[240][0]/P0001 , \wishbone_bd_ram_mem0_reg[240][1]/P0001 , \wishbone_bd_ram_mem0_reg[240][2]/P0001 , \wishbone_bd_ram_mem0_reg[240][3]/P0001 , \wishbone_bd_ram_mem0_reg[240][4]/P0001 , \wishbone_bd_ram_mem0_reg[240][5]/P0001 , \wishbone_bd_ram_mem0_reg[240][6]/P0001 , \wishbone_bd_ram_mem0_reg[240][7]/P0001 , \wishbone_bd_ram_mem0_reg[241][0]/P0001 , \wishbone_bd_ram_mem0_reg[241][1]/P0001 , \wishbone_bd_ram_mem0_reg[241][2]/P0001 , \wishbone_bd_ram_mem0_reg[241][3]/P0001 , \wishbone_bd_ram_mem0_reg[241][4]/P0001 , \wishbone_bd_ram_mem0_reg[241][5]/P0001 , \wishbone_bd_ram_mem0_reg[241][6]/P0001 , \wishbone_bd_ram_mem0_reg[241][7]/P0001 , \wishbone_bd_ram_mem0_reg[242][0]/P0001 , \wishbone_bd_ram_mem0_reg[242][1]/P0001 , \wishbone_bd_ram_mem0_reg[242][2]/P0001 , \wishbone_bd_ram_mem0_reg[242][3]/P0001 , \wishbone_bd_ram_mem0_reg[242][4]/P0001 , \wishbone_bd_ram_mem0_reg[242][5]/P0001 , \wishbone_bd_ram_mem0_reg[242][6]/P0001 , \wishbone_bd_ram_mem0_reg[242][7]/P0001 , \wishbone_bd_ram_mem0_reg[243][0]/P0001 , \wishbone_bd_ram_mem0_reg[243][1]/P0001 , \wishbone_bd_ram_mem0_reg[243][2]/P0001 , \wishbone_bd_ram_mem0_reg[243][3]/P0001 , \wishbone_bd_ram_mem0_reg[243][4]/P0001 , \wishbone_bd_ram_mem0_reg[243][5]/P0001 , \wishbone_bd_ram_mem0_reg[243][6]/P0001 , \wishbone_bd_ram_mem0_reg[243][7]/P0001 , \wishbone_bd_ram_mem0_reg[244][0]/P0001 , \wishbone_bd_ram_mem0_reg[244][1]/P0001 , \wishbone_bd_ram_mem0_reg[244][2]/P0001 , \wishbone_bd_ram_mem0_reg[244][3]/P0001 , \wishbone_bd_ram_mem0_reg[244][4]/P0001 , \wishbone_bd_ram_mem0_reg[244][5]/P0001 , \wishbone_bd_ram_mem0_reg[244][6]/P0001 , \wishbone_bd_ram_mem0_reg[244][7]/P0001 , \wishbone_bd_ram_mem0_reg[245][0]/P0001 , \wishbone_bd_ram_mem0_reg[245][1]/P0001 , \wishbone_bd_ram_mem0_reg[245][2]/P0001 , \wishbone_bd_ram_mem0_reg[245][3]/P0001 , \wishbone_bd_ram_mem0_reg[245][4]/P0001 , \wishbone_bd_ram_mem0_reg[245][5]/P0001 , \wishbone_bd_ram_mem0_reg[245][6]/P0001 , \wishbone_bd_ram_mem0_reg[245][7]/P0001 , \wishbone_bd_ram_mem0_reg[246][0]/P0001 , \wishbone_bd_ram_mem0_reg[246][1]/P0001 , \wishbone_bd_ram_mem0_reg[246][2]/P0001 , \wishbone_bd_ram_mem0_reg[246][3]/P0001 , \wishbone_bd_ram_mem0_reg[246][4]/P0001 , \wishbone_bd_ram_mem0_reg[246][5]/P0001 , \wishbone_bd_ram_mem0_reg[246][6]/P0001 , \wishbone_bd_ram_mem0_reg[246][7]/P0001 , \wishbone_bd_ram_mem0_reg[247][0]/P0001 , \wishbone_bd_ram_mem0_reg[247][1]/P0001 , \wishbone_bd_ram_mem0_reg[247][2]/P0001 , \wishbone_bd_ram_mem0_reg[247][3]/P0001 , \wishbone_bd_ram_mem0_reg[247][4]/P0001 , \wishbone_bd_ram_mem0_reg[247][5]/P0001 , \wishbone_bd_ram_mem0_reg[247][6]/P0001 , \wishbone_bd_ram_mem0_reg[247][7]/P0001 , \wishbone_bd_ram_mem0_reg[248][0]/P0001 , \wishbone_bd_ram_mem0_reg[248][1]/P0001 , \wishbone_bd_ram_mem0_reg[248][2]/P0001 , \wishbone_bd_ram_mem0_reg[248][3]/P0001 , \wishbone_bd_ram_mem0_reg[248][4]/P0001 , \wishbone_bd_ram_mem0_reg[248][5]/P0001 , \wishbone_bd_ram_mem0_reg[248][6]/P0001 , \wishbone_bd_ram_mem0_reg[248][7]/P0001 , \wishbone_bd_ram_mem0_reg[249][0]/P0001 , \wishbone_bd_ram_mem0_reg[249][1]/P0001 , \wishbone_bd_ram_mem0_reg[249][2]/P0001 , \wishbone_bd_ram_mem0_reg[249][3]/P0001 , \wishbone_bd_ram_mem0_reg[249][4]/P0001 , \wishbone_bd_ram_mem0_reg[249][5]/P0001 , \wishbone_bd_ram_mem0_reg[249][6]/P0001 , \wishbone_bd_ram_mem0_reg[249][7]/P0001 , \wishbone_bd_ram_mem0_reg[24][0]/P0001 , \wishbone_bd_ram_mem0_reg[24][1]/P0001 , \wishbone_bd_ram_mem0_reg[24][2]/P0001 , \wishbone_bd_ram_mem0_reg[24][3]/P0001 , \wishbone_bd_ram_mem0_reg[24][4]/P0001 , \wishbone_bd_ram_mem0_reg[24][5]/P0001 , \wishbone_bd_ram_mem0_reg[24][6]/P0001 , \wishbone_bd_ram_mem0_reg[24][7]/P0001 , \wishbone_bd_ram_mem0_reg[250][0]/P0001 , \wishbone_bd_ram_mem0_reg[250][1]/P0001 , \wishbone_bd_ram_mem0_reg[250][2]/P0001 , \wishbone_bd_ram_mem0_reg[250][3]/P0001 , \wishbone_bd_ram_mem0_reg[250][4]/P0001 , \wishbone_bd_ram_mem0_reg[250][5]/P0001 , \wishbone_bd_ram_mem0_reg[250][6]/P0001 , \wishbone_bd_ram_mem0_reg[250][7]/P0001 , \wishbone_bd_ram_mem0_reg[251][0]/P0001 , \wishbone_bd_ram_mem0_reg[251][1]/P0001 , \wishbone_bd_ram_mem0_reg[251][2]/P0001 , \wishbone_bd_ram_mem0_reg[251][3]/P0001 , \wishbone_bd_ram_mem0_reg[251][4]/P0001 , \wishbone_bd_ram_mem0_reg[251][5]/P0001 , \wishbone_bd_ram_mem0_reg[251][6]/P0001 , \wishbone_bd_ram_mem0_reg[251][7]/P0001 , \wishbone_bd_ram_mem0_reg[252][0]/P0001 , \wishbone_bd_ram_mem0_reg[252][1]/P0001 , \wishbone_bd_ram_mem0_reg[252][2]/P0001 , \wishbone_bd_ram_mem0_reg[252][3]/P0001 , \wishbone_bd_ram_mem0_reg[252][4]/P0001 , \wishbone_bd_ram_mem0_reg[252][5]/P0001 , \wishbone_bd_ram_mem0_reg[252][6]/P0001 , \wishbone_bd_ram_mem0_reg[252][7]/P0001 , \wishbone_bd_ram_mem0_reg[253][0]/P0001 , \wishbone_bd_ram_mem0_reg[253][1]/P0001 , \wishbone_bd_ram_mem0_reg[253][2]/P0001 , \wishbone_bd_ram_mem0_reg[253][3]/P0001 , \wishbone_bd_ram_mem0_reg[253][4]/P0001 , \wishbone_bd_ram_mem0_reg[253][5]/P0001 , \wishbone_bd_ram_mem0_reg[253][6]/P0001 , \wishbone_bd_ram_mem0_reg[253][7]/P0001 , \wishbone_bd_ram_mem0_reg[254][0]/P0001 , \wishbone_bd_ram_mem0_reg[254][1]/P0001 , \wishbone_bd_ram_mem0_reg[254][2]/P0001 , \wishbone_bd_ram_mem0_reg[254][3]/P0001 , \wishbone_bd_ram_mem0_reg[254][4]/P0001 , \wishbone_bd_ram_mem0_reg[254][5]/P0001 , \wishbone_bd_ram_mem0_reg[254][6]/P0001 , \wishbone_bd_ram_mem0_reg[254][7]/P0001 , \wishbone_bd_ram_mem0_reg[255][0]/P0001 , \wishbone_bd_ram_mem0_reg[255][1]/P0001 , \wishbone_bd_ram_mem0_reg[255][2]/P0001 , \wishbone_bd_ram_mem0_reg[255][3]/P0001 , \wishbone_bd_ram_mem0_reg[255][4]/P0001 , \wishbone_bd_ram_mem0_reg[255][5]/P0001 , \wishbone_bd_ram_mem0_reg[255][6]/P0001 , \wishbone_bd_ram_mem0_reg[255][7]/P0001 , \wishbone_bd_ram_mem0_reg[25][0]/P0001 , \wishbone_bd_ram_mem0_reg[25][1]/P0001 , \wishbone_bd_ram_mem0_reg[25][2]/P0001 , \wishbone_bd_ram_mem0_reg[25][3]/P0001 , \wishbone_bd_ram_mem0_reg[25][4]/P0001 , \wishbone_bd_ram_mem0_reg[25][5]/P0001 , \wishbone_bd_ram_mem0_reg[25][6]/P0001 , \wishbone_bd_ram_mem0_reg[25][7]/P0001 , \wishbone_bd_ram_mem0_reg[26][0]/P0001 , \wishbone_bd_ram_mem0_reg[26][1]/P0001 , \wishbone_bd_ram_mem0_reg[26][2]/P0001 , \wishbone_bd_ram_mem0_reg[26][3]/P0001 , \wishbone_bd_ram_mem0_reg[26][4]/P0001 , \wishbone_bd_ram_mem0_reg[26][5]/P0001 , \wishbone_bd_ram_mem0_reg[26][6]/P0001 , \wishbone_bd_ram_mem0_reg[26][7]/P0001 , \wishbone_bd_ram_mem0_reg[27][0]/P0001 , \wishbone_bd_ram_mem0_reg[27][1]/P0001 , \wishbone_bd_ram_mem0_reg[27][2]/P0001 , \wishbone_bd_ram_mem0_reg[27][3]/P0001 , \wishbone_bd_ram_mem0_reg[27][4]/P0001 , \wishbone_bd_ram_mem0_reg[27][5]/P0001 , \wishbone_bd_ram_mem0_reg[27][6]/P0001 , \wishbone_bd_ram_mem0_reg[27][7]/P0001 , \wishbone_bd_ram_mem0_reg[28][0]/P0001 , \wishbone_bd_ram_mem0_reg[28][1]/P0001 , \wishbone_bd_ram_mem0_reg[28][2]/P0001 , \wishbone_bd_ram_mem0_reg[28][3]/P0001 , \wishbone_bd_ram_mem0_reg[28][4]/P0001 , \wishbone_bd_ram_mem0_reg[28][5]/P0001 , \wishbone_bd_ram_mem0_reg[28][6]/P0001 , \wishbone_bd_ram_mem0_reg[28][7]/P0001 , \wishbone_bd_ram_mem0_reg[29][0]/P0001 , \wishbone_bd_ram_mem0_reg[29][1]/P0001 , \wishbone_bd_ram_mem0_reg[29][2]/P0001 , \wishbone_bd_ram_mem0_reg[29][3]/P0001 , \wishbone_bd_ram_mem0_reg[29][4]/P0001 , \wishbone_bd_ram_mem0_reg[29][5]/P0001 , \wishbone_bd_ram_mem0_reg[29][6]/P0001 , \wishbone_bd_ram_mem0_reg[29][7]/P0001 , \wishbone_bd_ram_mem0_reg[2][0]/P0001 , \wishbone_bd_ram_mem0_reg[2][1]/P0001 , \wishbone_bd_ram_mem0_reg[2][2]/P0001 , \wishbone_bd_ram_mem0_reg[2][3]/P0001 , \wishbone_bd_ram_mem0_reg[2][4]/P0001 , \wishbone_bd_ram_mem0_reg[2][5]/P0001 , \wishbone_bd_ram_mem0_reg[2][6]/P0001 , \wishbone_bd_ram_mem0_reg[2][7]/P0001 , \wishbone_bd_ram_mem0_reg[30][0]/P0001 , \wishbone_bd_ram_mem0_reg[30][1]/P0001 , \wishbone_bd_ram_mem0_reg[30][2]/P0001 , \wishbone_bd_ram_mem0_reg[30][3]/P0001 , \wishbone_bd_ram_mem0_reg[30][4]/P0001 , \wishbone_bd_ram_mem0_reg[30][5]/P0001 , \wishbone_bd_ram_mem0_reg[30][6]/P0001 , \wishbone_bd_ram_mem0_reg[30][7]/P0001 , \wishbone_bd_ram_mem0_reg[31][0]/P0001 , \wishbone_bd_ram_mem0_reg[31][1]/P0001 , \wishbone_bd_ram_mem0_reg[31][2]/P0001 , \wishbone_bd_ram_mem0_reg[31][3]/P0001 , \wishbone_bd_ram_mem0_reg[31][4]/P0001 , \wishbone_bd_ram_mem0_reg[31][5]/P0001 , \wishbone_bd_ram_mem0_reg[31][6]/P0001 , \wishbone_bd_ram_mem0_reg[31][7]/P0001 , \wishbone_bd_ram_mem0_reg[32][0]/P0001 , \wishbone_bd_ram_mem0_reg[32][1]/P0001 , \wishbone_bd_ram_mem0_reg[32][2]/P0001 , \wishbone_bd_ram_mem0_reg[32][3]/P0001 , \wishbone_bd_ram_mem0_reg[32][4]/P0001 , \wishbone_bd_ram_mem0_reg[32][5]/P0001 , \wishbone_bd_ram_mem0_reg[32][6]/P0001 , \wishbone_bd_ram_mem0_reg[32][7]/P0001 , \wishbone_bd_ram_mem0_reg[33][0]/P0001 , \wishbone_bd_ram_mem0_reg[33][1]/P0001 , \wishbone_bd_ram_mem0_reg[33][2]/P0001 , \wishbone_bd_ram_mem0_reg[33][3]/P0001 , \wishbone_bd_ram_mem0_reg[33][4]/P0001 , \wishbone_bd_ram_mem0_reg[33][5]/P0001 , \wishbone_bd_ram_mem0_reg[33][6]/P0001 , \wishbone_bd_ram_mem0_reg[33][7]/P0001 , \wishbone_bd_ram_mem0_reg[34][0]/P0001 , \wishbone_bd_ram_mem0_reg[34][1]/P0001 , \wishbone_bd_ram_mem0_reg[34][2]/P0001 , \wishbone_bd_ram_mem0_reg[34][3]/P0001 , \wishbone_bd_ram_mem0_reg[34][4]/P0001 , \wishbone_bd_ram_mem0_reg[34][5]/P0001 , \wishbone_bd_ram_mem0_reg[34][6]/P0001 , \wishbone_bd_ram_mem0_reg[34][7]/P0001 , \wishbone_bd_ram_mem0_reg[35][0]/P0001 , \wishbone_bd_ram_mem0_reg[35][1]/P0001 , \wishbone_bd_ram_mem0_reg[35][2]/P0001 , \wishbone_bd_ram_mem0_reg[35][3]/P0001 , \wishbone_bd_ram_mem0_reg[35][4]/P0001 , \wishbone_bd_ram_mem0_reg[35][5]/P0001 , \wishbone_bd_ram_mem0_reg[35][6]/P0001 , \wishbone_bd_ram_mem0_reg[35][7]/P0001 , \wishbone_bd_ram_mem0_reg[36][0]/P0001 , \wishbone_bd_ram_mem0_reg[36][1]/P0001 , \wishbone_bd_ram_mem0_reg[36][2]/P0001 , \wishbone_bd_ram_mem0_reg[36][3]/P0001 , \wishbone_bd_ram_mem0_reg[36][4]/P0001 , \wishbone_bd_ram_mem0_reg[36][5]/P0001 , \wishbone_bd_ram_mem0_reg[36][6]/P0001 , \wishbone_bd_ram_mem0_reg[36][7]/P0001 , \wishbone_bd_ram_mem0_reg[37][0]/P0001 , \wishbone_bd_ram_mem0_reg[37][1]/P0001 , \wishbone_bd_ram_mem0_reg[37][2]/P0001 , \wishbone_bd_ram_mem0_reg[37][3]/P0001 , \wishbone_bd_ram_mem0_reg[37][4]/P0001 , \wishbone_bd_ram_mem0_reg[37][5]/P0001 , \wishbone_bd_ram_mem0_reg[37][6]/P0001 , \wishbone_bd_ram_mem0_reg[37][7]/P0001 , \wishbone_bd_ram_mem0_reg[38][0]/P0001 , \wishbone_bd_ram_mem0_reg[38][1]/P0001 , \wishbone_bd_ram_mem0_reg[38][2]/P0001 , \wishbone_bd_ram_mem0_reg[38][3]/P0001 , \wishbone_bd_ram_mem0_reg[38][4]/P0001 , \wishbone_bd_ram_mem0_reg[38][5]/P0001 , \wishbone_bd_ram_mem0_reg[38][6]/P0001 , \wishbone_bd_ram_mem0_reg[38][7]/P0001 , \wishbone_bd_ram_mem0_reg[39][0]/P0001 , \wishbone_bd_ram_mem0_reg[39][1]/P0001 , \wishbone_bd_ram_mem0_reg[39][2]/P0001 , \wishbone_bd_ram_mem0_reg[39][3]/P0001 , \wishbone_bd_ram_mem0_reg[39][4]/P0001 , \wishbone_bd_ram_mem0_reg[39][5]/P0001 , \wishbone_bd_ram_mem0_reg[39][6]/P0001 , \wishbone_bd_ram_mem0_reg[39][7]/P0001 , \wishbone_bd_ram_mem0_reg[3][0]/P0001 , \wishbone_bd_ram_mem0_reg[3][1]/P0001 , \wishbone_bd_ram_mem0_reg[3][2]/P0001 , \wishbone_bd_ram_mem0_reg[3][3]/P0001 , \wishbone_bd_ram_mem0_reg[3][4]/P0001 , \wishbone_bd_ram_mem0_reg[3][5]/P0001 , \wishbone_bd_ram_mem0_reg[3][6]/P0001 , \wishbone_bd_ram_mem0_reg[3][7]/P0001 , \wishbone_bd_ram_mem0_reg[40][0]/P0001 , \wishbone_bd_ram_mem0_reg[40][1]/P0001 , \wishbone_bd_ram_mem0_reg[40][2]/P0001 , \wishbone_bd_ram_mem0_reg[40][3]/P0001 , \wishbone_bd_ram_mem0_reg[40][4]/P0001 , \wishbone_bd_ram_mem0_reg[40][5]/P0001 , \wishbone_bd_ram_mem0_reg[40][6]/P0001 , \wishbone_bd_ram_mem0_reg[40][7]/P0001 , \wishbone_bd_ram_mem0_reg[41][0]/P0001 , \wishbone_bd_ram_mem0_reg[41][1]/P0001 , \wishbone_bd_ram_mem0_reg[41][2]/P0001 , \wishbone_bd_ram_mem0_reg[41][3]/P0001 , \wishbone_bd_ram_mem0_reg[41][4]/P0001 , \wishbone_bd_ram_mem0_reg[41][5]/P0001 , \wishbone_bd_ram_mem0_reg[41][6]/P0001 , \wishbone_bd_ram_mem0_reg[41][7]/P0001 , \wishbone_bd_ram_mem0_reg[42][0]/P0001 , \wishbone_bd_ram_mem0_reg[42][1]/P0001 , \wishbone_bd_ram_mem0_reg[42][2]/P0001 , \wishbone_bd_ram_mem0_reg[42][3]/P0001 , \wishbone_bd_ram_mem0_reg[42][4]/P0001 , \wishbone_bd_ram_mem0_reg[42][5]/P0001 , \wishbone_bd_ram_mem0_reg[42][6]/P0001 , \wishbone_bd_ram_mem0_reg[42][7]/P0001 , \wishbone_bd_ram_mem0_reg[43][0]/P0001 , \wishbone_bd_ram_mem0_reg[43][1]/P0001 , \wishbone_bd_ram_mem0_reg[43][2]/P0001 , \wishbone_bd_ram_mem0_reg[43][3]/P0001 , \wishbone_bd_ram_mem0_reg[43][4]/P0001 , \wishbone_bd_ram_mem0_reg[43][5]/P0001 , \wishbone_bd_ram_mem0_reg[43][6]/P0001 , \wishbone_bd_ram_mem0_reg[43][7]/P0001 , \wishbone_bd_ram_mem0_reg[44][0]/P0001 , \wishbone_bd_ram_mem0_reg[44][1]/P0001 , \wishbone_bd_ram_mem0_reg[44][2]/P0001 , \wishbone_bd_ram_mem0_reg[44][3]/P0001 , \wishbone_bd_ram_mem0_reg[44][4]/P0001 , \wishbone_bd_ram_mem0_reg[44][5]/P0001 , \wishbone_bd_ram_mem0_reg[44][6]/P0001 , \wishbone_bd_ram_mem0_reg[44][7]/P0001 , \wishbone_bd_ram_mem0_reg[45][0]/P0001 , \wishbone_bd_ram_mem0_reg[45][1]/P0001 , \wishbone_bd_ram_mem0_reg[45][2]/P0001 , \wishbone_bd_ram_mem0_reg[45][3]/P0001 , \wishbone_bd_ram_mem0_reg[45][4]/P0001 , \wishbone_bd_ram_mem0_reg[45][5]/P0001 , \wishbone_bd_ram_mem0_reg[45][6]/P0001 , \wishbone_bd_ram_mem0_reg[45][7]/P0001 , \wishbone_bd_ram_mem0_reg[46][0]/P0001 , \wishbone_bd_ram_mem0_reg[46][1]/P0001 , \wishbone_bd_ram_mem0_reg[46][2]/P0001 , \wishbone_bd_ram_mem0_reg[46][3]/P0001 , \wishbone_bd_ram_mem0_reg[46][4]/P0001 , \wishbone_bd_ram_mem0_reg[46][5]/P0001 , \wishbone_bd_ram_mem0_reg[46][6]/P0001 , \wishbone_bd_ram_mem0_reg[46][7]/P0001 , \wishbone_bd_ram_mem0_reg[47][0]/P0001 , \wishbone_bd_ram_mem0_reg[47][1]/P0001 , \wishbone_bd_ram_mem0_reg[47][2]/P0001 , \wishbone_bd_ram_mem0_reg[47][3]/P0001 , \wishbone_bd_ram_mem0_reg[47][4]/P0001 , \wishbone_bd_ram_mem0_reg[47][5]/P0001 , \wishbone_bd_ram_mem0_reg[47][6]/P0001 , \wishbone_bd_ram_mem0_reg[47][7]/P0001 , \wishbone_bd_ram_mem0_reg[48][0]/P0001 , \wishbone_bd_ram_mem0_reg[48][1]/P0001 , \wishbone_bd_ram_mem0_reg[48][2]/P0001 , \wishbone_bd_ram_mem0_reg[48][3]/P0001 , \wishbone_bd_ram_mem0_reg[48][4]/P0001 , \wishbone_bd_ram_mem0_reg[48][5]/P0001 , \wishbone_bd_ram_mem0_reg[48][6]/P0001 , \wishbone_bd_ram_mem0_reg[48][7]/P0001 , \wishbone_bd_ram_mem0_reg[49][0]/P0001 , \wishbone_bd_ram_mem0_reg[49][1]/P0001 , \wishbone_bd_ram_mem0_reg[49][2]/P0001 , \wishbone_bd_ram_mem0_reg[49][3]/P0001 , \wishbone_bd_ram_mem0_reg[49][4]/P0001 , \wishbone_bd_ram_mem0_reg[49][5]/P0001 , \wishbone_bd_ram_mem0_reg[49][6]/P0001 , \wishbone_bd_ram_mem0_reg[49][7]/P0001 , \wishbone_bd_ram_mem0_reg[4][0]/P0001 , \wishbone_bd_ram_mem0_reg[4][1]/P0001 , \wishbone_bd_ram_mem0_reg[4][2]/P0001 , \wishbone_bd_ram_mem0_reg[4][3]/P0001 , \wishbone_bd_ram_mem0_reg[4][4]/P0001 , \wishbone_bd_ram_mem0_reg[4][5]/P0001 , \wishbone_bd_ram_mem0_reg[4][6]/P0001 , \wishbone_bd_ram_mem0_reg[4][7]/P0001 , \wishbone_bd_ram_mem0_reg[50][0]/P0001 , \wishbone_bd_ram_mem0_reg[50][1]/P0001 , \wishbone_bd_ram_mem0_reg[50][2]/P0001 , \wishbone_bd_ram_mem0_reg[50][3]/P0001 , \wishbone_bd_ram_mem0_reg[50][4]/P0001 , \wishbone_bd_ram_mem0_reg[50][5]/P0001 , \wishbone_bd_ram_mem0_reg[50][6]/P0001 , \wishbone_bd_ram_mem0_reg[50][7]/P0001 , \wishbone_bd_ram_mem0_reg[51][0]/P0001 , \wishbone_bd_ram_mem0_reg[51][1]/P0001 , \wishbone_bd_ram_mem0_reg[51][2]/P0001 , \wishbone_bd_ram_mem0_reg[51][3]/P0001 , \wishbone_bd_ram_mem0_reg[51][4]/P0001 , \wishbone_bd_ram_mem0_reg[51][5]/P0001 , \wishbone_bd_ram_mem0_reg[51][6]/P0001 , \wishbone_bd_ram_mem0_reg[51][7]/P0001 , \wishbone_bd_ram_mem0_reg[52][0]/P0001 , \wishbone_bd_ram_mem0_reg[52][1]/P0001 , \wishbone_bd_ram_mem0_reg[52][2]/P0001 , \wishbone_bd_ram_mem0_reg[52][3]/P0001 , \wishbone_bd_ram_mem0_reg[52][4]/P0001 , \wishbone_bd_ram_mem0_reg[52][5]/P0001 , \wishbone_bd_ram_mem0_reg[52][6]/P0001 , \wishbone_bd_ram_mem0_reg[52][7]/P0001 , \wishbone_bd_ram_mem0_reg[53][0]/P0001 , \wishbone_bd_ram_mem0_reg[53][1]/P0001 , \wishbone_bd_ram_mem0_reg[53][2]/P0001 , \wishbone_bd_ram_mem0_reg[53][3]/P0001 , \wishbone_bd_ram_mem0_reg[53][4]/P0001 , \wishbone_bd_ram_mem0_reg[53][5]/P0001 , \wishbone_bd_ram_mem0_reg[53][6]/P0001 , \wishbone_bd_ram_mem0_reg[53][7]/P0001 , \wishbone_bd_ram_mem0_reg[54][0]/P0001 , \wishbone_bd_ram_mem0_reg[54][1]/P0001 , \wishbone_bd_ram_mem0_reg[54][2]/P0001 , \wishbone_bd_ram_mem0_reg[54][3]/P0001 , \wishbone_bd_ram_mem0_reg[54][4]/P0001 , \wishbone_bd_ram_mem0_reg[54][5]/P0001 , \wishbone_bd_ram_mem0_reg[54][6]/P0001 , \wishbone_bd_ram_mem0_reg[54][7]/P0001 , \wishbone_bd_ram_mem0_reg[55][0]/P0001 , \wishbone_bd_ram_mem0_reg[55][1]/P0001 , \wishbone_bd_ram_mem0_reg[55][2]/P0001 , \wishbone_bd_ram_mem0_reg[55][3]/P0001 , \wishbone_bd_ram_mem0_reg[55][4]/P0001 , \wishbone_bd_ram_mem0_reg[55][5]/P0001 , \wishbone_bd_ram_mem0_reg[55][6]/P0001 , \wishbone_bd_ram_mem0_reg[55][7]/P0001 , \wishbone_bd_ram_mem0_reg[56][0]/P0001 , \wishbone_bd_ram_mem0_reg[56][1]/P0001 , \wishbone_bd_ram_mem0_reg[56][2]/P0001 , \wishbone_bd_ram_mem0_reg[56][3]/P0001 , \wishbone_bd_ram_mem0_reg[56][4]/P0001 , \wishbone_bd_ram_mem0_reg[56][5]/P0001 , \wishbone_bd_ram_mem0_reg[56][6]/P0001 , \wishbone_bd_ram_mem0_reg[56][7]/P0001 , \wishbone_bd_ram_mem0_reg[57][0]/P0001 , \wishbone_bd_ram_mem0_reg[57][1]/P0001 , \wishbone_bd_ram_mem0_reg[57][2]/P0001 , \wishbone_bd_ram_mem0_reg[57][3]/P0001 , \wishbone_bd_ram_mem0_reg[57][4]/P0001 , \wishbone_bd_ram_mem0_reg[57][5]/P0001 , \wishbone_bd_ram_mem0_reg[57][6]/P0001 , \wishbone_bd_ram_mem0_reg[57][7]/P0001 , \wishbone_bd_ram_mem0_reg[58][0]/P0001 , \wishbone_bd_ram_mem0_reg[58][1]/P0001 , \wishbone_bd_ram_mem0_reg[58][2]/P0001 , \wishbone_bd_ram_mem0_reg[58][3]/P0001 , \wishbone_bd_ram_mem0_reg[58][4]/P0001 , \wishbone_bd_ram_mem0_reg[58][5]/P0001 , \wishbone_bd_ram_mem0_reg[58][6]/P0001 , \wishbone_bd_ram_mem0_reg[58][7]/P0001 , \wishbone_bd_ram_mem0_reg[59][0]/P0001 , \wishbone_bd_ram_mem0_reg[59][1]/P0001 , \wishbone_bd_ram_mem0_reg[59][2]/P0001 , \wishbone_bd_ram_mem0_reg[59][3]/P0001 , \wishbone_bd_ram_mem0_reg[59][4]/P0001 , \wishbone_bd_ram_mem0_reg[59][5]/P0001 , \wishbone_bd_ram_mem0_reg[59][6]/P0001 , \wishbone_bd_ram_mem0_reg[59][7]/P0001 , \wishbone_bd_ram_mem0_reg[5][0]/P0001 , \wishbone_bd_ram_mem0_reg[5][1]/P0001 , \wishbone_bd_ram_mem0_reg[5][2]/P0001 , \wishbone_bd_ram_mem0_reg[5][3]/P0001 , \wishbone_bd_ram_mem0_reg[5][4]/P0001 , \wishbone_bd_ram_mem0_reg[5][5]/P0001 , \wishbone_bd_ram_mem0_reg[5][6]/P0001 , \wishbone_bd_ram_mem0_reg[5][7]/P0001 , \wishbone_bd_ram_mem0_reg[60][0]/P0001 , \wishbone_bd_ram_mem0_reg[60][1]/P0001 , \wishbone_bd_ram_mem0_reg[60][2]/P0001 , \wishbone_bd_ram_mem0_reg[60][3]/P0001 , \wishbone_bd_ram_mem0_reg[60][4]/P0001 , \wishbone_bd_ram_mem0_reg[60][5]/P0001 , \wishbone_bd_ram_mem0_reg[60][6]/P0001 , \wishbone_bd_ram_mem0_reg[60][7]/P0001 , \wishbone_bd_ram_mem0_reg[61][0]/P0001 , \wishbone_bd_ram_mem0_reg[61][1]/P0001 , \wishbone_bd_ram_mem0_reg[61][2]/P0001 , \wishbone_bd_ram_mem0_reg[61][3]/P0001 , \wishbone_bd_ram_mem0_reg[61][4]/P0001 , \wishbone_bd_ram_mem0_reg[61][5]/P0001 , \wishbone_bd_ram_mem0_reg[61][6]/P0001 , \wishbone_bd_ram_mem0_reg[61][7]/P0001 , \wishbone_bd_ram_mem0_reg[62][0]/P0001 , \wishbone_bd_ram_mem0_reg[62][1]/P0001 , \wishbone_bd_ram_mem0_reg[62][2]/P0001 , \wishbone_bd_ram_mem0_reg[62][3]/P0001 , \wishbone_bd_ram_mem0_reg[62][4]/P0001 , \wishbone_bd_ram_mem0_reg[62][5]/P0001 , \wishbone_bd_ram_mem0_reg[62][6]/P0001 , \wishbone_bd_ram_mem0_reg[62][7]/P0001 , \wishbone_bd_ram_mem0_reg[63][0]/P0001 , \wishbone_bd_ram_mem0_reg[63][1]/P0001 , \wishbone_bd_ram_mem0_reg[63][2]/P0001 , \wishbone_bd_ram_mem0_reg[63][3]/P0001 , \wishbone_bd_ram_mem0_reg[63][4]/P0001 , \wishbone_bd_ram_mem0_reg[63][5]/P0001 , \wishbone_bd_ram_mem0_reg[63][6]/P0001 , \wishbone_bd_ram_mem0_reg[63][7]/P0001 , \wishbone_bd_ram_mem0_reg[64][0]/P0001 , \wishbone_bd_ram_mem0_reg[64][1]/P0001 , \wishbone_bd_ram_mem0_reg[64][2]/P0001 , \wishbone_bd_ram_mem0_reg[64][3]/P0001 , \wishbone_bd_ram_mem0_reg[64][4]/P0001 , \wishbone_bd_ram_mem0_reg[64][5]/P0001 , \wishbone_bd_ram_mem0_reg[64][6]/P0001 , \wishbone_bd_ram_mem0_reg[64][7]/P0001 , \wishbone_bd_ram_mem0_reg[65][0]/P0001 , \wishbone_bd_ram_mem0_reg[65][1]/P0001 , \wishbone_bd_ram_mem0_reg[65][2]/P0001 , \wishbone_bd_ram_mem0_reg[65][3]/P0001 , \wishbone_bd_ram_mem0_reg[65][4]/P0001 , \wishbone_bd_ram_mem0_reg[65][5]/P0001 , \wishbone_bd_ram_mem0_reg[65][6]/P0001 , \wishbone_bd_ram_mem0_reg[65][7]/P0001 , \wishbone_bd_ram_mem0_reg[66][0]/P0001 , \wishbone_bd_ram_mem0_reg[66][1]/P0001 , \wishbone_bd_ram_mem0_reg[66][2]/P0001 , \wishbone_bd_ram_mem0_reg[66][3]/P0001 , \wishbone_bd_ram_mem0_reg[66][4]/P0001 , \wishbone_bd_ram_mem0_reg[66][5]/P0001 , \wishbone_bd_ram_mem0_reg[66][6]/P0001 , \wishbone_bd_ram_mem0_reg[66][7]/P0001 , \wishbone_bd_ram_mem0_reg[67][0]/P0001 , \wishbone_bd_ram_mem0_reg[67][1]/P0001 , \wishbone_bd_ram_mem0_reg[67][2]/P0001 , \wishbone_bd_ram_mem0_reg[67][3]/P0001 , \wishbone_bd_ram_mem0_reg[67][4]/P0001 , \wishbone_bd_ram_mem0_reg[67][5]/P0001 , \wishbone_bd_ram_mem0_reg[67][6]/P0001 , \wishbone_bd_ram_mem0_reg[67][7]/P0001 , \wishbone_bd_ram_mem0_reg[68][0]/P0001 , \wishbone_bd_ram_mem0_reg[68][1]/P0001 , \wishbone_bd_ram_mem0_reg[68][2]/P0001 , \wishbone_bd_ram_mem0_reg[68][3]/P0001 , \wishbone_bd_ram_mem0_reg[68][4]/P0001 , \wishbone_bd_ram_mem0_reg[68][5]/P0001 , \wishbone_bd_ram_mem0_reg[68][6]/P0001 , \wishbone_bd_ram_mem0_reg[68][7]/P0001 , \wishbone_bd_ram_mem0_reg[69][0]/P0001 , \wishbone_bd_ram_mem0_reg[69][1]/P0001 , \wishbone_bd_ram_mem0_reg[69][2]/P0001 , \wishbone_bd_ram_mem0_reg[69][3]/P0001 , \wishbone_bd_ram_mem0_reg[69][4]/P0001 , \wishbone_bd_ram_mem0_reg[69][5]/P0001 , \wishbone_bd_ram_mem0_reg[69][6]/P0001 , \wishbone_bd_ram_mem0_reg[69][7]/P0001 , \wishbone_bd_ram_mem0_reg[6][0]/P0001 , \wishbone_bd_ram_mem0_reg[6][1]/P0001 , \wishbone_bd_ram_mem0_reg[6][2]/P0001 , \wishbone_bd_ram_mem0_reg[6][3]/P0001 , \wishbone_bd_ram_mem0_reg[6][4]/P0001 , \wishbone_bd_ram_mem0_reg[6][5]/P0001 , \wishbone_bd_ram_mem0_reg[6][6]/P0001 , \wishbone_bd_ram_mem0_reg[6][7]/P0001 , \wishbone_bd_ram_mem0_reg[70][0]/P0001 , \wishbone_bd_ram_mem0_reg[70][1]/P0001 , \wishbone_bd_ram_mem0_reg[70][2]/P0001 , \wishbone_bd_ram_mem0_reg[70][3]/P0001 , \wishbone_bd_ram_mem0_reg[70][4]/P0001 , \wishbone_bd_ram_mem0_reg[70][5]/P0001 , \wishbone_bd_ram_mem0_reg[70][6]/P0001 , \wishbone_bd_ram_mem0_reg[70][7]/P0001 , \wishbone_bd_ram_mem0_reg[71][0]/P0001 , \wishbone_bd_ram_mem0_reg[71][1]/P0001 , \wishbone_bd_ram_mem0_reg[71][2]/P0001 , \wishbone_bd_ram_mem0_reg[71][3]/P0001 , \wishbone_bd_ram_mem0_reg[71][4]/P0001 , \wishbone_bd_ram_mem0_reg[71][5]/P0001 , \wishbone_bd_ram_mem0_reg[71][6]/P0001 , \wishbone_bd_ram_mem0_reg[71][7]/P0001 , \wishbone_bd_ram_mem0_reg[72][0]/P0001 , \wishbone_bd_ram_mem0_reg[72][1]/P0001 , \wishbone_bd_ram_mem0_reg[72][2]/P0001 , \wishbone_bd_ram_mem0_reg[72][3]/P0001 , \wishbone_bd_ram_mem0_reg[72][4]/P0001 , \wishbone_bd_ram_mem0_reg[72][5]/P0001 , \wishbone_bd_ram_mem0_reg[72][6]/P0001 , \wishbone_bd_ram_mem0_reg[72][7]/P0001 , \wishbone_bd_ram_mem0_reg[73][0]/P0001 , \wishbone_bd_ram_mem0_reg[73][1]/P0001 , \wishbone_bd_ram_mem0_reg[73][2]/P0001 , \wishbone_bd_ram_mem0_reg[73][3]/P0001 , \wishbone_bd_ram_mem0_reg[73][4]/P0001 , \wishbone_bd_ram_mem0_reg[73][5]/P0001 , \wishbone_bd_ram_mem0_reg[73][6]/P0001 , \wishbone_bd_ram_mem0_reg[73][7]/P0001 , \wishbone_bd_ram_mem0_reg[74][0]/P0001 , \wishbone_bd_ram_mem0_reg[74][1]/P0001 , \wishbone_bd_ram_mem0_reg[74][2]/P0001 , \wishbone_bd_ram_mem0_reg[74][3]/P0001 , \wishbone_bd_ram_mem0_reg[74][4]/P0001 , \wishbone_bd_ram_mem0_reg[74][5]/P0001 , \wishbone_bd_ram_mem0_reg[74][6]/P0001 , \wishbone_bd_ram_mem0_reg[74][7]/P0001 , \wishbone_bd_ram_mem0_reg[75][0]/P0001 , \wishbone_bd_ram_mem0_reg[75][1]/P0001 , \wishbone_bd_ram_mem0_reg[75][2]/P0001 , \wishbone_bd_ram_mem0_reg[75][3]/P0001 , \wishbone_bd_ram_mem0_reg[75][4]/P0001 , \wishbone_bd_ram_mem0_reg[75][5]/P0001 , \wishbone_bd_ram_mem0_reg[75][6]/P0001 , \wishbone_bd_ram_mem0_reg[75][7]/P0001 , \wishbone_bd_ram_mem0_reg[76][0]/P0001 , \wishbone_bd_ram_mem0_reg[76][1]/P0001 , \wishbone_bd_ram_mem0_reg[76][2]/P0001 , \wishbone_bd_ram_mem0_reg[76][3]/P0001 , \wishbone_bd_ram_mem0_reg[76][4]/P0001 , \wishbone_bd_ram_mem0_reg[76][5]/P0001 , \wishbone_bd_ram_mem0_reg[76][6]/P0001 , \wishbone_bd_ram_mem0_reg[76][7]/P0001 , \wishbone_bd_ram_mem0_reg[77][0]/P0001 , \wishbone_bd_ram_mem0_reg[77][1]/P0001 , \wishbone_bd_ram_mem0_reg[77][2]/P0001 , \wishbone_bd_ram_mem0_reg[77][3]/P0001 , \wishbone_bd_ram_mem0_reg[77][4]/P0001 , \wishbone_bd_ram_mem0_reg[77][5]/P0001 , \wishbone_bd_ram_mem0_reg[77][6]/P0001 , \wishbone_bd_ram_mem0_reg[77][7]/P0001 , \wishbone_bd_ram_mem0_reg[78][0]/P0001 , \wishbone_bd_ram_mem0_reg[78][1]/P0001 , \wishbone_bd_ram_mem0_reg[78][2]/P0001 , \wishbone_bd_ram_mem0_reg[78][3]/P0001 , \wishbone_bd_ram_mem0_reg[78][4]/P0001 , \wishbone_bd_ram_mem0_reg[78][5]/P0001 , \wishbone_bd_ram_mem0_reg[78][6]/P0001 , \wishbone_bd_ram_mem0_reg[78][7]/P0001 , \wishbone_bd_ram_mem0_reg[79][0]/P0001 , \wishbone_bd_ram_mem0_reg[79][1]/P0001 , \wishbone_bd_ram_mem0_reg[79][2]/P0001 , \wishbone_bd_ram_mem0_reg[79][3]/P0001 , \wishbone_bd_ram_mem0_reg[79][4]/P0001 , \wishbone_bd_ram_mem0_reg[79][5]/P0001 , \wishbone_bd_ram_mem0_reg[79][6]/P0001 , \wishbone_bd_ram_mem0_reg[79][7]/P0001 , \wishbone_bd_ram_mem0_reg[7][0]/P0001 , \wishbone_bd_ram_mem0_reg[7][1]/P0001 , \wishbone_bd_ram_mem0_reg[7][2]/P0001 , \wishbone_bd_ram_mem0_reg[7][3]/P0001 , \wishbone_bd_ram_mem0_reg[7][4]/P0001 , \wishbone_bd_ram_mem0_reg[7][5]/P0001 , \wishbone_bd_ram_mem0_reg[7][6]/P0001 , \wishbone_bd_ram_mem0_reg[7][7]/P0001 , \wishbone_bd_ram_mem0_reg[80][0]/P0001 , \wishbone_bd_ram_mem0_reg[80][1]/P0001 , \wishbone_bd_ram_mem0_reg[80][2]/P0001 , \wishbone_bd_ram_mem0_reg[80][3]/P0001 , \wishbone_bd_ram_mem0_reg[80][4]/P0001 , \wishbone_bd_ram_mem0_reg[80][5]/P0001 , \wishbone_bd_ram_mem0_reg[80][6]/P0001 , \wishbone_bd_ram_mem0_reg[80][7]/P0001 , \wishbone_bd_ram_mem0_reg[81][0]/P0001 , \wishbone_bd_ram_mem0_reg[81][1]/P0001 , \wishbone_bd_ram_mem0_reg[81][2]/P0001 , \wishbone_bd_ram_mem0_reg[81][3]/P0001 , \wishbone_bd_ram_mem0_reg[81][4]/P0001 , \wishbone_bd_ram_mem0_reg[81][5]/P0001 , \wishbone_bd_ram_mem0_reg[81][6]/P0001 , \wishbone_bd_ram_mem0_reg[81][7]/P0001 , \wishbone_bd_ram_mem0_reg[82][0]/P0001 , \wishbone_bd_ram_mem0_reg[82][1]/P0001 , \wishbone_bd_ram_mem0_reg[82][2]/P0001 , \wishbone_bd_ram_mem0_reg[82][3]/P0001 , \wishbone_bd_ram_mem0_reg[82][4]/P0001 , \wishbone_bd_ram_mem0_reg[82][5]/P0001 , \wishbone_bd_ram_mem0_reg[82][6]/P0001 , \wishbone_bd_ram_mem0_reg[82][7]/P0001 , \wishbone_bd_ram_mem0_reg[83][0]/P0001 , \wishbone_bd_ram_mem0_reg[83][1]/P0001 , \wishbone_bd_ram_mem0_reg[83][2]/P0001 , \wishbone_bd_ram_mem0_reg[83][3]/P0001 , \wishbone_bd_ram_mem0_reg[83][4]/P0001 , \wishbone_bd_ram_mem0_reg[83][5]/P0001 , \wishbone_bd_ram_mem0_reg[83][6]/P0001 , \wishbone_bd_ram_mem0_reg[83][7]/P0001 , \wishbone_bd_ram_mem0_reg[84][0]/P0001 , \wishbone_bd_ram_mem0_reg[84][1]/P0001 , \wishbone_bd_ram_mem0_reg[84][2]/P0001 , \wishbone_bd_ram_mem0_reg[84][3]/P0001 , \wishbone_bd_ram_mem0_reg[84][4]/P0001 , \wishbone_bd_ram_mem0_reg[84][5]/P0001 , \wishbone_bd_ram_mem0_reg[84][6]/P0001 , \wishbone_bd_ram_mem0_reg[84][7]/P0001 , \wishbone_bd_ram_mem0_reg[85][0]/P0001 , \wishbone_bd_ram_mem0_reg[85][1]/P0001 , \wishbone_bd_ram_mem0_reg[85][2]/P0001 , \wishbone_bd_ram_mem0_reg[85][3]/P0001 , \wishbone_bd_ram_mem0_reg[85][4]/P0001 , \wishbone_bd_ram_mem0_reg[85][5]/P0001 , \wishbone_bd_ram_mem0_reg[85][6]/P0001 , \wishbone_bd_ram_mem0_reg[85][7]/P0001 , \wishbone_bd_ram_mem0_reg[86][0]/P0001 , \wishbone_bd_ram_mem0_reg[86][1]/P0001 , \wishbone_bd_ram_mem0_reg[86][2]/P0001 , \wishbone_bd_ram_mem0_reg[86][3]/P0001 , \wishbone_bd_ram_mem0_reg[86][4]/P0001 , \wishbone_bd_ram_mem0_reg[86][5]/P0001 , \wishbone_bd_ram_mem0_reg[86][6]/P0001 , \wishbone_bd_ram_mem0_reg[86][7]/P0001 , \wishbone_bd_ram_mem0_reg[87][0]/P0001 , \wishbone_bd_ram_mem0_reg[87][1]/P0001 , \wishbone_bd_ram_mem0_reg[87][2]/P0001 , \wishbone_bd_ram_mem0_reg[87][3]/P0001 , \wishbone_bd_ram_mem0_reg[87][4]/P0001 , \wishbone_bd_ram_mem0_reg[87][5]/P0001 , \wishbone_bd_ram_mem0_reg[87][6]/P0001 , \wishbone_bd_ram_mem0_reg[87][7]/P0001 , \wishbone_bd_ram_mem0_reg[88][0]/P0001 , \wishbone_bd_ram_mem0_reg[88][1]/P0001 , \wishbone_bd_ram_mem0_reg[88][2]/P0001 , \wishbone_bd_ram_mem0_reg[88][3]/P0001 , \wishbone_bd_ram_mem0_reg[88][4]/P0001 , \wishbone_bd_ram_mem0_reg[88][5]/P0001 , \wishbone_bd_ram_mem0_reg[88][6]/P0001 , \wishbone_bd_ram_mem0_reg[88][7]/P0001 , \wishbone_bd_ram_mem0_reg[89][0]/P0001 , \wishbone_bd_ram_mem0_reg[89][1]/P0001 , \wishbone_bd_ram_mem0_reg[89][2]/P0001 , \wishbone_bd_ram_mem0_reg[89][3]/P0001 , \wishbone_bd_ram_mem0_reg[89][4]/P0001 , \wishbone_bd_ram_mem0_reg[89][5]/P0001 , \wishbone_bd_ram_mem0_reg[89][6]/P0001 , \wishbone_bd_ram_mem0_reg[89][7]/P0001 , \wishbone_bd_ram_mem0_reg[8][0]/P0001 , \wishbone_bd_ram_mem0_reg[8][1]/P0001 , \wishbone_bd_ram_mem0_reg[8][2]/P0001 , \wishbone_bd_ram_mem0_reg[8][3]/P0001 , \wishbone_bd_ram_mem0_reg[8][4]/P0001 , \wishbone_bd_ram_mem0_reg[8][5]/P0001 , \wishbone_bd_ram_mem0_reg[8][6]/P0001 , \wishbone_bd_ram_mem0_reg[8][7]/P0001 , \wishbone_bd_ram_mem0_reg[90][0]/P0001 , \wishbone_bd_ram_mem0_reg[90][1]/P0001 , \wishbone_bd_ram_mem0_reg[90][2]/P0001 , \wishbone_bd_ram_mem0_reg[90][3]/P0001 , \wishbone_bd_ram_mem0_reg[90][4]/P0001 , \wishbone_bd_ram_mem0_reg[90][5]/P0001 , \wishbone_bd_ram_mem0_reg[90][6]/P0001 , \wishbone_bd_ram_mem0_reg[90][7]/P0001 , \wishbone_bd_ram_mem0_reg[91][0]/P0001 , \wishbone_bd_ram_mem0_reg[91][1]/P0001 , \wishbone_bd_ram_mem0_reg[91][2]/P0001 , \wishbone_bd_ram_mem0_reg[91][3]/P0001 , \wishbone_bd_ram_mem0_reg[91][4]/P0001 , \wishbone_bd_ram_mem0_reg[91][5]/P0001 , \wishbone_bd_ram_mem0_reg[91][6]/P0001 , \wishbone_bd_ram_mem0_reg[91][7]/P0001 , \wishbone_bd_ram_mem0_reg[92][0]/P0001 , \wishbone_bd_ram_mem0_reg[92][1]/P0001 , \wishbone_bd_ram_mem0_reg[92][2]/P0001 , \wishbone_bd_ram_mem0_reg[92][3]/P0001 , \wishbone_bd_ram_mem0_reg[92][4]/P0001 , \wishbone_bd_ram_mem0_reg[92][5]/P0001 , \wishbone_bd_ram_mem0_reg[92][6]/P0001 , \wishbone_bd_ram_mem0_reg[92][7]/P0001 , \wishbone_bd_ram_mem0_reg[93][0]/P0001 , \wishbone_bd_ram_mem0_reg[93][1]/P0001 , \wishbone_bd_ram_mem0_reg[93][2]/P0001 , \wishbone_bd_ram_mem0_reg[93][3]/P0001 , \wishbone_bd_ram_mem0_reg[93][4]/P0001 , \wishbone_bd_ram_mem0_reg[93][5]/P0001 , \wishbone_bd_ram_mem0_reg[93][6]/P0001 , \wishbone_bd_ram_mem0_reg[93][7]/P0001 , \wishbone_bd_ram_mem0_reg[94][0]/P0001 , \wishbone_bd_ram_mem0_reg[94][1]/P0001 , \wishbone_bd_ram_mem0_reg[94][2]/P0001 , \wishbone_bd_ram_mem0_reg[94][3]/P0001 , \wishbone_bd_ram_mem0_reg[94][4]/P0001 , \wishbone_bd_ram_mem0_reg[94][5]/P0001 , \wishbone_bd_ram_mem0_reg[94][6]/P0001 , \wishbone_bd_ram_mem0_reg[94][7]/P0001 , \wishbone_bd_ram_mem0_reg[95][0]/P0001 , \wishbone_bd_ram_mem0_reg[95][1]/P0001 , \wishbone_bd_ram_mem0_reg[95][2]/P0001 , \wishbone_bd_ram_mem0_reg[95][3]/P0001 , \wishbone_bd_ram_mem0_reg[95][4]/P0001 , \wishbone_bd_ram_mem0_reg[95][5]/P0001 , \wishbone_bd_ram_mem0_reg[95][6]/P0001 , \wishbone_bd_ram_mem0_reg[95][7]/P0001 , \wishbone_bd_ram_mem0_reg[96][0]/P0001 , \wishbone_bd_ram_mem0_reg[96][1]/P0001 , \wishbone_bd_ram_mem0_reg[96][2]/P0001 , \wishbone_bd_ram_mem0_reg[96][3]/P0001 , \wishbone_bd_ram_mem0_reg[96][4]/P0001 , \wishbone_bd_ram_mem0_reg[96][5]/P0001 , \wishbone_bd_ram_mem0_reg[96][6]/P0001 , \wishbone_bd_ram_mem0_reg[96][7]/P0001 , \wishbone_bd_ram_mem0_reg[97][0]/P0001 , \wishbone_bd_ram_mem0_reg[97][1]/P0001 , \wishbone_bd_ram_mem0_reg[97][2]/P0001 , \wishbone_bd_ram_mem0_reg[97][3]/P0001 , \wishbone_bd_ram_mem0_reg[97][4]/P0001 , \wishbone_bd_ram_mem0_reg[97][5]/P0001 , \wishbone_bd_ram_mem0_reg[97][6]/P0001 , \wishbone_bd_ram_mem0_reg[97][7]/P0001 , \wishbone_bd_ram_mem0_reg[98][0]/P0001 , \wishbone_bd_ram_mem0_reg[98][1]/P0001 , \wishbone_bd_ram_mem0_reg[98][2]/P0001 , \wishbone_bd_ram_mem0_reg[98][3]/P0001 , \wishbone_bd_ram_mem0_reg[98][4]/P0001 , \wishbone_bd_ram_mem0_reg[98][5]/P0001 , \wishbone_bd_ram_mem0_reg[98][6]/P0001 , \wishbone_bd_ram_mem0_reg[98][7]/P0001 , \wishbone_bd_ram_mem0_reg[99][0]/P0001 , \wishbone_bd_ram_mem0_reg[99][1]/P0001 , \wishbone_bd_ram_mem0_reg[99][2]/P0001 , \wishbone_bd_ram_mem0_reg[99][3]/P0001 , \wishbone_bd_ram_mem0_reg[99][4]/P0001 , \wishbone_bd_ram_mem0_reg[99][5]/P0001 , \wishbone_bd_ram_mem0_reg[99][6]/P0001 , \wishbone_bd_ram_mem0_reg[99][7]/P0001 , \wishbone_bd_ram_mem0_reg[9][0]/P0001 , \wishbone_bd_ram_mem0_reg[9][1]/P0001 , \wishbone_bd_ram_mem0_reg[9][2]/P0001 , \wishbone_bd_ram_mem0_reg[9][3]/P0001 , \wishbone_bd_ram_mem0_reg[9][4]/P0001 , \wishbone_bd_ram_mem0_reg[9][5]/P0001 , \wishbone_bd_ram_mem0_reg[9][6]/P0001 , \wishbone_bd_ram_mem0_reg[9][7]/P0001 , \wishbone_bd_ram_mem1_reg[0][10]/P0001 , \wishbone_bd_ram_mem1_reg[0][11]/P0001 , \wishbone_bd_ram_mem1_reg[0][12]/P0001 , \wishbone_bd_ram_mem1_reg[0][13]/P0001 , \wishbone_bd_ram_mem1_reg[0][14]/P0001 , \wishbone_bd_ram_mem1_reg[0][15]/P0001 , \wishbone_bd_ram_mem1_reg[0][8]/P0001 , \wishbone_bd_ram_mem1_reg[0][9]/P0001 , \wishbone_bd_ram_mem1_reg[100][10]/P0001 , \wishbone_bd_ram_mem1_reg[100][11]/P0001 , \wishbone_bd_ram_mem1_reg[100][12]/P0001 , \wishbone_bd_ram_mem1_reg[100][13]/P0001 , \wishbone_bd_ram_mem1_reg[100][14]/P0001 , \wishbone_bd_ram_mem1_reg[100][15]/P0001 , \wishbone_bd_ram_mem1_reg[100][8]/P0001 , \wishbone_bd_ram_mem1_reg[100][9]/P0001 , \wishbone_bd_ram_mem1_reg[101][10]/P0001 , \wishbone_bd_ram_mem1_reg[101][11]/P0001 , \wishbone_bd_ram_mem1_reg[101][12]/P0001 , \wishbone_bd_ram_mem1_reg[101][13]/P0001 , \wishbone_bd_ram_mem1_reg[101][14]/P0001 , \wishbone_bd_ram_mem1_reg[101][15]/P0001 , \wishbone_bd_ram_mem1_reg[101][8]/P0001 , \wishbone_bd_ram_mem1_reg[101][9]/P0001 , \wishbone_bd_ram_mem1_reg[102][10]/P0001 , \wishbone_bd_ram_mem1_reg[102][11]/P0001 , \wishbone_bd_ram_mem1_reg[102][12]/P0001 , \wishbone_bd_ram_mem1_reg[102][13]/P0001 , \wishbone_bd_ram_mem1_reg[102][14]/P0001 , \wishbone_bd_ram_mem1_reg[102][15]/P0001 , \wishbone_bd_ram_mem1_reg[102][8]/P0001 , \wishbone_bd_ram_mem1_reg[102][9]/P0001 , \wishbone_bd_ram_mem1_reg[103][10]/P0001 , \wishbone_bd_ram_mem1_reg[103][11]/P0001 , \wishbone_bd_ram_mem1_reg[103][12]/P0001 , \wishbone_bd_ram_mem1_reg[103][13]/P0001 , \wishbone_bd_ram_mem1_reg[103][14]/P0001 , \wishbone_bd_ram_mem1_reg[103][15]/P0001 , \wishbone_bd_ram_mem1_reg[103][8]/P0001 , \wishbone_bd_ram_mem1_reg[103][9]/P0001 , \wishbone_bd_ram_mem1_reg[104][10]/P0001 , \wishbone_bd_ram_mem1_reg[104][11]/P0001 , \wishbone_bd_ram_mem1_reg[104][12]/P0001 , \wishbone_bd_ram_mem1_reg[104][13]/P0001 , \wishbone_bd_ram_mem1_reg[104][14]/P0001 , \wishbone_bd_ram_mem1_reg[104][15]/P0001 , \wishbone_bd_ram_mem1_reg[104][8]/P0001 , \wishbone_bd_ram_mem1_reg[104][9]/P0001 , \wishbone_bd_ram_mem1_reg[105][10]/P0001 , \wishbone_bd_ram_mem1_reg[105][11]/P0001 , \wishbone_bd_ram_mem1_reg[105][12]/P0001 , \wishbone_bd_ram_mem1_reg[105][13]/P0001 , \wishbone_bd_ram_mem1_reg[105][14]/P0001 , \wishbone_bd_ram_mem1_reg[105][15]/P0001 , \wishbone_bd_ram_mem1_reg[105][8]/P0001 , \wishbone_bd_ram_mem1_reg[105][9]/P0001 , \wishbone_bd_ram_mem1_reg[106][10]/P0001 , \wishbone_bd_ram_mem1_reg[106][11]/P0001 , \wishbone_bd_ram_mem1_reg[106][12]/P0001 , \wishbone_bd_ram_mem1_reg[106][13]/P0001 , \wishbone_bd_ram_mem1_reg[106][14]/P0001 , \wishbone_bd_ram_mem1_reg[106][15]/P0001 , \wishbone_bd_ram_mem1_reg[106][8]/P0001 , \wishbone_bd_ram_mem1_reg[106][9]/P0001 , \wishbone_bd_ram_mem1_reg[107][10]/P0001 , \wishbone_bd_ram_mem1_reg[107][11]/P0001 , \wishbone_bd_ram_mem1_reg[107][12]/P0001 , \wishbone_bd_ram_mem1_reg[107][13]/P0001 , \wishbone_bd_ram_mem1_reg[107][14]/P0001 , \wishbone_bd_ram_mem1_reg[107][15]/P0001 , \wishbone_bd_ram_mem1_reg[107][8]/P0001 , \wishbone_bd_ram_mem1_reg[107][9]/P0001 , \wishbone_bd_ram_mem1_reg[108][10]/P0001 , \wishbone_bd_ram_mem1_reg[108][11]/P0001 , \wishbone_bd_ram_mem1_reg[108][12]/P0001 , \wishbone_bd_ram_mem1_reg[108][13]/P0001 , \wishbone_bd_ram_mem1_reg[108][14]/P0001 , \wishbone_bd_ram_mem1_reg[108][15]/P0001 , \wishbone_bd_ram_mem1_reg[108][8]/P0001 , \wishbone_bd_ram_mem1_reg[108][9]/P0001 , \wishbone_bd_ram_mem1_reg[109][10]/P0001 , \wishbone_bd_ram_mem1_reg[109][11]/P0001 , \wishbone_bd_ram_mem1_reg[109][12]/P0001 , \wishbone_bd_ram_mem1_reg[109][13]/P0001 , \wishbone_bd_ram_mem1_reg[109][14]/P0001 , \wishbone_bd_ram_mem1_reg[109][15]/P0001 , \wishbone_bd_ram_mem1_reg[109][8]/P0001 , \wishbone_bd_ram_mem1_reg[109][9]/P0001 , \wishbone_bd_ram_mem1_reg[10][10]/P0001 , \wishbone_bd_ram_mem1_reg[10][11]/P0001 , \wishbone_bd_ram_mem1_reg[10][12]/P0001 , \wishbone_bd_ram_mem1_reg[10][13]/P0001 , \wishbone_bd_ram_mem1_reg[10][14]/P0001 , \wishbone_bd_ram_mem1_reg[10][15]/P0001 , \wishbone_bd_ram_mem1_reg[10][8]/P0001 , \wishbone_bd_ram_mem1_reg[10][9]/P0001 , \wishbone_bd_ram_mem1_reg[110][10]/P0001 , \wishbone_bd_ram_mem1_reg[110][11]/P0001 , \wishbone_bd_ram_mem1_reg[110][12]/P0001 , \wishbone_bd_ram_mem1_reg[110][13]/P0001 , \wishbone_bd_ram_mem1_reg[110][14]/P0001 , \wishbone_bd_ram_mem1_reg[110][15]/P0001 , \wishbone_bd_ram_mem1_reg[110][8]/P0001 , \wishbone_bd_ram_mem1_reg[110][9]/P0001 , \wishbone_bd_ram_mem1_reg[111][10]/P0001 , \wishbone_bd_ram_mem1_reg[111][11]/P0001 , \wishbone_bd_ram_mem1_reg[111][12]/P0001 , \wishbone_bd_ram_mem1_reg[111][13]/P0001 , \wishbone_bd_ram_mem1_reg[111][14]/P0001 , \wishbone_bd_ram_mem1_reg[111][15]/P0001 , \wishbone_bd_ram_mem1_reg[111][8]/P0001 , \wishbone_bd_ram_mem1_reg[111][9]/P0001 , \wishbone_bd_ram_mem1_reg[112][10]/P0001 , \wishbone_bd_ram_mem1_reg[112][11]/P0001 , \wishbone_bd_ram_mem1_reg[112][12]/P0001 , \wishbone_bd_ram_mem1_reg[112][13]/P0001 , \wishbone_bd_ram_mem1_reg[112][14]/P0001 , \wishbone_bd_ram_mem1_reg[112][15]/P0001 , \wishbone_bd_ram_mem1_reg[112][8]/P0001 , \wishbone_bd_ram_mem1_reg[112][9]/P0001 , \wishbone_bd_ram_mem1_reg[113][10]/P0001 , \wishbone_bd_ram_mem1_reg[113][11]/P0001 , \wishbone_bd_ram_mem1_reg[113][12]/P0001 , \wishbone_bd_ram_mem1_reg[113][13]/P0001 , \wishbone_bd_ram_mem1_reg[113][14]/P0001 , \wishbone_bd_ram_mem1_reg[113][15]/P0001 , \wishbone_bd_ram_mem1_reg[113][8]/P0001 , \wishbone_bd_ram_mem1_reg[113][9]/P0001 , \wishbone_bd_ram_mem1_reg[114][10]/P0001 , \wishbone_bd_ram_mem1_reg[114][11]/P0001 , \wishbone_bd_ram_mem1_reg[114][12]/P0001 , \wishbone_bd_ram_mem1_reg[114][13]/P0001 , \wishbone_bd_ram_mem1_reg[114][14]/P0001 , \wishbone_bd_ram_mem1_reg[114][15]/P0001 , \wishbone_bd_ram_mem1_reg[114][8]/P0001 , \wishbone_bd_ram_mem1_reg[114][9]/P0001 , \wishbone_bd_ram_mem1_reg[115][10]/P0001 , \wishbone_bd_ram_mem1_reg[115][11]/P0001 , \wishbone_bd_ram_mem1_reg[115][12]/P0001 , \wishbone_bd_ram_mem1_reg[115][13]/P0001 , \wishbone_bd_ram_mem1_reg[115][14]/P0001 , \wishbone_bd_ram_mem1_reg[115][15]/P0001 , \wishbone_bd_ram_mem1_reg[115][8]/P0001 , \wishbone_bd_ram_mem1_reg[115][9]/P0001 , \wishbone_bd_ram_mem1_reg[116][10]/P0001 , \wishbone_bd_ram_mem1_reg[116][11]/P0001 , \wishbone_bd_ram_mem1_reg[116][12]/P0001 , \wishbone_bd_ram_mem1_reg[116][13]/P0001 , \wishbone_bd_ram_mem1_reg[116][14]/P0001 , \wishbone_bd_ram_mem1_reg[116][15]/P0001 , \wishbone_bd_ram_mem1_reg[116][8]/P0001 , \wishbone_bd_ram_mem1_reg[116][9]/P0001 , \wishbone_bd_ram_mem1_reg[117][10]/P0001 , \wishbone_bd_ram_mem1_reg[117][11]/P0001 , \wishbone_bd_ram_mem1_reg[117][12]/P0001 , \wishbone_bd_ram_mem1_reg[117][13]/P0001 , \wishbone_bd_ram_mem1_reg[117][14]/P0001 , \wishbone_bd_ram_mem1_reg[117][15]/P0001 , \wishbone_bd_ram_mem1_reg[117][8]/P0001 , \wishbone_bd_ram_mem1_reg[117][9]/P0001 , \wishbone_bd_ram_mem1_reg[118][10]/P0001 , \wishbone_bd_ram_mem1_reg[118][11]/P0001 , \wishbone_bd_ram_mem1_reg[118][12]/P0001 , \wishbone_bd_ram_mem1_reg[118][13]/P0001 , \wishbone_bd_ram_mem1_reg[118][14]/P0001 , \wishbone_bd_ram_mem1_reg[118][15]/P0001 , \wishbone_bd_ram_mem1_reg[118][8]/P0001 , \wishbone_bd_ram_mem1_reg[118][9]/P0001 , \wishbone_bd_ram_mem1_reg[119][10]/P0001 , \wishbone_bd_ram_mem1_reg[119][11]/P0001 , \wishbone_bd_ram_mem1_reg[119][12]/P0001 , \wishbone_bd_ram_mem1_reg[119][13]/P0001 , \wishbone_bd_ram_mem1_reg[119][14]/P0001 , \wishbone_bd_ram_mem1_reg[119][15]/P0001 , \wishbone_bd_ram_mem1_reg[119][8]/P0001 , \wishbone_bd_ram_mem1_reg[119][9]/P0001 , \wishbone_bd_ram_mem1_reg[11][10]/P0001 , \wishbone_bd_ram_mem1_reg[11][11]/P0001 , \wishbone_bd_ram_mem1_reg[11][12]/P0001 , \wishbone_bd_ram_mem1_reg[11][13]/P0001 , \wishbone_bd_ram_mem1_reg[11][14]/P0001 , \wishbone_bd_ram_mem1_reg[11][15]/P0001 , \wishbone_bd_ram_mem1_reg[11][8]/P0001 , \wishbone_bd_ram_mem1_reg[11][9]/P0001 , \wishbone_bd_ram_mem1_reg[120][10]/P0001 , \wishbone_bd_ram_mem1_reg[120][11]/P0001 , \wishbone_bd_ram_mem1_reg[120][12]/P0001 , \wishbone_bd_ram_mem1_reg[120][13]/P0001 , \wishbone_bd_ram_mem1_reg[120][14]/P0001 , \wishbone_bd_ram_mem1_reg[120][15]/P0001 , \wishbone_bd_ram_mem1_reg[120][8]/P0001 , \wishbone_bd_ram_mem1_reg[120][9]/P0001 , \wishbone_bd_ram_mem1_reg[121][10]/P0001 , \wishbone_bd_ram_mem1_reg[121][11]/P0001 , \wishbone_bd_ram_mem1_reg[121][12]/P0001 , \wishbone_bd_ram_mem1_reg[121][13]/P0001 , \wishbone_bd_ram_mem1_reg[121][14]/P0001 , \wishbone_bd_ram_mem1_reg[121][15]/P0001 , \wishbone_bd_ram_mem1_reg[121][8]/P0001 , \wishbone_bd_ram_mem1_reg[121][9]/P0001 , \wishbone_bd_ram_mem1_reg[122][10]/P0001 , \wishbone_bd_ram_mem1_reg[122][11]/P0001 , \wishbone_bd_ram_mem1_reg[122][12]/P0001 , \wishbone_bd_ram_mem1_reg[122][13]/P0001 , \wishbone_bd_ram_mem1_reg[122][14]/P0001 , \wishbone_bd_ram_mem1_reg[122][15]/P0001 , \wishbone_bd_ram_mem1_reg[122][8]/P0001 , \wishbone_bd_ram_mem1_reg[122][9]/P0001 , \wishbone_bd_ram_mem1_reg[123][10]/P0001 , \wishbone_bd_ram_mem1_reg[123][11]/P0001 , \wishbone_bd_ram_mem1_reg[123][12]/P0001 , \wishbone_bd_ram_mem1_reg[123][13]/P0001 , \wishbone_bd_ram_mem1_reg[123][14]/P0001 , \wishbone_bd_ram_mem1_reg[123][15]/P0001 , \wishbone_bd_ram_mem1_reg[123][8]/P0001 , \wishbone_bd_ram_mem1_reg[123][9]/P0001 , \wishbone_bd_ram_mem1_reg[124][10]/P0001 , \wishbone_bd_ram_mem1_reg[124][11]/P0001 , \wishbone_bd_ram_mem1_reg[124][12]/P0001 , \wishbone_bd_ram_mem1_reg[124][13]/P0001 , \wishbone_bd_ram_mem1_reg[124][14]/P0001 , \wishbone_bd_ram_mem1_reg[124][15]/P0001 , \wishbone_bd_ram_mem1_reg[124][8]/P0001 , \wishbone_bd_ram_mem1_reg[124][9]/P0001 , \wishbone_bd_ram_mem1_reg[125][10]/P0001 , \wishbone_bd_ram_mem1_reg[125][11]/P0001 , \wishbone_bd_ram_mem1_reg[125][12]/P0001 , \wishbone_bd_ram_mem1_reg[125][13]/P0001 , \wishbone_bd_ram_mem1_reg[125][14]/P0001 , \wishbone_bd_ram_mem1_reg[125][15]/P0001 , \wishbone_bd_ram_mem1_reg[125][8]/P0001 , \wishbone_bd_ram_mem1_reg[125][9]/P0001 , \wishbone_bd_ram_mem1_reg[126][10]/P0001 , \wishbone_bd_ram_mem1_reg[126][11]/P0001 , \wishbone_bd_ram_mem1_reg[126][12]/P0001 , \wishbone_bd_ram_mem1_reg[126][13]/P0001 , \wishbone_bd_ram_mem1_reg[126][14]/P0001 , \wishbone_bd_ram_mem1_reg[126][15]/P0001 , \wishbone_bd_ram_mem1_reg[126][8]/P0001 , \wishbone_bd_ram_mem1_reg[126][9]/P0001 , \wishbone_bd_ram_mem1_reg[127][10]/P0001 , \wishbone_bd_ram_mem1_reg[127][11]/P0001 , \wishbone_bd_ram_mem1_reg[127][12]/P0001 , \wishbone_bd_ram_mem1_reg[127][13]/P0001 , \wishbone_bd_ram_mem1_reg[127][14]/P0001 , \wishbone_bd_ram_mem1_reg[127][15]/P0001 , \wishbone_bd_ram_mem1_reg[127][8]/P0001 , \wishbone_bd_ram_mem1_reg[127][9]/P0001 , \wishbone_bd_ram_mem1_reg[128][10]/P0001 , \wishbone_bd_ram_mem1_reg[128][11]/P0001 , \wishbone_bd_ram_mem1_reg[128][12]/P0001 , \wishbone_bd_ram_mem1_reg[128][13]/P0001 , \wishbone_bd_ram_mem1_reg[128][14]/P0001 , \wishbone_bd_ram_mem1_reg[128][15]/P0001 , \wishbone_bd_ram_mem1_reg[128][8]/P0001 , \wishbone_bd_ram_mem1_reg[128][9]/P0001 , \wishbone_bd_ram_mem1_reg[129][10]/P0001 , \wishbone_bd_ram_mem1_reg[129][11]/P0001 , \wishbone_bd_ram_mem1_reg[129][12]/P0001 , \wishbone_bd_ram_mem1_reg[129][13]/P0001 , \wishbone_bd_ram_mem1_reg[129][14]/P0001 , \wishbone_bd_ram_mem1_reg[129][15]/P0001 , \wishbone_bd_ram_mem1_reg[129][8]/P0001 , \wishbone_bd_ram_mem1_reg[129][9]/P0001 , \wishbone_bd_ram_mem1_reg[12][10]/P0001 , \wishbone_bd_ram_mem1_reg[12][11]/P0001 , \wishbone_bd_ram_mem1_reg[12][12]/P0001 , \wishbone_bd_ram_mem1_reg[12][13]/P0001 , \wishbone_bd_ram_mem1_reg[12][14]/P0001 , \wishbone_bd_ram_mem1_reg[12][15]/P0001 , \wishbone_bd_ram_mem1_reg[12][8]/P0001 , \wishbone_bd_ram_mem1_reg[12][9]/P0001 , \wishbone_bd_ram_mem1_reg[130][10]/P0001 , \wishbone_bd_ram_mem1_reg[130][11]/P0001 , \wishbone_bd_ram_mem1_reg[130][12]/P0001 , \wishbone_bd_ram_mem1_reg[130][13]/P0001 , \wishbone_bd_ram_mem1_reg[130][14]/P0001 , \wishbone_bd_ram_mem1_reg[130][15]/P0001 , \wishbone_bd_ram_mem1_reg[130][8]/P0001 , \wishbone_bd_ram_mem1_reg[130][9]/P0001 , \wishbone_bd_ram_mem1_reg[131][10]/P0001 , \wishbone_bd_ram_mem1_reg[131][11]/P0001 , \wishbone_bd_ram_mem1_reg[131][12]/P0001 , \wishbone_bd_ram_mem1_reg[131][13]/P0001 , \wishbone_bd_ram_mem1_reg[131][14]/P0001 , \wishbone_bd_ram_mem1_reg[131][15]/P0001 , \wishbone_bd_ram_mem1_reg[131][8]/P0001 , \wishbone_bd_ram_mem1_reg[131][9]/P0001 , \wishbone_bd_ram_mem1_reg[132][10]/P0001 , \wishbone_bd_ram_mem1_reg[132][11]/P0001 , \wishbone_bd_ram_mem1_reg[132][12]/P0001 , \wishbone_bd_ram_mem1_reg[132][13]/P0001 , \wishbone_bd_ram_mem1_reg[132][14]/P0001 , \wishbone_bd_ram_mem1_reg[132][15]/P0001 , \wishbone_bd_ram_mem1_reg[132][8]/P0001 , \wishbone_bd_ram_mem1_reg[132][9]/P0001 , \wishbone_bd_ram_mem1_reg[133][10]/P0001 , \wishbone_bd_ram_mem1_reg[133][11]/P0001 , \wishbone_bd_ram_mem1_reg[133][12]/P0001 , \wishbone_bd_ram_mem1_reg[133][13]/P0001 , \wishbone_bd_ram_mem1_reg[133][14]/P0001 , \wishbone_bd_ram_mem1_reg[133][15]/P0001 , \wishbone_bd_ram_mem1_reg[133][8]/P0001 , \wishbone_bd_ram_mem1_reg[133][9]/P0001 , \wishbone_bd_ram_mem1_reg[134][10]/P0001 , \wishbone_bd_ram_mem1_reg[134][11]/P0001 , \wishbone_bd_ram_mem1_reg[134][12]/P0001 , \wishbone_bd_ram_mem1_reg[134][13]/P0001 , \wishbone_bd_ram_mem1_reg[134][14]/P0001 , \wishbone_bd_ram_mem1_reg[134][15]/P0001 , \wishbone_bd_ram_mem1_reg[134][8]/P0001 , \wishbone_bd_ram_mem1_reg[134][9]/P0001 , \wishbone_bd_ram_mem1_reg[135][10]/P0001 , \wishbone_bd_ram_mem1_reg[135][11]/P0001 , \wishbone_bd_ram_mem1_reg[135][12]/P0001 , \wishbone_bd_ram_mem1_reg[135][13]/P0001 , \wishbone_bd_ram_mem1_reg[135][14]/P0001 , \wishbone_bd_ram_mem1_reg[135][15]/P0001 , \wishbone_bd_ram_mem1_reg[135][8]/P0001 , \wishbone_bd_ram_mem1_reg[135][9]/P0001 , \wishbone_bd_ram_mem1_reg[136][10]/P0001 , \wishbone_bd_ram_mem1_reg[136][11]/P0001 , \wishbone_bd_ram_mem1_reg[136][12]/P0001 , \wishbone_bd_ram_mem1_reg[136][13]/P0001 , \wishbone_bd_ram_mem1_reg[136][14]/P0001 , \wishbone_bd_ram_mem1_reg[136][15]/P0001 , \wishbone_bd_ram_mem1_reg[136][8]/P0001 , \wishbone_bd_ram_mem1_reg[136][9]/P0001 , \wishbone_bd_ram_mem1_reg[137][10]/P0001 , \wishbone_bd_ram_mem1_reg[137][11]/P0001 , \wishbone_bd_ram_mem1_reg[137][12]/P0001 , \wishbone_bd_ram_mem1_reg[137][13]/P0001 , \wishbone_bd_ram_mem1_reg[137][14]/P0001 , \wishbone_bd_ram_mem1_reg[137][15]/P0001 , \wishbone_bd_ram_mem1_reg[137][8]/P0001 , \wishbone_bd_ram_mem1_reg[137][9]/P0001 , \wishbone_bd_ram_mem1_reg[138][10]/P0001 , \wishbone_bd_ram_mem1_reg[138][11]/P0001 , \wishbone_bd_ram_mem1_reg[138][12]/P0001 , \wishbone_bd_ram_mem1_reg[138][13]/P0001 , \wishbone_bd_ram_mem1_reg[138][14]/P0001 , \wishbone_bd_ram_mem1_reg[138][15]/P0001 , \wishbone_bd_ram_mem1_reg[138][8]/P0001 , \wishbone_bd_ram_mem1_reg[138][9]/P0001 , \wishbone_bd_ram_mem1_reg[139][10]/P0001 , \wishbone_bd_ram_mem1_reg[139][11]/P0001 , \wishbone_bd_ram_mem1_reg[139][12]/P0001 , \wishbone_bd_ram_mem1_reg[139][13]/P0001 , \wishbone_bd_ram_mem1_reg[139][14]/P0001 , \wishbone_bd_ram_mem1_reg[139][15]/P0001 , \wishbone_bd_ram_mem1_reg[139][8]/P0001 , \wishbone_bd_ram_mem1_reg[139][9]/P0001 , \wishbone_bd_ram_mem1_reg[13][10]/P0001 , \wishbone_bd_ram_mem1_reg[13][11]/P0001 , \wishbone_bd_ram_mem1_reg[13][12]/P0001 , \wishbone_bd_ram_mem1_reg[13][13]/P0001 , \wishbone_bd_ram_mem1_reg[13][14]/P0001 , \wishbone_bd_ram_mem1_reg[13][15]/P0001 , \wishbone_bd_ram_mem1_reg[13][8]/P0001 , \wishbone_bd_ram_mem1_reg[13][9]/P0001 , \wishbone_bd_ram_mem1_reg[140][10]/P0001 , \wishbone_bd_ram_mem1_reg[140][11]/P0001 , \wishbone_bd_ram_mem1_reg[140][12]/P0001 , \wishbone_bd_ram_mem1_reg[140][13]/P0001 , \wishbone_bd_ram_mem1_reg[140][14]/P0001 , \wishbone_bd_ram_mem1_reg[140][15]/P0001 , \wishbone_bd_ram_mem1_reg[140][8]/P0001 , \wishbone_bd_ram_mem1_reg[140][9]/P0001 , \wishbone_bd_ram_mem1_reg[141][10]/P0001 , \wishbone_bd_ram_mem1_reg[141][11]/P0001 , \wishbone_bd_ram_mem1_reg[141][12]/P0001 , \wishbone_bd_ram_mem1_reg[141][13]/P0001 , \wishbone_bd_ram_mem1_reg[141][14]/P0001 , \wishbone_bd_ram_mem1_reg[141][15]/P0001 , \wishbone_bd_ram_mem1_reg[141][8]/P0001 , \wishbone_bd_ram_mem1_reg[141][9]/P0001 , \wishbone_bd_ram_mem1_reg[142][10]/P0001 , \wishbone_bd_ram_mem1_reg[142][11]/P0001 , \wishbone_bd_ram_mem1_reg[142][12]/P0001 , \wishbone_bd_ram_mem1_reg[142][13]/P0001 , \wishbone_bd_ram_mem1_reg[142][14]/P0001 , \wishbone_bd_ram_mem1_reg[142][15]/P0001 , \wishbone_bd_ram_mem1_reg[142][8]/P0001 , \wishbone_bd_ram_mem1_reg[142][9]/P0001 , \wishbone_bd_ram_mem1_reg[143][10]/P0001 , \wishbone_bd_ram_mem1_reg[143][11]/P0001 , \wishbone_bd_ram_mem1_reg[143][12]/P0001 , \wishbone_bd_ram_mem1_reg[143][13]/P0001 , \wishbone_bd_ram_mem1_reg[143][14]/P0001 , \wishbone_bd_ram_mem1_reg[143][15]/P0001 , \wishbone_bd_ram_mem1_reg[143][8]/P0001 , \wishbone_bd_ram_mem1_reg[143][9]/P0001 , \wishbone_bd_ram_mem1_reg[144][10]/P0001 , \wishbone_bd_ram_mem1_reg[144][11]/P0001 , \wishbone_bd_ram_mem1_reg[144][12]/P0001 , \wishbone_bd_ram_mem1_reg[144][13]/P0001 , \wishbone_bd_ram_mem1_reg[144][14]/P0001 , \wishbone_bd_ram_mem1_reg[144][15]/P0001 , \wishbone_bd_ram_mem1_reg[144][8]/P0001 , \wishbone_bd_ram_mem1_reg[144][9]/P0001 , \wishbone_bd_ram_mem1_reg[145][10]/P0001 , \wishbone_bd_ram_mem1_reg[145][11]/P0001 , \wishbone_bd_ram_mem1_reg[145][12]/P0001 , \wishbone_bd_ram_mem1_reg[145][13]/P0001 , \wishbone_bd_ram_mem1_reg[145][14]/P0001 , \wishbone_bd_ram_mem1_reg[145][15]/P0001 , \wishbone_bd_ram_mem1_reg[145][8]/P0001 , \wishbone_bd_ram_mem1_reg[145][9]/P0001 , \wishbone_bd_ram_mem1_reg[146][10]/P0001 , \wishbone_bd_ram_mem1_reg[146][11]/P0001 , \wishbone_bd_ram_mem1_reg[146][12]/P0001 , \wishbone_bd_ram_mem1_reg[146][13]/P0001 , \wishbone_bd_ram_mem1_reg[146][14]/P0001 , \wishbone_bd_ram_mem1_reg[146][15]/P0001 , \wishbone_bd_ram_mem1_reg[146][8]/P0001 , \wishbone_bd_ram_mem1_reg[146][9]/P0001 , \wishbone_bd_ram_mem1_reg[147][10]/P0001 , \wishbone_bd_ram_mem1_reg[147][11]/P0001 , \wishbone_bd_ram_mem1_reg[147][12]/P0001 , \wishbone_bd_ram_mem1_reg[147][13]/P0001 , \wishbone_bd_ram_mem1_reg[147][14]/P0001 , \wishbone_bd_ram_mem1_reg[147][15]/P0001 , \wishbone_bd_ram_mem1_reg[147][8]/P0001 , \wishbone_bd_ram_mem1_reg[147][9]/P0001 , \wishbone_bd_ram_mem1_reg[148][10]/P0001 , \wishbone_bd_ram_mem1_reg[148][11]/P0001 , \wishbone_bd_ram_mem1_reg[148][12]/P0001 , \wishbone_bd_ram_mem1_reg[148][13]/P0001 , \wishbone_bd_ram_mem1_reg[148][14]/P0001 , \wishbone_bd_ram_mem1_reg[148][15]/P0001 , \wishbone_bd_ram_mem1_reg[148][8]/P0001 , \wishbone_bd_ram_mem1_reg[148][9]/P0001 , \wishbone_bd_ram_mem1_reg[149][10]/P0001 , \wishbone_bd_ram_mem1_reg[149][11]/P0001 , \wishbone_bd_ram_mem1_reg[149][12]/P0001 , \wishbone_bd_ram_mem1_reg[149][13]/P0001 , \wishbone_bd_ram_mem1_reg[149][14]/P0001 , \wishbone_bd_ram_mem1_reg[149][15]/P0001 , \wishbone_bd_ram_mem1_reg[149][8]/P0001 , \wishbone_bd_ram_mem1_reg[149][9]/P0001 , \wishbone_bd_ram_mem1_reg[14][10]/P0001 , \wishbone_bd_ram_mem1_reg[14][11]/P0001 , \wishbone_bd_ram_mem1_reg[14][12]/P0001 , \wishbone_bd_ram_mem1_reg[14][13]/P0001 , \wishbone_bd_ram_mem1_reg[14][14]/P0001 , \wishbone_bd_ram_mem1_reg[14][15]/P0001 , \wishbone_bd_ram_mem1_reg[14][8]/P0001 , \wishbone_bd_ram_mem1_reg[14][9]/P0001 , \wishbone_bd_ram_mem1_reg[150][10]/P0001 , \wishbone_bd_ram_mem1_reg[150][11]/P0001 , \wishbone_bd_ram_mem1_reg[150][12]/P0001 , \wishbone_bd_ram_mem1_reg[150][13]/P0001 , \wishbone_bd_ram_mem1_reg[150][14]/P0001 , \wishbone_bd_ram_mem1_reg[150][15]/P0001 , \wishbone_bd_ram_mem1_reg[150][8]/P0001 , \wishbone_bd_ram_mem1_reg[150][9]/P0001 , \wishbone_bd_ram_mem1_reg[151][10]/P0001 , \wishbone_bd_ram_mem1_reg[151][11]/P0001 , \wishbone_bd_ram_mem1_reg[151][12]/P0001 , \wishbone_bd_ram_mem1_reg[151][13]/P0001 , \wishbone_bd_ram_mem1_reg[151][14]/P0001 , \wishbone_bd_ram_mem1_reg[151][15]/P0001 , \wishbone_bd_ram_mem1_reg[151][8]/P0001 , \wishbone_bd_ram_mem1_reg[151][9]/P0001 , \wishbone_bd_ram_mem1_reg[152][10]/P0001 , \wishbone_bd_ram_mem1_reg[152][11]/P0001 , \wishbone_bd_ram_mem1_reg[152][12]/P0001 , \wishbone_bd_ram_mem1_reg[152][13]/P0001 , \wishbone_bd_ram_mem1_reg[152][14]/P0001 , \wishbone_bd_ram_mem1_reg[152][15]/P0001 , \wishbone_bd_ram_mem1_reg[152][8]/P0001 , \wishbone_bd_ram_mem1_reg[152][9]/P0001 , \wishbone_bd_ram_mem1_reg[153][10]/P0001 , \wishbone_bd_ram_mem1_reg[153][11]/P0001 , \wishbone_bd_ram_mem1_reg[153][12]/P0001 , \wishbone_bd_ram_mem1_reg[153][13]/P0001 , \wishbone_bd_ram_mem1_reg[153][14]/P0001 , \wishbone_bd_ram_mem1_reg[153][15]/P0001 , \wishbone_bd_ram_mem1_reg[153][8]/P0001 , \wishbone_bd_ram_mem1_reg[153][9]/P0001 , \wishbone_bd_ram_mem1_reg[154][10]/P0001 , \wishbone_bd_ram_mem1_reg[154][11]/P0001 , \wishbone_bd_ram_mem1_reg[154][12]/P0001 , \wishbone_bd_ram_mem1_reg[154][13]/P0001 , \wishbone_bd_ram_mem1_reg[154][14]/P0001 , \wishbone_bd_ram_mem1_reg[154][15]/P0001 , \wishbone_bd_ram_mem1_reg[154][8]/P0001 , \wishbone_bd_ram_mem1_reg[154][9]/P0001 , \wishbone_bd_ram_mem1_reg[155][10]/P0001 , \wishbone_bd_ram_mem1_reg[155][11]/P0001 , \wishbone_bd_ram_mem1_reg[155][12]/P0001 , \wishbone_bd_ram_mem1_reg[155][13]/P0001 , \wishbone_bd_ram_mem1_reg[155][14]/P0001 , \wishbone_bd_ram_mem1_reg[155][15]/P0001 , \wishbone_bd_ram_mem1_reg[155][8]/P0001 , \wishbone_bd_ram_mem1_reg[155][9]/P0001 , \wishbone_bd_ram_mem1_reg[156][10]/P0001 , \wishbone_bd_ram_mem1_reg[156][11]/P0001 , \wishbone_bd_ram_mem1_reg[156][12]/P0001 , \wishbone_bd_ram_mem1_reg[156][13]/P0001 , \wishbone_bd_ram_mem1_reg[156][14]/P0001 , \wishbone_bd_ram_mem1_reg[156][15]/P0001 , \wishbone_bd_ram_mem1_reg[156][8]/P0001 , \wishbone_bd_ram_mem1_reg[156][9]/P0001 , \wishbone_bd_ram_mem1_reg[157][10]/P0001 , \wishbone_bd_ram_mem1_reg[157][11]/P0001 , \wishbone_bd_ram_mem1_reg[157][12]/P0001 , \wishbone_bd_ram_mem1_reg[157][13]/P0001 , \wishbone_bd_ram_mem1_reg[157][14]/P0001 , \wishbone_bd_ram_mem1_reg[157][15]/P0001 , \wishbone_bd_ram_mem1_reg[157][8]/P0001 , \wishbone_bd_ram_mem1_reg[157][9]/P0001 , \wishbone_bd_ram_mem1_reg[158][10]/P0001 , \wishbone_bd_ram_mem1_reg[158][11]/P0001 , \wishbone_bd_ram_mem1_reg[158][12]/P0001 , \wishbone_bd_ram_mem1_reg[158][13]/P0001 , \wishbone_bd_ram_mem1_reg[158][14]/P0001 , \wishbone_bd_ram_mem1_reg[158][15]/P0001 , \wishbone_bd_ram_mem1_reg[158][8]/P0001 , \wishbone_bd_ram_mem1_reg[158][9]/P0001 , \wishbone_bd_ram_mem1_reg[159][10]/P0001 , \wishbone_bd_ram_mem1_reg[159][11]/P0001 , \wishbone_bd_ram_mem1_reg[159][12]/P0001 , \wishbone_bd_ram_mem1_reg[159][13]/P0001 , \wishbone_bd_ram_mem1_reg[159][14]/P0001 , \wishbone_bd_ram_mem1_reg[159][15]/P0001 , \wishbone_bd_ram_mem1_reg[159][8]/P0001 , \wishbone_bd_ram_mem1_reg[159][9]/P0001 , \wishbone_bd_ram_mem1_reg[15][10]/P0001 , \wishbone_bd_ram_mem1_reg[15][11]/P0001 , \wishbone_bd_ram_mem1_reg[15][12]/P0001 , \wishbone_bd_ram_mem1_reg[15][13]/P0001 , \wishbone_bd_ram_mem1_reg[15][14]/P0001 , \wishbone_bd_ram_mem1_reg[15][15]/P0001 , \wishbone_bd_ram_mem1_reg[15][8]/P0001 , \wishbone_bd_ram_mem1_reg[15][9]/P0001 , \wishbone_bd_ram_mem1_reg[160][10]/P0001 , \wishbone_bd_ram_mem1_reg[160][11]/P0001 , \wishbone_bd_ram_mem1_reg[160][12]/P0001 , \wishbone_bd_ram_mem1_reg[160][13]/P0001 , \wishbone_bd_ram_mem1_reg[160][14]/P0001 , \wishbone_bd_ram_mem1_reg[160][15]/P0001 , \wishbone_bd_ram_mem1_reg[160][8]/P0001 , \wishbone_bd_ram_mem1_reg[160][9]/P0001 , \wishbone_bd_ram_mem1_reg[161][10]/P0001 , \wishbone_bd_ram_mem1_reg[161][11]/P0001 , \wishbone_bd_ram_mem1_reg[161][12]/P0001 , \wishbone_bd_ram_mem1_reg[161][13]/P0001 , \wishbone_bd_ram_mem1_reg[161][14]/P0001 , \wishbone_bd_ram_mem1_reg[161][15]/P0001 , \wishbone_bd_ram_mem1_reg[161][8]/P0001 , \wishbone_bd_ram_mem1_reg[161][9]/P0001 , \wishbone_bd_ram_mem1_reg[162][10]/P0001 , \wishbone_bd_ram_mem1_reg[162][11]/P0001 , \wishbone_bd_ram_mem1_reg[162][12]/P0001 , \wishbone_bd_ram_mem1_reg[162][13]/P0001 , \wishbone_bd_ram_mem1_reg[162][14]/P0001 , \wishbone_bd_ram_mem1_reg[162][15]/P0001 , \wishbone_bd_ram_mem1_reg[162][8]/P0001 , \wishbone_bd_ram_mem1_reg[162][9]/P0001 , \wishbone_bd_ram_mem1_reg[163][10]/P0001 , \wishbone_bd_ram_mem1_reg[163][11]/P0001 , \wishbone_bd_ram_mem1_reg[163][12]/P0001 , \wishbone_bd_ram_mem1_reg[163][13]/P0001 , \wishbone_bd_ram_mem1_reg[163][14]/P0001 , \wishbone_bd_ram_mem1_reg[163][15]/P0001 , \wishbone_bd_ram_mem1_reg[163][8]/P0001 , \wishbone_bd_ram_mem1_reg[163][9]/P0001 , \wishbone_bd_ram_mem1_reg[164][10]/P0001 , \wishbone_bd_ram_mem1_reg[164][11]/P0001 , \wishbone_bd_ram_mem1_reg[164][12]/P0001 , \wishbone_bd_ram_mem1_reg[164][13]/P0001 , \wishbone_bd_ram_mem1_reg[164][14]/P0001 , \wishbone_bd_ram_mem1_reg[164][15]/P0001 , \wishbone_bd_ram_mem1_reg[164][8]/P0001 , \wishbone_bd_ram_mem1_reg[164][9]/P0001 , \wishbone_bd_ram_mem1_reg[165][10]/P0001 , \wishbone_bd_ram_mem1_reg[165][11]/P0001 , \wishbone_bd_ram_mem1_reg[165][12]/P0001 , \wishbone_bd_ram_mem1_reg[165][13]/P0001 , \wishbone_bd_ram_mem1_reg[165][14]/P0001 , \wishbone_bd_ram_mem1_reg[165][15]/P0001 , \wishbone_bd_ram_mem1_reg[165][8]/P0001 , \wishbone_bd_ram_mem1_reg[165][9]/P0001 , \wishbone_bd_ram_mem1_reg[166][10]/P0001 , \wishbone_bd_ram_mem1_reg[166][11]/P0001 , \wishbone_bd_ram_mem1_reg[166][12]/P0001 , \wishbone_bd_ram_mem1_reg[166][13]/P0001 , \wishbone_bd_ram_mem1_reg[166][14]/P0001 , \wishbone_bd_ram_mem1_reg[166][15]/P0001 , \wishbone_bd_ram_mem1_reg[166][8]/P0001 , \wishbone_bd_ram_mem1_reg[166][9]/P0001 , \wishbone_bd_ram_mem1_reg[167][10]/P0001 , \wishbone_bd_ram_mem1_reg[167][11]/P0001 , \wishbone_bd_ram_mem1_reg[167][12]/P0001 , \wishbone_bd_ram_mem1_reg[167][13]/P0001 , \wishbone_bd_ram_mem1_reg[167][14]/P0001 , \wishbone_bd_ram_mem1_reg[167][15]/P0001 , \wishbone_bd_ram_mem1_reg[167][8]/P0001 , \wishbone_bd_ram_mem1_reg[167][9]/P0001 , \wishbone_bd_ram_mem1_reg[168][10]/P0001 , \wishbone_bd_ram_mem1_reg[168][11]/P0001 , \wishbone_bd_ram_mem1_reg[168][12]/P0001 , \wishbone_bd_ram_mem1_reg[168][13]/P0001 , \wishbone_bd_ram_mem1_reg[168][14]/P0001 , \wishbone_bd_ram_mem1_reg[168][15]/P0001 , \wishbone_bd_ram_mem1_reg[168][8]/P0001 , \wishbone_bd_ram_mem1_reg[168][9]/P0001 , \wishbone_bd_ram_mem1_reg[169][10]/P0001 , \wishbone_bd_ram_mem1_reg[169][11]/P0001 , \wishbone_bd_ram_mem1_reg[169][12]/P0001 , \wishbone_bd_ram_mem1_reg[169][13]/P0001 , \wishbone_bd_ram_mem1_reg[169][14]/P0001 , \wishbone_bd_ram_mem1_reg[169][15]/P0001 , \wishbone_bd_ram_mem1_reg[169][8]/P0001 , \wishbone_bd_ram_mem1_reg[169][9]/P0001 , \wishbone_bd_ram_mem1_reg[16][10]/P0001 , \wishbone_bd_ram_mem1_reg[16][11]/P0001 , \wishbone_bd_ram_mem1_reg[16][12]/P0001 , \wishbone_bd_ram_mem1_reg[16][13]/P0001 , \wishbone_bd_ram_mem1_reg[16][14]/P0001 , \wishbone_bd_ram_mem1_reg[16][15]/P0001 , \wishbone_bd_ram_mem1_reg[16][8]/P0001 , \wishbone_bd_ram_mem1_reg[16][9]/P0001 , \wishbone_bd_ram_mem1_reg[170][10]/P0001 , \wishbone_bd_ram_mem1_reg[170][11]/P0001 , \wishbone_bd_ram_mem1_reg[170][12]/P0001 , \wishbone_bd_ram_mem1_reg[170][13]/P0001 , \wishbone_bd_ram_mem1_reg[170][14]/P0001 , \wishbone_bd_ram_mem1_reg[170][15]/P0001 , \wishbone_bd_ram_mem1_reg[170][8]/P0001 , \wishbone_bd_ram_mem1_reg[170][9]/P0001 , \wishbone_bd_ram_mem1_reg[171][10]/P0001 , \wishbone_bd_ram_mem1_reg[171][11]/P0001 , \wishbone_bd_ram_mem1_reg[171][12]/P0001 , \wishbone_bd_ram_mem1_reg[171][13]/P0001 , \wishbone_bd_ram_mem1_reg[171][14]/P0001 , \wishbone_bd_ram_mem1_reg[171][15]/P0001 , \wishbone_bd_ram_mem1_reg[171][8]/P0001 , \wishbone_bd_ram_mem1_reg[171][9]/P0001 , \wishbone_bd_ram_mem1_reg[172][10]/P0001 , \wishbone_bd_ram_mem1_reg[172][11]/P0001 , \wishbone_bd_ram_mem1_reg[172][12]/P0001 , \wishbone_bd_ram_mem1_reg[172][13]/P0001 , \wishbone_bd_ram_mem1_reg[172][14]/P0001 , \wishbone_bd_ram_mem1_reg[172][15]/P0001 , \wishbone_bd_ram_mem1_reg[172][8]/P0001 , \wishbone_bd_ram_mem1_reg[172][9]/P0001 , \wishbone_bd_ram_mem1_reg[173][10]/P0001 , \wishbone_bd_ram_mem1_reg[173][11]/P0001 , \wishbone_bd_ram_mem1_reg[173][12]/P0001 , \wishbone_bd_ram_mem1_reg[173][13]/P0001 , \wishbone_bd_ram_mem1_reg[173][14]/P0001 , \wishbone_bd_ram_mem1_reg[173][15]/P0001 , \wishbone_bd_ram_mem1_reg[173][8]/P0001 , \wishbone_bd_ram_mem1_reg[173][9]/P0001 , \wishbone_bd_ram_mem1_reg[174][10]/P0001 , \wishbone_bd_ram_mem1_reg[174][11]/P0001 , \wishbone_bd_ram_mem1_reg[174][12]/P0001 , \wishbone_bd_ram_mem1_reg[174][13]/P0001 , \wishbone_bd_ram_mem1_reg[174][14]/P0001 , \wishbone_bd_ram_mem1_reg[174][15]/P0001 , \wishbone_bd_ram_mem1_reg[174][8]/P0001 , \wishbone_bd_ram_mem1_reg[174][9]/P0001 , \wishbone_bd_ram_mem1_reg[175][10]/P0001 , \wishbone_bd_ram_mem1_reg[175][11]/P0001 , \wishbone_bd_ram_mem1_reg[175][12]/P0001 , \wishbone_bd_ram_mem1_reg[175][13]/P0001 , \wishbone_bd_ram_mem1_reg[175][14]/P0001 , \wishbone_bd_ram_mem1_reg[175][15]/P0001 , \wishbone_bd_ram_mem1_reg[175][8]/P0001 , \wishbone_bd_ram_mem1_reg[175][9]/P0001 , \wishbone_bd_ram_mem1_reg[176][10]/P0001 , \wishbone_bd_ram_mem1_reg[176][11]/P0001 , \wishbone_bd_ram_mem1_reg[176][12]/P0001 , \wishbone_bd_ram_mem1_reg[176][13]/P0001 , \wishbone_bd_ram_mem1_reg[176][14]/P0001 , \wishbone_bd_ram_mem1_reg[176][15]/P0001 , \wishbone_bd_ram_mem1_reg[176][8]/P0001 , \wishbone_bd_ram_mem1_reg[176][9]/P0001 , \wishbone_bd_ram_mem1_reg[177][10]/P0001 , \wishbone_bd_ram_mem1_reg[177][11]/P0001 , \wishbone_bd_ram_mem1_reg[177][12]/P0001 , \wishbone_bd_ram_mem1_reg[177][13]/P0001 , \wishbone_bd_ram_mem1_reg[177][14]/P0001 , \wishbone_bd_ram_mem1_reg[177][15]/P0001 , \wishbone_bd_ram_mem1_reg[177][8]/P0001 , \wishbone_bd_ram_mem1_reg[177][9]/P0001 , \wishbone_bd_ram_mem1_reg[178][10]/P0001 , \wishbone_bd_ram_mem1_reg[178][11]/P0001 , \wishbone_bd_ram_mem1_reg[178][12]/P0001 , \wishbone_bd_ram_mem1_reg[178][13]/P0001 , \wishbone_bd_ram_mem1_reg[178][14]/P0001 , \wishbone_bd_ram_mem1_reg[178][15]/P0001 , \wishbone_bd_ram_mem1_reg[178][8]/P0001 , \wishbone_bd_ram_mem1_reg[178][9]/P0001 , \wishbone_bd_ram_mem1_reg[179][10]/P0001 , \wishbone_bd_ram_mem1_reg[179][11]/P0001 , \wishbone_bd_ram_mem1_reg[179][12]/P0001 , \wishbone_bd_ram_mem1_reg[179][13]/P0001 , \wishbone_bd_ram_mem1_reg[179][14]/P0001 , \wishbone_bd_ram_mem1_reg[179][15]/P0001 , \wishbone_bd_ram_mem1_reg[179][8]/P0001 , \wishbone_bd_ram_mem1_reg[179][9]/P0001 , \wishbone_bd_ram_mem1_reg[17][10]/P0001 , \wishbone_bd_ram_mem1_reg[17][11]/P0001 , \wishbone_bd_ram_mem1_reg[17][12]/P0001 , \wishbone_bd_ram_mem1_reg[17][13]/P0001 , \wishbone_bd_ram_mem1_reg[17][14]/P0001 , \wishbone_bd_ram_mem1_reg[17][15]/P0001 , \wishbone_bd_ram_mem1_reg[17][8]/P0001 , \wishbone_bd_ram_mem1_reg[17][9]/P0001 , \wishbone_bd_ram_mem1_reg[180][10]/P0001 , \wishbone_bd_ram_mem1_reg[180][11]/P0001 , \wishbone_bd_ram_mem1_reg[180][12]/P0001 , \wishbone_bd_ram_mem1_reg[180][13]/P0001 , \wishbone_bd_ram_mem1_reg[180][14]/P0001 , \wishbone_bd_ram_mem1_reg[180][15]/P0001 , \wishbone_bd_ram_mem1_reg[180][8]/P0001 , \wishbone_bd_ram_mem1_reg[180][9]/P0001 , \wishbone_bd_ram_mem1_reg[181][10]/P0001 , \wishbone_bd_ram_mem1_reg[181][11]/P0001 , \wishbone_bd_ram_mem1_reg[181][12]/P0001 , \wishbone_bd_ram_mem1_reg[181][13]/P0001 , \wishbone_bd_ram_mem1_reg[181][14]/P0001 , \wishbone_bd_ram_mem1_reg[181][15]/P0001 , \wishbone_bd_ram_mem1_reg[181][8]/P0001 , \wishbone_bd_ram_mem1_reg[181][9]/P0001 , \wishbone_bd_ram_mem1_reg[182][10]/P0001 , \wishbone_bd_ram_mem1_reg[182][11]/P0001 , \wishbone_bd_ram_mem1_reg[182][12]/P0001 , \wishbone_bd_ram_mem1_reg[182][13]/P0001 , \wishbone_bd_ram_mem1_reg[182][14]/P0001 , \wishbone_bd_ram_mem1_reg[182][15]/P0001 , \wishbone_bd_ram_mem1_reg[182][8]/P0001 , \wishbone_bd_ram_mem1_reg[182][9]/P0001 , \wishbone_bd_ram_mem1_reg[183][10]/P0001 , \wishbone_bd_ram_mem1_reg[183][11]/P0001 , \wishbone_bd_ram_mem1_reg[183][12]/P0001 , \wishbone_bd_ram_mem1_reg[183][13]/P0001 , \wishbone_bd_ram_mem1_reg[183][14]/P0001 , \wishbone_bd_ram_mem1_reg[183][15]/P0001 , \wishbone_bd_ram_mem1_reg[183][8]/P0001 , \wishbone_bd_ram_mem1_reg[183][9]/P0001 , \wishbone_bd_ram_mem1_reg[184][10]/P0001 , \wishbone_bd_ram_mem1_reg[184][11]/P0001 , \wishbone_bd_ram_mem1_reg[184][12]/P0001 , \wishbone_bd_ram_mem1_reg[184][13]/P0001 , \wishbone_bd_ram_mem1_reg[184][14]/P0001 , \wishbone_bd_ram_mem1_reg[184][15]/P0001 , \wishbone_bd_ram_mem1_reg[184][8]/P0001 , \wishbone_bd_ram_mem1_reg[184][9]/P0001 , \wishbone_bd_ram_mem1_reg[185][10]/P0001 , \wishbone_bd_ram_mem1_reg[185][11]/P0001 , \wishbone_bd_ram_mem1_reg[185][12]/P0001 , \wishbone_bd_ram_mem1_reg[185][13]/P0001 , \wishbone_bd_ram_mem1_reg[185][14]/P0001 , \wishbone_bd_ram_mem1_reg[185][15]/P0001 , \wishbone_bd_ram_mem1_reg[185][8]/P0001 , \wishbone_bd_ram_mem1_reg[185][9]/P0001 , \wishbone_bd_ram_mem1_reg[186][10]/P0001 , \wishbone_bd_ram_mem1_reg[186][11]/P0001 , \wishbone_bd_ram_mem1_reg[186][12]/P0001 , \wishbone_bd_ram_mem1_reg[186][13]/P0001 , \wishbone_bd_ram_mem1_reg[186][14]/P0001 , \wishbone_bd_ram_mem1_reg[186][15]/P0001 , \wishbone_bd_ram_mem1_reg[186][8]/P0001 , \wishbone_bd_ram_mem1_reg[186][9]/P0001 , \wishbone_bd_ram_mem1_reg[187][10]/P0001 , \wishbone_bd_ram_mem1_reg[187][11]/P0001 , \wishbone_bd_ram_mem1_reg[187][12]/P0001 , \wishbone_bd_ram_mem1_reg[187][13]/P0001 , \wishbone_bd_ram_mem1_reg[187][14]/P0001 , \wishbone_bd_ram_mem1_reg[187][15]/P0001 , \wishbone_bd_ram_mem1_reg[187][8]/P0001 , \wishbone_bd_ram_mem1_reg[187][9]/P0001 , \wishbone_bd_ram_mem1_reg[188][10]/P0001 , \wishbone_bd_ram_mem1_reg[188][11]/P0001 , \wishbone_bd_ram_mem1_reg[188][12]/P0001 , \wishbone_bd_ram_mem1_reg[188][13]/P0001 , \wishbone_bd_ram_mem1_reg[188][14]/P0001 , \wishbone_bd_ram_mem1_reg[188][15]/P0001 , \wishbone_bd_ram_mem1_reg[188][8]/P0001 , \wishbone_bd_ram_mem1_reg[188][9]/P0001 , \wishbone_bd_ram_mem1_reg[189][10]/P0001 , \wishbone_bd_ram_mem1_reg[189][11]/P0001 , \wishbone_bd_ram_mem1_reg[189][12]/P0001 , \wishbone_bd_ram_mem1_reg[189][13]/P0001 , \wishbone_bd_ram_mem1_reg[189][14]/P0001 , \wishbone_bd_ram_mem1_reg[189][15]/P0001 , \wishbone_bd_ram_mem1_reg[189][8]/P0001 , \wishbone_bd_ram_mem1_reg[189][9]/P0001 , \wishbone_bd_ram_mem1_reg[18][10]/P0001 , \wishbone_bd_ram_mem1_reg[18][11]/P0001 , \wishbone_bd_ram_mem1_reg[18][12]/P0001 , \wishbone_bd_ram_mem1_reg[18][13]/P0001 , \wishbone_bd_ram_mem1_reg[18][14]/P0001 , \wishbone_bd_ram_mem1_reg[18][15]/P0001 , \wishbone_bd_ram_mem1_reg[18][8]/P0001 , \wishbone_bd_ram_mem1_reg[18][9]/P0001 , \wishbone_bd_ram_mem1_reg[190][10]/P0001 , \wishbone_bd_ram_mem1_reg[190][11]/P0001 , \wishbone_bd_ram_mem1_reg[190][12]/P0001 , \wishbone_bd_ram_mem1_reg[190][13]/P0001 , \wishbone_bd_ram_mem1_reg[190][14]/P0001 , \wishbone_bd_ram_mem1_reg[190][15]/P0001 , \wishbone_bd_ram_mem1_reg[190][8]/P0001 , \wishbone_bd_ram_mem1_reg[190][9]/P0001 , \wishbone_bd_ram_mem1_reg[191][10]/P0001 , \wishbone_bd_ram_mem1_reg[191][11]/P0001 , \wishbone_bd_ram_mem1_reg[191][12]/P0001 , \wishbone_bd_ram_mem1_reg[191][13]/P0001 , \wishbone_bd_ram_mem1_reg[191][14]/P0001 , \wishbone_bd_ram_mem1_reg[191][15]/P0001 , \wishbone_bd_ram_mem1_reg[191][8]/P0001 , \wishbone_bd_ram_mem1_reg[191][9]/P0001 , \wishbone_bd_ram_mem1_reg[192][10]/P0001 , \wishbone_bd_ram_mem1_reg[192][11]/P0001 , \wishbone_bd_ram_mem1_reg[192][12]/P0001 , \wishbone_bd_ram_mem1_reg[192][13]/P0001 , \wishbone_bd_ram_mem1_reg[192][14]/P0001 , \wishbone_bd_ram_mem1_reg[192][15]/P0001 , \wishbone_bd_ram_mem1_reg[192][8]/P0001 , \wishbone_bd_ram_mem1_reg[192][9]/P0001 , \wishbone_bd_ram_mem1_reg[193][10]/P0001 , \wishbone_bd_ram_mem1_reg[193][11]/P0001 , \wishbone_bd_ram_mem1_reg[193][12]/P0001 , \wishbone_bd_ram_mem1_reg[193][13]/P0001 , \wishbone_bd_ram_mem1_reg[193][14]/P0001 , \wishbone_bd_ram_mem1_reg[193][15]/P0001 , \wishbone_bd_ram_mem1_reg[193][8]/P0001 , \wishbone_bd_ram_mem1_reg[193][9]/P0001 , \wishbone_bd_ram_mem1_reg[194][10]/P0001 , \wishbone_bd_ram_mem1_reg[194][11]/P0001 , \wishbone_bd_ram_mem1_reg[194][12]/P0001 , \wishbone_bd_ram_mem1_reg[194][13]/P0001 , \wishbone_bd_ram_mem1_reg[194][14]/P0001 , \wishbone_bd_ram_mem1_reg[194][15]/P0001 , \wishbone_bd_ram_mem1_reg[194][8]/P0001 , \wishbone_bd_ram_mem1_reg[194][9]/P0001 , \wishbone_bd_ram_mem1_reg[195][10]/P0001 , \wishbone_bd_ram_mem1_reg[195][11]/P0001 , \wishbone_bd_ram_mem1_reg[195][12]/P0001 , \wishbone_bd_ram_mem1_reg[195][13]/P0001 , \wishbone_bd_ram_mem1_reg[195][14]/P0001 , \wishbone_bd_ram_mem1_reg[195][15]/P0001 , \wishbone_bd_ram_mem1_reg[195][8]/P0001 , \wishbone_bd_ram_mem1_reg[195][9]/P0001 , \wishbone_bd_ram_mem1_reg[196][10]/P0001 , \wishbone_bd_ram_mem1_reg[196][11]/P0001 , \wishbone_bd_ram_mem1_reg[196][12]/P0001 , \wishbone_bd_ram_mem1_reg[196][13]/P0001 , \wishbone_bd_ram_mem1_reg[196][14]/P0001 , \wishbone_bd_ram_mem1_reg[196][15]/P0001 , \wishbone_bd_ram_mem1_reg[196][8]/P0001 , \wishbone_bd_ram_mem1_reg[196][9]/P0001 , \wishbone_bd_ram_mem1_reg[197][10]/P0001 , \wishbone_bd_ram_mem1_reg[197][11]/P0001 , \wishbone_bd_ram_mem1_reg[197][12]/P0001 , \wishbone_bd_ram_mem1_reg[197][13]/P0001 , \wishbone_bd_ram_mem1_reg[197][14]/P0001 , \wishbone_bd_ram_mem1_reg[197][15]/P0001 , \wishbone_bd_ram_mem1_reg[197][8]/P0001 , \wishbone_bd_ram_mem1_reg[197][9]/P0001 , \wishbone_bd_ram_mem1_reg[198][10]/P0001 , \wishbone_bd_ram_mem1_reg[198][11]/P0001 , \wishbone_bd_ram_mem1_reg[198][12]/P0001 , \wishbone_bd_ram_mem1_reg[198][13]/P0001 , \wishbone_bd_ram_mem1_reg[198][14]/P0001 , \wishbone_bd_ram_mem1_reg[198][15]/P0001 , \wishbone_bd_ram_mem1_reg[198][8]/P0001 , \wishbone_bd_ram_mem1_reg[198][9]/P0001 , \wishbone_bd_ram_mem1_reg[199][10]/P0001 , \wishbone_bd_ram_mem1_reg[199][11]/P0001 , \wishbone_bd_ram_mem1_reg[199][12]/P0001 , \wishbone_bd_ram_mem1_reg[199][13]/P0001 , \wishbone_bd_ram_mem1_reg[199][14]/P0001 , \wishbone_bd_ram_mem1_reg[199][15]/P0001 , \wishbone_bd_ram_mem1_reg[199][8]/P0001 , \wishbone_bd_ram_mem1_reg[199][9]/P0001 , \wishbone_bd_ram_mem1_reg[19][10]/P0001 , \wishbone_bd_ram_mem1_reg[19][11]/P0001 , \wishbone_bd_ram_mem1_reg[19][12]/P0001 , \wishbone_bd_ram_mem1_reg[19][13]/P0001 , \wishbone_bd_ram_mem1_reg[19][14]/P0001 , \wishbone_bd_ram_mem1_reg[19][15]/P0001 , \wishbone_bd_ram_mem1_reg[19][8]/P0001 , \wishbone_bd_ram_mem1_reg[19][9]/P0001 , \wishbone_bd_ram_mem1_reg[1][10]/P0001 , \wishbone_bd_ram_mem1_reg[1][11]/P0001 , \wishbone_bd_ram_mem1_reg[1][12]/P0001 , \wishbone_bd_ram_mem1_reg[1][13]/P0001 , \wishbone_bd_ram_mem1_reg[1][14]/P0001 , \wishbone_bd_ram_mem1_reg[1][15]/P0001 , \wishbone_bd_ram_mem1_reg[1][8]/P0001 , \wishbone_bd_ram_mem1_reg[1][9]/P0001 , \wishbone_bd_ram_mem1_reg[200][10]/P0001 , \wishbone_bd_ram_mem1_reg[200][11]/P0001 , \wishbone_bd_ram_mem1_reg[200][12]/P0001 , \wishbone_bd_ram_mem1_reg[200][13]/P0001 , \wishbone_bd_ram_mem1_reg[200][14]/P0001 , \wishbone_bd_ram_mem1_reg[200][15]/P0001 , \wishbone_bd_ram_mem1_reg[200][8]/P0001 , \wishbone_bd_ram_mem1_reg[200][9]/P0001 , \wishbone_bd_ram_mem1_reg[201][10]/P0001 , \wishbone_bd_ram_mem1_reg[201][11]/P0001 , \wishbone_bd_ram_mem1_reg[201][12]/P0001 , \wishbone_bd_ram_mem1_reg[201][13]/P0001 , \wishbone_bd_ram_mem1_reg[201][14]/P0001 , \wishbone_bd_ram_mem1_reg[201][15]/P0001 , \wishbone_bd_ram_mem1_reg[201][8]/P0001 , \wishbone_bd_ram_mem1_reg[201][9]/P0001 , \wishbone_bd_ram_mem1_reg[202][10]/P0001 , \wishbone_bd_ram_mem1_reg[202][11]/P0001 , \wishbone_bd_ram_mem1_reg[202][12]/P0001 , \wishbone_bd_ram_mem1_reg[202][13]/P0001 , \wishbone_bd_ram_mem1_reg[202][14]/P0001 , \wishbone_bd_ram_mem1_reg[202][15]/P0001 , \wishbone_bd_ram_mem1_reg[202][8]/P0001 , \wishbone_bd_ram_mem1_reg[202][9]/P0001 , \wishbone_bd_ram_mem1_reg[203][10]/P0001 , \wishbone_bd_ram_mem1_reg[203][11]/P0001 , \wishbone_bd_ram_mem1_reg[203][12]/P0001 , \wishbone_bd_ram_mem1_reg[203][13]/P0001 , \wishbone_bd_ram_mem1_reg[203][14]/P0001 , \wishbone_bd_ram_mem1_reg[203][15]/P0001 , \wishbone_bd_ram_mem1_reg[203][8]/P0001 , \wishbone_bd_ram_mem1_reg[203][9]/P0001 , \wishbone_bd_ram_mem1_reg[204][10]/P0001 , \wishbone_bd_ram_mem1_reg[204][11]/P0001 , \wishbone_bd_ram_mem1_reg[204][12]/P0001 , \wishbone_bd_ram_mem1_reg[204][13]/P0001 , \wishbone_bd_ram_mem1_reg[204][14]/P0001 , \wishbone_bd_ram_mem1_reg[204][15]/P0001 , \wishbone_bd_ram_mem1_reg[204][8]/P0001 , \wishbone_bd_ram_mem1_reg[204][9]/P0001 , \wishbone_bd_ram_mem1_reg[205][10]/P0001 , \wishbone_bd_ram_mem1_reg[205][11]/P0001 , \wishbone_bd_ram_mem1_reg[205][12]/P0001 , \wishbone_bd_ram_mem1_reg[205][13]/P0001 , \wishbone_bd_ram_mem1_reg[205][14]/P0001 , \wishbone_bd_ram_mem1_reg[205][15]/P0001 , \wishbone_bd_ram_mem1_reg[205][8]/P0001 , \wishbone_bd_ram_mem1_reg[205][9]/P0001 , \wishbone_bd_ram_mem1_reg[206][10]/P0001 , \wishbone_bd_ram_mem1_reg[206][11]/P0001 , \wishbone_bd_ram_mem1_reg[206][12]/P0001 , \wishbone_bd_ram_mem1_reg[206][13]/P0001 , \wishbone_bd_ram_mem1_reg[206][14]/P0001 , \wishbone_bd_ram_mem1_reg[206][15]/P0001 , \wishbone_bd_ram_mem1_reg[206][8]/P0001 , \wishbone_bd_ram_mem1_reg[206][9]/P0001 , \wishbone_bd_ram_mem1_reg[207][10]/P0001 , \wishbone_bd_ram_mem1_reg[207][11]/P0001 , \wishbone_bd_ram_mem1_reg[207][12]/P0001 , \wishbone_bd_ram_mem1_reg[207][13]/P0001 , \wishbone_bd_ram_mem1_reg[207][14]/P0001 , \wishbone_bd_ram_mem1_reg[207][15]/P0001 , \wishbone_bd_ram_mem1_reg[207][8]/P0001 , \wishbone_bd_ram_mem1_reg[207][9]/P0001 , \wishbone_bd_ram_mem1_reg[208][10]/P0001 , \wishbone_bd_ram_mem1_reg[208][11]/P0001 , \wishbone_bd_ram_mem1_reg[208][12]/P0001 , \wishbone_bd_ram_mem1_reg[208][13]/P0001 , \wishbone_bd_ram_mem1_reg[208][14]/P0001 , \wishbone_bd_ram_mem1_reg[208][15]/P0001 , \wishbone_bd_ram_mem1_reg[208][8]/P0001 , \wishbone_bd_ram_mem1_reg[208][9]/P0001 , \wishbone_bd_ram_mem1_reg[209][10]/P0001 , \wishbone_bd_ram_mem1_reg[209][11]/P0001 , \wishbone_bd_ram_mem1_reg[209][12]/P0001 , \wishbone_bd_ram_mem1_reg[209][13]/P0001 , \wishbone_bd_ram_mem1_reg[209][14]/P0001 , \wishbone_bd_ram_mem1_reg[209][15]/P0001 , \wishbone_bd_ram_mem1_reg[209][8]/P0001 , \wishbone_bd_ram_mem1_reg[209][9]/P0001 , \wishbone_bd_ram_mem1_reg[20][10]/P0001 , \wishbone_bd_ram_mem1_reg[20][11]/P0001 , \wishbone_bd_ram_mem1_reg[20][12]/P0001 , \wishbone_bd_ram_mem1_reg[20][13]/P0001 , \wishbone_bd_ram_mem1_reg[20][14]/P0001 , \wishbone_bd_ram_mem1_reg[20][15]/P0001 , \wishbone_bd_ram_mem1_reg[20][8]/P0001 , \wishbone_bd_ram_mem1_reg[20][9]/P0001 , \wishbone_bd_ram_mem1_reg[210][10]/P0001 , \wishbone_bd_ram_mem1_reg[210][11]/P0001 , \wishbone_bd_ram_mem1_reg[210][12]/P0001 , \wishbone_bd_ram_mem1_reg[210][13]/P0001 , \wishbone_bd_ram_mem1_reg[210][14]/P0001 , \wishbone_bd_ram_mem1_reg[210][15]/P0001 , \wishbone_bd_ram_mem1_reg[210][8]/P0001 , \wishbone_bd_ram_mem1_reg[210][9]/P0001 , \wishbone_bd_ram_mem1_reg[211][10]/P0001 , \wishbone_bd_ram_mem1_reg[211][11]/P0001 , \wishbone_bd_ram_mem1_reg[211][12]/P0001 , \wishbone_bd_ram_mem1_reg[211][13]/P0001 , \wishbone_bd_ram_mem1_reg[211][14]/P0001 , \wishbone_bd_ram_mem1_reg[211][15]/P0001 , \wishbone_bd_ram_mem1_reg[211][8]/P0001 , \wishbone_bd_ram_mem1_reg[211][9]/P0001 , \wishbone_bd_ram_mem1_reg[212][10]/P0001 , \wishbone_bd_ram_mem1_reg[212][11]/P0001 , \wishbone_bd_ram_mem1_reg[212][12]/P0001 , \wishbone_bd_ram_mem1_reg[212][13]/P0001 , \wishbone_bd_ram_mem1_reg[212][14]/P0001 , \wishbone_bd_ram_mem1_reg[212][15]/P0001 , \wishbone_bd_ram_mem1_reg[212][8]/P0001 , \wishbone_bd_ram_mem1_reg[212][9]/P0001 , \wishbone_bd_ram_mem1_reg[213][10]/P0001 , \wishbone_bd_ram_mem1_reg[213][11]/P0001 , \wishbone_bd_ram_mem1_reg[213][12]/P0001 , \wishbone_bd_ram_mem1_reg[213][13]/P0001 , \wishbone_bd_ram_mem1_reg[213][14]/P0001 , \wishbone_bd_ram_mem1_reg[213][15]/P0001 , \wishbone_bd_ram_mem1_reg[213][8]/P0001 , \wishbone_bd_ram_mem1_reg[213][9]/P0001 , \wishbone_bd_ram_mem1_reg[214][10]/P0001 , \wishbone_bd_ram_mem1_reg[214][11]/P0001 , \wishbone_bd_ram_mem1_reg[214][12]/P0001 , \wishbone_bd_ram_mem1_reg[214][13]/P0001 , \wishbone_bd_ram_mem1_reg[214][14]/P0001 , \wishbone_bd_ram_mem1_reg[214][15]/P0001 , \wishbone_bd_ram_mem1_reg[214][8]/P0001 , \wishbone_bd_ram_mem1_reg[214][9]/P0001 , \wishbone_bd_ram_mem1_reg[215][10]/P0001 , \wishbone_bd_ram_mem1_reg[215][11]/P0001 , \wishbone_bd_ram_mem1_reg[215][12]/P0001 , \wishbone_bd_ram_mem1_reg[215][13]/P0001 , \wishbone_bd_ram_mem1_reg[215][14]/P0001 , \wishbone_bd_ram_mem1_reg[215][15]/P0001 , \wishbone_bd_ram_mem1_reg[215][8]/P0001 , \wishbone_bd_ram_mem1_reg[215][9]/P0001 , \wishbone_bd_ram_mem1_reg[216][10]/P0001 , \wishbone_bd_ram_mem1_reg[216][11]/P0001 , \wishbone_bd_ram_mem1_reg[216][12]/P0001 , \wishbone_bd_ram_mem1_reg[216][13]/P0001 , \wishbone_bd_ram_mem1_reg[216][14]/P0001 , \wishbone_bd_ram_mem1_reg[216][15]/P0001 , \wishbone_bd_ram_mem1_reg[216][8]/P0001 , \wishbone_bd_ram_mem1_reg[216][9]/P0001 , \wishbone_bd_ram_mem1_reg[217][10]/P0001 , \wishbone_bd_ram_mem1_reg[217][11]/P0001 , \wishbone_bd_ram_mem1_reg[217][12]/P0001 , \wishbone_bd_ram_mem1_reg[217][13]/P0001 , \wishbone_bd_ram_mem1_reg[217][14]/P0001 , \wishbone_bd_ram_mem1_reg[217][15]/P0001 , \wishbone_bd_ram_mem1_reg[217][8]/P0001 , \wishbone_bd_ram_mem1_reg[217][9]/P0001 , \wishbone_bd_ram_mem1_reg[218][10]/P0001 , \wishbone_bd_ram_mem1_reg[218][11]/P0001 , \wishbone_bd_ram_mem1_reg[218][12]/P0001 , \wishbone_bd_ram_mem1_reg[218][13]/P0001 , \wishbone_bd_ram_mem1_reg[218][14]/P0001 , \wishbone_bd_ram_mem1_reg[218][15]/P0001 , \wishbone_bd_ram_mem1_reg[218][8]/P0001 , \wishbone_bd_ram_mem1_reg[218][9]/P0001 , \wishbone_bd_ram_mem1_reg[219][10]/P0001 , \wishbone_bd_ram_mem1_reg[219][11]/P0001 , \wishbone_bd_ram_mem1_reg[219][12]/P0001 , \wishbone_bd_ram_mem1_reg[219][13]/P0001 , \wishbone_bd_ram_mem1_reg[219][14]/P0001 , \wishbone_bd_ram_mem1_reg[219][15]/P0001 , \wishbone_bd_ram_mem1_reg[219][8]/P0001 , \wishbone_bd_ram_mem1_reg[219][9]/P0001 , \wishbone_bd_ram_mem1_reg[21][10]/P0001 , \wishbone_bd_ram_mem1_reg[21][11]/P0001 , \wishbone_bd_ram_mem1_reg[21][12]/P0001 , \wishbone_bd_ram_mem1_reg[21][13]/P0001 , \wishbone_bd_ram_mem1_reg[21][14]/P0001 , \wishbone_bd_ram_mem1_reg[21][15]/P0001 , \wishbone_bd_ram_mem1_reg[21][8]/P0001 , \wishbone_bd_ram_mem1_reg[21][9]/P0001 , \wishbone_bd_ram_mem1_reg[220][10]/P0001 , \wishbone_bd_ram_mem1_reg[220][11]/P0001 , \wishbone_bd_ram_mem1_reg[220][12]/P0001 , \wishbone_bd_ram_mem1_reg[220][13]/P0001 , \wishbone_bd_ram_mem1_reg[220][14]/P0001 , \wishbone_bd_ram_mem1_reg[220][15]/P0001 , \wishbone_bd_ram_mem1_reg[220][8]/P0001 , \wishbone_bd_ram_mem1_reg[220][9]/P0001 , \wishbone_bd_ram_mem1_reg[221][10]/P0001 , \wishbone_bd_ram_mem1_reg[221][11]/P0001 , \wishbone_bd_ram_mem1_reg[221][12]/P0001 , \wishbone_bd_ram_mem1_reg[221][13]/P0001 , \wishbone_bd_ram_mem1_reg[221][14]/P0001 , \wishbone_bd_ram_mem1_reg[221][15]/P0001 , \wishbone_bd_ram_mem1_reg[221][8]/P0001 , \wishbone_bd_ram_mem1_reg[221][9]/P0001 , \wishbone_bd_ram_mem1_reg[222][10]/P0001 , \wishbone_bd_ram_mem1_reg[222][11]/P0001 , \wishbone_bd_ram_mem1_reg[222][12]/P0001 , \wishbone_bd_ram_mem1_reg[222][13]/P0001 , \wishbone_bd_ram_mem1_reg[222][14]/P0001 , \wishbone_bd_ram_mem1_reg[222][15]/P0001 , \wishbone_bd_ram_mem1_reg[222][8]/P0001 , \wishbone_bd_ram_mem1_reg[222][9]/P0001 , \wishbone_bd_ram_mem1_reg[223][10]/P0001 , \wishbone_bd_ram_mem1_reg[223][11]/P0001 , \wishbone_bd_ram_mem1_reg[223][12]/P0001 , \wishbone_bd_ram_mem1_reg[223][13]/P0001 , \wishbone_bd_ram_mem1_reg[223][14]/P0001 , \wishbone_bd_ram_mem1_reg[223][15]/P0001 , \wishbone_bd_ram_mem1_reg[223][8]/P0001 , \wishbone_bd_ram_mem1_reg[223][9]/P0001 , \wishbone_bd_ram_mem1_reg[224][10]/P0001 , \wishbone_bd_ram_mem1_reg[224][11]/P0001 , \wishbone_bd_ram_mem1_reg[224][12]/P0001 , \wishbone_bd_ram_mem1_reg[224][13]/P0001 , \wishbone_bd_ram_mem1_reg[224][14]/P0001 , \wishbone_bd_ram_mem1_reg[224][15]/P0001 , \wishbone_bd_ram_mem1_reg[224][8]/P0001 , \wishbone_bd_ram_mem1_reg[224][9]/P0001 , \wishbone_bd_ram_mem1_reg[225][10]/P0001 , \wishbone_bd_ram_mem1_reg[225][11]/P0001 , \wishbone_bd_ram_mem1_reg[225][12]/P0001 , \wishbone_bd_ram_mem1_reg[225][13]/P0001 , \wishbone_bd_ram_mem1_reg[225][14]/P0001 , \wishbone_bd_ram_mem1_reg[225][15]/P0001 , \wishbone_bd_ram_mem1_reg[225][8]/P0001 , \wishbone_bd_ram_mem1_reg[225][9]/P0001 , \wishbone_bd_ram_mem1_reg[226][10]/P0001 , \wishbone_bd_ram_mem1_reg[226][11]/P0001 , \wishbone_bd_ram_mem1_reg[226][12]/P0001 , \wishbone_bd_ram_mem1_reg[226][13]/P0001 , \wishbone_bd_ram_mem1_reg[226][14]/P0001 , \wishbone_bd_ram_mem1_reg[226][15]/P0001 , \wishbone_bd_ram_mem1_reg[226][8]/P0001 , \wishbone_bd_ram_mem1_reg[226][9]/P0001 , \wishbone_bd_ram_mem1_reg[227][10]/P0001 , \wishbone_bd_ram_mem1_reg[227][11]/P0001 , \wishbone_bd_ram_mem1_reg[227][12]/P0001 , \wishbone_bd_ram_mem1_reg[227][13]/P0001 , \wishbone_bd_ram_mem1_reg[227][14]/P0001 , \wishbone_bd_ram_mem1_reg[227][15]/P0001 , \wishbone_bd_ram_mem1_reg[227][8]/P0001 , \wishbone_bd_ram_mem1_reg[227][9]/P0001 , \wishbone_bd_ram_mem1_reg[228][10]/P0001 , \wishbone_bd_ram_mem1_reg[228][11]/P0001 , \wishbone_bd_ram_mem1_reg[228][12]/P0001 , \wishbone_bd_ram_mem1_reg[228][13]/P0001 , \wishbone_bd_ram_mem1_reg[228][14]/P0001 , \wishbone_bd_ram_mem1_reg[228][15]/P0001 , \wishbone_bd_ram_mem1_reg[228][8]/P0001 , \wishbone_bd_ram_mem1_reg[228][9]/P0001 , \wishbone_bd_ram_mem1_reg[229][10]/P0001 , \wishbone_bd_ram_mem1_reg[229][11]/P0001 , \wishbone_bd_ram_mem1_reg[229][12]/P0001 , \wishbone_bd_ram_mem1_reg[229][13]/P0001 , \wishbone_bd_ram_mem1_reg[229][14]/P0001 , \wishbone_bd_ram_mem1_reg[229][15]/P0001 , \wishbone_bd_ram_mem1_reg[229][8]/P0001 , \wishbone_bd_ram_mem1_reg[229][9]/P0001 , \wishbone_bd_ram_mem1_reg[22][10]/P0001 , \wishbone_bd_ram_mem1_reg[22][11]/P0001 , \wishbone_bd_ram_mem1_reg[22][12]/P0001 , \wishbone_bd_ram_mem1_reg[22][13]/P0001 , \wishbone_bd_ram_mem1_reg[22][14]/P0001 , \wishbone_bd_ram_mem1_reg[22][15]/P0001 , \wishbone_bd_ram_mem1_reg[22][8]/P0001 , \wishbone_bd_ram_mem1_reg[22][9]/P0001 , \wishbone_bd_ram_mem1_reg[230][10]/P0001 , \wishbone_bd_ram_mem1_reg[230][11]/P0001 , \wishbone_bd_ram_mem1_reg[230][12]/P0001 , \wishbone_bd_ram_mem1_reg[230][13]/P0001 , \wishbone_bd_ram_mem1_reg[230][14]/P0001 , \wishbone_bd_ram_mem1_reg[230][15]/P0001 , \wishbone_bd_ram_mem1_reg[230][8]/P0001 , \wishbone_bd_ram_mem1_reg[230][9]/P0001 , \wishbone_bd_ram_mem1_reg[231][10]/P0001 , \wishbone_bd_ram_mem1_reg[231][11]/P0001 , \wishbone_bd_ram_mem1_reg[231][12]/P0001 , \wishbone_bd_ram_mem1_reg[231][13]/P0001 , \wishbone_bd_ram_mem1_reg[231][14]/P0001 , \wishbone_bd_ram_mem1_reg[231][15]/P0001 , \wishbone_bd_ram_mem1_reg[231][8]/P0001 , \wishbone_bd_ram_mem1_reg[231][9]/P0001 , \wishbone_bd_ram_mem1_reg[232][10]/P0001 , \wishbone_bd_ram_mem1_reg[232][11]/P0001 , \wishbone_bd_ram_mem1_reg[232][12]/P0001 , \wishbone_bd_ram_mem1_reg[232][13]/P0001 , \wishbone_bd_ram_mem1_reg[232][14]/P0001 , \wishbone_bd_ram_mem1_reg[232][15]/P0001 , \wishbone_bd_ram_mem1_reg[232][8]/P0001 , \wishbone_bd_ram_mem1_reg[232][9]/P0001 , \wishbone_bd_ram_mem1_reg[233][10]/P0001 , \wishbone_bd_ram_mem1_reg[233][11]/P0001 , \wishbone_bd_ram_mem1_reg[233][12]/P0001 , \wishbone_bd_ram_mem1_reg[233][13]/P0001 , \wishbone_bd_ram_mem1_reg[233][14]/P0001 , \wishbone_bd_ram_mem1_reg[233][15]/P0001 , \wishbone_bd_ram_mem1_reg[233][8]/P0001 , \wishbone_bd_ram_mem1_reg[233][9]/P0001 , \wishbone_bd_ram_mem1_reg[234][10]/P0001 , \wishbone_bd_ram_mem1_reg[234][11]/P0001 , \wishbone_bd_ram_mem1_reg[234][12]/P0001 , \wishbone_bd_ram_mem1_reg[234][13]/P0001 , \wishbone_bd_ram_mem1_reg[234][14]/P0001 , \wishbone_bd_ram_mem1_reg[234][15]/P0001 , \wishbone_bd_ram_mem1_reg[234][8]/P0001 , \wishbone_bd_ram_mem1_reg[234][9]/P0001 , \wishbone_bd_ram_mem1_reg[235][10]/P0001 , \wishbone_bd_ram_mem1_reg[235][11]/P0001 , \wishbone_bd_ram_mem1_reg[235][12]/P0001 , \wishbone_bd_ram_mem1_reg[235][13]/P0001 , \wishbone_bd_ram_mem1_reg[235][14]/P0001 , \wishbone_bd_ram_mem1_reg[235][15]/P0001 , \wishbone_bd_ram_mem1_reg[235][8]/P0001 , \wishbone_bd_ram_mem1_reg[235][9]/P0001 , \wishbone_bd_ram_mem1_reg[236][10]/P0001 , \wishbone_bd_ram_mem1_reg[236][11]/P0001 , \wishbone_bd_ram_mem1_reg[236][12]/P0001 , \wishbone_bd_ram_mem1_reg[236][13]/P0001 , \wishbone_bd_ram_mem1_reg[236][14]/P0001 , \wishbone_bd_ram_mem1_reg[236][15]/P0001 , \wishbone_bd_ram_mem1_reg[236][8]/P0001 , \wishbone_bd_ram_mem1_reg[236][9]/P0001 , \wishbone_bd_ram_mem1_reg[237][10]/P0001 , \wishbone_bd_ram_mem1_reg[237][11]/P0001 , \wishbone_bd_ram_mem1_reg[237][12]/P0001 , \wishbone_bd_ram_mem1_reg[237][13]/P0001 , \wishbone_bd_ram_mem1_reg[237][14]/P0001 , \wishbone_bd_ram_mem1_reg[237][15]/P0001 , \wishbone_bd_ram_mem1_reg[237][8]/P0001 , \wishbone_bd_ram_mem1_reg[237][9]/P0001 , \wishbone_bd_ram_mem1_reg[238][10]/P0001 , \wishbone_bd_ram_mem1_reg[238][11]/P0001 , \wishbone_bd_ram_mem1_reg[238][12]/P0001 , \wishbone_bd_ram_mem1_reg[238][13]/P0001 , \wishbone_bd_ram_mem1_reg[238][14]/P0001 , \wishbone_bd_ram_mem1_reg[238][15]/P0001 , \wishbone_bd_ram_mem1_reg[238][8]/P0001 , \wishbone_bd_ram_mem1_reg[238][9]/P0001 , \wishbone_bd_ram_mem1_reg[239][10]/P0001 , \wishbone_bd_ram_mem1_reg[239][11]/P0001 , \wishbone_bd_ram_mem1_reg[239][12]/P0001 , \wishbone_bd_ram_mem1_reg[239][13]/P0001 , \wishbone_bd_ram_mem1_reg[239][14]/P0001 , \wishbone_bd_ram_mem1_reg[239][15]/P0001 , \wishbone_bd_ram_mem1_reg[239][8]/P0001 , \wishbone_bd_ram_mem1_reg[239][9]/P0001 , \wishbone_bd_ram_mem1_reg[23][10]/P0001 , \wishbone_bd_ram_mem1_reg[23][11]/P0001 , \wishbone_bd_ram_mem1_reg[23][12]/P0001 , \wishbone_bd_ram_mem1_reg[23][13]/P0001 , \wishbone_bd_ram_mem1_reg[23][14]/P0001 , \wishbone_bd_ram_mem1_reg[23][15]/P0001 , \wishbone_bd_ram_mem1_reg[23][8]/P0001 , \wishbone_bd_ram_mem1_reg[23][9]/P0001 , \wishbone_bd_ram_mem1_reg[240][10]/P0001 , \wishbone_bd_ram_mem1_reg[240][11]/P0001 , \wishbone_bd_ram_mem1_reg[240][12]/P0001 , \wishbone_bd_ram_mem1_reg[240][13]/P0001 , \wishbone_bd_ram_mem1_reg[240][14]/P0001 , \wishbone_bd_ram_mem1_reg[240][15]/P0001 , \wishbone_bd_ram_mem1_reg[240][8]/P0001 , \wishbone_bd_ram_mem1_reg[240][9]/P0001 , \wishbone_bd_ram_mem1_reg[241][10]/P0001 , \wishbone_bd_ram_mem1_reg[241][11]/P0001 , \wishbone_bd_ram_mem1_reg[241][12]/P0001 , \wishbone_bd_ram_mem1_reg[241][13]/P0001 , \wishbone_bd_ram_mem1_reg[241][14]/P0001 , \wishbone_bd_ram_mem1_reg[241][15]/P0001 , \wishbone_bd_ram_mem1_reg[241][8]/P0001 , \wishbone_bd_ram_mem1_reg[241][9]/P0001 , \wishbone_bd_ram_mem1_reg[242][10]/P0001 , \wishbone_bd_ram_mem1_reg[242][11]/P0001 , \wishbone_bd_ram_mem1_reg[242][12]/P0001 , \wishbone_bd_ram_mem1_reg[242][13]/P0001 , \wishbone_bd_ram_mem1_reg[242][14]/P0001 , \wishbone_bd_ram_mem1_reg[242][15]/P0001 , \wishbone_bd_ram_mem1_reg[242][8]/P0001 , \wishbone_bd_ram_mem1_reg[242][9]/P0001 , \wishbone_bd_ram_mem1_reg[243][10]/P0001 , \wishbone_bd_ram_mem1_reg[243][11]/P0001 , \wishbone_bd_ram_mem1_reg[243][12]/P0001 , \wishbone_bd_ram_mem1_reg[243][13]/P0001 , \wishbone_bd_ram_mem1_reg[243][14]/P0001 , \wishbone_bd_ram_mem1_reg[243][15]/P0001 , \wishbone_bd_ram_mem1_reg[243][8]/P0001 , \wishbone_bd_ram_mem1_reg[243][9]/P0001 , \wishbone_bd_ram_mem1_reg[244][10]/P0001 , \wishbone_bd_ram_mem1_reg[244][11]/P0001 , \wishbone_bd_ram_mem1_reg[244][12]/P0001 , \wishbone_bd_ram_mem1_reg[244][13]/P0001 , \wishbone_bd_ram_mem1_reg[244][14]/P0001 , \wishbone_bd_ram_mem1_reg[244][15]/P0001 , \wishbone_bd_ram_mem1_reg[244][8]/P0001 , \wishbone_bd_ram_mem1_reg[244][9]/P0001 , \wishbone_bd_ram_mem1_reg[245][10]/P0001 , \wishbone_bd_ram_mem1_reg[245][11]/P0001 , \wishbone_bd_ram_mem1_reg[245][12]/P0001 , \wishbone_bd_ram_mem1_reg[245][13]/P0001 , \wishbone_bd_ram_mem1_reg[245][14]/P0001 , \wishbone_bd_ram_mem1_reg[245][15]/P0001 , \wishbone_bd_ram_mem1_reg[245][8]/P0001 , \wishbone_bd_ram_mem1_reg[245][9]/P0001 , \wishbone_bd_ram_mem1_reg[246][10]/P0001 , \wishbone_bd_ram_mem1_reg[246][11]/P0001 , \wishbone_bd_ram_mem1_reg[246][12]/P0001 , \wishbone_bd_ram_mem1_reg[246][13]/P0001 , \wishbone_bd_ram_mem1_reg[246][14]/P0001 , \wishbone_bd_ram_mem1_reg[246][15]/P0001 , \wishbone_bd_ram_mem1_reg[246][8]/P0001 , \wishbone_bd_ram_mem1_reg[246][9]/P0001 , \wishbone_bd_ram_mem1_reg[247][10]/P0001 , \wishbone_bd_ram_mem1_reg[247][11]/P0001 , \wishbone_bd_ram_mem1_reg[247][12]/P0001 , \wishbone_bd_ram_mem1_reg[247][13]/P0001 , \wishbone_bd_ram_mem1_reg[247][14]/P0001 , \wishbone_bd_ram_mem1_reg[247][15]/P0001 , \wishbone_bd_ram_mem1_reg[247][8]/P0001 , \wishbone_bd_ram_mem1_reg[247][9]/P0001 , \wishbone_bd_ram_mem1_reg[248][10]/P0001 , \wishbone_bd_ram_mem1_reg[248][11]/P0001 , \wishbone_bd_ram_mem1_reg[248][12]/P0001 , \wishbone_bd_ram_mem1_reg[248][13]/P0001 , \wishbone_bd_ram_mem1_reg[248][14]/P0001 , \wishbone_bd_ram_mem1_reg[248][15]/P0001 , \wishbone_bd_ram_mem1_reg[248][8]/P0001 , \wishbone_bd_ram_mem1_reg[248][9]/P0001 , \wishbone_bd_ram_mem1_reg[249][10]/P0001 , \wishbone_bd_ram_mem1_reg[249][11]/P0001 , \wishbone_bd_ram_mem1_reg[249][12]/P0001 , \wishbone_bd_ram_mem1_reg[249][13]/P0001 , \wishbone_bd_ram_mem1_reg[249][14]/P0001 , \wishbone_bd_ram_mem1_reg[249][15]/P0001 , \wishbone_bd_ram_mem1_reg[249][8]/P0001 , \wishbone_bd_ram_mem1_reg[249][9]/P0001 , \wishbone_bd_ram_mem1_reg[24][10]/P0001 , \wishbone_bd_ram_mem1_reg[24][11]/P0001 , \wishbone_bd_ram_mem1_reg[24][12]/P0001 , \wishbone_bd_ram_mem1_reg[24][13]/P0001 , \wishbone_bd_ram_mem1_reg[24][14]/P0001 , \wishbone_bd_ram_mem1_reg[24][15]/P0001 , \wishbone_bd_ram_mem1_reg[24][8]/P0001 , \wishbone_bd_ram_mem1_reg[24][9]/P0001 , \wishbone_bd_ram_mem1_reg[250][10]/P0001 , \wishbone_bd_ram_mem1_reg[250][11]/P0001 , \wishbone_bd_ram_mem1_reg[250][12]/P0001 , \wishbone_bd_ram_mem1_reg[250][13]/P0001 , \wishbone_bd_ram_mem1_reg[250][14]/P0001 , \wishbone_bd_ram_mem1_reg[250][15]/P0001 , \wishbone_bd_ram_mem1_reg[250][8]/P0001 , \wishbone_bd_ram_mem1_reg[250][9]/P0001 , \wishbone_bd_ram_mem1_reg[251][10]/P0001 , \wishbone_bd_ram_mem1_reg[251][11]/P0001 , \wishbone_bd_ram_mem1_reg[251][12]/P0001 , \wishbone_bd_ram_mem1_reg[251][13]/P0001 , \wishbone_bd_ram_mem1_reg[251][14]/P0001 , \wishbone_bd_ram_mem1_reg[251][15]/P0001 , \wishbone_bd_ram_mem1_reg[251][8]/P0001 , \wishbone_bd_ram_mem1_reg[251][9]/P0001 , \wishbone_bd_ram_mem1_reg[252][10]/P0001 , \wishbone_bd_ram_mem1_reg[252][11]/P0001 , \wishbone_bd_ram_mem1_reg[252][12]/P0001 , \wishbone_bd_ram_mem1_reg[252][13]/P0001 , \wishbone_bd_ram_mem1_reg[252][14]/P0001 , \wishbone_bd_ram_mem1_reg[252][15]/P0001 , \wishbone_bd_ram_mem1_reg[252][8]/P0001 , \wishbone_bd_ram_mem1_reg[252][9]/P0001 , \wishbone_bd_ram_mem1_reg[253][10]/P0001 , \wishbone_bd_ram_mem1_reg[253][11]/P0001 , \wishbone_bd_ram_mem1_reg[253][12]/P0001 , \wishbone_bd_ram_mem1_reg[253][13]/P0001 , \wishbone_bd_ram_mem1_reg[253][14]/P0001 , \wishbone_bd_ram_mem1_reg[253][15]/P0001 , \wishbone_bd_ram_mem1_reg[253][8]/P0001 , \wishbone_bd_ram_mem1_reg[253][9]/P0001 , \wishbone_bd_ram_mem1_reg[254][10]/P0001 , \wishbone_bd_ram_mem1_reg[254][11]/P0001 , \wishbone_bd_ram_mem1_reg[254][12]/P0001 , \wishbone_bd_ram_mem1_reg[254][13]/P0001 , \wishbone_bd_ram_mem1_reg[254][14]/P0001 , \wishbone_bd_ram_mem1_reg[254][15]/P0001 , \wishbone_bd_ram_mem1_reg[254][8]/P0001 , \wishbone_bd_ram_mem1_reg[254][9]/P0001 , \wishbone_bd_ram_mem1_reg[255][10]/P0001 , \wishbone_bd_ram_mem1_reg[255][11]/P0001 , \wishbone_bd_ram_mem1_reg[255][12]/P0001 , \wishbone_bd_ram_mem1_reg[255][13]/P0001 , \wishbone_bd_ram_mem1_reg[255][14]/P0001 , \wishbone_bd_ram_mem1_reg[255][15]/P0001 , \wishbone_bd_ram_mem1_reg[255][8]/P0001 , \wishbone_bd_ram_mem1_reg[255][9]/P0001 , \wishbone_bd_ram_mem1_reg[25][10]/P0001 , \wishbone_bd_ram_mem1_reg[25][11]/P0001 , \wishbone_bd_ram_mem1_reg[25][12]/P0001 , \wishbone_bd_ram_mem1_reg[25][13]/P0001 , \wishbone_bd_ram_mem1_reg[25][14]/P0001 , \wishbone_bd_ram_mem1_reg[25][15]/P0001 , \wishbone_bd_ram_mem1_reg[25][8]/P0001 , \wishbone_bd_ram_mem1_reg[25][9]/P0001 , \wishbone_bd_ram_mem1_reg[26][10]/P0001 , \wishbone_bd_ram_mem1_reg[26][11]/P0001 , \wishbone_bd_ram_mem1_reg[26][12]/P0001 , \wishbone_bd_ram_mem1_reg[26][13]/P0001 , \wishbone_bd_ram_mem1_reg[26][14]/P0001 , \wishbone_bd_ram_mem1_reg[26][15]/P0001 , \wishbone_bd_ram_mem1_reg[26][8]/P0001 , \wishbone_bd_ram_mem1_reg[26][9]/P0001 , \wishbone_bd_ram_mem1_reg[27][10]/P0001 , \wishbone_bd_ram_mem1_reg[27][11]/P0001 , \wishbone_bd_ram_mem1_reg[27][12]/P0001 , \wishbone_bd_ram_mem1_reg[27][13]/P0001 , \wishbone_bd_ram_mem1_reg[27][14]/P0001 , \wishbone_bd_ram_mem1_reg[27][15]/P0001 , \wishbone_bd_ram_mem1_reg[27][8]/P0001 , \wishbone_bd_ram_mem1_reg[27][9]/P0001 , \wishbone_bd_ram_mem1_reg[28][10]/P0001 , \wishbone_bd_ram_mem1_reg[28][11]/P0001 , \wishbone_bd_ram_mem1_reg[28][12]/P0001 , \wishbone_bd_ram_mem1_reg[28][13]/P0001 , \wishbone_bd_ram_mem1_reg[28][14]/P0001 , \wishbone_bd_ram_mem1_reg[28][15]/P0001 , \wishbone_bd_ram_mem1_reg[28][8]/P0001 , \wishbone_bd_ram_mem1_reg[28][9]/P0001 , \wishbone_bd_ram_mem1_reg[29][10]/P0001 , \wishbone_bd_ram_mem1_reg[29][11]/P0001 , \wishbone_bd_ram_mem1_reg[29][12]/P0001 , \wishbone_bd_ram_mem1_reg[29][13]/P0001 , \wishbone_bd_ram_mem1_reg[29][14]/P0001 , \wishbone_bd_ram_mem1_reg[29][15]/P0001 , \wishbone_bd_ram_mem1_reg[29][8]/P0001 , \wishbone_bd_ram_mem1_reg[29][9]/P0001 , \wishbone_bd_ram_mem1_reg[2][10]/P0001 , \wishbone_bd_ram_mem1_reg[2][11]/P0001 , \wishbone_bd_ram_mem1_reg[2][12]/P0001 , \wishbone_bd_ram_mem1_reg[2][13]/P0001 , \wishbone_bd_ram_mem1_reg[2][14]/P0001 , \wishbone_bd_ram_mem1_reg[2][15]/P0001 , \wishbone_bd_ram_mem1_reg[2][8]/P0001 , \wishbone_bd_ram_mem1_reg[2][9]/P0001 , \wishbone_bd_ram_mem1_reg[30][10]/P0001 , \wishbone_bd_ram_mem1_reg[30][11]/P0001 , \wishbone_bd_ram_mem1_reg[30][12]/P0001 , \wishbone_bd_ram_mem1_reg[30][13]/P0001 , \wishbone_bd_ram_mem1_reg[30][14]/P0001 , \wishbone_bd_ram_mem1_reg[30][15]/P0001 , \wishbone_bd_ram_mem1_reg[30][8]/P0001 , \wishbone_bd_ram_mem1_reg[30][9]/P0001 , \wishbone_bd_ram_mem1_reg[31][10]/P0001 , \wishbone_bd_ram_mem1_reg[31][11]/P0001 , \wishbone_bd_ram_mem1_reg[31][12]/P0001 , \wishbone_bd_ram_mem1_reg[31][13]/P0001 , \wishbone_bd_ram_mem1_reg[31][14]/P0001 , \wishbone_bd_ram_mem1_reg[31][15]/P0001 , \wishbone_bd_ram_mem1_reg[31][8]/P0001 , \wishbone_bd_ram_mem1_reg[31][9]/P0001 , \wishbone_bd_ram_mem1_reg[32][10]/P0001 , \wishbone_bd_ram_mem1_reg[32][11]/P0001 , \wishbone_bd_ram_mem1_reg[32][12]/P0001 , \wishbone_bd_ram_mem1_reg[32][13]/P0001 , \wishbone_bd_ram_mem1_reg[32][14]/P0001 , \wishbone_bd_ram_mem1_reg[32][15]/P0001 , \wishbone_bd_ram_mem1_reg[32][8]/P0001 , \wishbone_bd_ram_mem1_reg[32][9]/P0001 , \wishbone_bd_ram_mem1_reg[33][10]/P0001 , \wishbone_bd_ram_mem1_reg[33][11]/P0001 , \wishbone_bd_ram_mem1_reg[33][12]/P0001 , \wishbone_bd_ram_mem1_reg[33][13]/P0001 , \wishbone_bd_ram_mem1_reg[33][14]/P0001 , \wishbone_bd_ram_mem1_reg[33][15]/P0001 , \wishbone_bd_ram_mem1_reg[33][8]/P0001 , \wishbone_bd_ram_mem1_reg[33][9]/P0001 , \wishbone_bd_ram_mem1_reg[34][10]/P0001 , \wishbone_bd_ram_mem1_reg[34][11]/P0001 , \wishbone_bd_ram_mem1_reg[34][12]/P0001 , \wishbone_bd_ram_mem1_reg[34][13]/P0001 , \wishbone_bd_ram_mem1_reg[34][14]/P0001 , \wishbone_bd_ram_mem1_reg[34][15]/P0001 , \wishbone_bd_ram_mem1_reg[34][8]/P0001 , \wishbone_bd_ram_mem1_reg[34][9]/P0001 , \wishbone_bd_ram_mem1_reg[35][10]/P0001 , \wishbone_bd_ram_mem1_reg[35][11]/P0001 , \wishbone_bd_ram_mem1_reg[35][12]/P0001 , \wishbone_bd_ram_mem1_reg[35][13]/P0001 , \wishbone_bd_ram_mem1_reg[35][14]/P0001 , \wishbone_bd_ram_mem1_reg[35][15]/P0001 , \wishbone_bd_ram_mem1_reg[35][8]/P0001 , \wishbone_bd_ram_mem1_reg[35][9]/P0001 , \wishbone_bd_ram_mem1_reg[36][10]/P0001 , \wishbone_bd_ram_mem1_reg[36][11]/P0001 , \wishbone_bd_ram_mem1_reg[36][12]/P0001 , \wishbone_bd_ram_mem1_reg[36][13]/P0001 , \wishbone_bd_ram_mem1_reg[36][14]/P0001 , \wishbone_bd_ram_mem1_reg[36][15]/P0001 , \wishbone_bd_ram_mem1_reg[36][8]/P0001 , \wishbone_bd_ram_mem1_reg[36][9]/P0001 , \wishbone_bd_ram_mem1_reg[37][10]/P0001 , \wishbone_bd_ram_mem1_reg[37][11]/P0001 , \wishbone_bd_ram_mem1_reg[37][12]/P0001 , \wishbone_bd_ram_mem1_reg[37][13]/P0001 , \wishbone_bd_ram_mem1_reg[37][14]/P0001 , \wishbone_bd_ram_mem1_reg[37][15]/P0001 , \wishbone_bd_ram_mem1_reg[37][8]/P0001 , \wishbone_bd_ram_mem1_reg[37][9]/P0001 , \wishbone_bd_ram_mem1_reg[38][10]/P0001 , \wishbone_bd_ram_mem1_reg[38][11]/P0001 , \wishbone_bd_ram_mem1_reg[38][12]/P0001 , \wishbone_bd_ram_mem1_reg[38][13]/P0001 , \wishbone_bd_ram_mem1_reg[38][14]/P0001 , \wishbone_bd_ram_mem1_reg[38][15]/P0001 , \wishbone_bd_ram_mem1_reg[38][8]/P0001 , \wishbone_bd_ram_mem1_reg[38][9]/P0001 , \wishbone_bd_ram_mem1_reg[39][10]/P0001 , \wishbone_bd_ram_mem1_reg[39][11]/P0001 , \wishbone_bd_ram_mem1_reg[39][12]/P0001 , \wishbone_bd_ram_mem1_reg[39][13]/P0001 , \wishbone_bd_ram_mem1_reg[39][14]/P0001 , \wishbone_bd_ram_mem1_reg[39][15]/P0001 , \wishbone_bd_ram_mem1_reg[39][8]/P0001 , \wishbone_bd_ram_mem1_reg[39][9]/P0001 , \wishbone_bd_ram_mem1_reg[3][10]/P0001 , \wishbone_bd_ram_mem1_reg[3][11]/P0001 , \wishbone_bd_ram_mem1_reg[3][12]/P0001 , \wishbone_bd_ram_mem1_reg[3][13]/P0001 , \wishbone_bd_ram_mem1_reg[3][14]/P0001 , \wishbone_bd_ram_mem1_reg[3][15]/P0001 , \wishbone_bd_ram_mem1_reg[3][8]/P0001 , \wishbone_bd_ram_mem1_reg[3][9]/P0001 , \wishbone_bd_ram_mem1_reg[40][10]/P0001 , \wishbone_bd_ram_mem1_reg[40][11]/P0001 , \wishbone_bd_ram_mem1_reg[40][12]/P0001 , \wishbone_bd_ram_mem1_reg[40][13]/P0001 , \wishbone_bd_ram_mem1_reg[40][14]/P0001 , \wishbone_bd_ram_mem1_reg[40][15]/P0001 , \wishbone_bd_ram_mem1_reg[40][8]/P0001 , \wishbone_bd_ram_mem1_reg[40][9]/P0001 , \wishbone_bd_ram_mem1_reg[41][10]/P0001 , \wishbone_bd_ram_mem1_reg[41][11]/P0001 , \wishbone_bd_ram_mem1_reg[41][12]/P0001 , \wishbone_bd_ram_mem1_reg[41][13]/P0001 , \wishbone_bd_ram_mem1_reg[41][14]/P0001 , \wishbone_bd_ram_mem1_reg[41][15]/P0001 , \wishbone_bd_ram_mem1_reg[41][8]/P0001 , \wishbone_bd_ram_mem1_reg[41][9]/P0001 , \wishbone_bd_ram_mem1_reg[42][10]/P0001 , \wishbone_bd_ram_mem1_reg[42][11]/P0001 , \wishbone_bd_ram_mem1_reg[42][12]/P0001 , \wishbone_bd_ram_mem1_reg[42][13]/P0001 , \wishbone_bd_ram_mem1_reg[42][14]/P0001 , \wishbone_bd_ram_mem1_reg[42][15]/P0001 , \wishbone_bd_ram_mem1_reg[42][8]/P0001 , \wishbone_bd_ram_mem1_reg[42][9]/P0001 , \wishbone_bd_ram_mem1_reg[43][10]/P0001 , \wishbone_bd_ram_mem1_reg[43][11]/P0001 , \wishbone_bd_ram_mem1_reg[43][12]/P0001 , \wishbone_bd_ram_mem1_reg[43][13]/P0001 , \wishbone_bd_ram_mem1_reg[43][14]/P0001 , \wishbone_bd_ram_mem1_reg[43][15]/P0001 , \wishbone_bd_ram_mem1_reg[43][8]/P0001 , \wishbone_bd_ram_mem1_reg[43][9]/P0001 , \wishbone_bd_ram_mem1_reg[44][10]/P0001 , \wishbone_bd_ram_mem1_reg[44][11]/P0001 , \wishbone_bd_ram_mem1_reg[44][12]/P0001 , \wishbone_bd_ram_mem1_reg[44][13]/P0001 , \wishbone_bd_ram_mem1_reg[44][14]/P0001 , \wishbone_bd_ram_mem1_reg[44][15]/P0001 , \wishbone_bd_ram_mem1_reg[44][8]/P0001 , \wishbone_bd_ram_mem1_reg[44][9]/P0001 , \wishbone_bd_ram_mem1_reg[45][10]/P0001 , \wishbone_bd_ram_mem1_reg[45][11]/P0001 , \wishbone_bd_ram_mem1_reg[45][12]/P0001 , \wishbone_bd_ram_mem1_reg[45][13]/P0001 , \wishbone_bd_ram_mem1_reg[45][14]/P0001 , \wishbone_bd_ram_mem1_reg[45][15]/P0001 , \wishbone_bd_ram_mem1_reg[45][8]/P0001 , \wishbone_bd_ram_mem1_reg[45][9]/P0001 , \wishbone_bd_ram_mem1_reg[46][10]/P0001 , \wishbone_bd_ram_mem1_reg[46][11]/P0001 , \wishbone_bd_ram_mem1_reg[46][12]/P0001 , \wishbone_bd_ram_mem1_reg[46][13]/P0001 , \wishbone_bd_ram_mem1_reg[46][14]/P0001 , \wishbone_bd_ram_mem1_reg[46][15]/P0001 , \wishbone_bd_ram_mem1_reg[46][8]/P0001 , \wishbone_bd_ram_mem1_reg[46][9]/P0001 , \wishbone_bd_ram_mem1_reg[47][10]/P0001 , \wishbone_bd_ram_mem1_reg[47][11]/P0001 , \wishbone_bd_ram_mem1_reg[47][12]/P0001 , \wishbone_bd_ram_mem1_reg[47][13]/P0001 , \wishbone_bd_ram_mem1_reg[47][14]/P0001 , \wishbone_bd_ram_mem1_reg[47][15]/P0001 , \wishbone_bd_ram_mem1_reg[47][8]/P0001 , \wishbone_bd_ram_mem1_reg[47][9]/P0001 , \wishbone_bd_ram_mem1_reg[48][10]/P0001 , \wishbone_bd_ram_mem1_reg[48][11]/P0001 , \wishbone_bd_ram_mem1_reg[48][12]/P0001 , \wishbone_bd_ram_mem1_reg[48][13]/P0001 , \wishbone_bd_ram_mem1_reg[48][14]/P0001 , \wishbone_bd_ram_mem1_reg[48][15]/P0001 , \wishbone_bd_ram_mem1_reg[48][8]/P0001 , \wishbone_bd_ram_mem1_reg[48][9]/P0001 , \wishbone_bd_ram_mem1_reg[49][10]/P0001 , \wishbone_bd_ram_mem1_reg[49][11]/P0001 , \wishbone_bd_ram_mem1_reg[49][12]/P0001 , \wishbone_bd_ram_mem1_reg[49][13]/P0001 , \wishbone_bd_ram_mem1_reg[49][14]/P0001 , \wishbone_bd_ram_mem1_reg[49][15]/P0001 , \wishbone_bd_ram_mem1_reg[49][8]/P0001 , \wishbone_bd_ram_mem1_reg[49][9]/P0001 , \wishbone_bd_ram_mem1_reg[4][10]/P0001 , \wishbone_bd_ram_mem1_reg[4][11]/P0001 , \wishbone_bd_ram_mem1_reg[4][12]/P0001 , \wishbone_bd_ram_mem1_reg[4][13]/P0001 , \wishbone_bd_ram_mem1_reg[4][14]/P0001 , \wishbone_bd_ram_mem1_reg[4][15]/P0001 , \wishbone_bd_ram_mem1_reg[4][8]/P0001 , \wishbone_bd_ram_mem1_reg[4][9]/P0001 , \wishbone_bd_ram_mem1_reg[50][10]/P0001 , \wishbone_bd_ram_mem1_reg[50][11]/P0001 , \wishbone_bd_ram_mem1_reg[50][12]/P0001 , \wishbone_bd_ram_mem1_reg[50][13]/P0001 , \wishbone_bd_ram_mem1_reg[50][14]/P0001 , \wishbone_bd_ram_mem1_reg[50][15]/P0001 , \wishbone_bd_ram_mem1_reg[50][8]/P0001 , \wishbone_bd_ram_mem1_reg[50][9]/P0001 , \wishbone_bd_ram_mem1_reg[51][10]/P0001 , \wishbone_bd_ram_mem1_reg[51][11]/P0001 , \wishbone_bd_ram_mem1_reg[51][12]/P0001 , \wishbone_bd_ram_mem1_reg[51][13]/P0001 , \wishbone_bd_ram_mem1_reg[51][14]/P0001 , \wishbone_bd_ram_mem1_reg[51][15]/P0001 , \wishbone_bd_ram_mem1_reg[51][8]/P0001 , \wishbone_bd_ram_mem1_reg[51][9]/P0001 , \wishbone_bd_ram_mem1_reg[52][10]/P0001 , \wishbone_bd_ram_mem1_reg[52][11]/P0001 , \wishbone_bd_ram_mem1_reg[52][12]/P0001 , \wishbone_bd_ram_mem1_reg[52][13]/P0001 , \wishbone_bd_ram_mem1_reg[52][14]/P0001 , \wishbone_bd_ram_mem1_reg[52][15]/P0001 , \wishbone_bd_ram_mem1_reg[52][8]/P0001 , \wishbone_bd_ram_mem1_reg[52][9]/P0001 , \wishbone_bd_ram_mem1_reg[53][10]/P0001 , \wishbone_bd_ram_mem1_reg[53][11]/P0001 , \wishbone_bd_ram_mem1_reg[53][12]/P0001 , \wishbone_bd_ram_mem1_reg[53][13]/P0001 , \wishbone_bd_ram_mem1_reg[53][14]/P0001 , \wishbone_bd_ram_mem1_reg[53][15]/P0001 , \wishbone_bd_ram_mem1_reg[53][8]/P0001 , \wishbone_bd_ram_mem1_reg[53][9]/P0001 , \wishbone_bd_ram_mem1_reg[54][10]/P0001 , \wishbone_bd_ram_mem1_reg[54][11]/P0001 , \wishbone_bd_ram_mem1_reg[54][12]/P0001 , \wishbone_bd_ram_mem1_reg[54][13]/P0001 , \wishbone_bd_ram_mem1_reg[54][14]/P0001 , \wishbone_bd_ram_mem1_reg[54][15]/P0001 , \wishbone_bd_ram_mem1_reg[54][8]/P0001 , \wishbone_bd_ram_mem1_reg[54][9]/P0001 , \wishbone_bd_ram_mem1_reg[55][10]/P0001 , \wishbone_bd_ram_mem1_reg[55][11]/P0001 , \wishbone_bd_ram_mem1_reg[55][12]/P0001 , \wishbone_bd_ram_mem1_reg[55][13]/P0001 , \wishbone_bd_ram_mem1_reg[55][14]/P0001 , \wishbone_bd_ram_mem1_reg[55][15]/P0001 , \wishbone_bd_ram_mem1_reg[55][8]/P0001 , \wishbone_bd_ram_mem1_reg[55][9]/P0001 , \wishbone_bd_ram_mem1_reg[56][10]/P0001 , \wishbone_bd_ram_mem1_reg[56][11]/P0001 , \wishbone_bd_ram_mem1_reg[56][12]/P0001 , \wishbone_bd_ram_mem1_reg[56][13]/P0001 , \wishbone_bd_ram_mem1_reg[56][14]/P0001 , \wishbone_bd_ram_mem1_reg[56][15]/P0001 , \wishbone_bd_ram_mem1_reg[56][8]/P0001 , \wishbone_bd_ram_mem1_reg[56][9]/P0001 , \wishbone_bd_ram_mem1_reg[57][10]/P0001 , \wishbone_bd_ram_mem1_reg[57][11]/P0001 , \wishbone_bd_ram_mem1_reg[57][12]/P0001 , \wishbone_bd_ram_mem1_reg[57][13]/P0001 , \wishbone_bd_ram_mem1_reg[57][14]/P0001 , \wishbone_bd_ram_mem1_reg[57][15]/P0001 , \wishbone_bd_ram_mem1_reg[57][8]/P0001 , \wishbone_bd_ram_mem1_reg[57][9]/P0001 , \wishbone_bd_ram_mem1_reg[58][10]/P0001 , \wishbone_bd_ram_mem1_reg[58][11]/P0001 , \wishbone_bd_ram_mem1_reg[58][12]/P0001 , \wishbone_bd_ram_mem1_reg[58][13]/P0001 , \wishbone_bd_ram_mem1_reg[58][14]/P0001 , \wishbone_bd_ram_mem1_reg[58][15]/P0001 , \wishbone_bd_ram_mem1_reg[58][8]/P0001 , \wishbone_bd_ram_mem1_reg[58][9]/P0001 , \wishbone_bd_ram_mem1_reg[59][10]/P0001 , \wishbone_bd_ram_mem1_reg[59][11]/P0001 , \wishbone_bd_ram_mem1_reg[59][12]/P0001 , \wishbone_bd_ram_mem1_reg[59][13]/P0001 , \wishbone_bd_ram_mem1_reg[59][14]/P0001 , \wishbone_bd_ram_mem1_reg[59][15]/P0001 , \wishbone_bd_ram_mem1_reg[59][8]/P0001 , \wishbone_bd_ram_mem1_reg[59][9]/P0001 , \wishbone_bd_ram_mem1_reg[5][10]/P0001 , \wishbone_bd_ram_mem1_reg[5][11]/P0001 , \wishbone_bd_ram_mem1_reg[5][12]/P0001 , \wishbone_bd_ram_mem1_reg[5][13]/P0001 , \wishbone_bd_ram_mem1_reg[5][14]/P0001 , \wishbone_bd_ram_mem1_reg[5][15]/P0001 , \wishbone_bd_ram_mem1_reg[5][8]/P0001 , \wishbone_bd_ram_mem1_reg[5][9]/P0001 , \wishbone_bd_ram_mem1_reg[60][10]/P0001 , \wishbone_bd_ram_mem1_reg[60][11]/P0001 , \wishbone_bd_ram_mem1_reg[60][12]/P0001 , \wishbone_bd_ram_mem1_reg[60][13]/P0001 , \wishbone_bd_ram_mem1_reg[60][14]/P0001 , \wishbone_bd_ram_mem1_reg[60][15]/P0001 , \wishbone_bd_ram_mem1_reg[60][8]/P0001 , \wishbone_bd_ram_mem1_reg[60][9]/P0001 , \wishbone_bd_ram_mem1_reg[61][10]/P0001 , \wishbone_bd_ram_mem1_reg[61][11]/P0001 , \wishbone_bd_ram_mem1_reg[61][12]/P0001 , \wishbone_bd_ram_mem1_reg[61][13]/P0001 , \wishbone_bd_ram_mem1_reg[61][14]/P0001 , \wishbone_bd_ram_mem1_reg[61][15]/P0001 , \wishbone_bd_ram_mem1_reg[61][8]/P0001 , \wishbone_bd_ram_mem1_reg[61][9]/P0001 , \wishbone_bd_ram_mem1_reg[62][10]/P0001 , \wishbone_bd_ram_mem1_reg[62][11]/P0001 , \wishbone_bd_ram_mem1_reg[62][12]/P0001 , \wishbone_bd_ram_mem1_reg[62][13]/P0001 , \wishbone_bd_ram_mem1_reg[62][14]/P0001 , \wishbone_bd_ram_mem1_reg[62][15]/P0001 , \wishbone_bd_ram_mem1_reg[62][8]/P0001 , \wishbone_bd_ram_mem1_reg[62][9]/P0001 , \wishbone_bd_ram_mem1_reg[63][10]/P0001 , \wishbone_bd_ram_mem1_reg[63][11]/P0001 , \wishbone_bd_ram_mem1_reg[63][12]/P0001 , \wishbone_bd_ram_mem1_reg[63][13]/P0001 , \wishbone_bd_ram_mem1_reg[63][14]/P0001 , \wishbone_bd_ram_mem1_reg[63][15]/P0001 , \wishbone_bd_ram_mem1_reg[63][8]/P0001 , \wishbone_bd_ram_mem1_reg[63][9]/P0001 , \wishbone_bd_ram_mem1_reg[64][10]/P0001 , \wishbone_bd_ram_mem1_reg[64][11]/P0001 , \wishbone_bd_ram_mem1_reg[64][12]/P0001 , \wishbone_bd_ram_mem1_reg[64][13]/P0001 , \wishbone_bd_ram_mem1_reg[64][14]/P0001 , \wishbone_bd_ram_mem1_reg[64][15]/P0001 , \wishbone_bd_ram_mem1_reg[64][8]/P0001 , \wishbone_bd_ram_mem1_reg[64][9]/P0001 , \wishbone_bd_ram_mem1_reg[65][10]/P0001 , \wishbone_bd_ram_mem1_reg[65][11]/P0001 , \wishbone_bd_ram_mem1_reg[65][12]/P0001 , \wishbone_bd_ram_mem1_reg[65][13]/P0001 , \wishbone_bd_ram_mem1_reg[65][14]/P0001 , \wishbone_bd_ram_mem1_reg[65][15]/P0001 , \wishbone_bd_ram_mem1_reg[65][8]/P0001 , \wishbone_bd_ram_mem1_reg[65][9]/P0001 , \wishbone_bd_ram_mem1_reg[66][10]/P0001 , \wishbone_bd_ram_mem1_reg[66][11]/P0001 , \wishbone_bd_ram_mem1_reg[66][12]/P0001 , \wishbone_bd_ram_mem1_reg[66][13]/P0001 , \wishbone_bd_ram_mem1_reg[66][14]/P0001 , \wishbone_bd_ram_mem1_reg[66][15]/P0001 , \wishbone_bd_ram_mem1_reg[66][8]/P0001 , \wishbone_bd_ram_mem1_reg[66][9]/P0001 , \wishbone_bd_ram_mem1_reg[67][10]/P0001 , \wishbone_bd_ram_mem1_reg[67][11]/P0001 , \wishbone_bd_ram_mem1_reg[67][12]/P0001 , \wishbone_bd_ram_mem1_reg[67][13]/P0001 , \wishbone_bd_ram_mem1_reg[67][14]/P0001 , \wishbone_bd_ram_mem1_reg[67][15]/P0001 , \wishbone_bd_ram_mem1_reg[67][8]/P0001 , \wishbone_bd_ram_mem1_reg[67][9]/P0001 , \wishbone_bd_ram_mem1_reg[68][10]/P0001 , \wishbone_bd_ram_mem1_reg[68][11]/P0001 , \wishbone_bd_ram_mem1_reg[68][12]/P0001 , \wishbone_bd_ram_mem1_reg[68][13]/P0001 , \wishbone_bd_ram_mem1_reg[68][14]/P0001 , \wishbone_bd_ram_mem1_reg[68][15]/P0001 , \wishbone_bd_ram_mem1_reg[68][8]/P0001 , \wishbone_bd_ram_mem1_reg[68][9]/P0001 , \wishbone_bd_ram_mem1_reg[69][10]/P0001 , \wishbone_bd_ram_mem1_reg[69][11]/P0001 , \wishbone_bd_ram_mem1_reg[69][12]/P0001 , \wishbone_bd_ram_mem1_reg[69][13]/P0001 , \wishbone_bd_ram_mem1_reg[69][14]/P0001 , \wishbone_bd_ram_mem1_reg[69][15]/P0001 , \wishbone_bd_ram_mem1_reg[69][8]/P0001 , \wishbone_bd_ram_mem1_reg[69][9]/P0001 , \wishbone_bd_ram_mem1_reg[6][10]/P0001 , \wishbone_bd_ram_mem1_reg[6][11]/P0001 , \wishbone_bd_ram_mem1_reg[6][12]/P0001 , \wishbone_bd_ram_mem1_reg[6][13]/P0001 , \wishbone_bd_ram_mem1_reg[6][14]/P0001 , \wishbone_bd_ram_mem1_reg[6][15]/P0001 , \wishbone_bd_ram_mem1_reg[6][8]/P0001 , \wishbone_bd_ram_mem1_reg[6][9]/P0001 , \wishbone_bd_ram_mem1_reg[70][10]/P0001 , \wishbone_bd_ram_mem1_reg[70][11]/P0001 , \wishbone_bd_ram_mem1_reg[70][12]/P0001 , \wishbone_bd_ram_mem1_reg[70][13]/P0001 , \wishbone_bd_ram_mem1_reg[70][14]/P0001 , \wishbone_bd_ram_mem1_reg[70][15]/P0001 , \wishbone_bd_ram_mem1_reg[70][8]/P0001 , \wishbone_bd_ram_mem1_reg[70][9]/P0001 , \wishbone_bd_ram_mem1_reg[71][10]/P0001 , \wishbone_bd_ram_mem1_reg[71][11]/P0001 , \wishbone_bd_ram_mem1_reg[71][12]/P0001 , \wishbone_bd_ram_mem1_reg[71][13]/P0001 , \wishbone_bd_ram_mem1_reg[71][14]/P0001 , \wishbone_bd_ram_mem1_reg[71][15]/P0001 , \wishbone_bd_ram_mem1_reg[71][8]/P0001 , \wishbone_bd_ram_mem1_reg[71][9]/P0001 , \wishbone_bd_ram_mem1_reg[72][10]/P0001 , \wishbone_bd_ram_mem1_reg[72][11]/P0001 , \wishbone_bd_ram_mem1_reg[72][12]/P0001 , \wishbone_bd_ram_mem1_reg[72][13]/P0001 , \wishbone_bd_ram_mem1_reg[72][14]/P0001 , \wishbone_bd_ram_mem1_reg[72][15]/P0001 , \wishbone_bd_ram_mem1_reg[72][8]/P0001 , \wishbone_bd_ram_mem1_reg[72][9]/P0001 , \wishbone_bd_ram_mem1_reg[73][10]/P0001 , \wishbone_bd_ram_mem1_reg[73][11]/P0001 , \wishbone_bd_ram_mem1_reg[73][12]/P0001 , \wishbone_bd_ram_mem1_reg[73][13]/P0001 , \wishbone_bd_ram_mem1_reg[73][14]/P0001 , \wishbone_bd_ram_mem1_reg[73][15]/P0001 , \wishbone_bd_ram_mem1_reg[73][8]/P0001 , \wishbone_bd_ram_mem1_reg[73][9]/P0001 , \wishbone_bd_ram_mem1_reg[74][10]/P0001 , \wishbone_bd_ram_mem1_reg[74][11]/P0001 , \wishbone_bd_ram_mem1_reg[74][12]/P0001 , \wishbone_bd_ram_mem1_reg[74][13]/P0001 , \wishbone_bd_ram_mem1_reg[74][14]/P0001 , \wishbone_bd_ram_mem1_reg[74][15]/P0001 , \wishbone_bd_ram_mem1_reg[74][8]/P0001 , \wishbone_bd_ram_mem1_reg[74][9]/P0001 , \wishbone_bd_ram_mem1_reg[75][10]/P0001 , \wishbone_bd_ram_mem1_reg[75][11]/P0001 , \wishbone_bd_ram_mem1_reg[75][12]/P0001 , \wishbone_bd_ram_mem1_reg[75][13]/P0001 , \wishbone_bd_ram_mem1_reg[75][14]/P0001 , \wishbone_bd_ram_mem1_reg[75][15]/P0001 , \wishbone_bd_ram_mem1_reg[75][8]/P0001 , \wishbone_bd_ram_mem1_reg[75][9]/P0001 , \wishbone_bd_ram_mem1_reg[76][10]/P0001 , \wishbone_bd_ram_mem1_reg[76][11]/P0001 , \wishbone_bd_ram_mem1_reg[76][12]/P0001 , \wishbone_bd_ram_mem1_reg[76][13]/P0001 , \wishbone_bd_ram_mem1_reg[76][14]/P0001 , \wishbone_bd_ram_mem1_reg[76][15]/P0001 , \wishbone_bd_ram_mem1_reg[76][8]/P0001 , \wishbone_bd_ram_mem1_reg[76][9]/P0001 , \wishbone_bd_ram_mem1_reg[77][10]/P0001 , \wishbone_bd_ram_mem1_reg[77][11]/P0001 , \wishbone_bd_ram_mem1_reg[77][12]/P0001 , \wishbone_bd_ram_mem1_reg[77][13]/P0001 , \wishbone_bd_ram_mem1_reg[77][14]/P0001 , \wishbone_bd_ram_mem1_reg[77][15]/P0001 , \wishbone_bd_ram_mem1_reg[77][8]/P0001 , \wishbone_bd_ram_mem1_reg[77][9]/P0001 , \wishbone_bd_ram_mem1_reg[78][10]/P0001 , \wishbone_bd_ram_mem1_reg[78][11]/P0001 , \wishbone_bd_ram_mem1_reg[78][12]/P0001 , \wishbone_bd_ram_mem1_reg[78][13]/P0001 , \wishbone_bd_ram_mem1_reg[78][14]/P0001 , \wishbone_bd_ram_mem1_reg[78][15]/P0001 , \wishbone_bd_ram_mem1_reg[78][8]/P0001 , \wishbone_bd_ram_mem1_reg[78][9]/P0001 , \wishbone_bd_ram_mem1_reg[79][10]/P0001 , \wishbone_bd_ram_mem1_reg[79][11]/P0001 , \wishbone_bd_ram_mem1_reg[79][12]/P0001 , \wishbone_bd_ram_mem1_reg[79][13]/P0001 , \wishbone_bd_ram_mem1_reg[79][14]/P0001 , \wishbone_bd_ram_mem1_reg[79][15]/P0001 , \wishbone_bd_ram_mem1_reg[79][8]/P0001 , \wishbone_bd_ram_mem1_reg[79][9]/P0001 , \wishbone_bd_ram_mem1_reg[7][10]/P0001 , \wishbone_bd_ram_mem1_reg[7][11]/P0001 , \wishbone_bd_ram_mem1_reg[7][12]/P0001 , \wishbone_bd_ram_mem1_reg[7][13]/P0001 , \wishbone_bd_ram_mem1_reg[7][14]/P0001 , \wishbone_bd_ram_mem1_reg[7][15]/P0001 , \wishbone_bd_ram_mem1_reg[7][8]/P0001 , \wishbone_bd_ram_mem1_reg[7][9]/P0001 , \wishbone_bd_ram_mem1_reg[80][10]/P0001 , \wishbone_bd_ram_mem1_reg[80][11]/P0001 , \wishbone_bd_ram_mem1_reg[80][12]/P0001 , \wishbone_bd_ram_mem1_reg[80][13]/P0001 , \wishbone_bd_ram_mem1_reg[80][14]/P0001 , \wishbone_bd_ram_mem1_reg[80][15]/P0001 , \wishbone_bd_ram_mem1_reg[80][8]/P0001 , \wishbone_bd_ram_mem1_reg[80][9]/P0001 , \wishbone_bd_ram_mem1_reg[81][10]/P0001 , \wishbone_bd_ram_mem1_reg[81][11]/P0001 , \wishbone_bd_ram_mem1_reg[81][12]/P0001 , \wishbone_bd_ram_mem1_reg[81][13]/P0001 , \wishbone_bd_ram_mem1_reg[81][14]/P0001 , \wishbone_bd_ram_mem1_reg[81][15]/P0001 , \wishbone_bd_ram_mem1_reg[81][8]/P0001 , \wishbone_bd_ram_mem1_reg[81][9]/P0001 , \wishbone_bd_ram_mem1_reg[82][10]/P0001 , \wishbone_bd_ram_mem1_reg[82][11]/P0001 , \wishbone_bd_ram_mem1_reg[82][12]/P0001 , \wishbone_bd_ram_mem1_reg[82][13]/P0001 , \wishbone_bd_ram_mem1_reg[82][14]/P0001 , \wishbone_bd_ram_mem1_reg[82][15]/P0001 , \wishbone_bd_ram_mem1_reg[82][8]/P0001 , \wishbone_bd_ram_mem1_reg[82][9]/P0001 , \wishbone_bd_ram_mem1_reg[83][10]/P0001 , \wishbone_bd_ram_mem1_reg[83][11]/P0001 , \wishbone_bd_ram_mem1_reg[83][12]/P0001 , \wishbone_bd_ram_mem1_reg[83][13]/P0001 , \wishbone_bd_ram_mem1_reg[83][14]/P0001 , \wishbone_bd_ram_mem1_reg[83][15]/P0001 , \wishbone_bd_ram_mem1_reg[83][8]/P0001 , \wishbone_bd_ram_mem1_reg[83][9]/P0001 , \wishbone_bd_ram_mem1_reg[84][10]/P0001 , \wishbone_bd_ram_mem1_reg[84][11]/P0001 , \wishbone_bd_ram_mem1_reg[84][12]/P0001 , \wishbone_bd_ram_mem1_reg[84][13]/P0001 , \wishbone_bd_ram_mem1_reg[84][14]/P0001 , \wishbone_bd_ram_mem1_reg[84][15]/P0001 , \wishbone_bd_ram_mem1_reg[84][8]/P0001 , \wishbone_bd_ram_mem1_reg[84][9]/P0001 , \wishbone_bd_ram_mem1_reg[85][10]/P0001 , \wishbone_bd_ram_mem1_reg[85][11]/P0001 , \wishbone_bd_ram_mem1_reg[85][12]/P0001 , \wishbone_bd_ram_mem1_reg[85][13]/P0001 , \wishbone_bd_ram_mem1_reg[85][14]/P0001 , \wishbone_bd_ram_mem1_reg[85][15]/P0001 , \wishbone_bd_ram_mem1_reg[85][8]/P0001 , \wishbone_bd_ram_mem1_reg[85][9]/P0001 , \wishbone_bd_ram_mem1_reg[86][10]/P0001 , \wishbone_bd_ram_mem1_reg[86][11]/P0001 , \wishbone_bd_ram_mem1_reg[86][12]/P0001 , \wishbone_bd_ram_mem1_reg[86][13]/P0001 , \wishbone_bd_ram_mem1_reg[86][14]/P0001 , \wishbone_bd_ram_mem1_reg[86][15]/P0001 , \wishbone_bd_ram_mem1_reg[86][8]/P0001 , \wishbone_bd_ram_mem1_reg[86][9]/P0001 , \wishbone_bd_ram_mem1_reg[87][10]/P0001 , \wishbone_bd_ram_mem1_reg[87][11]/P0001 , \wishbone_bd_ram_mem1_reg[87][12]/P0001 , \wishbone_bd_ram_mem1_reg[87][13]/P0001 , \wishbone_bd_ram_mem1_reg[87][14]/P0001 , \wishbone_bd_ram_mem1_reg[87][15]/P0001 , \wishbone_bd_ram_mem1_reg[87][8]/P0001 , \wishbone_bd_ram_mem1_reg[87][9]/P0001 , \wishbone_bd_ram_mem1_reg[88][10]/P0001 , \wishbone_bd_ram_mem1_reg[88][11]/P0001 , \wishbone_bd_ram_mem1_reg[88][12]/P0001 , \wishbone_bd_ram_mem1_reg[88][13]/P0001 , \wishbone_bd_ram_mem1_reg[88][14]/P0001 , \wishbone_bd_ram_mem1_reg[88][15]/P0001 , \wishbone_bd_ram_mem1_reg[88][8]/P0001 , \wishbone_bd_ram_mem1_reg[88][9]/P0001 , \wishbone_bd_ram_mem1_reg[89][10]/P0001 , \wishbone_bd_ram_mem1_reg[89][11]/P0001 , \wishbone_bd_ram_mem1_reg[89][12]/P0001 , \wishbone_bd_ram_mem1_reg[89][13]/P0001 , \wishbone_bd_ram_mem1_reg[89][14]/P0001 , \wishbone_bd_ram_mem1_reg[89][15]/P0001 , \wishbone_bd_ram_mem1_reg[89][8]/P0001 , \wishbone_bd_ram_mem1_reg[89][9]/P0001 , \wishbone_bd_ram_mem1_reg[8][10]/P0001 , \wishbone_bd_ram_mem1_reg[8][11]/P0001 , \wishbone_bd_ram_mem1_reg[8][12]/P0001 , \wishbone_bd_ram_mem1_reg[8][13]/P0001 , \wishbone_bd_ram_mem1_reg[8][14]/P0001 , \wishbone_bd_ram_mem1_reg[8][15]/P0001 , \wishbone_bd_ram_mem1_reg[8][8]/P0001 , \wishbone_bd_ram_mem1_reg[8][9]/P0001 , \wishbone_bd_ram_mem1_reg[90][10]/P0001 , \wishbone_bd_ram_mem1_reg[90][11]/P0001 , \wishbone_bd_ram_mem1_reg[90][12]/P0001 , \wishbone_bd_ram_mem1_reg[90][13]/P0001 , \wishbone_bd_ram_mem1_reg[90][14]/P0001 , \wishbone_bd_ram_mem1_reg[90][15]/P0001 , \wishbone_bd_ram_mem1_reg[90][8]/P0001 , \wishbone_bd_ram_mem1_reg[90][9]/P0001 , \wishbone_bd_ram_mem1_reg[91][10]/P0001 , \wishbone_bd_ram_mem1_reg[91][11]/P0001 , \wishbone_bd_ram_mem1_reg[91][12]/P0001 , \wishbone_bd_ram_mem1_reg[91][13]/P0001 , \wishbone_bd_ram_mem1_reg[91][14]/P0001 , \wishbone_bd_ram_mem1_reg[91][15]/P0001 , \wishbone_bd_ram_mem1_reg[91][8]/P0001 , \wishbone_bd_ram_mem1_reg[91][9]/P0001 , \wishbone_bd_ram_mem1_reg[92][10]/P0001 , \wishbone_bd_ram_mem1_reg[92][11]/P0001 , \wishbone_bd_ram_mem1_reg[92][12]/P0001 , \wishbone_bd_ram_mem1_reg[92][13]/P0001 , \wishbone_bd_ram_mem1_reg[92][14]/P0001 , \wishbone_bd_ram_mem1_reg[92][15]/P0001 , \wishbone_bd_ram_mem1_reg[92][8]/P0001 , \wishbone_bd_ram_mem1_reg[92][9]/P0001 , \wishbone_bd_ram_mem1_reg[93][10]/P0001 , \wishbone_bd_ram_mem1_reg[93][11]/P0001 , \wishbone_bd_ram_mem1_reg[93][12]/P0001 , \wishbone_bd_ram_mem1_reg[93][13]/P0001 , \wishbone_bd_ram_mem1_reg[93][14]/P0001 , \wishbone_bd_ram_mem1_reg[93][15]/P0001 , \wishbone_bd_ram_mem1_reg[93][8]/P0001 , \wishbone_bd_ram_mem1_reg[93][9]/P0001 , \wishbone_bd_ram_mem1_reg[94][10]/P0001 , \wishbone_bd_ram_mem1_reg[94][11]/P0001 , \wishbone_bd_ram_mem1_reg[94][12]/P0001 , \wishbone_bd_ram_mem1_reg[94][13]/P0001 , \wishbone_bd_ram_mem1_reg[94][14]/P0001 , \wishbone_bd_ram_mem1_reg[94][15]/P0001 , \wishbone_bd_ram_mem1_reg[94][8]/P0001 , \wishbone_bd_ram_mem1_reg[94][9]/P0001 , \wishbone_bd_ram_mem1_reg[95][10]/P0001 , \wishbone_bd_ram_mem1_reg[95][11]/P0001 , \wishbone_bd_ram_mem1_reg[95][12]/P0001 , \wishbone_bd_ram_mem1_reg[95][13]/P0001 , \wishbone_bd_ram_mem1_reg[95][14]/P0001 , \wishbone_bd_ram_mem1_reg[95][15]/P0001 , \wishbone_bd_ram_mem1_reg[95][8]/P0001 , \wishbone_bd_ram_mem1_reg[95][9]/P0001 , \wishbone_bd_ram_mem1_reg[96][10]/P0001 , \wishbone_bd_ram_mem1_reg[96][11]/P0001 , \wishbone_bd_ram_mem1_reg[96][12]/P0001 , \wishbone_bd_ram_mem1_reg[96][13]/P0001 , \wishbone_bd_ram_mem1_reg[96][14]/P0001 , \wishbone_bd_ram_mem1_reg[96][15]/P0001 , \wishbone_bd_ram_mem1_reg[96][8]/P0001 , \wishbone_bd_ram_mem1_reg[96][9]/P0001 , \wishbone_bd_ram_mem1_reg[97][10]/P0001 , \wishbone_bd_ram_mem1_reg[97][11]/P0001 , \wishbone_bd_ram_mem1_reg[97][12]/P0001 , \wishbone_bd_ram_mem1_reg[97][13]/P0001 , \wishbone_bd_ram_mem1_reg[97][14]/P0001 , \wishbone_bd_ram_mem1_reg[97][15]/P0001 , \wishbone_bd_ram_mem1_reg[97][8]/P0001 , \wishbone_bd_ram_mem1_reg[97][9]/P0001 , \wishbone_bd_ram_mem1_reg[98][10]/P0001 , \wishbone_bd_ram_mem1_reg[98][11]/P0001 , \wishbone_bd_ram_mem1_reg[98][12]/P0001 , \wishbone_bd_ram_mem1_reg[98][13]/P0001 , \wishbone_bd_ram_mem1_reg[98][14]/P0001 , \wishbone_bd_ram_mem1_reg[98][15]/P0001 , \wishbone_bd_ram_mem1_reg[98][8]/P0001 , \wishbone_bd_ram_mem1_reg[98][9]/P0001 , \wishbone_bd_ram_mem1_reg[99][10]/P0001 , \wishbone_bd_ram_mem1_reg[99][11]/P0001 , \wishbone_bd_ram_mem1_reg[99][12]/P0001 , \wishbone_bd_ram_mem1_reg[99][13]/P0001 , \wishbone_bd_ram_mem1_reg[99][14]/P0001 , \wishbone_bd_ram_mem1_reg[99][15]/P0001 , \wishbone_bd_ram_mem1_reg[99][8]/P0001 , \wishbone_bd_ram_mem1_reg[99][9]/P0001 , \wishbone_bd_ram_mem1_reg[9][10]/P0001 , \wishbone_bd_ram_mem1_reg[9][11]/P0001 , \wishbone_bd_ram_mem1_reg[9][12]/P0001 , \wishbone_bd_ram_mem1_reg[9][13]/P0001 , \wishbone_bd_ram_mem1_reg[9][14]/P0001 , \wishbone_bd_ram_mem1_reg[9][15]/P0001 , \wishbone_bd_ram_mem1_reg[9][8]/P0001 , \wishbone_bd_ram_mem1_reg[9][9]/P0001 , \wishbone_bd_ram_mem2_reg[0][16]/P0001 , \wishbone_bd_ram_mem2_reg[0][17]/P0001 , \wishbone_bd_ram_mem2_reg[0][18]/P0001 , \wishbone_bd_ram_mem2_reg[0][19]/P0001 , \wishbone_bd_ram_mem2_reg[0][20]/P0001 , \wishbone_bd_ram_mem2_reg[0][21]/P0001 , \wishbone_bd_ram_mem2_reg[0][22]/P0001 , \wishbone_bd_ram_mem2_reg[0][23]/P0001 , \wishbone_bd_ram_mem2_reg[100][16]/P0001 , \wishbone_bd_ram_mem2_reg[100][17]/P0001 , \wishbone_bd_ram_mem2_reg[100][18]/P0001 , \wishbone_bd_ram_mem2_reg[100][19]/P0001 , \wishbone_bd_ram_mem2_reg[100][20]/P0001 , \wishbone_bd_ram_mem2_reg[100][21]/P0001 , \wishbone_bd_ram_mem2_reg[100][22]/P0001 , \wishbone_bd_ram_mem2_reg[100][23]/P0001 , \wishbone_bd_ram_mem2_reg[101][16]/P0001 , \wishbone_bd_ram_mem2_reg[101][17]/P0001 , \wishbone_bd_ram_mem2_reg[101][18]/P0001 , \wishbone_bd_ram_mem2_reg[101][19]/P0001 , \wishbone_bd_ram_mem2_reg[101][20]/P0001 , \wishbone_bd_ram_mem2_reg[101][21]/P0001 , \wishbone_bd_ram_mem2_reg[101][22]/P0001 , \wishbone_bd_ram_mem2_reg[101][23]/P0001 , \wishbone_bd_ram_mem2_reg[102][16]/P0001 , \wishbone_bd_ram_mem2_reg[102][17]/P0001 , \wishbone_bd_ram_mem2_reg[102][18]/P0001 , \wishbone_bd_ram_mem2_reg[102][19]/P0001 , \wishbone_bd_ram_mem2_reg[102][20]/P0001 , \wishbone_bd_ram_mem2_reg[102][21]/P0001 , \wishbone_bd_ram_mem2_reg[102][22]/P0001 , \wishbone_bd_ram_mem2_reg[102][23]/P0001 , \wishbone_bd_ram_mem2_reg[103][16]/P0001 , \wishbone_bd_ram_mem2_reg[103][17]/P0001 , \wishbone_bd_ram_mem2_reg[103][18]/P0001 , \wishbone_bd_ram_mem2_reg[103][19]/P0001 , \wishbone_bd_ram_mem2_reg[103][20]/P0001 , \wishbone_bd_ram_mem2_reg[103][21]/P0001 , \wishbone_bd_ram_mem2_reg[103][22]/P0001 , \wishbone_bd_ram_mem2_reg[103][23]/P0001 , \wishbone_bd_ram_mem2_reg[104][16]/P0001 , \wishbone_bd_ram_mem2_reg[104][17]/P0001 , \wishbone_bd_ram_mem2_reg[104][18]/P0001 , \wishbone_bd_ram_mem2_reg[104][19]/P0001 , \wishbone_bd_ram_mem2_reg[104][20]/P0001 , \wishbone_bd_ram_mem2_reg[104][21]/P0001 , \wishbone_bd_ram_mem2_reg[104][22]/P0001 , \wishbone_bd_ram_mem2_reg[104][23]/P0001 , \wishbone_bd_ram_mem2_reg[105][16]/P0001 , \wishbone_bd_ram_mem2_reg[105][17]/P0001 , \wishbone_bd_ram_mem2_reg[105][18]/P0001 , \wishbone_bd_ram_mem2_reg[105][19]/P0001 , \wishbone_bd_ram_mem2_reg[105][20]/P0001 , \wishbone_bd_ram_mem2_reg[105][21]/P0001 , \wishbone_bd_ram_mem2_reg[105][22]/P0001 , \wishbone_bd_ram_mem2_reg[105][23]/P0001 , \wishbone_bd_ram_mem2_reg[106][16]/P0001 , \wishbone_bd_ram_mem2_reg[106][17]/P0001 , \wishbone_bd_ram_mem2_reg[106][18]/P0001 , \wishbone_bd_ram_mem2_reg[106][19]/P0001 , \wishbone_bd_ram_mem2_reg[106][20]/P0001 , \wishbone_bd_ram_mem2_reg[106][21]/P0001 , \wishbone_bd_ram_mem2_reg[106][22]/P0001 , \wishbone_bd_ram_mem2_reg[106][23]/P0001 , \wishbone_bd_ram_mem2_reg[107][16]/P0001 , \wishbone_bd_ram_mem2_reg[107][17]/P0001 , \wishbone_bd_ram_mem2_reg[107][18]/P0001 , \wishbone_bd_ram_mem2_reg[107][19]/P0001 , \wishbone_bd_ram_mem2_reg[107][20]/P0001 , \wishbone_bd_ram_mem2_reg[107][21]/P0001 , \wishbone_bd_ram_mem2_reg[107][22]/P0001 , \wishbone_bd_ram_mem2_reg[107][23]/P0001 , \wishbone_bd_ram_mem2_reg[108][16]/P0001 , \wishbone_bd_ram_mem2_reg[108][17]/P0001 , \wishbone_bd_ram_mem2_reg[108][18]/P0001 , \wishbone_bd_ram_mem2_reg[108][19]/P0001 , \wishbone_bd_ram_mem2_reg[108][20]/P0001 , \wishbone_bd_ram_mem2_reg[108][21]/P0001 , \wishbone_bd_ram_mem2_reg[108][22]/P0001 , \wishbone_bd_ram_mem2_reg[108][23]/P0001 , \wishbone_bd_ram_mem2_reg[109][16]/P0001 , \wishbone_bd_ram_mem2_reg[109][17]/P0001 , \wishbone_bd_ram_mem2_reg[109][18]/P0001 , \wishbone_bd_ram_mem2_reg[109][19]/P0001 , \wishbone_bd_ram_mem2_reg[109][20]/P0001 , \wishbone_bd_ram_mem2_reg[109][21]/P0001 , \wishbone_bd_ram_mem2_reg[109][22]/P0001 , \wishbone_bd_ram_mem2_reg[109][23]/P0001 , \wishbone_bd_ram_mem2_reg[10][16]/P0001 , \wishbone_bd_ram_mem2_reg[10][17]/P0001 , \wishbone_bd_ram_mem2_reg[10][18]/P0001 , \wishbone_bd_ram_mem2_reg[10][19]/P0001 , \wishbone_bd_ram_mem2_reg[10][20]/P0001 , \wishbone_bd_ram_mem2_reg[10][21]/P0001 , \wishbone_bd_ram_mem2_reg[10][22]/P0001 , \wishbone_bd_ram_mem2_reg[10][23]/P0001 , \wishbone_bd_ram_mem2_reg[110][16]/P0001 , \wishbone_bd_ram_mem2_reg[110][17]/P0001 , \wishbone_bd_ram_mem2_reg[110][18]/P0001 , \wishbone_bd_ram_mem2_reg[110][19]/P0001 , \wishbone_bd_ram_mem2_reg[110][20]/P0001 , \wishbone_bd_ram_mem2_reg[110][21]/P0001 , \wishbone_bd_ram_mem2_reg[110][22]/P0001 , \wishbone_bd_ram_mem2_reg[110][23]/P0001 , \wishbone_bd_ram_mem2_reg[111][16]/P0001 , \wishbone_bd_ram_mem2_reg[111][17]/P0001 , \wishbone_bd_ram_mem2_reg[111][18]/P0001 , \wishbone_bd_ram_mem2_reg[111][19]/P0001 , \wishbone_bd_ram_mem2_reg[111][20]/P0001 , \wishbone_bd_ram_mem2_reg[111][21]/P0001 , \wishbone_bd_ram_mem2_reg[111][22]/P0001 , \wishbone_bd_ram_mem2_reg[111][23]/P0001 , \wishbone_bd_ram_mem2_reg[112][16]/P0001 , \wishbone_bd_ram_mem2_reg[112][17]/P0001 , \wishbone_bd_ram_mem2_reg[112][18]/P0001 , \wishbone_bd_ram_mem2_reg[112][19]/P0001 , \wishbone_bd_ram_mem2_reg[112][20]/P0001 , \wishbone_bd_ram_mem2_reg[112][21]/P0001 , \wishbone_bd_ram_mem2_reg[112][22]/P0001 , \wishbone_bd_ram_mem2_reg[112][23]/P0001 , \wishbone_bd_ram_mem2_reg[113][16]/P0001 , \wishbone_bd_ram_mem2_reg[113][17]/P0001 , \wishbone_bd_ram_mem2_reg[113][18]/P0001 , \wishbone_bd_ram_mem2_reg[113][19]/P0001 , \wishbone_bd_ram_mem2_reg[113][20]/P0001 , \wishbone_bd_ram_mem2_reg[113][21]/P0001 , \wishbone_bd_ram_mem2_reg[113][22]/P0001 , \wishbone_bd_ram_mem2_reg[113][23]/P0001 , \wishbone_bd_ram_mem2_reg[114][16]/P0001 , \wishbone_bd_ram_mem2_reg[114][17]/P0001 , \wishbone_bd_ram_mem2_reg[114][18]/P0001 , \wishbone_bd_ram_mem2_reg[114][19]/P0001 , \wishbone_bd_ram_mem2_reg[114][20]/P0001 , \wishbone_bd_ram_mem2_reg[114][21]/P0001 , \wishbone_bd_ram_mem2_reg[114][22]/P0001 , \wishbone_bd_ram_mem2_reg[114][23]/P0001 , \wishbone_bd_ram_mem2_reg[115][16]/P0001 , \wishbone_bd_ram_mem2_reg[115][17]/P0001 , \wishbone_bd_ram_mem2_reg[115][18]/P0001 , \wishbone_bd_ram_mem2_reg[115][19]/P0001 , \wishbone_bd_ram_mem2_reg[115][20]/P0001 , \wishbone_bd_ram_mem2_reg[115][21]/P0001 , \wishbone_bd_ram_mem2_reg[115][22]/P0001 , \wishbone_bd_ram_mem2_reg[115][23]/P0001 , \wishbone_bd_ram_mem2_reg[116][16]/P0001 , \wishbone_bd_ram_mem2_reg[116][17]/P0001 , \wishbone_bd_ram_mem2_reg[116][18]/P0001 , \wishbone_bd_ram_mem2_reg[116][19]/P0001 , \wishbone_bd_ram_mem2_reg[116][20]/P0001 , \wishbone_bd_ram_mem2_reg[116][21]/P0001 , \wishbone_bd_ram_mem2_reg[116][22]/P0001 , \wishbone_bd_ram_mem2_reg[116][23]/P0001 , \wishbone_bd_ram_mem2_reg[117][16]/P0001 , \wishbone_bd_ram_mem2_reg[117][17]/P0001 , \wishbone_bd_ram_mem2_reg[117][18]/P0001 , \wishbone_bd_ram_mem2_reg[117][19]/P0001 , \wishbone_bd_ram_mem2_reg[117][20]/P0001 , \wishbone_bd_ram_mem2_reg[117][21]/P0001 , \wishbone_bd_ram_mem2_reg[117][22]/P0001 , \wishbone_bd_ram_mem2_reg[117][23]/P0001 , \wishbone_bd_ram_mem2_reg[118][16]/P0001 , \wishbone_bd_ram_mem2_reg[118][17]/P0001 , \wishbone_bd_ram_mem2_reg[118][18]/P0001 , \wishbone_bd_ram_mem2_reg[118][19]/P0001 , \wishbone_bd_ram_mem2_reg[118][20]/P0001 , \wishbone_bd_ram_mem2_reg[118][21]/P0001 , \wishbone_bd_ram_mem2_reg[118][22]/P0001 , \wishbone_bd_ram_mem2_reg[118][23]/P0001 , \wishbone_bd_ram_mem2_reg[119][16]/P0001 , \wishbone_bd_ram_mem2_reg[119][17]/P0001 , \wishbone_bd_ram_mem2_reg[119][18]/P0001 , \wishbone_bd_ram_mem2_reg[119][19]/P0001 , \wishbone_bd_ram_mem2_reg[119][20]/P0001 , \wishbone_bd_ram_mem2_reg[119][21]/P0001 , \wishbone_bd_ram_mem2_reg[119][22]/P0001 , \wishbone_bd_ram_mem2_reg[119][23]/P0001 , \wishbone_bd_ram_mem2_reg[11][16]/P0001 , \wishbone_bd_ram_mem2_reg[11][17]/P0001 , \wishbone_bd_ram_mem2_reg[11][18]/P0001 , \wishbone_bd_ram_mem2_reg[11][19]/P0001 , \wishbone_bd_ram_mem2_reg[11][20]/P0001 , \wishbone_bd_ram_mem2_reg[11][21]/P0001 , \wishbone_bd_ram_mem2_reg[11][22]/P0001 , \wishbone_bd_ram_mem2_reg[11][23]/P0001 , \wishbone_bd_ram_mem2_reg[120][16]/P0001 , \wishbone_bd_ram_mem2_reg[120][17]/P0001 , \wishbone_bd_ram_mem2_reg[120][18]/P0001 , \wishbone_bd_ram_mem2_reg[120][19]/P0001 , \wishbone_bd_ram_mem2_reg[120][20]/P0001 , \wishbone_bd_ram_mem2_reg[120][21]/P0001 , \wishbone_bd_ram_mem2_reg[120][22]/P0001 , \wishbone_bd_ram_mem2_reg[120][23]/P0001 , \wishbone_bd_ram_mem2_reg[121][16]/P0001 , \wishbone_bd_ram_mem2_reg[121][17]/P0001 , \wishbone_bd_ram_mem2_reg[121][18]/P0001 , \wishbone_bd_ram_mem2_reg[121][19]/P0001 , \wishbone_bd_ram_mem2_reg[121][20]/P0001 , \wishbone_bd_ram_mem2_reg[121][21]/P0001 , \wishbone_bd_ram_mem2_reg[121][22]/P0001 , \wishbone_bd_ram_mem2_reg[121][23]/P0001 , \wishbone_bd_ram_mem2_reg[122][16]/P0001 , \wishbone_bd_ram_mem2_reg[122][17]/P0001 , \wishbone_bd_ram_mem2_reg[122][18]/P0001 , \wishbone_bd_ram_mem2_reg[122][19]/P0001 , \wishbone_bd_ram_mem2_reg[122][20]/P0001 , \wishbone_bd_ram_mem2_reg[122][21]/P0001 , \wishbone_bd_ram_mem2_reg[122][22]/P0001 , \wishbone_bd_ram_mem2_reg[122][23]/P0001 , \wishbone_bd_ram_mem2_reg[123][16]/P0001 , \wishbone_bd_ram_mem2_reg[123][17]/P0001 , \wishbone_bd_ram_mem2_reg[123][18]/P0001 , \wishbone_bd_ram_mem2_reg[123][19]/P0001 , \wishbone_bd_ram_mem2_reg[123][20]/P0001 , \wishbone_bd_ram_mem2_reg[123][21]/P0001 , \wishbone_bd_ram_mem2_reg[123][22]/P0001 , \wishbone_bd_ram_mem2_reg[123][23]/P0001 , \wishbone_bd_ram_mem2_reg[124][16]/P0001 , \wishbone_bd_ram_mem2_reg[124][17]/P0001 , \wishbone_bd_ram_mem2_reg[124][18]/P0001 , \wishbone_bd_ram_mem2_reg[124][19]/P0001 , \wishbone_bd_ram_mem2_reg[124][20]/P0001 , \wishbone_bd_ram_mem2_reg[124][21]/P0001 , \wishbone_bd_ram_mem2_reg[124][22]/P0001 , \wishbone_bd_ram_mem2_reg[124][23]/P0001 , \wishbone_bd_ram_mem2_reg[125][16]/P0001 , \wishbone_bd_ram_mem2_reg[125][17]/P0001 , \wishbone_bd_ram_mem2_reg[125][18]/P0001 , \wishbone_bd_ram_mem2_reg[125][19]/P0001 , \wishbone_bd_ram_mem2_reg[125][20]/P0001 , \wishbone_bd_ram_mem2_reg[125][21]/P0001 , \wishbone_bd_ram_mem2_reg[125][22]/P0001 , \wishbone_bd_ram_mem2_reg[125][23]/P0001 , \wishbone_bd_ram_mem2_reg[126][16]/P0001 , \wishbone_bd_ram_mem2_reg[126][17]/P0001 , \wishbone_bd_ram_mem2_reg[126][18]/P0001 , \wishbone_bd_ram_mem2_reg[126][19]/P0001 , \wishbone_bd_ram_mem2_reg[126][20]/P0001 , \wishbone_bd_ram_mem2_reg[126][21]/P0001 , \wishbone_bd_ram_mem2_reg[126][22]/P0001 , \wishbone_bd_ram_mem2_reg[126][23]/P0001 , \wishbone_bd_ram_mem2_reg[127][16]/P0001 , \wishbone_bd_ram_mem2_reg[127][17]/P0001 , \wishbone_bd_ram_mem2_reg[127][18]/P0001 , \wishbone_bd_ram_mem2_reg[127][19]/P0001 , \wishbone_bd_ram_mem2_reg[127][20]/P0001 , \wishbone_bd_ram_mem2_reg[127][21]/P0001 , \wishbone_bd_ram_mem2_reg[127][22]/P0001 , \wishbone_bd_ram_mem2_reg[127][23]/P0001 , \wishbone_bd_ram_mem2_reg[128][16]/P0001 , \wishbone_bd_ram_mem2_reg[128][17]/P0001 , \wishbone_bd_ram_mem2_reg[128][18]/P0001 , \wishbone_bd_ram_mem2_reg[128][19]/P0001 , \wishbone_bd_ram_mem2_reg[128][20]/P0001 , \wishbone_bd_ram_mem2_reg[128][21]/P0001 , \wishbone_bd_ram_mem2_reg[128][22]/P0001 , \wishbone_bd_ram_mem2_reg[128][23]/P0001 , \wishbone_bd_ram_mem2_reg[129][16]/P0001 , \wishbone_bd_ram_mem2_reg[129][17]/P0001 , \wishbone_bd_ram_mem2_reg[129][18]/P0001 , \wishbone_bd_ram_mem2_reg[129][19]/P0001 , \wishbone_bd_ram_mem2_reg[129][20]/P0001 , \wishbone_bd_ram_mem2_reg[129][21]/P0001 , \wishbone_bd_ram_mem2_reg[129][22]/P0001 , \wishbone_bd_ram_mem2_reg[129][23]/P0001 , \wishbone_bd_ram_mem2_reg[12][16]/P0001 , \wishbone_bd_ram_mem2_reg[12][17]/P0001 , \wishbone_bd_ram_mem2_reg[12][18]/P0001 , \wishbone_bd_ram_mem2_reg[12][19]/P0001 , \wishbone_bd_ram_mem2_reg[12][20]/P0001 , \wishbone_bd_ram_mem2_reg[12][21]/P0001 , \wishbone_bd_ram_mem2_reg[12][22]/P0001 , \wishbone_bd_ram_mem2_reg[12][23]/P0001 , \wishbone_bd_ram_mem2_reg[130][16]/P0001 , \wishbone_bd_ram_mem2_reg[130][17]/P0001 , \wishbone_bd_ram_mem2_reg[130][18]/P0001 , \wishbone_bd_ram_mem2_reg[130][19]/P0001 , \wishbone_bd_ram_mem2_reg[130][20]/P0001 , \wishbone_bd_ram_mem2_reg[130][21]/P0001 , \wishbone_bd_ram_mem2_reg[130][22]/P0001 , \wishbone_bd_ram_mem2_reg[130][23]/P0001 , \wishbone_bd_ram_mem2_reg[131][16]/P0001 , \wishbone_bd_ram_mem2_reg[131][17]/P0001 , \wishbone_bd_ram_mem2_reg[131][18]/P0001 , \wishbone_bd_ram_mem2_reg[131][19]/P0001 , \wishbone_bd_ram_mem2_reg[131][20]/P0001 , \wishbone_bd_ram_mem2_reg[131][21]/P0001 , \wishbone_bd_ram_mem2_reg[131][22]/P0001 , \wishbone_bd_ram_mem2_reg[131][23]/P0001 , \wishbone_bd_ram_mem2_reg[132][16]/P0001 , \wishbone_bd_ram_mem2_reg[132][17]/P0001 , \wishbone_bd_ram_mem2_reg[132][18]/P0001 , \wishbone_bd_ram_mem2_reg[132][19]/P0001 , \wishbone_bd_ram_mem2_reg[132][20]/P0001 , \wishbone_bd_ram_mem2_reg[132][21]/P0001 , \wishbone_bd_ram_mem2_reg[132][22]/P0001 , \wishbone_bd_ram_mem2_reg[132][23]/P0001 , \wishbone_bd_ram_mem2_reg[133][16]/P0001 , \wishbone_bd_ram_mem2_reg[133][17]/P0001 , \wishbone_bd_ram_mem2_reg[133][18]/P0001 , \wishbone_bd_ram_mem2_reg[133][19]/P0001 , \wishbone_bd_ram_mem2_reg[133][20]/P0001 , \wishbone_bd_ram_mem2_reg[133][21]/P0001 , \wishbone_bd_ram_mem2_reg[133][22]/P0001 , \wishbone_bd_ram_mem2_reg[133][23]/P0001 , \wishbone_bd_ram_mem2_reg[134][16]/P0001 , \wishbone_bd_ram_mem2_reg[134][17]/P0001 , \wishbone_bd_ram_mem2_reg[134][18]/P0001 , \wishbone_bd_ram_mem2_reg[134][19]/P0001 , \wishbone_bd_ram_mem2_reg[134][20]/P0001 , \wishbone_bd_ram_mem2_reg[134][21]/P0001 , \wishbone_bd_ram_mem2_reg[134][22]/P0001 , \wishbone_bd_ram_mem2_reg[134][23]/P0001 , \wishbone_bd_ram_mem2_reg[135][16]/P0001 , \wishbone_bd_ram_mem2_reg[135][17]/P0001 , \wishbone_bd_ram_mem2_reg[135][18]/P0001 , \wishbone_bd_ram_mem2_reg[135][19]/P0001 , \wishbone_bd_ram_mem2_reg[135][20]/P0001 , \wishbone_bd_ram_mem2_reg[135][21]/P0001 , \wishbone_bd_ram_mem2_reg[135][22]/P0001 , \wishbone_bd_ram_mem2_reg[135][23]/P0001 , \wishbone_bd_ram_mem2_reg[136][16]/P0001 , \wishbone_bd_ram_mem2_reg[136][17]/P0001 , \wishbone_bd_ram_mem2_reg[136][18]/P0001 , \wishbone_bd_ram_mem2_reg[136][19]/P0001 , \wishbone_bd_ram_mem2_reg[136][20]/P0001 , \wishbone_bd_ram_mem2_reg[136][21]/P0001 , \wishbone_bd_ram_mem2_reg[136][22]/P0001 , \wishbone_bd_ram_mem2_reg[136][23]/P0001 , \wishbone_bd_ram_mem2_reg[137][16]/P0001 , \wishbone_bd_ram_mem2_reg[137][17]/P0001 , \wishbone_bd_ram_mem2_reg[137][18]/P0001 , \wishbone_bd_ram_mem2_reg[137][19]/P0001 , \wishbone_bd_ram_mem2_reg[137][20]/P0001 , \wishbone_bd_ram_mem2_reg[137][21]/P0001 , \wishbone_bd_ram_mem2_reg[137][22]/P0001 , \wishbone_bd_ram_mem2_reg[137][23]/P0001 , \wishbone_bd_ram_mem2_reg[138][16]/P0001 , \wishbone_bd_ram_mem2_reg[138][17]/P0001 , \wishbone_bd_ram_mem2_reg[138][18]/P0001 , \wishbone_bd_ram_mem2_reg[138][19]/P0001 , \wishbone_bd_ram_mem2_reg[138][20]/P0001 , \wishbone_bd_ram_mem2_reg[138][21]/P0001 , \wishbone_bd_ram_mem2_reg[138][22]/P0001 , \wishbone_bd_ram_mem2_reg[138][23]/P0001 , \wishbone_bd_ram_mem2_reg[139][16]/P0001 , \wishbone_bd_ram_mem2_reg[139][17]/P0001 , \wishbone_bd_ram_mem2_reg[139][18]/P0001 , \wishbone_bd_ram_mem2_reg[139][19]/P0001 , \wishbone_bd_ram_mem2_reg[139][20]/P0001 , \wishbone_bd_ram_mem2_reg[139][21]/P0001 , \wishbone_bd_ram_mem2_reg[139][22]/P0001 , \wishbone_bd_ram_mem2_reg[139][23]/P0001 , \wishbone_bd_ram_mem2_reg[13][16]/P0001 , \wishbone_bd_ram_mem2_reg[13][17]/P0001 , \wishbone_bd_ram_mem2_reg[13][18]/P0001 , \wishbone_bd_ram_mem2_reg[13][19]/P0001 , \wishbone_bd_ram_mem2_reg[13][20]/P0001 , \wishbone_bd_ram_mem2_reg[13][21]/P0001 , \wishbone_bd_ram_mem2_reg[13][22]/P0001 , \wishbone_bd_ram_mem2_reg[13][23]/P0001 , \wishbone_bd_ram_mem2_reg[140][16]/P0001 , \wishbone_bd_ram_mem2_reg[140][17]/P0001 , \wishbone_bd_ram_mem2_reg[140][18]/P0001 , \wishbone_bd_ram_mem2_reg[140][19]/P0001 , \wishbone_bd_ram_mem2_reg[140][20]/P0001 , \wishbone_bd_ram_mem2_reg[140][21]/P0001 , \wishbone_bd_ram_mem2_reg[140][22]/P0001 , \wishbone_bd_ram_mem2_reg[140][23]/P0001 , \wishbone_bd_ram_mem2_reg[141][16]/P0001 , \wishbone_bd_ram_mem2_reg[141][17]/P0001 , \wishbone_bd_ram_mem2_reg[141][18]/P0001 , \wishbone_bd_ram_mem2_reg[141][19]/P0001 , \wishbone_bd_ram_mem2_reg[141][20]/P0001 , \wishbone_bd_ram_mem2_reg[141][21]/P0001 , \wishbone_bd_ram_mem2_reg[141][22]/P0001 , \wishbone_bd_ram_mem2_reg[141][23]/P0001 , \wishbone_bd_ram_mem2_reg[142][16]/P0001 , \wishbone_bd_ram_mem2_reg[142][17]/P0001 , \wishbone_bd_ram_mem2_reg[142][18]/P0001 , \wishbone_bd_ram_mem2_reg[142][19]/P0001 , \wishbone_bd_ram_mem2_reg[142][20]/P0001 , \wishbone_bd_ram_mem2_reg[142][21]/P0001 , \wishbone_bd_ram_mem2_reg[142][22]/P0001 , \wishbone_bd_ram_mem2_reg[142][23]/P0001 , \wishbone_bd_ram_mem2_reg[143][16]/P0001 , \wishbone_bd_ram_mem2_reg[143][17]/P0001 , \wishbone_bd_ram_mem2_reg[143][18]/P0001 , \wishbone_bd_ram_mem2_reg[143][19]/P0001 , \wishbone_bd_ram_mem2_reg[143][20]/P0001 , \wishbone_bd_ram_mem2_reg[143][21]/P0001 , \wishbone_bd_ram_mem2_reg[143][22]/P0001 , \wishbone_bd_ram_mem2_reg[143][23]/P0001 , \wishbone_bd_ram_mem2_reg[144][16]/P0001 , \wishbone_bd_ram_mem2_reg[144][17]/P0001 , \wishbone_bd_ram_mem2_reg[144][18]/P0001 , \wishbone_bd_ram_mem2_reg[144][19]/P0001 , \wishbone_bd_ram_mem2_reg[144][20]/P0001 , \wishbone_bd_ram_mem2_reg[144][21]/P0001 , \wishbone_bd_ram_mem2_reg[144][22]/P0001 , \wishbone_bd_ram_mem2_reg[144][23]/P0001 , \wishbone_bd_ram_mem2_reg[145][16]/P0001 , \wishbone_bd_ram_mem2_reg[145][17]/P0001 , \wishbone_bd_ram_mem2_reg[145][18]/P0001 , \wishbone_bd_ram_mem2_reg[145][19]/P0001 , \wishbone_bd_ram_mem2_reg[145][20]/P0001 , \wishbone_bd_ram_mem2_reg[145][21]/P0001 , \wishbone_bd_ram_mem2_reg[145][22]/P0001 , \wishbone_bd_ram_mem2_reg[145][23]/P0001 , \wishbone_bd_ram_mem2_reg[146][16]/P0001 , \wishbone_bd_ram_mem2_reg[146][17]/P0001 , \wishbone_bd_ram_mem2_reg[146][18]/P0001 , \wishbone_bd_ram_mem2_reg[146][19]/P0001 , \wishbone_bd_ram_mem2_reg[146][20]/P0001 , \wishbone_bd_ram_mem2_reg[146][21]/P0001 , \wishbone_bd_ram_mem2_reg[146][22]/P0001 , \wishbone_bd_ram_mem2_reg[146][23]/P0001 , \wishbone_bd_ram_mem2_reg[147][16]/P0001 , \wishbone_bd_ram_mem2_reg[147][17]/P0001 , \wishbone_bd_ram_mem2_reg[147][18]/P0001 , \wishbone_bd_ram_mem2_reg[147][19]/P0001 , \wishbone_bd_ram_mem2_reg[147][20]/P0001 , \wishbone_bd_ram_mem2_reg[147][21]/P0001 , \wishbone_bd_ram_mem2_reg[147][22]/P0001 , \wishbone_bd_ram_mem2_reg[147][23]/P0001 , \wishbone_bd_ram_mem2_reg[148][16]/P0001 , \wishbone_bd_ram_mem2_reg[148][17]/P0001 , \wishbone_bd_ram_mem2_reg[148][18]/P0001 , \wishbone_bd_ram_mem2_reg[148][19]/P0001 , \wishbone_bd_ram_mem2_reg[148][20]/P0001 , \wishbone_bd_ram_mem2_reg[148][21]/P0001 , \wishbone_bd_ram_mem2_reg[148][22]/P0001 , \wishbone_bd_ram_mem2_reg[148][23]/P0001 , \wishbone_bd_ram_mem2_reg[149][16]/P0001 , \wishbone_bd_ram_mem2_reg[149][17]/P0001 , \wishbone_bd_ram_mem2_reg[149][18]/P0001 , \wishbone_bd_ram_mem2_reg[149][19]/P0001 , \wishbone_bd_ram_mem2_reg[149][20]/P0001 , \wishbone_bd_ram_mem2_reg[149][21]/P0001 , \wishbone_bd_ram_mem2_reg[149][22]/P0001 , \wishbone_bd_ram_mem2_reg[149][23]/P0001 , \wishbone_bd_ram_mem2_reg[14][16]/P0001 , \wishbone_bd_ram_mem2_reg[14][17]/P0001 , \wishbone_bd_ram_mem2_reg[14][18]/P0001 , \wishbone_bd_ram_mem2_reg[14][19]/P0001 , \wishbone_bd_ram_mem2_reg[14][20]/P0001 , \wishbone_bd_ram_mem2_reg[14][21]/P0001 , \wishbone_bd_ram_mem2_reg[14][22]/P0001 , \wishbone_bd_ram_mem2_reg[14][23]/P0001 , \wishbone_bd_ram_mem2_reg[150][16]/P0001 , \wishbone_bd_ram_mem2_reg[150][17]/P0001 , \wishbone_bd_ram_mem2_reg[150][18]/P0001 , \wishbone_bd_ram_mem2_reg[150][19]/P0001 , \wishbone_bd_ram_mem2_reg[150][20]/P0001 , \wishbone_bd_ram_mem2_reg[150][21]/P0001 , \wishbone_bd_ram_mem2_reg[150][22]/P0001 , \wishbone_bd_ram_mem2_reg[150][23]/P0001 , \wishbone_bd_ram_mem2_reg[151][16]/P0001 , \wishbone_bd_ram_mem2_reg[151][17]/P0001 , \wishbone_bd_ram_mem2_reg[151][18]/P0001 , \wishbone_bd_ram_mem2_reg[151][19]/P0001 , \wishbone_bd_ram_mem2_reg[151][20]/P0001 , \wishbone_bd_ram_mem2_reg[151][21]/P0001 , \wishbone_bd_ram_mem2_reg[151][22]/P0001 , \wishbone_bd_ram_mem2_reg[151][23]/P0001 , \wishbone_bd_ram_mem2_reg[152][16]/P0001 , \wishbone_bd_ram_mem2_reg[152][17]/P0001 , \wishbone_bd_ram_mem2_reg[152][18]/P0001 , \wishbone_bd_ram_mem2_reg[152][19]/P0001 , \wishbone_bd_ram_mem2_reg[152][20]/P0001 , \wishbone_bd_ram_mem2_reg[152][21]/P0001 , \wishbone_bd_ram_mem2_reg[152][22]/P0001 , \wishbone_bd_ram_mem2_reg[152][23]/P0001 , \wishbone_bd_ram_mem2_reg[153][16]/P0001 , \wishbone_bd_ram_mem2_reg[153][17]/P0001 , \wishbone_bd_ram_mem2_reg[153][18]/P0001 , \wishbone_bd_ram_mem2_reg[153][19]/P0001 , \wishbone_bd_ram_mem2_reg[153][20]/P0001 , \wishbone_bd_ram_mem2_reg[153][21]/P0001 , \wishbone_bd_ram_mem2_reg[153][22]/P0001 , \wishbone_bd_ram_mem2_reg[153][23]/P0001 , \wishbone_bd_ram_mem2_reg[154][16]/P0001 , \wishbone_bd_ram_mem2_reg[154][17]/P0001 , \wishbone_bd_ram_mem2_reg[154][18]/P0001 , \wishbone_bd_ram_mem2_reg[154][19]/P0001 , \wishbone_bd_ram_mem2_reg[154][20]/P0001 , \wishbone_bd_ram_mem2_reg[154][21]/P0001 , \wishbone_bd_ram_mem2_reg[154][22]/P0001 , \wishbone_bd_ram_mem2_reg[154][23]/P0001 , \wishbone_bd_ram_mem2_reg[155][16]/P0001 , \wishbone_bd_ram_mem2_reg[155][17]/P0001 , \wishbone_bd_ram_mem2_reg[155][18]/P0001 , \wishbone_bd_ram_mem2_reg[155][19]/P0001 , \wishbone_bd_ram_mem2_reg[155][20]/P0001 , \wishbone_bd_ram_mem2_reg[155][21]/P0001 , \wishbone_bd_ram_mem2_reg[155][22]/P0001 , \wishbone_bd_ram_mem2_reg[155][23]/P0001 , \wishbone_bd_ram_mem2_reg[156][16]/P0001 , \wishbone_bd_ram_mem2_reg[156][17]/P0001 , \wishbone_bd_ram_mem2_reg[156][18]/P0001 , \wishbone_bd_ram_mem2_reg[156][19]/P0001 , \wishbone_bd_ram_mem2_reg[156][20]/P0001 , \wishbone_bd_ram_mem2_reg[156][21]/P0001 , \wishbone_bd_ram_mem2_reg[156][22]/P0001 , \wishbone_bd_ram_mem2_reg[156][23]/P0001 , \wishbone_bd_ram_mem2_reg[157][16]/P0001 , \wishbone_bd_ram_mem2_reg[157][17]/P0001 , \wishbone_bd_ram_mem2_reg[157][18]/P0001 , \wishbone_bd_ram_mem2_reg[157][19]/P0001 , \wishbone_bd_ram_mem2_reg[157][20]/P0001 , \wishbone_bd_ram_mem2_reg[157][21]/P0001 , \wishbone_bd_ram_mem2_reg[157][22]/P0001 , \wishbone_bd_ram_mem2_reg[157][23]/P0001 , \wishbone_bd_ram_mem2_reg[158][16]/P0001 , \wishbone_bd_ram_mem2_reg[158][17]/P0001 , \wishbone_bd_ram_mem2_reg[158][18]/P0001 , \wishbone_bd_ram_mem2_reg[158][19]/P0001 , \wishbone_bd_ram_mem2_reg[158][20]/P0001 , \wishbone_bd_ram_mem2_reg[158][21]/P0001 , \wishbone_bd_ram_mem2_reg[158][22]/P0001 , \wishbone_bd_ram_mem2_reg[158][23]/P0001 , \wishbone_bd_ram_mem2_reg[159][16]/P0001 , \wishbone_bd_ram_mem2_reg[159][17]/P0001 , \wishbone_bd_ram_mem2_reg[159][18]/P0001 , \wishbone_bd_ram_mem2_reg[159][19]/P0001 , \wishbone_bd_ram_mem2_reg[159][20]/P0001 , \wishbone_bd_ram_mem2_reg[159][21]/P0001 , \wishbone_bd_ram_mem2_reg[159][22]/P0001 , \wishbone_bd_ram_mem2_reg[159][23]/P0001 , \wishbone_bd_ram_mem2_reg[15][16]/P0001 , \wishbone_bd_ram_mem2_reg[15][17]/P0001 , \wishbone_bd_ram_mem2_reg[15][18]/P0001 , \wishbone_bd_ram_mem2_reg[15][19]/P0001 , \wishbone_bd_ram_mem2_reg[15][20]/P0001 , \wishbone_bd_ram_mem2_reg[15][21]/P0001 , \wishbone_bd_ram_mem2_reg[15][22]/P0001 , \wishbone_bd_ram_mem2_reg[15][23]/P0001 , \wishbone_bd_ram_mem2_reg[160][16]/P0001 , \wishbone_bd_ram_mem2_reg[160][17]/P0001 , \wishbone_bd_ram_mem2_reg[160][18]/P0001 , \wishbone_bd_ram_mem2_reg[160][19]/P0001 , \wishbone_bd_ram_mem2_reg[160][20]/P0001 , \wishbone_bd_ram_mem2_reg[160][21]/P0001 , \wishbone_bd_ram_mem2_reg[160][22]/P0001 , \wishbone_bd_ram_mem2_reg[160][23]/P0001 , \wishbone_bd_ram_mem2_reg[161][16]/P0001 , \wishbone_bd_ram_mem2_reg[161][17]/P0001 , \wishbone_bd_ram_mem2_reg[161][18]/P0001 , \wishbone_bd_ram_mem2_reg[161][19]/P0001 , \wishbone_bd_ram_mem2_reg[161][20]/P0001 , \wishbone_bd_ram_mem2_reg[161][21]/P0001 , \wishbone_bd_ram_mem2_reg[161][22]/P0001 , \wishbone_bd_ram_mem2_reg[161][23]/P0001 , \wishbone_bd_ram_mem2_reg[162][16]/P0001 , \wishbone_bd_ram_mem2_reg[162][17]/P0001 , \wishbone_bd_ram_mem2_reg[162][18]/P0001 , \wishbone_bd_ram_mem2_reg[162][19]/P0001 , \wishbone_bd_ram_mem2_reg[162][20]/P0001 , \wishbone_bd_ram_mem2_reg[162][21]/P0001 , \wishbone_bd_ram_mem2_reg[162][22]/P0001 , \wishbone_bd_ram_mem2_reg[162][23]/P0001 , \wishbone_bd_ram_mem2_reg[163][16]/P0001 , \wishbone_bd_ram_mem2_reg[163][17]/P0001 , \wishbone_bd_ram_mem2_reg[163][18]/P0001 , \wishbone_bd_ram_mem2_reg[163][19]/P0001 , \wishbone_bd_ram_mem2_reg[163][20]/P0001 , \wishbone_bd_ram_mem2_reg[163][21]/P0001 , \wishbone_bd_ram_mem2_reg[163][22]/P0001 , \wishbone_bd_ram_mem2_reg[163][23]/P0001 , \wishbone_bd_ram_mem2_reg[164][16]/P0001 , \wishbone_bd_ram_mem2_reg[164][17]/P0001 , \wishbone_bd_ram_mem2_reg[164][18]/P0001 , \wishbone_bd_ram_mem2_reg[164][19]/P0001 , \wishbone_bd_ram_mem2_reg[164][20]/P0001 , \wishbone_bd_ram_mem2_reg[164][21]/P0001 , \wishbone_bd_ram_mem2_reg[164][22]/P0001 , \wishbone_bd_ram_mem2_reg[164][23]/P0001 , \wishbone_bd_ram_mem2_reg[165][16]/P0001 , \wishbone_bd_ram_mem2_reg[165][17]/P0001 , \wishbone_bd_ram_mem2_reg[165][18]/P0001 , \wishbone_bd_ram_mem2_reg[165][19]/P0001 , \wishbone_bd_ram_mem2_reg[165][20]/P0001 , \wishbone_bd_ram_mem2_reg[165][21]/P0001 , \wishbone_bd_ram_mem2_reg[165][22]/P0001 , \wishbone_bd_ram_mem2_reg[165][23]/P0001 , \wishbone_bd_ram_mem2_reg[166][16]/P0001 , \wishbone_bd_ram_mem2_reg[166][17]/P0001 , \wishbone_bd_ram_mem2_reg[166][18]/P0001 , \wishbone_bd_ram_mem2_reg[166][19]/P0001 , \wishbone_bd_ram_mem2_reg[166][20]/P0001 , \wishbone_bd_ram_mem2_reg[166][21]/P0001 , \wishbone_bd_ram_mem2_reg[166][22]/P0001 , \wishbone_bd_ram_mem2_reg[166][23]/P0001 , \wishbone_bd_ram_mem2_reg[167][16]/P0001 , \wishbone_bd_ram_mem2_reg[167][17]/P0001 , \wishbone_bd_ram_mem2_reg[167][18]/P0001 , \wishbone_bd_ram_mem2_reg[167][19]/P0001 , \wishbone_bd_ram_mem2_reg[167][20]/P0001 , \wishbone_bd_ram_mem2_reg[167][21]/P0001 , \wishbone_bd_ram_mem2_reg[167][22]/P0001 , \wishbone_bd_ram_mem2_reg[167][23]/P0001 , \wishbone_bd_ram_mem2_reg[168][16]/P0001 , \wishbone_bd_ram_mem2_reg[168][17]/P0001 , \wishbone_bd_ram_mem2_reg[168][18]/P0001 , \wishbone_bd_ram_mem2_reg[168][19]/P0001 , \wishbone_bd_ram_mem2_reg[168][20]/P0001 , \wishbone_bd_ram_mem2_reg[168][21]/P0001 , \wishbone_bd_ram_mem2_reg[168][22]/P0001 , \wishbone_bd_ram_mem2_reg[168][23]/P0001 , \wishbone_bd_ram_mem2_reg[169][16]/P0001 , \wishbone_bd_ram_mem2_reg[169][17]/P0001 , \wishbone_bd_ram_mem2_reg[169][18]/P0001 , \wishbone_bd_ram_mem2_reg[169][19]/P0001 , \wishbone_bd_ram_mem2_reg[169][20]/P0001 , \wishbone_bd_ram_mem2_reg[169][21]/P0001 , \wishbone_bd_ram_mem2_reg[169][22]/P0001 , \wishbone_bd_ram_mem2_reg[169][23]/P0001 , \wishbone_bd_ram_mem2_reg[16][16]/P0001 , \wishbone_bd_ram_mem2_reg[16][17]/P0001 , \wishbone_bd_ram_mem2_reg[16][18]/P0001 , \wishbone_bd_ram_mem2_reg[16][19]/P0001 , \wishbone_bd_ram_mem2_reg[16][20]/P0001 , \wishbone_bd_ram_mem2_reg[16][21]/P0001 , \wishbone_bd_ram_mem2_reg[16][22]/P0001 , \wishbone_bd_ram_mem2_reg[16][23]/P0001 , \wishbone_bd_ram_mem2_reg[170][16]/P0001 , \wishbone_bd_ram_mem2_reg[170][17]/P0001 , \wishbone_bd_ram_mem2_reg[170][18]/P0001 , \wishbone_bd_ram_mem2_reg[170][19]/P0001 , \wishbone_bd_ram_mem2_reg[170][20]/P0001 , \wishbone_bd_ram_mem2_reg[170][21]/P0001 , \wishbone_bd_ram_mem2_reg[170][22]/P0001 , \wishbone_bd_ram_mem2_reg[170][23]/P0001 , \wishbone_bd_ram_mem2_reg[171][16]/P0001 , \wishbone_bd_ram_mem2_reg[171][17]/P0001 , \wishbone_bd_ram_mem2_reg[171][18]/P0001 , \wishbone_bd_ram_mem2_reg[171][19]/P0001 , \wishbone_bd_ram_mem2_reg[171][20]/P0001 , \wishbone_bd_ram_mem2_reg[171][21]/P0001 , \wishbone_bd_ram_mem2_reg[171][22]/P0001 , \wishbone_bd_ram_mem2_reg[171][23]/P0001 , \wishbone_bd_ram_mem2_reg[172][16]/P0001 , \wishbone_bd_ram_mem2_reg[172][17]/P0001 , \wishbone_bd_ram_mem2_reg[172][18]/P0001 , \wishbone_bd_ram_mem2_reg[172][19]/P0001 , \wishbone_bd_ram_mem2_reg[172][20]/P0001 , \wishbone_bd_ram_mem2_reg[172][21]/P0001 , \wishbone_bd_ram_mem2_reg[172][22]/P0001 , \wishbone_bd_ram_mem2_reg[172][23]/P0001 , \wishbone_bd_ram_mem2_reg[173][16]/P0001 , \wishbone_bd_ram_mem2_reg[173][17]/P0001 , \wishbone_bd_ram_mem2_reg[173][18]/P0001 , \wishbone_bd_ram_mem2_reg[173][19]/P0001 , \wishbone_bd_ram_mem2_reg[173][20]/P0001 , \wishbone_bd_ram_mem2_reg[173][21]/P0001 , \wishbone_bd_ram_mem2_reg[173][22]/P0001 , \wishbone_bd_ram_mem2_reg[173][23]/P0001 , \wishbone_bd_ram_mem2_reg[174][16]/P0001 , \wishbone_bd_ram_mem2_reg[174][17]/P0001 , \wishbone_bd_ram_mem2_reg[174][18]/P0001 , \wishbone_bd_ram_mem2_reg[174][19]/P0001 , \wishbone_bd_ram_mem2_reg[174][20]/P0001 , \wishbone_bd_ram_mem2_reg[174][21]/P0001 , \wishbone_bd_ram_mem2_reg[174][22]/P0001 , \wishbone_bd_ram_mem2_reg[174][23]/P0001 , \wishbone_bd_ram_mem2_reg[175][16]/P0001 , \wishbone_bd_ram_mem2_reg[175][17]/P0001 , \wishbone_bd_ram_mem2_reg[175][18]/P0001 , \wishbone_bd_ram_mem2_reg[175][19]/P0001 , \wishbone_bd_ram_mem2_reg[175][20]/P0001 , \wishbone_bd_ram_mem2_reg[175][21]/P0001 , \wishbone_bd_ram_mem2_reg[175][22]/P0001 , \wishbone_bd_ram_mem2_reg[175][23]/P0001 , \wishbone_bd_ram_mem2_reg[176][16]/P0001 , \wishbone_bd_ram_mem2_reg[176][17]/P0001 , \wishbone_bd_ram_mem2_reg[176][18]/P0001 , \wishbone_bd_ram_mem2_reg[176][19]/P0001 , \wishbone_bd_ram_mem2_reg[176][20]/P0001 , \wishbone_bd_ram_mem2_reg[176][21]/P0001 , \wishbone_bd_ram_mem2_reg[176][22]/P0001 , \wishbone_bd_ram_mem2_reg[176][23]/P0001 , \wishbone_bd_ram_mem2_reg[177][16]/P0001 , \wishbone_bd_ram_mem2_reg[177][17]/P0001 , \wishbone_bd_ram_mem2_reg[177][18]/P0001 , \wishbone_bd_ram_mem2_reg[177][19]/P0001 , \wishbone_bd_ram_mem2_reg[177][20]/P0001 , \wishbone_bd_ram_mem2_reg[177][21]/P0001 , \wishbone_bd_ram_mem2_reg[177][22]/P0001 , \wishbone_bd_ram_mem2_reg[177][23]/P0001 , \wishbone_bd_ram_mem2_reg[178][16]/P0001 , \wishbone_bd_ram_mem2_reg[178][17]/P0001 , \wishbone_bd_ram_mem2_reg[178][18]/P0001 , \wishbone_bd_ram_mem2_reg[178][19]/P0001 , \wishbone_bd_ram_mem2_reg[178][20]/P0001 , \wishbone_bd_ram_mem2_reg[178][21]/P0001 , \wishbone_bd_ram_mem2_reg[178][22]/P0001 , \wishbone_bd_ram_mem2_reg[178][23]/P0001 , \wishbone_bd_ram_mem2_reg[179][16]/P0001 , \wishbone_bd_ram_mem2_reg[179][17]/P0001 , \wishbone_bd_ram_mem2_reg[179][18]/P0001 , \wishbone_bd_ram_mem2_reg[179][19]/P0001 , \wishbone_bd_ram_mem2_reg[179][20]/P0001 , \wishbone_bd_ram_mem2_reg[179][21]/P0001 , \wishbone_bd_ram_mem2_reg[179][22]/P0001 , \wishbone_bd_ram_mem2_reg[179][23]/P0001 , \wishbone_bd_ram_mem2_reg[17][16]/P0001 , \wishbone_bd_ram_mem2_reg[17][17]/P0001 , \wishbone_bd_ram_mem2_reg[17][18]/P0001 , \wishbone_bd_ram_mem2_reg[17][19]/P0001 , \wishbone_bd_ram_mem2_reg[17][20]/P0001 , \wishbone_bd_ram_mem2_reg[17][21]/P0001 , \wishbone_bd_ram_mem2_reg[17][22]/P0001 , \wishbone_bd_ram_mem2_reg[17][23]/P0001 , \wishbone_bd_ram_mem2_reg[180][16]/P0001 , \wishbone_bd_ram_mem2_reg[180][17]/P0001 , \wishbone_bd_ram_mem2_reg[180][18]/P0001 , \wishbone_bd_ram_mem2_reg[180][19]/P0001 , \wishbone_bd_ram_mem2_reg[180][20]/P0001 , \wishbone_bd_ram_mem2_reg[180][21]/P0001 , \wishbone_bd_ram_mem2_reg[180][22]/P0001 , \wishbone_bd_ram_mem2_reg[180][23]/P0001 , \wishbone_bd_ram_mem2_reg[181][16]/P0001 , \wishbone_bd_ram_mem2_reg[181][17]/P0001 , \wishbone_bd_ram_mem2_reg[181][18]/P0001 , \wishbone_bd_ram_mem2_reg[181][19]/P0001 , \wishbone_bd_ram_mem2_reg[181][20]/P0001 , \wishbone_bd_ram_mem2_reg[181][21]/P0001 , \wishbone_bd_ram_mem2_reg[181][22]/P0001 , \wishbone_bd_ram_mem2_reg[181][23]/P0001 , \wishbone_bd_ram_mem2_reg[182][16]/P0001 , \wishbone_bd_ram_mem2_reg[182][17]/P0001 , \wishbone_bd_ram_mem2_reg[182][18]/P0001 , \wishbone_bd_ram_mem2_reg[182][19]/P0001 , \wishbone_bd_ram_mem2_reg[182][20]/P0001 , \wishbone_bd_ram_mem2_reg[182][21]/P0001 , \wishbone_bd_ram_mem2_reg[182][22]/P0001 , \wishbone_bd_ram_mem2_reg[182][23]/P0001 , \wishbone_bd_ram_mem2_reg[183][16]/P0001 , \wishbone_bd_ram_mem2_reg[183][17]/P0001 , \wishbone_bd_ram_mem2_reg[183][18]/P0001 , \wishbone_bd_ram_mem2_reg[183][19]/P0001 , \wishbone_bd_ram_mem2_reg[183][20]/P0001 , \wishbone_bd_ram_mem2_reg[183][21]/P0001 , \wishbone_bd_ram_mem2_reg[183][22]/P0001 , \wishbone_bd_ram_mem2_reg[183][23]/P0001 , \wishbone_bd_ram_mem2_reg[184][16]/P0001 , \wishbone_bd_ram_mem2_reg[184][17]/P0001 , \wishbone_bd_ram_mem2_reg[184][18]/P0001 , \wishbone_bd_ram_mem2_reg[184][19]/P0001 , \wishbone_bd_ram_mem2_reg[184][20]/P0001 , \wishbone_bd_ram_mem2_reg[184][21]/P0001 , \wishbone_bd_ram_mem2_reg[184][22]/P0001 , \wishbone_bd_ram_mem2_reg[184][23]/P0001 , \wishbone_bd_ram_mem2_reg[185][16]/P0001 , \wishbone_bd_ram_mem2_reg[185][17]/P0001 , \wishbone_bd_ram_mem2_reg[185][18]/P0001 , \wishbone_bd_ram_mem2_reg[185][19]/P0001 , \wishbone_bd_ram_mem2_reg[185][20]/P0001 , \wishbone_bd_ram_mem2_reg[185][21]/P0001 , \wishbone_bd_ram_mem2_reg[185][22]/P0001 , \wishbone_bd_ram_mem2_reg[185][23]/P0001 , \wishbone_bd_ram_mem2_reg[186][16]/P0001 , \wishbone_bd_ram_mem2_reg[186][17]/P0001 , \wishbone_bd_ram_mem2_reg[186][18]/P0001 , \wishbone_bd_ram_mem2_reg[186][19]/P0001 , \wishbone_bd_ram_mem2_reg[186][20]/P0001 , \wishbone_bd_ram_mem2_reg[186][21]/P0001 , \wishbone_bd_ram_mem2_reg[186][22]/P0001 , \wishbone_bd_ram_mem2_reg[186][23]/P0001 , \wishbone_bd_ram_mem2_reg[187][16]/P0001 , \wishbone_bd_ram_mem2_reg[187][17]/P0001 , \wishbone_bd_ram_mem2_reg[187][18]/P0001 , \wishbone_bd_ram_mem2_reg[187][19]/P0001 , \wishbone_bd_ram_mem2_reg[187][20]/P0001 , \wishbone_bd_ram_mem2_reg[187][21]/P0001 , \wishbone_bd_ram_mem2_reg[187][22]/P0001 , \wishbone_bd_ram_mem2_reg[187][23]/P0001 , \wishbone_bd_ram_mem2_reg[188][16]/P0001 , \wishbone_bd_ram_mem2_reg[188][17]/P0001 , \wishbone_bd_ram_mem2_reg[188][18]/P0001 , \wishbone_bd_ram_mem2_reg[188][19]/P0001 , \wishbone_bd_ram_mem2_reg[188][20]/P0001 , \wishbone_bd_ram_mem2_reg[188][21]/P0001 , \wishbone_bd_ram_mem2_reg[188][22]/P0001 , \wishbone_bd_ram_mem2_reg[188][23]/P0001 , \wishbone_bd_ram_mem2_reg[189][16]/P0001 , \wishbone_bd_ram_mem2_reg[189][17]/P0001 , \wishbone_bd_ram_mem2_reg[189][18]/P0001 , \wishbone_bd_ram_mem2_reg[189][19]/P0001 , \wishbone_bd_ram_mem2_reg[189][20]/P0001 , \wishbone_bd_ram_mem2_reg[189][21]/P0001 , \wishbone_bd_ram_mem2_reg[189][22]/P0001 , \wishbone_bd_ram_mem2_reg[189][23]/P0001 , \wishbone_bd_ram_mem2_reg[18][16]/P0001 , \wishbone_bd_ram_mem2_reg[18][17]/P0001 , \wishbone_bd_ram_mem2_reg[18][18]/P0001 , \wishbone_bd_ram_mem2_reg[18][19]/P0001 , \wishbone_bd_ram_mem2_reg[18][20]/P0001 , \wishbone_bd_ram_mem2_reg[18][21]/P0001 , \wishbone_bd_ram_mem2_reg[18][22]/P0001 , \wishbone_bd_ram_mem2_reg[18][23]/P0001 , \wishbone_bd_ram_mem2_reg[190][16]/P0001 , \wishbone_bd_ram_mem2_reg[190][17]/P0001 , \wishbone_bd_ram_mem2_reg[190][18]/P0001 , \wishbone_bd_ram_mem2_reg[190][19]/P0001 , \wishbone_bd_ram_mem2_reg[190][20]/P0001 , \wishbone_bd_ram_mem2_reg[190][21]/P0001 , \wishbone_bd_ram_mem2_reg[190][22]/P0001 , \wishbone_bd_ram_mem2_reg[190][23]/P0001 , \wishbone_bd_ram_mem2_reg[191][16]/P0001 , \wishbone_bd_ram_mem2_reg[191][17]/P0001 , \wishbone_bd_ram_mem2_reg[191][18]/P0001 , \wishbone_bd_ram_mem2_reg[191][19]/P0001 , \wishbone_bd_ram_mem2_reg[191][20]/P0001 , \wishbone_bd_ram_mem2_reg[191][21]/P0001 , \wishbone_bd_ram_mem2_reg[191][22]/P0001 , \wishbone_bd_ram_mem2_reg[191][23]/P0001 , \wishbone_bd_ram_mem2_reg[192][16]/P0001 , \wishbone_bd_ram_mem2_reg[192][17]/P0001 , \wishbone_bd_ram_mem2_reg[192][18]/P0001 , \wishbone_bd_ram_mem2_reg[192][19]/P0001 , \wishbone_bd_ram_mem2_reg[192][20]/P0001 , \wishbone_bd_ram_mem2_reg[192][21]/P0001 , \wishbone_bd_ram_mem2_reg[192][22]/P0001 , \wishbone_bd_ram_mem2_reg[192][23]/P0001 , \wishbone_bd_ram_mem2_reg[193][16]/P0001 , \wishbone_bd_ram_mem2_reg[193][17]/P0001 , \wishbone_bd_ram_mem2_reg[193][18]/P0001 , \wishbone_bd_ram_mem2_reg[193][19]/P0001 , \wishbone_bd_ram_mem2_reg[193][20]/P0001 , \wishbone_bd_ram_mem2_reg[193][21]/P0001 , \wishbone_bd_ram_mem2_reg[193][22]/P0001 , \wishbone_bd_ram_mem2_reg[193][23]/P0001 , \wishbone_bd_ram_mem2_reg[194][16]/P0001 , \wishbone_bd_ram_mem2_reg[194][17]/P0001 , \wishbone_bd_ram_mem2_reg[194][18]/P0001 , \wishbone_bd_ram_mem2_reg[194][19]/P0001 , \wishbone_bd_ram_mem2_reg[194][20]/P0001 , \wishbone_bd_ram_mem2_reg[194][21]/P0001 , \wishbone_bd_ram_mem2_reg[194][22]/P0001 , \wishbone_bd_ram_mem2_reg[194][23]/P0001 , \wishbone_bd_ram_mem2_reg[195][16]/P0001 , \wishbone_bd_ram_mem2_reg[195][17]/P0001 , \wishbone_bd_ram_mem2_reg[195][18]/P0001 , \wishbone_bd_ram_mem2_reg[195][19]/P0001 , \wishbone_bd_ram_mem2_reg[195][20]/P0001 , \wishbone_bd_ram_mem2_reg[195][21]/P0001 , \wishbone_bd_ram_mem2_reg[195][22]/P0001 , \wishbone_bd_ram_mem2_reg[195][23]/P0001 , \wishbone_bd_ram_mem2_reg[196][16]/P0001 , \wishbone_bd_ram_mem2_reg[196][17]/P0001 , \wishbone_bd_ram_mem2_reg[196][18]/P0001 , \wishbone_bd_ram_mem2_reg[196][19]/P0001 , \wishbone_bd_ram_mem2_reg[196][20]/P0001 , \wishbone_bd_ram_mem2_reg[196][21]/P0001 , \wishbone_bd_ram_mem2_reg[196][22]/P0001 , \wishbone_bd_ram_mem2_reg[196][23]/P0001 , \wishbone_bd_ram_mem2_reg[197][16]/P0001 , \wishbone_bd_ram_mem2_reg[197][17]/P0001 , \wishbone_bd_ram_mem2_reg[197][18]/P0001 , \wishbone_bd_ram_mem2_reg[197][19]/P0001 , \wishbone_bd_ram_mem2_reg[197][20]/P0001 , \wishbone_bd_ram_mem2_reg[197][21]/P0001 , \wishbone_bd_ram_mem2_reg[197][22]/P0001 , \wishbone_bd_ram_mem2_reg[197][23]/P0001 , \wishbone_bd_ram_mem2_reg[198][16]/P0001 , \wishbone_bd_ram_mem2_reg[198][17]/P0001 , \wishbone_bd_ram_mem2_reg[198][18]/P0001 , \wishbone_bd_ram_mem2_reg[198][19]/P0001 , \wishbone_bd_ram_mem2_reg[198][20]/P0001 , \wishbone_bd_ram_mem2_reg[198][21]/P0001 , \wishbone_bd_ram_mem2_reg[198][22]/P0001 , \wishbone_bd_ram_mem2_reg[198][23]/P0001 , \wishbone_bd_ram_mem2_reg[199][16]/P0001 , \wishbone_bd_ram_mem2_reg[199][17]/P0001 , \wishbone_bd_ram_mem2_reg[199][18]/P0001 , \wishbone_bd_ram_mem2_reg[199][19]/P0001 , \wishbone_bd_ram_mem2_reg[199][20]/P0001 , \wishbone_bd_ram_mem2_reg[199][21]/P0001 , \wishbone_bd_ram_mem2_reg[199][22]/P0001 , \wishbone_bd_ram_mem2_reg[199][23]/P0001 , \wishbone_bd_ram_mem2_reg[19][16]/P0001 , \wishbone_bd_ram_mem2_reg[19][17]/P0001 , \wishbone_bd_ram_mem2_reg[19][18]/P0001 , \wishbone_bd_ram_mem2_reg[19][19]/P0001 , \wishbone_bd_ram_mem2_reg[19][20]/P0001 , \wishbone_bd_ram_mem2_reg[19][21]/P0001 , \wishbone_bd_ram_mem2_reg[19][22]/P0001 , \wishbone_bd_ram_mem2_reg[19][23]/P0001 , \wishbone_bd_ram_mem2_reg[1][16]/P0001 , \wishbone_bd_ram_mem2_reg[1][17]/P0001 , \wishbone_bd_ram_mem2_reg[1][18]/P0001 , \wishbone_bd_ram_mem2_reg[1][19]/P0001 , \wishbone_bd_ram_mem2_reg[1][20]/P0001 , \wishbone_bd_ram_mem2_reg[1][21]/P0001 , \wishbone_bd_ram_mem2_reg[1][22]/P0001 , \wishbone_bd_ram_mem2_reg[1][23]/P0001 , \wishbone_bd_ram_mem2_reg[200][16]/P0001 , \wishbone_bd_ram_mem2_reg[200][17]/P0001 , \wishbone_bd_ram_mem2_reg[200][18]/P0001 , \wishbone_bd_ram_mem2_reg[200][19]/P0001 , \wishbone_bd_ram_mem2_reg[200][20]/P0001 , \wishbone_bd_ram_mem2_reg[200][21]/P0001 , \wishbone_bd_ram_mem2_reg[200][22]/P0001 , \wishbone_bd_ram_mem2_reg[200][23]/P0001 , \wishbone_bd_ram_mem2_reg[201][16]/P0001 , \wishbone_bd_ram_mem2_reg[201][17]/P0001 , \wishbone_bd_ram_mem2_reg[201][18]/P0001 , \wishbone_bd_ram_mem2_reg[201][19]/P0001 , \wishbone_bd_ram_mem2_reg[201][20]/P0001 , \wishbone_bd_ram_mem2_reg[201][21]/P0001 , \wishbone_bd_ram_mem2_reg[201][22]/P0001 , \wishbone_bd_ram_mem2_reg[201][23]/P0001 , \wishbone_bd_ram_mem2_reg[202][16]/P0001 , \wishbone_bd_ram_mem2_reg[202][17]/P0001 , \wishbone_bd_ram_mem2_reg[202][18]/P0001 , \wishbone_bd_ram_mem2_reg[202][19]/P0001 , \wishbone_bd_ram_mem2_reg[202][20]/P0001 , \wishbone_bd_ram_mem2_reg[202][21]/P0001 , \wishbone_bd_ram_mem2_reg[202][22]/P0001 , \wishbone_bd_ram_mem2_reg[202][23]/P0001 , \wishbone_bd_ram_mem2_reg[203][16]/P0001 , \wishbone_bd_ram_mem2_reg[203][17]/P0001 , \wishbone_bd_ram_mem2_reg[203][18]/P0001 , \wishbone_bd_ram_mem2_reg[203][19]/P0001 , \wishbone_bd_ram_mem2_reg[203][20]/P0001 , \wishbone_bd_ram_mem2_reg[203][21]/P0001 , \wishbone_bd_ram_mem2_reg[203][22]/P0001 , \wishbone_bd_ram_mem2_reg[203][23]/P0001 , \wishbone_bd_ram_mem2_reg[204][16]/P0001 , \wishbone_bd_ram_mem2_reg[204][17]/P0001 , \wishbone_bd_ram_mem2_reg[204][18]/P0001 , \wishbone_bd_ram_mem2_reg[204][19]/P0001 , \wishbone_bd_ram_mem2_reg[204][20]/P0001 , \wishbone_bd_ram_mem2_reg[204][21]/P0001 , \wishbone_bd_ram_mem2_reg[204][22]/P0001 , \wishbone_bd_ram_mem2_reg[204][23]/P0001 , \wishbone_bd_ram_mem2_reg[205][16]/P0001 , \wishbone_bd_ram_mem2_reg[205][17]/P0001 , \wishbone_bd_ram_mem2_reg[205][18]/P0001 , \wishbone_bd_ram_mem2_reg[205][19]/P0001 , \wishbone_bd_ram_mem2_reg[205][20]/P0001 , \wishbone_bd_ram_mem2_reg[205][21]/P0001 , \wishbone_bd_ram_mem2_reg[205][22]/P0001 , \wishbone_bd_ram_mem2_reg[205][23]/P0001 , \wishbone_bd_ram_mem2_reg[206][16]/P0001 , \wishbone_bd_ram_mem2_reg[206][17]/P0001 , \wishbone_bd_ram_mem2_reg[206][18]/P0001 , \wishbone_bd_ram_mem2_reg[206][19]/P0001 , \wishbone_bd_ram_mem2_reg[206][20]/P0001 , \wishbone_bd_ram_mem2_reg[206][21]/P0001 , \wishbone_bd_ram_mem2_reg[206][22]/P0001 , \wishbone_bd_ram_mem2_reg[206][23]/P0001 , \wishbone_bd_ram_mem2_reg[207][16]/P0001 , \wishbone_bd_ram_mem2_reg[207][17]/P0001 , \wishbone_bd_ram_mem2_reg[207][18]/P0001 , \wishbone_bd_ram_mem2_reg[207][19]/P0001 , \wishbone_bd_ram_mem2_reg[207][20]/P0001 , \wishbone_bd_ram_mem2_reg[207][21]/P0001 , \wishbone_bd_ram_mem2_reg[207][22]/P0001 , \wishbone_bd_ram_mem2_reg[207][23]/P0001 , \wishbone_bd_ram_mem2_reg[208][16]/P0001 , \wishbone_bd_ram_mem2_reg[208][17]/P0001 , \wishbone_bd_ram_mem2_reg[208][18]/P0001 , \wishbone_bd_ram_mem2_reg[208][19]/P0001 , \wishbone_bd_ram_mem2_reg[208][20]/P0001 , \wishbone_bd_ram_mem2_reg[208][21]/P0001 , \wishbone_bd_ram_mem2_reg[208][22]/P0001 , \wishbone_bd_ram_mem2_reg[208][23]/P0001 , \wishbone_bd_ram_mem2_reg[209][16]/P0001 , \wishbone_bd_ram_mem2_reg[209][17]/P0001 , \wishbone_bd_ram_mem2_reg[209][18]/P0001 , \wishbone_bd_ram_mem2_reg[209][19]/P0001 , \wishbone_bd_ram_mem2_reg[209][20]/P0001 , \wishbone_bd_ram_mem2_reg[209][21]/P0001 , \wishbone_bd_ram_mem2_reg[209][22]/P0001 , \wishbone_bd_ram_mem2_reg[209][23]/P0001 , \wishbone_bd_ram_mem2_reg[20][16]/P0001 , \wishbone_bd_ram_mem2_reg[20][17]/P0001 , \wishbone_bd_ram_mem2_reg[20][18]/P0001 , \wishbone_bd_ram_mem2_reg[20][19]/P0001 , \wishbone_bd_ram_mem2_reg[20][20]/P0001 , \wishbone_bd_ram_mem2_reg[20][21]/P0001 , \wishbone_bd_ram_mem2_reg[20][22]/P0001 , \wishbone_bd_ram_mem2_reg[20][23]/P0001 , \wishbone_bd_ram_mem2_reg[210][16]/P0001 , \wishbone_bd_ram_mem2_reg[210][17]/P0001 , \wishbone_bd_ram_mem2_reg[210][18]/P0001 , \wishbone_bd_ram_mem2_reg[210][19]/P0001 , \wishbone_bd_ram_mem2_reg[210][20]/P0001 , \wishbone_bd_ram_mem2_reg[210][21]/P0001 , \wishbone_bd_ram_mem2_reg[210][22]/P0001 , \wishbone_bd_ram_mem2_reg[210][23]/P0001 , \wishbone_bd_ram_mem2_reg[211][16]/P0001 , \wishbone_bd_ram_mem2_reg[211][17]/P0001 , \wishbone_bd_ram_mem2_reg[211][18]/P0001 , \wishbone_bd_ram_mem2_reg[211][19]/P0001 , \wishbone_bd_ram_mem2_reg[211][20]/P0001 , \wishbone_bd_ram_mem2_reg[211][21]/P0001 , \wishbone_bd_ram_mem2_reg[211][22]/P0001 , \wishbone_bd_ram_mem2_reg[211][23]/P0001 , \wishbone_bd_ram_mem2_reg[212][16]/P0001 , \wishbone_bd_ram_mem2_reg[212][17]/P0001 , \wishbone_bd_ram_mem2_reg[212][18]/P0001 , \wishbone_bd_ram_mem2_reg[212][19]/P0001 , \wishbone_bd_ram_mem2_reg[212][20]/P0001 , \wishbone_bd_ram_mem2_reg[212][21]/P0001 , \wishbone_bd_ram_mem2_reg[212][22]/P0001 , \wishbone_bd_ram_mem2_reg[212][23]/P0001 , \wishbone_bd_ram_mem2_reg[213][16]/P0001 , \wishbone_bd_ram_mem2_reg[213][17]/P0001 , \wishbone_bd_ram_mem2_reg[213][18]/P0001 , \wishbone_bd_ram_mem2_reg[213][19]/P0001 , \wishbone_bd_ram_mem2_reg[213][20]/P0001 , \wishbone_bd_ram_mem2_reg[213][21]/P0001 , \wishbone_bd_ram_mem2_reg[213][22]/P0001 , \wishbone_bd_ram_mem2_reg[213][23]/P0001 , \wishbone_bd_ram_mem2_reg[214][16]/P0001 , \wishbone_bd_ram_mem2_reg[214][17]/P0001 , \wishbone_bd_ram_mem2_reg[214][18]/P0001 , \wishbone_bd_ram_mem2_reg[214][19]/P0001 , \wishbone_bd_ram_mem2_reg[214][20]/P0001 , \wishbone_bd_ram_mem2_reg[214][21]/P0001 , \wishbone_bd_ram_mem2_reg[214][22]/P0001 , \wishbone_bd_ram_mem2_reg[214][23]/P0001 , \wishbone_bd_ram_mem2_reg[215][16]/P0001 , \wishbone_bd_ram_mem2_reg[215][17]/P0001 , \wishbone_bd_ram_mem2_reg[215][18]/P0001 , \wishbone_bd_ram_mem2_reg[215][19]/P0001 , \wishbone_bd_ram_mem2_reg[215][20]/P0001 , \wishbone_bd_ram_mem2_reg[215][21]/P0001 , \wishbone_bd_ram_mem2_reg[215][22]/P0001 , \wishbone_bd_ram_mem2_reg[215][23]/P0001 , \wishbone_bd_ram_mem2_reg[216][16]/P0001 , \wishbone_bd_ram_mem2_reg[216][17]/P0001 , \wishbone_bd_ram_mem2_reg[216][18]/P0001 , \wishbone_bd_ram_mem2_reg[216][19]/P0001 , \wishbone_bd_ram_mem2_reg[216][20]/P0001 , \wishbone_bd_ram_mem2_reg[216][21]/P0001 , \wishbone_bd_ram_mem2_reg[216][22]/P0001 , \wishbone_bd_ram_mem2_reg[216][23]/P0001 , \wishbone_bd_ram_mem2_reg[217][16]/P0001 , \wishbone_bd_ram_mem2_reg[217][17]/P0001 , \wishbone_bd_ram_mem2_reg[217][18]/P0001 , \wishbone_bd_ram_mem2_reg[217][19]/P0001 , \wishbone_bd_ram_mem2_reg[217][20]/P0001 , \wishbone_bd_ram_mem2_reg[217][21]/P0001 , \wishbone_bd_ram_mem2_reg[217][22]/P0001 , \wishbone_bd_ram_mem2_reg[217][23]/P0001 , \wishbone_bd_ram_mem2_reg[218][16]/P0001 , \wishbone_bd_ram_mem2_reg[218][17]/P0001 , \wishbone_bd_ram_mem2_reg[218][18]/P0001 , \wishbone_bd_ram_mem2_reg[218][19]/P0001 , \wishbone_bd_ram_mem2_reg[218][20]/P0001 , \wishbone_bd_ram_mem2_reg[218][21]/P0001 , \wishbone_bd_ram_mem2_reg[218][22]/P0001 , \wishbone_bd_ram_mem2_reg[218][23]/P0001 , \wishbone_bd_ram_mem2_reg[219][16]/P0001 , \wishbone_bd_ram_mem2_reg[219][17]/P0001 , \wishbone_bd_ram_mem2_reg[219][18]/P0001 , \wishbone_bd_ram_mem2_reg[219][19]/P0001 , \wishbone_bd_ram_mem2_reg[219][20]/P0001 , \wishbone_bd_ram_mem2_reg[219][21]/P0001 , \wishbone_bd_ram_mem2_reg[219][22]/P0001 , \wishbone_bd_ram_mem2_reg[219][23]/P0001 , \wishbone_bd_ram_mem2_reg[21][16]/P0001 , \wishbone_bd_ram_mem2_reg[21][17]/P0001 , \wishbone_bd_ram_mem2_reg[21][18]/P0001 , \wishbone_bd_ram_mem2_reg[21][19]/P0001 , \wishbone_bd_ram_mem2_reg[21][20]/P0001 , \wishbone_bd_ram_mem2_reg[21][21]/P0001 , \wishbone_bd_ram_mem2_reg[21][22]/P0001 , \wishbone_bd_ram_mem2_reg[21][23]/P0001 , \wishbone_bd_ram_mem2_reg[220][16]/P0001 , \wishbone_bd_ram_mem2_reg[220][17]/P0001 , \wishbone_bd_ram_mem2_reg[220][18]/P0001 , \wishbone_bd_ram_mem2_reg[220][19]/P0001 , \wishbone_bd_ram_mem2_reg[220][20]/P0001 , \wishbone_bd_ram_mem2_reg[220][21]/P0001 , \wishbone_bd_ram_mem2_reg[220][22]/P0001 , \wishbone_bd_ram_mem2_reg[220][23]/P0001 , \wishbone_bd_ram_mem2_reg[221][16]/P0001 , \wishbone_bd_ram_mem2_reg[221][17]/P0001 , \wishbone_bd_ram_mem2_reg[221][18]/P0001 , \wishbone_bd_ram_mem2_reg[221][19]/P0001 , \wishbone_bd_ram_mem2_reg[221][20]/P0001 , \wishbone_bd_ram_mem2_reg[221][21]/P0001 , \wishbone_bd_ram_mem2_reg[221][22]/P0001 , \wishbone_bd_ram_mem2_reg[221][23]/P0001 , \wishbone_bd_ram_mem2_reg[222][16]/P0001 , \wishbone_bd_ram_mem2_reg[222][17]/P0001 , \wishbone_bd_ram_mem2_reg[222][18]/P0001 , \wishbone_bd_ram_mem2_reg[222][19]/P0001 , \wishbone_bd_ram_mem2_reg[222][20]/P0001 , \wishbone_bd_ram_mem2_reg[222][21]/P0001 , \wishbone_bd_ram_mem2_reg[222][22]/P0001 , \wishbone_bd_ram_mem2_reg[222][23]/P0001 , \wishbone_bd_ram_mem2_reg[223][16]/P0001 , \wishbone_bd_ram_mem2_reg[223][17]/P0001 , \wishbone_bd_ram_mem2_reg[223][18]/P0001 , \wishbone_bd_ram_mem2_reg[223][19]/P0001 , \wishbone_bd_ram_mem2_reg[223][20]/P0001 , \wishbone_bd_ram_mem2_reg[223][21]/P0001 , \wishbone_bd_ram_mem2_reg[223][22]/P0001 , \wishbone_bd_ram_mem2_reg[223][23]/P0001 , \wishbone_bd_ram_mem2_reg[224][16]/P0001 , \wishbone_bd_ram_mem2_reg[224][17]/P0001 , \wishbone_bd_ram_mem2_reg[224][18]/P0001 , \wishbone_bd_ram_mem2_reg[224][19]/P0001 , \wishbone_bd_ram_mem2_reg[224][20]/P0001 , \wishbone_bd_ram_mem2_reg[224][21]/P0001 , \wishbone_bd_ram_mem2_reg[224][22]/P0001 , \wishbone_bd_ram_mem2_reg[224][23]/P0001 , \wishbone_bd_ram_mem2_reg[225][16]/P0001 , \wishbone_bd_ram_mem2_reg[225][17]/P0001 , \wishbone_bd_ram_mem2_reg[225][18]/P0001 , \wishbone_bd_ram_mem2_reg[225][19]/P0001 , \wishbone_bd_ram_mem2_reg[225][20]/P0001 , \wishbone_bd_ram_mem2_reg[225][21]/P0001 , \wishbone_bd_ram_mem2_reg[225][22]/P0001 , \wishbone_bd_ram_mem2_reg[225][23]/P0001 , \wishbone_bd_ram_mem2_reg[226][16]/P0001 , \wishbone_bd_ram_mem2_reg[226][17]/P0001 , \wishbone_bd_ram_mem2_reg[226][18]/P0001 , \wishbone_bd_ram_mem2_reg[226][19]/P0001 , \wishbone_bd_ram_mem2_reg[226][20]/P0001 , \wishbone_bd_ram_mem2_reg[226][21]/P0001 , \wishbone_bd_ram_mem2_reg[226][22]/P0001 , \wishbone_bd_ram_mem2_reg[226][23]/P0001 , \wishbone_bd_ram_mem2_reg[227][16]/P0001 , \wishbone_bd_ram_mem2_reg[227][17]/P0001 , \wishbone_bd_ram_mem2_reg[227][18]/P0001 , \wishbone_bd_ram_mem2_reg[227][19]/P0001 , \wishbone_bd_ram_mem2_reg[227][20]/P0001 , \wishbone_bd_ram_mem2_reg[227][21]/P0001 , \wishbone_bd_ram_mem2_reg[227][22]/P0001 , \wishbone_bd_ram_mem2_reg[227][23]/P0001 , \wishbone_bd_ram_mem2_reg[228][16]/P0001 , \wishbone_bd_ram_mem2_reg[228][17]/P0001 , \wishbone_bd_ram_mem2_reg[228][18]/P0001 , \wishbone_bd_ram_mem2_reg[228][19]/P0001 , \wishbone_bd_ram_mem2_reg[228][20]/P0001 , \wishbone_bd_ram_mem2_reg[228][21]/P0001 , \wishbone_bd_ram_mem2_reg[228][22]/P0001 , \wishbone_bd_ram_mem2_reg[228][23]/P0001 , \wishbone_bd_ram_mem2_reg[229][16]/P0001 , \wishbone_bd_ram_mem2_reg[229][17]/P0001 , \wishbone_bd_ram_mem2_reg[229][18]/P0001 , \wishbone_bd_ram_mem2_reg[229][19]/P0001 , \wishbone_bd_ram_mem2_reg[229][20]/P0001 , \wishbone_bd_ram_mem2_reg[229][21]/P0001 , \wishbone_bd_ram_mem2_reg[229][22]/P0001 , \wishbone_bd_ram_mem2_reg[229][23]/P0001 , \wishbone_bd_ram_mem2_reg[22][16]/P0001 , \wishbone_bd_ram_mem2_reg[22][17]/P0001 , \wishbone_bd_ram_mem2_reg[22][18]/P0001 , \wishbone_bd_ram_mem2_reg[22][19]/P0001 , \wishbone_bd_ram_mem2_reg[22][20]/P0001 , \wishbone_bd_ram_mem2_reg[22][21]/P0001 , \wishbone_bd_ram_mem2_reg[22][22]/P0001 , \wishbone_bd_ram_mem2_reg[22][23]/P0001 , \wishbone_bd_ram_mem2_reg[230][16]/P0001 , \wishbone_bd_ram_mem2_reg[230][17]/P0001 , \wishbone_bd_ram_mem2_reg[230][18]/P0001 , \wishbone_bd_ram_mem2_reg[230][19]/P0001 , \wishbone_bd_ram_mem2_reg[230][20]/P0001 , \wishbone_bd_ram_mem2_reg[230][21]/P0001 , \wishbone_bd_ram_mem2_reg[230][22]/P0001 , \wishbone_bd_ram_mem2_reg[230][23]/P0001 , \wishbone_bd_ram_mem2_reg[231][16]/P0001 , \wishbone_bd_ram_mem2_reg[231][17]/P0001 , \wishbone_bd_ram_mem2_reg[231][18]/P0001 , \wishbone_bd_ram_mem2_reg[231][19]/P0001 , \wishbone_bd_ram_mem2_reg[231][20]/P0001 , \wishbone_bd_ram_mem2_reg[231][21]/P0001 , \wishbone_bd_ram_mem2_reg[231][22]/P0001 , \wishbone_bd_ram_mem2_reg[231][23]/P0001 , \wishbone_bd_ram_mem2_reg[232][16]/P0001 , \wishbone_bd_ram_mem2_reg[232][17]/P0001 , \wishbone_bd_ram_mem2_reg[232][18]/P0001 , \wishbone_bd_ram_mem2_reg[232][19]/P0001 , \wishbone_bd_ram_mem2_reg[232][20]/P0001 , \wishbone_bd_ram_mem2_reg[232][21]/P0001 , \wishbone_bd_ram_mem2_reg[232][22]/P0001 , \wishbone_bd_ram_mem2_reg[232][23]/P0001 , \wishbone_bd_ram_mem2_reg[233][16]/P0001 , \wishbone_bd_ram_mem2_reg[233][17]/P0001 , \wishbone_bd_ram_mem2_reg[233][18]/P0001 , \wishbone_bd_ram_mem2_reg[233][19]/P0001 , \wishbone_bd_ram_mem2_reg[233][20]/P0001 , \wishbone_bd_ram_mem2_reg[233][21]/P0001 , \wishbone_bd_ram_mem2_reg[233][22]/P0001 , \wishbone_bd_ram_mem2_reg[233][23]/P0001 , \wishbone_bd_ram_mem2_reg[234][16]/P0001 , \wishbone_bd_ram_mem2_reg[234][17]/P0001 , \wishbone_bd_ram_mem2_reg[234][18]/P0001 , \wishbone_bd_ram_mem2_reg[234][19]/P0001 , \wishbone_bd_ram_mem2_reg[234][20]/P0001 , \wishbone_bd_ram_mem2_reg[234][21]/P0001 , \wishbone_bd_ram_mem2_reg[234][22]/P0001 , \wishbone_bd_ram_mem2_reg[234][23]/P0001 , \wishbone_bd_ram_mem2_reg[235][16]/P0001 , \wishbone_bd_ram_mem2_reg[235][17]/P0001 , \wishbone_bd_ram_mem2_reg[235][18]/P0001 , \wishbone_bd_ram_mem2_reg[235][19]/P0001 , \wishbone_bd_ram_mem2_reg[235][20]/P0001 , \wishbone_bd_ram_mem2_reg[235][21]/P0001 , \wishbone_bd_ram_mem2_reg[235][22]/P0001 , \wishbone_bd_ram_mem2_reg[235][23]/P0001 , \wishbone_bd_ram_mem2_reg[236][16]/P0001 , \wishbone_bd_ram_mem2_reg[236][17]/P0001 , \wishbone_bd_ram_mem2_reg[236][18]/P0001 , \wishbone_bd_ram_mem2_reg[236][19]/P0001 , \wishbone_bd_ram_mem2_reg[236][20]/P0001 , \wishbone_bd_ram_mem2_reg[236][21]/P0001 , \wishbone_bd_ram_mem2_reg[236][22]/P0001 , \wishbone_bd_ram_mem2_reg[236][23]/P0001 , \wishbone_bd_ram_mem2_reg[237][16]/P0001 , \wishbone_bd_ram_mem2_reg[237][17]/P0001 , \wishbone_bd_ram_mem2_reg[237][18]/P0001 , \wishbone_bd_ram_mem2_reg[237][19]/P0001 , \wishbone_bd_ram_mem2_reg[237][20]/P0001 , \wishbone_bd_ram_mem2_reg[237][21]/P0001 , \wishbone_bd_ram_mem2_reg[237][22]/P0001 , \wishbone_bd_ram_mem2_reg[237][23]/P0001 , \wishbone_bd_ram_mem2_reg[238][16]/P0001 , \wishbone_bd_ram_mem2_reg[238][17]/P0001 , \wishbone_bd_ram_mem2_reg[238][18]/P0001 , \wishbone_bd_ram_mem2_reg[238][19]/P0001 , \wishbone_bd_ram_mem2_reg[238][20]/P0001 , \wishbone_bd_ram_mem2_reg[238][21]/P0001 , \wishbone_bd_ram_mem2_reg[238][22]/P0001 , \wishbone_bd_ram_mem2_reg[238][23]/P0001 , \wishbone_bd_ram_mem2_reg[239][16]/P0001 , \wishbone_bd_ram_mem2_reg[239][17]/P0001 , \wishbone_bd_ram_mem2_reg[239][18]/P0001 , \wishbone_bd_ram_mem2_reg[239][19]/P0001 , \wishbone_bd_ram_mem2_reg[239][20]/P0001 , \wishbone_bd_ram_mem2_reg[239][21]/P0001 , \wishbone_bd_ram_mem2_reg[239][22]/P0001 , \wishbone_bd_ram_mem2_reg[239][23]/P0001 , \wishbone_bd_ram_mem2_reg[23][16]/P0001 , \wishbone_bd_ram_mem2_reg[23][17]/P0001 , \wishbone_bd_ram_mem2_reg[23][18]/P0001 , \wishbone_bd_ram_mem2_reg[23][19]/P0001 , \wishbone_bd_ram_mem2_reg[23][20]/P0001 , \wishbone_bd_ram_mem2_reg[23][21]/P0001 , \wishbone_bd_ram_mem2_reg[23][22]/P0001 , \wishbone_bd_ram_mem2_reg[23][23]/P0001 , \wishbone_bd_ram_mem2_reg[240][16]/P0001 , \wishbone_bd_ram_mem2_reg[240][17]/P0001 , \wishbone_bd_ram_mem2_reg[240][18]/P0001 , \wishbone_bd_ram_mem2_reg[240][19]/P0001 , \wishbone_bd_ram_mem2_reg[240][20]/P0001 , \wishbone_bd_ram_mem2_reg[240][21]/P0001 , \wishbone_bd_ram_mem2_reg[240][22]/P0001 , \wishbone_bd_ram_mem2_reg[240][23]/P0001 , \wishbone_bd_ram_mem2_reg[241][16]/P0001 , \wishbone_bd_ram_mem2_reg[241][17]/P0001 , \wishbone_bd_ram_mem2_reg[241][18]/P0001 , \wishbone_bd_ram_mem2_reg[241][19]/P0001 , \wishbone_bd_ram_mem2_reg[241][20]/P0001 , \wishbone_bd_ram_mem2_reg[241][21]/P0001 , \wishbone_bd_ram_mem2_reg[241][22]/P0001 , \wishbone_bd_ram_mem2_reg[241][23]/P0001 , \wishbone_bd_ram_mem2_reg[242][16]/P0001 , \wishbone_bd_ram_mem2_reg[242][17]/P0001 , \wishbone_bd_ram_mem2_reg[242][18]/P0001 , \wishbone_bd_ram_mem2_reg[242][19]/P0001 , \wishbone_bd_ram_mem2_reg[242][20]/P0001 , \wishbone_bd_ram_mem2_reg[242][21]/P0001 , \wishbone_bd_ram_mem2_reg[242][22]/P0001 , \wishbone_bd_ram_mem2_reg[242][23]/P0001 , \wishbone_bd_ram_mem2_reg[243][16]/P0001 , \wishbone_bd_ram_mem2_reg[243][17]/P0001 , \wishbone_bd_ram_mem2_reg[243][18]/P0001 , \wishbone_bd_ram_mem2_reg[243][19]/P0001 , \wishbone_bd_ram_mem2_reg[243][20]/P0001 , \wishbone_bd_ram_mem2_reg[243][21]/P0001 , \wishbone_bd_ram_mem2_reg[243][22]/P0001 , \wishbone_bd_ram_mem2_reg[243][23]/P0001 , \wishbone_bd_ram_mem2_reg[244][16]/P0001 , \wishbone_bd_ram_mem2_reg[244][17]/P0001 , \wishbone_bd_ram_mem2_reg[244][18]/P0001 , \wishbone_bd_ram_mem2_reg[244][19]/P0001 , \wishbone_bd_ram_mem2_reg[244][20]/P0001 , \wishbone_bd_ram_mem2_reg[244][21]/P0001 , \wishbone_bd_ram_mem2_reg[244][22]/P0001 , \wishbone_bd_ram_mem2_reg[244][23]/P0001 , \wishbone_bd_ram_mem2_reg[245][16]/P0001 , \wishbone_bd_ram_mem2_reg[245][17]/P0001 , \wishbone_bd_ram_mem2_reg[245][18]/P0001 , \wishbone_bd_ram_mem2_reg[245][19]/P0001 , \wishbone_bd_ram_mem2_reg[245][20]/P0001 , \wishbone_bd_ram_mem2_reg[245][21]/P0001 , \wishbone_bd_ram_mem2_reg[245][22]/P0001 , \wishbone_bd_ram_mem2_reg[245][23]/P0001 , \wishbone_bd_ram_mem2_reg[246][16]/P0001 , \wishbone_bd_ram_mem2_reg[246][17]/P0001 , \wishbone_bd_ram_mem2_reg[246][18]/P0001 , \wishbone_bd_ram_mem2_reg[246][19]/P0001 , \wishbone_bd_ram_mem2_reg[246][20]/P0001 , \wishbone_bd_ram_mem2_reg[246][21]/P0001 , \wishbone_bd_ram_mem2_reg[246][22]/P0001 , \wishbone_bd_ram_mem2_reg[246][23]/P0001 , \wishbone_bd_ram_mem2_reg[247][16]/P0001 , \wishbone_bd_ram_mem2_reg[247][17]/P0001 , \wishbone_bd_ram_mem2_reg[247][18]/P0001 , \wishbone_bd_ram_mem2_reg[247][19]/P0001 , \wishbone_bd_ram_mem2_reg[247][20]/P0001 , \wishbone_bd_ram_mem2_reg[247][21]/P0001 , \wishbone_bd_ram_mem2_reg[247][22]/P0001 , \wishbone_bd_ram_mem2_reg[247][23]/P0001 , \wishbone_bd_ram_mem2_reg[248][16]/P0001 , \wishbone_bd_ram_mem2_reg[248][17]/P0001 , \wishbone_bd_ram_mem2_reg[248][18]/P0001 , \wishbone_bd_ram_mem2_reg[248][19]/P0001 , \wishbone_bd_ram_mem2_reg[248][20]/P0001 , \wishbone_bd_ram_mem2_reg[248][21]/P0001 , \wishbone_bd_ram_mem2_reg[248][22]/P0001 , \wishbone_bd_ram_mem2_reg[248][23]/P0001 , \wishbone_bd_ram_mem2_reg[249][16]/P0001 , \wishbone_bd_ram_mem2_reg[249][17]/P0001 , \wishbone_bd_ram_mem2_reg[249][18]/P0001 , \wishbone_bd_ram_mem2_reg[249][19]/P0001 , \wishbone_bd_ram_mem2_reg[249][20]/P0001 , \wishbone_bd_ram_mem2_reg[249][21]/P0001 , \wishbone_bd_ram_mem2_reg[249][22]/P0001 , \wishbone_bd_ram_mem2_reg[249][23]/P0001 , \wishbone_bd_ram_mem2_reg[24][16]/P0001 , \wishbone_bd_ram_mem2_reg[24][17]/P0001 , \wishbone_bd_ram_mem2_reg[24][18]/P0001 , \wishbone_bd_ram_mem2_reg[24][19]/P0001 , \wishbone_bd_ram_mem2_reg[24][20]/P0001 , \wishbone_bd_ram_mem2_reg[24][21]/P0001 , \wishbone_bd_ram_mem2_reg[24][22]/P0001 , \wishbone_bd_ram_mem2_reg[24][23]/P0001 , \wishbone_bd_ram_mem2_reg[250][16]/P0001 , \wishbone_bd_ram_mem2_reg[250][17]/P0001 , \wishbone_bd_ram_mem2_reg[250][18]/P0001 , \wishbone_bd_ram_mem2_reg[250][19]/P0001 , \wishbone_bd_ram_mem2_reg[250][20]/P0001 , \wishbone_bd_ram_mem2_reg[250][21]/P0001 , \wishbone_bd_ram_mem2_reg[250][22]/P0001 , \wishbone_bd_ram_mem2_reg[250][23]/P0001 , \wishbone_bd_ram_mem2_reg[251][16]/P0001 , \wishbone_bd_ram_mem2_reg[251][17]/P0001 , \wishbone_bd_ram_mem2_reg[251][18]/P0001 , \wishbone_bd_ram_mem2_reg[251][19]/P0001 , \wishbone_bd_ram_mem2_reg[251][20]/P0001 , \wishbone_bd_ram_mem2_reg[251][21]/P0001 , \wishbone_bd_ram_mem2_reg[251][22]/P0001 , \wishbone_bd_ram_mem2_reg[251][23]/P0001 , \wishbone_bd_ram_mem2_reg[252][16]/P0001 , \wishbone_bd_ram_mem2_reg[252][17]/P0001 , \wishbone_bd_ram_mem2_reg[252][18]/P0001 , \wishbone_bd_ram_mem2_reg[252][19]/P0001 , \wishbone_bd_ram_mem2_reg[252][20]/P0001 , \wishbone_bd_ram_mem2_reg[252][21]/P0001 , \wishbone_bd_ram_mem2_reg[252][22]/P0001 , \wishbone_bd_ram_mem2_reg[252][23]/P0001 , \wishbone_bd_ram_mem2_reg[253][16]/P0001 , \wishbone_bd_ram_mem2_reg[253][17]/P0001 , \wishbone_bd_ram_mem2_reg[253][18]/P0001 , \wishbone_bd_ram_mem2_reg[253][19]/P0001 , \wishbone_bd_ram_mem2_reg[253][20]/P0001 , \wishbone_bd_ram_mem2_reg[253][21]/P0001 , \wishbone_bd_ram_mem2_reg[253][22]/P0001 , \wishbone_bd_ram_mem2_reg[253][23]/P0001 , \wishbone_bd_ram_mem2_reg[254][16]/P0001 , \wishbone_bd_ram_mem2_reg[254][17]/P0001 , \wishbone_bd_ram_mem2_reg[254][18]/P0001 , \wishbone_bd_ram_mem2_reg[254][19]/P0001 , \wishbone_bd_ram_mem2_reg[254][20]/P0001 , \wishbone_bd_ram_mem2_reg[254][21]/P0001 , \wishbone_bd_ram_mem2_reg[254][22]/P0001 , \wishbone_bd_ram_mem2_reg[254][23]/P0001 , \wishbone_bd_ram_mem2_reg[255][16]/P0001 , \wishbone_bd_ram_mem2_reg[255][17]/P0001 , \wishbone_bd_ram_mem2_reg[255][18]/P0001 , \wishbone_bd_ram_mem2_reg[255][19]/P0001 , \wishbone_bd_ram_mem2_reg[255][20]/P0001 , \wishbone_bd_ram_mem2_reg[255][21]/P0001 , \wishbone_bd_ram_mem2_reg[255][22]/P0001 , \wishbone_bd_ram_mem2_reg[255][23]/P0001 , \wishbone_bd_ram_mem2_reg[25][16]/P0001 , \wishbone_bd_ram_mem2_reg[25][17]/P0001 , \wishbone_bd_ram_mem2_reg[25][18]/P0001 , \wishbone_bd_ram_mem2_reg[25][19]/P0001 , \wishbone_bd_ram_mem2_reg[25][20]/P0001 , \wishbone_bd_ram_mem2_reg[25][21]/P0001 , \wishbone_bd_ram_mem2_reg[25][22]/P0001 , \wishbone_bd_ram_mem2_reg[25][23]/P0001 , \wishbone_bd_ram_mem2_reg[26][16]/P0001 , \wishbone_bd_ram_mem2_reg[26][17]/P0001 , \wishbone_bd_ram_mem2_reg[26][18]/P0001 , \wishbone_bd_ram_mem2_reg[26][19]/P0001 , \wishbone_bd_ram_mem2_reg[26][20]/P0001 , \wishbone_bd_ram_mem2_reg[26][21]/P0001 , \wishbone_bd_ram_mem2_reg[26][22]/P0001 , \wishbone_bd_ram_mem2_reg[26][23]/P0001 , \wishbone_bd_ram_mem2_reg[27][16]/P0001 , \wishbone_bd_ram_mem2_reg[27][17]/P0001 , \wishbone_bd_ram_mem2_reg[27][18]/P0001 , \wishbone_bd_ram_mem2_reg[27][19]/P0001 , \wishbone_bd_ram_mem2_reg[27][20]/P0001 , \wishbone_bd_ram_mem2_reg[27][21]/P0001 , \wishbone_bd_ram_mem2_reg[27][22]/P0001 , \wishbone_bd_ram_mem2_reg[27][23]/P0001 , \wishbone_bd_ram_mem2_reg[28][16]/P0001 , \wishbone_bd_ram_mem2_reg[28][17]/P0001 , \wishbone_bd_ram_mem2_reg[28][18]/P0001 , \wishbone_bd_ram_mem2_reg[28][19]/P0001 , \wishbone_bd_ram_mem2_reg[28][20]/P0001 , \wishbone_bd_ram_mem2_reg[28][21]/P0001 , \wishbone_bd_ram_mem2_reg[28][22]/P0001 , \wishbone_bd_ram_mem2_reg[28][23]/P0001 , \wishbone_bd_ram_mem2_reg[29][16]/P0001 , \wishbone_bd_ram_mem2_reg[29][17]/P0001 , \wishbone_bd_ram_mem2_reg[29][18]/P0001 , \wishbone_bd_ram_mem2_reg[29][19]/P0001 , \wishbone_bd_ram_mem2_reg[29][20]/P0001 , \wishbone_bd_ram_mem2_reg[29][21]/P0001 , \wishbone_bd_ram_mem2_reg[29][22]/P0001 , \wishbone_bd_ram_mem2_reg[29][23]/P0001 , \wishbone_bd_ram_mem2_reg[2][16]/P0001 , \wishbone_bd_ram_mem2_reg[2][17]/P0001 , \wishbone_bd_ram_mem2_reg[2][18]/P0001 , \wishbone_bd_ram_mem2_reg[2][19]/P0001 , \wishbone_bd_ram_mem2_reg[2][20]/P0001 , \wishbone_bd_ram_mem2_reg[2][21]/P0001 , \wishbone_bd_ram_mem2_reg[2][22]/P0001 , \wishbone_bd_ram_mem2_reg[2][23]/P0001 , \wishbone_bd_ram_mem2_reg[30][16]/P0001 , \wishbone_bd_ram_mem2_reg[30][17]/P0001 , \wishbone_bd_ram_mem2_reg[30][18]/P0001 , \wishbone_bd_ram_mem2_reg[30][19]/P0001 , \wishbone_bd_ram_mem2_reg[30][20]/P0001 , \wishbone_bd_ram_mem2_reg[30][21]/P0001 , \wishbone_bd_ram_mem2_reg[30][22]/P0001 , \wishbone_bd_ram_mem2_reg[30][23]/P0001 , \wishbone_bd_ram_mem2_reg[31][16]/P0001 , \wishbone_bd_ram_mem2_reg[31][17]/P0001 , \wishbone_bd_ram_mem2_reg[31][18]/P0001 , \wishbone_bd_ram_mem2_reg[31][19]/P0001 , \wishbone_bd_ram_mem2_reg[31][20]/P0001 , \wishbone_bd_ram_mem2_reg[31][21]/P0001 , \wishbone_bd_ram_mem2_reg[31][22]/P0001 , \wishbone_bd_ram_mem2_reg[31][23]/P0001 , \wishbone_bd_ram_mem2_reg[32][16]/P0001 , \wishbone_bd_ram_mem2_reg[32][17]/P0001 , \wishbone_bd_ram_mem2_reg[32][18]/P0001 , \wishbone_bd_ram_mem2_reg[32][19]/P0001 , \wishbone_bd_ram_mem2_reg[32][20]/P0001 , \wishbone_bd_ram_mem2_reg[32][21]/P0001 , \wishbone_bd_ram_mem2_reg[32][22]/P0001 , \wishbone_bd_ram_mem2_reg[32][23]/P0001 , \wishbone_bd_ram_mem2_reg[33][16]/P0001 , \wishbone_bd_ram_mem2_reg[33][17]/P0001 , \wishbone_bd_ram_mem2_reg[33][18]/P0001 , \wishbone_bd_ram_mem2_reg[33][19]/P0001 , \wishbone_bd_ram_mem2_reg[33][20]/P0001 , \wishbone_bd_ram_mem2_reg[33][21]/P0001 , \wishbone_bd_ram_mem2_reg[33][22]/P0001 , \wishbone_bd_ram_mem2_reg[33][23]/P0001 , \wishbone_bd_ram_mem2_reg[34][16]/P0001 , \wishbone_bd_ram_mem2_reg[34][17]/P0001 , \wishbone_bd_ram_mem2_reg[34][18]/P0001 , \wishbone_bd_ram_mem2_reg[34][19]/P0001 , \wishbone_bd_ram_mem2_reg[34][20]/P0001 , \wishbone_bd_ram_mem2_reg[34][21]/P0001 , \wishbone_bd_ram_mem2_reg[34][22]/P0001 , \wishbone_bd_ram_mem2_reg[34][23]/P0001 , \wishbone_bd_ram_mem2_reg[35][16]/P0001 , \wishbone_bd_ram_mem2_reg[35][17]/P0001 , \wishbone_bd_ram_mem2_reg[35][18]/P0001 , \wishbone_bd_ram_mem2_reg[35][19]/P0001 , \wishbone_bd_ram_mem2_reg[35][20]/P0001 , \wishbone_bd_ram_mem2_reg[35][21]/P0001 , \wishbone_bd_ram_mem2_reg[35][22]/P0001 , \wishbone_bd_ram_mem2_reg[35][23]/P0001 , \wishbone_bd_ram_mem2_reg[36][16]/P0001 , \wishbone_bd_ram_mem2_reg[36][17]/P0001 , \wishbone_bd_ram_mem2_reg[36][18]/P0001 , \wishbone_bd_ram_mem2_reg[36][19]/P0001 , \wishbone_bd_ram_mem2_reg[36][20]/P0001 , \wishbone_bd_ram_mem2_reg[36][21]/P0001 , \wishbone_bd_ram_mem2_reg[36][22]/P0001 , \wishbone_bd_ram_mem2_reg[36][23]/P0001 , \wishbone_bd_ram_mem2_reg[37][16]/P0001 , \wishbone_bd_ram_mem2_reg[37][17]/P0001 , \wishbone_bd_ram_mem2_reg[37][18]/P0001 , \wishbone_bd_ram_mem2_reg[37][19]/P0001 , \wishbone_bd_ram_mem2_reg[37][20]/P0001 , \wishbone_bd_ram_mem2_reg[37][21]/P0001 , \wishbone_bd_ram_mem2_reg[37][22]/P0001 , \wishbone_bd_ram_mem2_reg[37][23]/P0001 , \wishbone_bd_ram_mem2_reg[38][16]/P0001 , \wishbone_bd_ram_mem2_reg[38][17]/P0001 , \wishbone_bd_ram_mem2_reg[38][18]/P0001 , \wishbone_bd_ram_mem2_reg[38][19]/P0001 , \wishbone_bd_ram_mem2_reg[38][20]/P0001 , \wishbone_bd_ram_mem2_reg[38][21]/P0001 , \wishbone_bd_ram_mem2_reg[38][22]/P0001 , \wishbone_bd_ram_mem2_reg[38][23]/P0001 , \wishbone_bd_ram_mem2_reg[39][16]/P0001 , \wishbone_bd_ram_mem2_reg[39][17]/P0001 , \wishbone_bd_ram_mem2_reg[39][18]/P0001 , \wishbone_bd_ram_mem2_reg[39][19]/P0001 , \wishbone_bd_ram_mem2_reg[39][20]/P0001 , \wishbone_bd_ram_mem2_reg[39][21]/P0001 , \wishbone_bd_ram_mem2_reg[39][22]/P0001 , \wishbone_bd_ram_mem2_reg[39][23]/P0001 , \wishbone_bd_ram_mem2_reg[3][16]/P0001 , \wishbone_bd_ram_mem2_reg[3][17]/P0001 , \wishbone_bd_ram_mem2_reg[3][18]/P0001 , \wishbone_bd_ram_mem2_reg[3][19]/P0001 , \wishbone_bd_ram_mem2_reg[3][20]/P0001 , \wishbone_bd_ram_mem2_reg[3][21]/P0001 , \wishbone_bd_ram_mem2_reg[3][22]/P0001 , \wishbone_bd_ram_mem2_reg[3][23]/P0001 , \wishbone_bd_ram_mem2_reg[40][16]/P0001 , \wishbone_bd_ram_mem2_reg[40][17]/P0001 , \wishbone_bd_ram_mem2_reg[40][18]/P0001 , \wishbone_bd_ram_mem2_reg[40][19]/P0001 , \wishbone_bd_ram_mem2_reg[40][20]/P0001 , \wishbone_bd_ram_mem2_reg[40][21]/P0001 , \wishbone_bd_ram_mem2_reg[40][22]/P0001 , \wishbone_bd_ram_mem2_reg[40][23]/P0001 , \wishbone_bd_ram_mem2_reg[41][16]/P0001 , \wishbone_bd_ram_mem2_reg[41][17]/P0001 , \wishbone_bd_ram_mem2_reg[41][18]/P0001 , \wishbone_bd_ram_mem2_reg[41][19]/P0001 , \wishbone_bd_ram_mem2_reg[41][20]/P0001 , \wishbone_bd_ram_mem2_reg[41][21]/P0001 , \wishbone_bd_ram_mem2_reg[41][22]/P0001 , \wishbone_bd_ram_mem2_reg[41][23]/P0001 , \wishbone_bd_ram_mem2_reg[42][16]/P0001 , \wishbone_bd_ram_mem2_reg[42][17]/P0001 , \wishbone_bd_ram_mem2_reg[42][18]/P0001 , \wishbone_bd_ram_mem2_reg[42][19]/P0001 , \wishbone_bd_ram_mem2_reg[42][20]/P0001 , \wishbone_bd_ram_mem2_reg[42][21]/P0001 , \wishbone_bd_ram_mem2_reg[42][22]/P0001 , \wishbone_bd_ram_mem2_reg[42][23]/P0001 , \wishbone_bd_ram_mem2_reg[43][16]/P0001 , \wishbone_bd_ram_mem2_reg[43][17]/P0001 , \wishbone_bd_ram_mem2_reg[43][18]/P0001 , \wishbone_bd_ram_mem2_reg[43][19]/P0001 , \wishbone_bd_ram_mem2_reg[43][20]/P0001 , \wishbone_bd_ram_mem2_reg[43][21]/P0001 , \wishbone_bd_ram_mem2_reg[43][22]/P0001 , \wishbone_bd_ram_mem2_reg[43][23]/P0001 , \wishbone_bd_ram_mem2_reg[44][16]/P0001 , \wishbone_bd_ram_mem2_reg[44][17]/P0001 , \wishbone_bd_ram_mem2_reg[44][18]/P0001 , \wishbone_bd_ram_mem2_reg[44][19]/P0001 , \wishbone_bd_ram_mem2_reg[44][20]/P0001 , \wishbone_bd_ram_mem2_reg[44][21]/P0001 , \wishbone_bd_ram_mem2_reg[44][22]/P0001 , \wishbone_bd_ram_mem2_reg[44][23]/P0001 , \wishbone_bd_ram_mem2_reg[45][16]/P0001 , \wishbone_bd_ram_mem2_reg[45][17]/P0001 , \wishbone_bd_ram_mem2_reg[45][18]/P0001 , \wishbone_bd_ram_mem2_reg[45][19]/P0001 , \wishbone_bd_ram_mem2_reg[45][20]/P0001 , \wishbone_bd_ram_mem2_reg[45][21]/P0001 , \wishbone_bd_ram_mem2_reg[45][22]/P0001 , \wishbone_bd_ram_mem2_reg[45][23]/P0001 , \wishbone_bd_ram_mem2_reg[46][16]/P0001 , \wishbone_bd_ram_mem2_reg[46][17]/P0001 , \wishbone_bd_ram_mem2_reg[46][18]/P0001 , \wishbone_bd_ram_mem2_reg[46][19]/P0001 , \wishbone_bd_ram_mem2_reg[46][20]/P0001 , \wishbone_bd_ram_mem2_reg[46][21]/P0001 , \wishbone_bd_ram_mem2_reg[46][22]/P0001 , \wishbone_bd_ram_mem2_reg[46][23]/P0001 , \wishbone_bd_ram_mem2_reg[47][16]/P0001 , \wishbone_bd_ram_mem2_reg[47][17]/P0001 , \wishbone_bd_ram_mem2_reg[47][18]/P0001 , \wishbone_bd_ram_mem2_reg[47][19]/P0001 , \wishbone_bd_ram_mem2_reg[47][20]/P0001 , \wishbone_bd_ram_mem2_reg[47][21]/P0001 , \wishbone_bd_ram_mem2_reg[47][22]/P0001 , \wishbone_bd_ram_mem2_reg[47][23]/P0001 , \wishbone_bd_ram_mem2_reg[48][16]/P0001 , \wishbone_bd_ram_mem2_reg[48][17]/P0001 , \wishbone_bd_ram_mem2_reg[48][18]/P0001 , \wishbone_bd_ram_mem2_reg[48][19]/P0001 , \wishbone_bd_ram_mem2_reg[48][20]/P0001 , \wishbone_bd_ram_mem2_reg[48][21]/P0001 , \wishbone_bd_ram_mem2_reg[48][22]/P0001 , \wishbone_bd_ram_mem2_reg[48][23]/P0001 , \wishbone_bd_ram_mem2_reg[49][16]/P0001 , \wishbone_bd_ram_mem2_reg[49][17]/P0001 , \wishbone_bd_ram_mem2_reg[49][18]/P0001 , \wishbone_bd_ram_mem2_reg[49][19]/P0001 , \wishbone_bd_ram_mem2_reg[49][20]/P0001 , \wishbone_bd_ram_mem2_reg[49][21]/P0001 , \wishbone_bd_ram_mem2_reg[49][22]/P0001 , \wishbone_bd_ram_mem2_reg[49][23]/P0001 , \wishbone_bd_ram_mem2_reg[4][16]/P0001 , \wishbone_bd_ram_mem2_reg[4][17]/P0001 , \wishbone_bd_ram_mem2_reg[4][18]/P0001 , \wishbone_bd_ram_mem2_reg[4][19]/P0001 , \wishbone_bd_ram_mem2_reg[4][20]/P0001 , \wishbone_bd_ram_mem2_reg[4][21]/P0001 , \wishbone_bd_ram_mem2_reg[4][22]/P0001 , \wishbone_bd_ram_mem2_reg[4][23]/P0001 , \wishbone_bd_ram_mem2_reg[50][16]/P0001 , \wishbone_bd_ram_mem2_reg[50][17]/P0001 , \wishbone_bd_ram_mem2_reg[50][18]/P0001 , \wishbone_bd_ram_mem2_reg[50][19]/P0001 , \wishbone_bd_ram_mem2_reg[50][20]/P0001 , \wishbone_bd_ram_mem2_reg[50][21]/P0001 , \wishbone_bd_ram_mem2_reg[50][22]/P0001 , \wishbone_bd_ram_mem2_reg[50][23]/P0001 , \wishbone_bd_ram_mem2_reg[51][16]/P0001 , \wishbone_bd_ram_mem2_reg[51][17]/P0001 , \wishbone_bd_ram_mem2_reg[51][18]/P0001 , \wishbone_bd_ram_mem2_reg[51][19]/P0001 , \wishbone_bd_ram_mem2_reg[51][20]/P0001 , \wishbone_bd_ram_mem2_reg[51][21]/P0001 , \wishbone_bd_ram_mem2_reg[51][22]/P0001 , \wishbone_bd_ram_mem2_reg[51][23]/P0001 , \wishbone_bd_ram_mem2_reg[52][16]/P0001 , \wishbone_bd_ram_mem2_reg[52][17]/P0001 , \wishbone_bd_ram_mem2_reg[52][18]/P0001 , \wishbone_bd_ram_mem2_reg[52][19]/P0001 , \wishbone_bd_ram_mem2_reg[52][20]/P0001 , \wishbone_bd_ram_mem2_reg[52][21]/P0001 , \wishbone_bd_ram_mem2_reg[52][22]/P0001 , \wishbone_bd_ram_mem2_reg[52][23]/P0001 , \wishbone_bd_ram_mem2_reg[53][16]/P0001 , \wishbone_bd_ram_mem2_reg[53][17]/P0001 , \wishbone_bd_ram_mem2_reg[53][18]/P0001 , \wishbone_bd_ram_mem2_reg[53][19]/P0001 , \wishbone_bd_ram_mem2_reg[53][20]/P0001 , \wishbone_bd_ram_mem2_reg[53][21]/P0001 , \wishbone_bd_ram_mem2_reg[53][22]/P0001 , \wishbone_bd_ram_mem2_reg[53][23]/P0001 , \wishbone_bd_ram_mem2_reg[54][16]/P0001 , \wishbone_bd_ram_mem2_reg[54][17]/P0001 , \wishbone_bd_ram_mem2_reg[54][18]/P0001 , \wishbone_bd_ram_mem2_reg[54][19]/P0001 , \wishbone_bd_ram_mem2_reg[54][20]/P0001 , \wishbone_bd_ram_mem2_reg[54][21]/P0001 , \wishbone_bd_ram_mem2_reg[54][22]/P0001 , \wishbone_bd_ram_mem2_reg[54][23]/P0001 , \wishbone_bd_ram_mem2_reg[55][16]/P0001 , \wishbone_bd_ram_mem2_reg[55][17]/P0001 , \wishbone_bd_ram_mem2_reg[55][18]/P0001 , \wishbone_bd_ram_mem2_reg[55][19]/P0001 , \wishbone_bd_ram_mem2_reg[55][20]/P0001 , \wishbone_bd_ram_mem2_reg[55][21]/P0001 , \wishbone_bd_ram_mem2_reg[55][22]/P0001 , \wishbone_bd_ram_mem2_reg[55][23]/P0001 , \wishbone_bd_ram_mem2_reg[56][16]/P0001 , \wishbone_bd_ram_mem2_reg[56][17]/P0001 , \wishbone_bd_ram_mem2_reg[56][18]/P0001 , \wishbone_bd_ram_mem2_reg[56][19]/P0001 , \wishbone_bd_ram_mem2_reg[56][20]/P0001 , \wishbone_bd_ram_mem2_reg[56][21]/P0001 , \wishbone_bd_ram_mem2_reg[56][22]/P0001 , \wishbone_bd_ram_mem2_reg[56][23]/P0001 , \wishbone_bd_ram_mem2_reg[57][16]/P0001 , \wishbone_bd_ram_mem2_reg[57][17]/P0001 , \wishbone_bd_ram_mem2_reg[57][18]/P0001 , \wishbone_bd_ram_mem2_reg[57][19]/P0001 , \wishbone_bd_ram_mem2_reg[57][20]/P0001 , \wishbone_bd_ram_mem2_reg[57][21]/P0001 , \wishbone_bd_ram_mem2_reg[57][22]/P0001 , \wishbone_bd_ram_mem2_reg[57][23]/P0001 , \wishbone_bd_ram_mem2_reg[58][16]/P0001 , \wishbone_bd_ram_mem2_reg[58][17]/P0001 , \wishbone_bd_ram_mem2_reg[58][18]/P0001 , \wishbone_bd_ram_mem2_reg[58][19]/P0001 , \wishbone_bd_ram_mem2_reg[58][20]/P0001 , \wishbone_bd_ram_mem2_reg[58][21]/P0001 , \wishbone_bd_ram_mem2_reg[58][22]/P0001 , \wishbone_bd_ram_mem2_reg[58][23]/P0001 , \wishbone_bd_ram_mem2_reg[59][16]/P0001 , \wishbone_bd_ram_mem2_reg[59][17]/P0001 , \wishbone_bd_ram_mem2_reg[59][18]/P0001 , \wishbone_bd_ram_mem2_reg[59][19]/P0001 , \wishbone_bd_ram_mem2_reg[59][20]/P0001 , \wishbone_bd_ram_mem2_reg[59][21]/P0001 , \wishbone_bd_ram_mem2_reg[59][22]/P0001 , \wishbone_bd_ram_mem2_reg[59][23]/P0001 , \wishbone_bd_ram_mem2_reg[5][16]/P0001 , \wishbone_bd_ram_mem2_reg[5][17]/P0001 , \wishbone_bd_ram_mem2_reg[5][18]/P0001 , \wishbone_bd_ram_mem2_reg[5][19]/P0001 , \wishbone_bd_ram_mem2_reg[5][20]/P0001 , \wishbone_bd_ram_mem2_reg[5][21]/P0001 , \wishbone_bd_ram_mem2_reg[5][22]/P0001 , \wishbone_bd_ram_mem2_reg[5][23]/P0001 , \wishbone_bd_ram_mem2_reg[60][16]/P0001 , \wishbone_bd_ram_mem2_reg[60][17]/P0001 , \wishbone_bd_ram_mem2_reg[60][18]/P0001 , \wishbone_bd_ram_mem2_reg[60][19]/P0001 , \wishbone_bd_ram_mem2_reg[60][20]/P0001 , \wishbone_bd_ram_mem2_reg[60][21]/P0001 , \wishbone_bd_ram_mem2_reg[60][22]/P0001 , \wishbone_bd_ram_mem2_reg[60][23]/P0001 , \wishbone_bd_ram_mem2_reg[61][16]/P0001 , \wishbone_bd_ram_mem2_reg[61][17]/P0001 , \wishbone_bd_ram_mem2_reg[61][18]/P0001 , \wishbone_bd_ram_mem2_reg[61][19]/P0001 , \wishbone_bd_ram_mem2_reg[61][20]/P0001 , \wishbone_bd_ram_mem2_reg[61][21]/P0001 , \wishbone_bd_ram_mem2_reg[61][22]/P0001 , \wishbone_bd_ram_mem2_reg[61][23]/P0001 , \wishbone_bd_ram_mem2_reg[62][16]/P0001 , \wishbone_bd_ram_mem2_reg[62][17]/P0001 , \wishbone_bd_ram_mem2_reg[62][18]/P0001 , \wishbone_bd_ram_mem2_reg[62][19]/P0001 , \wishbone_bd_ram_mem2_reg[62][20]/P0001 , \wishbone_bd_ram_mem2_reg[62][21]/P0001 , \wishbone_bd_ram_mem2_reg[62][22]/P0001 , \wishbone_bd_ram_mem2_reg[62][23]/P0001 , \wishbone_bd_ram_mem2_reg[63][16]/P0001 , \wishbone_bd_ram_mem2_reg[63][17]/P0001 , \wishbone_bd_ram_mem2_reg[63][18]/P0001 , \wishbone_bd_ram_mem2_reg[63][19]/P0001 , \wishbone_bd_ram_mem2_reg[63][20]/P0001 , \wishbone_bd_ram_mem2_reg[63][21]/P0001 , \wishbone_bd_ram_mem2_reg[63][22]/P0001 , \wishbone_bd_ram_mem2_reg[63][23]/P0001 , \wishbone_bd_ram_mem2_reg[64][16]/P0001 , \wishbone_bd_ram_mem2_reg[64][17]/P0001 , \wishbone_bd_ram_mem2_reg[64][18]/P0001 , \wishbone_bd_ram_mem2_reg[64][19]/P0001 , \wishbone_bd_ram_mem2_reg[64][20]/P0001 , \wishbone_bd_ram_mem2_reg[64][21]/P0001 , \wishbone_bd_ram_mem2_reg[64][22]/P0001 , \wishbone_bd_ram_mem2_reg[64][23]/P0001 , \wishbone_bd_ram_mem2_reg[65][16]/P0001 , \wishbone_bd_ram_mem2_reg[65][17]/P0001 , \wishbone_bd_ram_mem2_reg[65][18]/P0001 , \wishbone_bd_ram_mem2_reg[65][19]/P0001 , \wishbone_bd_ram_mem2_reg[65][20]/P0001 , \wishbone_bd_ram_mem2_reg[65][21]/P0001 , \wishbone_bd_ram_mem2_reg[65][22]/P0001 , \wishbone_bd_ram_mem2_reg[65][23]/P0001 , \wishbone_bd_ram_mem2_reg[66][16]/P0001 , \wishbone_bd_ram_mem2_reg[66][17]/P0001 , \wishbone_bd_ram_mem2_reg[66][18]/P0001 , \wishbone_bd_ram_mem2_reg[66][19]/P0001 , \wishbone_bd_ram_mem2_reg[66][20]/P0001 , \wishbone_bd_ram_mem2_reg[66][21]/P0001 , \wishbone_bd_ram_mem2_reg[66][22]/P0001 , \wishbone_bd_ram_mem2_reg[66][23]/P0001 , \wishbone_bd_ram_mem2_reg[67][16]/P0001 , \wishbone_bd_ram_mem2_reg[67][17]/P0001 , \wishbone_bd_ram_mem2_reg[67][18]/P0001 , \wishbone_bd_ram_mem2_reg[67][19]/P0001 , \wishbone_bd_ram_mem2_reg[67][20]/P0001 , \wishbone_bd_ram_mem2_reg[67][21]/P0001 , \wishbone_bd_ram_mem2_reg[67][22]/P0001 , \wishbone_bd_ram_mem2_reg[67][23]/P0001 , \wishbone_bd_ram_mem2_reg[68][16]/P0001 , \wishbone_bd_ram_mem2_reg[68][17]/P0001 , \wishbone_bd_ram_mem2_reg[68][18]/P0001 , \wishbone_bd_ram_mem2_reg[68][19]/P0001 , \wishbone_bd_ram_mem2_reg[68][20]/P0001 , \wishbone_bd_ram_mem2_reg[68][21]/P0001 , \wishbone_bd_ram_mem2_reg[68][22]/P0001 , \wishbone_bd_ram_mem2_reg[68][23]/P0001 , \wishbone_bd_ram_mem2_reg[69][16]/P0001 , \wishbone_bd_ram_mem2_reg[69][17]/P0001 , \wishbone_bd_ram_mem2_reg[69][18]/P0001 , \wishbone_bd_ram_mem2_reg[69][19]/P0001 , \wishbone_bd_ram_mem2_reg[69][20]/P0001 , \wishbone_bd_ram_mem2_reg[69][21]/P0001 , \wishbone_bd_ram_mem2_reg[69][22]/P0001 , \wishbone_bd_ram_mem2_reg[69][23]/P0001 , \wishbone_bd_ram_mem2_reg[6][16]/P0001 , \wishbone_bd_ram_mem2_reg[6][17]/P0001 , \wishbone_bd_ram_mem2_reg[6][18]/P0001 , \wishbone_bd_ram_mem2_reg[6][19]/P0001 , \wishbone_bd_ram_mem2_reg[6][20]/P0001 , \wishbone_bd_ram_mem2_reg[6][21]/P0001 , \wishbone_bd_ram_mem2_reg[6][22]/P0001 , \wishbone_bd_ram_mem2_reg[6][23]/P0001 , \wishbone_bd_ram_mem2_reg[70][16]/P0001 , \wishbone_bd_ram_mem2_reg[70][17]/P0001 , \wishbone_bd_ram_mem2_reg[70][18]/P0001 , \wishbone_bd_ram_mem2_reg[70][19]/P0001 , \wishbone_bd_ram_mem2_reg[70][20]/P0001 , \wishbone_bd_ram_mem2_reg[70][21]/P0001 , \wishbone_bd_ram_mem2_reg[70][22]/P0001 , \wishbone_bd_ram_mem2_reg[70][23]/P0001 , \wishbone_bd_ram_mem2_reg[71][16]/P0001 , \wishbone_bd_ram_mem2_reg[71][17]/P0001 , \wishbone_bd_ram_mem2_reg[71][18]/P0001 , \wishbone_bd_ram_mem2_reg[71][19]/P0001 , \wishbone_bd_ram_mem2_reg[71][20]/P0001 , \wishbone_bd_ram_mem2_reg[71][21]/P0001 , \wishbone_bd_ram_mem2_reg[71][22]/P0001 , \wishbone_bd_ram_mem2_reg[71][23]/P0001 , \wishbone_bd_ram_mem2_reg[72][16]/P0001 , \wishbone_bd_ram_mem2_reg[72][17]/P0001 , \wishbone_bd_ram_mem2_reg[72][18]/P0001 , \wishbone_bd_ram_mem2_reg[72][19]/P0001 , \wishbone_bd_ram_mem2_reg[72][20]/P0001 , \wishbone_bd_ram_mem2_reg[72][21]/P0001 , \wishbone_bd_ram_mem2_reg[72][22]/P0001 , \wishbone_bd_ram_mem2_reg[72][23]/P0001 , \wishbone_bd_ram_mem2_reg[73][16]/P0001 , \wishbone_bd_ram_mem2_reg[73][17]/P0001 , \wishbone_bd_ram_mem2_reg[73][18]/P0001 , \wishbone_bd_ram_mem2_reg[73][19]/P0001 , \wishbone_bd_ram_mem2_reg[73][20]/P0001 , \wishbone_bd_ram_mem2_reg[73][21]/P0001 , \wishbone_bd_ram_mem2_reg[73][22]/P0001 , \wishbone_bd_ram_mem2_reg[73][23]/P0001 , \wishbone_bd_ram_mem2_reg[74][16]/P0001 , \wishbone_bd_ram_mem2_reg[74][17]/P0001 , \wishbone_bd_ram_mem2_reg[74][18]/P0001 , \wishbone_bd_ram_mem2_reg[74][19]/P0001 , \wishbone_bd_ram_mem2_reg[74][20]/P0001 , \wishbone_bd_ram_mem2_reg[74][21]/P0001 , \wishbone_bd_ram_mem2_reg[74][22]/P0001 , \wishbone_bd_ram_mem2_reg[74][23]/P0001 , \wishbone_bd_ram_mem2_reg[75][16]/P0001 , \wishbone_bd_ram_mem2_reg[75][17]/P0001 , \wishbone_bd_ram_mem2_reg[75][18]/P0001 , \wishbone_bd_ram_mem2_reg[75][19]/P0001 , \wishbone_bd_ram_mem2_reg[75][20]/P0001 , \wishbone_bd_ram_mem2_reg[75][21]/P0001 , \wishbone_bd_ram_mem2_reg[75][22]/P0001 , \wishbone_bd_ram_mem2_reg[75][23]/P0001 , \wishbone_bd_ram_mem2_reg[76][16]/P0001 , \wishbone_bd_ram_mem2_reg[76][17]/P0001 , \wishbone_bd_ram_mem2_reg[76][18]/P0001 , \wishbone_bd_ram_mem2_reg[76][19]/P0001 , \wishbone_bd_ram_mem2_reg[76][20]/P0001 , \wishbone_bd_ram_mem2_reg[76][21]/P0001 , \wishbone_bd_ram_mem2_reg[76][22]/P0001 , \wishbone_bd_ram_mem2_reg[76][23]/P0001 , \wishbone_bd_ram_mem2_reg[77][16]/P0001 , \wishbone_bd_ram_mem2_reg[77][17]/P0001 , \wishbone_bd_ram_mem2_reg[77][18]/P0001 , \wishbone_bd_ram_mem2_reg[77][19]/P0001 , \wishbone_bd_ram_mem2_reg[77][20]/P0001 , \wishbone_bd_ram_mem2_reg[77][21]/P0001 , \wishbone_bd_ram_mem2_reg[77][22]/P0001 , \wishbone_bd_ram_mem2_reg[77][23]/P0001 , \wishbone_bd_ram_mem2_reg[78][16]/P0001 , \wishbone_bd_ram_mem2_reg[78][17]/P0001 , \wishbone_bd_ram_mem2_reg[78][18]/P0001 , \wishbone_bd_ram_mem2_reg[78][19]/P0001 , \wishbone_bd_ram_mem2_reg[78][20]/P0001 , \wishbone_bd_ram_mem2_reg[78][21]/P0001 , \wishbone_bd_ram_mem2_reg[78][22]/P0001 , \wishbone_bd_ram_mem2_reg[78][23]/P0001 , \wishbone_bd_ram_mem2_reg[79][16]/P0001 , \wishbone_bd_ram_mem2_reg[79][17]/P0001 , \wishbone_bd_ram_mem2_reg[79][18]/P0001 , \wishbone_bd_ram_mem2_reg[79][19]/P0001 , \wishbone_bd_ram_mem2_reg[79][20]/P0001 , \wishbone_bd_ram_mem2_reg[79][21]/P0001 , \wishbone_bd_ram_mem2_reg[79][22]/P0001 , \wishbone_bd_ram_mem2_reg[79][23]/P0001 , \wishbone_bd_ram_mem2_reg[7][16]/P0001 , \wishbone_bd_ram_mem2_reg[7][17]/P0001 , \wishbone_bd_ram_mem2_reg[7][18]/P0001 , \wishbone_bd_ram_mem2_reg[7][19]/P0001 , \wishbone_bd_ram_mem2_reg[7][20]/P0001 , \wishbone_bd_ram_mem2_reg[7][21]/P0001 , \wishbone_bd_ram_mem2_reg[7][22]/P0001 , \wishbone_bd_ram_mem2_reg[7][23]/P0001 , \wishbone_bd_ram_mem2_reg[80][16]/P0001 , \wishbone_bd_ram_mem2_reg[80][17]/P0001 , \wishbone_bd_ram_mem2_reg[80][18]/P0001 , \wishbone_bd_ram_mem2_reg[80][19]/P0001 , \wishbone_bd_ram_mem2_reg[80][20]/P0001 , \wishbone_bd_ram_mem2_reg[80][21]/P0001 , \wishbone_bd_ram_mem2_reg[80][22]/P0001 , \wishbone_bd_ram_mem2_reg[80][23]/P0001 , \wishbone_bd_ram_mem2_reg[81][16]/P0001 , \wishbone_bd_ram_mem2_reg[81][17]/P0001 , \wishbone_bd_ram_mem2_reg[81][18]/P0001 , \wishbone_bd_ram_mem2_reg[81][19]/P0001 , \wishbone_bd_ram_mem2_reg[81][20]/P0001 , \wishbone_bd_ram_mem2_reg[81][21]/P0001 , \wishbone_bd_ram_mem2_reg[81][22]/P0001 , \wishbone_bd_ram_mem2_reg[81][23]/P0001 , \wishbone_bd_ram_mem2_reg[82][16]/P0001 , \wishbone_bd_ram_mem2_reg[82][17]/P0001 , \wishbone_bd_ram_mem2_reg[82][18]/P0001 , \wishbone_bd_ram_mem2_reg[82][19]/P0001 , \wishbone_bd_ram_mem2_reg[82][20]/P0001 , \wishbone_bd_ram_mem2_reg[82][21]/P0001 , \wishbone_bd_ram_mem2_reg[82][22]/P0001 , \wishbone_bd_ram_mem2_reg[82][23]/P0001 , \wishbone_bd_ram_mem2_reg[83][16]/P0001 , \wishbone_bd_ram_mem2_reg[83][17]/P0001 , \wishbone_bd_ram_mem2_reg[83][18]/P0001 , \wishbone_bd_ram_mem2_reg[83][19]/P0001 , \wishbone_bd_ram_mem2_reg[83][20]/P0001 , \wishbone_bd_ram_mem2_reg[83][21]/P0001 , \wishbone_bd_ram_mem2_reg[83][22]/P0001 , \wishbone_bd_ram_mem2_reg[83][23]/P0001 , \wishbone_bd_ram_mem2_reg[84][16]/P0001 , \wishbone_bd_ram_mem2_reg[84][17]/P0001 , \wishbone_bd_ram_mem2_reg[84][18]/P0001 , \wishbone_bd_ram_mem2_reg[84][19]/P0001 , \wishbone_bd_ram_mem2_reg[84][20]/P0001 , \wishbone_bd_ram_mem2_reg[84][21]/P0001 , \wishbone_bd_ram_mem2_reg[84][22]/P0001 , \wishbone_bd_ram_mem2_reg[84][23]/P0001 , \wishbone_bd_ram_mem2_reg[85][16]/P0001 , \wishbone_bd_ram_mem2_reg[85][17]/P0001 , \wishbone_bd_ram_mem2_reg[85][18]/P0001 , \wishbone_bd_ram_mem2_reg[85][19]/P0001 , \wishbone_bd_ram_mem2_reg[85][20]/P0001 , \wishbone_bd_ram_mem2_reg[85][21]/P0001 , \wishbone_bd_ram_mem2_reg[85][22]/P0001 , \wishbone_bd_ram_mem2_reg[85][23]/P0001 , \wishbone_bd_ram_mem2_reg[86][16]/P0001 , \wishbone_bd_ram_mem2_reg[86][17]/P0001 , \wishbone_bd_ram_mem2_reg[86][18]/P0001 , \wishbone_bd_ram_mem2_reg[86][19]/P0001 , \wishbone_bd_ram_mem2_reg[86][20]/P0001 , \wishbone_bd_ram_mem2_reg[86][21]/P0001 , \wishbone_bd_ram_mem2_reg[86][22]/P0001 , \wishbone_bd_ram_mem2_reg[86][23]/P0001 , \wishbone_bd_ram_mem2_reg[87][16]/P0001 , \wishbone_bd_ram_mem2_reg[87][17]/P0001 , \wishbone_bd_ram_mem2_reg[87][18]/P0001 , \wishbone_bd_ram_mem2_reg[87][19]/P0001 , \wishbone_bd_ram_mem2_reg[87][20]/P0001 , \wishbone_bd_ram_mem2_reg[87][21]/P0001 , \wishbone_bd_ram_mem2_reg[87][22]/P0001 , \wishbone_bd_ram_mem2_reg[87][23]/P0001 , \wishbone_bd_ram_mem2_reg[88][16]/P0001 , \wishbone_bd_ram_mem2_reg[88][17]/P0001 , \wishbone_bd_ram_mem2_reg[88][18]/P0001 , \wishbone_bd_ram_mem2_reg[88][19]/P0001 , \wishbone_bd_ram_mem2_reg[88][20]/P0001 , \wishbone_bd_ram_mem2_reg[88][21]/P0001 , \wishbone_bd_ram_mem2_reg[88][22]/P0001 , \wishbone_bd_ram_mem2_reg[88][23]/P0001 , \wishbone_bd_ram_mem2_reg[89][16]/P0001 , \wishbone_bd_ram_mem2_reg[89][17]/P0001 , \wishbone_bd_ram_mem2_reg[89][18]/P0001 , \wishbone_bd_ram_mem2_reg[89][19]/P0001 , \wishbone_bd_ram_mem2_reg[89][20]/P0001 , \wishbone_bd_ram_mem2_reg[89][21]/P0001 , \wishbone_bd_ram_mem2_reg[89][22]/P0001 , \wishbone_bd_ram_mem2_reg[89][23]/P0001 , \wishbone_bd_ram_mem2_reg[8][16]/P0001 , \wishbone_bd_ram_mem2_reg[8][17]/P0001 , \wishbone_bd_ram_mem2_reg[8][18]/P0001 , \wishbone_bd_ram_mem2_reg[8][19]/P0001 , \wishbone_bd_ram_mem2_reg[8][20]/P0001 , \wishbone_bd_ram_mem2_reg[8][21]/P0001 , \wishbone_bd_ram_mem2_reg[8][22]/P0001 , \wishbone_bd_ram_mem2_reg[8][23]/P0001 , \wishbone_bd_ram_mem2_reg[90][16]/P0001 , \wishbone_bd_ram_mem2_reg[90][17]/P0001 , \wishbone_bd_ram_mem2_reg[90][18]/P0001 , \wishbone_bd_ram_mem2_reg[90][19]/P0001 , \wishbone_bd_ram_mem2_reg[90][20]/P0001 , \wishbone_bd_ram_mem2_reg[90][21]/P0001 , \wishbone_bd_ram_mem2_reg[90][22]/P0001 , \wishbone_bd_ram_mem2_reg[90][23]/P0001 , \wishbone_bd_ram_mem2_reg[91][16]/P0001 , \wishbone_bd_ram_mem2_reg[91][17]/P0001 , \wishbone_bd_ram_mem2_reg[91][18]/P0001 , \wishbone_bd_ram_mem2_reg[91][19]/P0001 , \wishbone_bd_ram_mem2_reg[91][20]/P0001 , \wishbone_bd_ram_mem2_reg[91][21]/P0001 , \wishbone_bd_ram_mem2_reg[91][22]/P0001 , \wishbone_bd_ram_mem2_reg[91][23]/P0001 , \wishbone_bd_ram_mem2_reg[92][16]/P0001 , \wishbone_bd_ram_mem2_reg[92][17]/P0001 , \wishbone_bd_ram_mem2_reg[92][18]/P0001 , \wishbone_bd_ram_mem2_reg[92][19]/P0001 , \wishbone_bd_ram_mem2_reg[92][20]/P0001 , \wishbone_bd_ram_mem2_reg[92][21]/P0001 , \wishbone_bd_ram_mem2_reg[92][22]/P0001 , \wishbone_bd_ram_mem2_reg[92][23]/P0001 , \wishbone_bd_ram_mem2_reg[93][16]/P0001 , \wishbone_bd_ram_mem2_reg[93][17]/P0001 , \wishbone_bd_ram_mem2_reg[93][18]/P0001 , \wishbone_bd_ram_mem2_reg[93][19]/P0001 , \wishbone_bd_ram_mem2_reg[93][20]/P0001 , \wishbone_bd_ram_mem2_reg[93][21]/P0001 , \wishbone_bd_ram_mem2_reg[93][22]/P0001 , \wishbone_bd_ram_mem2_reg[93][23]/P0001 , \wishbone_bd_ram_mem2_reg[94][16]/P0001 , \wishbone_bd_ram_mem2_reg[94][17]/P0001 , \wishbone_bd_ram_mem2_reg[94][18]/P0001 , \wishbone_bd_ram_mem2_reg[94][19]/P0001 , \wishbone_bd_ram_mem2_reg[94][20]/P0001 , \wishbone_bd_ram_mem2_reg[94][21]/P0001 , \wishbone_bd_ram_mem2_reg[94][22]/P0001 , \wishbone_bd_ram_mem2_reg[94][23]/P0001 , \wishbone_bd_ram_mem2_reg[95][16]/P0001 , \wishbone_bd_ram_mem2_reg[95][17]/P0001 , \wishbone_bd_ram_mem2_reg[95][18]/P0001 , \wishbone_bd_ram_mem2_reg[95][19]/P0001 , \wishbone_bd_ram_mem2_reg[95][20]/P0001 , \wishbone_bd_ram_mem2_reg[95][21]/P0001 , \wishbone_bd_ram_mem2_reg[95][22]/P0001 , \wishbone_bd_ram_mem2_reg[95][23]/P0001 , \wishbone_bd_ram_mem2_reg[96][16]/P0001 , \wishbone_bd_ram_mem2_reg[96][17]/P0001 , \wishbone_bd_ram_mem2_reg[96][18]/P0001 , \wishbone_bd_ram_mem2_reg[96][19]/P0001 , \wishbone_bd_ram_mem2_reg[96][20]/P0001 , \wishbone_bd_ram_mem2_reg[96][21]/P0001 , \wishbone_bd_ram_mem2_reg[96][22]/P0001 , \wishbone_bd_ram_mem2_reg[96][23]/P0001 , \wishbone_bd_ram_mem2_reg[97][16]/P0001 , \wishbone_bd_ram_mem2_reg[97][17]/P0001 , \wishbone_bd_ram_mem2_reg[97][18]/P0001 , \wishbone_bd_ram_mem2_reg[97][19]/P0001 , \wishbone_bd_ram_mem2_reg[97][20]/P0001 , \wishbone_bd_ram_mem2_reg[97][21]/P0001 , \wishbone_bd_ram_mem2_reg[97][22]/P0001 , \wishbone_bd_ram_mem2_reg[97][23]/P0001 , \wishbone_bd_ram_mem2_reg[98][16]/P0001 , \wishbone_bd_ram_mem2_reg[98][17]/P0001 , \wishbone_bd_ram_mem2_reg[98][18]/P0001 , \wishbone_bd_ram_mem2_reg[98][19]/P0001 , \wishbone_bd_ram_mem2_reg[98][20]/P0001 , \wishbone_bd_ram_mem2_reg[98][21]/P0001 , \wishbone_bd_ram_mem2_reg[98][22]/P0001 , \wishbone_bd_ram_mem2_reg[98][23]/P0001 , \wishbone_bd_ram_mem2_reg[99][16]/P0001 , \wishbone_bd_ram_mem2_reg[99][17]/P0001 , \wishbone_bd_ram_mem2_reg[99][18]/P0001 , \wishbone_bd_ram_mem2_reg[99][19]/P0001 , \wishbone_bd_ram_mem2_reg[99][20]/P0001 , \wishbone_bd_ram_mem2_reg[99][21]/P0001 , \wishbone_bd_ram_mem2_reg[99][22]/P0001 , \wishbone_bd_ram_mem2_reg[99][23]/P0001 , \wishbone_bd_ram_mem2_reg[9][16]/P0001 , \wishbone_bd_ram_mem2_reg[9][17]/P0001 , \wishbone_bd_ram_mem2_reg[9][18]/P0001 , \wishbone_bd_ram_mem2_reg[9][19]/P0001 , \wishbone_bd_ram_mem2_reg[9][20]/P0001 , \wishbone_bd_ram_mem2_reg[9][21]/P0001 , \wishbone_bd_ram_mem2_reg[9][22]/P0001 , \wishbone_bd_ram_mem2_reg[9][23]/P0001 , \wishbone_bd_ram_mem3_reg[0][24]/P0001 , \wishbone_bd_ram_mem3_reg[0][25]/P0001 , \wishbone_bd_ram_mem3_reg[0][26]/P0001 , \wishbone_bd_ram_mem3_reg[0][27]/P0001 , \wishbone_bd_ram_mem3_reg[0][28]/P0001 , \wishbone_bd_ram_mem3_reg[0][29]/P0001 , \wishbone_bd_ram_mem3_reg[0][30]/P0001 , \wishbone_bd_ram_mem3_reg[0][31]/P0001 , \wishbone_bd_ram_mem3_reg[100][24]/P0001 , \wishbone_bd_ram_mem3_reg[100][25]/P0001 , \wishbone_bd_ram_mem3_reg[100][26]/P0001 , \wishbone_bd_ram_mem3_reg[100][27]/P0001 , \wishbone_bd_ram_mem3_reg[100][28]/P0001 , \wishbone_bd_ram_mem3_reg[100][29]/P0001 , \wishbone_bd_ram_mem3_reg[100][30]/P0001 , \wishbone_bd_ram_mem3_reg[100][31]/P0001 , \wishbone_bd_ram_mem3_reg[101][24]/P0001 , \wishbone_bd_ram_mem3_reg[101][25]/P0001 , \wishbone_bd_ram_mem3_reg[101][26]/P0001 , \wishbone_bd_ram_mem3_reg[101][27]/P0001 , \wishbone_bd_ram_mem3_reg[101][28]/P0001 , \wishbone_bd_ram_mem3_reg[101][29]/P0001 , \wishbone_bd_ram_mem3_reg[101][30]/P0001 , \wishbone_bd_ram_mem3_reg[101][31]/P0001 , \wishbone_bd_ram_mem3_reg[102][24]/P0001 , \wishbone_bd_ram_mem3_reg[102][25]/P0001 , \wishbone_bd_ram_mem3_reg[102][26]/P0001 , \wishbone_bd_ram_mem3_reg[102][27]/P0001 , \wishbone_bd_ram_mem3_reg[102][28]/P0001 , \wishbone_bd_ram_mem3_reg[102][29]/P0001 , \wishbone_bd_ram_mem3_reg[102][30]/P0001 , \wishbone_bd_ram_mem3_reg[102][31]/P0001 , \wishbone_bd_ram_mem3_reg[103][24]/P0001 , \wishbone_bd_ram_mem3_reg[103][25]/P0001 , \wishbone_bd_ram_mem3_reg[103][26]/P0001 , \wishbone_bd_ram_mem3_reg[103][27]/P0001 , \wishbone_bd_ram_mem3_reg[103][28]/P0001 , \wishbone_bd_ram_mem3_reg[103][29]/P0001 , \wishbone_bd_ram_mem3_reg[103][30]/P0001 , \wishbone_bd_ram_mem3_reg[103][31]/P0001 , \wishbone_bd_ram_mem3_reg[104][24]/P0001 , \wishbone_bd_ram_mem3_reg[104][25]/P0001 , \wishbone_bd_ram_mem3_reg[104][26]/P0001 , \wishbone_bd_ram_mem3_reg[104][27]/P0001 , \wishbone_bd_ram_mem3_reg[104][28]/P0001 , \wishbone_bd_ram_mem3_reg[104][29]/P0001 , \wishbone_bd_ram_mem3_reg[104][30]/P0001 , \wishbone_bd_ram_mem3_reg[104][31]/P0001 , \wishbone_bd_ram_mem3_reg[105][24]/P0001 , \wishbone_bd_ram_mem3_reg[105][25]/P0001 , \wishbone_bd_ram_mem3_reg[105][26]/P0001 , \wishbone_bd_ram_mem3_reg[105][27]/P0001 , \wishbone_bd_ram_mem3_reg[105][28]/P0001 , \wishbone_bd_ram_mem3_reg[105][29]/P0001 , \wishbone_bd_ram_mem3_reg[105][30]/P0001 , \wishbone_bd_ram_mem3_reg[105][31]/P0001 , \wishbone_bd_ram_mem3_reg[106][24]/P0001 , \wishbone_bd_ram_mem3_reg[106][25]/P0001 , \wishbone_bd_ram_mem3_reg[106][26]/P0001 , \wishbone_bd_ram_mem3_reg[106][27]/P0001 , \wishbone_bd_ram_mem3_reg[106][28]/P0001 , \wishbone_bd_ram_mem3_reg[106][29]/P0001 , \wishbone_bd_ram_mem3_reg[106][30]/P0001 , \wishbone_bd_ram_mem3_reg[106][31]/P0001 , \wishbone_bd_ram_mem3_reg[107][24]/P0001 , \wishbone_bd_ram_mem3_reg[107][25]/P0001 , \wishbone_bd_ram_mem3_reg[107][26]/P0001 , \wishbone_bd_ram_mem3_reg[107][27]/P0001 , \wishbone_bd_ram_mem3_reg[107][28]/P0001 , \wishbone_bd_ram_mem3_reg[107][29]/P0001 , \wishbone_bd_ram_mem3_reg[107][30]/P0001 , \wishbone_bd_ram_mem3_reg[107][31]/P0001 , \wishbone_bd_ram_mem3_reg[108][24]/P0001 , \wishbone_bd_ram_mem3_reg[108][25]/P0001 , \wishbone_bd_ram_mem3_reg[108][26]/P0001 , \wishbone_bd_ram_mem3_reg[108][27]/P0001 , \wishbone_bd_ram_mem3_reg[108][28]/P0001 , \wishbone_bd_ram_mem3_reg[108][29]/P0001 , \wishbone_bd_ram_mem3_reg[108][30]/P0001 , \wishbone_bd_ram_mem3_reg[108][31]/P0001 , \wishbone_bd_ram_mem3_reg[109][24]/P0001 , \wishbone_bd_ram_mem3_reg[109][25]/P0001 , \wishbone_bd_ram_mem3_reg[109][26]/P0001 , \wishbone_bd_ram_mem3_reg[109][27]/P0001 , \wishbone_bd_ram_mem3_reg[109][28]/P0001 , \wishbone_bd_ram_mem3_reg[109][29]/P0001 , \wishbone_bd_ram_mem3_reg[109][30]/P0001 , \wishbone_bd_ram_mem3_reg[109][31]/P0001 , \wishbone_bd_ram_mem3_reg[10][24]/P0001 , \wishbone_bd_ram_mem3_reg[10][25]/P0001 , \wishbone_bd_ram_mem3_reg[10][26]/P0001 , \wishbone_bd_ram_mem3_reg[10][27]/P0001 , \wishbone_bd_ram_mem3_reg[10][28]/P0001 , \wishbone_bd_ram_mem3_reg[10][29]/P0001 , \wishbone_bd_ram_mem3_reg[10][30]/P0001 , \wishbone_bd_ram_mem3_reg[10][31]/P0001 , \wishbone_bd_ram_mem3_reg[110][24]/P0001 , \wishbone_bd_ram_mem3_reg[110][25]/P0001 , \wishbone_bd_ram_mem3_reg[110][26]/P0001 , \wishbone_bd_ram_mem3_reg[110][27]/P0001 , \wishbone_bd_ram_mem3_reg[110][28]/P0001 , \wishbone_bd_ram_mem3_reg[110][29]/P0001 , \wishbone_bd_ram_mem3_reg[110][30]/P0001 , \wishbone_bd_ram_mem3_reg[110][31]/P0001 , \wishbone_bd_ram_mem3_reg[111][24]/P0001 , \wishbone_bd_ram_mem3_reg[111][25]/P0001 , \wishbone_bd_ram_mem3_reg[111][26]/P0001 , \wishbone_bd_ram_mem3_reg[111][27]/P0001 , \wishbone_bd_ram_mem3_reg[111][28]/P0001 , \wishbone_bd_ram_mem3_reg[111][29]/P0001 , \wishbone_bd_ram_mem3_reg[111][30]/P0001 , \wishbone_bd_ram_mem3_reg[111][31]/P0001 , \wishbone_bd_ram_mem3_reg[112][24]/P0001 , \wishbone_bd_ram_mem3_reg[112][25]/P0001 , \wishbone_bd_ram_mem3_reg[112][26]/P0001 , \wishbone_bd_ram_mem3_reg[112][27]/P0001 , \wishbone_bd_ram_mem3_reg[112][28]/P0001 , \wishbone_bd_ram_mem3_reg[112][29]/P0001 , \wishbone_bd_ram_mem3_reg[112][30]/P0001 , \wishbone_bd_ram_mem3_reg[112][31]/P0001 , \wishbone_bd_ram_mem3_reg[113][24]/P0001 , \wishbone_bd_ram_mem3_reg[113][25]/P0001 , \wishbone_bd_ram_mem3_reg[113][26]/P0001 , \wishbone_bd_ram_mem3_reg[113][27]/P0001 , \wishbone_bd_ram_mem3_reg[113][28]/P0001 , \wishbone_bd_ram_mem3_reg[113][29]/P0001 , \wishbone_bd_ram_mem3_reg[113][30]/P0001 , \wishbone_bd_ram_mem3_reg[113][31]/P0001 , \wishbone_bd_ram_mem3_reg[114][24]/P0001 , \wishbone_bd_ram_mem3_reg[114][25]/P0001 , \wishbone_bd_ram_mem3_reg[114][26]/P0001 , \wishbone_bd_ram_mem3_reg[114][27]/P0001 , \wishbone_bd_ram_mem3_reg[114][28]/P0001 , \wishbone_bd_ram_mem3_reg[114][29]/P0001 , \wishbone_bd_ram_mem3_reg[114][30]/P0001 , \wishbone_bd_ram_mem3_reg[114][31]/P0001 , \wishbone_bd_ram_mem3_reg[115][24]/P0001 , \wishbone_bd_ram_mem3_reg[115][25]/P0001 , \wishbone_bd_ram_mem3_reg[115][26]/P0001 , \wishbone_bd_ram_mem3_reg[115][27]/P0001 , \wishbone_bd_ram_mem3_reg[115][28]/P0001 , \wishbone_bd_ram_mem3_reg[115][29]/P0001 , \wishbone_bd_ram_mem3_reg[115][30]/P0001 , \wishbone_bd_ram_mem3_reg[115][31]/P0001 , \wishbone_bd_ram_mem3_reg[116][24]/P0001 , \wishbone_bd_ram_mem3_reg[116][25]/P0001 , \wishbone_bd_ram_mem3_reg[116][26]/P0001 , \wishbone_bd_ram_mem3_reg[116][27]/P0001 , \wishbone_bd_ram_mem3_reg[116][28]/P0001 , \wishbone_bd_ram_mem3_reg[116][29]/P0001 , \wishbone_bd_ram_mem3_reg[116][30]/P0001 , \wishbone_bd_ram_mem3_reg[116][31]/P0001 , \wishbone_bd_ram_mem3_reg[117][24]/P0001 , \wishbone_bd_ram_mem3_reg[117][25]/P0001 , \wishbone_bd_ram_mem3_reg[117][26]/P0001 , \wishbone_bd_ram_mem3_reg[117][27]/P0001 , \wishbone_bd_ram_mem3_reg[117][28]/P0001 , \wishbone_bd_ram_mem3_reg[117][29]/P0001 , \wishbone_bd_ram_mem3_reg[117][30]/P0001 , \wishbone_bd_ram_mem3_reg[117][31]/P0001 , \wishbone_bd_ram_mem3_reg[118][24]/P0001 , \wishbone_bd_ram_mem3_reg[118][25]/P0001 , \wishbone_bd_ram_mem3_reg[118][26]/P0001 , \wishbone_bd_ram_mem3_reg[118][27]/P0001 , \wishbone_bd_ram_mem3_reg[118][28]/P0001 , \wishbone_bd_ram_mem3_reg[118][29]/P0001 , \wishbone_bd_ram_mem3_reg[118][30]/P0001 , \wishbone_bd_ram_mem3_reg[118][31]/P0001 , \wishbone_bd_ram_mem3_reg[119][24]/P0001 , \wishbone_bd_ram_mem3_reg[119][25]/P0001 , \wishbone_bd_ram_mem3_reg[119][26]/P0001 , \wishbone_bd_ram_mem3_reg[119][27]/P0001 , \wishbone_bd_ram_mem3_reg[119][28]/P0001 , \wishbone_bd_ram_mem3_reg[119][29]/P0001 , \wishbone_bd_ram_mem3_reg[119][30]/P0001 , \wishbone_bd_ram_mem3_reg[119][31]/P0001 , \wishbone_bd_ram_mem3_reg[11][24]/P0001 , \wishbone_bd_ram_mem3_reg[11][25]/P0001 , \wishbone_bd_ram_mem3_reg[11][26]/P0001 , \wishbone_bd_ram_mem3_reg[11][27]/P0001 , \wishbone_bd_ram_mem3_reg[11][28]/P0001 , \wishbone_bd_ram_mem3_reg[11][29]/P0001 , \wishbone_bd_ram_mem3_reg[11][30]/P0001 , \wishbone_bd_ram_mem3_reg[11][31]/P0001 , \wishbone_bd_ram_mem3_reg[120][24]/P0001 , \wishbone_bd_ram_mem3_reg[120][25]/P0001 , \wishbone_bd_ram_mem3_reg[120][26]/P0001 , \wishbone_bd_ram_mem3_reg[120][27]/P0001 , \wishbone_bd_ram_mem3_reg[120][28]/P0001 , \wishbone_bd_ram_mem3_reg[120][29]/P0001 , \wishbone_bd_ram_mem3_reg[120][30]/P0001 , \wishbone_bd_ram_mem3_reg[120][31]/P0001 , \wishbone_bd_ram_mem3_reg[121][24]/P0001 , \wishbone_bd_ram_mem3_reg[121][25]/P0001 , \wishbone_bd_ram_mem3_reg[121][26]/P0001 , \wishbone_bd_ram_mem3_reg[121][27]/P0001 , \wishbone_bd_ram_mem3_reg[121][28]/P0001 , \wishbone_bd_ram_mem3_reg[121][29]/P0001 , \wishbone_bd_ram_mem3_reg[121][30]/P0001 , \wishbone_bd_ram_mem3_reg[121][31]/P0001 , \wishbone_bd_ram_mem3_reg[122][24]/P0001 , \wishbone_bd_ram_mem3_reg[122][25]/P0001 , \wishbone_bd_ram_mem3_reg[122][26]/P0001 , \wishbone_bd_ram_mem3_reg[122][27]/P0001 , \wishbone_bd_ram_mem3_reg[122][28]/P0001 , \wishbone_bd_ram_mem3_reg[122][29]/P0001 , \wishbone_bd_ram_mem3_reg[122][30]/P0001 , \wishbone_bd_ram_mem3_reg[122][31]/P0001 , \wishbone_bd_ram_mem3_reg[123][24]/P0001 , \wishbone_bd_ram_mem3_reg[123][25]/P0001 , \wishbone_bd_ram_mem3_reg[123][26]/P0001 , \wishbone_bd_ram_mem3_reg[123][27]/P0001 , \wishbone_bd_ram_mem3_reg[123][28]/P0001 , \wishbone_bd_ram_mem3_reg[123][29]/P0001 , \wishbone_bd_ram_mem3_reg[123][30]/P0001 , \wishbone_bd_ram_mem3_reg[123][31]/P0001 , \wishbone_bd_ram_mem3_reg[124][24]/P0001 , \wishbone_bd_ram_mem3_reg[124][25]/P0001 , \wishbone_bd_ram_mem3_reg[124][26]/P0001 , \wishbone_bd_ram_mem3_reg[124][27]/P0001 , \wishbone_bd_ram_mem3_reg[124][28]/P0001 , \wishbone_bd_ram_mem3_reg[124][29]/P0001 , \wishbone_bd_ram_mem3_reg[124][30]/P0001 , \wishbone_bd_ram_mem3_reg[124][31]/P0001 , \wishbone_bd_ram_mem3_reg[125][24]/P0001 , \wishbone_bd_ram_mem3_reg[125][25]/P0001 , \wishbone_bd_ram_mem3_reg[125][26]/P0001 , \wishbone_bd_ram_mem3_reg[125][27]/P0001 , \wishbone_bd_ram_mem3_reg[125][28]/P0001 , \wishbone_bd_ram_mem3_reg[125][29]/P0001 , \wishbone_bd_ram_mem3_reg[125][30]/P0001 , \wishbone_bd_ram_mem3_reg[125][31]/P0001 , \wishbone_bd_ram_mem3_reg[126][24]/P0001 , \wishbone_bd_ram_mem3_reg[126][25]/P0001 , \wishbone_bd_ram_mem3_reg[126][26]/P0001 , \wishbone_bd_ram_mem3_reg[126][27]/P0001 , \wishbone_bd_ram_mem3_reg[126][28]/P0001 , \wishbone_bd_ram_mem3_reg[126][29]/P0001 , \wishbone_bd_ram_mem3_reg[126][30]/P0001 , \wishbone_bd_ram_mem3_reg[126][31]/P0001 , \wishbone_bd_ram_mem3_reg[127][24]/P0001 , \wishbone_bd_ram_mem3_reg[127][25]/P0001 , \wishbone_bd_ram_mem3_reg[127][26]/P0001 , \wishbone_bd_ram_mem3_reg[127][27]/P0001 , \wishbone_bd_ram_mem3_reg[127][28]/P0001 , \wishbone_bd_ram_mem3_reg[127][29]/P0001 , \wishbone_bd_ram_mem3_reg[127][30]/P0001 , \wishbone_bd_ram_mem3_reg[127][31]/P0001 , \wishbone_bd_ram_mem3_reg[128][24]/P0001 , \wishbone_bd_ram_mem3_reg[128][25]/P0001 , \wishbone_bd_ram_mem3_reg[128][26]/P0001 , \wishbone_bd_ram_mem3_reg[128][27]/P0001 , \wishbone_bd_ram_mem3_reg[128][28]/P0001 , \wishbone_bd_ram_mem3_reg[128][29]/P0001 , \wishbone_bd_ram_mem3_reg[128][30]/P0001 , \wishbone_bd_ram_mem3_reg[128][31]/P0001 , \wishbone_bd_ram_mem3_reg[129][24]/P0001 , \wishbone_bd_ram_mem3_reg[129][25]/P0001 , \wishbone_bd_ram_mem3_reg[129][26]/P0001 , \wishbone_bd_ram_mem3_reg[129][27]/P0001 , \wishbone_bd_ram_mem3_reg[129][28]/P0001 , \wishbone_bd_ram_mem3_reg[129][29]/P0001 , \wishbone_bd_ram_mem3_reg[129][30]/P0001 , \wishbone_bd_ram_mem3_reg[129][31]/P0001 , \wishbone_bd_ram_mem3_reg[12][24]/P0001 , \wishbone_bd_ram_mem3_reg[12][25]/P0001 , \wishbone_bd_ram_mem3_reg[12][26]/P0001 , \wishbone_bd_ram_mem3_reg[12][27]/P0001 , \wishbone_bd_ram_mem3_reg[12][28]/P0001 , \wishbone_bd_ram_mem3_reg[12][29]/P0001 , \wishbone_bd_ram_mem3_reg[12][30]/P0001 , \wishbone_bd_ram_mem3_reg[12][31]/P0001 , \wishbone_bd_ram_mem3_reg[130][24]/P0001 , \wishbone_bd_ram_mem3_reg[130][25]/P0001 , \wishbone_bd_ram_mem3_reg[130][26]/P0001 , \wishbone_bd_ram_mem3_reg[130][27]/P0001 , \wishbone_bd_ram_mem3_reg[130][28]/P0001 , \wishbone_bd_ram_mem3_reg[130][29]/P0001 , \wishbone_bd_ram_mem3_reg[130][30]/P0001 , \wishbone_bd_ram_mem3_reg[130][31]/P0001 , \wishbone_bd_ram_mem3_reg[131][24]/P0001 , \wishbone_bd_ram_mem3_reg[131][25]/P0001 , \wishbone_bd_ram_mem3_reg[131][26]/P0001 , \wishbone_bd_ram_mem3_reg[131][27]/P0001 , \wishbone_bd_ram_mem3_reg[131][28]/P0001 , \wishbone_bd_ram_mem3_reg[131][29]/P0001 , \wishbone_bd_ram_mem3_reg[131][30]/P0001 , \wishbone_bd_ram_mem3_reg[131][31]/P0001 , \wishbone_bd_ram_mem3_reg[132][24]/P0001 , \wishbone_bd_ram_mem3_reg[132][25]/P0001 , \wishbone_bd_ram_mem3_reg[132][26]/P0001 , \wishbone_bd_ram_mem3_reg[132][27]/P0001 , \wishbone_bd_ram_mem3_reg[132][28]/P0001 , \wishbone_bd_ram_mem3_reg[132][29]/P0001 , \wishbone_bd_ram_mem3_reg[132][30]/P0001 , \wishbone_bd_ram_mem3_reg[132][31]/P0001 , \wishbone_bd_ram_mem3_reg[133][24]/P0001 , \wishbone_bd_ram_mem3_reg[133][25]/P0001 , \wishbone_bd_ram_mem3_reg[133][26]/P0001 , \wishbone_bd_ram_mem3_reg[133][27]/P0001 , \wishbone_bd_ram_mem3_reg[133][28]/P0001 , \wishbone_bd_ram_mem3_reg[133][29]/P0001 , \wishbone_bd_ram_mem3_reg[133][30]/P0001 , \wishbone_bd_ram_mem3_reg[133][31]/P0001 , \wishbone_bd_ram_mem3_reg[134][24]/P0001 , \wishbone_bd_ram_mem3_reg[134][25]/P0001 , \wishbone_bd_ram_mem3_reg[134][26]/P0001 , \wishbone_bd_ram_mem3_reg[134][27]/P0001 , \wishbone_bd_ram_mem3_reg[134][28]/P0001 , \wishbone_bd_ram_mem3_reg[134][29]/P0001 , \wishbone_bd_ram_mem3_reg[134][30]/P0001 , \wishbone_bd_ram_mem3_reg[134][31]/P0001 , \wishbone_bd_ram_mem3_reg[135][24]/P0001 , \wishbone_bd_ram_mem3_reg[135][25]/P0001 , \wishbone_bd_ram_mem3_reg[135][26]/P0001 , \wishbone_bd_ram_mem3_reg[135][27]/P0001 , \wishbone_bd_ram_mem3_reg[135][28]/P0001 , \wishbone_bd_ram_mem3_reg[135][29]/P0001 , \wishbone_bd_ram_mem3_reg[135][30]/P0001 , \wishbone_bd_ram_mem3_reg[135][31]/P0001 , \wishbone_bd_ram_mem3_reg[136][24]/P0001 , \wishbone_bd_ram_mem3_reg[136][25]/P0001 , \wishbone_bd_ram_mem3_reg[136][26]/P0001 , \wishbone_bd_ram_mem3_reg[136][27]/P0001 , \wishbone_bd_ram_mem3_reg[136][28]/P0001 , \wishbone_bd_ram_mem3_reg[136][29]/P0001 , \wishbone_bd_ram_mem3_reg[136][30]/P0001 , \wishbone_bd_ram_mem3_reg[136][31]/P0001 , \wishbone_bd_ram_mem3_reg[137][24]/P0001 , \wishbone_bd_ram_mem3_reg[137][25]/P0001 , \wishbone_bd_ram_mem3_reg[137][26]/P0001 , \wishbone_bd_ram_mem3_reg[137][27]/P0001 , \wishbone_bd_ram_mem3_reg[137][28]/P0001 , \wishbone_bd_ram_mem3_reg[137][29]/P0001 , \wishbone_bd_ram_mem3_reg[137][30]/P0001 , \wishbone_bd_ram_mem3_reg[137][31]/P0001 , \wishbone_bd_ram_mem3_reg[138][24]/P0001 , \wishbone_bd_ram_mem3_reg[138][25]/P0001 , \wishbone_bd_ram_mem3_reg[138][26]/P0001 , \wishbone_bd_ram_mem3_reg[138][27]/P0001 , \wishbone_bd_ram_mem3_reg[138][28]/P0001 , \wishbone_bd_ram_mem3_reg[138][29]/P0001 , \wishbone_bd_ram_mem3_reg[138][30]/P0001 , \wishbone_bd_ram_mem3_reg[138][31]/P0001 , \wishbone_bd_ram_mem3_reg[139][24]/P0001 , \wishbone_bd_ram_mem3_reg[139][25]/P0001 , \wishbone_bd_ram_mem3_reg[139][26]/P0001 , \wishbone_bd_ram_mem3_reg[139][27]/P0001 , \wishbone_bd_ram_mem3_reg[139][28]/P0001 , \wishbone_bd_ram_mem3_reg[139][29]/P0001 , \wishbone_bd_ram_mem3_reg[139][30]/P0001 , \wishbone_bd_ram_mem3_reg[139][31]/P0001 , \wishbone_bd_ram_mem3_reg[13][24]/P0001 , \wishbone_bd_ram_mem3_reg[13][25]/P0001 , \wishbone_bd_ram_mem3_reg[13][26]/P0001 , \wishbone_bd_ram_mem3_reg[13][27]/P0001 , \wishbone_bd_ram_mem3_reg[13][28]/P0001 , \wishbone_bd_ram_mem3_reg[13][29]/P0001 , \wishbone_bd_ram_mem3_reg[13][30]/P0001 , \wishbone_bd_ram_mem3_reg[13][31]/P0001 , \wishbone_bd_ram_mem3_reg[140][24]/P0001 , \wishbone_bd_ram_mem3_reg[140][25]/P0001 , \wishbone_bd_ram_mem3_reg[140][26]/P0001 , \wishbone_bd_ram_mem3_reg[140][27]/P0001 , \wishbone_bd_ram_mem3_reg[140][28]/P0001 , \wishbone_bd_ram_mem3_reg[140][29]/P0001 , \wishbone_bd_ram_mem3_reg[140][30]/P0001 , \wishbone_bd_ram_mem3_reg[140][31]/P0001 , \wishbone_bd_ram_mem3_reg[141][24]/P0001 , \wishbone_bd_ram_mem3_reg[141][25]/P0001 , \wishbone_bd_ram_mem3_reg[141][26]/P0001 , \wishbone_bd_ram_mem3_reg[141][27]/P0001 , \wishbone_bd_ram_mem3_reg[141][28]/P0001 , \wishbone_bd_ram_mem3_reg[141][29]/P0001 , \wishbone_bd_ram_mem3_reg[141][30]/P0001 , \wishbone_bd_ram_mem3_reg[141][31]/P0001 , \wishbone_bd_ram_mem3_reg[142][24]/P0001 , \wishbone_bd_ram_mem3_reg[142][25]/P0001 , \wishbone_bd_ram_mem3_reg[142][26]/P0001 , \wishbone_bd_ram_mem3_reg[142][27]/P0001 , \wishbone_bd_ram_mem3_reg[142][28]/P0001 , \wishbone_bd_ram_mem3_reg[142][29]/P0001 , \wishbone_bd_ram_mem3_reg[142][30]/P0001 , \wishbone_bd_ram_mem3_reg[142][31]/P0001 , \wishbone_bd_ram_mem3_reg[143][24]/P0001 , \wishbone_bd_ram_mem3_reg[143][25]/P0001 , \wishbone_bd_ram_mem3_reg[143][26]/P0001 , \wishbone_bd_ram_mem3_reg[143][27]/P0001 , \wishbone_bd_ram_mem3_reg[143][28]/P0001 , \wishbone_bd_ram_mem3_reg[143][29]/P0001 , \wishbone_bd_ram_mem3_reg[143][30]/P0001 , \wishbone_bd_ram_mem3_reg[143][31]/P0001 , \wishbone_bd_ram_mem3_reg[144][24]/P0001 , \wishbone_bd_ram_mem3_reg[144][25]/P0001 , \wishbone_bd_ram_mem3_reg[144][26]/P0001 , \wishbone_bd_ram_mem3_reg[144][27]/P0001 , \wishbone_bd_ram_mem3_reg[144][28]/P0001 , \wishbone_bd_ram_mem3_reg[144][29]/P0001 , \wishbone_bd_ram_mem3_reg[144][30]/P0001 , \wishbone_bd_ram_mem3_reg[144][31]/P0001 , \wishbone_bd_ram_mem3_reg[145][24]/P0001 , \wishbone_bd_ram_mem3_reg[145][25]/P0001 , \wishbone_bd_ram_mem3_reg[145][26]/P0001 , \wishbone_bd_ram_mem3_reg[145][27]/P0001 , \wishbone_bd_ram_mem3_reg[145][28]/P0001 , \wishbone_bd_ram_mem3_reg[145][29]/P0001 , \wishbone_bd_ram_mem3_reg[145][30]/P0001 , \wishbone_bd_ram_mem3_reg[145][31]/P0001 , \wishbone_bd_ram_mem3_reg[146][24]/P0001 , \wishbone_bd_ram_mem3_reg[146][25]/P0001 , \wishbone_bd_ram_mem3_reg[146][26]/P0001 , \wishbone_bd_ram_mem3_reg[146][27]/P0001 , \wishbone_bd_ram_mem3_reg[146][28]/P0001 , \wishbone_bd_ram_mem3_reg[146][29]/P0001 , \wishbone_bd_ram_mem3_reg[146][30]/P0001 , \wishbone_bd_ram_mem3_reg[146][31]/P0001 , \wishbone_bd_ram_mem3_reg[147][24]/P0001 , \wishbone_bd_ram_mem3_reg[147][25]/P0001 , \wishbone_bd_ram_mem3_reg[147][26]/P0001 , \wishbone_bd_ram_mem3_reg[147][27]/P0001 , \wishbone_bd_ram_mem3_reg[147][28]/P0001 , \wishbone_bd_ram_mem3_reg[147][29]/P0001 , \wishbone_bd_ram_mem3_reg[147][30]/P0001 , \wishbone_bd_ram_mem3_reg[147][31]/P0001 , \wishbone_bd_ram_mem3_reg[148][24]/P0001 , \wishbone_bd_ram_mem3_reg[148][25]/P0001 , \wishbone_bd_ram_mem3_reg[148][26]/P0001 , \wishbone_bd_ram_mem3_reg[148][27]/P0001 , \wishbone_bd_ram_mem3_reg[148][28]/P0001 , \wishbone_bd_ram_mem3_reg[148][29]/P0001 , \wishbone_bd_ram_mem3_reg[148][30]/P0001 , \wishbone_bd_ram_mem3_reg[148][31]/P0001 , \wishbone_bd_ram_mem3_reg[149][24]/P0001 , \wishbone_bd_ram_mem3_reg[149][25]/P0001 , \wishbone_bd_ram_mem3_reg[149][26]/P0001 , \wishbone_bd_ram_mem3_reg[149][27]/P0001 , \wishbone_bd_ram_mem3_reg[149][28]/P0001 , \wishbone_bd_ram_mem3_reg[149][29]/P0001 , \wishbone_bd_ram_mem3_reg[149][30]/P0001 , \wishbone_bd_ram_mem3_reg[149][31]/P0001 , \wishbone_bd_ram_mem3_reg[14][24]/P0001 , \wishbone_bd_ram_mem3_reg[14][25]/P0001 , \wishbone_bd_ram_mem3_reg[14][26]/P0001 , \wishbone_bd_ram_mem3_reg[14][27]/P0001 , \wishbone_bd_ram_mem3_reg[14][28]/P0001 , \wishbone_bd_ram_mem3_reg[14][29]/P0001 , \wishbone_bd_ram_mem3_reg[14][30]/P0001 , \wishbone_bd_ram_mem3_reg[14][31]/P0001 , \wishbone_bd_ram_mem3_reg[150][24]/P0001 , \wishbone_bd_ram_mem3_reg[150][25]/P0001 , \wishbone_bd_ram_mem3_reg[150][26]/P0001 , \wishbone_bd_ram_mem3_reg[150][27]/P0001 , \wishbone_bd_ram_mem3_reg[150][28]/P0001 , \wishbone_bd_ram_mem3_reg[150][29]/P0001 , \wishbone_bd_ram_mem3_reg[150][30]/P0001 , \wishbone_bd_ram_mem3_reg[150][31]/P0001 , \wishbone_bd_ram_mem3_reg[151][24]/P0001 , \wishbone_bd_ram_mem3_reg[151][25]/P0001 , \wishbone_bd_ram_mem3_reg[151][26]/P0001 , \wishbone_bd_ram_mem3_reg[151][27]/P0001 , \wishbone_bd_ram_mem3_reg[151][28]/P0001 , \wishbone_bd_ram_mem3_reg[151][29]/P0001 , \wishbone_bd_ram_mem3_reg[151][30]/P0001 , \wishbone_bd_ram_mem3_reg[151][31]/P0001 , \wishbone_bd_ram_mem3_reg[152][24]/P0001 , \wishbone_bd_ram_mem3_reg[152][25]/P0001 , \wishbone_bd_ram_mem3_reg[152][26]/P0001 , \wishbone_bd_ram_mem3_reg[152][27]/P0001 , \wishbone_bd_ram_mem3_reg[152][28]/P0001 , \wishbone_bd_ram_mem3_reg[152][29]/P0001 , \wishbone_bd_ram_mem3_reg[152][30]/P0001 , \wishbone_bd_ram_mem3_reg[152][31]/P0001 , \wishbone_bd_ram_mem3_reg[153][24]/P0001 , \wishbone_bd_ram_mem3_reg[153][25]/P0001 , \wishbone_bd_ram_mem3_reg[153][26]/P0001 , \wishbone_bd_ram_mem3_reg[153][27]/P0001 , \wishbone_bd_ram_mem3_reg[153][28]/P0001 , \wishbone_bd_ram_mem3_reg[153][29]/P0001 , \wishbone_bd_ram_mem3_reg[153][30]/P0001 , \wishbone_bd_ram_mem3_reg[153][31]/P0001 , \wishbone_bd_ram_mem3_reg[154][24]/P0001 , \wishbone_bd_ram_mem3_reg[154][25]/P0001 , \wishbone_bd_ram_mem3_reg[154][26]/P0001 , \wishbone_bd_ram_mem3_reg[154][27]/P0001 , \wishbone_bd_ram_mem3_reg[154][28]/P0001 , \wishbone_bd_ram_mem3_reg[154][29]/P0001 , \wishbone_bd_ram_mem3_reg[154][30]/P0001 , \wishbone_bd_ram_mem3_reg[154][31]/P0001 , \wishbone_bd_ram_mem3_reg[155][24]/P0001 , \wishbone_bd_ram_mem3_reg[155][25]/P0001 , \wishbone_bd_ram_mem3_reg[155][26]/P0001 , \wishbone_bd_ram_mem3_reg[155][27]/P0001 , \wishbone_bd_ram_mem3_reg[155][28]/P0001 , \wishbone_bd_ram_mem3_reg[155][29]/P0001 , \wishbone_bd_ram_mem3_reg[155][30]/P0001 , \wishbone_bd_ram_mem3_reg[155][31]/P0001 , \wishbone_bd_ram_mem3_reg[156][24]/P0001 , \wishbone_bd_ram_mem3_reg[156][25]/P0001 , \wishbone_bd_ram_mem3_reg[156][26]/P0001 , \wishbone_bd_ram_mem3_reg[156][27]/P0001 , \wishbone_bd_ram_mem3_reg[156][28]/P0001 , \wishbone_bd_ram_mem3_reg[156][29]/P0001 , \wishbone_bd_ram_mem3_reg[156][30]/P0001 , \wishbone_bd_ram_mem3_reg[156][31]/P0001 , \wishbone_bd_ram_mem3_reg[157][24]/P0001 , \wishbone_bd_ram_mem3_reg[157][25]/P0001 , \wishbone_bd_ram_mem3_reg[157][26]/P0001 , \wishbone_bd_ram_mem3_reg[157][27]/P0001 , \wishbone_bd_ram_mem3_reg[157][28]/P0001 , \wishbone_bd_ram_mem3_reg[157][29]/P0001 , \wishbone_bd_ram_mem3_reg[157][30]/P0001 , \wishbone_bd_ram_mem3_reg[157][31]/P0001 , \wishbone_bd_ram_mem3_reg[158][24]/P0001 , \wishbone_bd_ram_mem3_reg[158][25]/P0001 , \wishbone_bd_ram_mem3_reg[158][26]/P0001 , \wishbone_bd_ram_mem3_reg[158][27]/P0001 , \wishbone_bd_ram_mem3_reg[158][28]/P0001 , \wishbone_bd_ram_mem3_reg[158][29]/P0001 , \wishbone_bd_ram_mem3_reg[158][30]/P0001 , \wishbone_bd_ram_mem3_reg[158][31]/P0001 , \wishbone_bd_ram_mem3_reg[159][24]/P0001 , \wishbone_bd_ram_mem3_reg[159][25]/P0001 , \wishbone_bd_ram_mem3_reg[159][26]/P0001 , \wishbone_bd_ram_mem3_reg[159][27]/P0001 , \wishbone_bd_ram_mem3_reg[159][28]/P0001 , \wishbone_bd_ram_mem3_reg[159][29]/P0001 , \wishbone_bd_ram_mem3_reg[159][30]/P0001 , \wishbone_bd_ram_mem3_reg[159][31]/P0001 , \wishbone_bd_ram_mem3_reg[15][24]/P0001 , \wishbone_bd_ram_mem3_reg[15][25]/P0001 , \wishbone_bd_ram_mem3_reg[15][26]/P0001 , \wishbone_bd_ram_mem3_reg[15][27]/P0001 , \wishbone_bd_ram_mem3_reg[15][28]/P0001 , \wishbone_bd_ram_mem3_reg[15][29]/P0001 , \wishbone_bd_ram_mem3_reg[15][30]/P0001 , \wishbone_bd_ram_mem3_reg[15][31]/P0001 , \wishbone_bd_ram_mem3_reg[160][24]/P0001 , \wishbone_bd_ram_mem3_reg[160][25]/P0001 , \wishbone_bd_ram_mem3_reg[160][26]/P0001 , \wishbone_bd_ram_mem3_reg[160][27]/P0001 , \wishbone_bd_ram_mem3_reg[160][28]/P0001 , \wishbone_bd_ram_mem3_reg[160][29]/P0001 , \wishbone_bd_ram_mem3_reg[160][30]/P0001 , \wishbone_bd_ram_mem3_reg[160][31]/P0001 , \wishbone_bd_ram_mem3_reg[161][24]/P0001 , \wishbone_bd_ram_mem3_reg[161][25]/P0001 , \wishbone_bd_ram_mem3_reg[161][26]/P0001 , \wishbone_bd_ram_mem3_reg[161][27]/P0001 , \wishbone_bd_ram_mem3_reg[161][28]/P0001 , \wishbone_bd_ram_mem3_reg[161][29]/P0001 , \wishbone_bd_ram_mem3_reg[161][30]/P0001 , \wishbone_bd_ram_mem3_reg[161][31]/P0001 , \wishbone_bd_ram_mem3_reg[162][24]/P0001 , \wishbone_bd_ram_mem3_reg[162][25]/P0001 , \wishbone_bd_ram_mem3_reg[162][26]/P0001 , \wishbone_bd_ram_mem3_reg[162][27]/P0001 , \wishbone_bd_ram_mem3_reg[162][28]/P0001 , \wishbone_bd_ram_mem3_reg[162][29]/P0001 , \wishbone_bd_ram_mem3_reg[162][30]/P0001 , \wishbone_bd_ram_mem3_reg[162][31]/P0001 , \wishbone_bd_ram_mem3_reg[163][24]/P0001 , \wishbone_bd_ram_mem3_reg[163][25]/P0001 , \wishbone_bd_ram_mem3_reg[163][26]/P0001 , \wishbone_bd_ram_mem3_reg[163][27]/P0001 , \wishbone_bd_ram_mem3_reg[163][28]/P0001 , \wishbone_bd_ram_mem3_reg[163][29]/P0001 , \wishbone_bd_ram_mem3_reg[163][30]/P0001 , \wishbone_bd_ram_mem3_reg[163][31]/P0001 , \wishbone_bd_ram_mem3_reg[164][24]/P0001 , \wishbone_bd_ram_mem3_reg[164][25]/P0001 , \wishbone_bd_ram_mem3_reg[164][26]/P0001 , \wishbone_bd_ram_mem3_reg[164][27]/P0001 , \wishbone_bd_ram_mem3_reg[164][28]/P0001 , \wishbone_bd_ram_mem3_reg[164][29]/P0001 , \wishbone_bd_ram_mem3_reg[164][30]/P0001 , \wishbone_bd_ram_mem3_reg[164][31]/P0001 , \wishbone_bd_ram_mem3_reg[165][24]/P0001 , \wishbone_bd_ram_mem3_reg[165][25]/P0001 , \wishbone_bd_ram_mem3_reg[165][26]/P0001 , \wishbone_bd_ram_mem3_reg[165][27]/P0001 , \wishbone_bd_ram_mem3_reg[165][28]/P0001 , \wishbone_bd_ram_mem3_reg[165][29]/P0001 , \wishbone_bd_ram_mem3_reg[165][30]/P0001 , \wishbone_bd_ram_mem3_reg[165][31]/P0001 , \wishbone_bd_ram_mem3_reg[166][24]/P0001 , \wishbone_bd_ram_mem3_reg[166][25]/P0001 , \wishbone_bd_ram_mem3_reg[166][26]/P0001 , \wishbone_bd_ram_mem3_reg[166][27]/P0001 , \wishbone_bd_ram_mem3_reg[166][28]/P0001 , \wishbone_bd_ram_mem3_reg[166][29]/P0001 , \wishbone_bd_ram_mem3_reg[166][30]/P0001 , \wishbone_bd_ram_mem3_reg[166][31]/P0001 , \wishbone_bd_ram_mem3_reg[167][24]/P0001 , \wishbone_bd_ram_mem3_reg[167][25]/P0001 , \wishbone_bd_ram_mem3_reg[167][26]/P0001 , \wishbone_bd_ram_mem3_reg[167][27]/P0001 , \wishbone_bd_ram_mem3_reg[167][28]/P0001 , \wishbone_bd_ram_mem3_reg[167][29]/P0001 , \wishbone_bd_ram_mem3_reg[167][30]/P0001 , \wishbone_bd_ram_mem3_reg[167][31]/P0001 , \wishbone_bd_ram_mem3_reg[168][24]/P0001 , \wishbone_bd_ram_mem3_reg[168][25]/P0001 , \wishbone_bd_ram_mem3_reg[168][26]/P0001 , \wishbone_bd_ram_mem3_reg[168][27]/P0001 , \wishbone_bd_ram_mem3_reg[168][28]/P0001 , \wishbone_bd_ram_mem3_reg[168][29]/P0001 , \wishbone_bd_ram_mem3_reg[168][30]/P0001 , \wishbone_bd_ram_mem3_reg[168][31]/P0001 , \wishbone_bd_ram_mem3_reg[169][24]/P0001 , \wishbone_bd_ram_mem3_reg[169][25]/P0001 , \wishbone_bd_ram_mem3_reg[169][26]/P0001 , \wishbone_bd_ram_mem3_reg[169][27]/P0001 , \wishbone_bd_ram_mem3_reg[169][28]/P0001 , \wishbone_bd_ram_mem3_reg[169][29]/P0001 , \wishbone_bd_ram_mem3_reg[169][30]/P0001 , \wishbone_bd_ram_mem3_reg[169][31]/P0001 , \wishbone_bd_ram_mem3_reg[16][24]/P0001 , \wishbone_bd_ram_mem3_reg[16][25]/P0001 , \wishbone_bd_ram_mem3_reg[16][26]/P0001 , \wishbone_bd_ram_mem3_reg[16][27]/P0001 , \wishbone_bd_ram_mem3_reg[16][28]/P0001 , \wishbone_bd_ram_mem3_reg[16][29]/P0001 , \wishbone_bd_ram_mem3_reg[16][30]/P0001 , \wishbone_bd_ram_mem3_reg[16][31]/P0001 , \wishbone_bd_ram_mem3_reg[170][24]/P0001 , \wishbone_bd_ram_mem3_reg[170][25]/P0001 , \wishbone_bd_ram_mem3_reg[170][26]/P0001 , \wishbone_bd_ram_mem3_reg[170][27]/P0001 , \wishbone_bd_ram_mem3_reg[170][28]/P0001 , \wishbone_bd_ram_mem3_reg[170][29]/P0001 , \wishbone_bd_ram_mem3_reg[170][30]/P0001 , \wishbone_bd_ram_mem3_reg[170][31]/P0001 , \wishbone_bd_ram_mem3_reg[171][24]/P0001 , \wishbone_bd_ram_mem3_reg[171][25]/P0001 , \wishbone_bd_ram_mem3_reg[171][26]/P0001 , \wishbone_bd_ram_mem3_reg[171][27]/P0001 , \wishbone_bd_ram_mem3_reg[171][28]/P0001 , \wishbone_bd_ram_mem3_reg[171][29]/P0001 , \wishbone_bd_ram_mem3_reg[171][30]/P0001 , \wishbone_bd_ram_mem3_reg[171][31]/P0001 , \wishbone_bd_ram_mem3_reg[172][24]/P0001 , \wishbone_bd_ram_mem3_reg[172][25]/P0001 , \wishbone_bd_ram_mem3_reg[172][26]/P0001 , \wishbone_bd_ram_mem3_reg[172][27]/P0001 , \wishbone_bd_ram_mem3_reg[172][28]/P0001 , \wishbone_bd_ram_mem3_reg[172][29]/P0001 , \wishbone_bd_ram_mem3_reg[172][30]/P0001 , \wishbone_bd_ram_mem3_reg[172][31]/P0001 , \wishbone_bd_ram_mem3_reg[173][24]/P0001 , \wishbone_bd_ram_mem3_reg[173][25]/P0001 , \wishbone_bd_ram_mem3_reg[173][26]/P0001 , \wishbone_bd_ram_mem3_reg[173][27]/P0001 , \wishbone_bd_ram_mem3_reg[173][28]/P0001 , \wishbone_bd_ram_mem3_reg[173][29]/P0001 , \wishbone_bd_ram_mem3_reg[173][30]/P0001 , \wishbone_bd_ram_mem3_reg[173][31]/P0001 , \wishbone_bd_ram_mem3_reg[174][24]/P0001 , \wishbone_bd_ram_mem3_reg[174][25]/P0001 , \wishbone_bd_ram_mem3_reg[174][26]/P0001 , \wishbone_bd_ram_mem3_reg[174][27]/P0001 , \wishbone_bd_ram_mem3_reg[174][28]/P0001 , \wishbone_bd_ram_mem3_reg[174][29]/P0001 , \wishbone_bd_ram_mem3_reg[174][30]/P0001 , \wishbone_bd_ram_mem3_reg[174][31]/P0001 , \wishbone_bd_ram_mem3_reg[175][24]/P0001 , \wishbone_bd_ram_mem3_reg[175][25]/P0001 , \wishbone_bd_ram_mem3_reg[175][26]/P0001 , \wishbone_bd_ram_mem3_reg[175][27]/P0001 , \wishbone_bd_ram_mem3_reg[175][28]/P0001 , \wishbone_bd_ram_mem3_reg[175][29]/P0001 , \wishbone_bd_ram_mem3_reg[175][30]/P0001 , \wishbone_bd_ram_mem3_reg[175][31]/P0001 , \wishbone_bd_ram_mem3_reg[176][24]/P0001 , \wishbone_bd_ram_mem3_reg[176][25]/P0001 , \wishbone_bd_ram_mem3_reg[176][26]/P0001 , \wishbone_bd_ram_mem3_reg[176][27]/P0001 , \wishbone_bd_ram_mem3_reg[176][28]/P0001 , \wishbone_bd_ram_mem3_reg[176][29]/P0001 , \wishbone_bd_ram_mem3_reg[176][30]/P0001 , \wishbone_bd_ram_mem3_reg[176][31]/P0001 , \wishbone_bd_ram_mem3_reg[177][24]/P0001 , \wishbone_bd_ram_mem3_reg[177][25]/P0001 , \wishbone_bd_ram_mem3_reg[177][26]/P0001 , \wishbone_bd_ram_mem3_reg[177][27]/P0001 , \wishbone_bd_ram_mem3_reg[177][28]/P0001 , \wishbone_bd_ram_mem3_reg[177][29]/P0001 , \wishbone_bd_ram_mem3_reg[177][30]/P0001 , \wishbone_bd_ram_mem3_reg[177][31]/P0001 , \wishbone_bd_ram_mem3_reg[178][24]/P0001 , \wishbone_bd_ram_mem3_reg[178][25]/P0001 , \wishbone_bd_ram_mem3_reg[178][26]/P0001 , \wishbone_bd_ram_mem3_reg[178][27]/P0001 , \wishbone_bd_ram_mem3_reg[178][28]/P0001 , \wishbone_bd_ram_mem3_reg[178][29]/P0001 , \wishbone_bd_ram_mem3_reg[178][30]/P0001 , \wishbone_bd_ram_mem3_reg[178][31]/P0001 , \wishbone_bd_ram_mem3_reg[179][24]/P0001 , \wishbone_bd_ram_mem3_reg[179][25]/P0001 , \wishbone_bd_ram_mem3_reg[179][26]/P0001 , \wishbone_bd_ram_mem3_reg[179][27]/P0001 , \wishbone_bd_ram_mem3_reg[179][28]/P0001 , \wishbone_bd_ram_mem3_reg[179][29]/P0001 , \wishbone_bd_ram_mem3_reg[179][30]/P0001 , \wishbone_bd_ram_mem3_reg[179][31]/P0001 , \wishbone_bd_ram_mem3_reg[17][24]/P0001 , \wishbone_bd_ram_mem3_reg[17][25]/P0001 , \wishbone_bd_ram_mem3_reg[17][26]/P0001 , \wishbone_bd_ram_mem3_reg[17][27]/P0001 , \wishbone_bd_ram_mem3_reg[17][28]/P0001 , \wishbone_bd_ram_mem3_reg[17][29]/P0001 , \wishbone_bd_ram_mem3_reg[17][30]/P0001 , \wishbone_bd_ram_mem3_reg[17][31]/P0001 , \wishbone_bd_ram_mem3_reg[180][24]/P0001 , \wishbone_bd_ram_mem3_reg[180][25]/P0001 , \wishbone_bd_ram_mem3_reg[180][26]/P0001 , \wishbone_bd_ram_mem3_reg[180][27]/P0001 , \wishbone_bd_ram_mem3_reg[180][28]/P0001 , \wishbone_bd_ram_mem3_reg[180][29]/P0001 , \wishbone_bd_ram_mem3_reg[180][30]/P0001 , \wishbone_bd_ram_mem3_reg[180][31]/P0001 , \wishbone_bd_ram_mem3_reg[181][24]/P0001 , \wishbone_bd_ram_mem3_reg[181][25]/P0001 , \wishbone_bd_ram_mem3_reg[181][26]/P0001 , \wishbone_bd_ram_mem3_reg[181][27]/P0001 , \wishbone_bd_ram_mem3_reg[181][28]/P0001 , \wishbone_bd_ram_mem3_reg[181][29]/P0001 , \wishbone_bd_ram_mem3_reg[181][30]/P0001 , \wishbone_bd_ram_mem3_reg[181][31]/P0001 , \wishbone_bd_ram_mem3_reg[182][24]/P0001 , \wishbone_bd_ram_mem3_reg[182][25]/P0001 , \wishbone_bd_ram_mem3_reg[182][26]/P0001 , \wishbone_bd_ram_mem3_reg[182][27]/P0001 , \wishbone_bd_ram_mem3_reg[182][28]/P0001 , \wishbone_bd_ram_mem3_reg[182][29]/P0001 , \wishbone_bd_ram_mem3_reg[182][30]/P0001 , \wishbone_bd_ram_mem3_reg[182][31]/P0001 , \wishbone_bd_ram_mem3_reg[183][24]/P0001 , \wishbone_bd_ram_mem3_reg[183][25]/P0001 , \wishbone_bd_ram_mem3_reg[183][26]/P0001 , \wishbone_bd_ram_mem3_reg[183][27]/P0001 , \wishbone_bd_ram_mem3_reg[183][28]/P0001 , \wishbone_bd_ram_mem3_reg[183][29]/P0001 , \wishbone_bd_ram_mem3_reg[183][30]/P0001 , \wishbone_bd_ram_mem3_reg[183][31]/P0001 , \wishbone_bd_ram_mem3_reg[184][24]/P0001 , \wishbone_bd_ram_mem3_reg[184][25]/P0001 , \wishbone_bd_ram_mem3_reg[184][26]/P0001 , \wishbone_bd_ram_mem3_reg[184][27]/P0001 , \wishbone_bd_ram_mem3_reg[184][28]/P0001 , \wishbone_bd_ram_mem3_reg[184][29]/P0001 , \wishbone_bd_ram_mem3_reg[184][30]/P0001 , \wishbone_bd_ram_mem3_reg[184][31]/P0001 , \wishbone_bd_ram_mem3_reg[185][24]/P0001 , \wishbone_bd_ram_mem3_reg[185][25]/P0001 , \wishbone_bd_ram_mem3_reg[185][26]/P0001 , \wishbone_bd_ram_mem3_reg[185][27]/P0001 , \wishbone_bd_ram_mem3_reg[185][28]/P0001 , \wishbone_bd_ram_mem3_reg[185][29]/P0001 , \wishbone_bd_ram_mem3_reg[185][30]/P0001 , \wishbone_bd_ram_mem3_reg[185][31]/P0001 , \wishbone_bd_ram_mem3_reg[186][24]/P0001 , \wishbone_bd_ram_mem3_reg[186][25]/P0001 , \wishbone_bd_ram_mem3_reg[186][26]/P0001 , \wishbone_bd_ram_mem3_reg[186][27]/P0001 , \wishbone_bd_ram_mem3_reg[186][28]/P0001 , \wishbone_bd_ram_mem3_reg[186][29]/P0001 , \wishbone_bd_ram_mem3_reg[186][30]/P0001 , \wishbone_bd_ram_mem3_reg[186][31]/P0001 , \wishbone_bd_ram_mem3_reg[187][24]/P0001 , \wishbone_bd_ram_mem3_reg[187][25]/P0001 , \wishbone_bd_ram_mem3_reg[187][26]/P0001 , \wishbone_bd_ram_mem3_reg[187][27]/P0001 , \wishbone_bd_ram_mem3_reg[187][28]/P0001 , \wishbone_bd_ram_mem3_reg[187][29]/P0001 , \wishbone_bd_ram_mem3_reg[187][30]/P0001 , \wishbone_bd_ram_mem3_reg[187][31]/P0001 , \wishbone_bd_ram_mem3_reg[188][24]/P0001 , \wishbone_bd_ram_mem3_reg[188][25]/P0001 , \wishbone_bd_ram_mem3_reg[188][26]/P0001 , \wishbone_bd_ram_mem3_reg[188][27]/P0001 , \wishbone_bd_ram_mem3_reg[188][28]/P0001 , \wishbone_bd_ram_mem3_reg[188][29]/P0001 , \wishbone_bd_ram_mem3_reg[188][30]/P0001 , \wishbone_bd_ram_mem3_reg[188][31]/P0001 , \wishbone_bd_ram_mem3_reg[189][24]/P0001 , \wishbone_bd_ram_mem3_reg[189][25]/P0001 , \wishbone_bd_ram_mem3_reg[189][26]/P0001 , \wishbone_bd_ram_mem3_reg[189][27]/P0001 , \wishbone_bd_ram_mem3_reg[189][28]/P0001 , \wishbone_bd_ram_mem3_reg[189][29]/P0001 , \wishbone_bd_ram_mem3_reg[189][30]/P0001 , \wishbone_bd_ram_mem3_reg[189][31]/P0001 , \wishbone_bd_ram_mem3_reg[18][24]/P0001 , \wishbone_bd_ram_mem3_reg[18][25]/P0001 , \wishbone_bd_ram_mem3_reg[18][26]/P0001 , \wishbone_bd_ram_mem3_reg[18][27]/P0001 , \wishbone_bd_ram_mem3_reg[18][28]/P0001 , \wishbone_bd_ram_mem3_reg[18][29]/P0001 , \wishbone_bd_ram_mem3_reg[18][30]/P0001 , \wishbone_bd_ram_mem3_reg[18][31]/P0001 , \wishbone_bd_ram_mem3_reg[190][24]/P0001 , \wishbone_bd_ram_mem3_reg[190][25]/P0001 , \wishbone_bd_ram_mem3_reg[190][26]/P0001 , \wishbone_bd_ram_mem3_reg[190][27]/P0001 , \wishbone_bd_ram_mem3_reg[190][28]/P0001 , \wishbone_bd_ram_mem3_reg[190][29]/P0001 , \wishbone_bd_ram_mem3_reg[190][30]/P0001 , \wishbone_bd_ram_mem3_reg[190][31]/P0001 , \wishbone_bd_ram_mem3_reg[191][24]/P0001 , \wishbone_bd_ram_mem3_reg[191][25]/P0001 , \wishbone_bd_ram_mem3_reg[191][26]/P0001 , \wishbone_bd_ram_mem3_reg[191][27]/P0001 , \wishbone_bd_ram_mem3_reg[191][28]/P0001 , \wishbone_bd_ram_mem3_reg[191][29]/P0001 , \wishbone_bd_ram_mem3_reg[191][30]/P0001 , \wishbone_bd_ram_mem3_reg[191][31]/P0001 , \wishbone_bd_ram_mem3_reg[192][24]/P0001 , \wishbone_bd_ram_mem3_reg[192][25]/P0001 , \wishbone_bd_ram_mem3_reg[192][26]/P0001 , \wishbone_bd_ram_mem3_reg[192][27]/P0001 , \wishbone_bd_ram_mem3_reg[192][28]/P0001 , \wishbone_bd_ram_mem3_reg[192][29]/P0001 , \wishbone_bd_ram_mem3_reg[192][30]/P0001 , \wishbone_bd_ram_mem3_reg[192][31]/P0001 , \wishbone_bd_ram_mem3_reg[193][24]/P0001 , \wishbone_bd_ram_mem3_reg[193][25]/P0001 , \wishbone_bd_ram_mem3_reg[193][26]/P0001 , \wishbone_bd_ram_mem3_reg[193][27]/P0001 , \wishbone_bd_ram_mem3_reg[193][28]/P0001 , \wishbone_bd_ram_mem3_reg[193][29]/P0001 , \wishbone_bd_ram_mem3_reg[193][30]/P0001 , \wishbone_bd_ram_mem3_reg[193][31]/P0001 , \wishbone_bd_ram_mem3_reg[194][24]/P0001 , \wishbone_bd_ram_mem3_reg[194][25]/P0001 , \wishbone_bd_ram_mem3_reg[194][26]/P0001 , \wishbone_bd_ram_mem3_reg[194][27]/P0001 , \wishbone_bd_ram_mem3_reg[194][28]/P0001 , \wishbone_bd_ram_mem3_reg[194][29]/P0001 , \wishbone_bd_ram_mem3_reg[194][30]/P0001 , \wishbone_bd_ram_mem3_reg[194][31]/P0001 , \wishbone_bd_ram_mem3_reg[195][24]/P0001 , \wishbone_bd_ram_mem3_reg[195][25]/P0001 , \wishbone_bd_ram_mem3_reg[195][26]/P0001 , \wishbone_bd_ram_mem3_reg[195][27]/P0001 , \wishbone_bd_ram_mem3_reg[195][28]/P0001 , \wishbone_bd_ram_mem3_reg[195][29]/P0001 , \wishbone_bd_ram_mem3_reg[195][30]/P0001 , \wishbone_bd_ram_mem3_reg[195][31]/P0001 , \wishbone_bd_ram_mem3_reg[196][24]/P0001 , \wishbone_bd_ram_mem3_reg[196][25]/P0001 , \wishbone_bd_ram_mem3_reg[196][26]/P0001 , \wishbone_bd_ram_mem3_reg[196][27]/P0001 , \wishbone_bd_ram_mem3_reg[196][28]/P0001 , \wishbone_bd_ram_mem3_reg[196][29]/P0001 , \wishbone_bd_ram_mem3_reg[196][30]/P0001 , \wishbone_bd_ram_mem3_reg[196][31]/P0001 , \wishbone_bd_ram_mem3_reg[197][24]/P0001 , \wishbone_bd_ram_mem3_reg[197][25]/P0001 , \wishbone_bd_ram_mem3_reg[197][26]/P0001 , \wishbone_bd_ram_mem3_reg[197][27]/P0001 , \wishbone_bd_ram_mem3_reg[197][28]/P0001 , \wishbone_bd_ram_mem3_reg[197][29]/P0001 , \wishbone_bd_ram_mem3_reg[197][30]/P0001 , \wishbone_bd_ram_mem3_reg[197][31]/P0001 , \wishbone_bd_ram_mem3_reg[198][24]/P0001 , \wishbone_bd_ram_mem3_reg[198][25]/P0001 , \wishbone_bd_ram_mem3_reg[198][26]/P0001 , \wishbone_bd_ram_mem3_reg[198][27]/P0001 , \wishbone_bd_ram_mem3_reg[198][28]/P0001 , \wishbone_bd_ram_mem3_reg[198][29]/P0001 , \wishbone_bd_ram_mem3_reg[198][30]/P0001 , \wishbone_bd_ram_mem3_reg[198][31]/P0001 , \wishbone_bd_ram_mem3_reg[199][24]/P0001 , \wishbone_bd_ram_mem3_reg[199][25]/P0001 , \wishbone_bd_ram_mem3_reg[199][26]/P0001 , \wishbone_bd_ram_mem3_reg[199][27]/P0001 , \wishbone_bd_ram_mem3_reg[199][28]/P0001 , \wishbone_bd_ram_mem3_reg[199][29]/P0001 , \wishbone_bd_ram_mem3_reg[199][30]/P0001 , \wishbone_bd_ram_mem3_reg[199][31]/P0001 , \wishbone_bd_ram_mem3_reg[19][24]/P0001 , \wishbone_bd_ram_mem3_reg[19][25]/P0001 , \wishbone_bd_ram_mem3_reg[19][26]/P0001 , \wishbone_bd_ram_mem3_reg[19][27]/P0001 , \wishbone_bd_ram_mem3_reg[19][28]/P0001 , \wishbone_bd_ram_mem3_reg[19][29]/P0001 , \wishbone_bd_ram_mem3_reg[19][30]/P0001 , \wishbone_bd_ram_mem3_reg[19][31]/P0001 , \wishbone_bd_ram_mem3_reg[1][24]/P0001 , \wishbone_bd_ram_mem3_reg[1][25]/P0001 , \wishbone_bd_ram_mem3_reg[1][26]/P0001 , \wishbone_bd_ram_mem3_reg[1][27]/P0001 , \wishbone_bd_ram_mem3_reg[1][28]/P0001 , \wishbone_bd_ram_mem3_reg[1][29]/P0001 , \wishbone_bd_ram_mem3_reg[1][30]/P0001 , \wishbone_bd_ram_mem3_reg[1][31]/P0001 , \wishbone_bd_ram_mem3_reg[200][24]/P0001 , \wishbone_bd_ram_mem3_reg[200][25]/P0001 , \wishbone_bd_ram_mem3_reg[200][26]/P0001 , \wishbone_bd_ram_mem3_reg[200][27]/P0001 , \wishbone_bd_ram_mem3_reg[200][28]/P0001 , \wishbone_bd_ram_mem3_reg[200][29]/P0001 , \wishbone_bd_ram_mem3_reg[200][30]/P0001 , \wishbone_bd_ram_mem3_reg[200][31]/P0001 , \wishbone_bd_ram_mem3_reg[201][24]/P0001 , \wishbone_bd_ram_mem3_reg[201][25]/P0001 , \wishbone_bd_ram_mem3_reg[201][26]/P0001 , \wishbone_bd_ram_mem3_reg[201][27]/P0001 , \wishbone_bd_ram_mem3_reg[201][28]/P0001 , \wishbone_bd_ram_mem3_reg[201][29]/P0001 , \wishbone_bd_ram_mem3_reg[201][30]/P0001 , \wishbone_bd_ram_mem3_reg[201][31]/P0001 , \wishbone_bd_ram_mem3_reg[202][24]/P0001 , \wishbone_bd_ram_mem3_reg[202][25]/P0001 , \wishbone_bd_ram_mem3_reg[202][26]/P0001 , \wishbone_bd_ram_mem3_reg[202][27]/P0001 , \wishbone_bd_ram_mem3_reg[202][28]/P0001 , \wishbone_bd_ram_mem3_reg[202][29]/P0001 , \wishbone_bd_ram_mem3_reg[202][30]/P0001 , \wishbone_bd_ram_mem3_reg[202][31]/P0001 , \wishbone_bd_ram_mem3_reg[203][24]/P0001 , \wishbone_bd_ram_mem3_reg[203][25]/P0001 , \wishbone_bd_ram_mem3_reg[203][26]/P0001 , \wishbone_bd_ram_mem3_reg[203][27]/P0001 , \wishbone_bd_ram_mem3_reg[203][28]/P0001 , \wishbone_bd_ram_mem3_reg[203][29]/P0001 , \wishbone_bd_ram_mem3_reg[203][30]/P0001 , \wishbone_bd_ram_mem3_reg[203][31]/P0001 , \wishbone_bd_ram_mem3_reg[204][24]/P0001 , \wishbone_bd_ram_mem3_reg[204][25]/P0001 , \wishbone_bd_ram_mem3_reg[204][26]/P0001 , \wishbone_bd_ram_mem3_reg[204][27]/P0001 , \wishbone_bd_ram_mem3_reg[204][28]/P0001 , \wishbone_bd_ram_mem3_reg[204][29]/P0001 , \wishbone_bd_ram_mem3_reg[204][30]/P0001 , \wishbone_bd_ram_mem3_reg[204][31]/P0001 , \wishbone_bd_ram_mem3_reg[205][24]/P0001 , \wishbone_bd_ram_mem3_reg[205][25]/P0001 , \wishbone_bd_ram_mem3_reg[205][26]/P0001 , \wishbone_bd_ram_mem3_reg[205][27]/P0001 , \wishbone_bd_ram_mem3_reg[205][28]/P0001 , \wishbone_bd_ram_mem3_reg[205][29]/P0001 , \wishbone_bd_ram_mem3_reg[205][30]/P0001 , \wishbone_bd_ram_mem3_reg[205][31]/P0001 , \wishbone_bd_ram_mem3_reg[206][24]/P0001 , \wishbone_bd_ram_mem3_reg[206][25]/P0001 , \wishbone_bd_ram_mem3_reg[206][26]/P0001 , \wishbone_bd_ram_mem3_reg[206][27]/P0001 , \wishbone_bd_ram_mem3_reg[206][28]/P0001 , \wishbone_bd_ram_mem3_reg[206][29]/P0001 , \wishbone_bd_ram_mem3_reg[206][30]/P0001 , \wishbone_bd_ram_mem3_reg[206][31]/P0001 , \wishbone_bd_ram_mem3_reg[207][24]/P0001 , \wishbone_bd_ram_mem3_reg[207][25]/P0001 , \wishbone_bd_ram_mem3_reg[207][26]/P0001 , \wishbone_bd_ram_mem3_reg[207][27]/P0001 , \wishbone_bd_ram_mem3_reg[207][28]/P0001 , \wishbone_bd_ram_mem3_reg[207][29]/P0001 , \wishbone_bd_ram_mem3_reg[207][30]/P0001 , \wishbone_bd_ram_mem3_reg[207][31]/P0001 , \wishbone_bd_ram_mem3_reg[208][24]/P0001 , \wishbone_bd_ram_mem3_reg[208][25]/P0001 , \wishbone_bd_ram_mem3_reg[208][26]/P0001 , \wishbone_bd_ram_mem3_reg[208][27]/P0001 , \wishbone_bd_ram_mem3_reg[208][28]/P0001 , \wishbone_bd_ram_mem3_reg[208][29]/P0001 , \wishbone_bd_ram_mem3_reg[208][30]/P0001 , \wishbone_bd_ram_mem3_reg[208][31]/P0001 , \wishbone_bd_ram_mem3_reg[209][24]/P0001 , \wishbone_bd_ram_mem3_reg[209][25]/P0001 , \wishbone_bd_ram_mem3_reg[209][26]/P0001 , \wishbone_bd_ram_mem3_reg[209][27]/P0001 , \wishbone_bd_ram_mem3_reg[209][28]/P0001 , \wishbone_bd_ram_mem3_reg[209][29]/P0001 , \wishbone_bd_ram_mem3_reg[209][30]/P0001 , \wishbone_bd_ram_mem3_reg[209][31]/P0001 , \wishbone_bd_ram_mem3_reg[20][24]/P0001 , \wishbone_bd_ram_mem3_reg[20][25]/P0001 , \wishbone_bd_ram_mem3_reg[20][26]/P0001 , \wishbone_bd_ram_mem3_reg[20][27]/P0001 , \wishbone_bd_ram_mem3_reg[20][28]/P0001 , \wishbone_bd_ram_mem3_reg[20][29]/P0001 , \wishbone_bd_ram_mem3_reg[20][30]/P0001 , \wishbone_bd_ram_mem3_reg[20][31]/P0001 , \wishbone_bd_ram_mem3_reg[210][24]/P0001 , \wishbone_bd_ram_mem3_reg[210][25]/P0001 , \wishbone_bd_ram_mem3_reg[210][26]/P0001 , \wishbone_bd_ram_mem3_reg[210][27]/P0001 , \wishbone_bd_ram_mem3_reg[210][28]/P0001 , \wishbone_bd_ram_mem3_reg[210][29]/P0001 , \wishbone_bd_ram_mem3_reg[210][30]/P0001 , \wishbone_bd_ram_mem3_reg[210][31]/P0001 , \wishbone_bd_ram_mem3_reg[211][24]/P0001 , \wishbone_bd_ram_mem3_reg[211][25]/P0001 , \wishbone_bd_ram_mem3_reg[211][26]/P0001 , \wishbone_bd_ram_mem3_reg[211][27]/P0001 , \wishbone_bd_ram_mem3_reg[211][28]/P0001 , \wishbone_bd_ram_mem3_reg[211][29]/P0001 , \wishbone_bd_ram_mem3_reg[211][30]/P0001 , \wishbone_bd_ram_mem3_reg[211][31]/P0001 , \wishbone_bd_ram_mem3_reg[212][24]/P0001 , \wishbone_bd_ram_mem3_reg[212][25]/P0001 , \wishbone_bd_ram_mem3_reg[212][26]/P0001 , \wishbone_bd_ram_mem3_reg[212][27]/P0001 , \wishbone_bd_ram_mem3_reg[212][28]/P0001 , \wishbone_bd_ram_mem3_reg[212][29]/P0001 , \wishbone_bd_ram_mem3_reg[212][30]/P0001 , \wishbone_bd_ram_mem3_reg[212][31]/P0001 , \wishbone_bd_ram_mem3_reg[213][24]/P0001 , \wishbone_bd_ram_mem3_reg[213][25]/P0001 , \wishbone_bd_ram_mem3_reg[213][26]/P0001 , \wishbone_bd_ram_mem3_reg[213][27]/P0001 , \wishbone_bd_ram_mem3_reg[213][28]/P0001 , \wishbone_bd_ram_mem3_reg[213][29]/P0001 , \wishbone_bd_ram_mem3_reg[213][30]/P0001 , \wishbone_bd_ram_mem3_reg[213][31]/P0001 , \wishbone_bd_ram_mem3_reg[214][24]/P0001 , \wishbone_bd_ram_mem3_reg[214][25]/P0001 , \wishbone_bd_ram_mem3_reg[214][26]/P0001 , \wishbone_bd_ram_mem3_reg[214][27]/P0001 , \wishbone_bd_ram_mem3_reg[214][28]/P0001 , \wishbone_bd_ram_mem3_reg[214][29]/P0001 , \wishbone_bd_ram_mem3_reg[214][30]/P0001 , \wishbone_bd_ram_mem3_reg[214][31]/P0001 , \wishbone_bd_ram_mem3_reg[215][24]/P0001 , \wishbone_bd_ram_mem3_reg[215][25]/P0001 , \wishbone_bd_ram_mem3_reg[215][26]/P0001 , \wishbone_bd_ram_mem3_reg[215][27]/P0001 , \wishbone_bd_ram_mem3_reg[215][28]/P0001 , \wishbone_bd_ram_mem3_reg[215][29]/P0001 , \wishbone_bd_ram_mem3_reg[215][30]/P0001 , \wishbone_bd_ram_mem3_reg[215][31]/P0001 , \wishbone_bd_ram_mem3_reg[216][24]/P0001 , \wishbone_bd_ram_mem3_reg[216][25]/P0001 , \wishbone_bd_ram_mem3_reg[216][26]/P0001 , \wishbone_bd_ram_mem3_reg[216][27]/P0001 , \wishbone_bd_ram_mem3_reg[216][28]/P0001 , \wishbone_bd_ram_mem3_reg[216][29]/P0001 , \wishbone_bd_ram_mem3_reg[216][30]/P0001 , \wishbone_bd_ram_mem3_reg[216][31]/P0001 , \wishbone_bd_ram_mem3_reg[217][24]/P0001 , \wishbone_bd_ram_mem3_reg[217][25]/P0001 , \wishbone_bd_ram_mem3_reg[217][26]/P0001 , \wishbone_bd_ram_mem3_reg[217][27]/P0001 , \wishbone_bd_ram_mem3_reg[217][28]/P0001 , \wishbone_bd_ram_mem3_reg[217][29]/P0001 , \wishbone_bd_ram_mem3_reg[217][30]/P0001 , \wishbone_bd_ram_mem3_reg[217][31]/P0001 , \wishbone_bd_ram_mem3_reg[218][24]/P0001 , \wishbone_bd_ram_mem3_reg[218][25]/P0001 , \wishbone_bd_ram_mem3_reg[218][26]/P0001 , \wishbone_bd_ram_mem3_reg[218][27]/P0001 , \wishbone_bd_ram_mem3_reg[218][28]/P0001 , \wishbone_bd_ram_mem3_reg[218][29]/P0001 , \wishbone_bd_ram_mem3_reg[218][30]/P0001 , \wishbone_bd_ram_mem3_reg[218][31]/P0001 , \wishbone_bd_ram_mem3_reg[219][24]/P0001 , \wishbone_bd_ram_mem3_reg[219][25]/P0001 , \wishbone_bd_ram_mem3_reg[219][26]/P0001 , \wishbone_bd_ram_mem3_reg[219][27]/P0001 , \wishbone_bd_ram_mem3_reg[219][28]/P0001 , \wishbone_bd_ram_mem3_reg[219][29]/P0001 , \wishbone_bd_ram_mem3_reg[219][30]/P0001 , \wishbone_bd_ram_mem3_reg[219][31]/P0001 , \wishbone_bd_ram_mem3_reg[21][24]/P0001 , \wishbone_bd_ram_mem3_reg[21][25]/P0001 , \wishbone_bd_ram_mem3_reg[21][26]/P0001 , \wishbone_bd_ram_mem3_reg[21][27]/P0001 , \wishbone_bd_ram_mem3_reg[21][28]/P0001 , \wishbone_bd_ram_mem3_reg[21][29]/P0001 , \wishbone_bd_ram_mem3_reg[21][30]/P0001 , \wishbone_bd_ram_mem3_reg[21][31]/P0001 , \wishbone_bd_ram_mem3_reg[220][24]/P0001 , \wishbone_bd_ram_mem3_reg[220][25]/P0001 , \wishbone_bd_ram_mem3_reg[220][26]/P0001 , \wishbone_bd_ram_mem3_reg[220][27]/P0001 , \wishbone_bd_ram_mem3_reg[220][28]/P0001 , \wishbone_bd_ram_mem3_reg[220][29]/P0001 , \wishbone_bd_ram_mem3_reg[220][30]/P0001 , \wishbone_bd_ram_mem3_reg[220][31]/P0001 , \wishbone_bd_ram_mem3_reg[221][24]/P0001 , \wishbone_bd_ram_mem3_reg[221][25]/P0001 , \wishbone_bd_ram_mem3_reg[221][26]/P0001 , \wishbone_bd_ram_mem3_reg[221][27]/P0001 , \wishbone_bd_ram_mem3_reg[221][28]/P0001 , \wishbone_bd_ram_mem3_reg[221][29]/P0001 , \wishbone_bd_ram_mem3_reg[221][30]/P0001 , \wishbone_bd_ram_mem3_reg[221][31]/P0001 , \wishbone_bd_ram_mem3_reg[222][24]/P0001 , \wishbone_bd_ram_mem3_reg[222][25]/P0001 , \wishbone_bd_ram_mem3_reg[222][26]/P0001 , \wishbone_bd_ram_mem3_reg[222][27]/P0001 , \wishbone_bd_ram_mem3_reg[222][28]/P0001 , \wishbone_bd_ram_mem3_reg[222][29]/P0001 , \wishbone_bd_ram_mem3_reg[222][30]/P0001 , \wishbone_bd_ram_mem3_reg[222][31]/P0001 , \wishbone_bd_ram_mem3_reg[223][24]/P0001 , \wishbone_bd_ram_mem3_reg[223][25]/P0001 , \wishbone_bd_ram_mem3_reg[223][26]/P0001 , \wishbone_bd_ram_mem3_reg[223][27]/P0001 , \wishbone_bd_ram_mem3_reg[223][28]/P0001 , \wishbone_bd_ram_mem3_reg[223][29]/P0001 , \wishbone_bd_ram_mem3_reg[223][30]/P0001 , \wishbone_bd_ram_mem3_reg[223][31]/P0001 , \wishbone_bd_ram_mem3_reg[224][24]/P0001 , \wishbone_bd_ram_mem3_reg[224][25]/P0001 , \wishbone_bd_ram_mem3_reg[224][26]/P0001 , \wishbone_bd_ram_mem3_reg[224][27]/P0001 , \wishbone_bd_ram_mem3_reg[224][28]/P0001 , \wishbone_bd_ram_mem3_reg[224][29]/P0001 , \wishbone_bd_ram_mem3_reg[224][30]/P0001 , \wishbone_bd_ram_mem3_reg[224][31]/P0001 , \wishbone_bd_ram_mem3_reg[225][24]/P0001 , \wishbone_bd_ram_mem3_reg[225][25]/P0001 , \wishbone_bd_ram_mem3_reg[225][26]/P0001 , \wishbone_bd_ram_mem3_reg[225][27]/P0001 , \wishbone_bd_ram_mem3_reg[225][28]/P0001 , \wishbone_bd_ram_mem3_reg[225][29]/P0001 , \wishbone_bd_ram_mem3_reg[225][30]/P0001 , \wishbone_bd_ram_mem3_reg[225][31]/P0001 , \wishbone_bd_ram_mem3_reg[226][24]/P0001 , \wishbone_bd_ram_mem3_reg[226][25]/P0001 , \wishbone_bd_ram_mem3_reg[226][26]/P0001 , \wishbone_bd_ram_mem3_reg[226][27]/P0001 , \wishbone_bd_ram_mem3_reg[226][28]/P0001 , \wishbone_bd_ram_mem3_reg[226][29]/P0001 , \wishbone_bd_ram_mem3_reg[226][30]/P0001 , \wishbone_bd_ram_mem3_reg[226][31]/P0001 , \wishbone_bd_ram_mem3_reg[227][24]/P0001 , \wishbone_bd_ram_mem3_reg[227][25]/P0001 , \wishbone_bd_ram_mem3_reg[227][26]/P0001 , \wishbone_bd_ram_mem3_reg[227][27]/P0001 , \wishbone_bd_ram_mem3_reg[227][28]/P0001 , \wishbone_bd_ram_mem3_reg[227][29]/P0001 , \wishbone_bd_ram_mem3_reg[227][30]/P0001 , \wishbone_bd_ram_mem3_reg[227][31]/P0001 , \wishbone_bd_ram_mem3_reg[228][24]/P0001 , \wishbone_bd_ram_mem3_reg[228][25]/P0001 , \wishbone_bd_ram_mem3_reg[228][26]/P0001 , \wishbone_bd_ram_mem3_reg[228][27]/P0001 , \wishbone_bd_ram_mem3_reg[228][28]/P0001 , \wishbone_bd_ram_mem3_reg[228][29]/P0001 , \wishbone_bd_ram_mem3_reg[228][30]/P0001 , \wishbone_bd_ram_mem3_reg[228][31]/P0001 , \wishbone_bd_ram_mem3_reg[229][24]/P0001 , \wishbone_bd_ram_mem3_reg[229][25]/P0001 , \wishbone_bd_ram_mem3_reg[229][26]/P0001 , \wishbone_bd_ram_mem3_reg[229][27]/P0001 , \wishbone_bd_ram_mem3_reg[229][28]/P0001 , \wishbone_bd_ram_mem3_reg[229][29]/P0001 , \wishbone_bd_ram_mem3_reg[229][30]/P0001 , \wishbone_bd_ram_mem3_reg[229][31]/P0001 , \wishbone_bd_ram_mem3_reg[22][24]/P0001 , \wishbone_bd_ram_mem3_reg[22][25]/P0001 , \wishbone_bd_ram_mem3_reg[22][26]/P0001 , \wishbone_bd_ram_mem3_reg[22][27]/P0001 , \wishbone_bd_ram_mem3_reg[22][28]/P0001 , \wishbone_bd_ram_mem3_reg[22][29]/P0001 , \wishbone_bd_ram_mem3_reg[22][30]/P0001 , \wishbone_bd_ram_mem3_reg[22][31]/P0001 , \wishbone_bd_ram_mem3_reg[230][24]/P0001 , \wishbone_bd_ram_mem3_reg[230][25]/P0001 , \wishbone_bd_ram_mem3_reg[230][26]/P0001 , \wishbone_bd_ram_mem3_reg[230][27]/P0001 , \wishbone_bd_ram_mem3_reg[230][28]/P0001 , \wishbone_bd_ram_mem3_reg[230][29]/P0001 , \wishbone_bd_ram_mem3_reg[230][30]/P0001 , \wishbone_bd_ram_mem3_reg[230][31]/P0001 , \wishbone_bd_ram_mem3_reg[231][24]/P0001 , \wishbone_bd_ram_mem3_reg[231][25]/P0001 , \wishbone_bd_ram_mem3_reg[231][26]/P0001 , \wishbone_bd_ram_mem3_reg[231][27]/P0001 , \wishbone_bd_ram_mem3_reg[231][28]/P0001 , \wishbone_bd_ram_mem3_reg[231][29]/P0001 , \wishbone_bd_ram_mem3_reg[231][30]/P0001 , \wishbone_bd_ram_mem3_reg[231][31]/P0001 , \wishbone_bd_ram_mem3_reg[232][24]/P0001 , \wishbone_bd_ram_mem3_reg[232][25]/P0001 , \wishbone_bd_ram_mem3_reg[232][26]/P0001 , \wishbone_bd_ram_mem3_reg[232][27]/P0001 , \wishbone_bd_ram_mem3_reg[232][28]/P0001 , \wishbone_bd_ram_mem3_reg[232][29]/P0001 , \wishbone_bd_ram_mem3_reg[232][30]/P0001 , \wishbone_bd_ram_mem3_reg[232][31]/P0001 , \wishbone_bd_ram_mem3_reg[233][24]/P0001 , \wishbone_bd_ram_mem3_reg[233][25]/P0001 , \wishbone_bd_ram_mem3_reg[233][26]/P0001 , \wishbone_bd_ram_mem3_reg[233][27]/P0001 , \wishbone_bd_ram_mem3_reg[233][28]/P0001 , \wishbone_bd_ram_mem3_reg[233][29]/P0001 , \wishbone_bd_ram_mem3_reg[233][30]/P0001 , \wishbone_bd_ram_mem3_reg[233][31]/P0001 , \wishbone_bd_ram_mem3_reg[234][24]/P0001 , \wishbone_bd_ram_mem3_reg[234][25]/P0001 , \wishbone_bd_ram_mem3_reg[234][26]/P0001 , \wishbone_bd_ram_mem3_reg[234][27]/P0001 , \wishbone_bd_ram_mem3_reg[234][28]/P0001 , \wishbone_bd_ram_mem3_reg[234][29]/P0001 , \wishbone_bd_ram_mem3_reg[234][30]/P0001 , \wishbone_bd_ram_mem3_reg[234][31]/P0001 , \wishbone_bd_ram_mem3_reg[235][24]/P0001 , \wishbone_bd_ram_mem3_reg[235][25]/P0001 , \wishbone_bd_ram_mem3_reg[235][26]/P0001 , \wishbone_bd_ram_mem3_reg[235][27]/P0001 , \wishbone_bd_ram_mem3_reg[235][28]/P0001 , \wishbone_bd_ram_mem3_reg[235][29]/P0001 , \wishbone_bd_ram_mem3_reg[235][30]/P0001 , \wishbone_bd_ram_mem3_reg[235][31]/P0001 , \wishbone_bd_ram_mem3_reg[236][24]/P0001 , \wishbone_bd_ram_mem3_reg[236][25]/P0001 , \wishbone_bd_ram_mem3_reg[236][26]/P0001 , \wishbone_bd_ram_mem3_reg[236][27]/P0001 , \wishbone_bd_ram_mem3_reg[236][28]/P0001 , \wishbone_bd_ram_mem3_reg[236][29]/P0001 , \wishbone_bd_ram_mem3_reg[236][30]/P0001 , \wishbone_bd_ram_mem3_reg[236][31]/P0001 , \wishbone_bd_ram_mem3_reg[237][24]/P0001 , \wishbone_bd_ram_mem3_reg[237][25]/P0001 , \wishbone_bd_ram_mem3_reg[237][26]/P0001 , \wishbone_bd_ram_mem3_reg[237][27]/P0001 , \wishbone_bd_ram_mem3_reg[237][28]/P0001 , \wishbone_bd_ram_mem3_reg[237][29]/P0001 , \wishbone_bd_ram_mem3_reg[237][30]/P0001 , \wishbone_bd_ram_mem3_reg[237][31]/P0001 , \wishbone_bd_ram_mem3_reg[238][24]/P0001 , \wishbone_bd_ram_mem3_reg[238][25]/P0001 , \wishbone_bd_ram_mem3_reg[238][26]/P0001 , \wishbone_bd_ram_mem3_reg[238][27]/P0001 , \wishbone_bd_ram_mem3_reg[238][28]/P0001 , \wishbone_bd_ram_mem3_reg[238][29]/P0001 , \wishbone_bd_ram_mem3_reg[238][30]/P0001 , \wishbone_bd_ram_mem3_reg[238][31]/P0001 , \wishbone_bd_ram_mem3_reg[239][24]/P0001 , \wishbone_bd_ram_mem3_reg[239][25]/P0001 , \wishbone_bd_ram_mem3_reg[239][26]/P0001 , \wishbone_bd_ram_mem3_reg[239][27]/P0001 , \wishbone_bd_ram_mem3_reg[239][28]/P0001 , \wishbone_bd_ram_mem3_reg[239][29]/P0001 , \wishbone_bd_ram_mem3_reg[239][30]/P0001 , \wishbone_bd_ram_mem3_reg[239][31]/P0001 , \wishbone_bd_ram_mem3_reg[23][24]/P0001 , \wishbone_bd_ram_mem3_reg[23][25]/P0001 , \wishbone_bd_ram_mem3_reg[23][26]/P0001 , \wishbone_bd_ram_mem3_reg[23][27]/P0001 , \wishbone_bd_ram_mem3_reg[23][28]/P0001 , \wishbone_bd_ram_mem3_reg[23][29]/P0001 , \wishbone_bd_ram_mem3_reg[23][30]/P0001 , \wishbone_bd_ram_mem3_reg[23][31]/P0001 , \wishbone_bd_ram_mem3_reg[240][24]/P0001 , \wishbone_bd_ram_mem3_reg[240][25]/P0001 , \wishbone_bd_ram_mem3_reg[240][26]/P0001 , \wishbone_bd_ram_mem3_reg[240][27]/P0001 , \wishbone_bd_ram_mem3_reg[240][28]/P0001 , \wishbone_bd_ram_mem3_reg[240][29]/P0001 , \wishbone_bd_ram_mem3_reg[240][30]/P0001 , \wishbone_bd_ram_mem3_reg[240][31]/P0001 , \wishbone_bd_ram_mem3_reg[241][24]/P0001 , \wishbone_bd_ram_mem3_reg[241][25]/P0001 , \wishbone_bd_ram_mem3_reg[241][26]/P0001 , \wishbone_bd_ram_mem3_reg[241][27]/P0001 , \wishbone_bd_ram_mem3_reg[241][28]/P0001 , \wishbone_bd_ram_mem3_reg[241][29]/P0001 , \wishbone_bd_ram_mem3_reg[241][30]/P0001 , \wishbone_bd_ram_mem3_reg[241][31]/P0001 , \wishbone_bd_ram_mem3_reg[242][24]/P0001 , \wishbone_bd_ram_mem3_reg[242][25]/P0001 , \wishbone_bd_ram_mem3_reg[242][26]/P0001 , \wishbone_bd_ram_mem3_reg[242][27]/P0001 , \wishbone_bd_ram_mem3_reg[242][28]/P0001 , \wishbone_bd_ram_mem3_reg[242][29]/P0001 , \wishbone_bd_ram_mem3_reg[242][30]/P0001 , \wishbone_bd_ram_mem3_reg[242][31]/P0001 , \wishbone_bd_ram_mem3_reg[243][24]/P0001 , \wishbone_bd_ram_mem3_reg[243][25]/P0001 , \wishbone_bd_ram_mem3_reg[243][26]/P0001 , \wishbone_bd_ram_mem3_reg[243][27]/P0001 , \wishbone_bd_ram_mem3_reg[243][28]/P0001 , \wishbone_bd_ram_mem3_reg[243][29]/P0001 , \wishbone_bd_ram_mem3_reg[243][30]/P0001 , \wishbone_bd_ram_mem3_reg[243][31]/P0001 , \wishbone_bd_ram_mem3_reg[244][24]/P0001 , \wishbone_bd_ram_mem3_reg[244][25]/P0001 , \wishbone_bd_ram_mem3_reg[244][26]/P0001 , \wishbone_bd_ram_mem3_reg[244][27]/P0001 , \wishbone_bd_ram_mem3_reg[244][28]/P0001 , \wishbone_bd_ram_mem3_reg[244][29]/P0001 , \wishbone_bd_ram_mem3_reg[244][30]/P0001 , \wishbone_bd_ram_mem3_reg[244][31]/P0001 , \wishbone_bd_ram_mem3_reg[245][24]/P0001 , \wishbone_bd_ram_mem3_reg[245][25]/P0001 , \wishbone_bd_ram_mem3_reg[245][26]/P0001 , \wishbone_bd_ram_mem3_reg[245][27]/P0001 , \wishbone_bd_ram_mem3_reg[245][28]/P0001 , \wishbone_bd_ram_mem3_reg[245][29]/P0001 , \wishbone_bd_ram_mem3_reg[245][30]/P0001 , \wishbone_bd_ram_mem3_reg[245][31]/P0001 , \wishbone_bd_ram_mem3_reg[246][24]/P0001 , \wishbone_bd_ram_mem3_reg[246][25]/P0001 , \wishbone_bd_ram_mem3_reg[246][26]/P0001 , \wishbone_bd_ram_mem3_reg[246][27]/P0001 , \wishbone_bd_ram_mem3_reg[246][28]/P0001 , \wishbone_bd_ram_mem3_reg[246][29]/P0001 , \wishbone_bd_ram_mem3_reg[246][30]/P0001 , \wishbone_bd_ram_mem3_reg[246][31]/P0001 , \wishbone_bd_ram_mem3_reg[247][24]/P0001 , \wishbone_bd_ram_mem3_reg[247][25]/P0001 , \wishbone_bd_ram_mem3_reg[247][26]/P0001 , \wishbone_bd_ram_mem3_reg[247][27]/P0001 , \wishbone_bd_ram_mem3_reg[247][28]/P0001 , \wishbone_bd_ram_mem3_reg[247][29]/P0001 , \wishbone_bd_ram_mem3_reg[247][30]/P0001 , \wishbone_bd_ram_mem3_reg[247][31]/P0001 , \wishbone_bd_ram_mem3_reg[248][24]/P0001 , \wishbone_bd_ram_mem3_reg[248][25]/P0001 , \wishbone_bd_ram_mem3_reg[248][26]/P0001 , \wishbone_bd_ram_mem3_reg[248][27]/P0001 , \wishbone_bd_ram_mem3_reg[248][28]/P0001 , \wishbone_bd_ram_mem3_reg[248][29]/P0001 , \wishbone_bd_ram_mem3_reg[248][30]/P0001 , \wishbone_bd_ram_mem3_reg[248][31]/P0001 , \wishbone_bd_ram_mem3_reg[249][24]/P0001 , \wishbone_bd_ram_mem3_reg[249][25]/P0001 , \wishbone_bd_ram_mem3_reg[249][26]/P0001 , \wishbone_bd_ram_mem3_reg[249][27]/P0001 , \wishbone_bd_ram_mem3_reg[249][28]/P0001 , \wishbone_bd_ram_mem3_reg[249][29]/P0001 , \wishbone_bd_ram_mem3_reg[249][30]/P0001 , \wishbone_bd_ram_mem3_reg[249][31]/P0001 , \wishbone_bd_ram_mem3_reg[24][24]/P0001 , \wishbone_bd_ram_mem3_reg[24][25]/P0001 , \wishbone_bd_ram_mem3_reg[24][26]/P0001 , \wishbone_bd_ram_mem3_reg[24][27]/P0001 , \wishbone_bd_ram_mem3_reg[24][28]/P0001 , \wishbone_bd_ram_mem3_reg[24][29]/P0001 , \wishbone_bd_ram_mem3_reg[24][30]/P0001 , \wishbone_bd_ram_mem3_reg[24][31]/P0001 , \wishbone_bd_ram_mem3_reg[250][24]/P0001 , \wishbone_bd_ram_mem3_reg[250][25]/P0001 , \wishbone_bd_ram_mem3_reg[250][26]/P0001 , \wishbone_bd_ram_mem3_reg[250][27]/P0001 , \wishbone_bd_ram_mem3_reg[250][28]/P0001 , \wishbone_bd_ram_mem3_reg[250][29]/P0001 , \wishbone_bd_ram_mem3_reg[250][30]/P0001 , \wishbone_bd_ram_mem3_reg[250][31]/P0001 , \wishbone_bd_ram_mem3_reg[251][24]/P0001 , \wishbone_bd_ram_mem3_reg[251][25]/P0001 , \wishbone_bd_ram_mem3_reg[251][26]/P0001 , \wishbone_bd_ram_mem3_reg[251][27]/P0001 , \wishbone_bd_ram_mem3_reg[251][28]/P0001 , \wishbone_bd_ram_mem3_reg[251][29]/P0001 , \wishbone_bd_ram_mem3_reg[251][30]/P0001 , \wishbone_bd_ram_mem3_reg[251][31]/P0001 , \wishbone_bd_ram_mem3_reg[252][24]/P0001 , \wishbone_bd_ram_mem3_reg[252][25]/P0001 , \wishbone_bd_ram_mem3_reg[252][26]/P0001 , \wishbone_bd_ram_mem3_reg[252][27]/P0001 , \wishbone_bd_ram_mem3_reg[252][28]/P0001 , \wishbone_bd_ram_mem3_reg[252][29]/P0001 , \wishbone_bd_ram_mem3_reg[252][30]/P0001 , \wishbone_bd_ram_mem3_reg[252][31]/P0001 , \wishbone_bd_ram_mem3_reg[253][24]/P0001 , \wishbone_bd_ram_mem3_reg[253][25]/P0001 , \wishbone_bd_ram_mem3_reg[253][26]/P0001 , \wishbone_bd_ram_mem3_reg[253][27]/P0001 , \wishbone_bd_ram_mem3_reg[253][28]/P0001 , \wishbone_bd_ram_mem3_reg[253][29]/P0001 , \wishbone_bd_ram_mem3_reg[253][30]/P0001 , \wishbone_bd_ram_mem3_reg[253][31]/P0001 , \wishbone_bd_ram_mem3_reg[254][24]/P0001 , \wishbone_bd_ram_mem3_reg[254][25]/P0001 , \wishbone_bd_ram_mem3_reg[254][26]/P0001 , \wishbone_bd_ram_mem3_reg[254][27]/P0001 , \wishbone_bd_ram_mem3_reg[254][28]/P0001 , \wishbone_bd_ram_mem3_reg[254][29]/P0001 , \wishbone_bd_ram_mem3_reg[254][30]/P0001 , \wishbone_bd_ram_mem3_reg[254][31]/P0001 , \wishbone_bd_ram_mem3_reg[255][24]/P0001 , \wishbone_bd_ram_mem3_reg[255][25]/P0001 , \wishbone_bd_ram_mem3_reg[255][26]/P0001 , \wishbone_bd_ram_mem3_reg[255][27]/P0001 , \wishbone_bd_ram_mem3_reg[255][28]/P0001 , \wishbone_bd_ram_mem3_reg[255][29]/P0001 , \wishbone_bd_ram_mem3_reg[255][30]/P0001 , \wishbone_bd_ram_mem3_reg[255][31]/P0001 , \wishbone_bd_ram_mem3_reg[25][24]/P0001 , \wishbone_bd_ram_mem3_reg[25][25]/P0001 , \wishbone_bd_ram_mem3_reg[25][26]/P0001 , \wishbone_bd_ram_mem3_reg[25][27]/P0001 , \wishbone_bd_ram_mem3_reg[25][28]/P0001 , \wishbone_bd_ram_mem3_reg[25][29]/P0001 , \wishbone_bd_ram_mem3_reg[25][30]/P0001 , \wishbone_bd_ram_mem3_reg[25][31]/P0001 , \wishbone_bd_ram_mem3_reg[26][24]/P0001 , \wishbone_bd_ram_mem3_reg[26][25]/P0001 , \wishbone_bd_ram_mem3_reg[26][26]/P0001 , \wishbone_bd_ram_mem3_reg[26][27]/P0001 , \wishbone_bd_ram_mem3_reg[26][28]/P0001 , \wishbone_bd_ram_mem3_reg[26][29]/P0001 , \wishbone_bd_ram_mem3_reg[26][30]/P0001 , \wishbone_bd_ram_mem3_reg[26][31]/P0001 , \wishbone_bd_ram_mem3_reg[27][24]/P0001 , \wishbone_bd_ram_mem3_reg[27][25]/P0001 , \wishbone_bd_ram_mem3_reg[27][26]/P0001 , \wishbone_bd_ram_mem3_reg[27][27]/P0001 , \wishbone_bd_ram_mem3_reg[27][28]/P0001 , \wishbone_bd_ram_mem3_reg[27][29]/P0001 , \wishbone_bd_ram_mem3_reg[27][30]/P0001 , \wishbone_bd_ram_mem3_reg[27][31]/P0001 , \wishbone_bd_ram_mem3_reg[28][24]/P0001 , \wishbone_bd_ram_mem3_reg[28][25]/P0001 , \wishbone_bd_ram_mem3_reg[28][26]/P0001 , \wishbone_bd_ram_mem3_reg[28][27]/P0001 , \wishbone_bd_ram_mem3_reg[28][28]/P0001 , \wishbone_bd_ram_mem3_reg[28][29]/P0001 , \wishbone_bd_ram_mem3_reg[28][30]/P0001 , \wishbone_bd_ram_mem3_reg[28][31]/P0001 , \wishbone_bd_ram_mem3_reg[29][24]/P0001 , \wishbone_bd_ram_mem3_reg[29][25]/P0001 , \wishbone_bd_ram_mem3_reg[29][26]/P0001 , \wishbone_bd_ram_mem3_reg[29][27]/P0001 , \wishbone_bd_ram_mem3_reg[29][28]/P0001 , \wishbone_bd_ram_mem3_reg[29][29]/P0001 , \wishbone_bd_ram_mem3_reg[29][30]/P0001 , \wishbone_bd_ram_mem3_reg[29][31]/P0001 , \wishbone_bd_ram_mem3_reg[2][24]/P0001 , \wishbone_bd_ram_mem3_reg[2][25]/P0001 , \wishbone_bd_ram_mem3_reg[2][26]/P0001 , \wishbone_bd_ram_mem3_reg[2][27]/P0001 , \wishbone_bd_ram_mem3_reg[2][28]/P0001 , \wishbone_bd_ram_mem3_reg[2][29]/P0001 , \wishbone_bd_ram_mem3_reg[2][30]/P0001 , \wishbone_bd_ram_mem3_reg[2][31]/P0001 , \wishbone_bd_ram_mem3_reg[30][24]/P0001 , \wishbone_bd_ram_mem3_reg[30][25]/P0001 , \wishbone_bd_ram_mem3_reg[30][26]/P0001 , \wishbone_bd_ram_mem3_reg[30][27]/P0001 , \wishbone_bd_ram_mem3_reg[30][28]/P0001 , \wishbone_bd_ram_mem3_reg[30][29]/P0001 , \wishbone_bd_ram_mem3_reg[30][30]/P0001 , \wishbone_bd_ram_mem3_reg[30][31]/P0001 , \wishbone_bd_ram_mem3_reg[31][24]/P0001 , \wishbone_bd_ram_mem3_reg[31][25]/P0001 , \wishbone_bd_ram_mem3_reg[31][26]/P0001 , \wishbone_bd_ram_mem3_reg[31][27]/P0001 , \wishbone_bd_ram_mem3_reg[31][28]/P0001 , \wishbone_bd_ram_mem3_reg[31][29]/P0001 , \wishbone_bd_ram_mem3_reg[31][30]/P0001 , \wishbone_bd_ram_mem3_reg[31][31]/P0001 , \wishbone_bd_ram_mem3_reg[32][24]/P0001 , \wishbone_bd_ram_mem3_reg[32][25]/P0001 , \wishbone_bd_ram_mem3_reg[32][26]/P0001 , \wishbone_bd_ram_mem3_reg[32][27]/P0001 , \wishbone_bd_ram_mem3_reg[32][28]/P0001 , \wishbone_bd_ram_mem3_reg[32][29]/P0001 , \wishbone_bd_ram_mem3_reg[32][30]/P0001 , \wishbone_bd_ram_mem3_reg[32][31]/P0001 , \wishbone_bd_ram_mem3_reg[33][24]/P0001 , \wishbone_bd_ram_mem3_reg[33][25]/P0001 , \wishbone_bd_ram_mem3_reg[33][26]/P0001 , \wishbone_bd_ram_mem3_reg[33][27]/P0001 , \wishbone_bd_ram_mem3_reg[33][28]/P0001 , \wishbone_bd_ram_mem3_reg[33][29]/P0001 , \wishbone_bd_ram_mem3_reg[33][30]/P0001 , \wishbone_bd_ram_mem3_reg[33][31]/P0001 , \wishbone_bd_ram_mem3_reg[34][24]/P0001 , \wishbone_bd_ram_mem3_reg[34][25]/P0001 , \wishbone_bd_ram_mem3_reg[34][26]/P0001 , \wishbone_bd_ram_mem3_reg[34][27]/P0001 , \wishbone_bd_ram_mem3_reg[34][28]/P0001 , \wishbone_bd_ram_mem3_reg[34][29]/P0001 , \wishbone_bd_ram_mem3_reg[34][30]/P0001 , \wishbone_bd_ram_mem3_reg[34][31]/P0001 , \wishbone_bd_ram_mem3_reg[35][24]/P0001 , \wishbone_bd_ram_mem3_reg[35][25]/P0001 , \wishbone_bd_ram_mem3_reg[35][26]/P0001 , \wishbone_bd_ram_mem3_reg[35][27]/P0001 , \wishbone_bd_ram_mem3_reg[35][28]/P0001 , \wishbone_bd_ram_mem3_reg[35][29]/P0001 , \wishbone_bd_ram_mem3_reg[35][30]/P0001 , \wishbone_bd_ram_mem3_reg[35][31]/P0001 , \wishbone_bd_ram_mem3_reg[36][24]/P0001 , \wishbone_bd_ram_mem3_reg[36][25]/P0001 , \wishbone_bd_ram_mem3_reg[36][26]/P0001 , \wishbone_bd_ram_mem3_reg[36][27]/P0001 , \wishbone_bd_ram_mem3_reg[36][28]/P0001 , \wishbone_bd_ram_mem3_reg[36][29]/P0001 , \wishbone_bd_ram_mem3_reg[36][30]/P0001 , \wishbone_bd_ram_mem3_reg[36][31]/P0001 , \wishbone_bd_ram_mem3_reg[37][24]/P0001 , \wishbone_bd_ram_mem3_reg[37][25]/P0001 , \wishbone_bd_ram_mem3_reg[37][26]/P0001 , \wishbone_bd_ram_mem3_reg[37][27]/P0001 , \wishbone_bd_ram_mem3_reg[37][28]/P0001 , \wishbone_bd_ram_mem3_reg[37][29]/P0001 , \wishbone_bd_ram_mem3_reg[37][30]/P0001 , \wishbone_bd_ram_mem3_reg[37][31]/P0001 , \wishbone_bd_ram_mem3_reg[38][24]/P0001 , \wishbone_bd_ram_mem3_reg[38][25]/P0001 , \wishbone_bd_ram_mem3_reg[38][26]/P0001 , \wishbone_bd_ram_mem3_reg[38][27]/P0001 , \wishbone_bd_ram_mem3_reg[38][28]/P0001 , \wishbone_bd_ram_mem3_reg[38][29]/P0001 , \wishbone_bd_ram_mem3_reg[38][30]/P0001 , \wishbone_bd_ram_mem3_reg[38][31]/P0001 , \wishbone_bd_ram_mem3_reg[39][24]/P0001 , \wishbone_bd_ram_mem3_reg[39][25]/P0001 , \wishbone_bd_ram_mem3_reg[39][26]/P0001 , \wishbone_bd_ram_mem3_reg[39][27]/P0001 , \wishbone_bd_ram_mem3_reg[39][28]/P0001 , \wishbone_bd_ram_mem3_reg[39][29]/P0001 , \wishbone_bd_ram_mem3_reg[39][30]/P0001 , \wishbone_bd_ram_mem3_reg[39][31]/P0001 , \wishbone_bd_ram_mem3_reg[3][24]/P0001 , \wishbone_bd_ram_mem3_reg[3][25]/P0001 , \wishbone_bd_ram_mem3_reg[3][26]/P0001 , \wishbone_bd_ram_mem3_reg[3][27]/P0001 , \wishbone_bd_ram_mem3_reg[3][28]/P0001 , \wishbone_bd_ram_mem3_reg[3][29]/P0001 , \wishbone_bd_ram_mem3_reg[3][30]/P0001 , \wishbone_bd_ram_mem3_reg[3][31]/P0001 , \wishbone_bd_ram_mem3_reg[40][24]/P0001 , \wishbone_bd_ram_mem3_reg[40][25]/P0001 , \wishbone_bd_ram_mem3_reg[40][26]/P0001 , \wishbone_bd_ram_mem3_reg[40][27]/P0001 , \wishbone_bd_ram_mem3_reg[40][28]/P0001 , \wishbone_bd_ram_mem3_reg[40][29]/P0001 , \wishbone_bd_ram_mem3_reg[40][30]/P0001 , \wishbone_bd_ram_mem3_reg[40][31]/P0001 , \wishbone_bd_ram_mem3_reg[41][24]/P0001 , \wishbone_bd_ram_mem3_reg[41][25]/P0001 , \wishbone_bd_ram_mem3_reg[41][26]/P0001 , \wishbone_bd_ram_mem3_reg[41][27]/P0001 , \wishbone_bd_ram_mem3_reg[41][28]/P0001 , \wishbone_bd_ram_mem3_reg[41][29]/P0001 , \wishbone_bd_ram_mem3_reg[41][30]/P0001 , \wishbone_bd_ram_mem3_reg[41][31]/P0001 , \wishbone_bd_ram_mem3_reg[42][24]/P0001 , \wishbone_bd_ram_mem3_reg[42][25]/P0001 , \wishbone_bd_ram_mem3_reg[42][26]/P0001 , \wishbone_bd_ram_mem3_reg[42][27]/P0001 , \wishbone_bd_ram_mem3_reg[42][28]/P0001 , \wishbone_bd_ram_mem3_reg[42][29]/P0001 , \wishbone_bd_ram_mem3_reg[42][30]/P0001 , \wishbone_bd_ram_mem3_reg[42][31]/P0001 , \wishbone_bd_ram_mem3_reg[43][24]/P0001 , \wishbone_bd_ram_mem3_reg[43][25]/P0001 , \wishbone_bd_ram_mem3_reg[43][26]/P0001 , \wishbone_bd_ram_mem3_reg[43][27]/P0001 , \wishbone_bd_ram_mem3_reg[43][28]/P0001 , \wishbone_bd_ram_mem3_reg[43][29]/P0001 , \wishbone_bd_ram_mem3_reg[43][30]/P0001 , \wishbone_bd_ram_mem3_reg[43][31]/P0001 , \wishbone_bd_ram_mem3_reg[44][24]/P0001 , \wishbone_bd_ram_mem3_reg[44][25]/P0001 , \wishbone_bd_ram_mem3_reg[44][26]/P0001 , \wishbone_bd_ram_mem3_reg[44][27]/P0001 , \wishbone_bd_ram_mem3_reg[44][28]/P0001 , \wishbone_bd_ram_mem3_reg[44][29]/P0001 , \wishbone_bd_ram_mem3_reg[44][30]/P0001 , \wishbone_bd_ram_mem3_reg[44][31]/P0001 , \wishbone_bd_ram_mem3_reg[45][24]/P0001 , \wishbone_bd_ram_mem3_reg[45][25]/P0001 , \wishbone_bd_ram_mem3_reg[45][26]/P0001 , \wishbone_bd_ram_mem3_reg[45][27]/P0001 , \wishbone_bd_ram_mem3_reg[45][28]/P0001 , \wishbone_bd_ram_mem3_reg[45][29]/P0001 , \wishbone_bd_ram_mem3_reg[45][30]/P0001 , \wishbone_bd_ram_mem3_reg[45][31]/P0001 , \wishbone_bd_ram_mem3_reg[46][24]/P0001 , \wishbone_bd_ram_mem3_reg[46][25]/P0001 , \wishbone_bd_ram_mem3_reg[46][26]/P0001 , \wishbone_bd_ram_mem3_reg[46][27]/P0001 , \wishbone_bd_ram_mem3_reg[46][28]/P0001 , \wishbone_bd_ram_mem3_reg[46][29]/P0001 , \wishbone_bd_ram_mem3_reg[46][30]/P0001 , \wishbone_bd_ram_mem3_reg[46][31]/P0001 , \wishbone_bd_ram_mem3_reg[47][24]/P0001 , \wishbone_bd_ram_mem3_reg[47][25]/P0001 , \wishbone_bd_ram_mem3_reg[47][26]/P0001 , \wishbone_bd_ram_mem3_reg[47][27]/P0001 , \wishbone_bd_ram_mem3_reg[47][28]/P0001 , \wishbone_bd_ram_mem3_reg[47][29]/P0001 , \wishbone_bd_ram_mem3_reg[47][30]/P0001 , \wishbone_bd_ram_mem3_reg[47][31]/P0001 , \wishbone_bd_ram_mem3_reg[48][24]/P0001 , \wishbone_bd_ram_mem3_reg[48][25]/P0001 , \wishbone_bd_ram_mem3_reg[48][26]/P0001 , \wishbone_bd_ram_mem3_reg[48][27]/P0001 , \wishbone_bd_ram_mem3_reg[48][28]/P0001 , \wishbone_bd_ram_mem3_reg[48][29]/P0001 , \wishbone_bd_ram_mem3_reg[48][30]/P0001 , \wishbone_bd_ram_mem3_reg[48][31]/P0001 , \wishbone_bd_ram_mem3_reg[49][24]/P0001 , \wishbone_bd_ram_mem3_reg[49][25]/P0001 , \wishbone_bd_ram_mem3_reg[49][26]/P0001 , \wishbone_bd_ram_mem3_reg[49][27]/P0001 , \wishbone_bd_ram_mem3_reg[49][28]/P0001 , \wishbone_bd_ram_mem3_reg[49][29]/P0001 , \wishbone_bd_ram_mem3_reg[49][30]/P0001 , \wishbone_bd_ram_mem3_reg[49][31]/P0001 , \wishbone_bd_ram_mem3_reg[4][24]/P0001 , \wishbone_bd_ram_mem3_reg[4][25]/P0001 , \wishbone_bd_ram_mem3_reg[4][26]/P0001 , \wishbone_bd_ram_mem3_reg[4][27]/P0001 , \wishbone_bd_ram_mem3_reg[4][28]/P0001 , \wishbone_bd_ram_mem3_reg[4][29]/P0001 , \wishbone_bd_ram_mem3_reg[4][30]/P0001 , \wishbone_bd_ram_mem3_reg[4][31]/P0001 , \wishbone_bd_ram_mem3_reg[50][24]/P0001 , \wishbone_bd_ram_mem3_reg[50][25]/P0001 , \wishbone_bd_ram_mem3_reg[50][26]/P0001 , \wishbone_bd_ram_mem3_reg[50][27]/P0001 , \wishbone_bd_ram_mem3_reg[50][28]/P0001 , \wishbone_bd_ram_mem3_reg[50][29]/P0001 , \wishbone_bd_ram_mem3_reg[50][30]/P0001 , \wishbone_bd_ram_mem3_reg[50][31]/P0001 , \wishbone_bd_ram_mem3_reg[51][24]/P0001 , \wishbone_bd_ram_mem3_reg[51][25]/P0001 , \wishbone_bd_ram_mem3_reg[51][26]/P0001 , \wishbone_bd_ram_mem3_reg[51][27]/P0001 , \wishbone_bd_ram_mem3_reg[51][28]/P0001 , \wishbone_bd_ram_mem3_reg[51][29]/P0001 , \wishbone_bd_ram_mem3_reg[51][30]/P0001 , \wishbone_bd_ram_mem3_reg[51][31]/P0001 , \wishbone_bd_ram_mem3_reg[52][24]/P0001 , \wishbone_bd_ram_mem3_reg[52][25]/P0001 , \wishbone_bd_ram_mem3_reg[52][26]/P0001 , \wishbone_bd_ram_mem3_reg[52][27]/P0001 , \wishbone_bd_ram_mem3_reg[52][28]/P0001 , \wishbone_bd_ram_mem3_reg[52][29]/P0001 , \wishbone_bd_ram_mem3_reg[52][30]/P0001 , \wishbone_bd_ram_mem3_reg[52][31]/P0001 , \wishbone_bd_ram_mem3_reg[53][24]/P0001 , \wishbone_bd_ram_mem3_reg[53][25]/P0001 , \wishbone_bd_ram_mem3_reg[53][26]/P0001 , \wishbone_bd_ram_mem3_reg[53][27]/P0001 , \wishbone_bd_ram_mem3_reg[53][28]/P0001 , \wishbone_bd_ram_mem3_reg[53][29]/P0001 , \wishbone_bd_ram_mem3_reg[53][30]/P0001 , \wishbone_bd_ram_mem3_reg[53][31]/P0001 , \wishbone_bd_ram_mem3_reg[54][24]/P0001 , \wishbone_bd_ram_mem3_reg[54][25]/P0001 , \wishbone_bd_ram_mem3_reg[54][26]/P0001 , \wishbone_bd_ram_mem3_reg[54][27]/P0001 , \wishbone_bd_ram_mem3_reg[54][28]/P0001 , \wishbone_bd_ram_mem3_reg[54][29]/P0001 , \wishbone_bd_ram_mem3_reg[54][30]/P0001 , \wishbone_bd_ram_mem3_reg[54][31]/P0001 , \wishbone_bd_ram_mem3_reg[55][24]/P0001 , \wishbone_bd_ram_mem3_reg[55][25]/P0001 , \wishbone_bd_ram_mem3_reg[55][26]/P0001 , \wishbone_bd_ram_mem3_reg[55][27]/P0001 , \wishbone_bd_ram_mem3_reg[55][28]/P0001 , \wishbone_bd_ram_mem3_reg[55][29]/P0001 , \wishbone_bd_ram_mem3_reg[55][30]/P0001 , \wishbone_bd_ram_mem3_reg[55][31]/P0001 , \wishbone_bd_ram_mem3_reg[56][24]/P0001 , \wishbone_bd_ram_mem3_reg[56][25]/P0001 , \wishbone_bd_ram_mem3_reg[56][26]/P0001 , \wishbone_bd_ram_mem3_reg[56][27]/P0001 , \wishbone_bd_ram_mem3_reg[56][28]/P0001 , \wishbone_bd_ram_mem3_reg[56][29]/P0001 , \wishbone_bd_ram_mem3_reg[56][30]/P0001 , \wishbone_bd_ram_mem3_reg[56][31]/P0001 , \wishbone_bd_ram_mem3_reg[57][24]/P0001 , \wishbone_bd_ram_mem3_reg[57][25]/P0001 , \wishbone_bd_ram_mem3_reg[57][26]/P0001 , \wishbone_bd_ram_mem3_reg[57][27]/P0001 , \wishbone_bd_ram_mem3_reg[57][28]/P0001 , \wishbone_bd_ram_mem3_reg[57][29]/P0001 , \wishbone_bd_ram_mem3_reg[57][30]/P0001 , \wishbone_bd_ram_mem3_reg[57][31]/P0001 , \wishbone_bd_ram_mem3_reg[58][24]/P0001 , \wishbone_bd_ram_mem3_reg[58][25]/P0001 , \wishbone_bd_ram_mem3_reg[58][26]/P0001 , \wishbone_bd_ram_mem3_reg[58][27]/P0001 , \wishbone_bd_ram_mem3_reg[58][28]/P0001 , \wishbone_bd_ram_mem3_reg[58][29]/P0001 , \wishbone_bd_ram_mem3_reg[58][30]/P0001 , \wishbone_bd_ram_mem3_reg[58][31]/P0001 , \wishbone_bd_ram_mem3_reg[59][24]/P0001 , \wishbone_bd_ram_mem3_reg[59][25]/P0001 , \wishbone_bd_ram_mem3_reg[59][26]/P0001 , \wishbone_bd_ram_mem3_reg[59][27]/P0001 , \wishbone_bd_ram_mem3_reg[59][28]/P0001 , \wishbone_bd_ram_mem3_reg[59][29]/P0001 , \wishbone_bd_ram_mem3_reg[59][30]/P0001 , \wishbone_bd_ram_mem3_reg[59][31]/P0001 , \wishbone_bd_ram_mem3_reg[5][24]/P0001 , \wishbone_bd_ram_mem3_reg[5][25]/P0001 , \wishbone_bd_ram_mem3_reg[5][26]/P0001 , \wishbone_bd_ram_mem3_reg[5][27]/P0001 , \wishbone_bd_ram_mem3_reg[5][28]/P0001 , \wishbone_bd_ram_mem3_reg[5][29]/P0001 , \wishbone_bd_ram_mem3_reg[5][30]/P0001 , \wishbone_bd_ram_mem3_reg[5][31]/P0001 , \wishbone_bd_ram_mem3_reg[60][24]/P0001 , \wishbone_bd_ram_mem3_reg[60][25]/P0001 , \wishbone_bd_ram_mem3_reg[60][26]/P0001 , \wishbone_bd_ram_mem3_reg[60][27]/P0001 , \wishbone_bd_ram_mem3_reg[60][28]/P0001 , \wishbone_bd_ram_mem3_reg[60][29]/P0001 , \wishbone_bd_ram_mem3_reg[60][30]/P0001 , \wishbone_bd_ram_mem3_reg[60][31]/P0001 , \wishbone_bd_ram_mem3_reg[61][24]/P0001 , \wishbone_bd_ram_mem3_reg[61][25]/P0001 , \wishbone_bd_ram_mem3_reg[61][26]/P0001 , \wishbone_bd_ram_mem3_reg[61][27]/P0001 , \wishbone_bd_ram_mem3_reg[61][28]/P0001 , \wishbone_bd_ram_mem3_reg[61][29]/P0001 , \wishbone_bd_ram_mem3_reg[61][30]/P0001 , \wishbone_bd_ram_mem3_reg[61][31]/P0001 , \wishbone_bd_ram_mem3_reg[62][24]/P0001 , \wishbone_bd_ram_mem3_reg[62][25]/P0001 , \wishbone_bd_ram_mem3_reg[62][26]/P0001 , \wishbone_bd_ram_mem3_reg[62][27]/P0001 , \wishbone_bd_ram_mem3_reg[62][28]/P0001 , \wishbone_bd_ram_mem3_reg[62][29]/P0001 , \wishbone_bd_ram_mem3_reg[62][30]/P0001 , \wishbone_bd_ram_mem3_reg[62][31]/P0001 , \wishbone_bd_ram_mem3_reg[63][24]/P0001 , \wishbone_bd_ram_mem3_reg[63][25]/P0001 , \wishbone_bd_ram_mem3_reg[63][26]/P0001 , \wishbone_bd_ram_mem3_reg[63][27]/P0001 , \wishbone_bd_ram_mem3_reg[63][28]/P0001 , \wishbone_bd_ram_mem3_reg[63][29]/P0001 , \wishbone_bd_ram_mem3_reg[63][30]/P0001 , \wishbone_bd_ram_mem3_reg[63][31]/P0001 , \wishbone_bd_ram_mem3_reg[64][24]/P0001 , \wishbone_bd_ram_mem3_reg[64][25]/P0001 , \wishbone_bd_ram_mem3_reg[64][26]/P0001 , \wishbone_bd_ram_mem3_reg[64][27]/P0001 , \wishbone_bd_ram_mem3_reg[64][28]/P0001 , \wishbone_bd_ram_mem3_reg[64][29]/P0001 , \wishbone_bd_ram_mem3_reg[64][30]/P0001 , \wishbone_bd_ram_mem3_reg[64][31]/P0001 , \wishbone_bd_ram_mem3_reg[65][24]/P0001 , \wishbone_bd_ram_mem3_reg[65][25]/P0001 , \wishbone_bd_ram_mem3_reg[65][26]/P0001 , \wishbone_bd_ram_mem3_reg[65][27]/P0001 , \wishbone_bd_ram_mem3_reg[65][28]/P0001 , \wishbone_bd_ram_mem3_reg[65][29]/P0001 , \wishbone_bd_ram_mem3_reg[65][30]/P0001 , \wishbone_bd_ram_mem3_reg[65][31]/P0001 , \wishbone_bd_ram_mem3_reg[66][24]/P0001 , \wishbone_bd_ram_mem3_reg[66][25]/P0001 , \wishbone_bd_ram_mem3_reg[66][26]/P0001 , \wishbone_bd_ram_mem3_reg[66][27]/P0001 , \wishbone_bd_ram_mem3_reg[66][28]/P0001 , \wishbone_bd_ram_mem3_reg[66][29]/P0001 , \wishbone_bd_ram_mem3_reg[66][30]/P0001 , \wishbone_bd_ram_mem3_reg[66][31]/P0001 , \wishbone_bd_ram_mem3_reg[67][24]/P0001 , \wishbone_bd_ram_mem3_reg[67][25]/P0001 , \wishbone_bd_ram_mem3_reg[67][26]/P0001 , \wishbone_bd_ram_mem3_reg[67][27]/P0001 , \wishbone_bd_ram_mem3_reg[67][28]/P0001 , \wishbone_bd_ram_mem3_reg[67][29]/P0001 , \wishbone_bd_ram_mem3_reg[67][30]/P0001 , \wishbone_bd_ram_mem3_reg[67][31]/P0001 , \wishbone_bd_ram_mem3_reg[68][24]/P0001 , \wishbone_bd_ram_mem3_reg[68][25]/P0001 , \wishbone_bd_ram_mem3_reg[68][26]/P0001 , \wishbone_bd_ram_mem3_reg[68][27]/P0001 , \wishbone_bd_ram_mem3_reg[68][28]/P0001 , \wishbone_bd_ram_mem3_reg[68][29]/P0001 , \wishbone_bd_ram_mem3_reg[68][30]/P0001 , \wishbone_bd_ram_mem3_reg[68][31]/P0001 , \wishbone_bd_ram_mem3_reg[69][24]/P0001 , \wishbone_bd_ram_mem3_reg[69][25]/P0001 , \wishbone_bd_ram_mem3_reg[69][26]/P0001 , \wishbone_bd_ram_mem3_reg[69][27]/P0001 , \wishbone_bd_ram_mem3_reg[69][28]/P0001 , \wishbone_bd_ram_mem3_reg[69][29]/P0001 , \wishbone_bd_ram_mem3_reg[69][30]/P0001 , \wishbone_bd_ram_mem3_reg[69][31]/P0001 , \wishbone_bd_ram_mem3_reg[6][24]/P0001 , \wishbone_bd_ram_mem3_reg[6][25]/P0001 , \wishbone_bd_ram_mem3_reg[6][26]/P0001 , \wishbone_bd_ram_mem3_reg[6][27]/P0001 , \wishbone_bd_ram_mem3_reg[6][28]/P0001 , \wishbone_bd_ram_mem3_reg[6][29]/P0001 , \wishbone_bd_ram_mem3_reg[6][30]/P0001 , \wishbone_bd_ram_mem3_reg[6][31]/P0001 , \wishbone_bd_ram_mem3_reg[70][24]/P0001 , \wishbone_bd_ram_mem3_reg[70][25]/P0001 , \wishbone_bd_ram_mem3_reg[70][26]/P0001 , \wishbone_bd_ram_mem3_reg[70][27]/P0001 , \wishbone_bd_ram_mem3_reg[70][28]/P0001 , \wishbone_bd_ram_mem3_reg[70][29]/P0001 , \wishbone_bd_ram_mem3_reg[70][30]/P0001 , \wishbone_bd_ram_mem3_reg[70][31]/P0001 , \wishbone_bd_ram_mem3_reg[71][24]/P0001 , \wishbone_bd_ram_mem3_reg[71][25]/P0001 , \wishbone_bd_ram_mem3_reg[71][26]/P0001 , \wishbone_bd_ram_mem3_reg[71][27]/P0001 , \wishbone_bd_ram_mem3_reg[71][28]/P0001 , \wishbone_bd_ram_mem3_reg[71][29]/P0001 , \wishbone_bd_ram_mem3_reg[71][30]/P0001 , \wishbone_bd_ram_mem3_reg[71][31]/P0001 , \wishbone_bd_ram_mem3_reg[72][24]/P0001 , \wishbone_bd_ram_mem3_reg[72][25]/P0001 , \wishbone_bd_ram_mem3_reg[72][26]/P0001 , \wishbone_bd_ram_mem3_reg[72][27]/P0001 , \wishbone_bd_ram_mem3_reg[72][28]/P0001 , \wishbone_bd_ram_mem3_reg[72][29]/P0001 , \wishbone_bd_ram_mem3_reg[72][30]/P0001 , \wishbone_bd_ram_mem3_reg[72][31]/P0001 , \wishbone_bd_ram_mem3_reg[73][24]/P0001 , \wishbone_bd_ram_mem3_reg[73][25]/P0001 , \wishbone_bd_ram_mem3_reg[73][26]/P0001 , \wishbone_bd_ram_mem3_reg[73][27]/P0001 , \wishbone_bd_ram_mem3_reg[73][28]/P0001 , \wishbone_bd_ram_mem3_reg[73][29]/P0001 , \wishbone_bd_ram_mem3_reg[73][30]/P0001 , \wishbone_bd_ram_mem3_reg[73][31]/P0001 , \wishbone_bd_ram_mem3_reg[74][24]/P0001 , \wishbone_bd_ram_mem3_reg[74][25]/P0001 , \wishbone_bd_ram_mem3_reg[74][26]/P0001 , \wishbone_bd_ram_mem3_reg[74][27]/P0001 , \wishbone_bd_ram_mem3_reg[74][28]/P0001 , \wishbone_bd_ram_mem3_reg[74][29]/P0001 , \wishbone_bd_ram_mem3_reg[74][30]/P0001 , \wishbone_bd_ram_mem3_reg[74][31]/P0001 , \wishbone_bd_ram_mem3_reg[75][24]/P0001 , \wishbone_bd_ram_mem3_reg[75][25]/P0001 , \wishbone_bd_ram_mem3_reg[75][26]/P0001 , \wishbone_bd_ram_mem3_reg[75][27]/P0001 , \wishbone_bd_ram_mem3_reg[75][28]/P0001 , \wishbone_bd_ram_mem3_reg[75][29]/P0001 , \wishbone_bd_ram_mem3_reg[75][30]/P0001 , \wishbone_bd_ram_mem3_reg[75][31]/P0001 , \wishbone_bd_ram_mem3_reg[76][24]/P0001 , \wishbone_bd_ram_mem3_reg[76][25]/P0001 , \wishbone_bd_ram_mem3_reg[76][26]/P0001 , \wishbone_bd_ram_mem3_reg[76][27]/P0001 , \wishbone_bd_ram_mem3_reg[76][28]/P0001 , \wishbone_bd_ram_mem3_reg[76][29]/P0001 , \wishbone_bd_ram_mem3_reg[76][30]/P0001 , \wishbone_bd_ram_mem3_reg[76][31]/P0001 , \wishbone_bd_ram_mem3_reg[77][24]/P0001 , \wishbone_bd_ram_mem3_reg[77][25]/P0001 , \wishbone_bd_ram_mem3_reg[77][26]/P0001 , \wishbone_bd_ram_mem3_reg[77][27]/P0001 , \wishbone_bd_ram_mem3_reg[77][28]/P0001 , \wishbone_bd_ram_mem3_reg[77][29]/P0001 , \wishbone_bd_ram_mem3_reg[77][30]/P0001 , \wishbone_bd_ram_mem3_reg[77][31]/P0001 , \wishbone_bd_ram_mem3_reg[78][24]/P0001 , \wishbone_bd_ram_mem3_reg[78][25]/P0001 , \wishbone_bd_ram_mem3_reg[78][26]/P0001 , \wishbone_bd_ram_mem3_reg[78][27]/P0001 , \wishbone_bd_ram_mem3_reg[78][28]/P0001 , \wishbone_bd_ram_mem3_reg[78][29]/P0001 , \wishbone_bd_ram_mem3_reg[78][30]/P0001 , \wishbone_bd_ram_mem3_reg[78][31]/P0001 , \wishbone_bd_ram_mem3_reg[79][24]/P0001 , \wishbone_bd_ram_mem3_reg[79][25]/P0001 , \wishbone_bd_ram_mem3_reg[79][26]/P0001 , \wishbone_bd_ram_mem3_reg[79][27]/P0001 , \wishbone_bd_ram_mem3_reg[79][28]/P0001 , \wishbone_bd_ram_mem3_reg[79][29]/P0001 , \wishbone_bd_ram_mem3_reg[79][30]/P0001 , \wishbone_bd_ram_mem3_reg[79][31]/P0001 , \wishbone_bd_ram_mem3_reg[7][24]/P0001 , \wishbone_bd_ram_mem3_reg[7][25]/P0001 , \wishbone_bd_ram_mem3_reg[7][26]/P0001 , \wishbone_bd_ram_mem3_reg[7][27]/P0001 , \wishbone_bd_ram_mem3_reg[7][28]/P0001 , \wishbone_bd_ram_mem3_reg[7][29]/P0001 , \wishbone_bd_ram_mem3_reg[7][30]/P0001 , \wishbone_bd_ram_mem3_reg[7][31]/P0001 , \wishbone_bd_ram_mem3_reg[80][24]/P0001 , \wishbone_bd_ram_mem3_reg[80][25]/P0001 , \wishbone_bd_ram_mem3_reg[80][26]/P0001 , \wishbone_bd_ram_mem3_reg[80][27]/P0001 , \wishbone_bd_ram_mem3_reg[80][28]/P0001 , \wishbone_bd_ram_mem3_reg[80][29]/P0001 , \wishbone_bd_ram_mem3_reg[80][30]/P0001 , \wishbone_bd_ram_mem3_reg[80][31]/P0001 , \wishbone_bd_ram_mem3_reg[81][24]/P0001 , \wishbone_bd_ram_mem3_reg[81][25]/P0001 , \wishbone_bd_ram_mem3_reg[81][26]/P0001 , \wishbone_bd_ram_mem3_reg[81][27]/P0001 , \wishbone_bd_ram_mem3_reg[81][28]/P0001 , \wishbone_bd_ram_mem3_reg[81][29]/P0001 , \wishbone_bd_ram_mem3_reg[81][30]/P0001 , \wishbone_bd_ram_mem3_reg[81][31]/P0001 , \wishbone_bd_ram_mem3_reg[82][24]/P0001 , \wishbone_bd_ram_mem3_reg[82][25]/P0001 , \wishbone_bd_ram_mem3_reg[82][26]/P0001 , \wishbone_bd_ram_mem3_reg[82][27]/P0001 , \wishbone_bd_ram_mem3_reg[82][28]/P0001 , \wishbone_bd_ram_mem3_reg[82][29]/P0001 , \wishbone_bd_ram_mem3_reg[82][30]/P0001 , \wishbone_bd_ram_mem3_reg[82][31]/P0001 , \wishbone_bd_ram_mem3_reg[83][24]/P0001 , \wishbone_bd_ram_mem3_reg[83][25]/P0001 , \wishbone_bd_ram_mem3_reg[83][26]/P0001 , \wishbone_bd_ram_mem3_reg[83][27]/P0001 , \wishbone_bd_ram_mem3_reg[83][28]/P0001 , \wishbone_bd_ram_mem3_reg[83][29]/P0001 , \wishbone_bd_ram_mem3_reg[83][30]/P0001 , \wishbone_bd_ram_mem3_reg[83][31]/P0001 , \wishbone_bd_ram_mem3_reg[84][24]/P0001 , \wishbone_bd_ram_mem3_reg[84][25]/P0001 , \wishbone_bd_ram_mem3_reg[84][26]/P0001 , \wishbone_bd_ram_mem3_reg[84][27]/P0001 , \wishbone_bd_ram_mem3_reg[84][28]/P0001 , \wishbone_bd_ram_mem3_reg[84][29]/P0001 , \wishbone_bd_ram_mem3_reg[84][30]/P0001 , \wishbone_bd_ram_mem3_reg[84][31]/P0001 , \wishbone_bd_ram_mem3_reg[85][24]/P0001 , \wishbone_bd_ram_mem3_reg[85][25]/P0001 , \wishbone_bd_ram_mem3_reg[85][26]/P0001 , \wishbone_bd_ram_mem3_reg[85][27]/P0001 , \wishbone_bd_ram_mem3_reg[85][28]/P0001 , \wishbone_bd_ram_mem3_reg[85][29]/P0001 , \wishbone_bd_ram_mem3_reg[85][30]/P0001 , \wishbone_bd_ram_mem3_reg[85][31]/P0001 , \wishbone_bd_ram_mem3_reg[86][24]/P0001 , \wishbone_bd_ram_mem3_reg[86][25]/P0001 , \wishbone_bd_ram_mem3_reg[86][26]/P0001 , \wishbone_bd_ram_mem3_reg[86][27]/P0001 , \wishbone_bd_ram_mem3_reg[86][28]/P0001 , \wishbone_bd_ram_mem3_reg[86][29]/P0001 , \wishbone_bd_ram_mem3_reg[86][30]/P0001 , \wishbone_bd_ram_mem3_reg[86][31]/P0001 , \wishbone_bd_ram_mem3_reg[87][24]/P0001 , \wishbone_bd_ram_mem3_reg[87][25]/P0001 , \wishbone_bd_ram_mem3_reg[87][26]/P0001 , \wishbone_bd_ram_mem3_reg[87][27]/P0001 , \wishbone_bd_ram_mem3_reg[87][28]/P0001 , \wishbone_bd_ram_mem3_reg[87][29]/P0001 , \wishbone_bd_ram_mem3_reg[87][30]/P0001 , \wishbone_bd_ram_mem3_reg[87][31]/P0001 , \wishbone_bd_ram_mem3_reg[88][24]/P0001 , \wishbone_bd_ram_mem3_reg[88][25]/P0001 , \wishbone_bd_ram_mem3_reg[88][26]/P0001 , \wishbone_bd_ram_mem3_reg[88][27]/P0001 , \wishbone_bd_ram_mem3_reg[88][28]/P0001 , \wishbone_bd_ram_mem3_reg[88][29]/P0001 , \wishbone_bd_ram_mem3_reg[88][30]/P0001 , \wishbone_bd_ram_mem3_reg[88][31]/P0001 , \wishbone_bd_ram_mem3_reg[89][24]/P0001 , \wishbone_bd_ram_mem3_reg[89][25]/P0001 , \wishbone_bd_ram_mem3_reg[89][26]/P0001 , \wishbone_bd_ram_mem3_reg[89][27]/P0001 , \wishbone_bd_ram_mem3_reg[89][28]/P0001 , \wishbone_bd_ram_mem3_reg[89][29]/P0001 , \wishbone_bd_ram_mem3_reg[89][30]/P0001 , \wishbone_bd_ram_mem3_reg[89][31]/P0001 , \wishbone_bd_ram_mem3_reg[8][24]/P0001 , \wishbone_bd_ram_mem3_reg[8][25]/P0001 , \wishbone_bd_ram_mem3_reg[8][26]/P0001 , \wishbone_bd_ram_mem3_reg[8][27]/P0001 , \wishbone_bd_ram_mem3_reg[8][28]/P0001 , \wishbone_bd_ram_mem3_reg[8][29]/P0001 , \wishbone_bd_ram_mem3_reg[8][30]/P0001 , \wishbone_bd_ram_mem3_reg[8][31]/P0001 , \wishbone_bd_ram_mem3_reg[90][24]/P0001 , \wishbone_bd_ram_mem3_reg[90][25]/P0001 , \wishbone_bd_ram_mem3_reg[90][26]/P0001 , \wishbone_bd_ram_mem3_reg[90][27]/P0001 , \wishbone_bd_ram_mem3_reg[90][28]/P0001 , \wishbone_bd_ram_mem3_reg[90][29]/P0001 , \wishbone_bd_ram_mem3_reg[90][30]/P0001 , \wishbone_bd_ram_mem3_reg[90][31]/P0001 , \wishbone_bd_ram_mem3_reg[91][24]/P0001 , \wishbone_bd_ram_mem3_reg[91][25]/P0001 , \wishbone_bd_ram_mem3_reg[91][26]/P0001 , \wishbone_bd_ram_mem3_reg[91][27]/P0001 , \wishbone_bd_ram_mem3_reg[91][28]/P0001 , \wishbone_bd_ram_mem3_reg[91][29]/P0001 , \wishbone_bd_ram_mem3_reg[91][30]/P0001 , \wishbone_bd_ram_mem3_reg[91][31]/P0001 , \wishbone_bd_ram_mem3_reg[92][24]/P0001 , \wishbone_bd_ram_mem3_reg[92][25]/P0001 , \wishbone_bd_ram_mem3_reg[92][26]/P0001 , \wishbone_bd_ram_mem3_reg[92][27]/P0001 , \wishbone_bd_ram_mem3_reg[92][28]/P0001 , \wishbone_bd_ram_mem3_reg[92][29]/P0001 , \wishbone_bd_ram_mem3_reg[92][30]/P0001 , \wishbone_bd_ram_mem3_reg[92][31]/P0001 , \wishbone_bd_ram_mem3_reg[93][24]/P0001 , \wishbone_bd_ram_mem3_reg[93][25]/P0001 , \wishbone_bd_ram_mem3_reg[93][26]/P0001 , \wishbone_bd_ram_mem3_reg[93][27]/P0001 , \wishbone_bd_ram_mem3_reg[93][28]/P0001 , \wishbone_bd_ram_mem3_reg[93][29]/P0001 , \wishbone_bd_ram_mem3_reg[93][30]/P0001 , \wishbone_bd_ram_mem3_reg[93][31]/P0001 , \wishbone_bd_ram_mem3_reg[94][24]/P0001 , \wishbone_bd_ram_mem3_reg[94][25]/P0001 , \wishbone_bd_ram_mem3_reg[94][26]/P0001 , \wishbone_bd_ram_mem3_reg[94][27]/P0001 , \wishbone_bd_ram_mem3_reg[94][28]/P0001 , \wishbone_bd_ram_mem3_reg[94][29]/P0001 , \wishbone_bd_ram_mem3_reg[94][30]/P0001 , \wishbone_bd_ram_mem3_reg[94][31]/P0001 , \wishbone_bd_ram_mem3_reg[95][24]/P0001 , \wishbone_bd_ram_mem3_reg[95][25]/P0001 , \wishbone_bd_ram_mem3_reg[95][26]/P0001 , \wishbone_bd_ram_mem3_reg[95][27]/P0001 , \wishbone_bd_ram_mem3_reg[95][28]/P0001 , \wishbone_bd_ram_mem3_reg[95][29]/P0001 , \wishbone_bd_ram_mem3_reg[95][30]/P0001 , \wishbone_bd_ram_mem3_reg[95][31]/P0001 , \wishbone_bd_ram_mem3_reg[96][24]/P0001 , \wishbone_bd_ram_mem3_reg[96][25]/P0001 , \wishbone_bd_ram_mem3_reg[96][26]/P0001 , \wishbone_bd_ram_mem3_reg[96][27]/P0001 , \wishbone_bd_ram_mem3_reg[96][28]/P0001 , \wishbone_bd_ram_mem3_reg[96][29]/P0001 , \wishbone_bd_ram_mem3_reg[96][30]/P0001 , \wishbone_bd_ram_mem3_reg[96][31]/P0001 , \wishbone_bd_ram_mem3_reg[97][24]/P0001 , \wishbone_bd_ram_mem3_reg[97][25]/P0001 , \wishbone_bd_ram_mem3_reg[97][26]/P0001 , \wishbone_bd_ram_mem3_reg[97][27]/P0001 , \wishbone_bd_ram_mem3_reg[97][28]/P0001 , \wishbone_bd_ram_mem3_reg[97][29]/P0001 , \wishbone_bd_ram_mem3_reg[97][30]/P0001 , \wishbone_bd_ram_mem3_reg[97][31]/P0001 , \wishbone_bd_ram_mem3_reg[98][24]/P0001 , \wishbone_bd_ram_mem3_reg[98][25]/P0001 , \wishbone_bd_ram_mem3_reg[98][26]/P0001 , \wishbone_bd_ram_mem3_reg[98][27]/P0001 , \wishbone_bd_ram_mem3_reg[98][28]/P0001 , \wishbone_bd_ram_mem3_reg[98][29]/P0001 , \wishbone_bd_ram_mem3_reg[98][30]/P0001 , \wishbone_bd_ram_mem3_reg[98][31]/P0001 , \wishbone_bd_ram_mem3_reg[99][24]/P0001 , \wishbone_bd_ram_mem3_reg[99][25]/P0001 , \wishbone_bd_ram_mem3_reg[99][26]/P0001 , \wishbone_bd_ram_mem3_reg[99][27]/P0001 , \wishbone_bd_ram_mem3_reg[99][28]/P0001 , \wishbone_bd_ram_mem3_reg[99][29]/P0001 , \wishbone_bd_ram_mem3_reg[99][30]/P0001 , \wishbone_bd_ram_mem3_reg[99][31]/P0001 , \wishbone_bd_ram_mem3_reg[9][24]/P0001 , \wishbone_bd_ram_mem3_reg[9][25]/P0001 , \wishbone_bd_ram_mem3_reg[9][26]/P0001 , \wishbone_bd_ram_mem3_reg[9][27]/P0001 , \wishbone_bd_ram_mem3_reg[9][28]/P0001 , \wishbone_bd_ram_mem3_reg[9][29]/P0001 , \wishbone_bd_ram_mem3_reg[9][30]/P0001 , \wishbone_bd_ram_mem3_reg[9][31]/P0001 , \wishbone_bd_ram_raddr_reg[0]/P0001 , \wishbone_bd_ram_raddr_reg[1]/NET0131 , \wishbone_bd_ram_raddr_reg[2]/NET0131 , \wishbone_bd_ram_raddr_reg[3]/P0001 , \wishbone_bd_ram_raddr_reg[4]/NET0131 , \wishbone_bd_ram_raddr_reg[5]/NET0131 , \wishbone_bd_ram_raddr_reg[6]/NET0131 , \wishbone_bd_ram_raddr_reg[7]/NET0131 , \wishbone_cyc_cleared_reg/NET0131 , \wishbone_r_RxEn_q_reg/NET0131 , \wishbone_r_TxEn_q_reg/NET0131 , \wishbone_ram_addr_reg[0]/NET0131 , \wishbone_ram_addr_reg[1]/NET0131 , \wishbone_ram_addr_reg[2]/NET0131 , \wishbone_ram_addr_reg[3]/NET0131 , \wishbone_ram_addr_reg[4]/NET0131 , \wishbone_ram_addr_reg[5]/NET0131 , \wishbone_ram_addr_reg[6]/NET0131 , \wishbone_ram_addr_reg[7]/NET0131 , \wishbone_ram_di_reg[0]/NET0131 , \wishbone_ram_di_reg[10]/NET0131 , \wishbone_ram_di_reg[11]/NET0131 , \wishbone_ram_di_reg[12]/NET0131 , \wishbone_ram_di_reg[13]/NET0131 , \wishbone_ram_di_reg[14]/NET0131 , \wishbone_ram_di_reg[15]/NET0131 , \wishbone_ram_di_reg[16]/NET0131 , \wishbone_ram_di_reg[17]/NET0131 , \wishbone_ram_di_reg[18]/NET0131 , \wishbone_ram_di_reg[19]/NET0131 , \wishbone_ram_di_reg[1]/NET0131 , \wishbone_ram_di_reg[20]/NET0131 , \wishbone_ram_di_reg[21]/NET0131 , \wishbone_ram_di_reg[22]/NET0131 , \wishbone_ram_di_reg[23]/NET0131 , \wishbone_ram_di_reg[24]/NET0131 , \wishbone_ram_di_reg[25]/NET0131 , \wishbone_ram_di_reg[26]/NET0131 , \wishbone_ram_di_reg[27]/NET0131 , \wishbone_ram_di_reg[28]/NET0131 , \wishbone_ram_di_reg[29]/NET0131 , \wishbone_ram_di_reg[2]/NET0131 , \wishbone_ram_di_reg[30]/NET0131 , \wishbone_ram_di_reg[31]/NET0131 , \wishbone_ram_di_reg[3]/NET0131 , \wishbone_ram_di_reg[4]/NET0131 , \wishbone_ram_di_reg[5]/NET0131 , \wishbone_ram_di_reg[6]/NET0131 , \wishbone_ram_di_reg[7]/NET0131 , \wishbone_ram_di_reg[8]/NET0131 , \wishbone_ram_di_reg[9]/NET0131 , \wishbone_rx_burst_cnt_reg[0]/NET0131 , \wishbone_rx_burst_cnt_reg[1]/NET0131 , \wishbone_rx_burst_cnt_reg[2]/NET0131 , \wishbone_rx_burst_en_reg/NET0131 , \wishbone_rx_fifo_cnt_reg[0]/NET0131 , \wishbone_rx_fifo_cnt_reg[1]/NET0131 , \wishbone_rx_fifo_cnt_reg[2]/NET0131 , \wishbone_rx_fifo_cnt_reg[3]/NET0131 , \wishbone_rx_fifo_cnt_reg[4]/NET0131 , \wishbone_rx_fifo_fifo_reg[0][0]/P0001 , \wishbone_rx_fifo_fifo_reg[0][10]/P0001 , \wishbone_rx_fifo_fifo_reg[0][11]/P0001 , \wishbone_rx_fifo_fifo_reg[0][12]/P0001 , \wishbone_rx_fifo_fifo_reg[0][13]/P0001 , \wishbone_rx_fifo_fifo_reg[0][14]/P0001 , \wishbone_rx_fifo_fifo_reg[0][15]/P0001 , \wishbone_rx_fifo_fifo_reg[0][16]/P0001 , \wishbone_rx_fifo_fifo_reg[0][17]/P0001 , \wishbone_rx_fifo_fifo_reg[0][18]/P0001 , \wishbone_rx_fifo_fifo_reg[0][19]/P0001 , \wishbone_rx_fifo_fifo_reg[0][1]/P0001 , \wishbone_rx_fifo_fifo_reg[0][20]/P0001 , \wishbone_rx_fifo_fifo_reg[0][21]/P0001 , \wishbone_rx_fifo_fifo_reg[0][22]/P0001 , \wishbone_rx_fifo_fifo_reg[0][23]/P0001 , \wishbone_rx_fifo_fifo_reg[0][24]/P0001 , \wishbone_rx_fifo_fifo_reg[0][25]/P0001 , \wishbone_rx_fifo_fifo_reg[0][26]/P0001 , \wishbone_rx_fifo_fifo_reg[0][27]/P0001 , \wishbone_rx_fifo_fifo_reg[0][28]/P0001 , \wishbone_rx_fifo_fifo_reg[0][29]/P0001 , \wishbone_rx_fifo_fifo_reg[0][2]/P0001 , \wishbone_rx_fifo_fifo_reg[0][30]/P0001 , \wishbone_rx_fifo_fifo_reg[0][31]/P0001 , \wishbone_rx_fifo_fifo_reg[0][3]/P0001 , \wishbone_rx_fifo_fifo_reg[0][4]/P0001 , \wishbone_rx_fifo_fifo_reg[0][5]/P0001 , \wishbone_rx_fifo_fifo_reg[0][6]/P0001 , \wishbone_rx_fifo_fifo_reg[0][7]/P0001 , \wishbone_rx_fifo_fifo_reg[0][8]/P0001 , \wishbone_rx_fifo_fifo_reg[0][9]/P0001 , \wishbone_rx_fifo_fifo_reg[10][0]/P0001 , \wishbone_rx_fifo_fifo_reg[10][10]/P0001 , \wishbone_rx_fifo_fifo_reg[10][11]/P0001 , \wishbone_rx_fifo_fifo_reg[10][12]/P0001 , \wishbone_rx_fifo_fifo_reg[10][13]/P0001 , \wishbone_rx_fifo_fifo_reg[10][14]/P0001 , \wishbone_rx_fifo_fifo_reg[10][15]/P0001 , \wishbone_rx_fifo_fifo_reg[10][16]/P0001 , \wishbone_rx_fifo_fifo_reg[10][17]/P0001 , \wishbone_rx_fifo_fifo_reg[10][18]/P0001 , \wishbone_rx_fifo_fifo_reg[10][19]/P0001 , \wishbone_rx_fifo_fifo_reg[10][1]/P0001 , \wishbone_rx_fifo_fifo_reg[10][20]/P0001 , \wishbone_rx_fifo_fifo_reg[10][21]/P0001 , \wishbone_rx_fifo_fifo_reg[10][22]/P0001 , \wishbone_rx_fifo_fifo_reg[10][23]/P0001 , \wishbone_rx_fifo_fifo_reg[10][24]/P0001 , \wishbone_rx_fifo_fifo_reg[10][25]/P0001 , \wishbone_rx_fifo_fifo_reg[10][26]/P0001 , \wishbone_rx_fifo_fifo_reg[10][27]/P0001 , \wishbone_rx_fifo_fifo_reg[10][28]/P0001 , \wishbone_rx_fifo_fifo_reg[10][29]/P0001 , \wishbone_rx_fifo_fifo_reg[10][2]/P0001 , \wishbone_rx_fifo_fifo_reg[10][30]/P0001 , \wishbone_rx_fifo_fifo_reg[10][31]/P0001 , \wishbone_rx_fifo_fifo_reg[10][3]/P0001 , \wishbone_rx_fifo_fifo_reg[10][4]/P0001 , \wishbone_rx_fifo_fifo_reg[10][5]/P0001 , \wishbone_rx_fifo_fifo_reg[10][6]/P0001 , \wishbone_rx_fifo_fifo_reg[10][7]/P0001 , \wishbone_rx_fifo_fifo_reg[10][8]/P0001 , \wishbone_rx_fifo_fifo_reg[10][9]/P0001 , \wishbone_rx_fifo_fifo_reg[11][0]/P0001 , \wishbone_rx_fifo_fifo_reg[11][10]/P0001 , \wishbone_rx_fifo_fifo_reg[11][11]/P0001 , \wishbone_rx_fifo_fifo_reg[11][12]/P0001 , \wishbone_rx_fifo_fifo_reg[11][13]/P0001 , \wishbone_rx_fifo_fifo_reg[11][14]/P0001 , \wishbone_rx_fifo_fifo_reg[11][15]/P0001 , \wishbone_rx_fifo_fifo_reg[11][16]/P0001 , \wishbone_rx_fifo_fifo_reg[11][17]/P0001 , \wishbone_rx_fifo_fifo_reg[11][18]/P0001 , \wishbone_rx_fifo_fifo_reg[11][19]/P0001 , \wishbone_rx_fifo_fifo_reg[11][1]/P0001 , \wishbone_rx_fifo_fifo_reg[11][20]/P0001 , \wishbone_rx_fifo_fifo_reg[11][21]/P0001 , \wishbone_rx_fifo_fifo_reg[11][22]/P0001 , \wishbone_rx_fifo_fifo_reg[11][23]/P0001 , \wishbone_rx_fifo_fifo_reg[11][24]/P0001 , \wishbone_rx_fifo_fifo_reg[11][25]/P0001 , \wishbone_rx_fifo_fifo_reg[11][26]/P0001 , \wishbone_rx_fifo_fifo_reg[11][27]/P0001 , \wishbone_rx_fifo_fifo_reg[11][28]/P0001 , \wishbone_rx_fifo_fifo_reg[11][29]/P0001 , \wishbone_rx_fifo_fifo_reg[11][2]/P0001 , \wishbone_rx_fifo_fifo_reg[11][30]/P0001 , \wishbone_rx_fifo_fifo_reg[11][31]/P0001 , \wishbone_rx_fifo_fifo_reg[11][3]/P0001 , \wishbone_rx_fifo_fifo_reg[11][4]/P0001 , \wishbone_rx_fifo_fifo_reg[11][5]/P0001 , \wishbone_rx_fifo_fifo_reg[11][6]/P0001 , \wishbone_rx_fifo_fifo_reg[11][7]/P0001 , \wishbone_rx_fifo_fifo_reg[11][8]/P0001 , \wishbone_rx_fifo_fifo_reg[11][9]/P0001 , \wishbone_rx_fifo_fifo_reg[12][0]/P0001 , \wishbone_rx_fifo_fifo_reg[12][10]/P0001 , \wishbone_rx_fifo_fifo_reg[12][11]/P0001 , \wishbone_rx_fifo_fifo_reg[12][12]/P0001 , \wishbone_rx_fifo_fifo_reg[12][13]/P0001 , \wishbone_rx_fifo_fifo_reg[12][14]/P0001 , \wishbone_rx_fifo_fifo_reg[12][15]/P0001 , \wishbone_rx_fifo_fifo_reg[12][16]/P0001 , \wishbone_rx_fifo_fifo_reg[12][17]/P0001 , \wishbone_rx_fifo_fifo_reg[12][18]/P0001 , \wishbone_rx_fifo_fifo_reg[12][19]/P0001 , \wishbone_rx_fifo_fifo_reg[12][1]/P0001 , \wishbone_rx_fifo_fifo_reg[12][20]/P0001 , \wishbone_rx_fifo_fifo_reg[12][21]/P0001 , \wishbone_rx_fifo_fifo_reg[12][22]/P0001 , \wishbone_rx_fifo_fifo_reg[12][23]/P0001 , \wishbone_rx_fifo_fifo_reg[12][24]/P0001 , \wishbone_rx_fifo_fifo_reg[12][25]/P0001 , \wishbone_rx_fifo_fifo_reg[12][26]/P0001 , \wishbone_rx_fifo_fifo_reg[12][27]/P0001 , \wishbone_rx_fifo_fifo_reg[12][28]/P0001 , \wishbone_rx_fifo_fifo_reg[12][29]/P0001 , \wishbone_rx_fifo_fifo_reg[12][2]/P0001 , \wishbone_rx_fifo_fifo_reg[12][30]/P0001 , \wishbone_rx_fifo_fifo_reg[12][31]/P0001 , \wishbone_rx_fifo_fifo_reg[12][3]/P0001 , \wishbone_rx_fifo_fifo_reg[12][4]/P0001 , \wishbone_rx_fifo_fifo_reg[12][5]/P0001 , \wishbone_rx_fifo_fifo_reg[12][6]/P0001 , \wishbone_rx_fifo_fifo_reg[12][7]/P0001 , \wishbone_rx_fifo_fifo_reg[12][8]/P0001 , \wishbone_rx_fifo_fifo_reg[12][9]/P0001 , \wishbone_rx_fifo_fifo_reg[13][0]/P0001 , \wishbone_rx_fifo_fifo_reg[13][10]/P0001 , \wishbone_rx_fifo_fifo_reg[13][11]/P0001 , \wishbone_rx_fifo_fifo_reg[13][12]/P0001 , \wishbone_rx_fifo_fifo_reg[13][13]/P0001 , \wishbone_rx_fifo_fifo_reg[13][14]/P0001 , \wishbone_rx_fifo_fifo_reg[13][15]/P0001 , \wishbone_rx_fifo_fifo_reg[13][16]/P0001 , \wishbone_rx_fifo_fifo_reg[13][17]/P0001 , \wishbone_rx_fifo_fifo_reg[13][18]/P0001 , \wishbone_rx_fifo_fifo_reg[13][19]/P0001 , \wishbone_rx_fifo_fifo_reg[13][1]/P0001 , \wishbone_rx_fifo_fifo_reg[13][20]/P0001 , \wishbone_rx_fifo_fifo_reg[13][21]/P0001 , \wishbone_rx_fifo_fifo_reg[13][22]/P0001 , \wishbone_rx_fifo_fifo_reg[13][23]/P0001 , \wishbone_rx_fifo_fifo_reg[13][24]/P0001 , \wishbone_rx_fifo_fifo_reg[13][25]/P0001 , \wishbone_rx_fifo_fifo_reg[13][26]/P0001 , \wishbone_rx_fifo_fifo_reg[13][27]/P0001 , \wishbone_rx_fifo_fifo_reg[13][28]/P0001 , \wishbone_rx_fifo_fifo_reg[13][29]/P0001 , \wishbone_rx_fifo_fifo_reg[13][2]/P0001 , \wishbone_rx_fifo_fifo_reg[13][30]/P0001 , \wishbone_rx_fifo_fifo_reg[13][31]/P0001 , \wishbone_rx_fifo_fifo_reg[13][3]/P0001 , \wishbone_rx_fifo_fifo_reg[13][4]/P0001 , \wishbone_rx_fifo_fifo_reg[13][5]/P0001 , \wishbone_rx_fifo_fifo_reg[13][6]/P0001 , \wishbone_rx_fifo_fifo_reg[13][7]/P0001 , \wishbone_rx_fifo_fifo_reg[13][8]/P0001 , \wishbone_rx_fifo_fifo_reg[13][9]/P0001 , \wishbone_rx_fifo_fifo_reg[14][0]/P0001 , \wishbone_rx_fifo_fifo_reg[14][10]/P0001 , \wishbone_rx_fifo_fifo_reg[14][11]/P0001 , \wishbone_rx_fifo_fifo_reg[14][12]/P0001 , \wishbone_rx_fifo_fifo_reg[14][13]/P0001 , \wishbone_rx_fifo_fifo_reg[14][14]/P0001 , \wishbone_rx_fifo_fifo_reg[14][15]/P0001 , \wishbone_rx_fifo_fifo_reg[14][16]/P0001 , \wishbone_rx_fifo_fifo_reg[14][17]/P0001 , \wishbone_rx_fifo_fifo_reg[14][18]/P0001 , \wishbone_rx_fifo_fifo_reg[14][19]/P0001 , \wishbone_rx_fifo_fifo_reg[14][1]/P0001 , \wishbone_rx_fifo_fifo_reg[14][20]/P0001 , \wishbone_rx_fifo_fifo_reg[14][21]/P0001 , \wishbone_rx_fifo_fifo_reg[14][22]/P0001 , \wishbone_rx_fifo_fifo_reg[14][23]/P0001 , \wishbone_rx_fifo_fifo_reg[14][24]/P0001 , \wishbone_rx_fifo_fifo_reg[14][25]/P0001 , \wishbone_rx_fifo_fifo_reg[14][26]/P0001 , \wishbone_rx_fifo_fifo_reg[14][27]/P0001 , \wishbone_rx_fifo_fifo_reg[14][28]/P0001 , \wishbone_rx_fifo_fifo_reg[14][29]/P0001 , \wishbone_rx_fifo_fifo_reg[14][2]/P0001 , \wishbone_rx_fifo_fifo_reg[14][30]/P0001 , \wishbone_rx_fifo_fifo_reg[14][31]/P0001 , \wishbone_rx_fifo_fifo_reg[14][3]/P0001 , \wishbone_rx_fifo_fifo_reg[14][4]/P0001 , \wishbone_rx_fifo_fifo_reg[14][5]/P0001 , \wishbone_rx_fifo_fifo_reg[14][6]/P0001 , \wishbone_rx_fifo_fifo_reg[14][7]/P0001 , \wishbone_rx_fifo_fifo_reg[14][8]/P0001 , \wishbone_rx_fifo_fifo_reg[14][9]/P0001 , \wishbone_rx_fifo_fifo_reg[15][0]/P0001 , \wishbone_rx_fifo_fifo_reg[15][10]/P0001 , \wishbone_rx_fifo_fifo_reg[15][11]/P0001 , \wishbone_rx_fifo_fifo_reg[15][12]/P0001 , \wishbone_rx_fifo_fifo_reg[15][13]/P0001 , \wishbone_rx_fifo_fifo_reg[15][14]/P0001 , \wishbone_rx_fifo_fifo_reg[15][15]/P0001 , \wishbone_rx_fifo_fifo_reg[15][16]/P0001 , \wishbone_rx_fifo_fifo_reg[15][17]/P0001 , \wishbone_rx_fifo_fifo_reg[15][18]/P0001 , \wishbone_rx_fifo_fifo_reg[15][19]/P0001 , \wishbone_rx_fifo_fifo_reg[15][1]/P0001 , \wishbone_rx_fifo_fifo_reg[15][20]/P0001 , \wishbone_rx_fifo_fifo_reg[15][21]/P0001 , \wishbone_rx_fifo_fifo_reg[15][22]/P0001 , \wishbone_rx_fifo_fifo_reg[15][23]/P0001 , \wishbone_rx_fifo_fifo_reg[15][24]/P0001 , \wishbone_rx_fifo_fifo_reg[15][25]/P0001 , \wishbone_rx_fifo_fifo_reg[15][26]/P0001 , \wishbone_rx_fifo_fifo_reg[15][27]/P0001 , \wishbone_rx_fifo_fifo_reg[15][28]/P0001 , \wishbone_rx_fifo_fifo_reg[15][29]/P0001 , \wishbone_rx_fifo_fifo_reg[15][2]/P0001 , \wishbone_rx_fifo_fifo_reg[15][30]/P0001 , \wishbone_rx_fifo_fifo_reg[15][31]/P0001 , \wishbone_rx_fifo_fifo_reg[15][3]/P0001 , \wishbone_rx_fifo_fifo_reg[15][4]/P0001 , \wishbone_rx_fifo_fifo_reg[15][5]/P0001 , \wishbone_rx_fifo_fifo_reg[15][6]/P0001 , \wishbone_rx_fifo_fifo_reg[15][7]/P0001 , \wishbone_rx_fifo_fifo_reg[15][8]/P0001 , \wishbone_rx_fifo_fifo_reg[15][9]/P0001 , \wishbone_rx_fifo_fifo_reg[1][0]/P0001 , \wishbone_rx_fifo_fifo_reg[1][10]/P0001 , \wishbone_rx_fifo_fifo_reg[1][11]/P0001 , \wishbone_rx_fifo_fifo_reg[1][12]/P0001 , \wishbone_rx_fifo_fifo_reg[1][13]/P0001 , \wishbone_rx_fifo_fifo_reg[1][14]/P0001 , \wishbone_rx_fifo_fifo_reg[1][15]/P0001 , \wishbone_rx_fifo_fifo_reg[1][16]/P0001 , \wishbone_rx_fifo_fifo_reg[1][17]/P0001 , \wishbone_rx_fifo_fifo_reg[1][18]/P0001 , \wishbone_rx_fifo_fifo_reg[1][19]/P0001 , \wishbone_rx_fifo_fifo_reg[1][1]/P0001 , \wishbone_rx_fifo_fifo_reg[1][20]/P0001 , \wishbone_rx_fifo_fifo_reg[1][21]/P0001 , \wishbone_rx_fifo_fifo_reg[1][22]/P0001 , \wishbone_rx_fifo_fifo_reg[1][23]/P0001 , \wishbone_rx_fifo_fifo_reg[1][24]/P0001 , \wishbone_rx_fifo_fifo_reg[1][25]/P0001 , \wishbone_rx_fifo_fifo_reg[1][26]/P0001 , \wishbone_rx_fifo_fifo_reg[1][27]/P0001 , \wishbone_rx_fifo_fifo_reg[1][28]/P0001 , \wishbone_rx_fifo_fifo_reg[1][29]/P0001 , \wishbone_rx_fifo_fifo_reg[1][2]/P0001 , \wishbone_rx_fifo_fifo_reg[1][30]/P0001 , \wishbone_rx_fifo_fifo_reg[1][31]/P0001 , \wishbone_rx_fifo_fifo_reg[1][3]/P0001 , \wishbone_rx_fifo_fifo_reg[1][4]/P0001 , \wishbone_rx_fifo_fifo_reg[1][5]/P0001 , \wishbone_rx_fifo_fifo_reg[1][6]/P0001 , \wishbone_rx_fifo_fifo_reg[1][7]/P0001 , \wishbone_rx_fifo_fifo_reg[1][8]/P0001 , \wishbone_rx_fifo_fifo_reg[1][9]/P0001 , \wishbone_rx_fifo_fifo_reg[2][0]/P0001 , \wishbone_rx_fifo_fifo_reg[2][10]/P0001 , \wishbone_rx_fifo_fifo_reg[2][11]/P0001 , \wishbone_rx_fifo_fifo_reg[2][12]/P0001 , \wishbone_rx_fifo_fifo_reg[2][13]/P0001 , \wishbone_rx_fifo_fifo_reg[2][14]/P0001 , \wishbone_rx_fifo_fifo_reg[2][15]/P0001 , \wishbone_rx_fifo_fifo_reg[2][16]/P0001 , \wishbone_rx_fifo_fifo_reg[2][17]/P0001 , \wishbone_rx_fifo_fifo_reg[2][18]/P0001 , \wishbone_rx_fifo_fifo_reg[2][19]/P0001 , \wishbone_rx_fifo_fifo_reg[2][1]/P0001 , \wishbone_rx_fifo_fifo_reg[2][20]/P0001 , \wishbone_rx_fifo_fifo_reg[2][21]/P0001 , \wishbone_rx_fifo_fifo_reg[2][22]/P0001 , \wishbone_rx_fifo_fifo_reg[2][23]/P0001 , \wishbone_rx_fifo_fifo_reg[2][24]/P0001 , \wishbone_rx_fifo_fifo_reg[2][25]/P0001 , \wishbone_rx_fifo_fifo_reg[2][26]/P0001 , \wishbone_rx_fifo_fifo_reg[2][27]/P0001 , \wishbone_rx_fifo_fifo_reg[2][28]/P0001 , \wishbone_rx_fifo_fifo_reg[2][29]/P0001 , \wishbone_rx_fifo_fifo_reg[2][2]/P0001 , \wishbone_rx_fifo_fifo_reg[2][30]/P0001 , \wishbone_rx_fifo_fifo_reg[2][31]/P0001 , \wishbone_rx_fifo_fifo_reg[2][3]/P0001 , \wishbone_rx_fifo_fifo_reg[2][4]/P0001 , \wishbone_rx_fifo_fifo_reg[2][5]/P0001 , \wishbone_rx_fifo_fifo_reg[2][6]/P0001 , \wishbone_rx_fifo_fifo_reg[2][7]/P0001 , \wishbone_rx_fifo_fifo_reg[2][8]/P0001 , \wishbone_rx_fifo_fifo_reg[2][9]/P0001 , \wishbone_rx_fifo_fifo_reg[3][0]/P0001 , \wishbone_rx_fifo_fifo_reg[3][10]/P0001 , \wishbone_rx_fifo_fifo_reg[3][11]/P0001 , \wishbone_rx_fifo_fifo_reg[3][12]/P0001 , \wishbone_rx_fifo_fifo_reg[3][13]/P0001 , \wishbone_rx_fifo_fifo_reg[3][14]/P0001 , \wishbone_rx_fifo_fifo_reg[3][15]/P0001 , \wishbone_rx_fifo_fifo_reg[3][16]/P0001 , \wishbone_rx_fifo_fifo_reg[3][17]/P0001 , \wishbone_rx_fifo_fifo_reg[3][18]/P0001 , \wishbone_rx_fifo_fifo_reg[3][19]/P0001 , \wishbone_rx_fifo_fifo_reg[3][1]/P0001 , \wishbone_rx_fifo_fifo_reg[3][20]/P0001 , \wishbone_rx_fifo_fifo_reg[3][21]/P0001 , \wishbone_rx_fifo_fifo_reg[3][22]/P0001 , \wishbone_rx_fifo_fifo_reg[3][23]/P0001 , \wishbone_rx_fifo_fifo_reg[3][24]/P0001 , \wishbone_rx_fifo_fifo_reg[3][25]/P0001 , \wishbone_rx_fifo_fifo_reg[3][26]/P0001 , \wishbone_rx_fifo_fifo_reg[3][27]/P0001 , \wishbone_rx_fifo_fifo_reg[3][28]/P0001 , \wishbone_rx_fifo_fifo_reg[3][29]/P0001 , \wishbone_rx_fifo_fifo_reg[3][2]/P0001 , \wishbone_rx_fifo_fifo_reg[3][30]/P0001 , \wishbone_rx_fifo_fifo_reg[3][31]/P0001 , \wishbone_rx_fifo_fifo_reg[3][3]/P0001 , \wishbone_rx_fifo_fifo_reg[3][4]/P0001 , \wishbone_rx_fifo_fifo_reg[3][5]/P0001 , \wishbone_rx_fifo_fifo_reg[3][6]/P0001 , \wishbone_rx_fifo_fifo_reg[3][7]/P0001 , \wishbone_rx_fifo_fifo_reg[3][8]/P0001 , \wishbone_rx_fifo_fifo_reg[3][9]/P0001 , \wishbone_rx_fifo_fifo_reg[4][0]/P0001 , \wishbone_rx_fifo_fifo_reg[4][10]/P0001 , \wishbone_rx_fifo_fifo_reg[4][11]/P0001 , \wishbone_rx_fifo_fifo_reg[4][12]/P0001 , \wishbone_rx_fifo_fifo_reg[4][13]/P0001 , \wishbone_rx_fifo_fifo_reg[4][14]/P0001 , \wishbone_rx_fifo_fifo_reg[4][15]/P0001 , \wishbone_rx_fifo_fifo_reg[4][16]/P0001 , \wishbone_rx_fifo_fifo_reg[4][17]/P0001 , \wishbone_rx_fifo_fifo_reg[4][18]/P0001 , \wishbone_rx_fifo_fifo_reg[4][19]/P0001 , \wishbone_rx_fifo_fifo_reg[4][1]/P0001 , \wishbone_rx_fifo_fifo_reg[4][20]/P0001 , \wishbone_rx_fifo_fifo_reg[4][21]/P0001 , \wishbone_rx_fifo_fifo_reg[4][22]/P0001 , \wishbone_rx_fifo_fifo_reg[4][23]/P0001 , \wishbone_rx_fifo_fifo_reg[4][24]/P0001 , \wishbone_rx_fifo_fifo_reg[4][25]/P0001 , \wishbone_rx_fifo_fifo_reg[4][26]/P0001 , \wishbone_rx_fifo_fifo_reg[4][27]/P0001 , \wishbone_rx_fifo_fifo_reg[4][28]/P0001 , \wishbone_rx_fifo_fifo_reg[4][29]/P0001 , \wishbone_rx_fifo_fifo_reg[4][2]/P0001 , \wishbone_rx_fifo_fifo_reg[4][30]/P0001 , \wishbone_rx_fifo_fifo_reg[4][31]/P0001 , \wishbone_rx_fifo_fifo_reg[4][3]/P0001 , \wishbone_rx_fifo_fifo_reg[4][4]/P0001 , \wishbone_rx_fifo_fifo_reg[4][5]/P0001 , \wishbone_rx_fifo_fifo_reg[4][6]/P0001 , \wishbone_rx_fifo_fifo_reg[4][7]/P0001 , \wishbone_rx_fifo_fifo_reg[4][8]/P0001 , \wishbone_rx_fifo_fifo_reg[4][9]/P0001 , \wishbone_rx_fifo_fifo_reg[5][0]/P0001 , \wishbone_rx_fifo_fifo_reg[5][10]/P0001 , \wishbone_rx_fifo_fifo_reg[5][11]/P0001 , \wishbone_rx_fifo_fifo_reg[5][12]/P0001 , \wishbone_rx_fifo_fifo_reg[5][13]/P0001 , \wishbone_rx_fifo_fifo_reg[5][14]/P0001 , \wishbone_rx_fifo_fifo_reg[5][15]/P0001 , \wishbone_rx_fifo_fifo_reg[5][16]/P0001 , \wishbone_rx_fifo_fifo_reg[5][17]/P0001 , \wishbone_rx_fifo_fifo_reg[5][18]/P0001 , \wishbone_rx_fifo_fifo_reg[5][19]/P0001 , \wishbone_rx_fifo_fifo_reg[5][1]/P0001 , \wishbone_rx_fifo_fifo_reg[5][20]/P0001 , \wishbone_rx_fifo_fifo_reg[5][21]/P0001 , \wishbone_rx_fifo_fifo_reg[5][22]/P0001 , \wishbone_rx_fifo_fifo_reg[5][23]/P0001 , \wishbone_rx_fifo_fifo_reg[5][24]/P0001 , \wishbone_rx_fifo_fifo_reg[5][25]/P0001 , \wishbone_rx_fifo_fifo_reg[5][26]/P0001 , \wishbone_rx_fifo_fifo_reg[5][27]/P0001 , \wishbone_rx_fifo_fifo_reg[5][28]/P0001 , \wishbone_rx_fifo_fifo_reg[5][29]/P0001 , \wishbone_rx_fifo_fifo_reg[5][2]/P0001 , \wishbone_rx_fifo_fifo_reg[5][30]/P0001 , \wishbone_rx_fifo_fifo_reg[5][31]/P0001 , \wishbone_rx_fifo_fifo_reg[5][3]/P0001 , \wishbone_rx_fifo_fifo_reg[5][4]/P0001 , \wishbone_rx_fifo_fifo_reg[5][5]/P0001 , \wishbone_rx_fifo_fifo_reg[5][6]/P0001 , \wishbone_rx_fifo_fifo_reg[5][7]/P0001 , \wishbone_rx_fifo_fifo_reg[5][8]/P0001 , \wishbone_rx_fifo_fifo_reg[5][9]/P0001 , \wishbone_rx_fifo_fifo_reg[6][0]/P0001 , \wishbone_rx_fifo_fifo_reg[6][10]/P0001 , \wishbone_rx_fifo_fifo_reg[6][11]/P0001 , \wishbone_rx_fifo_fifo_reg[6][12]/P0001 , \wishbone_rx_fifo_fifo_reg[6][13]/P0001 , \wishbone_rx_fifo_fifo_reg[6][14]/P0001 , \wishbone_rx_fifo_fifo_reg[6][15]/P0001 , \wishbone_rx_fifo_fifo_reg[6][16]/P0001 , \wishbone_rx_fifo_fifo_reg[6][17]/P0001 , \wishbone_rx_fifo_fifo_reg[6][18]/P0001 , \wishbone_rx_fifo_fifo_reg[6][19]/P0001 , \wishbone_rx_fifo_fifo_reg[6][1]/P0001 , \wishbone_rx_fifo_fifo_reg[6][20]/P0001 , \wishbone_rx_fifo_fifo_reg[6][21]/P0001 , \wishbone_rx_fifo_fifo_reg[6][22]/P0001 , \wishbone_rx_fifo_fifo_reg[6][23]/P0001 , \wishbone_rx_fifo_fifo_reg[6][24]/P0001 , \wishbone_rx_fifo_fifo_reg[6][25]/P0001 , \wishbone_rx_fifo_fifo_reg[6][26]/P0001 , \wishbone_rx_fifo_fifo_reg[6][27]/P0001 , \wishbone_rx_fifo_fifo_reg[6][28]/P0001 , \wishbone_rx_fifo_fifo_reg[6][29]/P0001 , \wishbone_rx_fifo_fifo_reg[6][2]/P0001 , \wishbone_rx_fifo_fifo_reg[6][30]/P0001 , \wishbone_rx_fifo_fifo_reg[6][31]/P0001 , \wishbone_rx_fifo_fifo_reg[6][3]/P0001 , \wishbone_rx_fifo_fifo_reg[6][4]/P0001 , \wishbone_rx_fifo_fifo_reg[6][5]/P0001 , \wishbone_rx_fifo_fifo_reg[6][6]/P0001 , \wishbone_rx_fifo_fifo_reg[6][7]/P0001 , \wishbone_rx_fifo_fifo_reg[6][8]/P0001 , \wishbone_rx_fifo_fifo_reg[6][9]/P0001 , \wishbone_rx_fifo_fifo_reg[7][0]/P0001 , \wishbone_rx_fifo_fifo_reg[7][10]/P0001 , \wishbone_rx_fifo_fifo_reg[7][11]/P0001 , \wishbone_rx_fifo_fifo_reg[7][12]/P0001 , \wishbone_rx_fifo_fifo_reg[7][13]/P0001 , \wishbone_rx_fifo_fifo_reg[7][14]/P0001 , \wishbone_rx_fifo_fifo_reg[7][15]/P0001 , \wishbone_rx_fifo_fifo_reg[7][16]/P0001 , \wishbone_rx_fifo_fifo_reg[7][17]/P0001 , \wishbone_rx_fifo_fifo_reg[7][18]/P0001 , \wishbone_rx_fifo_fifo_reg[7][19]/P0001 , \wishbone_rx_fifo_fifo_reg[7][1]/P0001 , \wishbone_rx_fifo_fifo_reg[7][20]/P0001 , \wishbone_rx_fifo_fifo_reg[7][21]/P0001 , \wishbone_rx_fifo_fifo_reg[7][22]/P0001 , \wishbone_rx_fifo_fifo_reg[7][23]/P0001 , \wishbone_rx_fifo_fifo_reg[7][24]/P0001 , \wishbone_rx_fifo_fifo_reg[7][25]/P0001 , \wishbone_rx_fifo_fifo_reg[7][26]/P0001 , \wishbone_rx_fifo_fifo_reg[7][27]/P0001 , \wishbone_rx_fifo_fifo_reg[7][28]/P0001 , \wishbone_rx_fifo_fifo_reg[7][29]/P0001 , \wishbone_rx_fifo_fifo_reg[7][2]/P0001 , \wishbone_rx_fifo_fifo_reg[7][30]/P0001 , \wishbone_rx_fifo_fifo_reg[7][31]/P0001 , \wishbone_rx_fifo_fifo_reg[7][3]/P0001 , \wishbone_rx_fifo_fifo_reg[7][4]/P0001 , \wishbone_rx_fifo_fifo_reg[7][5]/P0001 , \wishbone_rx_fifo_fifo_reg[7][6]/P0001 , \wishbone_rx_fifo_fifo_reg[7][7]/P0001 , \wishbone_rx_fifo_fifo_reg[7][8]/P0001 , \wishbone_rx_fifo_fifo_reg[7][9]/P0001 , \wishbone_rx_fifo_fifo_reg[8][0]/P0001 , \wishbone_rx_fifo_fifo_reg[8][10]/P0001 , \wishbone_rx_fifo_fifo_reg[8][11]/P0001 , \wishbone_rx_fifo_fifo_reg[8][12]/P0001 , \wishbone_rx_fifo_fifo_reg[8][13]/P0001 , \wishbone_rx_fifo_fifo_reg[8][14]/P0001 , \wishbone_rx_fifo_fifo_reg[8][15]/P0001 , \wishbone_rx_fifo_fifo_reg[8][16]/P0001 , \wishbone_rx_fifo_fifo_reg[8][17]/P0001 , \wishbone_rx_fifo_fifo_reg[8][18]/P0001 , \wishbone_rx_fifo_fifo_reg[8][19]/P0001 , \wishbone_rx_fifo_fifo_reg[8][1]/P0001 , \wishbone_rx_fifo_fifo_reg[8][20]/P0001 , \wishbone_rx_fifo_fifo_reg[8][21]/P0001 , \wishbone_rx_fifo_fifo_reg[8][22]/P0001 , \wishbone_rx_fifo_fifo_reg[8][23]/P0001 , \wishbone_rx_fifo_fifo_reg[8][24]/P0001 , \wishbone_rx_fifo_fifo_reg[8][25]/P0001 , \wishbone_rx_fifo_fifo_reg[8][26]/P0001 , \wishbone_rx_fifo_fifo_reg[8][27]/P0001 , \wishbone_rx_fifo_fifo_reg[8][28]/P0001 , \wishbone_rx_fifo_fifo_reg[8][29]/P0001 , \wishbone_rx_fifo_fifo_reg[8][2]/P0001 , \wishbone_rx_fifo_fifo_reg[8][30]/P0001 , \wishbone_rx_fifo_fifo_reg[8][31]/P0001 , \wishbone_rx_fifo_fifo_reg[8][3]/P0001 , \wishbone_rx_fifo_fifo_reg[8][4]/P0001 , \wishbone_rx_fifo_fifo_reg[8][5]/P0001 , \wishbone_rx_fifo_fifo_reg[8][6]/P0001 , \wishbone_rx_fifo_fifo_reg[8][7]/P0001 , \wishbone_rx_fifo_fifo_reg[8][8]/P0001 , \wishbone_rx_fifo_fifo_reg[8][9]/P0001 , \wishbone_rx_fifo_fifo_reg[9][0]/P0001 , \wishbone_rx_fifo_fifo_reg[9][10]/P0001 , \wishbone_rx_fifo_fifo_reg[9][11]/P0001 , \wishbone_rx_fifo_fifo_reg[9][12]/P0001 , \wishbone_rx_fifo_fifo_reg[9][13]/P0001 , \wishbone_rx_fifo_fifo_reg[9][14]/P0001 , \wishbone_rx_fifo_fifo_reg[9][15]/P0001 , \wishbone_rx_fifo_fifo_reg[9][16]/P0001 , \wishbone_rx_fifo_fifo_reg[9][17]/P0001 , \wishbone_rx_fifo_fifo_reg[9][18]/P0001 , \wishbone_rx_fifo_fifo_reg[9][19]/P0001 , \wishbone_rx_fifo_fifo_reg[9][1]/P0001 , \wishbone_rx_fifo_fifo_reg[9][20]/P0001 , \wishbone_rx_fifo_fifo_reg[9][21]/P0001 , \wishbone_rx_fifo_fifo_reg[9][22]/P0001 , \wishbone_rx_fifo_fifo_reg[9][23]/P0001 , \wishbone_rx_fifo_fifo_reg[9][24]/P0001 , \wishbone_rx_fifo_fifo_reg[9][25]/P0001 , \wishbone_rx_fifo_fifo_reg[9][26]/P0001 , \wishbone_rx_fifo_fifo_reg[9][27]/P0001 , \wishbone_rx_fifo_fifo_reg[9][28]/P0001 , \wishbone_rx_fifo_fifo_reg[9][29]/P0001 , \wishbone_rx_fifo_fifo_reg[9][2]/P0001 , \wishbone_rx_fifo_fifo_reg[9][30]/P0001 , \wishbone_rx_fifo_fifo_reg[9][31]/P0001 , \wishbone_rx_fifo_fifo_reg[9][3]/P0001 , \wishbone_rx_fifo_fifo_reg[9][4]/P0001 , \wishbone_rx_fifo_fifo_reg[9][5]/P0001 , \wishbone_rx_fifo_fifo_reg[9][6]/P0001 , \wishbone_rx_fifo_fifo_reg[9][7]/P0001 , \wishbone_rx_fifo_fifo_reg[9][8]/P0001 , \wishbone_rx_fifo_fifo_reg[9][9]/P0001 , \wishbone_rx_fifo_read_pointer_reg[0]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[1]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[2]/NET0131 , \wishbone_rx_fifo_read_pointer_reg[3]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[0]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[1]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[2]/NET0131 , \wishbone_rx_fifo_write_pointer_reg[3]/NET0131 , \wishbone_tx_burst_cnt_reg[0]/NET0131 , \wishbone_tx_burst_cnt_reg[1]/NET0131 , \wishbone_tx_burst_cnt_reg[2]/NET0131 , \wishbone_tx_burst_en_reg/NET0131 , \wishbone_tx_fifo_cnt_reg[0]/NET0131 , \wishbone_tx_fifo_cnt_reg[1]/NET0131 , \wishbone_tx_fifo_cnt_reg[2]/NET0131 , \wishbone_tx_fifo_cnt_reg[3]/NET0131 , \wishbone_tx_fifo_cnt_reg[4]/NET0131 , \wishbone_tx_fifo_data_out_reg[0]/P0001 , \wishbone_tx_fifo_data_out_reg[10]/P0001 , \wishbone_tx_fifo_data_out_reg[11]/P0001 , \wishbone_tx_fifo_data_out_reg[12]/P0001 , \wishbone_tx_fifo_data_out_reg[13]/P0001 , \wishbone_tx_fifo_data_out_reg[14]/P0001 , \wishbone_tx_fifo_data_out_reg[15]/P0001 , \wishbone_tx_fifo_data_out_reg[16]/P0001 , \wishbone_tx_fifo_data_out_reg[17]/P0001 , \wishbone_tx_fifo_data_out_reg[18]/P0001 , \wishbone_tx_fifo_data_out_reg[19]/P0001 , \wishbone_tx_fifo_data_out_reg[1]/P0001 , \wishbone_tx_fifo_data_out_reg[20]/P0001 , \wishbone_tx_fifo_data_out_reg[21]/P0001 , \wishbone_tx_fifo_data_out_reg[22]/P0001 , \wishbone_tx_fifo_data_out_reg[23]/P0001 , \wishbone_tx_fifo_data_out_reg[24]/P0001 , \wishbone_tx_fifo_data_out_reg[25]/P0001 , \wishbone_tx_fifo_data_out_reg[26]/P0001 , \wishbone_tx_fifo_data_out_reg[27]/P0001 , \wishbone_tx_fifo_data_out_reg[28]/P0001 , \wishbone_tx_fifo_data_out_reg[29]/P0001 , \wishbone_tx_fifo_data_out_reg[2]/P0001 , \wishbone_tx_fifo_data_out_reg[30]/P0001 , \wishbone_tx_fifo_data_out_reg[31]/P0001 , \wishbone_tx_fifo_data_out_reg[3]/P0001 , \wishbone_tx_fifo_data_out_reg[4]/P0001 , \wishbone_tx_fifo_data_out_reg[5]/P0001 , \wishbone_tx_fifo_data_out_reg[6]/P0001 , \wishbone_tx_fifo_data_out_reg[7]/P0001 , \wishbone_tx_fifo_data_out_reg[8]/P0001 , \wishbone_tx_fifo_data_out_reg[9]/P0001 , \wishbone_tx_fifo_fifo_reg[0][0]/P0001 , \wishbone_tx_fifo_fifo_reg[0][10]/P0001 , \wishbone_tx_fifo_fifo_reg[0][11]/P0001 , \wishbone_tx_fifo_fifo_reg[0][12]/P0001 , \wishbone_tx_fifo_fifo_reg[0][13]/P0001 , \wishbone_tx_fifo_fifo_reg[0][14]/P0001 , \wishbone_tx_fifo_fifo_reg[0][15]/P0001 , \wishbone_tx_fifo_fifo_reg[0][16]/P0001 , \wishbone_tx_fifo_fifo_reg[0][17]/P0001 , \wishbone_tx_fifo_fifo_reg[0][18]/P0001 , \wishbone_tx_fifo_fifo_reg[0][19]/P0001 , \wishbone_tx_fifo_fifo_reg[0][1]/P0001 , \wishbone_tx_fifo_fifo_reg[0][20]/P0001 , \wishbone_tx_fifo_fifo_reg[0][21]/P0001 , \wishbone_tx_fifo_fifo_reg[0][22]/P0001 , \wishbone_tx_fifo_fifo_reg[0][23]/P0001 , \wishbone_tx_fifo_fifo_reg[0][24]/P0001 , \wishbone_tx_fifo_fifo_reg[0][25]/P0001 , \wishbone_tx_fifo_fifo_reg[0][26]/P0001 , \wishbone_tx_fifo_fifo_reg[0][27]/P0001 , \wishbone_tx_fifo_fifo_reg[0][28]/P0001 , \wishbone_tx_fifo_fifo_reg[0][29]/P0001 , \wishbone_tx_fifo_fifo_reg[0][2]/P0001 , \wishbone_tx_fifo_fifo_reg[0][30]/P0001 , \wishbone_tx_fifo_fifo_reg[0][31]/P0001 , \wishbone_tx_fifo_fifo_reg[0][3]/P0001 , \wishbone_tx_fifo_fifo_reg[0][4]/P0001 , \wishbone_tx_fifo_fifo_reg[0][5]/P0001 , \wishbone_tx_fifo_fifo_reg[0][6]/P0001 , \wishbone_tx_fifo_fifo_reg[0][7]/P0001 , \wishbone_tx_fifo_fifo_reg[0][8]/P0001 , \wishbone_tx_fifo_fifo_reg[0][9]/P0001 , \wishbone_tx_fifo_fifo_reg[10][0]/P0001 , \wishbone_tx_fifo_fifo_reg[10][10]/P0001 , \wishbone_tx_fifo_fifo_reg[10][11]/P0001 , \wishbone_tx_fifo_fifo_reg[10][12]/P0001 , \wishbone_tx_fifo_fifo_reg[10][13]/P0001 , \wishbone_tx_fifo_fifo_reg[10][14]/P0001 , \wishbone_tx_fifo_fifo_reg[10][15]/P0001 , \wishbone_tx_fifo_fifo_reg[10][16]/P0001 , \wishbone_tx_fifo_fifo_reg[10][17]/P0001 , \wishbone_tx_fifo_fifo_reg[10][18]/P0001 , \wishbone_tx_fifo_fifo_reg[10][19]/P0001 , \wishbone_tx_fifo_fifo_reg[10][1]/P0001 , \wishbone_tx_fifo_fifo_reg[10][20]/P0001 , \wishbone_tx_fifo_fifo_reg[10][21]/P0001 , \wishbone_tx_fifo_fifo_reg[10][22]/P0001 , \wishbone_tx_fifo_fifo_reg[10][23]/P0001 , \wishbone_tx_fifo_fifo_reg[10][24]/P0001 , \wishbone_tx_fifo_fifo_reg[10][25]/P0001 , \wishbone_tx_fifo_fifo_reg[10][26]/P0001 , \wishbone_tx_fifo_fifo_reg[10][27]/P0001 , \wishbone_tx_fifo_fifo_reg[10][28]/P0001 , \wishbone_tx_fifo_fifo_reg[10][29]/P0001 , \wishbone_tx_fifo_fifo_reg[10][2]/P0001 , \wishbone_tx_fifo_fifo_reg[10][30]/P0001 , \wishbone_tx_fifo_fifo_reg[10][31]/P0001 , \wishbone_tx_fifo_fifo_reg[10][3]/P0001 , \wishbone_tx_fifo_fifo_reg[10][4]/P0001 , \wishbone_tx_fifo_fifo_reg[10][5]/P0001 , \wishbone_tx_fifo_fifo_reg[10][6]/P0001 , \wishbone_tx_fifo_fifo_reg[10][7]/P0001 , \wishbone_tx_fifo_fifo_reg[10][8]/P0001 , \wishbone_tx_fifo_fifo_reg[10][9]/P0001 , \wishbone_tx_fifo_fifo_reg[11][0]/P0001 , \wishbone_tx_fifo_fifo_reg[11][10]/P0001 , \wishbone_tx_fifo_fifo_reg[11][11]/P0001 , \wishbone_tx_fifo_fifo_reg[11][12]/P0001 , \wishbone_tx_fifo_fifo_reg[11][13]/P0001 , \wishbone_tx_fifo_fifo_reg[11][14]/P0001 , \wishbone_tx_fifo_fifo_reg[11][15]/P0001 , \wishbone_tx_fifo_fifo_reg[11][16]/P0001 , \wishbone_tx_fifo_fifo_reg[11][17]/P0001 , \wishbone_tx_fifo_fifo_reg[11][18]/P0001 , \wishbone_tx_fifo_fifo_reg[11][19]/P0001 , \wishbone_tx_fifo_fifo_reg[11][1]/P0001 , \wishbone_tx_fifo_fifo_reg[11][20]/P0001 , \wishbone_tx_fifo_fifo_reg[11][21]/P0001 , \wishbone_tx_fifo_fifo_reg[11][22]/P0001 , \wishbone_tx_fifo_fifo_reg[11][23]/P0001 , \wishbone_tx_fifo_fifo_reg[11][24]/P0001 , \wishbone_tx_fifo_fifo_reg[11][25]/P0001 , \wishbone_tx_fifo_fifo_reg[11][26]/P0001 , \wishbone_tx_fifo_fifo_reg[11][27]/P0001 , \wishbone_tx_fifo_fifo_reg[11][28]/P0001 , \wishbone_tx_fifo_fifo_reg[11][29]/P0001 , \wishbone_tx_fifo_fifo_reg[11][2]/P0001 , \wishbone_tx_fifo_fifo_reg[11][30]/P0001 , \wishbone_tx_fifo_fifo_reg[11][31]/P0001 , \wishbone_tx_fifo_fifo_reg[11][3]/P0001 , \wishbone_tx_fifo_fifo_reg[11][4]/P0001 , \wishbone_tx_fifo_fifo_reg[11][5]/P0001 , \wishbone_tx_fifo_fifo_reg[11][6]/P0001 , \wishbone_tx_fifo_fifo_reg[11][7]/P0001 , \wishbone_tx_fifo_fifo_reg[11][8]/P0001 , \wishbone_tx_fifo_fifo_reg[11][9]/P0001 , \wishbone_tx_fifo_fifo_reg[12][0]/P0001 , \wishbone_tx_fifo_fifo_reg[12][10]/P0001 , \wishbone_tx_fifo_fifo_reg[12][11]/P0001 , \wishbone_tx_fifo_fifo_reg[12][12]/P0001 , \wishbone_tx_fifo_fifo_reg[12][13]/P0001 , \wishbone_tx_fifo_fifo_reg[12][14]/P0001 , \wishbone_tx_fifo_fifo_reg[12][15]/P0001 , \wishbone_tx_fifo_fifo_reg[12][16]/P0001 , \wishbone_tx_fifo_fifo_reg[12][17]/P0001 , \wishbone_tx_fifo_fifo_reg[12][18]/P0001 , \wishbone_tx_fifo_fifo_reg[12][19]/P0001 , \wishbone_tx_fifo_fifo_reg[12][1]/P0001 , \wishbone_tx_fifo_fifo_reg[12][20]/P0001 , \wishbone_tx_fifo_fifo_reg[12][21]/P0001 , \wishbone_tx_fifo_fifo_reg[12][22]/P0001 , \wishbone_tx_fifo_fifo_reg[12][23]/P0001 , \wishbone_tx_fifo_fifo_reg[12][24]/P0001 , \wishbone_tx_fifo_fifo_reg[12][25]/P0001 , \wishbone_tx_fifo_fifo_reg[12][26]/P0001 , \wishbone_tx_fifo_fifo_reg[12][27]/P0001 , \wishbone_tx_fifo_fifo_reg[12][28]/P0001 , \wishbone_tx_fifo_fifo_reg[12][29]/P0001 , \wishbone_tx_fifo_fifo_reg[12][2]/P0001 , \wishbone_tx_fifo_fifo_reg[12][30]/P0001 , \wishbone_tx_fifo_fifo_reg[12][31]/P0001 , \wishbone_tx_fifo_fifo_reg[12][3]/P0001 , \wishbone_tx_fifo_fifo_reg[12][4]/P0001 , \wishbone_tx_fifo_fifo_reg[12][5]/P0001 , \wishbone_tx_fifo_fifo_reg[12][6]/P0001 , \wishbone_tx_fifo_fifo_reg[12][7]/P0001 , \wishbone_tx_fifo_fifo_reg[12][8]/P0001 , \wishbone_tx_fifo_fifo_reg[12][9]/P0001 , \wishbone_tx_fifo_fifo_reg[13][0]/P0001 , \wishbone_tx_fifo_fifo_reg[13][10]/P0001 , \wishbone_tx_fifo_fifo_reg[13][11]/P0001 , \wishbone_tx_fifo_fifo_reg[13][12]/P0001 , \wishbone_tx_fifo_fifo_reg[13][13]/P0001 , \wishbone_tx_fifo_fifo_reg[13][14]/P0001 , \wishbone_tx_fifo_fifo_reg[13][15]/P0001 , \wishbone_tx_fifo_fifo_reg[13][16]/P0001 , \wishbone_tx_fifo_fifo_reg[13][17]/P0001 , \wishbone_tx_fifo_fifo_reg[13][18]/P0001 , \wishbone_tx_fifo_fifo_reg[13][19]/P0001 , \wishbone_tx_fifo_fifo_reg[13][1]/P0001 , \wishbone_tx_fifo_fifo_reg[13][20]/P0001 , \wishbone_tx_fifo_fifo_reg[13][21]/P0001 , \wishbone_tx_fifo_fifo_reg[13][22]/P0001 , \wishbone_tx_fifo_fifo_reg[13][23]/P0001 , \wishbone_tx_fifo_fifo_reg[13][24]/P0001 , \wishbone_tx_fifo_fifo_reg[13][25]/P0001 , \wishbone_tx_fifo_fifo_reg[13][26]/P0001 , \wishbone_tx_fifo_fifo_reg[13][27]/P0001 , \wishbone_tx_fifo_fifo_reg[13][28]/P0001 , \wishbone_tx_fifo_fifo_reg[13][29]/P0001 , \wishbone_tx_fifo_fifo_reg[13][2]/P0001 , \wishbone_tx_fifo_fifo_reg[13][30]/P0001 , \wishbone_tx_fifo_fifo_reg[13][31]/P0001 , \wishbone_tx_fifo_fifo_reg[13][3]/P0001 , \wishbone_tx_fifo_fifo_reg[13][4]/P0001 , \wishbone_tx_fifo_fifo_reg[13][5]/P0001 , \wishbone_tx_fifo_fifo_reg[13][6]/P0001 , \wishbone_tx_fifo_fifo_reg[13][7]/P0001 , \wishbone_tx_fifo_fifo_reg[13][8]/P0001 , \wishbone_tx_fifo_fifo_reg[13][9]/P0001 , \wishbone_tx_fifo_fifo_reg[14][0]/P0001 , \wishbone_tx_fifo_fifo_reg[14][10]/P0001 , \wishbone_tx_fifo_fifo_reg[14][11]/P0001 , \wishbone_tx_fifo_fifo_reg[14][12]/P0001 , \wishbone_tx_fifo_fifo_reg[14][13]/P0001 , \wishbone_tx_fifo_fifo_reg[14][14]/P0001 , \wishbone_tx_fifo_fifo_reg[14][15]/P0001 , \wishbone_tx_fifo_fifo_reg[14][16]/P0001 , \wishbone_tx_fifo_fifo_reg[14][17]/P0001 , \wishbone_tx_fifo_fifo_reg[14][18]/P0001 , \wishbone_tx_fifo_fifo_reg[14][19]/P0001 , \wishbone_tx_fifo_fifo_reg[14][1]/P0001 , \wishbone_tx_fifo_fifo_reg[14][20]/P0001 , \wishbone_tx_fifo_fifo_reg[14][21]/P0001 , \wishbone_tx_fifo_fifo_reg[14][22]/P0001 , \wishbone_tx_fifo_fifo_reg[14][23]/P0001 , \wishbone_tx_fifo_fifo_reg[14][24]/P0001 , \wishbone_tx_fifo_fifo_reg[14][25]/P0001 , \wishbone_tx_fifo_fifo_reg[14][26]/P0001 , \wishbone_tx_fifo_fifo_reg[14][27]/P0001 , \wishbone_tx_fifo_fifo_reg[14][28]/P0001 , \wishbone_tx_fifo_fifo_reg[14][29]/P0001 , \wishbone_tx_fifo_fifo_reg[14][2]/P0001 , \wishbone_tx_fifo_fifo_reg[14][30]/P0001 , \wishbone_tx_fifo_fifo_reg[14][31]/P0001 , \wishbone_tx_fifo_fifo_reg[14][3]/P0001 , \wishbone_tx_fifo_fifo_reg[14][4]/P0001 , \wishbone_tx_fifo_fifo_reg[14][5]/P0001 , \wishbone_tx_fifo_fifo_reg[14][6]/P0001 , \wishbone_tx_fifo_fifo_reg[14][7]/P0001 , \wishbone_tx_fifo_fifo_reg[14][8]/P0001 , \wishbone_tx_fifo_fifo_reg[14][9]/P0001 , \wishbone_tx_fifo_fifo_reg[15][0]/P0001 , \wishbone_tx_fifo_fifo_reg[15][10]/P0001 , \wishbone_tx_fifo_fifo_reg[15][11]/P0001 , \wishbone_tx_fifo_fifo_reg[15][12]/P0001 , \wishbone_tx_fifo_fifo_reg[15][13]/P0001 , \wishbone_tx_fifo_fifo_reg[15][14]/P0001 , \wishbone_tx_fifo_fifo_reg[15][15]/P0001 , \wishbone_tx_fifo_fifo_reg[15][16]/P0001 , \wishbone_tx_fifo_fifo_reg[15][17]/P0001 , \wishbone_tx_fifo_fifo_reg[15][18]/P0001 , \wishbone_tx_fifo_fifo_reg[15][19]/P0001 , \wishbone_tx_fifo_fifo_reg[15][1]/P0001 , \wishbone_tx_fifo_fifo_reg[15][20]/P0001 , \wishbone_tx_fifo_fifo_reg[15][21]/P0001 , \wishbone_tx_fifo_fifo_reg[15][22]/P0001 , \wishbone_tx_fifo_fifo_reg[15][23]/P0001 , \wishbone_tx_fifo_fifo_reg[15][24]/P0001 , \wishbone_tx_fifo_fifo_reg[15][25]/P0001 , \wishbone_tx_fifo_fifo_reg[15][26]/P0001 , \wishbone_tx_fifo_fifo_reg[15][27]/P0001 , \wishbone_tx_fifo_fifo_reg[15][28]/P0001 , \wishbone_tx_fifo_fifo_reg[15][29]/P0001 , \wishbone_tx_fifo_fifo_reg[15][2]/P0001 , \wishbone_tx_fifo_fifo_reg[15][30]/P0001 , \wishbone_tx_fifo_fifo_reg[15][31]/P0001 , \wishbone_tx_fifo_fifo_reg[15][3]/P0001 , \wishbone_tx_fifo_fifo_reg[15][4]/P0001 , \wishbone_tx_fifo_fifo_reg[15][5]/P0001 , \wishbone_tx_fifo_fifo_reg[15][6]/P0001 , \wishbone_tx_fifo_fifo_reg[15][7]/P0001 , \wishbone_tx_fifo_fifo_reg[15][8]/P0001 , \wishbone_tx_fifo_fifo_reg[15][9]/P0001 , \wishbone_tx_fifo_fifo_reg[1][0]/P0001 , \wishbone_tx_fifo_fifo_reg[1][10]/P0001 , \wishbone_tx_fifo_fifo_reg[1][11]/P0001 , \wishbone_tx_fifo_fifo_reg[1][12]/P0001 , \wishbone_tx_fifo_fifo_reg[1][13]/P0001 , \wishbone_tx_fifo_fifo_reg[1][14]/P0001 , \wishbone_tx_fifo_fifo_reg[1][15]/P0001 , \wishbone_tx_fifo_fifo_reg[1][16]/P0001 , \wishbone_tx_fifo_fifo_reg[1][17]/P0001 , \wishbone_tx_fifo_fifo_reg[1][18]/P0001 , \wishbone_tx_fifo_fifo_reg[1][19]/P0001 , \wishbone_tx_fifo_fifo_reg[1][1]/P0001 , \wishbone_tx_fifo_fifo_reg[1][20]/P0001 , \wishbone_tx_fifo_fifo_reg[1][21]/P0001 , \wishbone_tx_fifo_fifo_reg[1][22]/P0001 , \wishbone_tx_fifo_fifo_reg[1][23]/P0001 , \wishbone_tx_fifo_fifo_reg[1][24]/P0001 , \wishbone_tx_fifo_fifo_reg[1][25]/P0001 , \wishbone_tx_fifo_fifo_reg[1][26]/P0001 , \wishbone_tx_fifo_fifo_reg[1][27]/P0001 , \wishbone_tx_fifo_fifo_reg[1][28]/P0001 , \wishbone_tx_fifo_fifo_reg[1][29]/P0001 , \wishbone_tx_fifo_fifo_reg[1][2]/P0001 , \wishbone_tx_fifo_fifo_reg[1][30]/P0001 , \wishbone_tx_fifo_fifo_reg[1][31]/P0001 , \wishbone_tx_fifo_fifo_reg[1][3]/P0001 , \wishbone_tx_fifo_fifo_reg[1][4]/P0001 , \wishbone_tx_fifo_fifo_reg[1][5]/P0001 , \wishbone_tx_fifo_fifo_reg[1][6]/P0001 , \wishbone_tx_fifo_fifo_reg[1][7]/P0001 , \wishbone_tx_fifo_fifo_reg[1][8]/P0001 , \wishbone_tx_fifo_fifo_reg[1][9]/P0001 , \wishbone_tx_fifo_fifo_reg[2][0]/P0001 , \wishbone_tx_fifo_fifo_reg[2][10]/P0001 , \wishbone_tx_fifo_fifo_reg[2][11]/P0001 , \wishbone_tx_fifo_fifo_reg[2][12]/P0001 , \wishbone_tx_fifo_fifo_reg[2][13]/P0001 , \wishbone_tx_fifo_fifo_reg[2][14]/P0001 , \wishbone_tx_fifo_fifo_reg[2][15]/P0001 , \wishbone_tx_fifo_fifo_reg[2][16]/P0001 , \wishbone_tx_fifo_fifo_reg[2][17]/P0001 , \wishbone_tx_fifo_fifo_reg[2][18]/P0001 , \wishbone_tx_fifo_fifo_reg[2][19]/P0001 , \wishbone_tx_fifo_fifo_reg[2][1]/P0001 , \wishbone_tx_fifo_fifo_reg[2][20]/P0001 , \wishbone_tx_fifo_fifo_reg[2][21]/P0001 , \wishbone_tx_fifo_fifo_reg[2][22]/P0001 , \wishbone_tx_fifo_fifo_reg[2][23]/P0001 , \wishbone_tx_fifo_fifo_reg[2][24]/P0001 , \wishbone_tx_fifo_fifo_reg[2][25]/P0001 , \wishbone_tx_fifo_fifo_reg[2][26]/P0001 , \wishbone_tx_fifo_fifo_reg[2][27]/P0001 , \wishbone_tx_fifo_fifo_reg[2][28]/P0001 , \wishbone_tx_fifo_fifo_reg[2][29]/P0001 , \wishbone_tx_fifo_fifo_reg[2][2]/P0001 , \wishbone_tx_fifo_fifo_reg[2][30]/P0001 , \wishbone_tx_fifo_fifo_reg[2][31]/P0001 , \wishbone_tx_fifo_fifo_reg[2][3]/P0001 , \wishbone_tx_fifo_fifo_reg[2][4]/P0001 , \wishbone_tx_fifo_fifo_reg[2][5]/P0001 , \wishbone_tx_fifo_fifo_reg[2][6]/P0001 , \wishbone_tx_fifo_fifo_reg[2][7]/P0001 , \wishbone_tx_fifo_fifo_reg[2][8]/P0001 , \wishbone_tx_fifo_fifo_reg[2][9]/P0001 , \wishbone_tx_fifo_fifo_reg[3][0]/P0001 , \wishbone_tx_fifo_fifo_reg[3][10]/P0001 , \wishbone_tx_fifo_fifo_reg[3][11]/P0001 , \wishbone_tx_fifo_fifo_reg[3][12]/P0001 , \wishbone_tx_fifo_fifo_reg[3][13]/P0001 , \wishbone_tx_fifo_fifo_reg[3][14]/P0001 , \wishbone_tx_fifo_fifo_reg[3][15]/P0001 , \wishbone_tx_fifo_fifo_reg[3][16]/P0001 , \wishbone_tx_fifo_fifo_reg[3][17]/P0001 , \wishbone_tx_fifo_fifo_reg[3][18]/P0001 , \wishbone_tx_fifo_fifo_reg[3][19]/P0001 , \wishbone_tx_fifo_fifo_reg[3][1]/P0001 , \wishbone_tx_fifo_fifo_reg[3][20]/P0001 , \wishbone_tx_fifo_fifo_reg[3][21]/P0001 , \wishbone_tx_fifo_fifo_reg[3][22]/P0001 , \wishbone_tx_fifo_fifo_reg[3][23]/P0001 , \wishbone_tx_fifo_fifo_reg[3][24]/P0001 , \wishbone_tx_fifo_fifo_reg[3][25]/P0001 , \wishbone_tx_fifo_fifo_reg[3][26]/P0001 , \wishbone_tx_fifo_fifo_reg[3][27]/P0001 , \wishbone_tx_fifo_fifo_reg[3][28]/P0001 , \wishbone_tx_fifo_fifo_reg[3][29]/P0001 , \wishbone_tx_fifo_fifo_reg[3][2]/P0001 , \wishbone_tx_fifo_fifo_reg[3][30]/P0001 , \wishbone_tx_fifo_fifo_reg[3][31]/P0001 , \wishbone_tx_fifo_fifo_reg[3][3]/P0001 , \wishbone_tx_fifo_fifo_reg[3][4]/P0001 , \wishbone_tx_fifo_fifo_reg[3][5]/P0001 , \wishbone_tx_fifo_fifo_reg[3][6]/P0001 , \wishbone_tx_fifo_fifo_reg[3][7]/P0001 , \wishbone_tx_fifo_fifo_reg[3][8]/P0001 , \wishbone_tx_fifo_fifo_reg[3][9]/P0001 , \wishbone_tx_fifo_fifo_reg[4][0]/P0001 , \wishbone_tx_fifo_fifo_reg[4][10]/P0001 , \wishbone_tx_fifo_fifo_reg[4][11]/P0001 , \wishbone_tx_fifo_fifo_reg[4][12]/P0001 , \wishbone_tx_fifo_fifo_reg[4][13]/P0001 , \wishbone_tx_fifo_fifo_reg[4][14]/P0001 , \wishbone_tx_fifo_fifo_reg[4][15]/P0001 , \wishbone_tx_fifo_fifo_reg[4][16]/P0001 , \wishbone_tx_fifo_fifo_reg[4][17]/P0001 , \wishbone_tx_fifo_fifo_reg[4][18]/P0001 , \wishbone_tx_fifo_fifo_reg[4][19]/P0001 , \wishbone_tx_fifo_fifo_reg[4][1]/P0001 , \wishbone_tx_fifo_fifo_reg[4][20]/P0001 , \wishbone_tx_fifo_fifo_reg[4][21]/P0001 , \wishbone_tx_fifo_fifo_reg[4][22]/P0001 , \wishbone_tx_fifo_fifo_reg[4][23]/P0001 , \wishbone_tx_fifo_fifo_reg[4][24]/P0001 , \wishbone_tx_fifo_fifo_reg[4][25]/P0001 , \wishbone_tx_fifo_fifo_reg[4][26]/P0001 , \wishbone_tx_fifo_fifo_reg[4][27]/P0001 , \wishbone_tx_fifo_fifo_reg[4][28]/P0001 , \wishbone_tx_fifo_fifo_reg[4][29]/P0001 , \wishbone_tx_fifo_fifo_reg[4][2]/P0001 , \wishbone_tx_fifo_fifo_reg[4][30]/P0001 , \wishbone_tx_fifo_fifo_reg[4][31]/P0001 , \wishbone_tx_fifo_fifo_reg[4][3]/P0001 , \wishbone_tx_fifo_fifo_reg[4][4]/P0001 , \wishbone_tx_fifo_fifo_reg[4][5]/P0001 , \wishbone_tx_fifo_fifo_reg[4][6]/P0001 , \wishbone_tx_fifo_fifo_reg[4][7]/P0001 , \wishbone_tx_fifo_fifo_reg[4][8]/P0001 , \wishbone_tx_fifo_fifo_reg[4][9]/P0001 , \wishbone_tx_fifo_fifo_reg[5][0]/P0001 , \wishbone_tx_fifo_fifo_reg[5][10]/P0001 , \wishbone_tx_fifo_fifo_reg[5][11]/P0001 , \wishbone_tx_fifo_fifo_reg[5][12]/P0001 , \wishbone_tx_fifo_fifo_reg[5][13]/P0001 , \wishbone_tx_fifo_fifo_reg[5][14]/P0001 , \wishbone_tx_fifo_fifo_reg[5][15]/P0001 , \wishbone_tx_fifo_fifo_reg[5][16]/P0001 , \wishbone_tx_fifo_fifo_reg[5][17]/P0001 , \wishbone_tx_fifo_fifo_reg[5][18]/P0001 , \wishbone_tx_fifo_fifo_reg[5][19]/P0001 , \wishbone_tx_fifo_fifo_reg[5][1]/P0001 , \wishbone_tx_fifo_fifo_reg[5][20]/P0001 , \wishbone_tx_fifo_fifo_reg[5][21]/P0001 , \wishbone_tx_fifo_fifo_reg[5][22]/P0001 , \wishbone_tx_fifo_fifo_reg[5][23]/P0001 , \wishbone_tx_fifo_fifo_reg[5][24]/P0001 , \wishbone_tx_fifo_fifo_reg[5][25]/P0001 , \wishbone_tx_fifo_fifo_reg[5][26]/P0001 , \wishbone_tx_fifo_fifo_reg[5][27]/P0001 , \wishbone_tx_fifo_fifo_reg[5][28]/P0001 , \wishbone_tx_fifo_fifo_reg[5][29]/P0001 , \wishbone_tx_fifo_fifo_reg[5][2]/P0001 , \wishbone_tx_fifo_fifo_reg[5][30]/P0001 , \wishbone_tx_fifo_fifo_reg[5][31]/P0001 , \wishbone_tx_fifo_fifo_reg[5][3]/P0001 , \wishbone_tx_fifo_fifo_reg[5][4]/P0001 , \wishbone_tx_fifo_fifo_reg[5][5]/P0001 , \wishbone_tx_fifo_fifo_reg[5][6]/P0001 , \wishbone_tx_fifo_fifo_reg[5][7]/P0001 , \wishbone_tx_fifo_fifo_reg[5][8]/P0001 , \wishbone_tx_fifo_fifo_reg[5][9]/P0001 , \wishbone_tx_fifo_fifo_reg[6][0]/P0001 , \wishbone_tx_fifo_fifo_reg[6][10]/P0001 , \wishbone_tx_fifo_fifo_reg[6][11]/P0001 , \wishbone_tx_fifo_fifo_reg[6][12]/P0001 , \wishbone_tx_fifo_fifo_reg[6][13]/P0001 , \wishbone_tx_fifo_fifo_reg[6][14]/P0001 , \wishbone_tx_fifo_fifo_reg[6][15]/P0001 , \wishbone_tx_fifo_fifo_reg[6][16]/P0001 , \wishbone_tx_fifo_fifo_reg[6][17]/P0001 , \wishbone_tx_fifo_fifo_reg[6][18]/P0001 , \wishbone_tx_fifo_fifo_reg[6][19]/P0001 , \wishbone_tx_fifo_fifo_reg[6][1]/P0001 , \wishbone_tx_fifo_fifo_reg[6][20]/P0001 , \wishbone_tx_fifo_fifo_reg[6][21]/P0001 , \wishbone_tx_fifo_fifo_reg[6][22]/P0001 , \wishbone_tx_fifo_fifo_reg[6][23]/P0001 , \wishbone_tx_fifo_fifo_reg[6][24]/P0001 , \wishbone_tx_fifo_fifo_reg[6][25]/P0001 , \wishbone_tx_fifo_fifo_reg[6][26]/P0001 , \wishbone_tx_fifo_fifo_reg[6][27]/P0001 , \wishbone_tx_fifo_fifo_reg[6][28]/P0001 , \wishbone_tx_fifo_fifo_reg[6][29]/P0001 , \wishbone_tx_fifo_fifo_reg[6][2]/P0001 , \wishbone_tx_fifo_fifo_reg[6][30]/P0001 , \wishbone_tx_fifo_fifo_reg[6][31]/P0001 , \wishbone_tx_fifo_fifo_reg[6][3]/P0001 , \wishbone_tx_fifo_fifo_reg[6][4]/P0001 , \wishbone_tx_fifo_fifo_reg[6][5]/P0001 , \wishbone_tx_fifo_fifo_reg[6][6]/P0001 , \wishbone_tx_fifo_fifo_reg[6][7]/P0001 , \wishbone_tx_fifo_fifo_reg[6][8]/P0001 , \wishbone_tx_fifo_fifo_reg[6][9]/P0001 , \wishbone_tx_fifo_fifo_reg[7][0]/P0001 , \wishbone_tx_fifo_fifo_reg[7][10]/P0001 , \wishbone_tx_fifo_fifo_reg[7][11]/P0001 , \wishbone_tx_fifo_fifo_reg[7][12]/P0001 , \wishbone_tx_fifo_fifo_reg[7][13]/P0001 , \wishbone_tx_fifo_fifo_reg[7][14]/P0001 , \wishbone_tx_fifo_fifo_reg[7][15]/P0001 , \wishbone_tx_fifo_fifo_reg[7][16]/P0001 , \wishbone_tx_fifo_fifo_reg[7][17]/P0001 , \wishbone_tx_fifo_fifo_reg[7][18]/P0001 , \wishbone_tx_fifo_fifo_reg[7][19]/P0001 , \wishbone_tx_fifo_fifo_reg[7][1]/P0001 , \wishbone_tx_fifo_fifo_reg[7][20]/P0001 , \wishbone_tx_fifo_fifo_reg[7][21]/P0001 , \wishbone_tx_fifo_fifo_reg[7][22]/P0001 , \wishbone_tx_fifo_fifo_reg[7][23]/P0001 , \wishbone_tx_fifo_fifo_reg[7][24]/P0001 , \wishbone_tx_fifo_fifo_reg[7][25]/P0001 , \wishbone_tx_fifo_fifo_reg[7][26]/P0001 , \wishbone_tx_fifo_fifo_reg[7][27]/P0001 , \wishbone_tx_fifo_fifo_reg[7][28]/P0001 , \wishbone_tx_fifo_fifo_reg[7][29]/P0001 , \wishbone_tx_fifo_fifo_reg[7][2]/P0001 , \wishbone_tx_fifo_fifo_reg[7][30]/P0001 , \wishbone_tx_fifo_fifo_reg[7][31]/P0001 , \wishbone_tx_fifo_fifo_reg[7][3]/P0001 , \wishbone_tx_fifo_fifo_reg[7][4]/P0001 , \wishbone_tx_fifo_fifo_reg[7][5]/P0001 , \wishbone_tx_fifo_fifo_reg[7][6]/P0001 , \wishbone_tx_fifo_fifo_reg[7][7]/P0001 , \wishbone_tx_fifo_fifo_reg[7][8]/P0001 , \wishbone_tx_fifo_fifo_reg[7][9]/P0001 , \wishbone_tx_fifo_fifo_reg[8][0]/P0001 , \wishbone_tx_fifo_fifo_reg[8][10]/P0001 , \wishbone_tx_fifo_fifo_reg[8][11]/P0001 , \wishbone_tx_fifo_fifo_reg[8][12]/P0001 , \wishbone_tx_fifo_fifo_reg[8][13]/P0001 , \wishbone_tx_fifo_fifo_reg[8][14]/P0001 , \wishbone_tx_fifo_fifo_reg[8][15]/P0001 , \wishbone_tx_fifo_fifo_reg[8][16]/P0001 , \wishbone_tx_fifo_fifo_reg[8][17]/P0001 , \wishbone_tx_fifo_fifo_reg[8][18]/P0001 , \wishbone_tx_fifo_fifo_reg[8][19]/P0001 , \wishbone_tx_fifo_fifo_reg[8][1]/P0001 , \wishbone_tx_fifo_fifo_reg[8][20]/P0001 , \wishbone_tx_fifo_fifo_reg[8][21]/P0001 , \wishbone_tx_fifo_fifo_reg[8][22]/P0001 , \wishbone_tx_fifo_fifo_reg[8][23]/P0001 , \wishbone_tx_fifo_fifo_reg[8][24]/P0001 , \wishbone_tx_fifo_fifo_reg[8][25]/P0001 , \wishbone_tx_fifo_fifo_reg[8][26]/P0001 , \wishbone_tx_fifo_fifo_reg[8][27]/P0001 , \wishbone_tx_fifo_fifo_reg[8][28]/P0001 , \wishbone_tx_fifo_fifo_reg[8][29]/P0001 , \wishbone_tx_fifo_fifo_reg[8][2]/P0001 , \wishbone_tx_fifo_fifo_reg[8][30]/P0001 , \wishbone_tx_fifo_fifo_reg[8][31]/P0001 , \wishbone_tx_fifo_fifo_reg[8][3]/P0001 , \wishbone_tx_fifo_fifo_reg[8][4]/P0001 , \wishbone_tx_fifo_fifo_reg[8][5]/P0001 , \wishbone_tx_fifo_fifo_reg[8][6]/P0001 , \wishbone_tx_fifo_fifo_reg[8][7]/P0001 , \wishbone_tx_fifo_fifo_reg[8][8]/P0001 , \wishbone_tx_fifo_fifo_reg[8][9]/P0001 , \wishbone_tx_fifo_fifo_reg[9][0]/P0001 , \wishbone_tx_fifo_fifo_reg[9][10]/P0001 , \wishbone_tx_fifo_fifo_reg[9][11]/P0001 , \wishbone_tx_fifo_fifo_reg[9][12]/P0001 , \wishbone_tx_fifo_fifo_reg[9][13]/P0001 , \wishbone_tx_fifo_fifo_reg[9][14]/P0001 , \wishbone_tx_fifo_fifo_reg[9][15]/P0001 , \wishbone_tx_fifo_fifo_reg[9][16]/P0001 , \wishbone_tx_fifo_fifo_reg[9][17]/P0001 , \wishbone_tx_fifo_fifo_reg[9][18]/P0001 , \wishbone_tx_fifo_fifo_reg[9][19]/P0001 , \wishbone_tx_fifo_fifo_reg[9][1]/P0001 , \wishbone_tx_fifo_fifo_reg[9][20]/P0001 , \wishbone_tx_fifo_fifo_reg[9][21]/P0001 , \wishbone_tx_fifo_fifo_reg[9][22]/P0001 , \wishbone_tx_fifo_fifo_reg[9][23]/P0001 , \wishbone_tx_fifo_fifo_reg[9][24]/P0001 , \wishbone_tx_fifo_fifo_reg[9][25]/P0001 , \wishbone_tx_fifo_fifo_reg[9][26]/P0001 , \wishbone_tx_fifo_fifo_reg[9][27]/P0001 , \wishbone_tx_fifo_fifo_reg[9][28]/P0001 , \wishbone_tx_fifo_fifo_reg[9][29]/P0001 , \wishbone_tx_fifo_fifo_reg[9][2]/P0001 , \wishbone_tx_fifo_fifo_reg[9][30]/P0001 , \wishbone_tx_fifo_fifo_reg[9][31]/P0001 , \wishbone_tx_fifo_fifo_reg[9][3]/P0001 , \wishbone_tx_fifo_fifo_reg[9][4]/P0001 , \wishbone_tx_fifo_fifo_reg[9][5]/P0001 , \wishbone_tx_fifo_fifo_reg[9][6]/P0001 , \wishbone_tx_fifo_fifo_reg[9][7]/P0001 , \wishbone_tx_fifo_fifo_reg[9][8]/P0001 , \wishbone_tx_fifo_fifo_reg[9][9]/P0001 , \wishbone_tx_fifo_read_pointer_reg[0]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[1]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[2]/NET0131 , \wishbone_tx_fifo_read_pointer_reg[3]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[0]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[1]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[2]/NET0131 , \wishbone_tx_fifo_write_pointer_reg[3]/NET0131 , \_al_n1 , \g215539/_0_ , \g215543/_0_ , \g215547/_0_ , \g215551/_0_ , \g215552/_0_ , \g215578/_0_ , \g215587/_1_ , \g215589/_1_ , \g215591/_1_ , \g215593/_1_ , \g215595/_1_ , \g215597/_1_ , \g215599/_1_ , \g215601/_1_ , \g215603/_1_ , \g215605/_1_ , \g215607/_1_ , \g215609/_1_ , \g215611/_1_ , \g215613/_1_ , \g215615/_1_ , \g215617/_1_ , \g215618/_0_ , \g215619/_0_ , \g215620/_0_ , \g215632/_1_ , \g215634/_0_ , \g215635/_0_ , \g215636/_0_ , \g215637/_0_ , \g215638/_0_ , \g215639/_0_ , \g215655/_1_ , \g215657/_1_ , \g215659/_1_ , \g215661/_1_ , \g215662/_0_ , \g215663/_0_ , \g215664/_0_ , \g215665/_0_ , \g215668/_0_ , \g215674/_0_ , \g215677/_0_ , \g215686/_0_ , \g215695/_0_ , \g215696/_0_ , \g215702/_1__syn_2 , \g215705/_0_ , \g215706/_0_ , \g215716/_0_ , \g215717/_0_ , \g215718/_0_ , \g215726/_0_ , \g215727/_0_ , \g215728/_0_ , \g215760/_0_ , \g215764/_0_ , \g215765/_0_ , \g215766/_0_ , \g215767/_3_ , \g215768/_3_ , \g215769/_3_ , \g215770/_3_ , \g215771/_3_ , \g215772/_3_ , \g215773/_3_ , \g215774/_3_ , \g215775/_3_ , \g215776/_3_ , \g215777/_3_ , \g215778/_3_ , \g215779/_3_ , \g215780/_3_ , \g215790/_0_ , \g215791/_0_ , \g215792/_0_ , \g215793/_0_ , \g215801/_0_ , \g215802/_0_ , \g215803/_0_ , \g215804/_0_ , \g215812/_0_ , \g215813/_0_ , \g215821/_0_ , \g215823/_0_ , \g215831/_0_ , \g215832/_0_ , \g215833/_0_ , \g215845/_0_ , \g215846/_0_ , \g215847/_0_ , \g215872/_0_ , \g215873/_0_ , \g215874/_0_ , \g215904/_0_ , \g215905/_0_ , \g215906/_0_ , \g215907/_0_ , \g215908/_0_ , \g215909/_0_ , \g215910/_0_ , \g215911/_0_ , \g215912/_0_ , \g215913/_0_ , \g215914/_0_ , \g215915/_0_ , \g215916/_0_ , \g215917/_0_ , \g215918/_0_ , \g215919/_0_ , \g215920/_0_ , \g215923/_0_ , \g215926/_0_ , \g215941/_0_ , \g215942/_0_ , \g215943/_0_ , \g215944/_0_ , \g215945/_0_ , \g215946/_0_ , \g215947/_0_ , \g215948/_0_ , \g215949/_0_ , \g215950/_0_ , \g215951/_0_ , \g215952/_0_ , \g215953/_0_ , \g215954/_0_ , \g215955/_0_ , \g215956/_0_ , \g215957/_0_ , \g215959/_00_ , \g215960/_0_ , \g215962/_0_ , \g215964/_0_ , \g215966/_0_ , \g215972/_0_ , \g216035/_0_ , \g216037/_0_ , \g216038/_0_ , \g216039/_0_ , \g216040/_0_ , \g216041/_0_ , \g216042/_0_ , \g216046/_0_ , \g216048/_0_ , \g216057/_0_ , \g216263/_0_ , \g216264/_0_ , \g216265/_0_ , \g216266/_0_ , \g216267/_0_ , \g216268/_0_ , \g216269/_0_ , \g216270/_0_ , \g216271/_0_ , \g216272/_0_ , \g216273/_0_ , \g216284/_0_ , \g216289/_0_ , \g216290/_0_ , \g216292/_0_ , \g216296/_0_ , \g216297/_0_ , \g216300/_0_ , \g216301/_0_ , \g216302/_0_ , \g216303/_0_ , \g216304/_0_ , \g216305/_0_ , \g216306/_0_ , \g216307/_0_ , \g216310/_3_ , \g216311/_3_ , \g216314/u3_syn_7 , \g216322/_3_ , \g216323/_3_ , \g216324/_3_ , \g216325/_3_ , \g216326/_3_ , \g216327/_3_ , \g216328/_3_ , \g216329/_3_ , \g216369/_0_ , \g216370/_0_ , \g216371/_0_ , \g216372/_0_ , \g216373/_0_ , \g216374/_0_ , \g216375/_0_ , \g216376/_0_ , \g216379/_0_ , \g216380/_0_ , \g216381/_0_ , \g216385/_0_ , \g216389/_0_ , \g216390/_0_ , \g216402/_0_ , \g216404/_0_ , \g216405/_0_ , \g216406/_0_ , \g216407/_0_ , \g216408/_0_ , \g216409/_0_ , \g216410/_0_ , \g216411/_0_ , \g216412/_0_ , \g216413/_0_ , \g216414/_0_ , \g216415/_0_ , \g216416/_0_ , \g216417/_0_ , \g216418/_0_ , \g216419/_0_ , \g216420/_0_ , \g216421/_0_ , \g216422/_0_ , \g216423/_0_ , \g216424/_0_ , \g216425/_0_ , \g216426/_0_ , \g216427/_0_ , \g216428/_0_ , \g216429/_0_ , \g216430/_0_ , \g216431/_0_ , \g216432/_0_ , \g216433/_0_ , \g216434/_0_ , \g216435/_0_ , \g216436/_0_ , \g216437/_0_ , \g216438/_0_ , \g216439/_3_ , \g216447/_3_ , \g216448/_3_ , \g216452/_0_ , \g216453/_0_ , \g216454/_0_ , \g216455/_0_ , \g216456/_0_ , \g216457/_0_ , \g216458/_3_ , \g216459/_3_ , \g216461/_3_ , \g216462/_3_ , \g216463/_3_ , \g216464/_3_ , \g216465/_3_ , \g216466/_0_ , \g216467/_3_ , \g216468/_3_ , \g216469/_3_ , \g216470/_3_ , \g216471/_3_ , \g216473/_3_ , \g216474/_3_ , \g216475/_3_ , \g216476/_3_ , \g216477/_3_ , \g216478/_0_ , \g216479/_3_ , \g216480/_3_ , \g216481/_3_ , \g216492/_0_ , \g216494/_0_ , \g216495/_3_ , \g216496/_3_ , \g216498/_3_ , \g216499/_3_ , \g216500/_3_ , \g216513/_3_ , \g216514/_3_ , \g216515/_3_ , \g216516/_3_ , \g216517/_3_ , \g216518/_3_ , \g216519/_3_ , \g216520/_3_ , \g216521/_3_ , \g216522/_3_ , \g216523/_3_ , \g216524/_3_ , \g216525/_3_ , \g216526/_3_ , \g216527/_3_ , \g216528/_3_ , \g216529/_3_ , \g216530/_3_ , \g216531/_3_ , \g216532/_3_ , \g216533/_3_ , \g216534/_3_ , \g216535/_3_ , \g216536/_3_ , \g216537/_3_ , \g216538/_3_ , \g216555/_3_ , \g216556/_3_ , \g216557/_3_ , \g216560/_3_ , \g216561/_3_ , \g216562/_3_ , \g216563/_3_ , \g216564/_3_ , \g216565/_3_ , \g216566/_3_ , \g216567/_3_ , \g216568/_3_ , \g216569/_3_ , \g216570/_3_ , \g216571/_3_ , \g216575/_3_ , \g216576/_3_ , \g216577/_3_ , \g216578/_3_ , \g216579/_3_ , \g216580/_3_ , \g216581/_3_ , \g216582/_3_ , \g216583/_3_ , \g216586/_3_ , \g216587/_3_ , \g216588/_3_ , \g216589/_3_ , \g216590/_3_ , \g216591/_3_ , \g216592/_3_ , \g216593/_3_ , \g216594/_3_ , \g216595/_3_ , \g216600/_3_ , \g216683/_0_ , \g216689/_0_ , \g216693/_0_ , \g216694/_0_ , \g216727/_0_ , \g216728/_0_ , \g216729/_0_ , \g216732/_0_ , \g216733/_0_ , \g216734/_0_ , \g216735/_0_ , \g216736/_0_ , \g216737/_0_ , \g216738/_0_ , \g216739/_0_ , \g216740/_0_ , \g216741/_0_ , \g216742/_0_ , \g216743/_0_ , \g216744/_0_ , \g216745/_0_ , \g216746/_0_ , \g216748/_0_ , \g216751/_0_ , \g216754/_0_ , \g216762/_0_ , \g216934/_2_ , \g216952/_0_ , \g216955/_0_ , \g216969/_0_ , \g216979/_0_ , \g216984/_0_ , \g216996/_0_ , \g217002/_0_ , \g217014/_0_ , \g217015/_0_ , \g217016/_0_ , \g217017/_0_ , \g217018/_0_ , \g217019/_0_ , \g217023/_0_ , \g217116/_0_ , \g217146/_3_ , \g217149/_0_ , \g217151/_0_ , \g217160/_0_ , \g217167/_0_ , \g217168/_0_ , \g217169/_0_ , \g217170/_0_ , \g217171/_0_ , \g217172/_0_ , \g217173/_0_ , \g217174/_0_ , \g217175/_0_ , \g217176/_0_ , \g217177/_0_ , \g217178/_0_ , \g217179/_0_ , \g217180/_0_ , \g217181/_0_ , \g217182/_0_ , \g217183/_0_ , \g217187/_0_ , \g217188/_0_ , \g217189/_0_ , \g217193/_0_ , \g217194/_0_ , \g217195/_0_ , \g217196/_0_ , \g217202/_0_ , \g217205/_0_ , \g217206/_0_ , \g217207/_0_ , \g217208/_0_ , \g217209/_0_ , \g217210/_0_ , \g217211/_0_ , \g217212/_0_ , \g217213/_0_ , \g217214/_0_ , \g217215/_0_ , \g217216/_0_ , \g217217/_0_ , \g217218/_0_ , \g217219/_0_ , \g217220/_0_ , \g217223/_0_ , \g217231/_0_ , \g217237/_0_ , \g217238/_0_ , \g217242/_0_ , \g217243/_0_ , \g217250/_3_ , \g217251/_3_ , \g217252/_3_ , \g217253/_3_ , \g217254/_3_ , \g217255/_3_ , \g217256/_3_ , \g217257/_3_ , \g217258/_3_ , \g217259/_3_ , \g217260/_3_ , \g217261/_3_ , \g217262/_3_ , \g217263/_3_ , \g217264/_3_ , \g217265/_3_ , \g217266/_3_ , \g217267/_3_ , \g217268/_3_ , \g217269/_3_ , \g217270/_3_ , \g217271/_3_ , \g217272/_3_ , \g217273/_3_ , \g217274/_3_ , \g217275/_3_ , \g217276/_3_ , \g217277/_3_ , \g217278/_3_ , \g217279/_3_ , \g217280/_3_ , \g217281/_3_ , \g217282/_3_ , \g217283/_3_ , \g217284/_3_ , \g217285/_3_ , \g217286/_3_ , \g217287/_3_ , \g217288/_3_ , \g217289/_3_ , \g217290/_3_ , \g217291/_3_ , \g217292/_3_ , \g217293/_3_ , \g217294/_3_ , \g217295/_3_ , \g217296/_3_ , \g217297/_3_ , \g217298/_3_ , \g217299/_3_ , \g217300/_3_ , \g217301/_3_ , \g217302/_3_ , \g217303/_3_ , \g217304/_3_ , \g217305/_3_ , \g217306/_3_ , \g217307/_3_ , \g217308/_3_ , \g217309/_3_ , \g217310/_3_ , \g217311/_3_ , \g217312/_3_ , \g217313/_3_ , \g217318/_0_ , \g217662/_0_ , \g217663/_0_ , \g217682/_0_ , \g217697/_0_ , \g217698/_0_ , \g217699/_0_ , \g217700/_0_ , \g217701/_0_ , \g217705/_0_ , \g217711/_0_ , \g217747/_0_ , \g217753/_00_ , \g217775/_0_ , \g217781/_0_ , \g217784/_0_ , \g217785/_0_ , \g217786/_0_ , \g217787/_0_ , \g217788/_0_ , \g217790/_0_ , \g217815/_0_ , \g217817/_0_ , \g218145/_0_ , \g218148/_0_ , \g218150/_0_ , \g218167/_0_ , \g218168/_0_ , \g218234/_0_ , \g218235/_0_ , \g218236/_0_ , \g218238/_0_ , \g218242/_0_ , \g218332/_0_ , \g218335/_0_ , \g218336/_0_ , \g218337/_0_ , \g218338/_0_ , \g218339/_0_ , \g218340/_0_ , \g218341/_0_ , \g218342/_0_ , \g218343/_0_ , \g218344/_0_ , \g218345/_0_ , \g218346/_0_ , \g218347/_0_ , \g218348/_0_ , \g218349/_0_ , \g218350/_0_ , \g218351/_0_ , \g218352/_0_ , \g218353/_0_ , \g218354/_0_ , \g218355/_0_ , \g218356/_0_ , \g218357/_0_ , \g218358/_0_ , \g218359/_0_ , \g218360/_0_ , \g218398/_3_ , \g218430/_0_ , \g218440/_0_ , \g218452/u3_syn_4 , \g218495/u3_syn_4 , \g218517/u3_syn_4 , \g218554/u3_syn_4 , \g218575/u3_syn_4 , \g218600/u3_syn_4 , \g218621/u3_syn_4 , \g218638/u3_syn_4 , \g218659/u3_syn_4 , \g218673/u3_syn_4 , \g218707/u3_syn_4 , \g218735/_3_ , \g219186/_0_ , \g219187/_0_ , \g219188/_0_ , \g219189/_0_ , \g219190/_0_ , \g219196/_0_ , \g219198/_0_ , \g219199/_0_ , \g219200/_0_ , \g219308/_0_ , \g219314/_0_ , \g219326/_0_ , \g219328/_0_ , \g219348/_0_ , \g219351/_0_ , \g219363/_0_ , \g219364/_0_ , \g219365/_0_ , \g219366/_0_ , \g219367/_0_ , \g219368/_0_ , \g219369/_0_ , \g219376/_0_ , \g219381/_0_ , \g219382/_0_ , \g219384/_0_ , \g219385/_0_ , \g219391/_0_ , \g219394/_0_ , \g219395/_0_ , \g219396/_0_ , \g219397/_0_ , \g219398/_0_ , \g219399/_0_ , \g219400/_0_ , \g219401/_0_ , \g219402/_0_ , \g219403/_0_ , \g219404/_0_ , \g219405/_0_ , \g219406/_0_ , \g219407/_0_ , \g219408/_0_ , \g219409/_0_ , \g219410/_0_ , \g219411/_0_ , \g219412/_0_ , \g219413/_0_ , \g219414/_0_ , \g219415/_0_ , \g219416/_0_ , \g219417/_0_ , \g219418/_0_ , \g219419/_0_ , \g219420/_0_ , \g219421/_0_ , \g219422/_0_ , \g219423/_0_ , \g219424/_0_ , \g219425/_0_ , \g219426/_0_ , \g219427/_0_ , \g219428/_0_ , \g219429/_0_ , \g219430/_0_ , \g219431/_0_ , \g219432/_0_ , \g219433/_0_ , \g219434/_0_ , \g219435/_0_ , \g219436/_0_ , \g219437/_0_ , \g219438/_0_ , \g219439/_0_ , \g219440/_0_ , \g219441/_0_ , \g219442/_0_ , \g219443/_0_ , \g219444/_0_ , \g219445/_0_ , \g219446/_0_ , \g219447/_0_ , \g219449/_0_ , \g219450/_0_ , \g219451/_0_ , \g219452/_0_ , \g219453/_0_ , \g219454/_0_ , \g219455/_0_ , \g219456/_0_ , \g219457/_0_ , \g219458/_0_ , \g219464/u3_syn_7 , \g219496/u3_syn_4 , \g219512/u3_syn_4 , \g219526/u3_syn_4 , \g219549/u3_syn_4 , \g219571/u3_syn_4 , \g219588/u3_syn_4 , \g219603/u3_syn_4 , \g219621/u3_syn_4 , \g219636/_3_ , \g219652/u3_syn_4 , \g219676/_3_ , \g219686/_0_ , \g219689/_0_ , \g219694/_3_ , \g220062/_0_ , \g220068/_0_ , \g220069/_0_ , \g220072/_0_ , \g220084/_0_ , \g220149/_0_ , \g220162/_0_ , \g220317/_0_ , \g220360/_2_ , \g220368/_2_ , \g220369/_0_ , \g220370/_0_ , \g220371/_0_ , \g220372/_0_ , \g220376/_0_ , \g220390/_0_ , \g220395/_0_ , \g220499/_0_ , \g220500/_0_ , \g220501/_0_ , \g220502/_0_ , \g220503/_0_ , \g220504/_0_ , \g220505/_0_ , \g220506/_0_ , \g220507/_0_ , \g220508/_0_ , \g220509/_0_ , \g220510/_0_ , \g220511/_0_ , \g220512/_0_ , \g220513/_0_ , \g220514/_0_ , \g220515/_0_ , \g220516/_0_ , \g220517/_0_ , \g220518/_0_ , \g220519/_0_ , \g220520/_0_ , \g220521/_0_ , \g220522/_0_ , \g220523/_0_ , \g220524/_0_ , \g220525/_0_ , \g220526/_0_ , \g220527/_0_ , \g220528/_0_ , \g220529/_0_ , \g220530/_0_ , \g220531/_0_ , \g220532/_0_ , \g220533/_0_ , \g220534/_0_ , \g220535/_0_ , \g220557/_0_ , \g220558/_0_ , \g220559/_0_ , \g220560/_0_ , \g220561/_0_ , \g220562/_0_ , \g220563/_0_ , \g220564/_0_ , \g220565/_0_ , \g220566/_0_ , \g220567/_0_ , \g220568/_0_ , \g220569/_0_ , \g220570/_0_ , \g220571/_0_ , \g220572/_0_ , \g220573/_0_ , \g220574/_0_ , \g220575/_0_ , \g220576/_0_ , \g220577/_0_ , \g220578/_0_ , \g220579/_0_ , \g220580/_0_ , \g220581/_0_ , \g220582/_0_ , \g220583/_0_ , \g220584/_0_ , \g220585/_0_ , \g220586/_0_ , \g220587/_0_ , \g220588/_0_ , \g220589/_0_ , \g220590/_0_ , \g220591/_0_ , \g220592/_0_ , \g220593/_0_ , \g220594/_0_ , \g220595/_0_ , \g220596/_0_ , \g220597/_0_ , \g220598/_0_ , \g220599/_0_ , \g220600/_0_ , \g220601/_0_ , \g220602/_0_ , \g220603/_0_ , \g220604/_0_ , \g220605/_0_ , \g220606/_0_ , \g220607/_0_ , \g220608/_0_ , \g220609/_0_ , \g220610/_0_ , \g220611/_0_ , \g220612/_0_ , \g220613/_0_ , \g220614/_0_ , \g220615/_0_ , \g220616/_0_ , \g220617/_0_ , \g220618/_0_ , \g220619/_0_ , \g220620/_0_ , \g220621/_0_ , \g220622/_0_ , \g220623/_0_ , \g220624/_0_ , \g220625/_0_ , \g220626/_0_ , \g220627/_0_ , \g220628/_0_ , \g220629/_0_ , \g220630/_0_ , \g220631/_0_ , \g220632/_0_ , \g220633/_0_ , \g220634/_0_ , \g220635/_0_ , \g220636/_0_ , \g220637/_0_ , \g220638/_0_ , \g220639/_0_ , \g220640/_0_ , \g220641/_0_ , \g220642/_0_ , \g220643/_0_ , \g220644/_0_ , \g220645/_0_ , \g220646/_0_ , \g220647/_0_ , \g220648/_0_ , \g220649/_0_ , \g220650/_0_ , \g220651/_0_ , \g220652/_0_ , \g220653/_0_ , \g220654/_0_ , \g220655/_0_ , \g220656/_0_ , \g220657/_0_ , \g220658/_0_ , \g220659/_0_ , \g220660/_0_ , \g220661/_0_ , \g220662/_0_ , \g220663/_0_ , \g220664/_0_ , \g220665/_0_ , \g220666/_0_ , \g220674/_0_ , \g220679/u3_syn_7 , \g220711/u3_syn_4 , \g220726/u3_syn_4 , \g220739/u3_syn_4 , \g220751/u3_syn_4 , \g220759/u3_syn_4 , \g220773/u3_syn_4 , \g220782/u3_syn_4 , \g220805/u3_syn_4 , \g220828/u3_syn_4 , \g220921/_0_ , \g220930/u3_syn_4 , \g220949/_3_ , \g220994/_3_ , \g221207/_0_ , \g221213/_0_ , \g221223/_0_ , \g221224/_0_ , \g221225/_0_ , \g221226/_0_ , \g221231/_0_ , \g221232/_0_ , \g221234/_0_ , \g221235/_0_ , \g221246/_2_ , \g221249/_2_ , \g221265/_0_ , \g221287/_0_ , \g221325/_0_ , \g221326/_0_ , \g221447/_0_ , \g221449/_0_ , \g221452/_0_ , \g221469/_0_ , \g221473/_0_ , \g221503/_0_ , \g221510/_0_ , \g221512/_0_ , \g221516/_0_ , \g221517/_0_ , \g221524/_0_ , \g221530/_0_ , \g221592/_0_ , \g221593/_0_ , \g221634/u3_syn_4 , \g221669/u3_syn_4 , \g221789/u3_syn_4 , \g221813/u3_syn_4 , \g221829/u3_syn_4 , \g221861/u3_syn_4 , \g221876/_0_ , \g221935/_0_ , \g221944/_3_ , \g230200/_0_ , \g230201/_0_ , \g230205/_0_ , \g230295/_0_ , \g230297/_0_ , \g230298/_0_ , \g230300/_0_ , \g230302/_0_ , \g230303/_0_ , \g230343/_0_ , \g230368/_0_ , \g230511/_0_ , \g230531/_0_ , \g230635/_2_ , \g230661/_0_ , \g230715/_1__syn_2 , \g230731/_0_ , \g230766/_0_ , \g230784/_0_ , \g230785/_0_ , \g230786/_0_ , \g230787/_0_ , \g230797/_0_ , \g230798/_0_ , \g230803/_0_ , \g230804/_00_ , \g230805/_00_ , \g230806/_00_ , \g230807/_00_ , \g230808/_00_ , \g230809/_00_ , \g230815/_0_ , \g230816/_2_ , \g230817/_2_ , \g230829/_0_ , \g230834/_0_ , \g230835/_0_ , \g230836/_0_ , \g230837/_0_ , \g230844/_0_ , \g230863/_3_ , \g230864/_3_ , \g230870/_0_ , \g230988/_3_ , \g231010/_3_ , \g231016/_3_ , \g231042/_3_ , \g231471/_0_ , \g231472/_0_ , \g231476/_3_ , \g231480/_3_ , \g231484/_3_ , \g231504/_0_ , \g231532/_0_ , \g231542/_0_ , \g231560/_1_ , \g231578/_1_ , \g231580/_0_ , \g231590/_1__syn_2 , \g231615/_0_ , \g231623/_1_ , \g231634/_2_ , \g231635/_0_ , \g231638/_2_ , \g231640/_0_ , \g231653/_2_ , \g231787/_0_ , \g231931/_0_ , \g231939/_3_ , \g231940/_0_ , \g231951/_0_ , \g231955/_0_ , \g231956/_0_ , \g231959/_2_ , \g231960/_0_ , \g231964/_0_ , \g231965/_0_ , \g231975/_0_ , \g231986/_1_ , \g231987/_1_ , \g231989/_1_ , \g231990/_1_ , \g231991/_0_ , \g231992/_0_ , \g231995/_0_ , \g231998/_0_ , \g231999/_0_ , \g232002/_3_ , \g232035/u3_syn_4 , \g232038/u3_syn_4 , \g232046/u3_syn_4 , \g232054/u3_syn_4 , \g232062/u3_syn_4 , \g232070/u3_syn_4 , \g232078/u3_syn_4 , \g232079/u3_syn_4 , \g232087/u3_syn_4 , \g232096/u3_syn_4 , \g232104/u3_syn_4 , \g232112/u3_syn_4 , \g232120/u3_syn_4 , \g232128/u3_syn_4 , \g232136/u3_syn_4 , \g232144/u3_syn_4 , \g232152/u3_syn_4 , \g232161/u3_syn_4 , \g232169/u3_syn_4 , \g232177/u3_syn_4 , \g232185/u3_syn_4 , \g232186/u3_syn_4 , \g232194/u3_syn_4 , \g232202/u3_syn_4 , \g232210/u3_syn_4 , \g232218/u3_syn_4 , \g232226/u3_syn_4 , \g232234/u3_syn_4 , \g232242/u3_syn_4 , \g232251/u3_syn_4 , \g232259/u3_syn_4 , \g232267/u3_syn_4 , \g232275/u3_syn_4 , \g232283/u3_syn_4 , \g232291/u3_syn_4 , \g232299/u3_syn_4 , \g232307/u3_syn_4 , \g232315/u3_syn_4 , \g232324/u3_syn_4 , \g232332/u3_syn_4 , \g232341/u3_syn_4 , \g232349/u3_syn_4 , \g232357/u3_syn_4 , \g232366/u3_syn_4 , \g232374/u3_syn_4 , \g232382/u3_syn_4 , \g232390/u3_syn_4 , \g232398/u3_syn_4 , \g232406/u3_syn_4 , \g232414/u3_syn_4 , \g232422/u3_syn_4 , \g232427/u3_syn_4 , \g232431/u3_syn_4 , \g232439/u3_syn_4 , \g232444/u3_syn_4 , \g232452/u3_syn_4 , \g232461/u3_syn_4 , \g232471/u3_syn_4 , \g232479/u3_syn_4 , \g232487/u3_syn_4 , \g232495/u3_syn_4 , \g232503/u3_syn_4 , \g232506/u3_syn_4 , \g232514/u3_syn_4 , \g232527/u3_syn_4 , \g232530/u3_syn_4 , \g232536/u3_syn_4 , \g232544/u3_syn_4 , \g232551/u3_syn_4 , \g232557/u3_syn_4 , \g232568/u3_syn_4 , \g232576/u3_syn_4 , \g232585/u3_syn_4 , \g232593/u3_syn_4 , \g232597/u3_syn_4 , \g232609/u3_syn_4 , \g232617/u3_syn_4 , \g232625/u3_syn_4 , \g232633/u3_syn_4 , \g232641/u3_syn_4 , \g232649/u3_syn_4 , \g232657/u3_syn_4 , \g232665/u3_syn_4 , \g232673/u3_syn_4 , \g232681/u3_syn_4 , \g232689/u3_syn_4 , \g232697/u3_syn_4 , \g232705/u3_syn_4 , \g232713/u3_syn_4 , \g232717/u3_syn_4 , \g232729/u3_syn_4 , \g232737/u3_syn_4 , \g232745/u3_syn_4 , \g232749/u3_syn_4 , \g232761/u3_syn_4 , \g232768/u3_syn_4 , \g232777/u3_syn_4 , \g232785/u3_syn_4 , \g232793/u3_syn_4 , \g232801/u3_syn_4 , \g232809/u3_syn_4 , \g232815/u3_syn_4 , \g232823/u3_syn_4 , \g232833/u3_syn_4 , \g232841/u3_syn_4 , \g232846/u3_syn_4 , \g232851/u3_syn_4 , \g232865/u3_syn_4 , \g232873/u3_syn_4 , \g232881/u3_syn_4 , \g232882/u3_syn_4 , \g232895/u3_syn_4 , \g232904/u3_syn_4 , \g232913/u3_syn_4 , \g232921/u3_syn_4 , \g232928/u3_syn_4 , \g232934/u3_syn_4 , \g232945/u3_syn_4 , \g232953/u3_syn_4 , \g232954/u3_syn_4 , \g232969/u3_syn_4 , \g232977/u3_syn_4 , \g232981/u3_syn_4 , \g232993/u3_syn_4 , \g232995/u3_syn_4 , \g233009/u3_syn_4 , \g233017/u3_syn_4 , \g233025/u3_syn_4 , \g233033/u3_syn_4 , \g233041/u3_syn_4 , \g233047/u3_syn_4 , \g233057/u3_syn_4 , \g233065/u3_syn_4 , \g233073/u3_syn_4 , \g233081/u3_syn_4 , \g233087/u3_syn_4 , \g233097/u3_syn_4 , \g233105/u3_syn_4 , \g233113/u3_syn_4 , \g233121/u3_syn_4 , \g233128/u3_syn_4 , \g233134/u3_syn_4 , \g233144/u3_syn_4 , \g233153/u3_syn_4 , \g233161/u3_syn_4 , \g233169/u3_syn_4 , \g233177/u3_syn_4 , \g233185/u3_syn_4 , \g233193/u3_syn_4 , \g233201/u3_syn_4 , \g233209/u3_syn_4 , \g233217/u3_syn_4 , \g233219/u3_syn_4 , \g233229/u3_syn_4 , \g233241/u3_syn_4 , \g233249/u3_syn_4 , \g233257/u3_syn_4 , \g233265/u3_syn_4 , \g233273/u3_syn_4 , \g233281/u3_syn_4 , \g233289/u3_syn_4 , \g233297/u3_syn_4 , \g233305/u3_syn_4 , \g233313/u3_syn_4 , \g233321/u3_syn_4 , \g233329/u3_syn_4 , \g233337/u3_syn_4 , \g233345/u3_syn_4 , \g233353/u3_syn_4 , \g233361/u3_syn_4 , \g233369/u3_syn_4 , \g233377/u3_syn_4 , \g233382/u3_syn_4 , \g233392/u3_syn_4 , \g233394/u3_syn_4 , \g233409/u3_syn_4 , \g233417/u3_syn_4 , \g233425/u3_syn_4 , \g233433/u3_syn_4 , \g233441/u3_syn_4 , \g233449/u3_syn_4 , \g233453/u3_syn_4 , \g233465/u3_syn_4 , \g233473/u3_syn_4 , \g233481/u3_syn_4 , \g233489/u3_syn_4 , \g233497/u3_syn_4 , \g233505/u3_syn_4 , \g233513/u3_syn_4 , \g233516/u3_syn_4 , \g233529/u3_syn_4 , \g233531/u3_syn_4 , \g233546/u3_syn_4 , \g233554/u3_syn_4 , \g233562/u3_syn_4 , \g233570/u3_syn_4 , \g233578/u3_syn_4 , \g233586/u3_syn_4 , \g233594/u3_syn_4 , \g233602/u3_syn_4 , \g233603/u3_syn_4 , \g233618/u3_syn_4 , \g233626/u3_syn_4 , \g233634/u3_syn_4 , \g233642/u3_syn_4 , \g233650/u3_syn_4 , \g233658/u3_syn_4 , \g233666/u3_syn_4 , \g233674/u3_syn_4 , \g233682/u3_syn_4 , \g233690/u3_syn_4 , \g233698/u3_syn_4 , \g233706/u3_syn_4 , \g233714/u3_syn_4 , \g233722/u3_syn_4 , \g233730/u3_syn_4 , \g233738/u3_syn_4 , \g233746/u3_syn_4 , \g233754/u3_syn_4 , \g233762/u3_syn_4 , \g233770/u3_syn_4 , \g233778/u3_syn_4 , \g233783/u3_syn_4 , \g233794/u3_syn_4 , \g233802/u3_syn_4 , \g233806/u3_syn_4 , \g233818/u3_syn_4 , \g233826/u3_syn_4 , \g233828/u3_syn_4 , \g233838/u3_syn_4 , \g233850/u3_syn_4 , \g233858/u3_syn_4 , \g233860/u3_syn_4 , \g233870/u3_syn_4 , \g233881/u3_syn_4 , \g233890/u3_syn_4 , \g233899/u3_syn_4 , \g233908/u3_syn_4 , \g233917/u3_syn_4 , \g233919/u3_syn_4 , \g233927/u3_syn_4 , \g233935/u3_syn_4 , \g233943/u3_syn_4 , \g233945/u3_syn_4 , \g233953/u3_syn_4 , \g233961/u3_syn_4 , \g233969/u3_syn_4 , \g233977/u3_syn_4 , \g233985/u3_syn_4 , \g233993/u3_syn_4 , \g234001/u3_syn_4 , \g234008/u3_syn_4 , \g234009/u3_syn_4 , \g234024/u3_syn_4 , \g234032/u3_syn_4 , \g234038/u3_syn_4 , \g234056/u3_syn_4 , \g234063/u3_syn_4 , \g234071/u3_syn_4 , \g234079/u3_syn_4 , \g234098/u3_syn_4 , \g234106/u3_syn_4 , \g234114/u3_syn_4 , \g234122/u3_syn_4 , \g234130/u3_syn_4 , \g234138/u3_syn_4 , \g234145/u3_syn_4 , \g234156/u3_syn_4 , \g234162/u3_syn_4 , \g234171/u3_syn_4 , \g234183/u3_syn_4 , \g234248/u3_syn_4 , \g234265/u3_syn_4 , \g234273/u3_syn_4 , \g234281/u3_syn_4 , \g234289/u3_syn_4 , \g234297/u3_syn_4 , \g234306/u3_syn_4 , \g234314/u3_syn_4 , \g234322/u3_syn_4 , \g234331/u3_syn_4 , \g234339/u3_syn_4 , \g234347/u3_syn_4 , \g234355/u3_syn_4 , \g234363/u3_syn_4 , \g234371/u3_syn_4 , \g234379/u3_syn_4 , \g234387/u3_syn_4 , \g234395/u3_syn_4 , \g234403/u3_syn_4 , \g234411/u3_syn_4 , \g234419/u3_syn_4 , \g234427/u3_syn_4 , \g234435/u3_syn_4 , \g234443/u3_syn_4 , \g234451/u3_syn_4 , \g234459/u3_syn_4 , \g234467/u3_syn_4 , \g234475/u3_syn_4 , \g234483/u3_syn_4 , \g234491/u3_syn_4 , \g234499/u3_syn_4 , \g234507/u3_syn_4 , \g234515/u3_syn_4 , \g234523/u3_syn_4 , \g234531/u3_syn_4 , \g234539/u3_syn_4 , \g234547/u3_syn_4 , \g234555/u3_syn_4 , \g234563/u3_syn_4 , \g234571/u3_syn_4 , \g234579/u3_syn_4 , \g234587/u3_syn_4 , \g234595/u3_syn_4 , \g234604/u3_syn_4 , \g234612/u3_syn_4 , \g234620/u3_syn_4 , \g234628/u3_syn_4 , \g234636/u3_syn_4 , \g234644/u3_syn_4 , \g234652/u3_syn_4 , \g234660/u3_syn_4 , \g234668/u3_syn_4 , \g234676/u3_syn_4 , \g234684/u3_syn_4 , \g234692/u3_syn_4 , \g234700/u3_syn_4 , \g234708/u3_syn_4 , \g234716/u3_syn_4 , \g234725/u3_syn_4 , \g234733/u3_syn_4 , \g234741/u3_syn_4 , \g234749/u3_syn_4 , \g234757/u3_syn_4 , \g234765/u3_syn_4 , \g234773/u3_syn_4 , \g234781/u3_syn_4 , \g234789/u3_syn_4 , \g234798/u3_syn_4 , \g234806/u3_syn_4 , \g234814/u3_syn_4 , \g234822/u3_syn_4 , \g234830/u3_syn_4 , \g234838/u3_syn_4 , \g235911/u3_syn_4 , \g235912/u3_syn_4 , \g235920/u3_syn_4 , \g235928/u3_syn_4 , \g235936/u3_syn_4 , \g235944/u3_syn_4 , \g235952/u3_syn_4 , \g235960/u3_syn_4 , \g235968/u3_syn_4 , \g235976/u3_syn_4 , \g235984/u3_syn_4 , \g235992/u3_syn_4 , \g236000/u3_syn_4 , \g236008/u3_syn_4 , \g236016/u3_syn_4 , \g236021/u3_syn_4 , \g236025/u3_syn_4 , \g236033/u3_syn_4 , \g236041/u3_syn_4 , \g236049/u3_syn_4 , \g236057/u3_syn_4 , \g236065/u3_syn_4 , \g236073/u3_syn_4 , \g236081/u3_syn_4 , \g236089/u3_syn_4 , \g236097/u3_syn_4 , \g236105/u3_syn_4 , \g236113/u3_syn_4 , \g236121/u3_syn_4 , \g236129/u3_syn_4 , \g236137/u3_syn_4 , \g236145/u3_syn_4 , \g236153/u3_syn_4 , \g236161/u3_syn_4 , \g236169/u3_syn_4 , \g236177/u3_syn_4 , \g236185/u3_syn_4 , \g236193/u3_syn_4 , \g236196/u3_syn_4 , \g236198/u3_syn_4 , \g236203/u3_syn_4 , \g236211/u3_syn_4 , \g236219/u3_syn_4 , \g236220/u3_syn_4 , \g236229/u3_syn_4 , \g236232/u3_syn_4 , \g236238/u3_syn_4 , \g236246/u3_syn_4 , \g236255/u3_syn_4 , \g236263/u3_syn_4 , \g236271/u3_syn_4 , \g236275/u3_syn_4 , \g236280/u3_syn_4 , \g236288/u3_syn_4 , \g236296/u3_syn_4 , \g236304/u3_syn_4 , \g236305/u3_syn_4 , \g236306/u3_syn_4 , \g236315/u3_syn_4 , \g236323/u3_syn_4 , \g236331/u3_syn_4 , \g236334/u3_syn_4 , \g236340/u3_syn_4 , \g236348/u3_syn_4 , \g236357/u3_syn_4 , \g236359/u3_syn_4 , \g236367/u3_syn_4 , \g236374/u3_syn_4 , \g236376/u3_syn_4 , \g236377/u3_syn_4 , \g236385/u3_syn_4 , \g236393/u3_syn_4 , \g236402/u3_syn_4 , \g236410/u3_syn_4 , \g236419/u3_syn_4 , \g236427/u3_syn_4 , \g236433/u3_syn_4 , \g236436/u3_syn_4 , \g236444/u3_syn_4 , \g236452/u3_syn_4 , \g236460/u3_syn_4 , \g236468/u3_syn_4 , \g236476/u3_syn_4 , \g236484/u3_syn_4 , \g236492/u3_syn_4 , \g236500/u3_syn_4 , \g236508/u3_syn_4 , \g236516/u3_syn_4 , \g236518/u3_syn_4 , \g236525/u3_syn_4 , \g236533/u3_syn_4 , \g236542/u3_syn_4 , \g236550/u3_syn_4 , \g236559/u3_syn_4 , \g236567/u3_syn_4 , \g236575/u3_syn_4 , \g236583/u3_syn_4 , \g236591/u3_syn_4 , \g236599/u3_syn_4 , \g236607/u3_syn_4 , \g236608/u3_syn_4 , \g236616/u3_syn_4 , \g236624/u3_syn_4 , \g236632/u3_syn_4 , \g236640/u3_syn_4 , \g236647/u3_syn_4 , \g236649/u3_syn_4 , \g236659/u3_syn_4 , \g236671/u3_syn_4 , \g236677/u3_syn_4 , \g236688/u3_syn_4 , \g236696/u3_syn_4 , \g236705/u3_syn_4 , \g236712/u3_syn_4 , \g236718/u3_syn_4 , \g236729/u3_syn_4 , \g236732/u3_syn_4 , \g236745/u3_syn_4 , \g236753/u3_syn_4 , \g236761/u3_syn_4 , \g236769/u3_syn_4 , \g236777/u3_syn_4 , \g236779/u3_syn_4 , \g236788/u3_syn_4 , \g236800/u3_syn_4 , \g236802/u3_syn_4 , \g236805/u3_syn_4 , \g236813/u3_syn_4 , \g236825/u3_syn_4 , \g236829/u3_syn_4 , \g236837/u3_syn_4 , \g236849/u3_syn_4 , \g236854/u3_syn_4 , \g236860/u3_syn_4 , \g236872/u3_syn_4 , \g236878/u3_syn_4 , \g236884/u3_syn_4 , \g236896/u3_syn_4 , \g236903/u3_syn_4 , \g236908/u3_syn_4 , \g236920/u3_syn_4 , \g236930/u3_syn_4 , \g236939/u3_syn_4 , \g236947/u3_syn_4 , \g236949/u3_syn_4 , \g236956/u3_syn_4 , \g236962/u3_syn_4 , \g236965/u3_syn_4 , \g236980/u3_syn_4 , \g236988/u3_syn_4 , \g236989/u3_syn_4 , \g237004/u3_syn_4 , \g237005/u3_syn_4 , \g237020/u3_syn_4 , \g237021/u3_syn_4 , \g237033/u3_syn_4 , \g237044/u3_syn_4 , \g237045/u3_syn_4 , \g237056/u3_syn_4 , \g237068/u3_syn_4 , \g237076/u3_syn_4 , \g237084/u3_syn_4 , \g237092/u3_syn_4 , \g237095/u3_syn_4 , \g237107/u3_syn_4 , \g237110/u3_syn_4 , \g237119/u3_syn_4 , \g237131/u3_syn_4 , \g237135/u3_syn_4 , \g237148/u3_syn_4 , \g237152/u3_syn_4 , \g237165/u3_syn_4 , \g237168/u3_syn_4 , \g237180/u3_syn_4 , \g237185/u3_syn_4 , \g237192/u3_syn_4 , \g237204/u3_syn_4 , \g237209/u3_syn_4 , \g237215/u3_syn_4 , \g237229/u3_syn_4 , \g237231/u3_syn_4 , \g237245/u3_syn_4 , \g237251/u3_syn_4 , \g237260/u3_syn_4 , \g237262/u3_syn_4 , \g237277/u3_syn_4 , \g237281/u3_syn_4 , \g237293/u3_syn_4 , \g237294/u3_syn_4 , \g237310/u3_syn_4 , \g237311/u3_syn_4 , \g237323/u3_syn_4 , \g237334/u3_syn_4 , \g237342/u3_syn_4 , \g237350/u3_syn_4 , \g237353/u3_syn_4 , \g237359/u3_syn_4 , \g237367/u3_syn_4 , \g237368/u3_syn_4 , \g237378/u3_syn_4 , \g237391/u3_syn_4 , \g237392/u3_syn_4 , \g237403/u3_syn_4 , \g237415/u3_syn_4 , \g237417/u3_syn_4 , \g237431/u3_syn_4 , \g237439/u3_syn_4 , \g237440/u3_syn_4 , \g237454/u3_syn_4 , \g237457/u3_syn_4 , \g237472/u3_syn_4 , \g237480/u3_syn_4 , \g237488/u3_syn_4 , \g237496/u3_syn_4 , \g237499/u3_syn_4 , \g237512/u3_syn_4 , \g237515/u3_syn_4 , \g237525/u3_syn_4 , \g237529/u3_syn_4 , \g237535/u3_syn_4 , \g237541/u3_syn_4 , \g237553/u3_syn_4 , \g237561/u3_syn_4 , \g237569/u3_syn_4 , \g237575/u3_syn_4 , \g237578/u3_syn_4 , \g237581/u3_syn_4 , \g237591/u3_syn_4 , \g237602/u3_syn_4 , \g237610/u3_syn_4 , \g237617/u3_syn_4 , \g237623/u3_syn_4 , \g237633/u3_syn_4 , \g237635/u3_syn_4 , \g237648/u3_syn_4 , \g237658/u3_syn_4 , \g237659/u3_syn_4 , \g237660/u3_syn_4 , \g237668/u3_syn_4 , \g237675/u3_syn_4 , \g237684/u3_syn_4 , \g237692/u3_syn_4 , \g237693/u3_syn_4 , \g237705/u3_syn_4 , \g237716/u3_syn_4 , \g237717/u3_syn_4 , \g237729/u3_syn_4 , \g237740/u3_syn_4 , \g237741/u3_syn_4 , \g237756/u3_syn_4 , \g237764/u3_syn_4 , \g237768/u3_syn_4 , \g237780/u3_syn_4 , \g237782/u3_syn_4 , \g237792/u3_syn_4 , \g237804/u3_syn_4 , \g237812/u3_syn_4 , \g237820/u3_syn_4 , \g237828/u3_syn_4 , \g237836/u3_syn_4 , \g237844/u3_syn_4 , \g237852/u3_syn_4 , \g237860/u3_syn_4 , \g237868/u3_syn_4 , \g237876/u3_syn_4 , \g237884/u3_syn_4 , \g237888/u3_syn_4 , \g237895/u3_syn_4 , \g237907/u3_syn_4 , \g237916/u3_syn_4 , \g237924/u3_syn_4 , \g237931/u3_syn_4 , \g237940/u3_syn_4 , \g237949/u3_syn_4 , \g237950/u3_syn_4 , \g237955/u3_syn_4 , \g237961/u3_syn_4 , \g237965/u3_syn_4 , \g237975/u3_syn_4 , \g237983/u3_syn_4 , \g237989/u3_syn_4 , \g237999/u3_syn_4 , \g238007/u3_syn_4 , \g238015/u3_syn_4 , \g238017/u3_syn_4 , \g238033/u3_syn_4 , \g238035/u3_syn_4 , \g238049/u3_syn_4 , \g238057/u3_syn_4 , \g238065/u3_syn_4 , \g238072/u3_syn_4 , \g238081/u3_syn_4 , \g238082/u3_syn_4 , \g238097/u3_syn_4 , \g238105/u3_syn_4 , \g238113/u3_syn_4 , \g238114/u3_syn_4 , \g238129/u3_syn_4 , \g238137/u3_syn_4 , \g238145/u3_syn_4 , \g238153/u3_syn_4 , \g238161/u3_syn_4 , \g238163/u3_syn_4 , \g238177/u3_syn_4 , \g238179/u3_syn_4 , \g238194/u3_syn_4 , \g238197/u3_syn_4 , \g238209/u3_syn_4 , \g238213/u3_syn_4 , \g238225/u3_syn_4 , \g238229/u3_syn_4 , \g238237/u3_syn_4 , \g238250/u3_syn_4 , \g238257/u3_syn_4 , \g238263/u3_syn_4 , \g238269/u3_syn_4 , \g238282/u3_syn_4 , \g238285/u3_syn_4 , \g238298/u3_syn_4 , \g238301/u3_syn_4 , \g238314/u3_syn_4 , \g238316/u3_syn_4 , \g238329/u3_syn_4 , \g238338/u3_syn_4 , \g238346/u3_syn_4 , \g238351/u3_syn_4 , \g238356/u3_syn_4 , \g238368/u3_syn_4 , \g238378/u3_syn_4 , \g238386/u3_syn_4 , \g238394/u3_syn_4 , \g238402/u3_syn_4 , \g238409/u3_syn_4 , \g238412/u3_syn_4 , \g238427/u3_syn_4 , \g238429/u3_syn_4 , \g238443/u3_syn_4 , \g238448/u3_syn_4 , \g238457/u3_syn_4 , \g238460/u3_syn_4 , \g238472/u3_syn_4 , \g238484/u3_syn_4 , \g238492/u3_syn_4 , \g238500/u3_syn_4 , \g238505/u3_syn_4 , \g238516/u3_syn_4 , \g238524/u3_syn_4 , \g238532/u3_syn_4 , \g238534/u3_syn_4 , \g238544/u3_syn_4 , \g238549/u3_syn_4 , \g238550/u3_syn_4 , \g238565/u3_syn_4 , \g238566/u3_syn_4 , \g238582/u3_syn_4 , \g238583/u3_syn_4 , \g238594/u3_syn_4 , \g238606/u3_syn_4 , \g238614/u3_syn_4 , \g238615/u3_syn_4 , \g238619/u3_syn_4 , \g238631/u3_syn_4 , \g238639/u3_syn_4 , \g238647/u3_syn_4 , \g238649/u3_syn_4 , \g238659/u3_syn_4 , \g238670/u3_syn_4 , \g238671/u3_syn_4 , \g238680/u3_syn_4 , \g238688/u3_syn_4 , \g238691/u3_syn_4 , \g238696/u3_syn_4 , \g238705/u3_syn_4 , \g238708/u3_syn_4 , \g238721/u3_syn_4 , \g238724/u3_syn_4 , \g238736/u3_syn_4 , \g238745/u3_syn_4 , \g238753/u3_syn_4 , \g238757/u3_syn_4 , \g238764/u3_syn_4 , \g238776/u3_syn_4 , \g238781/u3_syn_4 , \g238787/u3_syn_4 , \g238799/u3_syn_4 , \g238807/u3_syn_4 , \g238811/u3_syn_4 , \g238824/u3_syn_4 , \g238830/u3_syn_4 , \g238841/u3_syn_4 , \g238843/u3_syn_4 , \g238855/u3_syn_4 , \g238859/u3_syn_4 , \g238863/u3_syn_4 , \g238868/u3_syn_4 , \g238880/u3_syn_4 , \g238888/u3_syn_4 , \g238892/u3_syn_4 , \g238903/u3_syn_4 , \g238911/u3_syn_4 , \g238915/u3_syn_4 , \g238927/u3_syn_4 , \g238937/u3_syn_4 , \g238945/u3_syn_4 , \g238953/u3_syn_4 , \g238961/u3_syn_4 , \g238970/u3_syn_4 , \g238971/u3_syn_4 , \g238983/u3_syn_4 , \g238994/u3_syn_4 , \g239002/u3_syn_4 , \g239009/u3_syn_4 , \g239015/u3_syn_4 , \g239025/u3_syn_4 , \g239030/u3_syn_4 , \g239041/u3_syn_4 , \g239048/u3_syn_4 , \g239053/u3_syn_4 , \g239065/u3_syn_4 , \g239073/u3_syn_4 , \g239081/u3_syn_4 , \g239082/u3_syn_4 , \g239093/u3_syn_4 , \g239105/u3_syn_4 , \g239108/u3_syn_4 , \g239117/u3_syn_4 , \g239129/u3_syn_4 , \g239137/u3_syn_4 , \g239139/u3_syn_4 , \g239148/u3_syn_4 , \g239160/u3_syn_4 , \g239162/u3_syn_4 , \g239172/u3_syn_4 , \g239184/u3_syn_4 , \g239187/u3_syn_4 , \g239189/u3_syn_4 , \g239201/u3_syn_4 , \g239208/u3_syn_4 , \g239217/u3_syn_4 , \g239219/u3_syn_4 , \g239226/u3_syn_4 , \g239234/u3_syn_4 , \g239242/u3_syn_4 , \g239246/u3_syn_4 , \g239257/u3_syn_4 , \g239258/u3_syn_4 , \g239263/u3_syn_4 , \g239275/u3_syn_4 , \g239277/u3_syn_4 , \g239291/u3_syn_4 , \g239296/u3_syn_4 , \g239308/u3_syn_4 , \g239311/u3_syn_4 , \g239322/u3_syn_4 , \g239329/u3_syn_4 , \g239338/u3_syn_4 , \g239339/u3_syn_4 , \g239346/u3_syn_4 , \g239351/u3_syn_4 , \g239363/u3_syn_4 , \g239370/u3_syn_4 , \g239375/u3_syn_4 , \g239387/u3_syn_4 , \g239395/u3_syn_4 , \g239418/u3_syn_4 , \g239439/u3_syn_4 , \g239442/u3_syn_4 , \g239454/u3_syn_4 , \g239464/u3_syn_4 , \g239470/u3_syn_4 , \g239481/u3_syn_4 , \g239487/u3_syn_4 , \g239497/u3_syn_4 , \g239520/u3_syn_4 , \g239532/u3_syn_4 , \g239543/u3_syn_4 , \g239551/u3_syn_4 , \g239552/u3_syn_4 , \g239567/u3_syn_4 , \g239575/u3_syn_4 , \g239579/u3_syn_4 , \g239592/u3_syn_4 , \g239594/u3_syn_4 , \g239608/u3_syn_4 , \g239626/u3_syn_4 , \g239634/u3_syn_4 , \g239646/u3_syn_4 , \g239649/u3_syn_4 , \g239657/u3_syn_4 , \g239670/u3_syn_4 , \g239673/u3_syn_4 , \g239686/u3_syn_4 , \g239694/u3_syn_4 , \g239695/u3_syn_4 , \g239701/u3_syn_4 , \g239705/u3_syn_4 , \g239709/u3_syn_4 , \g239715/u3_syn_4 , \g239717/u3_syn_4 , \g239726/u3_syn_4 , \g239734/u3_syn_4 , \g239735/u3_syn_4 , \g239743/u3_syn_4 , \g239760/u3_syn_4 , \g239768/u3_syn_4 , \g239776/u3_syn_4 , \g239784/u3_syn_4 , \g239793/u3_syn_4 , \g239801/u3_syn_4 , \g239817/u3_syn_4 , \g239818/u3_syn_4 , \g239848/u3_syn_4 , \g239856/u3_syn_4 , \g239872/u3_syn_4 , \g239880/u3_syn_4 , \g239888/u3_syn_4 , \g239896/u3_syn_4 , \g239904/u3_syn_4 , \g239912/u3_syn_4 , \g239920/u3_syn_4 , \g239928/u3_syn_4 , \g239936/u3_syn_4 , \g239951/u3_syn_4 , \g239963/u3_syn_4 , \g239979/u3_syn_4 , \g239986/u3_syn_4 , \g239999/u3_syn_4 , \g240000/u3_syn_4 , \g240008/u3_syn_4 , \g240012/u3_syn_4 , \g240018/u3_syn_4 , \g240026/u3_syn_4 , \g240034/u3_syn_4 , \g240042/u3_syn_4 , \g240050/u3_syn_4 , \g240074/u3_syn_4 , \g240091/u3_syn_4 , \g240122/u3_syn_4 , \g240147/u3_syn_4 , \g240209/u3_syn_4 , \g240219/u3_syn_4 , \g240259/u3_syn_4 , \g240334/u3_syn_4 , \g240406/u3_syn_4 , \g240416/u3_syn_4 , \g240424/u3_syn_4 , \g240432/u3_syn_4 , \g240440/u3_syn_4 , \g240448/u3_syn_4 , \g240456/u3_syn_4 , \g240464/u3_syn_4 , \g240472/u3_syn_4 , \g240480/u3_syn_4 , \g240488/u3_syn_4 , \g240496/u3_syn_4 , \g240504/u3_syn_4 , \g240512/u3_syn_4 , \g240520/u3_syn_4 , \g240530/u3_syn_4 , \g240538/u3_syn_4 , \g240547/u3_syn_4 , \g240555/u3_syn_4 , \g240563/u3_syn_4 , \g240571/u3_syn_4 , \g240579/u3_syn_4 , \g240587/u3_syn_4 , \g240595/u3_syn_4 , \g240603/u3_syn_4 , \g240611/u3_syn_4 , \g240619/u3_syn_4 , \g240627/u3_syn_4 , \g240635/u3_syn_4 , \g240643/u3_syn_4 , \g240651/u3_syn_4 , \g240659/u3_syn_4 , \g240667/u3_syn_4 , \g240675/u3_syn_4 , \g240683/u3_syn_4 , \g240691/u3_syn_4 , \g240699/u3_syn_4 , \g240707/u3_syn_4 , \g240715/u3_syn_4 , \g240723/u3_syn_4 , \g240731/u3_syn_4 , \g240739/u3_syn_4 , \g240747/u3_syn_4 , \g240755/u3_syn_4 , \g240763/u3_syn_4 , \g240771/u3_syn_4 , \g240779/u3_syn_4 , \g240787/u3_syn_4 , \g240795/u3_syn_4 , \g240803/u3_syn_4 , \g240811/u3_syn_4 , \g240819/u3_syn_4 , \g240827/u3_syn_4 , \g240835/u3_syn_4 , \g240843/u3_syn_4 , \g240851/u3_syn_4 , \g240859/u3_syn_4 , \g240867/u3_syn_4 , \g240875/u3_syn_4 , \g240883/u3_syn_4 , \g240891/u3_syn_4 , \g240899/u3_syn_4 , \g240907/u3_syn_4 , \g240915/u3_syn_4 , \g240923/u3_syn_4 , \g240931/u3_syn_4 , \g240939/u3_syn_4 , \g240947/u3_syn_4 , \g240955/u3_syn_4 , \g240963/u3_syn_4 , \g240971/u3_syn_4 , \g240979/u3_syn_4 , \g240987/u3_syn_4 , \g240995/u3_syn_4 , \g241003/u3_syn_4 , \g241011/u3_syn_4 , \g241019/u3_syn_4 , \g241027/u3_syn_4 , \g241036/u3_syn_4 , \g241044/u3_syn_4 , \g241052/u3_syn_4 , \g241060/u3_syn_4 , \g241068/u3_syn_4 , \g241076/u3_syn_4 , \g241084/u3_syn_4 , \g241092/u3_syn_4 , \g241100/u3_syn_4 , \g241108/u3_syn_4 , \g241116/u3_syn_4 , \g241124/u3_syn_4 , \g241132/u3_syn_4 , \g241140/u3_syn_4 , \g241148/u3_syn_4 , \g241156/u3_syn_4 , \g241164/u3_syn_4 , \g241172/u3_syn_4 , \g241180/u3_syn_4 , \g241188/u3_syn_4 , \g241196/u3_syn_4 , \g241205/u3_syn_4 , \g241213/u3_syn_4 , \g241221/u3_syn_4 , \g241229/u3_syn_4 , \g241237/u3_syn_4 , \g241245/u3_syn_4 , \g241253/u3_syn_4 , \g241261/u3_syn_4 , \g241269/u3_syn_4 , \g241277/u3_syn_4 , \g241285/u3_syn_4 , \g241293/u3_syn_4 , \g241301/u3_syn_4 , \g241309/u3_syn_4 , \g241317/u3_syn_4 , \g241325/u3_syn_4 , \g241333/u3_syn_4 , \g241341/u3_syn_4 , \g241349/u3_syn_4 , \g241358/u3_syn_4 , \g241366/u3_syn_4 , \g241374/u3_syn_4 , \g241382/u3_syn_4 , \g241390/u3_syn_4 , \g241398/u3_syn_4 , \g241406/u3_syn_4 , \g241415/u3_syn_4 , \g241424/u3_syn_4 , \g241433/u3_syn_4 , \g241441/u3_syn_4 , \g241449/u3_syn_4 , \g241459/u3_syn_4 , \g241470/u3_syn_4 , \g241480/u3_syn_4 , \g241489/u3_syn_4 , \g241497/u3_syn_4 , \g241505/u3_syn_4 , \g241513/u3_syn_4 , \g241545/_3_ , \g241580/_00_ , \g241737/_0_ , \g241752/_0_ , \g241755/_0_ , \g241767/_2__syn_2 , \g241781/_1__syn_2 , \g241782/_0_ , \g241803/_1__syn_2 , \g241805/_0_ , \g241812/_1__syn_2 , \g241814/_1__syn_2 , \g241816/_1__syn_2 , \g241819/_1__syn_2 , \g241822/_1__syn_2 , \g241823/_0_ , \g241833/_1__syn_2 , \g241843/_1__syn_2 , \g241844/_1__syn_2 , \g241848/_1__syn_2 , \g241855/_1__syn_2 , \g241868/_1__syn_2 , \g242013/_1__syn_2 , \g242015/_1__syn_2 , \g242017/_1__syn_2 , \g242021/_1__syn_2 , \g242039/_1__syn_2 , \g242081/_0_ , \g242086/_0_ , \g242101/_3_ , \g242116/_0_ , \g242135/_2_ , \g242147/_0_ , \g242158/_0_ , \g242196/_0_ , \g242202/_0_ , \g242203/_0_ , \g242204/_0_ , \g242212/_0_ , \g242226/_01_ , \g242281/_0_ , \g242407/_0_ , \g242410/_0_ , \g242426/_0_ , \g242438/_2_ , \g242466/_0_ , \g242530/_0_ , \g242532/_0_ , \g243397/_0_ , \g245925/_0_ , \g245932/_0_ , \g245933/_0_ , \g245986/_3_ , \g250157/_3_ , \g250202/_0_ , \g250246/_1_ , \g250248/_0_ , \g250250/_0_ , \g250305/_0_ , \g250323/_0_ , \g250373/_0_ , \g250377/_0_ , \g250412/_0_ , \g250413/_0_ , \g250418/_0_ , \g250419/_0_ , \g250421/_0_ , \g250433/_0_ , \g250448/_3_ , \g250567/_3_ , \g258965/_0_ , \g259006/_0_ , \g259471/_0_ , \g259473/_2_ , \g260557/_0_ , \g261035/_0_ , \g261095/_3_ , \g261207/_2__syn_2 , \g261754/_0_ , \g262017/_0_ , \g262045/_0_ , \g262046/_0_ , \g262100/_3_ , \g263539/_1_ , \g263574/_0_ , \g263858/_0_ , \g264104/_1_ , \g264107/_1_ , \g264117/_0_ , \g264282/_0_ , \g264511/_0_ , \g264541/_0_ , \g264562/_0_ , \g264618/_0_ , \g264660/_0_ , \g264681/_3_ , \g264727/_0_ , \g265013/_0_ , \g265084/_0_ , \g265378/_0_ , \g265413/_0_ , \g265446/_0_ , \g265486/_0_ , \g265524/_3_ , \g265528/_3_ , \g265548/_3_ , \g265579/_0_ , \g265768/_0_ , \g265801/_0_ , \g265819/_1_ , \g265853/_0_ , \g265933/_0_ , \g266022/_0_ , \g266183/_1_ , \g281909/_0_ , \g281965/_1_ , \g282284/_1_ , \g282639/_1_ , \g283047/_0_ , \g283157/_1_ , \g283184/_0_ , \g283334/_3_ , int_o_pad, \m_wb_adr_o[0]_pad , \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2 , \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3 , \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3 );
	input \CarrierSense_Tx2_reg/NET0131  ;
	input \Collision_Tx1_reg/NET0131  ;
	input \Collision_Tx2_reg/NET0131  ;
	input \RstTxPauseRq_reg/NET0131  ;
	input \RxAbortRst_reg/NET0131  ;
	input \RxAbort_latch_reg/NET0131  ;
	input \RxAbort_wb_reg/NET0131  ;
	input \RxEnSync_reg/NET0131  ;
	input \TPauseRq_reg/NET0131  ;
	input \TxPauseRq_sync2_reg/NET0131  ;
	input \TxPauseRq_sync3_reg/NET0131  ;
	input \WillSendControlFrame_sync2_reg/NET0131  ;
	input \WillSendControlFrame_sync3_reg/NET0131  ;
	input \WillTransmit_q2_reg/P0001  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGR1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGR2_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_IPGT_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131  ;
	input \ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MODER_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_MODER_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_MODER_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131  ;
	input \ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131  ;
	input \ethreg1_ResetRxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_ResetRxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_ResetTxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_rxclk_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetRxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_sync2_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_sync3_reg/NET0131  ;
	input \ethreg1_SetTxCIrq_txclk_reg/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131  ;
	input \ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131  ;
	input \ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131  ;
	input \ethreg1_irq_busy_reg/NET0131  ;
	input \ethreg1_irq_rxb_reg/NET0131  ;
	input \ethreg1_irq_rxc_reg/NET0131  ;
	input \ethreg1_irq_rxe_reg/NET0131  ;
	input \ethreg1_irq_txb_reg/NET0131  ;
	input \ethreg1_irq_txc_reg/NET0131  ;
	input \ethreg1_irq_txe_reg/NET0131  ;
	input m_wb_ack_i_pad ;
	input \m_wb_adr_o[10]_pad  ;
	input \m_wb_adr_o[11]_pad  ;
	input \m_wb_adr_o[12]_pad  ;
	input \m_wb_adr_o[13]_pad  ;
	input \m_wb_adr_o[14]_pad  ;
	input \m_wb_adr_o[15]_pad  ;
	input \m_wb_adr_o[16]_pad  ;
	input \m_wb_adr_o[17]_pad  ;
	input \m_wb_adr_o[18]_pad  ;
	input \m_wb_adr_o[19]_pad  ;
	input \m_wb_adr_o[20]_pad  ;
	input \m_wb_adr_o[21]_pad  ;
	input \m_wb_adr_o[22]_pad  ;
	input \m_wb_adr_o[23]_pad  ;
	input \m_wb_adr_o[24]_pad  ;
	input \m_wb_adr_o[25]_pad  ;
	input \m_wb_adr_o[26]_pad  ;
	input \m_wb_adr_o[27]_pad  ;
	input \m_wb_adr_o[28]_pad  ;
	input \m_wb_adr_o[29]_pad  ;
	input \m_wb_adr_o[2]_pad  ;
	input \m_wb_adr_o[30]_pad  ;
	input \m_wb_adr_o[31]_pad  ;
	input \m_wb_adr_o[3]_pad  ;
	input \m_wb_adr_o[4]_pad  ;
	input \m_wb_adr_o[5]_pad  ;
	input \m_wb_adr_o[6]_pad  ;
	input \m_wb_adr_o[7]_pad  ;
	input \m_wb_adr_o[8]_pad  ;
	input \m_wb_adr_o[9]_pad  ;
	input \m_wb_dat_i[10]_pad  ;
	input \m_wb_dat_i[11]_pad  ;
	input \m_wb_dat_i[12]_pad  ;
	input \m_wb_dat_i[13]_pad  ;
	input \m_wb_dat_i[14]_pad  ;
	input \m_wb_dat_i[15]_pad  ;
	input \m_wb_dat_i[16]_pad  ;
	input \m_wb_dat_i[17]_pad  ;
	input \m_wb_dat_i[18]_pad  ;
	input \m_wb_dat_i[19]_pad  ;
	input \m_wb_dat_i[1]_pad  ;
	input \m_wb_dat_i[20]_pad  ;
	input \m_wb_dat_i[22]_pad  ;
	input \m_wb_dat_i[23]_pad  ;
	input \m_wb_dat_i[24]_pad  ;
	input \m_wb_dat_i[25]_pad  ;
	input \m_wb_dat_i[26]_pad  ;
	input \m_wb_dat_i[27]_pad  ;
	input \m_wb_dat_i[28]_pad  ;
	input \m_wb_dat_i[29]_pad  ;
	input \m_wb_dat_i[2]_pad  ;
	input \m_wb_dat_i[30]_pad  ;
	input \m_wb_dat_i[31]_pad  ;
	input \m_wb_dat_i[3]_pad  ;
	input \m_wb_dat_i[4]_pad  ;
	input \m_wb_dat_i[5]_pad  ;
	input \m_wb_dat_i[6]_pad  ;
	input \m_wb_dat_i[7]_pad  ;
	input \m_wb_dat_i[8]_pad  ;
	input m_wb_err_i_pad ;
	input \m_wb_sel_o[0]_pad  ;
	input \m_wb_sel_o[1]_pad  ;
	input \m_wb_sel_o[2]_pad  ;
	input \m_wb_sel_o[3]_pad  ;
	input m_wb_stb_o_pad ;
	input m_wb_we_o_pad ;
	input \maccontrol1_MuxedAbort_reg/NET0131  ;
	input \maccontrol1_MuxedDone_reg/NET0131  ;
	input \maccontrol1_TxAbortInLatched_reg/NET0131  ;
	input \maccontrol1_TxDoneInLatched_reg/NET0131  ;
	input \maccontrol1_TxUsedDataOutDetected_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_AddressOK_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_Divider2_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131  ;
	input \maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131  ;
	input \maccontrol1_receivecontrol1_Pause_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131  ;
	input \maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131  ;
	input \maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131  ;
	input \maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001  ;
	input \maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131  ;
	input \maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131  ;
	input \maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001  ;
	input \maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131  ;
	input \maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131  ;
	input \macstatus1_CarrierSenseLost_reg/NET0131  ;
	input \macstatus1_DeferLatched_reg/NET0131  ;
	input \macstatus1_DribbleNibble_reg/NET0131  ;
	input \macstatus1_InvalidSymbol_reg/NET0131  ;
	input \macstatus1_LatchedCrcError_reg/NET0131  ;
	input \macstatus1_LatchedMRxErr_reg/NET0131  ;
	input \macstatus1_LateCollLatched_reg/P0002  ;
	input \macstatus1_LoadRxStatus_reg/NET0131  ;
	input \macstatus1_ReceiveEnd_reg/NET0131  ;
	input \macstatus1_ReceivedPacketTooBig_reg/NET0131  ;
	input \macstatus1_RetryCntLatched_reg[0]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[1]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[2]/P0002  ;
	input \macstatus1_RetryCntLatched_reg[3]/P0002  ;
	input \macstatus1_RetryLimit_reg/P0002  ;
	input \macstatus1_RxColWindow_reg/NET0131  ;
	input \macstatus1_RxLateCollision_reg/NET0131  ;
	input \macstatus1_ShortFrame_reg/NET0131  ;
	input mcoll_pad_i_pad ;
	input md_pad_i_pad ;
	input mdc_pad_o_pad ;
	input \miim1_BitCounter_reg[0]/NET0131  ;
	input \miim1_BitCounter_reg[1]/NET0131  ;
	input \miim1_BitCounter_reg[2]/NET0131  ;
	input \miim1_BitCounter_reg[3]/NET0131  ;
	input \miim1_BitCounter_reg[4]/NET0131  ;
	input \miim1_BitCounter_reg[5]/NET0131  ;
	input \miim1_BitCounter_reg[6]/NET0131  ;
	input \miim1_EndBusy_reg/NET0131  ;
	input \miim1_InProgress_q1_reg/NET0131  ;
	input \miim1_InProgress_q2_reg/NET0131  ;
	input \miim1_InProgress_q3_reg/NET0131  ;
	input \miim1_InProgress_reg/NET0131  ;
	input \miim1_LatchByte0_d_reg/NET0131  ;
	input \miim1_LatchByte1_d_reg/NET0131  ;
	input \miim1_LatchByte_reg[0]/NET0131  ;
	input \miim1_LatchByte_reg[1]/NET0131  ;
	input \miim1_Nvalid_reg/NET0131  ;
	input \miim1_RStatStart_q1_reg/NET0131  ;
	input \miim1_RStatStart_q2_reg/NET0131  ;
	input \miim1_RStatStart_reg/NET0131  ;
	input \miim1_RStat_q2_reg/NET0131  ;
	input \miim1_RStat_q3_reg/NET0131  ;
	input \miim1_ScanStat_q2_reg/NET0131  ;
	input \miim1_SyncStatMdcEn_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q1_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q2_reg/NET0131  ;
	input \miim1_WCtrlDataStart_q_reg/NET0131  ;
	input \miim1_WCtrlDataStart_reg/NET0131  ;
	input \miim1_WCtrlData_q2_reg/NET0131  ;
	input \miim1_WCtrlData_q3_reg/NET0131  ;
	input \miim1_WriteOp_reg/NET0131  ;
	input \miim1_clkgen_Counter_reg[0]/NET0131  ;
	input \miim1_clkgen_Counter_reg[1]/NET0131  ;
	input \miim1_clkgen_Counter_reg[2]/NET0131  ;
	input \miim1_clkgen_Counter_reg[3]/NET0131  ;
	input \miim1_clkgen_Counter_reg[4]/NET0131  ;
	input \miim1_clkgen_Counter_reg[5]/NET0131  ;
	input \miim1_clkgen_Counter_reg[6]/NET0131  ;
	input \miim1_outctrl_Mdo_2d_reg/NET0131  ;
	input \miim1_shftrg_LinkFail_reg/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[0]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[1]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[2]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[3]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[4]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[5]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[6]/NET0131  ;
	input \miim1_shftrg_ShiftReg_reg[7]/NET0131  ;
	input \mrxd_pad_i[0]_pad  ;
	input \mrxd_pad_i[1]_pad  ;
	input \mrxd_pad_i[2]_pad  ;
	input \mrxd_pad_i[3]_pad  ;
	input mrxdv_pad_i_pad ;
	input mrxerr_pad_i_pad ;
	input \mtxd_pad_o[0]_pad  ;
	input \mtxd_pad_o[1]_pad  ;
	input \mtxd_pad_o[2]_pad  ;
	input \mtxd_pad_o[3]_pad  ;
	input mtxen_pad_o_pad ;
	input mtxerr_pad_o_pad ;
	input \rxethmac1_Broadcast_reg/NET0131  ;
	input \rxethmac1_CrcHashGood_reg/P0001  ;
	input \rxethmac1_CrcHash_reg[0]/P0001  ;
	input \rxethmac1_CrcHash_reg[1]/P0001  ;
	input \rxethmac1_CrcHash_reg[2]/P0001  ;
	input \rxethmac1_CrcHash_reg[3]/P0001  ;
	input \rxethmac1_CrcHash_reg[4]/P0001  ;
	input \rxethmac1_CrcHash_reg[5]/P0001  ;
	input \rxethmac1_DelayData_reg/NET0131  ;
	input \rxethmac1_LatchedByte_reg[0]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[1]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[2]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[3]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[4]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[5]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[6]/NET0131  ;
	input \rxethmac1_LatchedByte_reg[7]/NET0131  ;
	input \rxethmac1_Multicast_reg/NET0131  ;
	input \rxethmac1_RxData_d_reg[0]/NET0131  ;
	input \rxethmac1_RxData_d_reg[1]/NET0131  ;
	input \rxethmac1_RxData_d_reg[2]/NET0131  ;
	input \rxethmac1_RxData_d_reg[3]/NET0131  ;
	input \rxethmac1_RxData_d_reg[4]/NET0131  ;
	input \rxethmac1_RxData_d_reg[5]/NET0131  ;
	input \rxethmac1_RxData_d_reg[6]/NET0131  ;
	input \rxethmac1_RxData_d_reg[7]/NET0131  ;
	input \rxethmac1_RxData_reg[0]/NET0131  ;
	input \rxethmac1_RxData_reg[1]/NET0131  ;
	input \rxethmac1_RxData_reg[2]/NET0131  ;
	input \rxethmac1_RxData_reg[3]/NET0131  ;
	input \rxethmac1_RxData_reg[4]/NET0131  ;
	input \rxethmac1_RxData_reg[5]/NET0131  ;
	input \rxethmac1_RxData_reg[6]/NET0131  ;
	input \rxethmac1_RxData_reg[7]/NET0131  ;
	input \rxethmac1_RxEndFrm_d_reg/NET0131  ;
	input \rxethmac1_RxEndFrm_reg/NET0131  ;
	input \rxethmac1_RxStartFrm_reg/NET0131  ;
	input \rxethmac1_RxValid_reg/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[0]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[10]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[11]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[12]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[13]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[14]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[15]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[16]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[17]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[18]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[19]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[1]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[20]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[21]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[22]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[23]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[24]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[25]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[26]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[27]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[28]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[29]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[2]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[30]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[31]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[3]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[4]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[5]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[6]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[7]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[8]/NET0131  ;
	input \rxethmac1_crcrx_Crc_reg[9]/NET0131  ;
	input \rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131  ;
	input \rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131  ;
	input \rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131  ;
	input \rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131  ;
	input \rxethmac1_rxstatem1_StateData0_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateData1_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateDrop_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateIdle_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StatePreamble_reg/NET0131  ;
	input \rxethmac1_rxstatem1_StateSFD_reg/NET0131  ;
	input \txethmac1_ColWindow_reg/NET0131  ;
	input \txethmac1_PacketFinished_q_reg/NET0131  ;
	input \txethmac1_RetryCnt_reg[0]/NET0131  ;
	input \txethmac1_RetryCnt_reg[1]/NET0131  ;
	input \txethmac1_RetryCnt_reg[2]/NET0131  ;
	input \txethmac1_RetryCnt_reg[3]/NET0131  ;
	input \txethmac1_StatusLatch_reg/NET0131  ;
	input \txethmac1_StopExcessiveDeferOccured_reg/NET0131  ;
	input \txethmac1_TxAbort_reg/NET0131  ;
	input \txethmac1_TxDone_reg/NET0131  ;
	input \txethmac1_TxRetry_reg/NET0131  ;
	input \txethmac1_TxUsedData_reg/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[0]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[1]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[2]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[3]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[4]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[5]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[6]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[7]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[8]/NET0131  ;
	input \txethmac1_random1_RandomLatched_reg[9]/NET0131  ;
	input \txethmac1_random1_x_reg[1]/NET0131  ;
	input \txethmac1_random1_x_reg[2]/NET0131  ;
	input \txethmac1_random1_x_reg[3]/NET0131  ;
	input \txethmac1_random1_x_reg[4]/NET0131  ;
	input \txethmac1_random1_x_reg[5]/NET0131  ;
	input \txethmac1_random1_x_reg[6]/NET0131  ;
	input \txethmac1_random1_x_reg[7]/NET0131  ;
	input \txethmac1_random1_x_reg[8]/NET0131  ;
	input \txethmac1_random1_x_reg[9]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[10]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[11]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[12]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[13]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[14]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[15]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[3]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[4]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[5]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[6]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[7]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[8]/NET0131  ;
	input \txethmac1_txcounters1_ByteCnt_reg[9]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[0]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[10]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[11]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[12]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[13]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[14]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[15]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[1]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[2]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[3]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[4]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[5]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[6]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[7]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[8]/NET0131  ;
	input \txethmac1_txcounters1_NibCnt_reg[9]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[0]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[10]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[11]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[12]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[13]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[14]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[15]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[16]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[17]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[18]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[19]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[1]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[20]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[21]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[22]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[23]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[24]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[25]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[26]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[27]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[28]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[29]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[2]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[30]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[31]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[3]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[4]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[5]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[6]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[7]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[8]/NET0131  ;
	input \txethmac1_txcrc_Crc_reg[9]/NET0131  ;
	input \txethmac1_txstatem1_Rule1_reg/NET0131  ;
	input \txethmac1_txstatem1_StateBackOff_reg/NET0131  ;
	input \txethmac1_txstatem1_StateData_reg[0]/NET0131  ;
	input \txethmac1_txstatem1_StateData_reg[1]/NET0131  ;
	input \txethmac1_txstatem1_StateDefer_reg/NET0131  ;
	input \txethmac1_txstatem1_StateFCS_reg/NET0131  ;
	input \txethmac1_txstatem1_StateIPG_reg/NET0131  ;
	input \txethmac1_txstatem1_StateIdle_reg/NET0131  ;
	input \txethmac1_txstatem1_StateJam_q_reg/NET0131  ;
	input \txethmac1_txstatem1_StateJam_reg/NET0131  ;
	input \txethmac1_txstatem1_StatePAD_reg/NET0131  ;
	input \txethmac1_txstatem1_StatePreamble_reg/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_adr_i[10]_pad  ;
	input \wb_adr_i[11]_pad  ;
	input \wb_adr_i[2]_pad  ;
	input \wb_adr_i[3]_pad  ;
	input \wb_adr_i[4]_pad  ;
	input \wb_adr_i[5]_pad  ;
	input \wb_adr_i[6]_pad  ;
	input \wb_adr_i[7]_pad  ;
	input \wb_adr_i[8]_pad  ;
	input \wb_adr_i[9]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_dat_i[0]_pad  ;
	input \wb_dat_i[10]_pad  ;
	input \wb_dat_i[11]_pad  ;
	input \wb_dat_i[12]_pad  ;
	input \wb_dat_i[13]_pad  ;
	input \wb_dat_i[14]_pad  ;
	input \wb_dat_i[15]_pad  ;
	input \wb_dat_i[16]_pad  ;
	input \wb_dat_i[17]_pad  ;
	input \wb_dat_i[18]_pad  ;
	input \wb_dat_i[19]_pad  ;
	input \wb_dat_i[1]_pad  ;
	input \wb_dat_i[20]_pad  ;
	input \wb_dat_i[21]_pad  ;
	input \wb_dat_i[22]_pad  ;
	input \wb_dat_i[23]_pad  ;
	input \wb_dat_i[24]_pad  ;
	input \wb_dat_i[25]_pad  ;
	input \wb_dat_i[26]_pad  ;
	input \wb_dat_i[27]_pad  ;
	input \wb_dat_i[28]_pad  ;
	input \wb_dat_i[29]_pad  ;
	input \wb_dat_i[2]_pad  ;
	input \wb_dat_i[30]_pad  ;
	input \wb_dat_i[31]_pad  ;
	input \wb_dat_i[3]_pad  ;
	input \wb_dat_i[4]_pad  ;
	input \wb_dat_i[5]_pad  ;
	input \wb_dat_i[6]_pad  ;
	input \wb_dat_i[7]_pad  ;
	input \wb_dat_i[8]_pad  ;
	input \wb_dat_i[9]_pad  ;
	input wb_err_o_pad ;
	input wb_rst_i_pad ;
	input \wb_sel_i[0]_pad  ;
	input \wb_sel_i[1]_pad  ;
	input \wb_sel_i[2]_pad  ;
	input \wb_sel_i[3]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	input \wishbone_BDRead_reg/NET0131  ;
	input \wishbone_BDWrite_reg[0]/NET0131  ;
	input \wishbone_BDWrite_reg[1]/NET0131  ;
	input \wishbone_BDWrite_reg[2]/NET0131  ;
	input \wishbone_BDWrite_reg[3]/NET0131  ;
	input \wishbone_BlockReadTxDataFromMemory_reg/NET0131  ;
	input \wishbone_BlockingIncrementTxPointer_reg/NET0131  ;
	input \wishbone_BlockingTxBDRead_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_sync2_reg/NET0131  ;
	input \wishbone_BlockingTxStatusWrite_sync3_reg/NET0131  ;
	input \wishbone_Busy_IRQ_rck_reg/NET0131  ;
	input \wishbone_Busy_IRQ_sync2_reg/P0001  ;
	input \wishbone_Busy_IRQ_sync3_reg/P0001  ;
	input \wishbone_Busy_IRQ_syncb2_reg/P0001  ;
	input \wishbone_Flop_reg/NET0131  ;
	input \wishbone_IncrTxPointer_reg/NET0131  ;
	input \wishbone_LastByteIn_reg/NET0131  ;
	input \wishbone_LastWord_reg/NET0131  ;
	input \wishbone_LatchValidBytes_q_reg/NET0131  ;
	input \wishbone_LatchValidBytes_reg/NET0131  ;
	input \wishbone_LatchedRxLength_reg[0]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[10]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[11]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[12]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[13]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[14]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[15]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[1]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[2]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[3]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[4]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[5]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[6]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[7]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[8]/NET0131  ;
	input \wishbone_LatchedRxLength_reg[9]/NET0131  ;
	input \wishbone_LatchedRxStartFrm_reg/NET0131  ;
	input \wishbone_LatchedTxLength_reg[0]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[10]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[11]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[12]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[13]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[14]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[15]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[1]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[2]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[3]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[4]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[5]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[6]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[7]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[8]/NET0131  ;
	input \wishbone_LatchedTxLength_reg[9]/NET0131  ;
	input \wishbone_MasterWbRX_reg/NET0131  ;
	input \wishbone_MasterWbTX_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_sync2_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_sync3_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131  ;
	input \wishbone_ReadTxDataFromFifo_tck_reg/NET0131  ;
	input \wishbone_ReadTxDataFromMemory_reg/NET0131  ;
	input \wishbone_RxAbortLatched_reg/NET0131  ;
	input \wishbone_RxAbortSync2_reg/NET0131  ;
	input \wishbone_RxAbortSync3_reg/NET0131  ;
	input \wishbone_RxAbortSync4_reg/NET0131  ;
	input \wishbone_RxAbortSyncb2_reg/NET0131  ;
	input \wishbone_RxBDAddress_reg[1]/NET0131  ;
	input \wishbone_RxBDAddress_reg[2]/NET0131  ;
	input \wishbone_RxBDAddress_reg[3]/NET0131  ;
	input \wishbone_RxBDAddress_reg[4]/NET0131  ;
	input \wishbone_RxBDAddress_reg[5]/NET0131  ;
	input \wishbone_RxBDAddress_reg[6]/NET0131  ;
	input \wishbone_RxBDAddress_reg[7]/NET0131  ;
	input \wishbone_RxBDRead_reg/NET0131  ;
	input \wishbone_RxBDReady_reg/NET0131  ;
	input \wishbone_RxB_IRQ_reg/NET0131  ;
	input \wishbone_RxByteCnt_reg[0]/NET0131  ;
	input \wishbone_RxByteCnt_reg[1]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[10]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[11]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[12]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[13]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[14]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[15]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[16]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[17]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[18]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[19]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[20]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[21]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[22]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[23]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[24]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[25]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[26]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[27]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[28]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[29]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[30]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[31]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[8]/NET0131  ;
	input \wishbone_RxDataLatched1_reg[9]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[0]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[10]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[11]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[12]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[13]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[14]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[15]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[16]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[17]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[18]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[19]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[1]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[20]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[21]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[22]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[23]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[24]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[25]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[26]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[27]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[28]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[29]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[2]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[30]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[31]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[3]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[4]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[5]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[6]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[7]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[8]/NET0131  ;
	input \wishbone_RxDataLatched2_reg[9]/NET0131  ;
	input \wishbone_RxE_IRQ_reg/NET0131  ;
	input \wishbone_RxEn_needed_reg/NET0131  ;
	input \wishbone_RxEn_q_reg/NET0131  ;
	input \wishbone_RxEn_reg/NET0131  ;
	input \wishbone_RxEnableWindow_reg/NET0131  ;
	input \wishbone_RxOverrun_reg/NET0131  ;
	input \wishbone_RxPointerLSB_rst_reg[0]/NET0131  ;
	input \wishbone_RxPointerLSB_rst_reg[1]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[10]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[11]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[12]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[13]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[14]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[15]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[16]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[17]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[18]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[19]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[20]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[21]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[22]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[23]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[24]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[25]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[26]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[27]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[28]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[29]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[2]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[30]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[31]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[3]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[4]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[5]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[6]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[7]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[8]/NET0131  ;
	input \wishbone_RxPointerMSB_reg[9]/NET0131  ;
	input \wishbone_RxPointerRead_reg/NET0131  ;
	input \wishbone_RxReady_reg/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[0]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[1]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[2]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[3]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[4]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[5]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[6]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[7]/NET0131  ;
	input \wishbone_RxStatusInLatched_reg[8]/NET0131  ;
	input \wishbone_RxStatusWriteLatched_reg/NET0131  ;
	input \wishbone_RxStatusWriteLatched_sync2_reg/NET0131  ;
	input \wishbone_RxStatusWriteLatched_syncb2_reg/NET0131  ;
	input \wishbone_RxStatus_reg[13]/NET0131  ;
	input \wishbone_RxStatus_reg[14]/NET0131  ;
	input \wishbone_RxValidBytes_reg[0]/NET0131  ;
	input \wishbone_RxValidBytes_reg[1]/NET0131  ;
	input \wishbone_ShiftEndedSync1_reg/NET0131  ;
	input \wishbone_ShiftEndedSync2_reg/NET0131  ;
	input \wishbone_ShiftEndedSync3_reg/NET0131  ;
	input \wishbone_ShiftEndedSync_c1_reg/NET0131  ;
	input \wishbone_ShiftEndedSync_c2_reg/NET0131  ;
	input \wishbone_ShiftEnded_rck_reg/NET0131  ;
	input \wishbone_ShiftEnded_reg/NET0131  ;
	input \wishbone_ShiftWillEnd_reg/NET0131  ;
	input \wishbone_StartOccured_reg/NET0131  ;
	input \wishbone_SyncRxStartFrm_q2_reg/NET0131  ;
	input \wishbone_SyncRxStartFrm_q_reg/NET0131  ;
	input \wishbone_TxAbortPacketBlocked_reg/NET0131  ;
	input \wishbone_TxAbortPacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxAbortPacket_reg/NET0131  ;
	input \wishbone_TxAbort_q_reg/NET0131  ;
	input \wishbone_TxAbort_wb_q_reg/NET0131  ;
	input \wishbone_TxAbort_wb_reg/NET0131  ;
	input \wishbone_TxBDAddress_reg[1]/NET0131  ;
	input \wishbone_TxBDAddress_reg[2]/NET0131  ;
	input \wishbone_TxBDAddress_reg[3]/NET0131  ;
	input \wishbone_TxBDAddress_reg[4]/NET0131  ;
	input \wishbone_TxBDAddress_reg[5]/NET0131  ;
	input \wishbone_TxBDAddress_reg[6]/NET0131  ;
	input \wishbone_TxBDAddress_reg[7]/NET0131  ;
	input \wishbone_TxBDRead_reg/NET0131  ;
	input \wishbone_TxBDReady_reg/NET0131  ;
	input \wishbone_TxB_IRQ_reg/NET0131  ;
	input \wishbone_TxByteCnt_reg[0]/NET0131  ;
	input \wishbone_TxByteCnt_reg[1]/NET0131  ;
	input \wishbone_TxDataLatched_reg[0]/NET0131  ;
	input \wishbone_TxDataLatched_reg[10]/NET0131  ;
	input \wishbone_TxDataLatched_reg[11]/NET0131  ;
	input \wishbone_TxDataLatched_reg[12]/NET0131  ;
	input \wishbone_TxDataLatched_reg[13]/NET0131  ;
	input \wishbone_TxDataLatched_reg[14]/NET0131  ;
	input \wishbone_TxDataLatched_reg[15]/NET0131  ;
	input \wishbone_TxDataLatched_reg[16]/NET0131  ;
	input \wishbone_TxDataLatched_reg[17]/NET0131  ;
	input \wishbone_TxDataLatched_reg[18]/NET0131  ;
	input \wishbone_TxDataLatched_reg[19]/NET0131  ;
	input \wishbone_TxDataLatched_reg[1]/NET0131  ;
	input \wishbone_TxDataLatched_reg[20]/NET0131  ;
	input \wishbone_TxDataLatched_reg[21]/NET0131  ;
	input \wishbone_TxDataLatched_reg[22]/NET0131  ;
	input \wishbone_TxDataLatched_reg[23]/NET0131  ;
	input \wishbone_TxDataLatched_reg[24]/NET0131  ;
	input \wishbone_TxDataLatched_reg[25]/NET0131  ;
	input \wishbone_TxDataLatched_reg[26]/NET0131  ;
	input \wishbone_TxDataLatched_reg[27]/NET0131  ;
	input \wishbone_TxDataLatched_reg[28]/NET0131  ;
	input \wishbone_TxDataLatched_reg[29]/NET0131  ;
	input \wishbone_TxDataLatched_reg[2]/NET0131  ;
	input \wishbone_TxDataLatched_reg[30]/NET0131  ;
	input \wishbone_TxDataLatched_reg[31]/NET0131  ;
	input \wishbone_TxDataLatched_reg[3]/NET0131  ;
	input \wishbone_TxDataLatched_reg[4]/NET0131  ;
	input \wishbone_TxDataLatched_reg[5]/NET0131  ;
	input \wishbone_TxDataLatched_reg[6]/NET0131  ;
	input \wishbone_TxDataLatched_reg[7]/NET0131  ;
	input \wishbone_TxDataLatched_reg[8]/NET0131  ;
	input \wishbone_TxDataLatched_reg[9]/NET0131  ;
	input \wishbone_TxData_reg[0]/NET0131  ;
	input \wishbone_TxData_reg[1]/NET0131  ;
	input \wishbone_TxData_reg[2]/NET0131  ;
	input \wishbone_TxData_reg[3]/NET0131  ;
	input \wishbone_TxData_reg[4]/NET0131  ;
	input \wishbone_TxData_reg[5]/NET0131  ;
	input \wishbone_TxData_reg[6]/NET0131  ;
	input \wishbone_TxData_reg[7]/NET0131  ;
	input \wishbone_TxDonePacketBlocked_reg/NET0131  ;
	input \wishbone_TxDonePacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxDonePacket_reg/NET0131  ;
	input \wishbone_TxDone_wb_q_reg/NET0131  ;
	input \wishbone_TxDone_wb_reg/NET0131  ;
	input \wishbone_TxE_IRQ_reg/NET0131  ;
	input \wishbone_TxEn_needed_reg/NET0131  ;
	input \wishbone_TxEn_q_reg/NET0131  ;
	input \wishbone_TxEn_reg/NET0131  ;
	input \wishbone_TxEndFrm_reg/NET0131  ;
	input \wishbone_TxEndFrm_wb_reg/NET0131  ;
	input \wishbone_TxLength_reg[0]/NET0131  ;
	input \wishbone_TxLength_reg[10]/NET0131  ;
	input \wishbone_TxLength_reg[11]/NET0131  ;
	input \wishbone_TxLength_reg[12]/NET0131  ;
	input \wishbone_TxLength_reg[13]/NET0131  ;
	input \wishbone_TxLength_reg[14]/NET0131  ;
	input \wishbone_TxLength_reg[15]/NET0131  ;
	input \wishbone_TxLength_reg[1]/NET0131  ;
	input \wishbone_TxLength_reg[2]/NET0131  ;
	input \wishbone_TxLength_reg[3]/NET0131  ;
	input \wishbone_TxLength_reg[4]/NET0131  ;
	input \wishbone_TxLength_reg[5]/NET0131  ;
	input \wishbone_TxLength_reg[6]/NET0131  ;
	input \wishbone_TxLength_reg[7]/NET0131  ;
	input \wishbone_TxLength_reg[8]/NET0131  ;
	input \wishbone_TxLength_reg[9]/NET0131  ;
	input \wishbone_TxPointerLSB_reg[0]/NET0131  ;
	input \wishbone_TxPointerLSB_reg[1]/NET0131  ;
	input \wishbone_TxPointerLSB_rst_reg[0]/NET0131  ;
	input \wishbone_TxPointerLSB_rst_reg[1]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[10]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[11]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[12]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[13]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[14]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[15]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[16]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[17]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[18]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[19]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[20]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[21]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[22]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[23]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[24]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[25]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[26]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[27]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[28]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[29]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[2]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[30]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[31]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[3]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[4]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[5]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[6]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[7]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[8]/NET0131  ;
	input \wishbone_TxPointerMSB_reg[9]/NET0131  ;
	input \wishbone_TxPointerRead_reg/NET0131  ;
	input \wishbone_TxRetryPacketBlocked_reg/NET0131  ;
	input \wishbone_TxRetryPacket_NotCleared_reg/NET0131  ;
	input \wishbone_TxRetryPacket_reg/NET0131  ;
	input \wishbone_TxRetry_q_reg/NET0131  ;
	input \wishbone_TxRetry_wb_q_reg/NET0131  ;
	input \wishbone_TxRetry_wb_reg/NET0131  ;
	input \wishbone_TxStartFrm_reg/NET0131  ;
	input \wishbone_TxStartFrm_sync2_reg/NET0131  ;
	input \wishbone_TxStartFrm_syncb2_reg/NET0131  ;
	input \wishbone_TxStartFrm_wb_reg/NET0131  ;
	input \wishbone_TxStatus_reg[11]/NET0131  ;
	input \wishbone_TxStatus_reg[12]/NET0131  ;
	input \wishbone_TxStatus_reg[13]/NET0131  ;
	input \wishbone_TxStatus_reg[14]/NET0131  ;
	input \wishbone_TxUnderRun_reg/NET0131  ;
	input \wishbone_TxUnderRun_sync1_reg/NET0131  ;
	input \wishbone_TxUnderRun_wb_reg/NET0131  ;
	input \wishbone_TxUsedData_q_reg/NET0131  ;
	input \wishbone_TxValidBytesLatched_reg[0]/NET0131  ;
	input \wishbone_TxValidBytesLatched_reg[1]/NET0131  ;
	input \wishbone_WB_ACK_O_reg/P0001  ;
	input \wishbone_WbEn_q_reg/NET0131  ;
	input \wishbone_WbEn_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifoSync2_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifoSync3_reg/NET0131  ;
	input \wishbone_WriteRxDataToFifo_reg/NET0131  ;
	input \wishbone_bd_ram_mem0_reg[0][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[0][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[100][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[101][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[102][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[103][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[104][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[105][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[106][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[107][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[108][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[109][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[10][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[110][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[111][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[112][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[113][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[114][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[115][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[116][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[117][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[118][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[119][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[11][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[120][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[121][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[122][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[123][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[124][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[125][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[126][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[127][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[128][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[129][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[12][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[130][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[131][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[132][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[133][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[134][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[135][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[136][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[137][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[138][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[139][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[13][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[140][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[141][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[142][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[143][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[144][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[145][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[146][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[147][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[148][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[149][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[14][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[150][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[151][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[152][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[153][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[154][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[155][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[156][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[157][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[158][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[159][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[15][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[160][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[161][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[162][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[163][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[164][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[165][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[166][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[167][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[168][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[169][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[16][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[170][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[171][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[172][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[173][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[174][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[175][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[176][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[177][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[178][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[179][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[17][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[180][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[181][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[182][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[183][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[184][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[185][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[186][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[187][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[188][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[189][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[18][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[190][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[191][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[192][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[193][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[194][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[195][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[196][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[197][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[198][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[199][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[19][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[1][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[200][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[201][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[202][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[203][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[204][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[205][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[206][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[207][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[208][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[209][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[20][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[210][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[211][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[212][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[213][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[214][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[215][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[216][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[217][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[218][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[219][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[21][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[220][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[221][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[222][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[223][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[224][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[225][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[226][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[227][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[228][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[229][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[22][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[230][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[231][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[232][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[233][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[234][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[235][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[236][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[237][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[238][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[239][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[23][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[240][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[241][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[242][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[243][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[244][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[245][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[246][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[247][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[248][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[249][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[24][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[250][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[251][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[252][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[253][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[254][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[255][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[25][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[26][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[27][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[28][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[29][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[2][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[30][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[31][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[32][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[33][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[34][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[35][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[36][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[37][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[38][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[39][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[3][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[40][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[41][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[42][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[43][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[44][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[45][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[46][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[47][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[48][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[49][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[4][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[50][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[51][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[52][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[53][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[54][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[55][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[56][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[57][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[58][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[59][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[5][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[60][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[61][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[62][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[63][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[64][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[65][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[66][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[67][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[68][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[69][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[6][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[70][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[71][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[72][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[73][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[74][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[75][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[76][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[77][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[78][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[79][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[7][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[80][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[81][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[82][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[83][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[84][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[85][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[86][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[87][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[88][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[89][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[8][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[90][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[91][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[92][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[93][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[94][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[95][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[96][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[97][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[98][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[99][7]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][0]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][1]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][2]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][3]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][4]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][5]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][6]/P0001  ;
	input \wishbone_bd_ram_mem0_reg[9][7]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[0][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[100][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[101][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[102][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[103][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[104][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[105][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[106][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[107][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[108][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[109][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[10][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[110][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[111][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[112][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[113][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[114][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[115][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[116][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[117][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[118][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[119][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[11][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[120][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[121][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[122][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[123][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[124][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[125][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[126][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[127][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[128][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[129][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[12][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[130][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[131][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[132][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[133][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[134][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[135][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[136][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[137][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[138][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[139][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[13][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[140][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[141][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[142][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[143][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[144][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[145][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[146][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[147][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[148][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[149][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[14][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[150][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[151][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[152][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[153][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[154][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[155][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[156][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[157][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[158][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[159][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[15][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[160][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[161][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[162][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[163][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[164][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[165][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[166][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[167][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[168][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[169][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[16][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[170][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[171][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[172][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[173][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[174][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[175][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[176][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[177][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[178][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[179][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[17][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[180][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[181][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[182][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[183][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[184][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[185][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[186][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[187][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[188][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[189][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[18][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[190][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[191][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[192][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[193][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[194][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[195][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[196][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[197][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[198][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[199][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[19][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[1][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[200][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[201][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[202][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[203][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[204][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[205][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[206][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[207][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[208][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[209][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[20][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[210][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[211][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[212][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[213][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[214][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[215][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[216][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[217][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[218][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[219][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[21][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[220][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[221][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[222][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[223][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[224][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[225][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[226][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[227][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[228][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[229][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[22][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[230][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[231][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[232][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[233][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[234][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[235][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[236][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[237][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[238][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[239][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[23][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[240][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[241][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[242][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[243][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[244][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[245][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[246][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[247][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[248][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[249][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[24][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[250][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[251][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[252][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[253][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[254][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[255][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[25][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[26][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[27][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[28][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[29][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[2][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[30][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[31][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[32][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[33][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[34][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[35][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[36][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[37][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[38][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[39][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[3][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[40][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[41][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[42][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[43][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[44][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[45][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[46][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[47][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[48][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[49][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[4][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[50][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[51][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[52][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[53][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[54][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[55][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[56][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[57][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[58][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[59][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[5][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[60][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[61][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[62][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[63][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[64][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[65][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[66][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[67][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[68][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[69][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[6][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[70][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[71][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[72][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[73][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[74][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[75][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[76][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[77][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[78][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[79][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[7][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[80][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[81][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[82][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[83][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[84][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[85][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[86][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[87][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[88][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[89][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[8][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[90][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[91][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[92][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[93][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[94][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[95][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[96][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[97][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[98][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[99][9]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][10]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][11]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][12]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][13]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][14]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][15]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][8]/P0001  ;
	input \wishbone_bd_ram_mem1_reg[9][9]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[0][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[100][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[101][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[102][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[103][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[104][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[105][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[106][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[107][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[108][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[109][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[10][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[110][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[111][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[112][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[113][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[114][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[115][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[116][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[117][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[118][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[119][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[11][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[120][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[121][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[122][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[123][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[124][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[125][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[126][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[127][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[128][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[129][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[12][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[130][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[131][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[132][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[133][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[134][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[135][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[136][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[137][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[138][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[139][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[13][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[140][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[141][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[142][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[143][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[144][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[145][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[146][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[147][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[148][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[149][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[14][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[150][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[151][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[152][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[153][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[154][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[155][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[156][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[157][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[158][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[159][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[15][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[160][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[161][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[162][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[163][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[164][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[165][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[166][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[167][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[168][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[169][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[16][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[170][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[171][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[172][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[173][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[174][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[175][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[176][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[177][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[178][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[179][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[17][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[180][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[181][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[182][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[183][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[184][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[185][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[186][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[187][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[188][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[189][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[18][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[190][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[191][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[192][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[193][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[194][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[195][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[196][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[197][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[198][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[199][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[19][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[1][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[200][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[201][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[202][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[203][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[204][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[205][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[206][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[207][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[208][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[209][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[20][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[210][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[211][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[212][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[213][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[214][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[215][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[216][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[217][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[218][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[219][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[21][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[220][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[221][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[222][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[223][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[224][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[225][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[226][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[227][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[228][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[229][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[22][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[230][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[231][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[232][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[233][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[234][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[235][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[236][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[237][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[238][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[239][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[23][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[240][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[241][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[242][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[243][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[244][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[245][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[246][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[247][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[248][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[249][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[24][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[250][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[251][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[252][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[253][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[254][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[255][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[25][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[26][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[27][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[28][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[29][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[2][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[30][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[31][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[32][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[33][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[34][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[35][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[36][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[37][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[38][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[39][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[3][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[40][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[41][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[42][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[43][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[44][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[45][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[46][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[47][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[48][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[49][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[4][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[50][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[51][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[52][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[53][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[54][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[55][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[56][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[57][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[58][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[59][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[5][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[60][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[61][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[62][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[63][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[64][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[65][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[66][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[67][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[68][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[69][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[6][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[70][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[71][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[72][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[73][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[74][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[75][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[76][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[77][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[78][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[79][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[7][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[80][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[81][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[82][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[83][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[84][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[85][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[86][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[87][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[88][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[89][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[8][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[90][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[91][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[92][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[93][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[94][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[95][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[96][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[97][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[98][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[99][23]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][16]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][17]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][18]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][19]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][20]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][21]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][22]/P0001  ;
	input \wishbone_bd_ram_mem2_reg[9][23]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[0][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[100][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[101][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[102][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[103][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[104][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[105][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[106][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[107][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[108][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[109][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[10][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[110][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[111][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[112][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[113][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[114][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[115][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[116][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[117][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[118][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[119][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[11][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[120][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[121][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[122][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[123][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[124][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[125][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[126][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[127][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[128][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[129][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[12][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[130][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[131][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[132][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[133][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[134][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[135][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[136][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[137][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[138][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[139][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[13][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[140][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[141][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[142][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[143][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[144][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[145][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[146][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[147][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[148][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[149][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[14][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[150][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[151][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[152][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[153][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[154][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[155][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[156][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[157][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[158][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[159][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[15][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[160][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[161][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[162][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[163][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[164][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[165][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[166][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[167][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[168][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[169][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[16][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[170][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[171][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[172][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[173][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[174][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[175][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[176][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[177][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[178][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[179][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[17][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[180][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[181][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[182][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[183][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[184][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[185][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[186][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[187][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[188][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[189][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[18][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[190][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[191][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[192][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[193][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[194][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[195][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[196][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[197][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[198][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[199][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[19][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[1][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[200][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[201][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[202][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[203][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[204][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[205][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[206][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[207][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[208][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[209][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[20][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[210][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[211][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[212][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[213][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[214][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[215][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[216][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[217][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[218][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[219][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[21][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[220][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[221][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[222][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[223][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[224][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[225][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[226][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[227][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[228][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[229][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[22][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[230][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[231][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[232][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[233][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[234][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[235][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[236][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[237][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[238][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[239][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[23][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[240][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[241][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[242][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[243][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[244][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[245][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[246][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[247][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[248][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[249][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[24][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[250][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[251][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[252][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[253][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[254][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[255][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[25][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[26][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[27][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[28][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[29][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[2][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[30][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[31][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[32][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[33][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[34][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[35][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[36][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[37][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[38][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[39][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[3][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[40][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[41][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[42][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[43][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[44][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[45][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[46][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[47][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[48][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[49][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[4][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[50][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[51][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[52][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[53][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[54][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[55][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[56][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[57][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[58][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[59][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[5][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[60][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[61][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[62][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[63][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[64][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[65][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[66][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[67][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[68][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[69][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[6][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[70][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[71][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[72][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[73][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[74][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[75][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[76][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[77][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[78][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[79][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[7][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[80][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[81][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[82][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[83][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[84][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[85][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[86][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[87][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[88][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[89][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[8][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[90][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[91][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[92][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[93][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[94][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[95][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[96][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[97][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[98][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[99][31]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][24]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][25]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][26]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][27]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][28]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][29]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][30]/P0001  ;
	input \wishbone_bd_ram_mem3_reg[9][31]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[0]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[1]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[2]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[3]/P0001  ;
	input \wishbone_bd_ram_raddr_reg[4]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[5]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[6]/NET0131  ;
	input \wishbone_bd_ram_raddr_reg[7]/NET0131  ;
	input \wishbone_cyc_cleared_reg/NET0131  ;
	input \wishbone_r_RxEn_q_reg/NET0131  ;
	input \wishbone_r_TxEn_q_reg/NET0131  ;
	input \wishbone_ram_addr_reg[0]/NET0131  ;
	input \wishbone_ram_addr_reg[1]/NET0131  ;
	input \wishbone_ram_addr_reg[2]/NET0131  ;
	input \wishbone_ram_addr_reg[3]/NET0131  ;
	input \wishbone_ram_addr_reg[4]/NET0131  ;
	input \wishbone_ram_addr_reg[5]/NET0131  ;
	input \wishbone_ram_addr_reg[6]/NET0131  ;
	input \wishbone_ram_addr_reg[7]/NET0131  ;
	input \wishbone_ram_di_reg[0]/NET0131  ;
	input \wishbone_ram_di_reg[10]/NET0131  ;
	input \wishbone_ram_di_reg[11]/NET0131  ;
	input \wishbone_ram_di_reg[12]/NET0131  ;
	input \wishbone_ram_di_reg[13]/NET0131  ;
	input \wishbone_ram_di_reg[14]/NET0131  ;
	input \wishbone_ram_di_reg[15]/NET0131  ;
	input \wishbone_ram_di_reg[16]/NET0131  ;
	input \wishbone_ram_di_reg[17]/NET0131  ;
	input \wishbone_ram_di_reg[18]/NET0131  ;
	input \wishbone_ram_di_reg[19]/NET0131  ;
	input \wishbone_ram_di_reg[1]/NET0131  ;
	input \wishbone_ram_di_reg[20]/NET0131  ;
	input \wishbone_ram_di_reg[21]/NET0131  ;
	input \wishbone_ram_di_reg[22]/NET0131  ;
	input \wishbone_ram_di_reg[23]/NET0131  ;
	input \wishbone_ram_di_reg[24]/NET0131  ;
	input \wishbone_ram_di_reg[25]/NET0131  ;
	input \wishbone_ram_di_reg[26]/NET0131  ;
	input \wishbone_ram_di_reg[27]/NET0131  ;
	input \wishbone_ram_di_reg[28]/NET0131  ;
	input \wishbone_ram_di_reg[29]/NET0131  ;
	input \wishbone_ram_di_reg[2]/NET0131  ;
	input \wishbone_ram_di_reg[30]/NET0131  ;
	input \wishbone_ram_di_reg[31]/NET0131  ;
	input \wishbone_ram_di_reg[3]/NET0131  ;
	input \wishbone_ram_di_reg[4]/NET0131  ;
	input \wishbone_ram_di_reg[5]/NET0131  ;
	input \wishbone_ram_di_reg[6]/NET0131  ;
	input \wishbone_ram_di_reg[7]/NET0131  ;
	input \wishbone_ram_di_reg[8]/NET0131  ;
	input \wishbone_ram_di_reg[9]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[0]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[1]/NET0131  ;
	input \wishbone_rx_burst_cnt_reg[2]/NET0131  ;
	input \wishbone_rx_burst_en_reg/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[3]/NET0131  ;
	input \wishbone_rx_fifo_cnt_reg[4]/NET0131  ;
	input \wishbone_rx_fifo_fifo_reg[0][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[0][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[10][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[11][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[12][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[13][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[14][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[15][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[1][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[2][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[3][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[4][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[5][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[6][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[7][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[8][9]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][0]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][10]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][11]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][12]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][13]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][14]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][15]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][16]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][17]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][18]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][19]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][1]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][20]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][21]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][22]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][23]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][24]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][25]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][26]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][27]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][28]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][29]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][2]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][30]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][31]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][3]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][4]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][5]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][6]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][7]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][8]/P0001  ;
	input \wishbone_rx_fifo_fifo_reg[9][9]/P0001  ;
	input \wishbone_rx_fifo_read_pointer_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_read_pointer_reg[3]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[0]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[1]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[2]/NET0131  ;
	input \wishbone_rx_fifo_write_pointer_reg[3]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[0]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[1]/NET0131  ;
	input \wishbone_tx_burst_cnt_reg[2]/NET0131  ;
	input \wishbone_tx_burst_en_reg/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[3]/NET0131  ;
	input \wishbone_tx_fifo_cnt_reg[4]/NET0131  ;
	input \wishbone_tx_fifo_data_out_reg[0]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[10]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[11]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[12]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[13]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[14]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[15]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[16]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[17]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[18]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[19]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[1]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[20]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[21]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[22]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[23]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[24]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[25]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[26]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[27]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[28]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[29]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[2]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[30]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[31]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[3]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[4]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[5]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[6]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[7]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[8]/P0001  ;
	input \wishbone_tx_fifo_data_out_reg[9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[0][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[10][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[11][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[12][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[13][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[14][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[15][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[1][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[2][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[3][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[4][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[5][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[6][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[7][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[8][9]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][0]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][10]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][11]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][12]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][13]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][14]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][15]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][16]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][17]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][18]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][19]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][1]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][20]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][21]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][22]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][23]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][24]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][25]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][26]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][27]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][28]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][29]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][2]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][30]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][31]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][3]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][4]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][5]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][6]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][7]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][8]/P0001  ;
	input \wishbone_tx_fifo_fifo_reg[9][9]/P0001  ;
	input \wishbone_tx_fifo_read_pointer_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_read_pointer_reg[3]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[0]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[1]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[2]/NET0131  ;
	input \wishbone_tx_fifo_write_pointer_reg[3]/NET0131  ;
	output \_al_n1  ;
	output \g215539/_0_  ;
	output \g215543/_0_  ;
	output \g215547/_0_  ;
	output \g215551/_0_  ;
	output \g215552/_0_  ;
	output \g215578/_0_  ;
	output \g215587/_1_  ;
	output \g215589/_1_  ;
	output \g215591/_1_  ;
	output \g215593/_1_  ;
	output \g215595/_1_  ;
	output \g215597/_1_  ;
	output \g215599/_1_  ;
	output \g215601/_1_  ;
	output \g215603/_1_  ;
	output \g215605/_1_  ;
	output \g215607/_1_  ;
	output \g215609/_1_  ;
	output \g215611/_1_  ;
	output \g215613/_1_  ;
	output \g215615/_1_  ;
	output \g215617/_1_  ;
	output \g215618/_0_  ;
	output \g215619/_0_  ;
	output \g215620/_0_  ;
	output \g215632/_1_  ;
	output \g215634/_0_  ;
	output \g215635/_0_  ;
	output \g215636/_0_  ;
	output \g215637/_0_  ;
	output \g215638/_0_  ;
	output \g215639/_0_  ;
	output \g215655/_1_  ;
	output \g215657/_1_  ;
	output \g215659/_1_  ;
	output \g215661/_1_  ;
	output \g215662/_0_  ;
	output \g215663/_0_  ;
	output \g215664/_0_  ;
	output \g215665/_0_  ;
	output \g215668/_0_  ;
	output \g215674/_0_  ;
	output \g215677/_0_  ;
	output \g215686/_0_  ;
	output \g215695/_0_  ;
	output \g215696/_0_  ;
	output \g215702/_1__syn_2  ;
	output \g215705/_0_  ;
	output \g215706/_0_  ;
	output \g215716/_0_  ;
	output \g215717/_0_  ;
	output \g215718/_0_  ;
	output \g215726/_0_  ;
	output \g215727/_0_  ;
	output \g215728/_0_  ;
	output \g215760/_0_  ;
	output \g215764/_0_  ;
	output \g215765/_0_  ;
	output \g215766/_0_  ;
	output \g215767/_3_  ;
	output \g215768/_3_  ;
	output \g215769/_3_  ;
	output \g215770/_3_  ;
	output \g215771/_3_  ;
	output \g215772/_3_  ;
	output \g215773/_3_  ;
	output \g215774/_3_  ;
	output \g215775/_3_  ;
	output \g215776/_3_  ;
	output \g215777/_3_  ;
	output \g215778/_3_  ;
	output \g215779/_3_  ;
	output \g215780/_3_  ;
	output \g215790/_0_  ;
	output \g215791/_0_  ;
	output \g215792/_0_  ;
	output \g215793/_0_  ;
	output \g215801/_0_  ;
	output \g215802/_0_  ;
	output \g215803/_0_  ;
	output \g215804/_0_  ;
	output \g215812/_0_  ;
	output \g215813/_0_  ;
	output \g215821/_0_  ;
	output \g215823/_0_  ;
	output \g215831/_0_  ;
	output \g215832/_0_  ;
	output \g215833/_0_  ;
	output \g215845/_0_  ;
	output \g215846/_0_  ;
	output \g215847/_0_  ;
	output \g215872/_0_  ;
	output \g215873/_0_  ;
	output \g215874/_0_  ;
	output \g215904/_0_  ;
	output \g215905/_0_  ;
	output \g215906/_0_  ;
	output \g215907/_0_  ;
	output \g215908/_0_  ;
	output \g215909/_0_  ;
	output \g215910/_0_  ;
	output \g215911/_0_  ;
	output \g215912/_0_  ;
	output \g215913/_0_  ;
	output \g215914/_0_  ;
	output \g215915/_0_  ;
	output \g215916/_0_  ;
	output \g215917/_0_  ;
	output \g215918/_0_  ;
	output \g215919/_0_  ;
	output \g215920/_0_  ;
	output \g215923/_0_  ;
	output \g215926/_0_  ;
	output \g215941/_0_  ;
	output \g215942/_0_  ;
	output \g215943/_0_  ;
	output \g215944/_0_  ;
	output \g215945/_0_  ;
	output \g215946/_0_  ;
	output \g215947/_0_  ;
	output \g215948/_0_  ;
	output \g215949/_0_  ;
	output \g215950/_0_  ;
	output \g215951/_0_  ;
	output \g215952/_0_  ;
	output \g215953/_0_  ;
	output \g215954/_0_  ;
	output \g215955/_0_  ;
	output \g215956/_0_  ;
	output \g215957/_0_  ;
	output \g215959/_00_  ;
	output \g215960/_0_  ;
	output \g215962/_0_  ;
	output \g215964/_0_  ;
	output \g215966/_0_  ;
	output \g215972/_0_  ;
	output \g216035/_0_  ;
	output \g216037/_0_  ;
	output \g216038/_0_  ;
	output \g216039/_0_  ;
	output \g216040/_0_  ;
	output \g216041/_0_  ;
	output \g216042/_0_  ;
	output \g216046/_0_  ;
	output \g216048/_0_  ;
	output \g216057/_0_  ;
	output \g216263/_0_  ;
	output \g216264/_0_  ;
	output \g216265/_0_  ;
	output \g216266/_0_  ;
	output \g216267/_0_  ;
	output \g216268/_0_  ;
	output \g216269/_0_  ;
	output \g216270/_0_  ;
	output \g216271/_0_  ;
	output \g216272/_0_  ;
	output \g216273/_0_  ;
	output \g216284/_0_  ;
	output \g216289/_0_  ;
	output \g216290/_0_  ;
	output \g216292/_0_  ;
	output \g216296/_0_  ;
	output \g216297/_0_  ;
	output \g216300/_0_  ;
	output \g216301/_0_  ;
	output \g216302/_0_  ;
	output \g216303/_0_  ;
	output \g216304/_0_  ;
	output \g216305/_0_  ;
	output \g216306/_0_  ;
	output \g216307/_0_  ;
	output \g216310/_3_  ;
	output \g216311/_3_  ;
	output \g216314/u3_syn_7  ;
	output \g216322/_3_  ;
	output \g216323/_3_  ;
	output \g216324/_3_  ;
	output \g216325/_3_  ;
	output \g216326/_3_  ;
	output \g216327/_3_  ;
	output \g216328/_3_  ;
	output \g216329/_3_  ;
	output \g216369/_0_  ;
	output \g216370/_0_  ;
	output \g216371/_0_  ;
	output \g216372/_0_  ;
	output \g216373/_0_  ;
	output \g216374/_0_  ;
	output \g216375/_0_  ;
	output \g216376/_0_  ;
	output \g216379/_0_  ;
	output \g216380/_0_  ;
	output \g216381/_0_  ;
	output \g216385/_0_  ;
	output \g216389/_0_  ;
	output \g216390/_0_  ;
	output \g216402/_0_  ;
	output \g216404/_0_  ;
	output \g216405/_0_  ;
	output \g216406/_0_  ;
	output \g216407/_0_  ;
	output \g216408/_0_  ;
	output \g216409/_0_  ;
	output \g216410/_0_  ;
	output \g216411/_0_  ;
	output \g216412/_0_  ;
	output \g216413/_0_  ;
	output \g216414/_0_  ;
	output \g216415/_0_  ;
	output \g216416/_0_  ;
	output \g216417/_0_  ;
	output \g216418/_0_  ;
	output \g216419/_0_  ;
	output \g216420/_0_  ;
	output \g216421/_0_  ;
	output \g216422/_0_  ;
	output \g216423/_0_  ;
	output \g216424/_0_  ;
	output \g216425/_0_  ;
	output \g216426/_0_  ;
	output \g216427/_0_  ;
	output \g216428/_0_  ;
	output \g216429/_0_  ;
	output \g216430/_0_  ;
	output \g216431/_0_  ;
	output \g216432/_0_  ;
	output \g216433/_0_  ;
	output \g216434/_0_  ;
	output \g216435/_0_  ;
	output \g216436/_0_  ;
	output \g216437/_0_  ;
	output \g216438/_0_  ;
	output \g216439/_3_  ;
	output \g216447/_3_  ;
	output \g216448/_3_  ;
	output \g216452/_0_  ;
	output \g216453/_0_  ;
	output \g216454/_0_  ;
	output \g216455/_0_  ;
	output \g216456/_0_  ;
	output \g216457/_0_  ;
	output \g216458/_3_  ;
	output \g216459/_3_  ;
	output \g216461/_3_  ;
	output \g216462/_3_  ;
	output \g216463/_3_  ;
	output \g216464/_3_  ;
	output \g216465/_3_  ;
	output \g216466/_0_  ;
	output \g216467/_3_  ;
	output \g216468/_3_  ;
	output \g216469/_3_  ;
	output \g216470/_3_  ;
	output \g216471/_3_  ;
	output \g216473/_3_  ;
	output \g216474/_3_  ;
	output \g216475/_3_  ;
	output \g216476/_3_  ;
	output \g216477/_3_  ;
	output \g216478/_0_  ;
	output \g216479/_3_  ;
	output \g216480/_3_  ;
	output \g216481/_3_  ;
	output \g216492/_0_  ;
	output \g216494/_0_  ;
	output \g216495/_3_  ;
	output \g216496/_3_  ;
	output \g216498/_3_  ;
	output \g216499/_3_  ;
	output \g216500/_3_  ;
	output \g216513/_3_  ;
	output \g216514/_3_  ;
	output \g216515/_3_  ;
	output \g216516/_3_  ;
	output \g216517/_3_  ;
	output \g216518/_3_  ;
	output \g216519/_3_  ;
	output \g216520/_3_  ;
	output \g216521/_3_  ;
	output \g216522/_3_  ;
	output \g216523/_3_  ;
	output \g216524/_3_  ;
	output \g216525/_3_  ;
	output \g216526/_3_  ;
	output \g216527/_3_  ;
	output \g216528/_3_  ;
	output \g216529/_3_  ;
	output \g216530/_3_  ;
	output \g216531/_3_  ;
	output \g216532/_3_  ;
	output \g216533/_3_  ;
	output \g216534/_3_  ;
	output \g216535/_3_  ;
	output \g216536/_3_  ;
	output \g216537/_3_  ;
	output \g216538/_3_  ;
	output \g216555/_3_  ;
	output \g216556/_3_  ;
	output \g216557/_3_  ;
	output \g216560/_3_  ;
	output \g216561/_3_  ;
	output \g216562/_3_  ;
	output \g216563/_3_  ;
	output \g216564/_3_  ;
	output \g216565/_3_  ;
	output \g216566/_3_  ;
	output \g216567/_3_  ;
	output \g216568/_3_  ;
	output \g216569/_3_  ;
	output \g216570/_3_  ;
	output \g216571/_3_  ;
	output \g216575/_3_  ;
	output \g216576/_3_  ;
	output \g216577/_3_  ;
	output \g216578/_3_  ;
	output \g216579/_3_  ;
	output \g216580/_3_  ;
	output \g216581/_3_  ;
	output \g216582/_3_  ;
	output \g216583/_3_  ;
	output \g216586/_3_  ;
	output \g216587/_3_  ;
	output \g216588/_3_  ;
	output \g216589/_3_  ;
	output \g216590/_3_  ;
	output \g216591/_3_  ;
	output \g216592/_3_  ;
	output \g216593/_3_  ;
	output \g216594/_3_  ;
	output \g216595/_3_  ;
	output \g216600/_3_  ;
	output \g216683/_0_  ;
	output \g216689/_0_  ;
	output \g216693/_0_  ;
	output \g216694/_0_  ;
	output \g216727/_0_  ;
	output \g216728/_0_  ;
	output \g216729/_0_  ;
	output \g216732/_0_  ;
	output \g216733/_0_  ;
	output \g216734/_0_  ;
	output \g216735/_0_  ;
	output \g216736/_0_  ;
	output \g216737/_0_  ;
	output \g216738/_0_  ;
	output \g216739/_0_  ;
	output \g216740/_0_  ;
	output \g216741/_0_  ;
	output \g216742/_0_  ;
	output \g216743/_0_  ;
	output \g216744/_0_  ;
	output \g216745/_0_  ;
	output \g216746/_0_  ;
	output \g216748/_0_  ;
	output \g216751/_0_  ;
	output \g216754/_0_  ;
	output \g216762/_0_  ;
	output \g216934/_2_  ;
	output \g216952/_0_  ;
	output \g216955/_0_  ;
	output \g216969/_0_  ;
	output \g216979/_0_  ;
	output \g216984/_0_  ;
	output \g216996/_0_  ;
	output \g217002/_0_  ;
	output \g217014/_0_  ;
	output \g217015/_0_  ;
	output \g217016/_0_  ;
	output \g217017/_0_  ;
	output \g217018/_0_  ;
	output \g217019/_0_  ;
	output \g217023/_0_  ;
	output \g217116/_0_  ;
	output \g217146/_3_  ;
	output \g217149/_0_  ;
	output \g217151/_0_  ;
	output \g217160/_0_  ;
	output \g217167/_0_  ;
	output \g217168/_0_  ;
	output \g217169/_0_  ;
	output \g217170/_0_  ;
	output \g217171/_0_  ;
	output \g217172/_0_  ;
	output \g217173/_0_  ;
	output \g217174/_0_  ;
	output \g217175/_0_  ;
	output \g217176/_0_  ;
	output \g217177/_0_  ;
	output \g217178/_0_  ;
	output \g217179/_0_  ;
	output \g217180/_0_  ;
	output \g217181/_0_  ;
	output \g217182/_0_  ;
	output \g217183/_0_  ;
	output \g217187/_0_  ;
	output \g217188/_0_  ;
	output \g217189/_0_  ;
	output \g217193/_0_  ;
	output \g217194/_0_  ;
	output \g217195/_0_  ;
	output \g217196/_0_  ;
	output \g217202/_0_  ;
	output \g217205/_0_  ;
	output \g217206/_0_  ;
	output \g217207/_0_  ;
	output \g217208/_0_  ;
	output \g217209/_0_  ;
	output \g217210/_0_  ;
	output \g217211/_0_  ;
	output \g217212/_0_  ;
	output \g217213/_0_  ;
	output \g217214/_0_  ;
	output \g217215/_0_  ;
	output \g217216/_0_  ;
	output \g217217/_0_  ;
	output \g217218/_0_  ;
	output \g217219/_0_  ;
	output \g217220/_0_  ;
	output \g217223/_0_  ;
	output \g217231/_0_  ;
	output \g217237/_0_  ;
	output \g217238/_0_  ;
	output \g217242/_0_  ;
	output \g217243/_0_  ;
	output \g217250/_3_  ;
	output \g217251/_3_  ;
	output \g217252/_3_  ;
	output \g217253/_3_  ;
	output \g217254/_3_  ;
	output \g217255/_3_  ;
	output \g217256/_3_  ;
	output \g217257/_3_  ;
	output \g217258/_3_  ;
	output \g217259/_3_  ;
	output \g217260/_3_  ;
	output \g217261/_3_  ;
	output \g217262/_3_  ;
	output \g217263/_3_  ;
	output \g217264/_3_  ;
	output \g217265/_3_  ;
	output \g217266/_3_  ;
	output \g217267/_3_  ;
	output \g217268/_3_  ;
	output \g217269/_3_  ;
	output \g217270/_3_  ;
	output \g217271/_3_  ;
	output \g217272/_3_  ;
	output \g217273/_3_  ;
	output \g217274/_3_  ;
	output \g217275/_3_  ;
	output \g217276/_3_  ;
	output \g217277/_3_  ;
	output \g217278/_3_  ;
	output \g217279/_3_  ;
	output \g217280/_3_  ;
	output \g217281/_3_  ;
	output \g217282/_3_  ;
	output \g217283/_3_  ;
	output \g217284/_3_  ;
	output \g217285/_3_  ;
	output \g217286/_3_  ;
	output \g217287/_3_  ;
	output \g217288/_3_  ;
	output \g217289/_3_  ;
	output \g217290/_3_  ;
	output \g217291/_3_  ;
	output \g217292/_3_  ;
	output \g217293/_3_  ;
	output \g217294/_3_  ;
	output \g217295/_3_  ;
	output \g217296/_3_  ;
	output \g217297/_3_  ;
	output \g217298/_3_  ;
	output \g217299/_3_  ;
	output \g217300/_3_  ;
	output \g217301/_3_  ;
	output \g217302/_3_  ;
	output \g217303/_3_  ;
	output \g217304/_3_  ;
	output \g217305/_3_  ;
	output \g217306/_3_  ;
	output \g217307/_3_  ;
	output \g217308/_3_  ;
	output \g217309/_3_  ;
	output \g217310/_3_  ;
	output \g217311/_3_  ;
	output \g217312/_3_  ;
	output \g217313/_3_  ;
	output \g217318/_0_  ;
	output \g217662/_0_  ;
	output \g217663/_0_  ;
	output \g217682/_0_  ;
	output \g217697/_0_  ;
	output \g217698/_0_  ;
	output \g217699/_0_  ;
	output \g217700/_0_  ;
	output \g217701/_0_  ;
	output \g217705/_0_  ;
	output \g217711/_0_  ;
	output \g217747/_0_  ;
	output \g217753/_00_  ;
	output \g217775/_0_  ;
	output \g217781/_0_  ;
	output \g217784/_0_  ;
	output \g217785/_0_  ;
	output \g217786/_0_  ;
	output \g217787/_0_  ;
	output \g217788/_0_  ;
	output \g217790/_0_  ;
	output \g217815/_0_  ;
	output \g217817/_0_  ;
	output \g218145/_0_  ;
	output \g218148/_0_  ;
	output \g218150/_0_  ;
	output \g218167/_0_  ;
	output \g218168/_0_  ;
	output \g218234/_0_  ;
	output \g218235/_0_  ;
	output \g218236/_0_  ;
	output \g218238/_0_  ;
	output \g218242/_0_  ;
	output \g218332/_0_  ;
	output \g218335/_0_  ;
	output \g218336/_0_  ;
	output \g218337/_0_  ;
	output \g218338/_0_  ;
	output \g218339/_0_  ;
	output \g218340/_0_  ;
	output \g218341/_0_  ;
	output \g218342/_0_  ;
	output \g218343/_0_  ;
	output \g218344/_0_  ;
	output \g218345/_0_  ;
	output \g218346/_0_  ;
	output \g218347/_0_  ;
	output \g218348/_0_  ;
	output \g218349/_0_  ;
	output \g218350/_0_  ;
	output \g218351/_0_  ;
	output \g218352/_0_  ;
	output \g218353/_0_  ;
	output \g218354/_0_  ;
	output \g218355/_0_  ;
	output \g218356/_0_  ;
	output \g218357/_0_  ;
	output \g218358/_0_  ;
	output \g218359/_0_  ;
	output \g218360/_0_  ;
	output \g218398/_3_  ;
	output \g218430/_0_  ;
	output \g218440/_0_  ;
	output \g218452/u3_syn_4  ;
	output \g218495/u3_syn_4  ;
	output \g218517/u3_syn_4  ;
	output \g218554/u3_syn_4  ;
	output \g218575/u3_syn_4  ;
	output \g218600/u3_syn_4  ;
	output \g218621/u3_syn_4  ;
	output \g218638/u3_syn_4  ;
	output \g218659/u3_syn_4  ;
	output \g218673/u3_syn_4  ;
	output \g218707/u3_syn_4  ;
	output \g218735/_3_  ;
	output \g219186/_0_  ;
	output \g219187/_0_  ;
	output \g219188/_0_  ;
	output \g219189/_0_  ;
	output \g219190/_0_  ;
	output \g219196/_0_  ;
	output \g219198/_0_  ;
	output \g219199/_0_  ;
	output \g219200/_0_  ;
	output \g219308/_0_  ;
	output \g219314/_0_  ;
	output \g219326/_0_  ;
	output \g219328/_0_  ;
	output \g219348/_0_  ;
	output \g219351/_0_  ;
	output \g219363/_0_  ;
	output \g219364/_0_  ;
	output \g219365/_0_  ;
	output \g219366/_0_  ;
	output \g219367/_0_  ;
	output \g219368/_0_  ;
	output \g219369/_0_  ;
	output \g219376/_0_  ;
	output \g219381/_0_  ;
	output \g219382/_0_  ;
	output \g219384/_0_  ;
	output \g219385/_0_  ;
	output \g219391/_0_  ;
	output \g219394/_0_  ;
	output \g219395/_0_  ;
	output \g219396/_0_  ;
	output \g219397/_0_  ;
	output \g219398/_0_  ;
	output \g219399/_0_  ;
	output \g219400/_0_  ;
	output \g219401/_0_  ;
	output \g219402/_0_  ;
	output \g219403/_0_  ;
	output \g219404/_0_  ;
	output \g219405/_0_  ;
	output \g219406/_0_  ;
	output \g219407/_0_  ;
	output \g219408/_0_  ;
	output \g219409/_0_  ;
	output \g219410/_0_  ;
	output \g219411/_0_  ;
	output \g219412/_0_  ;
	output \g219413/_0_  ;
	output \g219414/_0_  ;
	output \g219415/_0_  ;
	output \g219416/_0_  ;
	output \g219417/_0_  ;
	output \g219418/_0_  ;
	output \g219419/_0_  ;
	output \g219420/_0_  ;
	output \g219421/_0_  ;
	output \g219422/_0_  ;
	output \g219423/_0_  ;
	output \g219424/_0_  ;
	output \g219425/_0_  ;
	output \g219426/_0_  ;
	output \g219427/_0_  ;
	output \g219428/_0_  ;
	output \g219429/_0_  ;
	output \g219430/_0_  ;
	output \g219431/_0_  ;
	output \g219432/_0_  ;
	output \g219433/_0_  ;
	output \g219434/_0_  ;
	output \g219435/_0_  ;
	output \g219436/_0_  ;
	output \g219437/_0_  ;
	output \g219438/_0_  ;
	output \g219439/_0_  ;
	output \g219440/_0_  ;
	output \g219441/_0_  ;
	output \g219442/_0_  ;
	output \g219443/_0_  ;
	output \g219444/_0_  ;
	output \g219445/_0_  ;
	output \g219446/_0_  ;
	output \g219447/_0_  ;
	output \g219449/_0_  ;
	output \g219450/_0_  ;
	output \g219451/_0_  ;
	output \g219452/_0_  ;
	output \g219453/_0_  ;
	output \g219454/_0_  ;
	output \g219455/_0_  ;
	output \g219456/_0_  ;
	output \g219457/_0_  ;
	output \g219458/_0_  ;
	output \g219464/u3_syn_7  ;
	output \g219496/u3_syn_4  ;
	output \g219512/u3_syn_4  ;
	output \g219526/u3_syn_4  ;
	output \g219549/u3_syn_4  ;
	output \g219571/u3_syn_4  ;
	output \g219588/u3_syn_4  ;
	output \g219603/u3_syn_4  ;
	output \g219621/u3_syn_4  ;
	output \g219636/_3_  ;
	output \g219652/u3_syn_4  ;
	output \g219676/_3_  ;
	output \g219686/_0_  ;
	output \g219689/_0_  ;
	output \g219694/_3_  ;
	output \g220062/_0_  ;
	output \g220068/_0_  ;
	output \g220069/_0_  ;
	output \g220072/_0_  ;
	output \g220084/_0_  ;
	output \g220149/_0_  ;
	output \g220162/_0_  ;
	output \g220317/_0_  ;
	output \g220360/_2_  ;
	output \g220368/_2_  ;
	output \g220369/_0_  ;
	output \g220370/_0_  ;
	output \g220371/_0_  ;
	output \g220372/_0_  ;
	output \g220376/_0_  ;
	output \g220390/_0_  ;
	output \g220395/_0_  ;
	output \g220499/_0_  ;
	output \g220500/_0_  ;
	output \g220501/_0_  ;
	output \g220502/_0_  ;
	output \g220503/_0_  ;
	output \g220504/_0_  ;
	output \g220505/_0_  ;
	output \g220506/_0_  ;
	output \g220507/_0_  ;
	output \g220508/_0_  ;
	output \g220509/_0_  ;
	output \g220510/_0_  ;
	output \g220511/_0_  ;
	output \g220512/_0_  ;
	output \g220513/_0_  ;
	output \g220514/_0_  ;
	output \g220515/_0_  ;
	output \g220516/_0_  ;
	output \g220517/_0_  ;
	output \g220518/_0_  ;
	output \g220519/_0_  ;
	output \g220520/_0_  ;
	output \g220521/_0_  ;
	output \g220522/_0_  ;
	output \g220523/_0_  ;
	output \g220524/_0_  ;
	output \g220525/_0_  ;
	output \g220526/_0_  ;
	output \g220527/_0_  ;
	output \g220528/_0_  ;
	output \g220529/_0_  ;
	output \g220530/_0_  ;
	output \g220531/_0_  ;
	output \g220532/_0_  ;
	output \g220533/_0_  ;
	output \g220534/_0_  ;
	output \g220535/_0_  ;
	output \g220557/_0_  ;
	output \g220558/_0_  ;
	output \g220559/_0_  ;
	output \g220560/_0_  ;
	output \g220561/_0_  ;
	output \g220562/_0_  ;
	output \g220563/_0_  ;
	output \g220564/_0_  ;
	output \g220565/_0_  ;
	output \g220566/_0_  ;
	output \g220567/_0_  ;
	output \g220568/_0_  ;
	output \g220569/_0_  ;
	output \g220570/_0_  ;
	output \g220571/_0_  ;
	output \g220572/_0_  ;
	output \g220573/_0_  ;
	output \g220574/_0_  ;
	output \g220575/_0_  ;
	output \g220576/_0_  ;
	output \g220577/_0_  ;
	output \g220578/_0_  ;
	output \g220579/_0_  ;
	output \g220580/_0_  ;
	output \g220581/_0_  ;
	output \g220582/_0_  ;
	output \g220583/_0_  ;
	output \g220584/_0_  ;
	output \g220585/_0_  ;
	output \g220586/_0_  ;
	output \g220587/_0_  ;
	output \g220588/_0_  ;
	output \g220589/_0_  ;
	output \g220590/_0_  ;
	output \g220591/_0_  ;
	output \g220592/_0_  ;
	output \g220593/_0_  ;
	output \g220594/_0_  ;
	output \g220595/_0_  ;
	output \g220596/_0_  ;
	output \g220597/_0_  ;
	output \g220598/_0_  ;
	output \g220599/_0_  ;
	output \g220600/_0_  ;
	output \g220601/_0_  ;
	output \g220602/_0_  ;
	output \g220603/_0_  ;
	output \g220604/_0_  ;
	output \g220605/_0_  ;
	output \g220606/_0_  ;
	output \g220607/_0_  ;
	output \g220608/_0_  ;
	output \g220609/_0_  ;
	output \g220610/_0_  ;
	output \g220611/_0_  ;
	output \g220612/_0_  ;
	output \g220613/_0_  ;
	output \g220614/_0_  ;
	output \g220615/_0_  ;
	output \g220616/_0_  ;
	output \g220617/_0_  ;
	output \g220618/_0_  ;
	output \g220619/_0_  ;
	output \g220620/_0_  ;
	output \g220621/_0_  ;
	output \g220622/_0_  ;
	output \g220623/_0_  ;
	output \g220624/_0_  ;
	output \g220625/_0_  ;
	output \g220626/_0_  ;
	output \g220627/_0_  ;
	output \g220628/_0_  ;
	output \g220629/_0_  ;
	output \g220630/_0_  ;
	output \g220631/_0_  ;
	output \g220632/_0_  ;
	output \g220633/_0_  ;
	output \g220634/_0_  ;
	output \g220635/_0_  ;
	output \g220636/_0_  ;
	output \g220637/_0_  ;
	output \g220638/_0_  ;
	output \g220639/_0_  ;
	output \g220640/_0_  ;
	output \g220641/_0_  ;
	output \g220642/_0_  ;
	output \g220643/_0_  ;
	output \g220644/_0_  ;
	output \g220645/_0_  ;
	output \g220646/_0_  ;
	output \g220647/_0_  ;
	output \g220648/_0_  ;
	output \g220649/_0_  ;
	output \g220650/_0_  ;
	output \g220651/_0_  ;
	output \g220652/_0_  ;
	output \g220653/_0_  ;
	output \g220654/_0_  ;
	output \g220655/_0_  ;
	output \g220656/_0_  ;
	output \g220657/_0_  ;
	output \g220658/_0_  ;
	output \g220659/_0_  ;
	output \g220660/_0_  ;
	output \g220661/_0_  ;
	output \g220662/_0_  ;
	output \g220663/_0_  ;
	output \g220664/_0_  ;
	output \g220665/_0_  ;
	output \g220666/_0_  ;
	output \g220674/_0_  ;
	output \g220679/u3_syn_7  ;
	output \g220711/u3_syn_4  ;
	output \g220726/u3_syn_4  ;
	output \g220739/u3_syn_4  ;
	output \g220751/u3_syn_4  ;
	output \g220759/u3_syn_4  ;
	output \g220773/u3_syn_4  ;
	output \g220782/u3_syn_4  ;
	output \g220805/u3_syn_4  ;
	output \g220828/u3_syn_4  ;
	output \g220921/_0_  ;
	output \g220930/u3_syn_4  ;
	output \g220949/_3_  ;
	output \g220994/_3_  ;
	output \g221207/_0_  ;
	output \g221213/_0_  ;
	output \g221223/_0_  ;
	output \g221224/_0_  ;
	output \g221225/_0_  ;
	output \g221226/_0_  ;
	output \g221231/_0_  ;
	output \g221232/_0_  ;
	output \g221234/_0_  ;
	output \g221235/_0_  ;
	output \g221246/_2_  ;
	output \g221249/_2_  ;
	output \g221265/_0_  ;
	output \g221287/_0_  ;
	output \g221325/_0_  ;
	output \g221326/_0_  ;
	output \g221447/_0_  ;
	output \g221449/_0_  ;
	output \g221452/_0_  ;
	output \g221469/_0_  ;
	output \g221473/_0_  ;
	output \g221503/_0_  ;
	output \g221510/_0_  ;
	output \g221512/_0_  ;
	output \g221516/_0_  ;
	output \g221517/_0_  ;
	output \g221524/_0_  ;
	output \g221530/_0_  ;
	output \g221592/_0_  ;
	output \g221593/_0_  ;
	output \g221634/u3_syn_4  ;
	output \g221669/u3_syn_4  ;
	output \g221789/u3_syn_4  ;
	output \g221813/u3_syn_4  ;
	output \g221829/u3_syn_4  ;
	output \g221861/u3_syn_4  ;
	output \g221876/_0_  ;
	output \g221935/_0_  ;
	output \g221944/_3_  ;
	output \g230200/_0_  ;
	output \g230201/_0_  ;
	output \g230205/_0_  ;
	output \g230295/_0_  ;
	output \g230297/_0_  ;
	output \g230298/_0_  ;
	output \g230300/_0_  ;
	output \g230302/_0_  ;
	output \g230303/_0_  ;
	output \g230343/_0_  ;
	output \g230368/_0_  ;
	output \g230511/_0_  ;
	output \g230531/_0_  ;
	output \g230635/_2_  ;
	output \g230661/_0_  ;
	output \g230715/_1__syn_2  ;
	output \g230731/_0_  ;
	output \g230766/_0_  ;
	output \g230784/_0_  ;
	output \g230785/_0_  ;
	output \g230786/_0_  ;
	output \g230787/_0_  ;
	output \g230797/_0_  ;
	output \g230798/_0_  ;
	output \g230803/_0_  ;
	output \g230804/_00_  ;
	output \g230805/_00_  ;
	output \g230806/_00_  ;
	output \g230807/_00_  ;
	output \g230808/_00_  ;
	output \g230809/_00_  ;
	output \g230815/_0_  ;
	output \g230816/_2_  ;
	output \g230817/_2_  ;
	output \g230829/_0_  ;
	output \g230834/_0_  ;
	output \g230835/_0_  ;
	output \g230836/_0_  ;
	output \g230837/_0_  ;
	output \g230844/_0_  ;
	output \g230863/_3_  ;
	output \g230864/_3_  ;
	output \g230870/_0_  ;
	output \g230988/_3_  ;
	output \g231010/_3_  ;
	output \g231016/_3_  ;
	output \g231042/_3_  ;
	output \g231471/_0_  ;
	output \g231472/_0_  ;
	output \g231476/_3_  ;
	output \g231480/_3_  ;
	output \g231484/_3_  ;
	output \g231504/_0_  ;
	output \g231532/_0_  ;
	output \g231542/_0_  ;
	output \g231560/_1_  ;
	output \g231578/_1_  ;
	output \g231580/_0_  ;
	output \g231590/_1__syn_2  ;
	output \g231615/_0_  ;
	output \g231623/_1_  ;
	output \g231634/_2_  ;
	output \g231635/_0_  ;
	output \g231638/_2_  ;
	output \g231640/_0_  ;
	output \g231653/_2_  ;
	output \g231787/_0_  ;
	output \g231931/_0_  ;
	output \g231939/_3_  ;
	output \g231940/_0_  ;
	output \g231951/_0_  ;
	output \g231955/_0_  ;
	output \g231956/_0_  ;
	output \g231959/_2_  ;
	output \g231960/_0_  ;
	output \g231964/_0_  ;
	output \g231965/_0_  ;
	output \g231975/_0_  ;
	output \g231986/_1_  ;
	output \g231987/_1_  ;
	output \g231989/_1_  ;
	output \g231990/_1_  ;
	output \g231991/_0_  ;
	output \g231992/_0_  ;
	output \g231995/_0_  ;
	output \g231998/_0_  ;
	output \g231999/_0_  ;
	output \g232002/_3_  ;
	output \g232035/u3_syn_4  ;
	output \g232038/u3_syn_4  ;
	output \g232046/u3_syn_4  ;
	output \g232054/u3_syn_4  ;
	output \g232062/u3_syn_4  ;
	output \g232070/u3_syn_4  ;
	output \g232078/u3_syn_4  ;
	output \g232079/u3_syn_4  ;
	output \g232087/u3_syn_4  ;
	output \g232096/u3_syn_4  ;
	output \g232104/u3_syn_4  ;
	output \g232112/u3_syn_4  ;
	output \g232120/u3_syn_4  ;
	output \g232128/u3_syn_4  ;
	output \g232136/u3_syn_4  ;
	output \g232144/u3_syn_4  ;
	output \g232152/u3_syn_4  ;
	output \g232161/u3_syn_4  ;
	output \g232169/u3_syn_4  ;
	output \g232177/u3_syn_4  ;
	output \g232185/u3_syn_4  ;
	output \g232186/u3_syn_4  ;
	output \g232194/u3_syn_4  ;
	output \g232202/u3_syn_4  ;
	output \g232210/u3_syn_4  ;
	output \g232218/u3_syn_4  ;
	output \g232226/u3_syn_4  ;
	output \g232234/u3_syn_4  ;
	output \g232242/u3_syn_4  ;
	output \g232251/u3_syn_4  ;
	output \g232259/u3_syn_4  ;
	output \g232267/u3_syn_4  ;
	output \g232275/u3_syn_4  ;
	output \g232283/u3_syn_4  ;
	output \g232291/u3_syn_4  ;
	output \g232299/u3_syn_4  ;
	output \g232307/u3_syn_4  ;
	output \g232315/u3_syn_4  ;
	output \g232324/u3_syn_4  ;
	output \g232332/u3_syn_4  ;
	output \g232341/u3_syn_4  ;
	output \g232349/u3_syn_4  ;
	output \g232357/u3_syn_4  ;
	output \g232366/u3_syn_4  ;
	output \g232374/u3_syn_4  ;
	output \g232382/u3_syn_4  ;
	output \g232390/u3_syn_4  ;
	output \g232398/u3_syn_4  ;
	output \g232406/u3_syn_4  ;
	output \g232414/u3_syn_4  ;
	output \g232422/u3_syn_4  ;
	output \g232427/u3_syn_4  ;
	output \g232431/u3_syn_4  ;
	output \g232439/u3_syn_4  ;
	output \g232444/u3_syn_4  ;
	output \g232452/u3_syn_4  ;
	output \g232461/u3_syn_4  ;
	output \g232471/u3_syn_4  ;
	output \g232479/u3_syn_4  ;
	output \g232487/u3_syn_4  ;
	output \g232495/u3_syn_4  ;
	output \g232503/u3_syn_4  ;
	output \g232506/u3_syn_4  ;
	output \g232514/u3_syn_4  ;
	output \g232527/u3_syn_4  ;
	output \g232530/u3_syn_4  ;
	output \g232536/u3_syn_4  ;
	output \g232544/u3_syn_4  ;
	output \g232551/u3_syn_4  ;
	output \g232557/u3_syn_4  ;
	output \g232568/u3_syn_4  ;
	output \g232576/u3_syn_4  ;
	output \g232585/u3_syn_4  ;
	output \g232593/u3_syn_4  ;
	output \g232597/u3_syn_4  ;
	output \g232609/u3_syn_4  ;
	output \g232617/u3_syn_4  ;
	output \g232625/u3_syn_4  ;
	output \g232633/u3_syn_4  ;
	output \g232641/u3_syn_4  ;
	output \g232649/u3_syn_4  ;
	output \g232657/u3_syn_4  ;
	output \g232665/u3_syn_4  ;
	output \g232673/u3_syn_4  ;
	output \g232681/u3_syn_4  ;
	output \g232689/u3_syn_4  ;
	output \g232697/u3_syn_4  ;
	output \g232705/u3_syn_4  ;
	output \g232713/u3_syn_4  ;
	output \g232717/u3_syn_4  ;
	output \g232729/u3_syn_4  ;
	output \g232737/u3_syn_4  ;
	output \g232745/u3_syn_4  ;
	output \g232749/u3_syn_4  ;
	output \g232761/u3_syn_4  ;
	output \g232768/u3_syn_4  ;
	output \g232777/u3_syn_4  ;
	output \g232785/u3_syn_4  ;
	output \g232793/u3_syn_4  ;
	output \g232801/u3_syn_4  ;
	output \g232809/u3_syn_4  ;
	output \g232815/u3_syn_4  ;
	output \g232823/u3_syn_4  ;
	output \g232833/u3_syn_4  ;
	output \g232841/u3_syn_4  ;
	output \g232846/u3_syn_4  ;
	output \g232851/u3_syn_4  ;
	output \g232865/u3_syn_4  ;
	output \g232873/u3_syn_4  ;
	output \g232881/u3_syn_4  ;
	output \g232882/u3_syn_4  ;
	output \g232895/u3_syn_4  ;
	output \g232904/u3_syn_4  ;
	output \g232913/u3_syn_4  ;
	output \g232921/u3_syn_4  ;
	output \g232928/u3_syn_4  ;
	output \g232934/u3_syn_4  ;
	output \g232945/u3_syn_4  ;
	output \g232953/u3_syn_4  ;
	output \g232954/u3_syn_4  ;
	output \g232969/u3_syn_4  ;
	output \g232977/u3_syn_4  ;
	output \g232981/u3_syn_4  ;
	output \g232993/u3_syn_4  ;
	output \g232995/u3_syn_4  ;
	output \g233009/u3_syn_4  ;
	output \g233017/u3_syn_4  ;
	output \g233025/u3_syn_4  ;
	output \g233033/u3_syn_4  ;
	output \g233041/u3_syn_4  ;
	output \g233047/u3_syn_4  ;
	output \g233057/u3_syn_4  ;
	output \g233065/u3_syn_4  ;
	output \g233073/u3_syn_4  ;
	output \g233081/u3_syn_4  ;
	output \g233087/u3_syn_4  ;
	output \g233097/u3_syn_4  ;
	output \g233105/u3_syn_4  ;
	output \g233113/u3_syn_4  ;
	output \g233121/u3_syn_4  ;
	output \g233128/u3_syn_4  ;
	output \g233134/u3_syn_4  ;
	output \g233144/u3_syn_4  ;
	output \g233153/u3_syn_4  ;
	output \g233161/u3_syn_4  ;
	output \g233169/u3_syn_4  ;
	output \g233177/u3_syn_4  ;
	output \g233185/u3_syn_4  ;
	output \g233193/u3_syn_4  ;
	output \g233201/u3_syn_4  ;
	output \g233209/u3_syn_4  ;
	output \g233217/u3_syn_4  ;
	output \g233219/u3_syn_4  ;
	output \g233229/u3_syn_4  ;
	output \g233241/u3_syn_4  ;
	output \g233249/u3_syn_4  ;
	output \g233257/u3_syn_4  ;
	output \g233265/u3_syn_4  ;
	output \g233273/u3_syn_4  ;
	output \g233281/u3_syn_4  ;
	output \g233289/u3_syn_4  ;
	output \g233297/u3_syn_4  ;
	output \g233305/u3_syn_4  ;
	output \g233313/u3_syn_4  ;
	output \g233321/u3_syn_4  ;
	output \g233329/u3_syn_4  ;
	output \g233337/u3_syn_4  ;
	output \g233345/u3_syn_4  ;
	output \g233353/u3_syn_4  ;
	output \g233361/u3_syn_4  ;
	output \g233369/u3_syn_4  ;
	output \g233377/u3_syn_4  ;
	output \g233382/u3_syn_4  ;
	output \g233392/u3_syn_4  ;
	output \g233394/u3_syn_4  ;
	output \g233409/u3_syn_4  ;
	output \g233417/u3_syn_4  ;
	output \g233425/u3_syn_4  ;
	output \g233433/u3_syn_4  ;
	output \g233441/u3_syn_4  ;
	output \g233449/u3_syn_4  ;
	output \g233453/u3_syn_4  ;
	output \g233465/u3_syn_4  ;
	output \g233473/u3_syn_4  ;
	output \g233481/u3_syn_4  ;
	output \g233489/u3_syn_4  ;
	output \g233497/u3_syn_4  ;
	output \g233505/u3_syn_4  ;
	output \g233513/u3_syn_4  ;
	output \g233516/u3_syn_4  ;
	output \g233529/u3_syn_4  ;
	output \g233531/u3_syn_4  ;
	output \g233546/u3_syn_4  ;
	output \g233554/u3_syn_4  ;
	output \g233562/u3_syn_4  ;
	output \g233570/u3_syn_4  ;
	output \g233578/u3_syn_4  ;
	output \g233586/u3_syn_4  ;
	output \g233594/u3_syn_4  ;
	output \g233602/u3_syn_4  ;
	output \g233603/u3_syn_4  ;
	output \g233618/u3_syn_4  ;
	output \g233626/u3_syn_4  ;
	output \g233634/u3_syn_4  ;
	output \g233642/u3_syn_4  ;
	output \g233650/u3_syn_4  ;
	output \g233658/u3_syn_4  ;
	output \g233666/u3_syn_4  ;
	output \g233674/u3_syn_4  ;
	output \g233682/u3_syn_4  ;
	output \g233690/u3_syn_4  ;
	output \g233698/u3_syn_4  ;
	output \g233706/u3_syn_4  ;
	output \g233714/u3_syn_4  ;
	output \g233722/u3_syn_4  ;
	output \g233730/u3_syn_4  ;
	output \g233738/u3_syn_4  ;
	output \g233746/u3_syn_4  ;
	output \g233754/u3_syn_4  ;
	output \g233762/u3_syn_4  ;
	output \g233770/u3_syn_4  ;
	output \g233778/u3_syn_4  ;
	output \g233783/u3_syn_4  ;
	output \g233794/u3_syn_4  ;
	output \g233802/u3_syn_4  ;
	output \g233806/u3_syn_4  ;
	output \g233818/u3_syn_4  ;
	output \g233826/u3_syn_4  ;
	output \g233828/u3_syn_4  ;
	output \g233838/u3_syn_4  ;
	output \g233850/u3_syn_4  ;
	output \g233858/u3_syn_4  ;
	output \g233860/u3_syn_4  ;
	output \g233870/u3_syn_4  ;
	output \g233881/u3_syn_4  ;
	output \g233890/u3_syn_4  ;
	output \g233899/u3_syn_4  ;
	output \g233908/u3_syn_4  ;
	output \g233917/u3_syn_4  ;
	output \g233919/u3_syn_4  ;
	output \g233927/u3_syn_4  ;
	output \g233935/u3_syn_4  ;
	output \g233943/u3_syn_4  ;
	output \g233945/u3_syn_4  ;
	output \g233953/u3_syn_4  ;
	output \g233961/u3_syn_4  ;
	output \g233969/u3_syn_4  ;
	output \g233977/u3_syn_4  ;
	output \g233985/u3_syn_4  ;
	output \g233993/u3_syn_4  ;
	output \g234001/u3_syn_4  ;
	output \g234008/u3_syn_4  ;
	output \g234009/u3_syn_4  ;
	output \g234024/u3_syn_4  ;
	output \g234032/u3_syn_4  ;
	output \g234038/u3_syn_4  ;
	output \g234056/u3_syn_4  ;
	output \g234063/u3_syn_4  ;
	output \g234071/u3_syn_4  ;
	output \g234079/u3_syn_4  ;
	output \g234098/u3_syn_4  ;
	output \g234106/u3_syn_4  ;
	output \g234114/u3_syn_4  ;
	output \g234122/u3_syn_4  ;
	output \g234130/u3_syn_4  ;
	output \g234138/u3_syn_4  ;
	output \g234145/u3_syn_4  ;
	output \g234156/u3_syn_4  ;
	output \g234162/u3_syn_4  ;
	output \g234171/u3_syn_4  ;
	output \g234183/u3_syn_4  ;
	output \g234248/u3_syn_4  ;
	output \g234265/u3_syn_4  ;
	output \g234273/u3_syn_4  ;
	output \g234281/u3_syn_4  ;
	output \g234289/u3_syn_4  ;
	output \g234297/u3_syn_4  ;
	output \g234306/u3_syn_4  ;
	output \g234314/u3_syn_4  ;
	output \g234322/u3_syn_4  ;
	output \g234331/u3_syn_4  ;
	output \g234339/u3_syn_4  ;
	output \g234347/u3_syn_4  ;
	output \g234355/u3_syn_4  ;
	output \g234363/u3_syn_4  ;
	output \g234371/u3_syn_4  ;
	output \g234379/u3_syn_4  ;
	output \g234387/u3_syn_4  ;
	output \g234395/u3_syn_4  ;
	output \g234403/u3_syn_4  ;
	output \g234411/u3_syn_4  ;
	output \g234419/u3_syn_4  ;
	output \g234427/u3_syn_4  ;
	output \g234435/u3_syn_4  ;
	output \g234443/u3_syn_4  ;
	output \g234451/u3_syn_4  ;
	output \g234459/u3_syn_4  ;
	output \g234467/u3_syn_4  ;
	output \g234475/u3_syn_4  ;
	output \g234483/u3_syn_4  ;
	output \g234491/u3_syn_4  ;
	output \g234499/u3_syn_4  ;
	output \g234507/u3_syn_4  ;
	output \g234515/u3_syn_4  ;
	output \g234523/u3_syn_4  ;
	output \g234531/u3_syn_4  ;
	output \g234539/u3_syn_4  ;
	output \g234547/u3_syn_4  ;
	output \g234555/u3_syn_4  ;
	output \g234563/u3_syn_4  ;
	output \g234571/u3_syn_4  ;
	output \g234579/u3_syn_4  ;
	output \g234587/u3_syn_4  ;
	output \g234595/u3_syn_4  ;
	output \g234604/u3_syn_4  ;
	output \g234612/u3_syn_4  ;
	output \g234620/u3_syn_4  ;
	output \g234628/u3_syn_4  ;
	output \g234636/u3_syn_4  ;
	output \g234644/u3_syn_4  ;
	output \g234652/u3_syn_4  ;
	output \g234660/u3_syn_4  ;
	output \g234668/u3_syn_4  ;
	output \g234676/u3_syn_4  ;
	output \g234684/u3_syn_4  ;
	output \g234692/u3_syn_4  ;
	output \g234700/u3_syn_4  ;
	output \g234708/u3_syn_4  ;
	output \g234716/u3_syn_4  ;
	output \g234725/u3_syn_4  ;
	output \g234733/u3_syn_4  ;
	output \g234741/u3_syn_4  ;
	output \g234749/u3_syn_4  ;
	output \g234757/u3_syn_4  ;
	output \g234765/u3_syn_4  ;
	output \g234773/u3_syn_4  ;
	output \g234781/u3_syn_4  ;
	output \g234789/u3_syn_4  ;
	output \g234798/u3_syn_4  ;
	output \g234806/u3_syn_4  ;
	output \g234814/u3_syn_4  ;
	output \g234822/u3_syn_4  ;
	output \g234830/u3_syn_4  ;
	output \g234838/u3_syn_4  ;
	output \g235911/u3_syn_4  ;
	output \g235912/u3_syn_4  ;
	output \g235920/u3_syn_4  ;
	output \g235928/u3_syn_4  ;
	output \g235936/u3_syn_4  ;
	output \g235944/u3_syn_4  ;
	output \g235952/u3_syn_4  ;
	output \g235960/u3_syn_4  ;
	output \g235968/u3_syn_4  ;
	output \g235976/u3_syn_4  ;
	output \g235984/u3_syn_4  ;
	output \g235992/u3_syn_4  ;
	output \g236000/u3_syn_4  ;
	output \g236008/u3_syn_4  ;
	output \g236016/u3_syn_4  ;
	output \g236021/u3_syn_4  ;
	output \g236025/u3_syn_4  ;
	output \g236033/u3_syn_4  ;
	output \g236041/u3_syn_4  ;
	output \g236049/u3_syn_4  ;
	output \g236057/u3_syn_4  ;
	output \g236065/u3_syn_4  ;
	output \g236073/u3_syn_4  ;
	output \g236081/u3_syn_4  ;
	output \g236089/u3_syn_4  ;
	output \g236097/u3_syn_4  ;
	output \g236105/u3_syn_4  ;
	output \g236113/u3_syn_4  ;
	output \g236121/u3_syn_4  ;
	output \g236129/u3_syn_4  ;
	output \g236137/u3_syn_4  ;
	output \g236145/u3_syn_4  ;
	output \g236153/u3_syn_4  ;
	output \g236161/u3_syn_4  ;
	output \g236169/u3_syn_4  ;
	output \g236177/u3_syn_4  ;
	output \g236185/u3_syn_4  ;
	output \g236193/u3_syn_4  ;
	output \g236196/u3_syn_4  ;
	output \g236198/u3_syn_4  ;
	output \g236203/u3_syn_4  ;
	output \g236211/u3_syn_4  ;
	output \g236219/u3_syn_4  ;
	output \g236220/u3_syn_4  ;
	output \g236229/u3_syn_4  ;
	output \g236232/u3_syn_4  ;
	output \g236238/u3_syn_4  ;
	output \g236246/u3_syn_4  ;
	output \g236255/u3_syn_4  ;
	output \g236263/u3_syn_4  ;
	output \g236271/u3_syn_4  ;
	output \g236275/u3_syn_4  ;
	output \g236280/u3_syn_4  ;
	output \g236288/u3_syn_4  ;
	output \g236296/u3_syn_4  ;
	output \g236304/u3_syn_4  ;
	output \g236305/u3_syn_4  ;
	output \g236306/u3_syn_4  ;
	output \g236315/u3_syn_4  ;
	output \g236323/u3_syn_4  ;
	output \g236331/u3_syn_4  ;
	output \g236334/u3_syn_4  ;
	output \g236340/u3_syn_4  ;
	output \g236348/u3_syn_4  ;
	output \g236357/u3_syn_4  ;
	output \g236359/u3_syn_4  ;
	output \g236367/u3_syn_4  ;
	output \g236374/u3_syn_4  ;
	output \g236376/u3_syn_4  ;
	output \g236377/u3_syn_4  ;
	output \g236385/u3_syn_4  ;
	output \g236393/u3_syn_4  ;
	output \g236402/u3_syn_4  ;
	output \g236410/u3_syn_4  ;
	output \g236419/u3_syn_4  ;
	output \g236427/u3_syn_4  ;
	output \g236433/u3_syn_4  ;
	output \g236436/u3_syn_4  ;
	output \g236444/u3_syn_4  ;
	output \g236452/u3_syn_4  ;
	output \g236460/u3_syn_4  ;
	output \g236468/u3_syn_4  ;
	output \g236476/u3_syn_4  ;
	output \g236484/u3_syn_4  ;
	output \g236492/u3_syn_4  ;
	output \g236500/u3_syn_4  ;
	output \g236508/u3_syn_4  ;
	output \g236516/u3_syn_4  ;
	output \g236518/u3_syn_4  ;
	output \g236525/u3_syn_4  ;
	output \g236533/u3_syn_4  ;
	output \g236542/u3_syn_4  ;
	output \g236550/u3_syn_4  ;
	output \g236559/u3_syn_4  ;
	output \g236567/u3_syn_4  ;
	output \g236575/u3_syn_4  ;
	output \g236583/u3_syn_4  ;
	output \g236591/u3_syn_4  ;
	output \g236599/u3_syn_4  ;
	output \g236607/u3_syn_4  ;
	output \g236608/u3_syn_4  ;
	output \g236616/u3_syn_4  ;
	output \g236624/u3_syn_4  ;
	output \g236632/u3_syn_4  ;
	output \g236640/u3_syn_4  ;
	output \g236647/u3_syn_4  ;
	output \g236649/u3_syn_4  ;
	output \g236659/u3_syn_4  ;
	output \g236671/u3_syn_4  ;
	output \g236677/u3_syn_4  ;
	output \g236688/u3_syn_4  ;
	output \g236696/u3_syn_4  ;
	output \g236705/u3_syn_4  ;
	output \g236712/u3_syn_4  ;
	output \g236718/u3_syn_4  ;
	output \g236729/u3_syn_4  ;
	output \g236732/u3_syn_4  ;
	output \g236745/u3_syn_4  ;
	output \g236753/u3_syn_4  ;
	output \g236761/u3_syn_4  ;
	output \g236769/u3_syn_4  ;
	output \g236777/u3_syn_4  ;
	output \g236779/u3_syn_4  ;
	output \g236788/u3_syn_4  ;
	output \g236800/u3_syn_4  ;
	output \g236802/u3_syn_4  ;
	output \g236805/u3_syn_4  ;
	output \g236813/u3_syn_4  ;
	output \g236825/u3_syn_4  ;
	output \g236829/u3_syn_4  ;
	output \g236837/u3_syn_4  ;
	output \g236849/u3_syn_4  ;
	output \g236854/u3_syn_4  ;
	output \g236860/u3_syn_4  ;
	output \g236872/u3_syn_4  ;
	output \g236878/u3_syn_4  ;
	output \g236884/u3_syn_4  ;
	output \g236896/u3_syn_4  ;
	output \g236903/u3_syn_4  ;
	output \g236908/u3_syn_4  ;
	output \g236920/u3_syn_4  ;
	output \g236930/u3_syn_4  ;
	output \g236939/u3_syn_4  ;
	output \g236947/u3_syn_4  ;
	output \g236949/u3_syn_4  ;
	output \g236956/u3_syn_4  ;
	output \g236962/u3_syn_4  ;
	output \g236965/u3_syn_4  ;
	output \g236980/u3_syn_4  ;
	output \g236988/u3_syn_4  ;
	output \g236989/u3_syn_4  ;
	output \g237004/u3_syn_4  ;
	output \g237005/u3_syn_4  ;
	output \g237020/u3_syn_4  ;
	output \g237021/u3_syn_4  ;
	output \g237033/u3_syn_4  ;
	output \g237044/u3_syn_4  ;
	output \g237045/u3_syn_4  ;
	output \g237056/u3_syn_4  ;
	output \g237068/u3_syn_4  ;
	output \g237076/u3_syn_4  ;
	output \g237084/u3_syn_4  ;
	output \g237092/u3_syn_4  ;
	output \g237095/u3_syn_4  ;
	output \g237107/u3_syn_4  ;
	output \g237110/u3_syn_4  ;
	output \g237119/u3_syn_4  ;
	output \g237131/u3_syn_4  ;
	output \g237135/u3_syn_4  ;
	output \g237148/u3_syn_4  ;
	output \g237152/u3_syn_4  ;
	output \g237165/u3_syn_4  ;
	output \g237168/u3_syn_4  ;
	output \g237180/u3_syn_4  ;
	output \g237185/u3_syn_4  ;
	output \g237192/u3_syn_4  ;
	output \g237204/u3_syn_4  ;
	output \g237209/u3_syn_4  ;
	output \g237215/u3_syn_4  ;
	output \g237229/u3_syn_4  ;
	output \g237231/u3_syn_4  ;
	output \g237245/u3_syn_4  ;
	output \g237251/u3_syn_4  ;
	output \g237260/u3_syn_4  ;
	output \g237262/u3_syn_4  ;
	output \g237277/u3_syn_4  ;
	output \g237281/u3_syn_4  ;
	output \g237293/u3_syn_4  ;
	output \g237294/u3_syn_4  ;
	output \g237310/u3_syn_4  ;
	output \g237311/u3_syn_4  ;
	output \g237323/u3_syn_4  ;
	output \g237334/u3_syn_4  ;
	output \g237342/u3_syn_4  ;
	output \g237350/u3_syn_4  ;
	output \g237353/u3_syn_4  ;
	output \g237359/u3_syn_4  ;
	output \g237367/u3_syn_4  ;
	output \g237368/u3_syn_4  ;
	output \g237378/u3_syn_4  ;
	output \g237391/u3_syn_4  ;
	output \g237392/u3_syn_4  ;
	output \g237403/u3_syn_4  ;
	output \g237415/u3_syn_4  ;
	output \g237417/u3_syn_4  ;
	output \g237431/u3_syn_4  ;
	output \g237439/u3_syn_4  ;
	output \g237440/u3_syn_4  ;
	output \g237454/u3_syn_4  ;
	output \g237457/u3_syn_4  ;
	output \g237472/u3_syn_4  ;
	output \g237480/u3_syn_4  ;
	output \g237488/u3_syn_4  ;
	output \g237496/u3_syn_4  ;
	output \g237499/u3_syn_4  ;
	output \g237512/u3_syn_4  ;
	output \g237515/u3_syn_4  ;
	output \g237525/u3_syn_4  ;
	output \g237529/u3_syn_4  ;
	output \g237535/u3_syn_4  ;
	output \g237541/u3_syn_4  ;
	output \g237553/u3_syn_4  ;
	output \g237561/u3_syn_4  ;
	output \g237569/u3_syn_4  ;
	output \g237575/u3_syn_4  ;
	output \g237578/u3_syn_4  ;
	output \g237581/u3_syn_4  ;
	output \g237591/u3_syn_4  ;
	output \g237602/u3_syn_4  ;
	output \g237610/u3_syn_4  ;
	output \g237617/u3_syn_4  ;
	output \g237623/u3_syn_4  ;
	output \g237633/u3_syn_4  ;
	output \g237635/u3_syn_4  ;
	output \g237648/u3_syn_4  ;
	output \g237658/u3_syn_4  ;
	output \g237659/u3_syn_4  ;
	output \g237660/u3_syn_4  ;
	output \g237668/u3_syn_4  ;
	output \g237675/u3_syn_4  ;
	output \g237684/u3_syn_4  ;
	output \g237692/u3_syn_4  ;
	output \g237693/u3_syn_4  ;
	output \g237705/u3_syn_4  ;
	output \g237716/u3_syn_4  ;
	output \g237717/u3_syn_4  ;
	output \g237729/u3_syn_4  ;
	output \g237740/u3_syn_4  ;
	output \g237741/u3_syn_4  ;
	output \g237756/u3_syn_4  ;
	output \g237764/u3_syn_4  ;
	output \g237768/u3_syn_4  ;
	output \g237780/u3_syn_4  ;
	output \g237782/u3_syn_4  ;
	output \g237792/u3_syn_4  ;
	output \g237804/u3_syn_4  ;
	output \g237812/u3_syn_4  ;
	output \g237820/u3_syn_4  ;
	output \g237828/u3_syn_4  ;
	output \g237836/u3_syn_4  ;
	output \g237844/u3_syn_4  ;
	output \g237852/u3_syn_4  ;
	output \g237860/u3_syn_4  ;
	output \g237868/u3_syn_4  ;
	output \g237876/u3_syn_4  ;
	output \g237884/u3_syn_4  ;
	output \g237888/u3_syn_4  ;
	output \g237895/u3_syn_4  ;
	output \g237907/u3_syn_4  ;
	output \g237916/u3_syn_4  ;
	output \g237924/u3_syn_4  ;
	output \g237931/u3_syn_4  ;
	output \g237940/u3_syn_4  ;
	output \g237949/u3_syn_4  ;
	output \g237950/u3_syn_4  ;
	output \g237955/u3_syn_4  ;
	output \g237961/u3_syn_4  ;
	output \g237965/u3_syn_4  ;
	output \g237975/u3_syn_4  ;
	output \g237983/u3_syn_4  ;
	output \g237989/u3_syn_4  ;
	output \g237999/u3_syn_4  ;
	output \g238007/u3_syn_4  ;
	output \g238015/u3_syn_4  ;
	output \g238017/u3_syn_4  ;
	output \g238033/u3_syn_4  ;
	output \g238035/u3_syn_4  ;
	output \g238049/u3_syn_4  ;
	output \g238057/u3_syn_4  ;
	output \g238065/u3_syn_4  ;
	output \g238072/u3_syn_4  ;
	output \g238081/u3_syn_4  ;
	output \g238082/u3_syn_4  ;
	output \g238097/u3_syn_4  ;
	output \g238105/u3_syn_4  ;
	output \g238113/u3_syn_4  ;
	output \g238114/u3_syn_4  ;
	output \g238129/u3_syn_4  ;
	output \g238137/u3_syn_4  ;
	output \g238145/u3_syn_4  ;
	output \g238153/u3_syn_4  ;
	output \g238161/u3_syn_4  ;
	output \g238163/u3_syn_4  ;
	output \g238177/u3_syn_4  ;
	output \g238179/u3_syn_4  ;
	output \g238194/u3_syn_4  ;
	output \g238197/u3_syn_4  ;
	output \g238209/u3_syn_4  ;
	output \g238213/u3_syn_4  ;
	output \g238225/u3_syn_4  ;
	output \g238229/u3_syn_4  ;
	output \g238237/u3_syn_4  ;
	output \g238250/u3_syn_4  ;
	output \g238257/u3_syn_4  ;
	output \g238263/u3_syn_4  ;
	output \g238269/u3_syn_4  ;
	output \g238282/u3_syn_4  ;
	output \g238285/u3_syn_4  ;
	output \g238298/u3_syn_4  ;
	output \g238301/u3_syn_4  ;
	output \g238314/u3_syn_4  ;
	output \g238316/u3_syn_4  ;
	output \g238329/u3_syn_4  ;
	output \g238338/u3_syn_4  ;
	output \g238346/u3_syn_4  ;
	output \g238351/u3_syn_4  ;
	output \g238356/u3_syn_4  ;
	output \g238368/u3_syn_4  ;
	output \g238378/u3_syn_4  ;
	output \g238386/u3_syn_4  ;
	output \g238394/u3_syn_4  ;
	output \g238402/u3_syn_4  ;
	output \g238409/u3_syn_4  ;
	output \g238412/u3_syn_4  ;
	output \g238427/u3_syn_4  ;
	output \g238429/u3_syn_4  ;
	output \g238443/u3_syn_4  ;
	output \g238448/u3_syn_4  ;
	output \g238457/u3_syn_4  ;
	output \g238460/u3_syn_4  ;
	output \g238472/u3_syn_4  ;
	output \g238484/u3_syn_4  ;
	output \g238492/u3_syn_4  ;
	output \g238500/u3_syn_4  ;
	output \g238505/u3_syn_4  ;
	output \g238516/u3_syn_4  ;
	output \g238524/u3_syn_4  ;
	output \g238532/u3_syn_4  ;
	output \g238534/u3_syn_4  ;
	output \g238544/u3_syn_4  ;
	output \g238549/u3_syn_4  ;
	output \g238550/u3_syn_4  ;
	output \g238565/u3_syn_4  ;
	output \g238566/u3_syn_4  ;
	output \g238582/u3_syn_4  ;
	output \g238583/u3_syn_4  ;
	output \g238594/u3_syn_4  ;
	output \g238606/u3_syn_4  ;
	output \g238614/u3_syn_4  ;
	output \g238615/u3_syn_4  ;
	output \g238619/u3_syn_4  ;
	output \g238631/u3_syn_4  ;
	output \g238639/u3_syn_4  ;
	output \g238647/u3_syn_4  ;
	output \g238649/u3_syn_4  ;
	output \g238659/u3_syn_4  ;
	output \g238670/u3_syn_4  ;
	output \g238671/u3_syn_4  ;
	output \g238680/u3_syn_4  ;
	output \g238688/u3_syn_4  ;
	output \g238691/u3_syn_4  ;
	output \g238696/u3_syn_4  ;
	output \g238705/u3_syn_4  ;
	output \g238708/u3_syn_4  ;
	output \g238721/u3_syn_4  ;
	output \g238724/u3_syn_4  ;
	output \g238736/u3_syn_4  ;
	output \g238745/u3_syn_4  ;
	output \g238753/u3_syn_4  ;
	output \g238757/u3_syn_4  ;
	output \g238764/u3_syn_4  ;
	output \g238776/u3_syn_4  ;
	output \g238781/u3_syn_4  ;
	output \g238787/u3_syn_4  ;
	output \g238799/u3_syn_4  ;
	output \g238807/u3_syn_4  ;
	output \g238811/u3_syn_4  ;
	output \g238824/u3_syn_4  ;
	output \g238830/u3_syn_4  ;
	output \g238841/u3_syn_4  ;
	output \g238843/u3_syn_4  ;
	output \g238855/u3_syn_4  ;
	output \g238859/u3_syn_4  ;
	output \g238863/u3_syn_4  ;
	output \g238868/u3_syn_4  ;
	output \g238880/u3_syn_4  ;
	output \g238888/u3_syn_4  ;
	output \g238892/u3_syn_4  ;
	output \g238903/u3_syn_4  ;
	output \g238911/u3_syn_4  ;
	output \g238915/u3_syn_4  ;
	output \g238927/u3_syn_4  ;
	output \g238937/u3_syn_4  ;
	output \g238945/u3_syn_4  ;
	output \g238953/u3_syn_4  ;
	output \g238961/u3_syn_4  ;
	output \g238970/u3_syn_4  ;
	output \g238971/u3_syn_4  ;
	output \g238983/u3_syn_4  ;
	output \g238994/u3_syn_4  ;
	output \g239002/u3_syn_4  ;
	output \g239009/u3_syn_4  ;
	output \g239015/u3_syn_4  ;
	output \g239025/u3_syn_4  ;
	output \g239030/u3_syn_4  ;
	output \g239041/u3_syn_4  ;
	output \g239048/u3_syn_4  ;
	output \g239053/u3_syn_4  ;
	output \g239065/u3_syn_4  ;
	output \g239073/u3_syn_4  ;
	output \g239081/u3_syn_4  ;
	output \g239082/u3_syn_4  ;
	output \g239093/u3_syn_4  ;
	output \g239105/u3_syn_4  ;
	output \g239108/u3_syn_4  ;
	output \g239117/u3_syn_4  ;
	output \g239129/u3_syn_4  ;
	output \g239137/u3_syn_4  ;
	output \g239139/u3_syn_4  ;
	output \g239148/u3_syn_4  ;
	output \g239160/u3_syn_4  ;
	output \g239162/u3_syn_4  ;
	output \g239172/u3_syn_4  ;
	output \g239184/u3_syn_4  ;
	output \g239187/u3_syn_4  ;
	output \g239189/u3_syn_4  ;
	output \g239201/u3_syn_4  ;
	output \g239208/u3_syn_4  ;
	output \g239217/u3_syn_4  ;
	output \g239219/u3_syn_4  ;
	output \g239226/u3_syn_4  ;
	output \g239234/u3_syn_4  ;
	output \g239242/u3_syn_4  ;
	output \g239246/u3_syn_4  ;
	output \g239257/u3_syn_4  ;
	output \g239258/u3_syn_4  ;
	output \g239263/u3_syn_4  ;
	output \g239275/u3_syn_4  ;
	output \g239277/u3_syn_4  ;
	output \g239291/u3_syn_4  ;
	output \g239296/u3_syn_4  ;
	output \g239308/u3_syn_4  ;
	output \g239311/u3_syn_4  ;
	output \g239322/u3_syn_4  ;
	output \g239329/u3_syn_4  ;
	output \g239338/u3_syn_4  ;
	output \g239339/u3_syn_4  ;
	output \g239346/u3_syn_4  ;
	output \g239351/u3_syn_4  ;
	output \g239363/u3_syn_4  ;
	output \g239370/u3_syn_4  ;
	output \g239375/u3_syn_4  ;
	output \g239387/u3_syn_4  ;
	output \g239395/u3_syn_4  ;
	output \g239418/u3_syn_4  ;
	output \g239439/u3_syn_4  ;
	output \g239442/u3_syn_4  ;
	output \g239454/u3_syn_4  ;
	output \g239464/u3_syn_4  ;
	output \g239470/u3_syn_4  ;
	output \g239481/u3_syn_4  ;
	output \g239487/u3_syn_4  ;
	output \g239497/u3_syn_4  ;
	output \g239520/u3_syn_4  ;
	output \g239532/u3_syn_4  ;
	output \g239543/u3_syn_4  ;
	output \g239551/u3_syn_4  ;
	output \g239552/u3_syn_4  ;
	output \g239567/u3_syn_4  ;
	output \g239575/u3_syn_4  ;
	output \g239579/u3_syn_4  ;
	output \g239592/u3_syn_4  ;
	output \g239594/u3_syn_4  ;
	output \g239608/u3_syn_4  ;
	output \g239626/u3_syn_4  ;
	output \g239634/u3_syn_4  ;
	output \g239646/u3_syn_4  ;
	output \g239649/u3_syn_4  ;
	output \g239657/u3_syn_4  ;
	output \g239670/u3_syn_4  ;
	output \g239673/u3_syn_4  ;
	output \g239686/u3_syn_4  ;
	output \g239694/u3_syn_4  ;
	output \g239695/u3_syn_4  ;
	output \g239701/u3_syn_4  ;
	output \g239705/u3_syn_4  ;
	output \g239709/u3_syn_4  ;
	output \g239715/u3_syn_4  ;
	output \g239717/u3_syn_4  ;
	output \g239726/u3_syn_4  ;
	output \g239734/u3_syn_4  ;
	output \g239735/u3_syn_4  ;
	output \g239743/u3_syn_4  ;
	output \g239760/u3_syn_4  ;
	output \g239768/u3_syn_4  ;
	output \g239776/u3_syn_4  ;
	output \g239784/u3_syn_4  ;
	output \g239793/u3_syn_4  ;
	output \g239801/u3_syn_4  ;
	output \g239817/u3_syn_4  ;
	output \g239818/u3_syn_4  ;
	output \g239848/u3_syn_4  ;
	output \g239856/u3_syn_4  ;
	output \g239872/u3_syn_4  ;
	output \g239880/u3_syn_4  ;
	output \g239888/u3_syn_4  ;
	output \g239896/u3_syn_4  ;
	output \g239904/u3_syn_4  ;
	output \g239912/u3_syn_4  ;
	output \g239920/u3_syn_4  ;
	output \g239928/u3_syn_4  ;
	output \g239936/u3_syn_4  ;
	output \g239951/u3_syn_4  ;
	output \g239963/u3_syn_4  ;
	output \g239979/u3_syn_4  ;
	output \g239986/u3_syn_4  ;
	output \g239999/u3_syn_4  ;
	output \g240000/u3_syn_4  ;
	output \g240008/u3_syn_4  ;
	output \g240012/u3_syn_4  ;
	output \g240018/u3_syn_4  ;
	output \g240026/u3_syn_4  ;
	output \g240034/u3_syn_4  ;
	output \g240042/u3_syn_4  ;
	output \g240050/u3_syn_4  ;
	output \g240074/u3_syn_4  ;
	output \g240091/u3_syn_4  ;
	output \g240122/u3_syn_4  ;
	output \g240147/u3_syn_4  ;
	output \g240209/u3_syn_4  ;
	output \g240219/u3_syn_4  ;
	output \g240259/u3_syn_4  ;
	output \g240334/u3_syn_4  ;
	output \g240406/u3_syn_4  ;
	output \g240416/u3_syn_4  ;
	output \g240424/u3_syn_4  ;
	output \g240432/u3_syn_4  ;
	output \g240440/u3_syn_4  ;
	output \g240448/u3_syn_4  ;
	output \g240456/u3_syn_4  ;
	output \g240464/u3_syn_4  ;
	output \g240472/u3_syn_4  ;
	output \g240480/u3_syn_4  ;
	output \g240488/u3_syn_4  ;
	output \g240496/u3_syn_4  ;
	output \g240504/u3_syn_4  ;
	output \g240512/u3_syn_4  ;
	output \g240520/u3_syn_4  ;
	output \g240530/u3_syn_4  ;
	output \g240538/u3_syn_4  ;
	output \g240547/u3_syn_4  ;
	output \g240555/u3_syn_4  ;
	output \g240563/u3_syn_4  ;
	output \g240571/u3_syn_4  ;
	output \g240579/u3_syn_4  ;
	output \g240587/u3_syn_4  ;
	output \g240595/u3_syn_4  ;
	output \g240603/u3_syn_4  ;
	output \g240611/u3_syn_4  ;
	output \g240619/u3_syn_4  ;
	output \g240627/u3_syn_4  ;
	output \g240635/u3_syn_4  ;
	output \g240643/u3_syn_4  ;
	output \g240651/u3_syn_4  ;
	output \g240659/u3_syn_4  ;
	output \g240667/u3_syn_4  ;
	output \g240675/u3_syn_4  ;
	output \g240683/u3_syn_4  ;
	output \g240691/u3_syn_4  ;
	output \g240699/u3_syn_4  ;
	output \g240707/u3_syn_4  ;
	output \g240715/u3_syn_4  ;
	output \g240723/u3_syn_4  ;
	output \g240731/u3_syn_4  ;
	output \g240739/u3_syn_4  ;
	output \g240747/u3_syn_4  ;
	output \g240755/u3_syn_4  ;
	output \g240763/u3_syn_4  ;
	output \g240771/u3_syn_4  ;
	output \g240779/u3_syn_4  ;
	output \g240787/u3_syn_4  ;
	output \g240795/u3_syn_4  ;
	output \g240803/u3_syn_4  ;
	output \g240811/u3_syn_4  ;
	output \g240819/u3_syn_4  ;
	output \g240827/u3_syn_4  ;
	output \g240835/u3_syn_4  ;
	output \g240843/u3_syn_4  ;
	output \g240851/u3_syn_4  ;
	output \g240859/u3_syn_4  ;
	output \g240867/u3_syn_4  ;
	output \g240875/u3_syn_4  ;
	output \g240883/u3_syn_4  ;
	output \g240891/u3_syn_4  ;
	output \g240899/u3_syn_4  ;
	output \g240907/u3_syn_4  ;
	output \g240915/u3_syn_4  ;
	output \g240923/u3_syn_4  ;
	output \g240931/u3_syn_4  ;
	output \g240939/u3_syn_4  ;
	output \g240947/u3_syn_4  ;
	output \g240955/u3_syn_4  ;
	output \g240963/u3_syn_4  ;
	output \g240971/u3_syn_4  ;
	output \g240979/u3_syn_4  ;
	output \g240987/u3_syn_4  ;
	output \g240995/u3_syn_4  ;
	output \g241003/u3_syn_4  ;
	output \g241011/u3_syn_4  ;
	output \g241019/u3_syn_4  ;
	output \g241027/u3_syn_4  ;
	output \g241036/u3_syn_4  ;
	output \g241044/u3_syn_4  ;
	output \g241052/u3_syn_4  ;
	output \g241060/u3_syn_4  ;
	output \g241068/u3_syn_4  ;
	output \g241076/u3_syn_4  ;
	output \g241084/u3_syn_4  ;
	output \g241092/u3_syn_4  ;
	output \g241100/u3_syn_4  ;
	output \g241108/u3_syn_4  ;
	output \g241116/u3_syn_4  ;
	output \g241124/u3_syn_4  ;
	output \g241132/u3_syn_4  ;
	output \g241140/u3_syn_4  ;
	output \g241148/u3_syn_4  ;
	output \g241156/u3_syn_4  ;
	output \g241164/u3_syn_4  ;
	output \g241172/u3_syn_4  ;
	output \g241180/u3_syn_4  ;
	output \g241188/u3_syn_4  ;
	output \g241196/u3_syn_4  ;
	output \g241205/u3_syn_4  ;
	output \g241213/u3_syn_4  ;
	output \g241221/u3_syn_4  ;
	output \g241229/u3_syn_4  ;
	output \g241237/u3_syn_4  ;
	output \g241245/u3_syn_4  ;
	output \g241253/u3_syn_4  ;
	output \g241261/u3_syn_4  ;
	output \g241269/u3_syn_4  ;
	output \g241277/u3_syn_4  ;
	output \g241285/u3_syn_4  ;
	output \g241293/u3_syn_4  ;
	output \g241301/u3_syn_4  ;
	output \g241309/u3_syn_4  ;
	output \g241317/u3_syn_4  ;
	output \g241325/u3_syn_4  ;
	output \g241333/u3_syn_4  ;
	output \g241341/u3_syn_4  ;
	output \g241349/u3_syn_4  ;
	output \g241358/u3_syn_4  ;
	output \g241366/u3_syn_4  ;
	output \g241374/u3_syn_4  ;
	output \g241382/u3_syn_4  ;
	output \g241390/u3_syn_4  ;
	output \g241398/u3_syn_4  ;
	output \g241406/u3_syn_4  ;
	output \g241415/u3_syn_4  ;
	output \g241424/u3_syn_4  ;
	output \g241433/u3_syn_4  ;
	output \g241441/u3_syn_4  ;
	output \g241449/u3_syn_4  ;
	output \g241459/u3_syn_4  ;
	output \g241470/u3_syn_4  ;
	output \g241480/u3_syn_4  ;
	output \g241489/u3_syn_4  ;
	output \g241497/u3_syn_4  ;
	output \g241505/u3_syn_4  ;
	output \g241513/u3_syn_4  ;
	output \g241545/_3_  ;
	output \g241580/_00_  ;
	output \g241737/_0_  ;
	output \g241752/_0_  ;
	output \g241755/_0_  ;
	output \g241767/_2__syn_2  ;
	output \g241781/_1__syn_2  ;
	output \g241782/_0_  ;
	output \g241803/_1__syn_2  ;
	output \g241805/_0_  ;
	output \g241812/_1__syn_2  ;
	output \g241814/_1__syn_2  ;
	output \g241816/_1__syn_2  ;
	output \g241819/_1__syn_2  ;
	output \g241822/_1__syn_2  ;
	output \g241823/_0_  ;
	output \g241833/_1__syn_2  ;
	output \g241843/_1__syn_2  ;
	output \g241844/_1__syn_2  ;
	output \g241848/_1__syn_2  ;
	output \g241855/_1__syn_2  ;
	output \g241868/_1__syn_2  ;
	output \g242013/_1__syn_2  ;
	output \g242015/_1__syn_2  ;
	output \g242017/_1__syn_2  ;
	output \g242021/_1__syn_2  ;
	output \g242039/_1__syn_2  ;
	output \g242081/_0_  ;
	output \g242086/_0_  ;
	output \g242101/_3_  ;
	output \g242116/_0_  ;
	output \g242135/_2_  ;
	output \g242147/_0_  ;
	output \g242158/_0_  ;
	output \g242196/_0_  ;
	output \g242202/_0_  ;
	output \g242203/_0_  ;
	output \g242204/_0_  ;
	output \g242212/_0_  ;
	output \g242226/_01_  ;
	output \g242281/_0_  ;
	output \g242407/_0_  ;
	output \g242410/_0_  ;
	output \g242426/_0_  ;
	output \g242438/_2_  ;
	output \g242466/_0_  ;
	output \g242530/_0_  ;
	output \g242532/_0_  ;
	output \g243397/_0_  ;
	output \g245925/_0_  ;
	output \g245932/_0_  ;
	output \g245933/_0_  ;
	output \g245986/_3_  ;
	output \g250157/_3_  ;
	output \g250202/_0_  ;
	output \g250246/_1_  ;
	output \g250248/_0_  ;
	output \g250250/_0_  ;
	output \g250305/_0_  ;
	output \g250323/_0_  ;
	output \g250373/_0_  ;
	output \g250377/_0_  ;
	output \g250412/_0_  ;
	output \g250413/_0_  ;
	output \g250418/_0_  ;
	output \g250419/_0_  ;
	output \g250421/_0_  ;
	output \g250433/_0_  ;
	output \g250448/_3_  ;
	output \g250567/_3_  ;
	output \g258965/_0_  ;
	output \g259006/_0_  ;
	output \g259471/_0_  ;
	output \g259473/_2_  ;
	output \g260557/_0_  ;
	output \g261035/_0_  ;
	output \g261095/_3_  ;
	output \g261207/_2__syn_2  ;
	output \g261754/_0_  ;
	output \g262017/_0_  ;
	output \g262045/_0_  ;
	output \g262046/_0_  ;
	output \g262100/_3_  ;
	output \g263539/_1_  ;
	output \g263574/_0_  ;
	output \g263858/_0_  ;
	output \g264104/_1_  ;
	output \g264107/_1_  ;
	output \g264117/_0_  ;
	output \g264282/_0_  ;
	output \g264511/_0_  ;
	output \g264541/_0_  ;
	output \g264562/_0_  ;
	output \g264618/_0_  ;
	output \g264660/_0_  ;
	output \g264681/_3_  ;
	output \g264727/_0_  ;
	output \g265013/_0_  ;
	output \g265084/_0_  ;
	output \g265378/_0_  ;
	output \g265413/_0_  ;
	output \g265446/_0_  ;
	output \g265486/_0_  ;
	output \g265524/_3_  ;
	output \g265528/_3_  ;
	output \g265548/_3_  ;
	output \g265579/_0_  ;
	output \g265768/_0_  ;
	output \g265801/_0_  ;
	output \g265819/_1_  ;
	output \g265853/_0_  ;
	output \g265933/_0_  ;
	output \g266022/_0_  ;
	output \g266183/_1_  ;
	output \g281909/_0_  ;
	output \g281965/_1_  ;
	output \g282284/_1_  ;
	output \g282639/_1_  ;
	output \g283047/_0_  ;
	output \g283157/_1_  ;
	output \g283184/_0_  ;
	output \g283334/_3_  ;
	output int_o_pad ;
	output \m_wb_adr_o[0]_pad  ;
	output \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  ;
	output \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  ;
	output \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  ;
	wire _w37836_ ;
	wire _w37835_ ;
	wire _w37834_ ;
	wire _w37833_ ;
	wire _w37832_ ;
	wire _w37831_ ;
	wire _w37830_ ;
	wire _w37829_ ;
	wire _w37828_ ;
	wire _w37827_ ;
	wire _w37826_ ;
	wire _w37825_ ;
	wire _w37824_ ;
	wire _w37823_ ;
	wire _w37822_ ;
	wire _w37821_ ;
	wire _w37820_ ;
	wire _w37819_ ;
	wire _w37818_ ;
	wire _w37817_ ;
	wire _w37816_ ;
	wire _w37815_ ;
	wire _w37814_ ;
	wire _w37813_ ;
	wire _w37812_ ;
	wire _w37811_ ;
	wire _w37810_ ;
	wire _w37809_ ;
	wire _w37808_ ;
	wire _w37807_ ;
	wire _w37806_ ;
	wire _w37805_ ;
	wire _w37804_ ;
	wire _w37803_ ;
	wire _w37802_ ;
	wire _w37801_ ;
	wire _w37800_ ;
	wire _w37799_ ;
	wire _w37798_ ;
	wire _w37797_ ;
	wire _w37796_ ;
	wire _w37795_ ;
	wire _w37794_ ;
	wire _w37793_ ;
	wire _w37792_ ;
	wire _w37791_ ;
	wire _w37790_ ;
	wire _w37789_ ;
	wire _w37788_ ;
	wire _w37787_ ;
	wire _w37786_ ;
	wire _w37785_ ;
	wire _w37784_ ;
	wire _w37783_ ;
	wire _w37782_ ;
	wire _w37781_ ;
	wire _w37780_ ;
	wire _w37779_ ;
	wire _w37778_ ;
	wire _w37777_ ;
	wire _w37776_ ;
	wire _w37775_ ;
	wire _w37774_ ;
	wire _w37773_ ;
	wire _w37772_ ;
	wire _w37771_ ;
	wire _w37770_ ;
	wire _w37769_ ;
	wire _w37768_ ;
	wire _w37767_ ;
	wire _w37766_ ;
	wire _w37765_ ;
	wire _w37764_ ;
	wire _w37763_ ;
	wire _w37762_ ;
	wire _w37761_ ;
	wire _w37760_ ;
	wire _w37759_ ;
	wire _w37758_ ;
	wire _w37757_ ;
	wire _w37756_ ;
	wire _w37755_ ;
	wire _w37754_ ;
	wire _w37753_ ;
	wire _w37752_ ;
	wire _w37751_ ;
	wire _w37750_ ;
	wire _w37749_ ;
	wire _w37748_ ;
	wire _w37747_ ;
	wire _w37746_ ;
	wire _w37745_ ;
	wire _w37744_ ;
	wire _w37743_ ;
	wire _w37742_ ;
	wire _w37741_ ;
	wire _w37740_ ;
	wire _w37739_ ;
	wire _w37738_ ;
	wire _w37737_ ;
	wire _w37736_ ;
	wire _w37735_ ;
	wire _w37734_ ;
	wire _w37733_ ;
	wire _w37732_ ;
	wire _w37731_ ;
	wire _w37730_ ;
	wire _w37729_ ;
	wire _w37728_ ;
	wire _w37727_ ;
	wire _w37726_ ;
	wire _w37725_ ;
	wire _w37724_ ;
	wire _w37723_ ;
	wire _w37722_ ;
	wire _w37721_ ;
	wire _w37720_ ;
	wire _w37719_ ;
	wire _w37718_ ;
	wire _w37717_ ;
	wire _w37716_ ;
	wire _w37715_ ;
	wire _w37714_ ;
	wire _w37713_ ;
	wire _w37712_ ;
	wire _w37711_ ;
	wire _w37710_ ;
	wire _w37709_ ;
	wire _w37708_ ;
	wire _w37707_ ;
	wire _w37706_ ;
	wire _w37705_ ;
	wire _w37704_ ;
	wire _w37703_ ;
	wire _w37702_ ;
	wire _w37701_ ;
	wire _w37700_ ;
	wire _w37699_ ;
	wire _w37698_ ;
	wire _w37697_ ;
	wire _w37696_ ;
	wire _w37695_ ;
	wire _w37694_ ;
	wire _w37693_ ;
	wire _w37692_ ;
	wire _w37691_ ;
	wire _w37690_ ;
	wire _w37689_ ;
	wire _w37688_ ;
	wire _w37687_ ;
	wire _w37686_ ;
	wire _w37685_ ;
	wire _w37684_ ;
	wire _w37683_ ;
	wire _w37682_ ;
	wire _w37681_ ;
	wire _w37680_ ;
	wire _w37679_ ;
	wire _w37678_ ;
	wire _w37677_ ;
	wire _w37676_ ;
	wire _w37675_ ;
	wire _w37674_ ;
	wire _w37673_ ;
	wire _w37672_ ;
	wire _w37671_ ;
	wire _w37670_ ;
	wire _w37669_ ;
	wire _w37668_ ;
	wire _w37667_ ;
	wire _w37666_ ;
	wire _w37665_ ;
	wire _w37664_ ;
	wire _w37663_ ;
	wire _w37662_ ;
	wire _w37661_ ;
	wire _w37660_ ;
	wire _w37659_ ;
	wire _w37658_ ;
	wire _w37657_ ;
	wire _w37656_ ;
	wire _w37655_ ;
	wire _w37654_ ;
	wire _w37653_ ;
	wire _w37652_ ;
	wire _w37651_ ;
	wire _w37650_ ;
	wire _w37649_ ;
	wire _w37648_ ;
	wire _w37647_ ;
	wire _w37646_ ;
	wire _w37645_ ;
	wire _w37644_ ;
	wire _w37643_ ;
	wire _w37642_ ;
	wire _w37641_ ;
	wire _w37640_ ;
	wire _w37639_ ;
	wire _w37638_ ;
	wire _w37637_ ;
	wire _w37636_ ;
	wire _w37635_ ;
	wire _w37634_ ;
	wire _w37633_ ;
	wire _w37632_ ;
	wire _w37631_ ;
	wire _w37630_ ;
	wire _w37629_ ;
	wire _w37628_ ;
	wire _w37627_ ;
	wire _w37626_ ;
	wire _w37625_ ;
	wire _w37624_ ;
	wire _w37623_ ;
	wire _w37622_ ;
	wire _w37621_ ;
	wire _w37620_ ;
	wire _w37619_ ;
	wire _w37618_ ;
	wire _w37617_ ;
	wire _w37616_ ;
	wire _w37615_ ;
	wire _w37614_ ;
	wire _w37613_ ;
	wire _w37612_ ;
	wire _w37611_ ;
	wire _w37610_ ;
	wire _w37609_ ;
	wire _w37608_ ;
	wire _w37607_ ;
	wire _w37606_ ;
	wire _w37605_ ;
	wire _w37604_ ;
	wire _w37603_ ;
	wire _w37602_ ;
	wire _w37601_ ;
	wire _w37600_ ;
	wire _w37599_ ;
	wire _w37598_ ;
	wire _w37597_ ;
	wire _w37596_ ;
	wire _w37595_ ;
	wire _w37594_ ;
	wire _w37593_ ;
	wire _w37592_ ;
	wire _w37591_ ;
	wire _w37590_ ;
	wire _w37589_ ;
	wire _w37588_ ;
	wire _w37587_ ;
	wire _w37586_ ;
	wire _w37585_ ;
	wire _w37584_ ;
	wire _w37583_ ;
	wire _w37582_ ;
	wire _w37581_ ;
	wire _w37580_ ;
	wire _w37579_ ;
	wire _w37578_ ;
	wire _w37577_ ;
	wire _w37576_ ;
	wire _w37575_ ;
	wire _w37574_ ;
	wire _w37573_ ;
	wire _w37572_ ;
	wire _w37571_ ;
	wire _w37570_ ;
	wire _w37569_ ;
	wire _w37568_ ;
	wire _w37567_ ;
	wire _w37566_ ;
	wire _w37565_ ;
	wire _w37564_ ;
	wire _w37563_ ;
	wire _w37562_ ;
	wire _w37561_ ;
	wire _w37560_ ;
	wire _w37559_ ;
	wire _w37558_ ;
	wire _w37557_ ;
	wire _w37556_ ;
	wire _w37555_ ;
	wire _w37554_ ;
	wire _w37553_ ;
	wire _w37552_ ;
	wire _w37551_ ;
	wire _w37550_ ;
	wire _w37549_ ;
	wire _w37548_ ;
	wire _w37547_ ;
	wire _w37546_ ;
	wire _w37545_ ;
	wire _w37544_ ;
	wire _w37543_ ;
	wire _w37542_ ;
	wire _w37541_ ;
	wire _w37540_ ;
	wire _w37539_ ;
	wire _w37538_ ;
	wire _w37537_ ;
	wire _w37536_ ;
	wire _w37535_ ;
	wire _w37534_ ;
	wire _w37533_ ;
	wire _w37532_ ;
	wire _w37531_ ;
	wire _w37530_ ;
	wire _w37529_ ;
	wire _w37528_ ;
	wire _w37527_ ;
	wire _w37526_ ;
	wire _w37525_ ;
	wire _w37524_ ;
	wire _w37523_ ;
	wire _w37522_ ;
	wire _w37521_ ;
	wire _w37520_ ;
	wire _w37519_ ;
	wire _w37518_ ;
	wire _w37517_ ;
	wire _w37516_ ;
	wire _w37515_ ;
	wire _w37514_ ;
	wire _w37513_ ;
	wire _w37512_ ;
	wire _w37511_ ;
	wire _w37510_ ;
	wire _w37509_ ;
	wire _w37508_ ;
	wire _w37507_ ;
	wire _w37506_ ;
	wire _w37505_ ;
	wire _w37504_ ;
	wire _w37503_ ;
	wire _w37502_ ;
	wire _w37501_ ;
	wire _w37500_ ;
	wire _w37499_ ;
	wire _w37498_ ;
	wire _w37497_ ;
	wire _w37496_ ;
	wire _w37495_ ;
	wire _w37494_ ;
	wire _w37493_ ;
	wire _w37492_ ;
	wire _w37491_ ;
	wire _w37490_ ;
	wire _w37489_ ;
	wire _w37488_ ;
	wire _w37487_ ;
	wire _w37486_ ;
	wire _w37485_ ;
	wire _w37484_ ;
	wire _w37483_ ;
	wire _w37482_ ;
	wire _w37481_ ;
	wire _w37480_ ;
	wire _w37479_ ;
	wire _w37478_ ;
	wire _w37477_ ;
	wire _w37476_ ;
	wire _w37475_ ;
	wire _w37474_ ;
	wire _w37473_ ;
	wire _w37472_ ;
	wire _w37471_ ;
	wire _w37470_ ;
	wire _w37469_ ;
	wire _w37468_ ;
	wire _w37467_ ;
	wire _w37466_ ;
	wire _w37465_ ;
	wire _w37464_ ;
	wire _w37463_ ;
	wire _w37462_ ;
	wire _w37461_ ;
	wire _w37460_ ;
	wire _w37459_ ;
	wire _w37458_ ;
	wire _w37457_ ;
	wire _w37456_ ;
	wire _w37455_ ;
	wire _w37454_ ;
	wire _w37453_ ;
	wire _w37452_ ;
	wire _w37451_ ;
	wire _w37450_ ;
	wire _w37449_ ;
	wire _w37448_ ;
	wire _w37447_ ;
	wire _w37446_ ;
	wire _w37445_ ;
	wire _w37444_ ;
	wire _w37443_ ;
	wire _w37442_ ;
	wire _w37441_ ;
	wire _w37440_ ;
	wire _w37439_ ;
	wire _w37438_ ;
	wire _w37437_ ;
	wire _w37436_ ;
	wire _w37435_ ;
	wire _w37434_ ;
	wire _w37433_ ;
	wire _w37432_ ;
	wire _w37431_ ;
	wire _w37430_ ;
	wire _w37429_ ;
	wire _w37428_ ;
	wire _w37427_ ;
	wire _w37426_ ;
	wire _w37425_ ;
	wire _w37424_ ;
	wire _w37423_ ;
	wire _w37422_ ;
	wire _w37421_ ;
	wire _w37420_ ;
	wire _w37419_ ;
	wire _w37418_ ;
	wire _w37417_ ;
	wire _w37416_ ;
	wire _w37415_ ;
	wire _w37414_ ;
	wire _w37413_ ;
	wire _w37412_ ;
	wire _w37411_ ;
	wire _w37410_ ;
	wire _w37409_ ;
	wire _w37408_ ;
	wire _w37407_ ;
	wire _w37406_ ;
	wire _w37405_ ;
	wire _w37404_ ;
	wire _w37403_ ;
	wire _w37402_ ;
	wire _w37401_ ;
	wire _w37400_ ;
	wire _w37399_ ;
	wire _w37398_ ;
	wire _w37397_ ;
	wire _w37396_ ;
	wire _w37395_ ;
	wire _w37394_ ;
	wire _w37393_ ;
	wire _w37392_ ;
	wire _w37391_ ;
	wire _w37390_ ;
	wire _w37389_ ;
	wire _w37388_ ;
	wire _w37387_ ;
	wire _w37386_ ;
	wire _w37385_ ;
	wire _w37384_ ;
	wire _w37383_ ;
	wire _w37382_ ;
	wire _w37381_ ;
	wire _w37380_ ;
	wire _w37379_ ;
	wire _w37378_ ;
	wire _w37377_ ;
	wire _w37376_ ;
	wire _w37375_ ;
	wire _w37374_ ;
	wire _w37373_ ;
	wire _w37372_ ;
	wire _w37371_ ;
	wire _w37370_ ;
	wire _w37369_ ;
	wire _w37368_ ;
	wire _w37367_ ;
	wire _w37366_ ;
	wire _w37365_ ;
	wire _w37364_ ;
	wire _w37363_ ;
	wire _w37362_ ;
	wire _w37361_ ;
	wire _w37360_ ;
	wire _w37359_ ;
	wire _w37358_ ;
	wire _w37357_ ;
	wire _w37356_ ;
	wire _w37355_ ;
	wire _w37354_ ;
	wire _w37353_ ;
	wire _w37352_ ;
	wire _w37351_ ;
	wire _w37350_ ;
	wire _w37349_ ;
	wire _w37348_ ;
	wire _w37347_ ;
	wire _w37346_ ;
	wire _w37345_ ;
	wire _w37344_ ;
	wire _w37343_ ;
	wire _w37342_ ;
	wire _w37341_ ;
	wire _w37340_ ;
	wire _w37339_ ;
	wire _w37338_ ;
	wire _w37337_ ;
	wire _w37336_ ;
	wire _w37335_ ;
	wire _w37334_ ;
	wire _w37333_ ;
	wire _w37332_ ;
	wire _w37331_ ;
	wire _w37330_ ;
	wire _w37329_ ;
	wire _w37328_ ;
	wire _w37327_ ;
	wire _w37326_ ;
	wire _w37325_ ;
	wire _w37324_ ;
	wire _w37323_ ;
	wire _w37322_ ;
	wire _w37321_ ;
	wire _w37320_ ;
	wire _w37319_ ;
	wire _w37318_ ;
	wire _w37317_ ;
	wire _w37316_ ;
	wire _w37315_ ;
	wire _w37314_ ;
	wire _w37313_ ;
	wire _w37312_ ;
	wire _w37311_ ;
	wire _w37310_ ;
	wire _w37309_ ;
	wire _w37308_ ;
	wire _w37307_ ;
	wire _w37306_ ;
	wire _w37305_ ;
	wire _w37304_ ;
	wire _w37303_ ;
	wire _w37302_ ;
	wire _w37301_ ;
	wire _w37300_ ;
	wire _w37299_ ;
	wire _w37298_ ;
	wire _w37297_ ;
	wire _w37296_ ;
	wire _w37295_ ;
	wire _w37294_ ;
	wire _w37293_ ;
	wire _w37292_ ;
	wire _w37291_ ;
	wire _w37290_ ;
	wire _w37289_ ;
	wire _w37288_ ;
	wire _w37287_ ;
	wire _w37286_ ;
	wire _w37285_ ;
	wire _w37284_ ;
	wire _w37283_ ;
	wire _w37282_ ;
	wire _w37281_ ;
	wire _w37280_ ;
	wire _w37279_ ;
	wire _w37278_ ;
	wire _w37277_ ;
	wire _w37276_ ;
	wire _w37275_ ;
	wire _w37274_ ;
	wire _w37273_ ;
	wire _w37272_ ;
	wire _w37271_ ;
	wire _w37270_ ;
	wire _w37269_ ;
	wire _w37268_ ;
	wire _w37267_ ;
	wire _w37266_ ;
	wire _w37265_ ;
	wire _w37264_ ;
	wire _w37263_ ;
	wire _w37262_ ;
	wire _w37261_ ;
	wire _w37260_ ;
	wire _w37259_ ;
	wire _w37258_ ;
	wire _w37257_ ;
	wire _w37256_ ;
	wire _w37255_ ;
	wire _w37254_ ;
	wire _w37253_ ;
	wire _w37252_ ;
	wire _w37251_ ;
	wire _w37250_ ;
	wire _w37249_ ;
	wire _w37248_ ;
	wire _w37247_ ;
	wire _w37246_ ;
	wire _w37245_ ;
	wire _w37244_ ;
	wire _w37243_ ;
	wire _w37242_ ;
	wire _w37241_ ;
	wire _w37240_ ;
	wire _w37239_ ;
	wire _w37238_ ;
	wire _w37237_ ;
	wire _w37236_ ;
	wire _w37235_ ;
	wire _w37234_ ;
	wire _w37233_ ;
	wire _w37232_ ;
	wire _w37231_ ;
	wire _w37230_ ;
	wire _w37229_ ;
	wire _w37228_ ;
	wire _w37227_ ;
	wire _w37226_ ;
	wire _w37225_ ;
	wire _w37224_ ;
	wire _w37223_ ;
	wire _w37222_ ;
	wire _w37221_ ;
	wire _w37220_ ;
	wire _w37219_ ;
	wire _w37218_ ;
	wire _w37217_ ;
	wire _w37216_ ;
	wire _w37215_ ;
	wire _w37214_ ;
	wire _w37213_ ;
	wire _w37212_ ;
	wire _w37211_ ;
	wire _w37210_ ;
	wire _w37209_ ;
	wire _w37208_ ;
	wire _w37207_ ;
	wire _w37206_ ;
	wire _w37205_ ;
	wire _w37204_ ;
	wire _w37203_ ;
	wire _w37202_ ;
	wire _w37201_ ;
	wire _w37200_ ;
	wire _w37199_ ;
	wire _w37198_ ;
	wire _w37197_ ;
	wire _w37196_ ;
	wire _w37195_ ;
	wire _w37194_ ;
	wire _w37193_ ;
	wire _w37192_ ;
	wire _w37191_ ;
	wire _w37190_ ;
	wire _w37189_ ;
	wire _w37188_ ;
	wire _w37187_ ;
	wire _w37186_ ;
	wire _w37185_ ;
	wire _w37184_ ;
	wire _w37183_ ;
	wire _w37182_ ;
	wire _w37181_ ;
	wire _w37180_ ;
	wire _w37179_ ;
	wire _w37178_ ;
	wire _w37177_ ;
	wire _w37176_ ;
	wire _w37175_ ;
	wire _w37174_ ;
	wire _w37173_ ;
	wire _w37172_ ;
	wire _w37171_ ;
	wire _w37170_ ;
	wire _w37169_ ;
	wire _w37168_ ;
	wire _w37167_ ;
	wire _w37166_ ;
	wire _w37165_ ;
	wire _w37164_ ;
	wire _w37163_ ;
	wire _w37162_ ;
	wire _w37161_ ;
	wire _w37160_ ;
	wire _w37159_ ;
	wire _w37158_ ;
	wire _w37157_ ;
	wire _w37156_ ;
	wire _w37155_ ;
	wire _w37154_ ;
	wire _w37153_ ;
	wire _w37152_ ;
	wire _w37151_ ;
	wire _w37150_ ;
	wire _w37149_ ;
	wire _w37148_ ;
	wire _w37147_ ;
	wire _w37146_ ;
	wire _w37145_ ;
	wire _w37144_ ;
	wire _w37143_ ;
	wire _w37142_ ;
	wire _w37141_ ;
	wire _w37140_ ;
	wire _w37139_ ;
	wire _w37138_ ;
	wire _w37137_ ;
	wire _w37136_ ;
	wire _w37135_ ;
	wire _w37134_ ;
	wire _w37133_ ;
	wire _w37132_ ;
	wire _w37131_ ;
	wire _w37130_ ;
	wire _w37129_ ;
	wire _w37128_ ;
	wire _w37127_ ;
	wire _w37126_ ;
	wire _w37125_ ;
	wire _w37124_ ;
	wire _w37123_ ;
	wire _w37122_ ;
	wire _w37121_ ;
	wire _w37120_ ;
	wire _w37119_ ;
	wire _w37118_ ;
	wire _w37117_ ;
	wire _w37116_ ;
	wire _w37115_ ;
	wire _w37114_ ;
	wire _w37113_ ;
	wire _w37112_ ;
	wire _w37111_ ;
	wire _w37110_ ;
	wire _w37109_ ;
	wire _w37108_ ;
	wire _w37107_ ;
	wire _w37106_ ;
	wire _w37105_ ;
	wire _w37104_ ;
	wire _w37103_ ;
	wire _w37102_ ;
	wire _w37101_ ;
	wire _w37100_ ;
	wire _w37099_ ;
	wire _w37098_ ;
	wire _w37097_ ;
	wire _w37096_ ;
	wire _w37095_ ;
	wire _w37094_ ;
	wire _w37093_ ;
	wire _w37092_ ;
	wire _w37091_ ;
	wire _w37090_ ;
	wire _w37089_ ;
	wire _w37088_ ;
	wire _w37087_ ;
	wire _w37086_ ;
	wire _w37085_ ;
	wire _w37084_ ;
	wire _w37083_ ;
	wire _w37082_ ;
	wire _w37081_ ;
	wire _w37080_ ;
	wire _w37079_ ;
	wire _w37078_ ;
	wire _w37077_ ;
	wire _w37076_ ;
	wire _w37075_ ;
	wire _w37074_ ;
	wire _w37073_ ;
	wire _w37072_ ;
	wire _w37071_ ;
	wire _w37070_ ;
	wire _w37069_ ;
	wire _w37068_ ;
	wire _w37067_ ;
	wire _w37066_ ;
	wire _w37065_ ;
	wire _w37064_ ;
	wire _w37063_ ;
	wire _w37062_ ;
	wire _w37061_ ;
	wire _w37060_ ;
	wire _w37059_ ;
	wire _w37058_ ;
	wire _w37057_ ;
	wire _w37056_ ;
	wire _w37055_ ;
	wire _w37054_ ;
	wire _w37053_ ;
	wire _w37052_ ;
	wire _w37051_ ;
	wire _w37050_ ;
	wire _w37049_ ;
	wire _w37048_ ;
	wire _w37047_ ;
	wire _w37046_ ;
	wire _w37045_ ;
	wire _w37044_ ;
	wire _w37043_ ;
	wire _w37042_ ;
	wire _w37041_ ;
	wire _w37040_ ;
	wire _w37039_ ;
	wire _w37038_ ;
	wire _w37037_ ;
	wire _w37036_ ;
	wire _w37035_ ;
	wire _w37034_ ;
	wire _w37033_ ;
	wire _w37032_ ;
	wire _w37031_ ;
	wire _w37030_ ;
	wire _w37029_ ;
	wire _w37028_ ;
	wire _w37027_ ;
	wire _w37026_ ;
	wire _w37025_ ;
	wire _w37024_ ;
	wire _w37023_ ;
	wire _w37022_ ;
	wire _w37021_ ;
	wire _w37020_ ;
	wire _w37019_ ;
	wire _w37018_ ;
	wire _w37017_ ;
	wire _w37016_ ;
	wire _w37015_ ;
	wire _w37014_ ;
	wire _w37013_ ;
	wire _w37012_ ;
	wire _w37011_ ;
	wire _w37010_ ;
	wire _w37009_ ;
	wire _w37008_ ;
	wire _w37007_ ;
	wire _w37006_ ;
	wire _w37005_ ;
	wire _w37004_ ;
	wire _w37003_ ;
	wire _w37002_ ;
	wire _w37001_ ;
	wire _w37000_ ;
	wire _w36999_ ;
	wire _w36998_ ;
	wire _w36997_ ;
	wire _w36996_ ;
	wire _w36995_ ;
	wire _w36994_ ;
	wire _w36993_ ;
	wire _w36992_ ;
	wire _w36991_ ;
	wire _w36990_ ;
	wire _w36989_ ;
	wire _w36988_ ;
	wire _w36987_ ;
	wire _w36986_ ;
	wire _w36985_ ;
	wire _w36984_ ;
	wire _w36983_ ;
	wire _w36982_ ;
	wire _w36981_ ;
	wire _w36980_ ;
	wire _w36979_ ;
	wire _w36978_ ;
	wire _w36977_ ;
	wire _w36976_ ;
	wire _w36975_ ;
	wire _w36974_ ;
	wire _w36973_ ;
	wire _w36972_ ;
	wire _w36971_ ;
	wire _w36970_ ;
	wire _w36969_ ;
	wire _w36968_ ;
	wire _w36967_ ;
	wire _w36966_ ;
	wire _w36965_ ;
	wire _w36964_ ;
	wire _w36963_ ;
	wire _w36962_ ;
	wire _w36961_ ;
	wire _w36960_ ;
	wire _w36959_ ;
	wire _w36958_ ;
	wire _w36957_ ;
	wire _w36956_ ;
	wire _w36955_ ;
	wire _w36954_ ;
	wire _w36953_ ;
	wire _w36952_ ;
	wire _w36951_ ;
	wire _w36950_ ;
	wire _w36949_ ;
	wire _w36948_ ;
	wire _w36947_ ;
	wire _w36946_ ;
	wire _w36945_ ;
	wire _w36944_ ;
	wire _w36943_ ;
	wire _w36942_ ;
	wire _w36941_ ;
	wire _w36940_ ;
	wire _w36939_ ;
	wire _w36938_ ;
	wire _w36937_ ;
	wire _w36936_ ;
	wire _w36935_ ;
	wire _w36934_ ;
	wire _w36933_ ;
	wire _w36932_ ;
	wire _w36931_ ;
	wire _w36930_ ;
	wire _w36929_ ;
	wire _w36928_ ;
	wire _w36927_ ;
	wire _w36926_ ;
	wire _w36925_ ;
	wire _w36924_ ;
	wire _w36923_ ;
	wire _w36922_ ;
	wire _w36921_ ;
	wire _w36920_ ;
	wire _w36919_ ;
	wire _w36918_ ;
	wire _w36917_ ;
	wire _w36916_ ;
	wire _w36915_ ;
	wire _w36914_ ;
	wire _w36913_ ;
	wire _w36912_ ;
	wire _w36911_ ;
	wire _w36910_ ;
	wire _w36909_ ;
	wire _w36908_ ;
	wire _w36907_ ;
	wire _w36906_ ;
	wire _w36905_ ;
	wire _w36904_ ;
	wire _w36903_ ;
	wire _w36902_ ;
	wire _w36901_ ;
	wire _w36900_ ;
	wire _w36899_ ;
	wire _w36898_ ;
	wire _w36897_ ;
	wire _w36896_ ;
	wire _w36895_ ;
	wire _w36894_ ;
	wire _w36893_ ;
	wire _w36892_ ;
	wire _w36891_ ;
	wire _w36890_ ;
	wire _w36889_ ;
	wire _w36888_ ;
	wire _w36887_ ;
	wire _w36886_ ;
	wire _w36885_ ;
	wire _w36884_ ;
	wire _w36883_ ;
	wire _w36882_ ;
	wire _w36881_ ;
	wire _w36880_ ;
	wire _w36879_ ;
	wire _w36878_ ;
	wire _w36877_ ;
	wire _w36876_ ;
	wire _w36875_ ;
	wire _w36874_ ;
	wire _w36873_ ;
	wire _w36872_ ;
	wire _w36871_ ;
	wire _w36870_ ;
	wire _w36869_ ;
	wire _w36868_ ;
	wire _w36867_ ;
	wire _w36866_ ;
	wire _w36865_ ;
	wire _w36864_ ;
	wire _w36863_ ;
	wire _w36862_ ;
	wire _w36861_ ;
	wire _w36860_ ;
	wire _w36859_ ;
	wire _w36858_ ;
	wire _w36857_ ;
	wire _w36856_ ;
	wire _w36855_ ;
	wire _w36854_ ;
	wire _w36853_ ;
	wire _w36852_ ;
	wire _w36851_ ;
	wire _w36850_ ;
	wire _w36849_ ;
	wire _w36848_ ;
	wire _w36847_ ;
	wire _w36846_ ;
	wire _w36845_ ;
	wire _w36844_ ;
	wire _w36843_ ;
	wire _w36842_ ;
	wire _w36841_ ;
	wire _w36840_ ;
	wire _w36839_ ;
	wire _w36838_ ;
	wire _w36837_ ;
	wire _w36836_ ;
	wire _w36835_ ;
	wire _w36834_ ;
	wire _w36833_ ;
	wire _w36832_ ;
	wire _w36831_ ;
	wire _w36830_ ;
	wire _w36829_ ;
	wire _w36828_ ;
	wire _w36827_ ;
	wire _w36826_ ;
	wire _w36825_ ;
	wire _w36824_ ;
	wire _w36823_ ;
	wire _w36822_ ;
	wire _w36821_ ;
	wire _w36820_ ;
	wire _w36819_ ;
	wire _w36818_ ;
	wire _w36817_ ;
	wire _w36816_ ;
	wire _w36815_ ;
	wire _w36814_ ;
	wire _w36813_ ;
	wire _w36812_ ;
	wire _w36811_ ;
	wire _w36810_ ;
	wire _w36809_ ;
	wire _w36808_ ;
	wire _w36807_ ;
	wire _w36806_ ;
	wire _w36805_ ;
	wire _w36804_ ;
	wire _w36803_ ;
	wire _w36802_ ;
	wire _w36801_ ;
	wire _w36800_ ;
	wire _w36799_ ;
	wire _w36798_ ;
	wire _w36797_ ;
	wire _w36796_ ;
	wire _w36795_ ;
	wire _w36794_ ;
	wire _w36793_ ;
	wire _w36792_ ;
	wire _w36791_ ;
	wire _w36790_ ;
	wire _w36789_ ;
	wire _w36788_ ;
	wire _w36787_ ;
	wire _w36786_ ;
	wire _w36785_ ;
	wire _w36784_ ;
	wire _w36783_ ;
	wire _w36782_ ;
	wire _w36781_ ;
	wire _w36780_ ;
	wire _w36779_ ;
	wire _w36778_ ;
	wire _w36777_ ;
	wire _w36776_ ;
	wire _w36775_ ;
	wire _w36774_ ;
	wire _w36773_ ;
	wire _w36772_ ;
	wire _w36771_ ;
	wire _w36770_ ;
	wire _w36769_ ;
	wire _w36768_ ;
	wire _w36767_ ;
	wire _w36766_ ;
	wire _w36765_ ;
	wire _w36764_ ;
	wire _w36763_ ;
	wire _w36762_ ;
	wire _w36761_ ;
	wire _w36760_ ;
	wire _w36759_ ;
	wire _w36758_ ;
	wire _w36757_ ;
	wire _w36756_ ;
	wire _w36755_ ;
	wire _w36754_ ;
	wire _w36753_ ;
	wire _w36752_ ;
	wire _w36751_ ;
	wire _w36750_ ;
	wire _w36749_ ;
	wire _w36748_ ;
	wire _w36747_ ;
	wire _w36746_ ;
	wire _w36745_ ;
	wire _w36744_ ;
	wire _w36743_ ;
	wire _w36742_ ;
	wire _w36741_ ;
	wire _w36740_ ;
	wire _w36739_ ;
	wire _w36738_ ;
	wire _w36737_ ;
	wire _w36736_ ;
	wire _w36735_ ;
	wire _w36734_ ;
	wire _w36733_ ;
	wire _w36732_ ;
	wire _w36731_ ;
	wire _w36730_ ;
	wire _w36729_ ;
	wire _w36728_ ;
	wire _w36727_ ;
	wire _w36726_ ;
	wire _w36725_ ;
	wire _w36724_ ;
	wire _w36723_ ;
	wire _w36722_ ;
	wire _w36721_ ;
	wire _w36720_ ;
	wire _w36719_ ;
	wire _w36718_ ;
	wire _w36717_ ;
	wire _w36716_ ;
	wire _w36715_ ;
	wire _w36714_ ;
	wire _w36713_ ;
	wire _w36712_ ;
	wire _w36711_ ;
	wire _w36710_ ;
	wire _w36709_ ;
	wire _w36708_ ;
	wire _w36707_ ;
	wire _w36706_ ;
	wire _w36705_ ;
	wire _w36704_ ;
	wire _w36703_ ;
	wire _w36702_ ;
	wire _w36701_ ;
	wire _w36700_ ;
	wire _w36699_ ;
	wire _w36698_ ;
	wire _w36697_ ;
	wire _w36696_ ;
	wire _w36695_ ;
	wire _w36694_ ;
	wire _w36693_ ;
	wire _w36692_ ;
	wire _w36691_ ;
	wire _w36690_ ;
	wire _w36689_ ;
	wire _w36688_ ;
	wire _w36687_ ;
	wire _w36686_ ;
	wire _w36685_ ;
	wire _w36684_ ;
	wire _w36683_ ;
	wire _w36682_ ;
	wire _w36681_ ;
	wire _w36680_ ;
	wire _w36679_ ;
	wire _w36678_ ;
	wire _w36677_ ;
	wire _w36676_ ;
	wire _w36675_ ;
	wire _w36674_ ;
	wire _w36673_ ;
	wire _w36672_ ;
	wire _w36671_ ;
	wire _w36670_ ;
	wire _w36669_ ;
	wire _w36668_ ;
	wire _w36667_ ;
	wire _w36666_ ;
	wire _w36665_ ;
	wire _w36664_ ;
	wire _w36663_ ;
	wire _w36662_ ;
	wire _w36661_ ;
	wire _w36660_ ;
	wire _w36659_ ;
	wire _w36658_ ;
	wire _w36657_ ;
	wire _w36656_ ;
	wire _w36655_ ;
	wire _w36654_ ;
	wire _w36653_ ;
	wire _w36652_ ;
	wire _w36651_ ;
	wire _w36650_ ;
	wire _w36649_ ;
	wire _w36648_ ;
	wire _w36647_ ;
	wire _w36646_ ;
	wire _w36645_ ;
	wire _w36644_ ;
	wire _w36643_ ;
	wire _w36642_ ;
	wire _w36641_ ;
	wire _w36640_ ;
	wire _w36639_ ;
	wire _w36638_ ;
	wire _w36637_ ;
	wire _w36636_ ;
	wire _w36635_ ;
	wire _w36634_ ;
	wire _w36633_ ;
	wire _w36632_ ;
	wire _w36631_ ;
	wire _w36630_ ;
	wire _w36629_ ;
	wire _w36628_ ;
	wire _w36627_ ;
	wire _w36626_ ;
	wire _w36625_ ;
	wire _w36624_ ;
	wire _w36623_ ;
	wire _w36622_ ;
	wire _w36621_ ;
	wire _w36620_ ;
	wire _w36619_ ;
	wire _w36618_ ;
	wire _w36617_ ;
	wire _w36616_ ;
	wire _w36615_ ;
	wire _w36614_ ;
	wire _w36613_ ;
	wire _w36612_ ;
	wire _w36611_ ;
	wire _w36610_ ;
	wire _w36609_ ;
	wire _w36608_ ;
	wire _w36607_ ;
	wire _w36606_ ;
	wire _w36605_ ;
	wire _w36604_ ;
	wire _w36603_ ;
	wire _w36602_ ;
	wire _w36601_ ;
	wire _w36600_ ;
	wire _w36599_ ;
	wire _w36598_ ;
	wire _w36597_ ;
	wire _w36596_ ;
	wire _w36595_ ;
	wire _w36594_ ;
	wire _w36593_ ;
	wire _w36592_ ;
	wire _w36591_ ;
	wire _w36590_ ;
	wire _w36589_ ;
	wire _w36588_ ;
	wire _w36587_ ;
	wire _w36586_ ;
	wire _w36585_ ;
	wire _w36584_ ;
	wire _w36583_ ;
	wire _w36582_ ;
	wire _w36581_ ;
	wire _w36580_ ;
	wire _w36579_ ;
	wire _w36578_ ;
	wire _w36577_ ;
	wire _w36576_ ;
	wire _w36575_ ;
	wire _w36574_ ;
	wire _w36573_ ;
	wire _w36572_ ;
	wire _w36571_ ;
	wire _w36570_ ;
	wire _w36569_ ;
	wire _w36568_ ;
	wire _w36567_ ;
	wire _w36566_ ;
	wire _w36565_ ;
	wire _w36564_ ;
	wire _w36563_ ;
	wire _w36562_ ;
	wire _w36561_ ;
	wire _w36560_ ;
	wire _w36559_ ;
	wire _w36558_ ;
	wire _w36557_ ;
	wire _w36556_ ;
	wire _w36555_ ;
	wire _w36554_ ;
	wire _w36553_ ;
	wire _w36552_ ;
	wire _w36551_ ;
	wire _w36550_ ;
	wire _w36549_ ;
	wire _w36548_ ;
	wire _w36547_ ;
	wire _w36546_ ;
	wire _w36545_ ;
	wire _w36544_ ;
	wire _w36543_ ;
	wire _w36542_ ;
	wire _w36541_ ;
	wire _w36540_ ;
	wire _w36539_ ;
	wire _w36538_ ;
	wire _w36537_ ;
	wire _w36536_ ;
	wire _w36535_ ;
	wire _w36534_ ;
	wire _w36533_ ;
	wire _w36532_ ;
	wire _w36531_ ;
	wire _w36530_ ;
	wire _w36529_ ;
	wire _w36528_ ;
	wire _w36527_ ;
	wire _w36526_ ;
	wire _w36525_ ;
	wire _w36524_ ;
	wire _w36523_ ;
	wire _w36522_ ;
	wire _w36521_ ;
	wire _w36520_ ;
	wire _w36519_ ;
	wire _w36518_ ;
	wire _w36517_ ;
	wire _w36516_ ;
	wire _w36515_ ;
	wire _w36514_ ;
	wire _w36513_ ;
	wire _w36512_ ;
	wire _w36511_ ;
	wire _w36510_ ;
	wire _w36509_ ;
	wire _w36508_ ;
	wire _w36507_ ;
	wire _w36506_ ;
	wire _w36505_ ;
	wire _w36504_ ;
	wire _w36503_ ;
	wire _w36502_ ;
	wire _w36501_ ;
	wire _w36500_ ;
	wire _w36499_ ;
	wire _w36498_ ;
	wire _w36497_ ;
	wire _w36496_ ;
	wire _w36495_ ;
	wire _w36494_ ;
	wire _w36493_ ;
	wire _w36492_ ;
	wire _w36491_ ;
	wire _w36490_ ;
	wire _w36489_ ;
	wire _w36488_ ;
	wire _w36487_ ;
	wire _w36486_ ;
	wire _w36485_ ;
	wire _w36484_ ;
	wire _w36483_ ;
	wire _w36482_ ;
	wire _w36481_ ;
	wire _w36480_ ;
	wire _w36479_ ;
	wire _w36478_ ;
	wire _w36477_ ;
	wire _w36476_ ;
	wire _w36475_ ;
	wire _w36474_ ;
	wire _w36473_ ;
	wire _w36472_ ;
	wire _w36471_ ;
	wire _w36470_ ;
	wire _w36469_ ;
	wire _w36468_ ;
	wire _w36467_ ;
	wire _w36466_ ;
	wire _w36465_ ;
	wire _w36464_ ;
	wire _w36463_ ;
	wire _w36462_ ;
	wire _w36461_ ;
	wire _w36460_ ;
	wire _w36459_ ;
	wire _w36458_ ;
	wire _w36457_ ;
	wire _w36456_ ;
	wire _w36455_ ;
	wire _w36454_ ;
	wire _w36453_ ;
	wire _w36452_ ;
	wire _w36451_ ;
	wire _w36450_ ;
	wire _w36449_ ;
	wire _w36448_ ;
	wire _w36447_ ;
	wire _w36446_ ;
	wire _w36445_ ;
	wire _w36444_ ;
	wire _w36443_ ;
	wire _w36442_ ;
	wire _w36441_ ;
	wire _w36440_ ;
	wire _w36439_ ;
	wire _w36438_ ;
	wire _w36437_ ;
	wire _w36436_ ;
	wire _w36435_ ;
	wire _w36434_ ;
	wire _w36433_ ;
	wire _w36432_ ;
	wire _w36431_ ;
	wire _w36430_ ;
	wire _w36429_ ;
	wire _w36428_ ;
	wire _w36427_ ;
	wire _w36426_ ;
	wire _w36425_ ;
	wire _w36424_ ;
	wire _w36423_ ;
	wire _w36422_ ;
	wire _w36421_ ;
	wire _w36420_ ;
	wire _w36419_ ;
	wire _w36418_ ;
	wire _w36417_ ;
	wire _w36416_ ;
	wire _w36415_ ;
	wire _w36414_ ;
	wire _w36413_ ;
	wire _w36412_ ;
	wire _w36411_ ;
	wire _w36410_ ;
	wire _w36409_ ;
	wire _w36408_ ;
	wire _w36407_ ;
	wire _w36406_ ;
	wire _w36405_ ;
	wire _w36404_ ;
	wire _w36403_ ;
	wire _w36402_ ;
	wire _w36401_ ;
	wire _w36400_ ;
	wire _w36399_ ;
	wire _w36398_ ;
	wire _w36397_ ;
	wire _w36396_ ;
	wire _w36395_ ;
	wire _w36394_ ;
	wire _w36393_ ;
	wire _w36392_ ;
	wire _w36391_ ;
	wire _w36390_ ;
	wire _w36389_ ;
	wire _w36388_ ;
	wire _w36387_ ;
	wire _w36386_ ;
	wire _w36385_ ;
	wire _w36384_ ;
	wire _w36383_ ;
	wire _w36382_ ;
	wire _w36381_ ;
	wire _w36380_ ;
	wire _w36379_ ;
	wire _w36378_ ;
	wire _w36377_ ;
	wire _w36376_ ;
	wire _w36375_ ;
	wire _w36374_ ;
	wire _w36373_ ;
	wire _w36372_ ;
	wire _w36371_ ;
	wire _w36370_ ;
	wire _w36369_ ;
	wire _w36368_ ;
	wire _w36367_ ;
	wire _w36366_ ;
	wire _w36365_ ;
	wire _w36364_ ;
	wire _w36363_ ;
	wire _w36362_ ;
	wire _w36361_ ;
	wire _w36360_ ;
	wire _w36359_ ;
	wire _w36358_ ;
	wire _w36357_ ;
	wire _w36356_ ;
	wire _w36355_ ;
	wire _w36354_ ;
	wire _w36353_ ;
	wire _w36352_ ;
	wire _w36351_ ;
	wire _w36350_ ;
	wire _w36349_ ;
	wire _w36348_ ;
	wire _w36347_ ;
	wire _w36346_ ;
	wire _w36345_ ;
	wire _w36344_ ;
	wire _w36343_ ;
	wire _w36342_ ;
	wire _w36341_ ;
	wire _w36340_ ;
	wire _w36339_ ;
	wire _w36338_ ;
	wire _w36337_ ;
	wire _w36336_ ;
	wire _w36335_ ;
	wire _w36334_ ;
	wire _w36333_ ;
	wire _w36332_ ;
	wire _w36331_ ;
	wire _w36330_ ;
	wire _w36329_ ;
	wire _w36328_ ;
	wire _w36327_ ;
	wire _w36326_ ;
	wire _w36325_ ;
	wire _w36324_ ;
	wire _w36323_ ;
	wire _w36322_ ;
	wire _w36321_ ;
	wire _w36320_ ;
	wire _w36319_ ;
	wire _w36318_ ;
	wire _w36317_ ;
	wire _w36316_ ;
	wire _w36315_ ;
	wire _w36314_ ;
	wire _w36313_ ;
	wire _w36312_ ;
	wire _w36311_ ;
	wire _w36310_ ;
	wire _w36309_ ;
	wire _w36308_ ;
	wire _w36307_ ;
	wire _w36306_ ;
	wire _w36305_ ;
	wire _w36304_ ;
	wire _w36303_ ;
	wire _w36302_ ;
	wire _w36301_ ;
	wire _w36300_ ;
	wire _w36299_ ;
	wire _w36298_ ;
	wire _w36297_ ;
	wire _w36296_ ;
	wire _w36295_ ;
	wire _w36294_ ;
	wire _w36293_ ;
	wire _w36292_ ;
	wire _w36291_ ;
	wire _w36290_ ;
	wire _w36289_ ;
	wire _w36288_ ;
	wire _w36287_ ;
	wire _w36286_ ;
	wire _w36285_ ;
	wire _w36284_ ;
	wire _w36283_ ;
	wire _w36282_ ;
	wire _w36281_ ;
	wire _w36280_ ;
	wire _w36279_ ;
	wire _w36278_ ;
	wire _w36277_ ;
	wire _w36276_ ;
	wire _w36275_ ;
	wire _w36274_ ;
	wire _w36273_ ;
	wire _w36272_ ;
	wire _w36271_ ;
	wire _w36270_ ;
	wire _w36269_ ;
	wire _w36268_ ;
	wire _w36267_ ;
	wire _w36266_ ;
	wire _w36265_ ;
	wire _w36264_ ;
	wire _w36263_ ;
	wire _w36262_ ;
	wire _w36261_ ;
	wire _w36260_ ;
	wire _w36259_ ;
	wire _w36258_ ;
	wire _w36257_ ;
	wire _w36256_ ;
	wire _w36255_ ;
	wire _w36254_ ;
	wire _w36253_ ;
	wire _w36252_ ;
	wire _w36251_ ;
	wire _w36250_ ;
	wire _w36249_ ;
	wire _w36248_ ;
	wire _w36247_ ;
	wire _w36246_ ;
	wire _w36245_ ;
	wire _w36244_ ;
	wire _w36243_ ;
	wire _w36242_ ;
	wire _w36241_ ;
	wire _w36240_ ;
	wire _w36239_ ;
	wire _w36238_ ;
	wire _w36237_ ;
	wire _w36236_ ;
	wire _w36235_ ;
	wire _w36234_ ;
	wire _w36233_ ;
	wire _w36232_ ;
	wire _w36231_ ;
	wire _w36230_ ;
	wire _w36229_ ;
	wire _w36228_ ;
	wire _w36227_ ;
	wire _w36226_ ;
	wire _w36225_ ;
	wire _w36224_ ;
	wire _w36223_ ;
	wire _w36222_ ;
	wire _w36221_ ;
	wire _w36220_ ;
	wire _w36219_ ;
	wire _w36218_ ;
	wire _w36217_ ;
	wire _w36216_ ;
	wire _w36215_ ;
	wire _w36214_ ;
	wire _w36213_ ;
	wire _w36212_ ;
	wire _w36211_ ;
	wire _w36210_ ;
	wire _w36209_ ;
	wire _w36208_ ;
	wire _w36207_ ;
	wire _w36206_ ;
	wire _w36205_ ;
	wire _w36204_ ;
	wire _w36203_ ;
	wire _w36202_ ;
	wire _w36201_ ;
	wire _w36200_ ;
	wire _w36199_ ;
	wire _w36198_ ;
	wire _w36197_ ;
	wire _w36196_ ;
	wire _w36195_ ;
	wire _w36194_ ;
	wire _w36193_ ;
	wire _w36192_ ;
	wire _w36191_ ;
	wire _w36190_ ;
	wire _w36189_ ;
	wire _w36188_ ;
	wire _w36187_ ;
	wire _w36186_ ;
	wire _w36185_ ;
	wire _w36184_ ;
	wire _w36183_ ;
	wire _w36182_ ;
	wire _w36181_ ;
	wire _w36180_ ;
	wire _w36179_ ;
	wire _w36178_ ;
	wire _w36177_ ;
	wire _w36176_ ;
	wire _w36175_ ;
	wire _w36174_ ;
	wire _w36173_ ;
	wire _w36172_ ;
	wire _w36171_ ;
	wire _w36170_ ;
	wire _w36169_ ;
	wire _w36168_ ;
	wire _w36167_ ;
	wire _w36166_ ;
	wire _w36165_ ;
	wire _w36164_ ;
	wire _w36163_ ;
	wire _w36162_ ;
	wire _w36161_ ;
	wire _w36160_ ;
	wire _w36159_ ;
	wire _w36158_ ;
	wire _w36157_ ;
	wire _w36156_ ;
	wire _w36155_ ;
	wire _w36154_ ;
	wire _w36153_ ;
	wire _w36152_ ;
	wire _w36151_ ;
	wire _w36150_ ;
	wire _w36149_ ;
	wire _w36148_ ;
	wire _w36147_ ;
	wire _w36146_ ;
	wire _w36145_ ;
	wire _w36144_ ;
	wire _w36143_ ;
	wire _w36142_ ;
	wire _w36141_ ;
	wire _w36140_ ;
	wire _w36139_ ;
	wire _w36138_ ;
	wire _w36137_ ;
	wire _w36136_ ;
	wire _w36135_ ;
	wire _w36134_ ;
	wire _w36133_ ;
	wire _w36132_ ;
	wire _w36131_ ;
	wire _w36130_ ;
	wire _w36129_ ;
	wire _w36128_ ;
	wire _w36127_ ;
	wire _w36126_ ;
	wire _w36125_ ;
	wire _w36124_ ;
	wire _w36123_ ;
	wire _w36122_ ;
	wire _w36121_ ;
	wire _w36120_ ;
	wire _w36119_ ;
	wire _w36118_ ;
	wire _w36117_ ;
	wire _w36116_ ;
	wire _w36115_ ;
	wire _w36114_ ;
	wire _w36113_ ;
	wire _w36112_ ;
	wire _w36111_ ;
	wire _w36110_ ;
	wire _w36109_ ;
	wire _w36108_ ;
	wire _w36107_ ;
	wire _w36106_ ;
	wire _w36105_ ;
	wire _w36104_ ;
	wire _w36103_ ;
	wire _w36102_ ;
	wire _w36101_ ;
	wire _w36100_ ;
	wire _w36099_ ;
	wire _w36098_ ;
	wire _w36097_ ;
	wire _w36096_ ;
	wire _w36095_ ;
	wire _w36094_ ;
	wire _w36093_ ;
	wire _w36092_ ;
	wire _w36091_ ;
	wire _w36090_ ;
	wire _w36089_ ;
	wire _w36088_ ;
	wire _w36087_ ;
	wire _w36086_ ;
	wire _w36085_ ;
	wire _w36084_ ;
	wire _w36083_ ;
	wire _w36082_ ;
	wire _w36081_ ;
	wire _w36080_ ;
	wire _w36079_ ;
	wire _w36078_ ;
	wire _w36077_ ;
	wire _w36076_ ;
	wire _w36075_ ;
	wire _w36074_ ;
	wire _w36073_ ;
	wire _w36072_ ;
	wire _w36071_ ;
	wire _w36070_ ;
	wire _w36069_ ;
	wire _w36068_ ;
	wire _w36067_ ;
	wire _w36066_ ;
	wire _w36065_ ;
	wire _w36064_ ;
	wire _w36063_ ;
	wire _w36062_ ;
	wire _w36061_ ;
	wire _w36060_ ;
	wire _w36059_ ;
	wire _w36058_ ;
	wire _w36057_ ;
	wire _w36056_ ;
	wire _w36055_ ;
	wire _w36054_ ;
	wire _w36053_ ;
	wire _w36052_ ;
	wire _w36051_ ;
	wire _w36050_ ;
	wire _w36049_ ;
	wire _w36048_ ;
	wire _w36047_ ;
	wire _w36046_ ;
	wire _w36045_ ;
	wire _w36044_ ;
	wire _w36043_ ;
	wire _w36042_ ;
	wire _w36041_ ;
	wire _w36040_ ;
	wire _w36039_ ;
	wire _w36038_ ;
	wire _w36037_ ;
	wire _w36036_ ;
	wire _w36035_ ;
	wire _w36034_ ;
	wire _w36033_ ;
	wire _w36032_ ;
	wire _w36031_ ;
	wire _w36030_ ;
	wire _w36029_ ;
	wire _w36028_ ;
	wire _w36027_ ;
	wire _w36026_ ;
	wire _w36025_ ;
	wire _w36024_ ;
	wire _w36023_ ;
	wire _w36022_ ;
	wire _w36021_ ;
	wire _w36020_ ;
	wire _w36019_ ;
	wire _w36018_ ;
	wire _w36017_ ;
	wire _w36016_ ;
	wire _w36015_ ;
	wire _w36014_ ;
	wire _w36013_ ;
	wire _w36012_ ;
	wire _w36011_ ;
	wire _w36010_ ;
	wire _w36009_ ;
	wire _w36008_ ;
	wire _w36007_ ;
	wire _w36006_ ;
	wire _w36005_ ;
	wire _w36004_ ;
	wire _w36003_ ;
	wire _w36002_ ;
	wire _w36001_ ;
	wire _w36000_ ;
	wire _w35999_ ;
	wire _w35998_ ;
	wire _w35997_ ;
	wire _w35996_ ;
	wire _w35995_ ;
	wire _w35994_ ;
	wire _w35993_ ;
	wire _w35992_ ;
	wire _w35991_ ;
	wire _w35990_ ;
	wire _w35989_ ;
	wire _w35988_ ;
	wire _w35987_ ;
	wire _w35986_ ;
	wire _w35985_ ;
	wire _w35984_ ;
	wire _w35983_ ;
	wire _w35982_ ;
	wire _w35981_ ;
	wire _w35980_ ;
	wire _w35979_ ;
	wire _w35978_ ;
	wire _w35977_ ;
	wire _w35976_ ;
	wire _w35975_ ;
	wire _w35974_ ;
	wire _w35973_ ;
	wire _w35972_ ;
	wire _w35971_ ;
	wire _w35970_ ;
	wire _w35969_ ;
	wire _w35968_ ;
	wire _w35967_ ;
	wire _w35966_ ;
	wire _w35965_ ;
	wire _w35964_ ;
	wire _w35963_ ;
	wire _w35962_ ;
	wire _w35961_ ;
	wire _w35960_ ;
	wire _w35959_ ;
	wire _w35958_ ;
	wire _w35957_ ;
	wire _w35956_ ;
	wire _w35955_ ;
	wire _w35954_ ;
	wire _w35953_ ;
	wire _w35952_ ;
	wire _w35951_ ;
	wire _w35950_ ;
	wire _w35949_ ;
	wire _w35948_ ;
	wire _w35947_ ;
	wire _w35946_ ;
	wire _w35945_ ;
	wire _w35944_ ;
	wire _w35943_ ;
	wire _w35942_ ;
	wire _w35941_ ;
	wire _w35940_ ;
	wire _w35939_ ;
	wire _w35938_ ;
	wire _w35937_ ;
	wire _w35936_ ;
	wire _w35935_ ;
	wire _w35934_ ;
	wire _w35933_ ;
	wire _w35932_ ;
	wire _w35931_ ;
	wire _w35930_ ;
	wire _w35929_ ;
	wire _w35928_ ;
	wire _w35927_ ;
	wire _w35926_ ;
	wire _w35925_ ;
	wire _w35924_ ;
	wire _w35923_ ;
	wire _w35922_ ;
	wire _w35921_ ;
	wire _w35920_ ;
	wire _w35919_ ;
	wire _w35918_ ;
	wire _w35917_ ;
	wire _w35916_ ;
	wire _w35915_ ;
	wire _w35914_ ;
	wire _w35913_ ;
	wire _w35912_ ;
	wire _w35911_ ;
	wire _w35910_ ;
	wire _w35909_ ;
	wire _w35908_ ;
	wire _w35907_ ;
	wire _w35906_ ;
	wire _w35905_ ;
	wire _w35904_ ;
	wire _w35903_ ;
	wire _w35902_ ;
	wire _w35901_ ;
	wire _w35900_ ;
	wire _w35899_ ;
	wire _w35898_ ;
	wire _w35897_ ;
	wire _w35896_ ;
	wire _w35895_ ;
	wire _w35894_ ;
	wire _w35893_ ;
	wire _w35892_ ;
	wire _w35891_ ;
	wire _w35890_ ;
	wire _w35889_ ;
	wire _w35888_ ;
	wire _w35887_ ;
	wire _w35886_ ;
	wire _w35885_ ;
	wire _w35884_ ;
	wire _w35883_ ;
	wire _w35882_ ;
	wire _w35881_ ;
	wire _w35880_ ;
	wire _w35879_ ;
	wire _w35878_ ;
	wire _w35877_ ;
	wire _w35876_ ;
	wire _w35875_ ;
	wire _w35874_ ;
	wire _w35873_ ;
	wire _w35872_ ;
	wire _w35871_ ;
	wire _w35870_ ;
	wire _w35869_ ;
	wire _w35868_ ;
	wire _w35867_ ;
	wire _w35866_ ;
	wire _w35865_ ;
	wire _w35864_ ;
	wire _w35863_ ;
	wire _w35862_ ;
	wire _w35861_ ;
	wire _w35860_ ;
	wire _w35859_ ;
	wire _w35858_ ;
	wire _w35857_ ;
	wire _w35856_ ;
	wire _w35855_ ;
	wire _w35854_ ;
	wire _w35853_ ;
	wire _w35852_ ;
	wire _w35851_ ;
	wire _w35850_ ;
	wire _w35849_ ;
	wire _w35848_ ;
	wire _w35847_ ;
	wire _w35846_ ;
	wire _w35845_ ;
	wire _w35844_ ;
	wire _w35843_ ;
	wire _w35842_ ;
	wire _w35841_ ;
	wire _w35840_ ;
	wire _w35839_ ;
	wire _w35838_ ;
	wire _w35837_ ;
	wire _w35836_ ;
	wire _w35835_ ;
	wire _w35834_ ;
	wire _w35833_ ;
	wire _w35832_ ;
	wire _w35831_ ;
	wire _w35830_ ;
	wire _w35829_ ;
	wire _w35828_ ;
	wire _w35827_ ;
	wire _w35826_ ;
	wire _w35825_ ;
	wire _w35824_ ;
	wire _w35823_ ;
	wire _w35822_ ;
	wire _w35821_ ;
	wire _w35820_ ;
	wire _w35819_ ;
	wire _w35818_ ;
	wire _w35817_ ;
	wire _w35816_ ;
	wire _w35815_ ;
	wire _w35814_ ;
	wire _w35813_ ;
	wire _w35812_ ;
	wire _w35811_ ;
	wire _w35810_ ;
	wire _w35809_ ;
	wire _w35808_ ;
	wire _w35807_ ;
	wire _w35806_ ;
	wire _w35805_ ;
	wire _w35804_ ;
	wire _w35803_ ;
	wire _w35802_ ;
	wire _w35801_ ;
	wire _w35800_ ;
	wire _w35799_ ;
	wire _w35798_ ;
	wire _w35797_ ;
	wire _w35796_ ;
	wire _w35795_ ;
	wire _w35794_ ;
	wire _w35793_ ;
	wire _w35792_ ;
	wire _w35791_ ;
	wire _w35790_ ;
	wire _w35789_ ;
	wire _w35788_ ;
	wire _w35787_ ;
	wire _w35786_ ;
	wire _w35785_ ;
	wire _w35784_ ;
	wire _w35783_ ;
	wire _w35782_ ;
	wire _w35781_ ;
	wire _w35780_ ;
	wire _w35779_ ;
	wire _w35778_ ;
	wire _w35777_ ;
	wire _w35776_ ;
	wire _w35775_ ;
	wire _w35774_ ;
	wire _w35773_ ;
	wire _w35772_ ;
	wire _w35771_ ;
	wire _w35770_ ;
	wire _w35769_ ;
	wire _w35768_ ;
	wire _w35767_ ;
	wire _w35766_ ;
	wire _w35765_ ;
	wire _w35764_ ;
	wire _w35763_ ;
	wire _w35762_ ;
	wire _w35761_ ;
	wire _w35760_ ;
	wire _w35759_ ;
	wire _w35758_ ;
	wire _w35757_ ;
	wire _w35756_ ;
	wire _w35755_ ;
	wire _w35754_ ;
	wire _w35753_ ;
	wire _w35752_ ;
	wire _w35751_ ;
	wire _w35750_ ;
	wire _w35749_ ;
	wire _w35748_ ;
	wire _w35747_ ;
	wire _w35746_ ;
	wire _w35745_ ;
	wire _w35744_ ;
	wire _w35743_ ;
	wire _w35742_ ;
	wire _w35741_ ;
	wire _w35740_ ;
	wire _w35739_ ;
	wire _w35738_ ;
	wire _w35737_ ;
	wire _w35736_ ;
	wire _w35735_ ;
	wire _w35734_ ;
	wire _w35733_ ;
	wire _w35732_ ;
	wire _w35731_ ;
	wire _w35730_ ;
	wire _w35729_ ;
	wire _w35728_ ;
	wire _w35727_ ;
	wire _w35726_ ;
	wire _w35725_ ;
	wire _w35724_ ;
	wire _w35723_ ;
	wire _w35722_ ;
	wire _w35721_ ;
	wire _w35720_ ;
	wire _w35719_ ;
	wire _w35718_ ;
	wire _w35717_ ;
	wire _w35716_ ;
	wire _w35715_ ;
	wire _w35714_ ;
	wire _w35713_ ;
	wire _w35712_ ;
	wire _w35711_ ;
	wire _w35710_ ;
	wire _w35709_ ;
	wire _w35708_ ;
	wire _w35707_ ;
	wire _w35706_ ;
	wire _w35705_ ;
	wire _w35704_ ;
	wire _w35703_ ;
	wire _w35702_ ;
	wire _w35701_ ;
	wire _w35700_ ;
	wire _w35699_ ;
	wire _w35698_ ;
	wire _w35697_ ;
	wire _w35696_ ;
	wire _w35695_ ;
	wire _w35694_ ;
	wire _w35693_ ;
	wire _w35692_ ;
	wire _w35691_ ;
	wire _w35690_ ;
	wire _w35689_ ;
	wire _w35688_ ;
	wire _w35687_ ;
	wire _w35686_ ;
	wire _w35685_ ;
	wire _w35684_ ;
	wire _w35683_ ;
	wire _w35682_ ;
	wire _w35681_ ;
	wire _w35680_ ;
	wire _w35679_ ;
	wire _w35678_ ;
	wire _w35677_ ;
	wire _w35676_ ;
	wire _w35675_ ;
	wire _w35674_ ;
	wire _w35673_ ;
	wire _w35672_ ;
	wire _w35671_ ;
	wire _w35670_ ;
	wire _w35669_ ;
	wire _w35668_ ;
	wire _w35667_ ;
	wire _w35666_ ;
	wire _w35665_ ;
	wire _w35664_ ;
	wire _w35663_ ;
	wire _w35662_ ;
	wire _w35661_ ;
	wire _w35660_ ;
	wire _w35659_ ;
	wire _w35658_ ;
	wire _w35657_ ;
	wire _w35656_ ;
	wire _w35655_ ;
	wire _w35654_ ;
	wire _w35653_ ;
	wire _w35652_ ;
	wire _w35651_ ;
	wire _w35650_ ;
	wire _w35649_ ;
	wire _w35648_ ;
	wire _w35647_ ;
	wire _w35646_ ;
	wire _w35645_ ;
	wire _w35644_ ;
	wire _w35643_ ;
	wire _w35642_ ;
	wire _w35641_ ;
	wire _w35640_ ;
	wire _w35639_ ;
	wire _w35638_ ;
	wire _w35637_ ;
	wire _w35636_ ;
	wire _w35635_ ;
	wire _w35634_ ;
	wire _w35633_ ;
	wire _w35632_ ;
	wire _w35631_ ;
	wire _w35630_ ;
	wire _w35629_ ;
	wire _w35628_ ;
	wire _w35627_ ;
	wire _w35626_ ;
	wire _w35625_ ;
	wire _w35624_ ;
	wire _w35623_ ;
	wire _w35622_ ;
	wire _w35621_ ;
	wire _w35620_ ;
	wire _w35619_ ;
	wire _w35618_ ;
	wire _w35617_ ;
	wire _w35616_ ;
	wire _w35615_ ;
	wire _w35614_ ;
	wire _w35613_ ;
	wire _w35612_ ;
	wire _w35611_ ;
	wire _w35610_ ;
	wire _w35609_ ;
	wire _w35608_ ;
	wire _w35607_ ;
	wire _w35606_ ;
	wire _w35605_ ;
	wire _w35604_ ;
	wire _w35603_ ;
	wire _w35602_ ;
	wire _w35601_ ;
	wire _w35600_ ;
	wire _w35599_ ;
	wire _w35598_ ;
	wire _w35597_ ;
	wire _w35596_ ;
	wire _w35595_ ;
	wire _w35594_ ;
	wire _w35593_ ;
	wire _w35592_ ;
	wire _w35591_ ;
	wire _w35590_ ;
	wire _w35589_ ;
	wire _w35588_ ;
	wire _w35587_ ;
	wire _w35586_ ;
	wire _w35585_ ;
	wire _w35584_ ;
	wire _w35583_ ;
	wire _w35582_ ;
	wire _w35581_ ;
	wire _w35580_ ;
	wire _w35579_ ;
	wire _w35578_ ;
	wire _w35577_ ;
	wire _w35576_ ;
	wire _w35575_ ;
	wire _w35574_ ;
	wire _w35573_ ;
	wire _w35572_ ;
	wire _w35571_ ;
	wire _w35570_ ;
	wire _w35569_ ;
	wire _w35568_ ;
	wire _w35567_ ;
	wire _w35566_ ;
	wire _w35565_ ;
	wire _w35564_ ;
	wire _w35563_ ;
	wire _w35562_ ;
	wire _w35561_ ;
	wire _w35560_ ;
	wire _w35559_ ;
	wire _w35558_ ;
	wire _w35557_ ;
	wire _w35556_ ;
	wire _w35555_ ;
	wire _w35554_ ;
	wire _w35553_ ;
	wire _w35552_ ;
	wire _w35551_ ;
	wire _w35550_ ;
	wire _w35549_ ;
	wire _w35548_ ;
	wire _w35547_ ;
	wire _w35546_ ;
	wire _w35545_ ;
	wire _w35544_ ;
	wire _w35543_ ;
	wire _w35542_ ;
	wire _w35541_ ;
	wire _w35540_ ;
	wire _w35539_ ;
	wire _w35538_ ;
	wire _w35537_ ;
	wire _w35536_ ;
	wire _w35535_ ;
	wire _w35534_ ;
	wire _w35533_ ;
	wire _w35532_ ;
	wire _w35531_ ;
	wire _w35530_ ;
	wire _w35529_ ;
	wire _w35528_ ;
	wire _w35527_ ;
	wire _w35526_ ;
	wire _w35525_ ;
	wire _w35524_ ;
	wire _w35523_ ;
	wire _w35522_ ;
	wire _w35521_ ;
	wire _w35520_ ;
	wire _w35519_ ;
	wire _w35518_ ;
	wire _w35517_ ;
	wire _w35516_ ;
	wire _w35515_ ;
	wire _w35514_ ;
	wire _w35513_ ;
	wire _w35512_ ;
	wire _w35511_ ;
	wire _w35510_ ;
	wire _w35509_ ;
	wire _w35508_ ;
	wire _w35507_ ;
	wire _w35506_ ;
	wire _w35505_ ;
	wire _w35504_ ;
	wire _w35503_ ;
	wire _w35502_ ;
	wire _w35501_ ;
	wire _w35500_ ;
	wire _w35499_ ;
	wire _w35498_ ;
	wire _w35497_ ;
	wire _w35496_ ;
	wire _w35495_ ;
	wire _w35494_ ;
	wire _w35493_ ;
	wire _w35492_ ;
	wire _w35491_ ;
	wire _w35490_ ;
	wire _w35489_ ;
	wire _w35488_ ;
	wire _w35487_ ;
	wire _w35486_ ;
	wire _w35485_ ;
	wire _w35484_ ;
	wire _w35483_ ;
	wire _w35482_ ;
	wire _w35481_ ;
	wire _w35480_ ;
	wire _w35479_ ;
	wire _w35478_ ;
	wire _w35477_ ;
	wire _w35476_ ;
	wire _w35475_ ;
	wire _w35474_ ;
	wire _w35473_ ;
	wire _w35472_ ;
	wire _w35471_ ;
	wire _w35470_ ;
	wire _w35469_ ;
	wire _w35468_ ;
	wire _w35467_ ;
	wire _w35466_ ;
	wire _w35465_ ;
	wire _w35464_ ;
	wire _w35463_ ;
	wire _w35462_ ;
	wire _w35461_ ;
	wire _w35460_ ;
	wire _w35459_ ;
	wire _w35458_ ;
	wire _w35457_ ;
	wire _w35456_ ;
	wire _w35455_ ;
	wire _w35454_ ;
	wire _w35453_ ;
	wire _w35452_ ;
	wire _w35451_ ;
	wire _w35450_ ;
	wire _w35449_ ;
	wire _w35448_ ;
	wire _w35447_ ;
	wire _w35446_ ;
	wire _w35445_ ;
	wire _w35444_ ;
	wire _w35443_ ;
	wire _w35442_ ;
	wire _w35441_ ;
	wire _w35440_ ;
	wire _w35439_ ;
	wire _w35438_ ;
	wire _w35437_ ;
	wire _w35436_ ;
	wire _w35435_ ;
	wire _w35434_ ;
	wire _w35433_ ;
	wire _w35432_ ;
	wire _w35431_ ;
	wire _w35430_ ;
	wire _w35429_ ;
	wire _w35428_ ;
	wire _w35427_ ;
	wire _w35426_ ;
	wire _w35425_ ;
	wire _w35424_ ;
	wire _w35423_ ;
	wire _w35422_ ;
	wire _w35421_ ;
	wire _w35420_ ;
	wire _w35419_ ;
	wire _w35418_ ;
	wire _w35417_ ;
	wire _w35416_ ;
	wire _w35415_ ;
	wire _w35414_ ;
	wire _w35413_ ;
	wire _w35412_ ;
	wire _w35411_ ;
	wire _w35410_ ;
	wire _w35409_ ;
	wire _w35408_ ;
	wire _w35407_ ;
	wire _w35406_ ;
	wire _w35405_ ;
	wire _w35404_ ;
	wire _w35403_ ;
	wire _w35402_ ;
	wire _w35401_ ;
	wire _w35400_ ;
	wire _w35399_ ;
	wire _w35398_ ;
	wire _w35397_ ;
	wire _w35396_ ;
	wire _w35395_ ;
	wire _w35394_ ;
	wire _w35393_ ;
	wire _w35392_ ;
	wire _w35391_ ;
	wire _w35390_ ;
	wire _w35389_ ;
	wire _w35388_ ;
	wire _w35387_ ;
	wire _w35386_ ;
	wire _w35385_ ;
	wire _w35384_ ;
	wire _w35383_ ;
	wire _w35382_ ;
	wire _w35381_ ;
	wire _w35380_ ;
	wire _w35379_ ;
	wire _w35378_ ;
	wire _w35377_ ;
	wire _w35376_ ;
	wire _w35375_ ;
	wire _w35374_ ;
	wire _w35373_ ;
	wire _w35372_ ;
	wire _w35371_ ;
	wire _w35370_ ;
	wire _w35369_ ;
	wire _w35368_ ;
	wire _w35367_ ;
	wire _w35366_ ;
	wire _w35365_ ;
	wire _w35364_ ;
	wire _w35363_ ;
	wire _w35362_ ;
	wire _w35361_ ;
	wire _w35360_ ;
	wire _w35359_ ;
	wire _w35358_ ;
	wire _w35357_ ;
	wire _w35356_ ;
	wire _w35355_ ;
	wire _w35354_ ;
	wire _w35353_ ;
	wire _w35352_ ;
	wire _w35351_ ;
	wire _w35350_ ;
	wire _w35349_ ;
	wire _w35348_ ;
	wire _w35347_ ;
	wire _w35346_ ;
	wire _w35345_ ;
	wire _w35344_ ;
	wire _w35343_ ;
	wire _w35342_ ;
	wire _w35341_ ;
	wire _w35340_ ;
	wire _w35339_ ;
	wire _w35338_ ;
	wire _w35337_ ;
	wire _w35336_ ;
	wire _w35335_ ;
	wire _w35334_ ;
	wire _w35333_ ;
	wire _w35332_ ;
	wire _w35331_ ;
	wire _w35330_ ;
	wire _w35329_ ;
	wire _w35328_ ;
	wire _w35327_ ;
	wire _w35326_ ;
	wire _w35325_ ;
	wire _w35324_ ;
	wire _w35323_ ;
	wire _w35322_ ;
	wire _w35321_ ;
	wire _w35320_ ;
	wire _w35319_ ;
	wire _w35318_ ;
	wire _w35317_ ;
	wire _w35316_ ;
	wire _w35315_ ;
	wire _w35314_ ;
	wire _w35313_ ;
	wire _w35312_ ;
	wire _w35311_ ;
	wire _w35310_ ;
	wire _w35309_ ;
	wire _w35308_ ;
	wire _w35307_ ;
	wire _w35306_ ;
	wire _w35305_ ;
	wire _w35304_ ;
	wire _w35303_ ;
	wire _w35302_ ;
	wire _w35301_ ;
	wire _w35300_ ;
	wire _w35299_ ;
	wire _w35298_ ;
	wire _w35297_ ;
	wire _w35296_ ;
	wire _w35295_ ;
	wire _w35294_ ;
	wire _w35293_ ;
	wire _w35292_ ;
	wire _w35291_ ;
	wire _w35290_ ;
	wire _w35289_ ;
	wire _w35288_ ;
	wire _w35287_ ;
	wire _w35286_ ;
	wire _w35285_ ;
	wire _w35284_ ;
	wire _w35283_ ;
	wire _w35282_ ;
	wire _w35281_ ;
	wire _w35280_ ;
	wire _w35279_ ;
	wire _w35278_ ;
	wire _w35277_ ;
	wire _w35276_ ;
	wire _w35275_ ;
	wire _w35274_ ;
	wire _w35273_ ;
	wire _w35272_ ;
	wire _w35271_ ;
	wire _w35270_ ;
	wire _w35269_ ;
	wire _w35268_ ;
	wire _w35267_ ;
	wire _w35266_ ;
	wire _w35265_ ;
	wire _w35264_ ;
	wire _w35263_ ;
	wire _w35262_ ;
	wire _w35261_ ;
	wire _w35260_ ;
	wire _w35259_ ;
	wire _w35258_ ;
	wire _w35257_ ;
	wire _w35256_ ;
	wire _w35255_ ;
	wire _w35254_ ;
	wire _w35253_ ;
	wire _w35252_ ;
	wire _w35251_ ;
	wire _w35250_ ;
	wire _w35249_ ;
	wire _w35248_ ;
	wire _w35247_ ;
	wire _w35246_ ;
	wire _w35245_ ;
	wire _w35244_ ;
	wire _w35243_ ;
	wire _w35242_ ;
	wire _w35241_ ;
	wire _w35240_ ;
	wire _w35239_ ;
	wire _w35238_ ;
	wire _w35237_ ;
	wire _w35236_ ;
	wire _w35235_ ;
	wire _w35234_ ;
	wire _w35233_ ;
	wire _w35232_ ;
	wire _w35231_ ;
	wire _w35230_ ;
	wire _w35229_ ;
	wire _w35228_ ;
	wire _w35227_ ;
	wire _w35226_ ;
	wire _w35225_ ;
	wire _w35224_ ;
	wire _w35223_ ;
	wire _w35222_ ;
	wire _w35221_ ;
	wire _w35220_ ;
	wire _w35219_ ;
	wire _w35218_ ;
	wire _w35217_ ;
	wire _w35216_ ;
	wire _w35215_ ;
	wire _w35214_ ;
	wire _w35213_ ;
	wire _w35212_ ;
	wire _w35211_ ;
	wire _w35210_ ;
	wire _w35209_ ;
	wire _w35208_ ;
	wire _w35207_ ;
	wire _w35206_ ;
	wire _w35205_ ;
	wire _w35204_ ;
	wire _w35203_ ;
	wire _w35202_ ;
	wire _w35201_ ;
	wire _w35200_ ;
	wire _w35199_ ;
	wire _w35198_ ;
	wire _w35197_ ;
	wire _w35196_ ;
	wire _w35195_ ;
	wire _w35194_ ;
	wire _w35193_ ;
	wire _w35192_ ;
	wire _w35191_ ;
	wire _w35190_ ;
	wire _w35189_ ;
	wire _w35188_ ;
	wire _w35187_ ;
	wire _w35186_ ;
	wire _w35185_ ;
	wire _w35184_ ;
	wire _w35183_ ;
	wire _w35182_ ;
	wire _w35181_ ;
	wire _w35180_ ;
	wire _w35179_ ;
	wire _w35178_ ;
	wire _w35177_ ;
	wire _w35176_ ;
	wire _w35175_ ;
	wire _w35174_ ;
	wire _w35173_ ;
	wire _w35172_ ;
	wire _w35171_ ;
	wire _w35170_ ;
	wire _w35169_ ;
	wire _w35168_ ;
	wire _w35167_ ;
	wire _w35166_ ;
	wire _w35165_ ;
	wire _w35164_ ;
	wire _w35163_ ;
	wire _w35162_ ;
	wire _w35161_ ;
	wire _w35160_ ;
	wire _w35159_ ;
	wire _w35158_ ;
	wire _w35157_ ;
	wire _w35156_ ;
	wire _w35155_ ;
	wire _w35154_ ;
	wire _w35153_ ;
	wire _w35152_ ;
	wire _w35151_ ;
	wire _w35150_ ;
	wire _w35149_ ;
	wire _w35148_ ;
	wire _w35147_ ;
	wire _w35146_ ;
	wire _w35145_ ;
	wire _w35144_ ;
	wire _w35143_ ;
	wire _w35142_ ;
	wire _w35141_ ;
	wire _w35140_ ;
	wire _w35139_ ;
	wire _w35138_ ;
	wire _w35137_ ;
	wire _w35136_ ;
	wire _w35135_ ;
	wire _w35134_ ;
	wire _w35133_ ;
	wire _w35132_ ;
	wire _w35131_ ;
	wire _w35130_ ;
	wire _w35129_ ;
	wire _w35128_ ;
	wire _w35127_ ;
	wire _w35126_ ;
	wire _w35125_ ;
	wire _w35124_ ;
	wire _w35123_ ;
	wire _w35122_ ;
	wire _w35121_ ;
	wire _w35120_ ;
	wire _w35119_ ;
	wire _w35118_ ;
	wire _w35117_ ;
	wire _w35116_ ;
	wire _w35115_ ;
	wire _w35114_ ;
	wire _w35113_ ;
	wire _w35112_ ;
	wire _w35111_ ;
	wire _w35110_ ;
	wire _w35109_ ;
	wire _w35108_ ;
	wire _w35107_ ;
	wire _w35106_ ;
	wire _w35105_ ;
	wire _w35104_ ;
	wire _w35103_ ;
	wire _w35102_ ;
	wire _w35101_ ;
	wire _w35100_ ;
	wire _w35099_ ;
	wire _w35098_ ;
	wire _w35097_ ;
	wire _w35096_ ;
	wire _w35095_ ;
	wire _w35094_ ;
	wire _w35093_ ;
	wire _w35092_ ;
	wire _w35091_ ;
	wire _w35090_ ;
	wire _w35089_ ;
	wire _w35088_ ;
	wire _w35087_ ;
	wire _w35086_ ;
	wire _w35085_ ;
	wire _w35084_ ;
	wire _w35083_ ;
	wire _w35082_ ;
	wire _w35081_ ;
	wire _w35080_ ;
	wire _w35079_ ;
	wire _w35078_ ;
	wire _w35077_ ;
	wire _w35076_ ;
	wire _w35075_ ;
	wire _w35074_ ;
	wire _w35073_ ;
	wire _w35072_ ;
	wire _w35071_ ;
	wire _w35070_ ;
	wire _w35069_ ;
	wire _w35068_ ;
	wire _w35067_ ;
	wire _w35066_ ;
	wire _w35065_ ;
	wire _w35064_ ;
	wire _w35063_ ;
	wire _w35062_ ;
	wire _w35061_ ;
	wire _w35060_ ;
	wire _w35059_ ;
	wire _w35058_ ;
	wire _w35057_ ;
	wire _w35056_ ;
	wire _w35055_ ;
	wire _w35054_ ;
	wire _w35053_ ;
	wire _w35052_ ;
	wire _w35051_ ;
	wire _w35050_ ;
	wire _w35049_ ;
	wire _w35048_ ;
	wire _w35047_ ;
	wire _w35046_ ;
	wire _w35045_ ;
	wire _w35044_ ;
	wire _w35043_ ;
	wire _w35042_ ;
	wire _w35041_ ;
	wire _w35040_ ;
	wire _w35039_ ;
	wire _w35038_ ;
	wire _w35037_ ;
	wire _w35036_ ;
	wire _w35035_ ;
	wire _w35034_ ;
	wire _w35033_ ;
	wire _w35032_ ;
	wire _w35031_ ;
	wire _w35030_ ;
	wire _w35029_ ;
	wire _w35028_ ;
	wire _w35027_ ;
	wire _w35026_ ;
	wire _w35025_ ;
	wire _w35024_ ;
	wire _w35023_ ;
	wire _w35022_ ;
	wire _w35021_ ;
	wire _w35020_ ;
	wire _w35019_ ;
	wire _w35018_ ;
	wire _w35017_ ;
	wire _w35016_ ;
	wire _w35015_ ;
	wire _w35014_ ;
	wire _w35013_ ;
	wire _w35012_ ;
	wire _w35011_ ;
	wire _w35010_ ;
	wire _w35009_ ;
	wire _w35008_ ;
	wire _w35007_ ;
	wire _w35006_ ;
	wire _w35005_ ;
	wire _w35004_ ;
	wire _w35003_ ;
	wire _w35002_ ;
	wire _w35001_ ;
	wire _w35000_ ;
	wire _w34999_ ;
	wire _w34998_ ;
	wire _w34997_ ;
	wire _w34996_ ;
	wire _w34995_ ;
	wire _w34994_ ;
	wire _w34993_ ;
	wire _w34992_ ;
	wire _w34991_ ;
	wire _w34990_ ;
	wire _w34989_ ;
	wire _w34988_ ;
	wire _w34987_ ;
	wire _w34986_ ;
	wire _w34985_ ;
	wire _w34984_ ;
	wire _w34983_ ;
	wire _w34982_ ;
	wire _w34981_ ;
	wire _w34980_ ;
	wire _w34979_ ;
	wire _w34978_ ;
	wire _w34977_ ;
	wire _w34976_ ;
	wire _w34975_ ;
	wire _w34974_ ;
	wire _w34973_ ;
	wire _w34972_ ;
	wire _w34971_ ;
	wire _w34970_ ;
	wire _w34969_ ;
	wire _w34968_ ;
	wire _w34967_ ;
	wire _w34966_ ;
	wire _w34965_ ;
	wire _w34964_ ;
	wire _w34963_ ;
	wire _w34962_ ;
	wire _w34961_ ;
	wire _w34960_ ;
	wire _w34959_ ;
	wire _w34958_ ;
	wire _w34957_ ;
	wire _w34956_ ;
	wire _w34955_ ;
	wire _w34954_ ;
	wire _w34953_ ;
	wire _w34952_ ;
	wire _w34951_ ;
	wire _w34950_ ;
	wire _w34949_ ;
	wire _w34948_ ;
	wire _w34947_ ;
	wire _w34946_ ;
	wire _w34945_ ;
	wire _w34944_ ;
	wire _w34943_ ;
	wire _w34942_ ;
	wire _w34941_ ;
	wire _w34940_ ;
	wire _w34939_ ;
	wire _w34938_ ;
	wire _w34937_ ;
	wire _w34936_ ;
	wire _w34935_ ;
	wire _w34934_ ;
	wire _w34933_ ;
	wire _w34932_ ;
	wire _w34931_ ;
	wire _w34930_ ;
	wire _w34929_ ;
	wire _w34928_ ;
	wire _w34927_ ;
	wire _w34926_ ;
	wire _w34925_ ;
	wire _w34924_ ;
	wire _w34923_ ;
	wire _w34922_ ;
	wire _w34921_ ;
	wire _w34920_ ;
	wire _w34919_ ;
	wire _w34918_ ;
	wire _w34917_ ;
	wire _w34916_ ;
	wire _w34915_ ;
	wire _w34914_ ;
	wire _w34913_ ;
	wire _w34912_ ;
	wire _w34911_ ;
	wire _w34910_ ;
	wire _w34909_ ;
	wire _w34908_ ;
	wire _w34907_ ;
	wire _w34906_ ;
	wire _w34905_ ;
	wire _w34904_ ;
	wire _w34903_ ;
	wire _w34902_ ;
	wire _w34901_ ;
	wire _w34900_ ;
	wire _w34899_ ;
	wire _w34898_ ;
	wire _w34897_ ;
	wire _w34896_ ;
	wire _w34895_ ;
	wire _w34894_ ;
	wire _w34893_ ;
	wire _w34892_ ;
	wire _w34891_ ;
	wire _w34890_ ;
	wire _w34889_ ;
	wire _w34888_ ;
	wire _w34887_ ;
	wire _w34886_ ;
	wire _w34885_ ;
	wire _w34884_ ;
	wire _w34883_ ;
	wire _w34882_ ;
	wire _w34881_ ;
	wire _w34880_ ;
	wire _w34879_ ;
	wire _w34878_ ;
	wire _w34877_ ;
	wire _w34876_ ;
	wire _w34875_ ;
	wire _w34874_ ;
	wire _w34873_ ;
	wire _w34872_ ;
	wire _w34871_ ;
	wire _w34870_ ;
	wire _w34869_ ;
	wire _w34868_ ;
	wire _w34867_ ;
	wire _w34866_ ;
	wire _w34865_ ;
	wire _w34864_ ;
	wire _w34863_ ;
	wire _w34862_ ;
	wire _w34861_ ;
	wire _w34860_ ;
	wire _w34859_ ;
	wire _w34858_ ;
	wire _w34857_ ;
	wire _w34856_ ;
	wire _w34855_ ;
	wire _w34854_ ;
	wire _w34853_ ;
	wire _w34852_ ;
	wire _w34851_ ;
	wire _w34850_ ;
	wire _w34849_ ;
	wire _w34848_ ;
	wire _w34847_ ;
	wire _w34846_ ;
	wire _w34845_ ;
	wire _w34844_ ;
	wire _w34843_ ;
	wire _w34842_ ;
	wire _w34841_ ;
	wire _w34840_ ;
	wire _w34839_ ;
	wire _w34838_ ;
	wire _w34837_ ;
	wire _w34836_ ;
	wire _w34835_ ;
	wire _w34834_ ;
	wire _w34833_ ;
	wire _w34832_ ;
	wire _w34831_ ;
	wire _w34830_ ;
	wire _w34829_ ;
	wire _w34828_ ;
	wire _w34827_ ;
	wire _w34826_ ;
	wire _w34825_ ;
	wire _w34824_ ;
	wire _w34823_ ;
	wire _w34822_ ;
	wire _w34821_ ;
	wire _w34820_ ;
	wire _w34819_ ;
	wire _w34818_ ;
	wire _w34817_ ;
	wire _w34816_ ;
	wire _w34815_ ;
	wire _w34814_ ;
	wire _w34813_ ;
	wire _w34812_ ;
	wire _w34811_ ;
	wire _w34810_ ;
	wire _w34809_ ;
	wire _w34808_ ;
	wire _w34807_ ;
	wire _w34806_ ;
	wire _w34805_ ;
	wire _w34804_ ;
	wire _w34803_ ;
	wire _w34802_ ;
	wire _w34801_ ;
	wire _w34800_ ;
	wire _w34799_ ;
	wire _w34798_ ;
	wire _w34797_ ;
	wire _w34796_ ;
	wire _w34795_ ;
	wire _w34794_ ;
	wire _w34793_ ;
	wire _w34792_ ;
	wire _w34791_ ;
	wire _w34790_ ;
	wire _w34789_ ;
	wire _w34788_ ;
	wire _w34787_ ;
	wire _w34786_ ;
	wire _w34785_ ;
	wire _w34784_ ;
	wire _w34783_ ;
	wire _w34782_ ;
	wire _w34781_ ;
	wire _w34780_ ;
	wire _w34779_ ;
	wire _w34778_ ;
	wire _w34777_ ;
	wire _w34776_ ;
	wire _w34775_ ;
	wire _w34774_ ;
	wire _w34773_ ;
	wire _w34772_ ;
	wire _w34771_ ;
	wire _w34770_ ;
	wire _w34769_ ;
	wire _w34768_ ;
	wire _w34767_ ;
	wire _w34766_ ;
	wire _w34765_ ;
	wire _w34764_ ;
	wire _w34763_ ;
	wire _w34762_ ;
	wire _w34761_ ;
	wire _w34760_ ;
	wire _w34759_ ;
	wire _w34758_ ;
	wire _w34757_ ;
	wire _w34756_ ;
	wire _w34755_ ;
	wire _w34754_ ;
	wire _w34753_ ;
	wire _w34752_ ;
	wire _w34751_ ;
	wire _w34750_ ;
	wire _w34749_ ;
	wire _w34748_ ;
	wire _w34747_ ;
	wire _w34746_ ;
	wire _w34745_ ;
	wire _w34744_ ;
	wire _w34743_ ;
	wire _w34742_ ;
	wire _w34741_ ;
	wire _w34740_ ;
	wire _w34739_ ;
	wire _w34738_ ;
	wire _w34737_ ;
	wire _w34736_ ;
	wire _w34735_ ;
	wire _w34734_ ;
	wire _w34733_ ;
	wire _w34732_ ;
	wire _w34731_ ;
	wire _w34730_ ;
	wire _w34729_ ;
	wire _w34728_ ;
	wire _w34727_ ;
	wire _w34726_ ;
	wire _w34725_ ;
	wire _w34724_ ;
	wire _w34723_ ;
	wire _w34722_ ;
	wire _w34721_ ;
	wire _w34720_ ;
	wire _w34719_ ;
	wire _w34718_ ;
	wire _w34717_ ;
	wire _w34716_ ;
	wire _w34715_ ;
	wire _w34714_ ;
	wire _w34713_ ;
	wire _w34712_ ;
	wire _w34711_ ;
	wire _w34710_ ;
	wire _w34709_ ;
	wire _w34708_ ;
	wire _w34707_ ;
	wire _w34706_ ;
	wire _w34705_ ;
	wire _w34704_ ;
	wire _w34703_ ;
	wire _w34702_ ;
	wire _w34701_ ;
	wire _w34700_ ;
	wire _w34699_ ;
	wire _w34698_ ;
	wire _w34697_ ;
	wire _w34696_ ;
	wire _w34695_ ;
	wire _w34694_ ;
	wire _w34693_ ;
	wire _w34692_ ;
	wire _w34691_ ;
	wire _w34690_ ;
	wire _w34689_ ;
	wire _w34688_ ;
	wire _w34687_ ;
	wire _w34686_ ;
	wire _w34685_ ;
	wire _w34684_ ;
	wire _w34683_ ;
	wire _w34682_ ;
	wire _w34681_ ;
	wire _w34680_ ;
	wire _w34679_ ;
	wire _w34678_ ;
	wire _w34677_ ;
	wire _w34676_ ;
	wire _w34675_ ;
	wire _w34674_ ;
	wire _w34673_ ;
	wire _w34672_ ;
	wire _w34671_ ;
	wire _w34670_ ;
	wire _w34669_ ;
	wire _w34668_ ;
	wire _w34667_ ;
	wire _w34666_ ;
	wire _w34665_ ;
	wire _w34664_ ;
	wire _w34663_ ;
	wire _w34662_ ;
	wire _w34661_ ;
	wire _w34660_ ;
	wire _w34659_ ;
	wire _w34658_ ;
	wire _w34657_ ;
	wire _w34656_ ;
	wire _w34655_ ;
	wire _w34654_ ;
	wire _w34653_ ;
	wire _w34652_ ;
	wire _w34651_ ;
	wire _w34650_ ;
	wire _w34649_ ;
	wire _w34648_ ;
	wire _w34647_ ;
	wire _w34646_ ;
	wire _w34645_ ;
	wire _w34644_ ;
	wire _w34643_ ;
	wire _w34642_ ;
	wire _w34641_ ;
	wire _w34640_ ;
	wire _w34639_ ;
	wire _w34638_ ;
	wire _w34637_ ;
	wire _w34636_ ;
	wire _w34635_ ;
	wire _w34634_ ;
	wire _w34633_ ;
	wire _w34632_ ;
	wire _w34631_ ;
	wire _w34630_ ;
	wire _w34629_ ;
	wire _w34628_ ;
	wire _w34627_ ;
	wire _w34626_ ;
	wire _w34625_ ;
	wire _w34624_ ;
	wire _w34623_ ;
	wire _w34622_ ;
	wire _w34621_ ;
	wire _w34620_ ;
	wire _w34619_ ;
	wire _w34618_ ;
	wire _w34617_ ;
	wire _w34616_ ;
	wire _w34615_ ;
	wire _w34614_ ;
	wire _w34613_ ;
	wire _w34612_ ;
	wire _w34611_ ;
	wire _w34610_ ;
	wire _w34609_ ;
	wire _w34608_ ;
	wire _w34607_ ;
	wire _w34606_ ;
	wire _w34605_ ;
	wire _w34604_ ;
	wire _w34603_ ;
	wire _w34602_ ;
	wire _w34601_ ;
	wire _w34600_ ;
	wire _w34599_ ;
	wire _w34598_ ;
	wire _w34597_ ;
	wire _w34596_ ;
	wire _w34595_ ;
	wire _w34594_ ;
	wire _w34593_ ;
	wire _w34592_ ;
	wire _w34591_ ;
	wire _w34590_ ;
	wire _w34589_ ;
	wire _w34588_ ;
	wire _w34587_ ;
	wire _w34586_ ;
	wire _w34585_ ;
	wire _w34584_ ;
	wire _w34583_ ;
	wire _w34582_ ;
	wire _w34581_ ;
	wire _w34580_ ;
	wire _w34579_ ;
	wire _w34578_ ;
	wire _w34577_ ;
	wire _w34576_ ;
	wire _w34575_ ;
	wire _w34574_ ;
	wire _w34573_ ;
	wire _w34572_ ;
	wire _w34571_ ;
	wire _w34570_ ;
	wire _w34569_ ;
	wire _w34568_ ;
	wire _w34567_ ;
	wire _w34566_ ;
	wire _w34565_ ;
	wire _w34564_ ;
	wire _w34563_ ;
	wire _w34562_ ;
	wire _w34561_ ;
	wire _w34560_ ;
	wire _w34559_ ;
	wire _w34558_ ;
	wire _w34557_ ;
	wire _w34556_ ;
	wire _w34555_ ;
	wire _w34554_ ;
	wire _w34553_ ;
	wire _w34552_ ;
	wire _w34551_ ;
	wire _w34550_ ;
	wire _w34549_ ;
	wire _w34548_ ;
	wire _w34547_ ;
	wire _w34546_ ;
	wire _w34545_ ;
	wire _w34544_ ;
	wire _w34543_ ;
	wire _w34542_ ;
	wire _w34541_ ;
	wire _w34540_ ;
	wire _w34539_ ;
	wire _w34538_ ;
	wire _w34537_ ;
	wire _w34536_ ;
	wire _w34535_ ;
	wire _w34534_ ;
	wire _w34533_ ;
	wire _w34532_ ;
	wire _w34531_ ;
	wire _w34530_ ;
	wire _w34529_ ;
	wire _w34528_ ;
	wire _w34527_ ;
	wire _w34526_ ;
	wire _w34525_ ;
	wire _w34524_ ;
	wire _w34523_ ;
	wire _w34522_ ;
	wire _w34521_ ;
	wire _w34520_ ;
	wire _w34519_ ;
	wire _w34518_ ;
	wire _w34517_ ;
	wire _w34516_ ;
	wire _w34515_ ;
	wire _w34514_ ;
	wire _w34513_ ;
	wire _w34512_ ;
	wire _w34511_ ;
	wire _w34510_ ;
	wire _w34509_ ;
	wire _w34508_ ;
	wire _w34507_ ;
	wire _w34506_ ;
	wire _w34505_ ;
	wire _w34504_ ;
	wire _w34503_ ;
	wire _w34502_ ;
	wire _w34501_ ;
	wire _w34500_ ;
	wire _w34499_ ;
	wire _w34498_ ;
	wire _w34497_ ;
	wire _w34496_ ;
	wire _w34495_ ;
	wire _w34494_ ;
	wire _w34493_ ;
	wire _w34492_ ;
	wire _w34491_ ;
	wire _w34490_ ;
	wire _w34489_ ;
	wire _w34488_ ;
	wire _w34487_ ;
	wire _w34486_ ;
	wire _w34485_ ;
	wire _w34484_ ;
	wire _w34483_ ;
	wire _w34482_ ;
	wire _w34481_ ;
	wire _w34480_ ;
	wire _w34479_ ;
	wire _w34478_ ;
	wire _w34477_ ;
	wire _w34476_ ;
	wire _w34475_ ;
	wire _w34474_ ;
	wire _w34473_ ;
	wire _w34472_ ;
	wire _w34471_ ;
	wire _w34470_ ;
	wire _w34469_ ;
	wire _w34468_ ;
	wire _w34467_ ;
	wire _w34466_ ;
	wire _w34465_ ;
	wire _w34464_ ;
	wire _w34463_ ;
	wire _w34462_ ;
	wire _w34461_ ;
	wire _w34460_ ;
	wire _w34459_ ;
	wire _w34458_ ;
	wire _w34457_ ;
	wire _w34456_ ;
	wire _w34455_ ;
	wire _w34454_ ;
	wire _w34453_ ;
	wire _w34452_ ;
	wire _w34451_ ;
	wire _w34450_ ;
	wire _w34449_ ;
	wire _w34448_ ;
	wire _w34447_ ;
	wire _w34446_ ;
	wire _w34445_ ;
	wire _w34444_ ;
	wire _w34443_ ;
	wire _w34442_ ;
	wire _w34441_ ;
	wire _w34440_ ;
	wire _w34439_ ;
	wire _w34438_ ;
	wire _w34437_ ;
	wire _w34436_ ;
	wire _w34435_ ;
	wire _w34434_ ;
	wire _w34433_ ;
	wire _w34432_ ;
	wire _w34431_ ;
	wire _w34430_ ;
	wire _w34429_ ;
	wire _w34428_ ;
	wire _w34427_ ;
	wire _w34426_ ;
	wire _w34425_ ;
	wire _w34424_ ;
	wire _w34423_ ;
	wire _w34422_ ;
	wire _w34421_ ;
	wire _w34420_ ;
	wire _w34419_ ;
	wire _w34418_ ;
	wire _w34417_ ;
	wire _w34416_ ;
	wire _w34415_ ;
	wire _w34414_ ;
	wire _w34413_ ;
	wire _w34412_ ;
	wire _w34411_ ;
	wire _w34410_ ;
	wire _w34409_ ;
	wire _w34408_ ;
	wire _w34407_ ;
	wire _w34406_ ;
	wire _w34405_ ;
	wire _w34404_ ;
	wire _w34403_ ;
	wire _w34402_ ;
	wire _w34401_ ;
	wire _w34400_ ;
	wire _w34399_ ;
	wire _w34398_ ;
	wire _w34397_ ;
	wire _w34396_ ;
	wire _w34395_ ;
	wire _w34394_ ;
	wire _w34393_ ;
	wire _w34392_ ;
	wire _w34391_ ;
	wire _w34390_ ;
	wire _w34389_ ;
	wire _w34388_ ;
	wire _w34387_ ;
	wire _w34386_ ;
	wire _w34385_ ;
	wire _w34384_ ;
	wire _w34383_ ;
	wire _w34382_ ;
	wire _w34381_ ;
	wire _w34380_ ;
	wire _w34379_ ;
	wire _w34378_ ;
	wire _w34377_ ;
	wire _w34376_ ;
	wire _w34375_ ;
	wire _w34374_ ;
	wire _w34373_ ;
	wire _w34372_ ;
	wire _w34371_ ;
	wire _w34370_ ;
	wire _w34369_ ;
	wire _w34368_ ;
	wire _w34367_ ;
	wire _w34366_ ;
	wire _w34365_ ;
	wire _w34364_ ;
	wire _w34363_ ;
	wire _w34362_ ;
	wire _w34361_ ;
	wire _w34360_ ;
	wire _w34359_ ;
	wire _w34358_ ;
	wire _w34357_ ;
	wire _w34356_ ;
	wire _w34355_ ;
	wire _w34354_ ;
	wire _w34353_ ;
	wire _w34352_ ;
	wire _w34351_ ;
	wire _w34350_ ;
	wire _w34349_ ;
	wire _w34348_ ;
	wire _w34347_ ;
	wire _w34346_ ;
	wire _w34345_ ;
	wire _w34344_ ;
	wire _w34343_ ;
	wire _w34342_ ;
	wire _w34341_ ;
	wire _w34340_ ;
	wire _w34339_ ;
	wire _w34338_ ;
	wire _w34337_ ;
	wire _w34336_ ;
	wire _w34335_ ;
	wire _w34334_ ;
	wire _w34333_ ;
	wire _w34332_ ;
	wire _w34331_ ;
	wire _w34330_ ;
	wire _w34329_ ;
	wire _w34328_ ;
	wire _w34327_ ;
	wire _w34326_ ;
	wire _w34325_ ;
	wire _w34324_ ;
	wire _w34323_ ;
	wire _w34322_ ;
	wire _w34321_ ;
	wire _w34320_ ;
	wire _w34319_ ;
	wire _w34318_ ;
	wire _w34317_ ;
	wire _w34316_ ;
	wire _w34315_ ;
	wire _w34314_ ;
	wire _w34313_ ;
	wire _w34312_ ;
	wire _w34311_ ;
	wire _w34310_ ;
	wire _w34309_ ;
	wire _w34308_ ;
	wire _w34307_ ;
	wire _w34306_ ;
	wire _w34305_ ;
	wire _w34304_ ;
	wire _w34303_ ;
	wire _w34302_ ;
	wire _w34301_ ;
	wire _w34300_ ;
	wire _w34299_ ;
	wire _w34298_ ;
	wire _w34297_ ;
	wire _w34296_ ;
	wire _w34295_ ;
	wire _w34294_ ;
	wire _w34293_ ;
	wire _w34292_ ;
	wire _w34291_ ;
	wire _w34290_ ;
	wire _w34289_ ;
	wire _w34288_ ;
	wire _w34287_ ;
	wire _w34286_ ;
	wire _w34285_ ;
	wire _w34284_ ;
	wire _w34283_ ;
	wire _w34282_ ;
	wire _w34281_ ;
	wire _w34280_ ;
	wire _w34279_ ;
	wire _w34278_ ;
	wire _w34277_ ;
	wire _w34276_ ;
	wire _w34275_ ;
	wire _w34274_ ;
	wire _w34273_ ;
	wire _w34272_ ;
	wire _w34271_ ;
	wire _w34270_ ;
	wire _w34269_ ;
	wire _w34268_ ;
	wire _w34267_ ;
	wire _w34266_ ;
	wire _w34265_ ;
	wire _w34264_ ;
	wire _w34263_ ;
	wire _w34262_ ;
	wire _w34261_ ;
	wire _w34260_ ;
	wire _w34259_ ;
	wire _w34258_ ;
	wire _w34257_ ;
	wire _w34256_ ;
	wire _w34255_ ;
	wire _w34254_ ;
	wire _w34253_ ;
	wire _w34252_ ;
	wire _w34251_ ;
	wire _w34250_ ;
	wire _w34249_ ;
	wire _w34248_ ;
	wire _w34247_ ;
	wire _w34246_ ;
	wire _w34245_ ;
	wire _w34244_ ;
	wire _w34243_ ;
	wire _w34242_ ;
	wire _w34241_ ;
	wire _w34240_ ;
	wire _w34239_ ;
	wire _w34238_ ;
	wire _w34237_ ;
	wire _w34236_ ;
	wire _w34235_ ;
	wire _w34234_ ;
	wire _w34233_ ;
	wire _w34232_ ;
	wire _w34231_ ;
	wire _w34230_ ;
	wire _w34229_ ;
	wire _w34228_ ;
	wire _w34227_ ;
	wire _w34226_ ;
	wire _w34225_ ;
	wire _w34224_ ;
	wire _w34223_ ;
	wire _w34222_ ;
	wire _w34221_ ;
	wire _w34220_ ;
	wire _w34219_ ;
	wire _w34218_ ;
	wire _w34217_ ;
	wire _w34216_ ;
	wire _w34215_ ;
	wire _w34214_ ;
	wire _w34213_ ;
	wire _w34212_ ;
	wire _w34211_ ;
	wire _w34210_ ;
	wire _w34209_ ;
	wire _w34208_ ;
	wire _w34207_ ;
	wire _w34206_ ;
	wire _w34205_ ;
	wire _w34204_ ;
	wire _w34203_ ;
	wire _w34202_ ;
	wire _w34201_ ;
	wire _w34200_ ;
	wire _w34199_ ;
	wire _w34198_ ;
	wire _w34197_ ;
	wire _w34196_ ;
	wire _w34195_ ;
	wire _w34194_ ;
	wire _w34193_ ;
	wire _w34192_ ;
	wire _w34191_ ;
	wire _w34190_ ;
	wire _w34189_ ;
	wire _w34188_ ;
	wire _w34187_ ;
	wire _w34186_ ;
	wire _w34185_ ;
	wire _w34184_ ;
	wire _w34183_ ;
	wire _w34182_ ;
	wire _w34181_ ;
	wire _w34180_ ;
	wire _w34179_ ;
	wire _w34178_ ;
	wire _w34177_ ;
	wire _w34176_ ;
	wire _w34175_ ;
	wire _w34174_ ;
	wire _w34173_ ;
	wire _w34172_ ;
	wire _w34171_ ;
	wire _w34170_ ;
	wire _w34169_ ;
	wire _w34168_ ;
	wire _w34167_ ;
	wire _w34166_ ;
	wire _w34165_ ;
	wire _w34164_ ;
	wire _w34163_ ;
	wire _w34162_ ;
	wire _w34161_ ;
	wire _w34160_ ;
	wire _w34159_ ;
	wire _w34158_ ;
	wire _w34157_ ;
	wire _w34156_ ;
	wire _w34155_ ;
	wire _w34154_ ;
	wire _w34153_ ;
	wire _w34152_ ;
	wire _w34151_ ;
	wire _w34150_ ;
	wire _w34149_ ;
	wire _w34148_ ;
	wire _w34147_ ;
	wire _w34146_ ;
	wire _w34145_ ;
	wire _w34144_ ;
	wire _w34143_ ;
	wire _w34142_ ;
	wire _w34141_ ;
	wire _w34140_ ;
	wire _w34139_ ;
	wire _w34138_ ;
	wire _w34137_ ;
	wire _w34136_ ;
	wire _w34135_ ;
	wire _w34134_ ;
	wire _w34133_ ;
	wire _w34132_ ;
	wire _w34131_ ;
	wire _w34130_ ;
	wire _w34129_ ;
	wire _w34128_ ;
	wire _w34127_ ;
	wire _w34126_ ;
	wire _w34125_ ;
	wire _w34124_ ;
	wire _w34123_ ;
	wire _w34122_ ;
	wire _w34121_ ;
	wire _w34120_ ;
	wire _w34119_ ;
	wire _w34118_ ;
	wire _w34117_ ;
	wire _w34116_ ;
	wire _w34115_ ;
	wire _w34114_ ;
	wire _w34113_ ;
	wire _w34112_ ;
	wire _w34111_ ;
	wire _w34110_ ;
	wire _w34109_ ;
	wire _w34108_ ;
	wire _w34107_ ;
	wire _w34106_ ;
	wire _w34105_ ;
	wire _w34104_ ;
	wire _w34103_ ;
	wire _w34102_ ;
	wire _w34101_ ;
	wire _w34100_ ;
	wire _w34099_ ;
	wire _w34098_ ;
	wire _w34097_ ;
	wire _w34096_ ;
	wire _w34095_ ;
	wire _w34094_ ;
	wire _w34093_ ;
	wire _w34092_ ;
	wire _w34091_ ;
	wire _w34090_ ;
	wire _w34089_ ;
	wire _w34088_ ;
	wire _w34087_ ;
	wire _w34086_ ;
	wire _w34085_ ;
	wire _w34084_ ;
	wire _w34083_ ;
	wire _w34082_ ;
	wire _w34081_ ;
	wire _w34080_ ;
	wire _w34079_ ;
	wire _w34078_ ;
	wire _w34077_ ;
	wire _w34076_ ;
	wire _w34075_ ;
	wire _w34074_ ;
	wire _w34073_ ;
	wire _w34072_ ;
	wire _w34071_ ;
	wire _w34070_ ;
	wire _w34069_ ;
	wire _w34068_ ;
	wire _w34067_ ;
	wire _w34066_ ;
	wire _w34065_ ;
	wire _w34064_ ;
	wire _w34063_ ;
	wire _w34062_ ;
	wire _w34061_ ;
	wire _w34060_ ;
	wire _w34059_ ;
	wire _w34058_ ;
	wire _w34057_ ;
	wire _w34056_ ;
	wire _w34055_ ;
	wire _w34054_ ;
	wire _w34053_ ;
	wire _w34052_ ;
	wire _w34051_ ;
	wire _w34050_ ;
	wire _w34049_ ;
	wire _w34048_ ;
	wire _w34047_ ;
	wire _w34046_ ;
	wire _w34045_ ;
	wire _w34044_ ;
	wire _w34043_ ;
	wire _w34042_ ;
	wire _w34041_ ;
	wire _w34040_ ;
	wire _w34039_ ;
	wire _w34038_ ;
	wire _w34037_ ;
	wire _w34036_ ;
	wire _w34035_ ;
	wire _w34034_ ;
	wire _w34033_ ;
	wire _w34032_ ;
	wire _w34031_ ;
	wire _w34030_ ;
	wire _w34029_ ;
	wire _w34028_ ;
	wire _w34027_ ;
	wire _w34026_ ;
	wire _w34025_ ;
	wire _w34024_ ;
	wire _w34023_ ;
	wire _w34022_ ;
	wire _w34021_ ;
	wire _w34020_ ;
	wire _w34019_ ;
	wire _w34018_ ;
	wire _w34017_ ;
	wire _w34016_ ;
	wire _w34015_ ;
	wire _w34014_ ;
	wire _w34013_ ;
	wire _w34012_ ;
	wire _w34011_ ;
	wire _w34010_ ;
	wire _w34009_ ;
	wire _w34008_ ;
	wire _w34007_ ;
	wire _w34006_ ;
	wire _w34005_ ;
	wire _w34004_ ;
	wire _w34003_ ;
	wire _w34002_ ;
	wire _w34001_ ;
	wire _w34000_ ;
	wire _w33999_ ;
	wire _w33998_ ;
	wire _w33997_ ;
	wire _w33996_ ;
	wire _w33995_ ;
	wire _w33994_ ;
	wire _w33993_ ;
	wire _w33992_ ;
	wire _w33991_ ;
	wire _w33990_ ;
	wire _w33989_ ;
	wire _w33988_ ;
	wire _w33987_ ;
	wire _w33986_ ;
	wire _w33985_ ;
	wire _w33984_ ;
	wire _w33983_ ;
	wire _w33982_ ;
	wire _w33981_ ;
	wire _w33980_ ;
	wire _w33979_ ;
	wire _w33978_ ;
	wire _w33977_ ;
	wire _w33976_ ;
	wire _w33975_ ;
	wire _w33974_ ;
	wire _w33973_ ;
	wire _w33972_ ;
	wire _w33971_ ;
	wire _w33970_ ;
	wire _w33969_ ;
	wire _w33968_ ;
	wire _w33967_ ;
	wire _w33966_ ;
	wire _w33965_ ;
	wire _w33964_ ;
	wire _w33963_ ;
	wire _w33962_ ;
	wire _w33961_ ;
	wire _w33960_ ;
	wire _w33959_ ;
	wire _w33958_ ;
	wire _w33957_ ;
	wire _w33956_ ;
	wire _w33955_ ;
	wire _w33954_ ;
	wire _w33953_ ;
	wire _w33952_ ;
	wire _w33951_ ;
	wire _w33950_ ;
	wire _w33949_ ;
	wire _w33948_ ;
	wire _w33947_ ;
	wire _w33946_ ;
	wire _w33945_ ;
	wire _w33944_ ;
	wire _w33943_ ;
	wire _w33942_ ;
	wire _w33941_ ;
	wire _w33940_ ;
	wire _w33939_ ;
	wire _w33938_ ;
	wire _w33937_ ;
	wire _w33936_ ;
	wire _w33935_ ;
	wire _w33934_ ;
	wire _w33933_ ;
	wire _w33932_ ;
	wire _w33931_ ;
	wire _w33930_ ;
	wire _w33929_ ;
	wire _w33928_ ;
	wire _w33927_ ;
	wire _w33926_ ;
	wire _w33925_ ;
	wire _w33924_ ;
	wire _w33923_ ;
	wire _w33922_ ;
	wire _w33921_ ;
	wire _w33920_ ;
	wire _w33919_ ;
	wire _w33918_ ;
	wire _w33917_ ;
	wire _w33916_ ;
	wire _w33915_ ;
	wire _w33914_ ;
	wire _w33913_ ;
	wire _w33912_ ;
	wire _w33911_ ;
	wire _w33910_ ;
	wire _w33909_ ;
	wire _w33908_ ;
	wire _w33907_ ;
	wire _w33906_ ;
	wire _w33905_ ;
	wire _w33904_ ;
	wire _w33903_ ;
	wire _w33902_ ;
	wire _w33901_ ;
	wire _w33900_ ;
	wire _w33899_ ;
	wire _w33898_ ;
	wire _w33897_ ;
	wire _w33896_ ;
	wire _w33895_ ;
	wire _w33894_ ;
	wire _w33893_ ;
	wire _w33892_ ;
	wire _w33891_ ;
	wire _w33890_ ;
	wire _w33889_ ;
	wire _w33888_ ;
	wire _w33887_ ;
	wire _w33886_ ;
	wire _w33885_ ;
	wire _w33884_ ;
	wire _w33883_ ;
	wire _w33882_ ;
	wire _w33881_ ;
	wire _w33880_ ;
	wire _w33879_ ;
	wire _w33878_ ;
	wire _w33877_ ;
	wire _w33876_ ;
	wire _w33875_ ;
	wire _w33874_ ;
	wire _w33873_ ;
	wire _w33872_ ;
	wire _w33871_ ;
	wire _w33870_ ;
	wire _w33869_ ;
	wire _w33868_ ;
	wire _w33867_ ;
	wire _w33866_ ;
	wire _w33865_ ;
	wire _w33864_ ;
	wire _w33863_ ;
	wire _w33862_ ;
	wire _w33861_ ;
	wire _w33860_ ;
	wire _w33859_ ;
	wire _w33858_ ;
	wire _w33857_ ;
	wire _w33856_ ;
	wire _w33855_ ;
	wire _w33854_ ;
	wire _w33853_ ;
	wire _w33852_ ;
	wire _w33851_ ;
	wire _w33850_ ;
	wire _w33849_ ;
	wire _w33848_ ;
	wire _w33847_ ;
	wire _w33846_ ;
	wire _w33845_ ;
	wire _w33844_ ;
	wire _w33843_ ;
	wire _w33842_ ;
	wire _w33841_ ;
	wire _w33840_ ;
	wire _w33839_ ;
	wire _w33838_ ;
	wire _w33837_ ;
	wire _w33836_ ;
	wire _w33835_ ;
	wire _w33834_ ;
	wire _w33833_ ;
	wire _w33832_ ;
	wire _w33831_ ;
	wire _w33830_ ;
	wire _w33829_ ;
	wire _w33828_ ;
	wire _w33827_ ;
	wire _w33826_ ;
	wire _w33825_ ;
	wire _w33824_ ;
	wire _w33823_ ;
	wire _w33822_ ;
	wire _w33821_ ;
	wire _w33820_ ;
	wire _w33819_ ;
	wire _w33818_ ;
	wire _w33817_ ;
	wire _w33816_ ;
	wire _w33815_ ;
	wire _w33814_ ;
	wire _w33813_ ;
	wire _w33812_ ;
	wire _w33811_ ;
	wire _w33810_ ;
	wire _w33809_ ;
	wire _w33808_ ;
	wire _w33807_ ;
	wire _w33806_ ;
	wire _w33805_ ;
	wire _w33804_ ;
	wire _w33803_ ;
	wire _w33802_ ;
	wire _w33801_ ;
	wire _w33800_ ;
	wire _w33799_ ;
	wire _w33798_ ;
	wire _w33797_ ;
	wire _w33796_ ;
	wire _w33795_ ;
	wire _w33794_ ;
	wire _w33793_ ;
	wire _w33792_ ;
	wire _w33791_ ;
	wire _w33790_ ;
	wire _w33789_ ;
	wire _w33788_ ;
	wire _w33787_ ;
	wire _w33786_ ;
	wire _w33785_ ;
	wire _w33784_ ;
	wire _w33783_ ;
	wire _w33782_ ;
	wire _w33781_ ;
	wire _w33780_ ;
	wire _w33779_ ;
	wire _w33778_ ;
	wire _w33777_ ;
	wire _w33776_ ;
	wire _w33775_ ;
	wire _w33774_ ;
	wire _w33773_ ;
	wire _w33772_ ;
	wire _w33771_ ;
	wire _w33770_ ;
	wire _w33769_ ;
	wire _w33768_ ;
	wire _w33767_ ;
	wire _w33766_ ;
	wire _w33765_ ;
	wire _w33764_ ;
	wire _w33763_ ;
	wire _w33762_ ;
	wire _w33761_ ;
	wire _w33760_ ;
	wire _w33759_ ;
	wire _w33758_ ;
	wire _w33757_ ;
	wire _w33756_ ;
	wire _w33755_ ;
	wire _w33754_ ;
	wire _w33753_ ;
	wire _w33752_ ;
	wire _w33751_ ;
	wire _w33750_ ;
	wire _w33749_ ;
	wire _w33748_ ;
	wire _w33747_ ;
	wire _w33746_ ;
	wire _w33745_ ;
	wire _w33744_ ;
	wire _w33743_ ;
	wire _w33742_ ;
	wire _w33741_ ;
	wire _w33740_ ;
	wire _w33739_ ;
	wire _w33738_ ;
	wire _w33737_ ;
	wire _w33736_ ;
	wire _w33735_ ;
	wire _w33734_ ;
	wire _w33733_ ;
	wire _w33732_ ;
	wire _w33731_ ;
	wire _w33730_ ;
	wire _w33729_ ;
	wire _w33728_ ;
	wire _w33727_ ;
	wire _w33726_ ;
	wire _w33725_ ;
	wire _w33724_ ;
	wire _w33723_ ;
	wire _w33722_ ;
	wire _w33721_ ;
	wire _w33720_ ;
	wire _w33719_ ;
	wire _w33718_ ;
	wire _w33717_ ;
	wire _w33716_ ;
	wire _w33715_ ;
	wire _w33714_ ;
	wire _w33713_ ;
	wire _w33712_ ;
	wire _w33711_ ;
	wire _w33710_ ;
	wire _w33709_ ;
	wire _w33708_ ;
	wire _w33707_ ;
	wire _w33706_ ;
	wire _w33705_ ;
	wire _w33704_ ;
	wire _w33703_ ;
	wire _w33702_ ;
	wire _w33701_ ;
	wire _w33700_ ;
	wire _w33699_ ;
	wire _w33698_ ;
	wire _w33697_ ;
	wire _w33696_ ;
	wire _w33695_ ;
	wire _w33694_ ;
	wire _w33693_ ;
	wire _w33692_ ;
	wire _w33691_ ;
	wire _w33690_ ;
	wire _w33689_ ;
	wire _w33688_ ;
	wire _w33687_ ;
	wire _w33686_ ;
	wire _w33685_ ;
	wire _w33684_ ;
	wire _w33683_ ;
	wire _w33682_ ;
	wire _w33681_ ;
	wire _w33680_ ;
	wire _w33679_ ;
	wire _w33678_ ;
	wire _w33677_ ;
	wire _w33676_ ;
	wire _w33675_ ;
	wire _w33674_ ;
	wire _w33673_ ;
	wire _w33672_ ;
	wire _w33671_ ;
	wire _w33670_ ;
	wire _w33669_ ;
	wire _w33668_ ;
	wire _w33667_ ;
	wire _w33666_ ;
	wire _w33665_ ;
	wire _w33664_ ;
	wire _w33663_ ;
	wire _w33662_ ;
	wire _w33661_ ;
	wire _w33660_ ;
	wire _w33659_ ;
	wire _w33658_ ;
	wire _w33657_ ;
	wire _w33656_ ;
	wire _w33655_ ;
	wire _w33654_ ;
	wire _w33653_ ;
	wire _w33652_ ;
	wire _w33651_ ;
	wire _w33650_ ;
	wire _w33649_ ;
	wire _w33648_ ;
	wire _w33647_ ;
	wire _w33646_ ;
	wire _w33645_ ;
	wire _w33644_ ;
	wire _w33643_ ;
	wire _w33642_ ;
	wire _w33641_ ;
	wire _w33640_ ;
	wire _w33639_ ;
	wire _w33638_ ;
	wire _w33637_ ;
	wire _w33636_ ;
	wire _w33635_ ;
	wire _w33634_ ;
	wire _w33633_ ;
	wire _w33632_ ;
	wire _w33631_ ;
	wire _w33630_ ;
	wire _w33629_ ;
	wire _w33628_ ;
	wire _w33627_ ;
	wire _w33626_ ;
	wire _w33625_ ;
	wire _w33624_ ;
	wire _w33623_ ;
	wire _w33622_ ;
	wire _w33621_ ;
	wire _w33620_ ;
	wire _w33619_ ;
	wire _w33618_ ;
	wire _w33617_ ;
	wire _w33616_ ;
	wire _w33615_ ;
	wire _w33614_ ;
	wire _w33613_ ;
	wire _w33612_ ;
	wire _w33611_ ;
	wire _w33610_ ;
	wire _w33609_ ;
	wire _w33608_ ;
	wire _w33607_ ;
	wire _w33606_ ;
	wire _w33605_ ;
	wire _w33604_ ;
	wire _w33603_ ;
	wire _w33602_ ;
	wire _w33601_ ;
	wire _w33600_ ;
	wire _w33599_ ;
	wire _w33598_ ;
	wire _w33597_ ;
	wire _w33596_ ;
	wire _w33595_ ;
	wire _w33594_ ;
	wire _w33593_ ;
	wire _w33592_ ;
	wire _w33591_ ;
	wire _w33590_ ;
	wire _w33589_ ;
	wire _w33588_ ;
	wire _w33587_ ;
	wire _w33586_ ;
	wire _w33585_ ;
	wire _w33584_ ;
	wire _w33583_ ;
	wire _w33582_ ;
	wire _w33581_ ;
	wire _w33580_ ;
	wire _w33579_ ;
	wire _w33578_ ;
	wire _w33577_ ;
	wire _w33576_ ;
	wire _w33575_ ;
	wire _w33574_ ;
	wire _w33573_ ;
	wire _w33572_ ;
	wire _w33571_ ;
	wire _w33570_ ;
	wire _w33569_ ;
	wire _w33568_ ;
	wire _w33567_ ;
	wire _w33566_ ;
	wire _w33565_ ;
	wire _w33564_ ;
	wire _w33563_ ;
	wire _w33562_ ;
	wire _w33561_ ;
	wire _w33560_ ;
	wire _w33559_ ;
	wire _w33558_ ;
	wire _w33557_ ;
	wire _w33556_ ;
	wire _w33555_ ;
	wire _w33554_ ;
	wire _w33553_ ;
	wire _w33552_ ;
	wire _w33551_ ;
	wire _w33550_ ;
	wire _w33549_ ;
	wire _w33548_ ;
	wire _w33547_ ;
	wire _w33546_ ;
	wire _w33545_ ;
	wire _w33544_ ;
	wire _w33543_ ;
	wire _w33542_ ;
	wire _w33541_ ;
	wire _w33540_ ;
	wire _w33539_ ;
	wire _w33538_ ;
	wire _w33537_ ;
	wire _w33536_ ;
	wire _w33535_ ;
	wire _w33534_ ;
	wire _w33533_ ;
	wire _w33532_ ;
	wire _w33531_ ;
	wire _w33530_ ;
	wire _w33529_ ;
	wire _w33528_ ;
	wire _w33527_ ;
	wire _w33526_ ;
	wire _w33525_ ;
	wire _w33524_ ;
	wire _w33523_ ;
	wire _w33522_ ;
	wire _w33521_ ;
	wire _w33520_ ;
	wire _w33519_ ;
	wire _w33518_ ;
	wire _w33517_ ;
	wire _w33516_ ;
	wire _w33515_ ;
	wire _w33514_ ;
	wire _w33513_ ;
	wire _w33512_ ;
	wire _w33511_ ;
	wire _w33510_ ;
	wire _w33509_ ;
	wire _w33508_ ;
	wire _w33507_ ;
	wire _w33506_ ;
	wire _w33505_ ;
	wire _w33504_ ;
	wire _w33503_ ;
	wire _w33502_ ;
	wire _w33501_ ;
	wire _w33500_ ;
	wire _w33499_ ;
	wire _w33498_ ;
	wire _w33497_ ;
	wire _w33496_ ;
	wire _w33495_ ;
	wire _w33494_ ;
	wire _w33493_ ;
	wire _w33492_ ;
	wire _w33491_ ;
	wire _w33490_ ;
	wire _w33489_ ;
	wire _w33488_ ;
	wire _w33487_ ;
	wire _w33486_ ;
	wire _w33485_ ;
	wire _w33484_ ;
	wire _w33483_ ;
	wire _w33482_ ;
	wire _w33481_ ;
	wire _w33480_ ;
	wire _w33479_ ;
	wire _w33478_ ;
	wire _w33477_ ;
	wire _w33476_ ;
	wire _w33475_ ;
	wire _w33474_ ;
	wire _w33473_ ;
	wire _w33472_ ;
	wire _w33471_ ;
	wire _w33470_ ;
	wire _w33469_ ;
	wire _w33468_ ;
	wire _w33467_ ;
	wire _w33466_ ;
	wire _w33465_ ;
	wire _w33464_ ;
	wire _w33463_ ;
	wire _w33462_ ;
	wire _w33461_ ;
	wire _w33460_ ;
	wire _w33459_ ;
	wire _w33458_ ;
	wire _w33457_ ;
	wire _w33456_ ;
	wire _w33455_ ;
	wire _w33454_ ;
	wire _w33453_ ;
	wire _w33452_ ;
	wire _w33451_ ;
	wire _w33450_ ;
	wire _w33449_ ;
	wire _w33448_ ;
	wire _w33447_ ;
	wire _w33446_ ;
	wire _w33445_ ;
	wire _w33444_ ;
	wire _w33443_ ;
	wire _w33442_ ;
	wire _w33441_ ;
	wire _w33440_ ;
	wire _w33439_ ;
	wire _w33438_ ;
	wire _w33437_ ;
	wire _w33436_ ;
	wire _w33435_ ;
	wire _w33434_ ;
	wire _w33433_ ;
	wire _w33432_ ;
	wire _w33431_ ;
	wire _w33430_ ;
	wire _w33429_ ;
	wire _w33428_ ;
	wire _w33427_ ;
	wire _w33426_ ;
	wire _w33425_ ;
	wire _w33424_ ;
	wire _w33423_ ;
	wire _w33422_ ;
	wire _w33421_ ;
	wire _w33420_ ;
	wire _w33419_ ;
	wire _w33418_ ;
	wire _w33417_ ;
	wire _w33416_ ;
	wire _w33415_ ;
	wire _w33414_ ;
	wire _w33413_ ;
	wire _w33412_ ;
	wire _w33411_ ;
	wire _w33410_ ;
	wire _w33409_ ;
	wire _w33408_ ;
	wire _w33407_ ;
	wire _w33406_ ;
	wire _w33405_ ;
	wire _w33404_ ;
	wire _w33403_ ;
	wire _w33402_ ;
	wire _w33401_ ;
	wire _w33400_ ;
	wire _w33399_ ;
	wire _w33398_ ;
	wire _w33397_ ;
	wire _w33396_ ;
	wire _w33395_ ;
	wire _w33394_ ;
	wire _w33393_ ;
	wire _w33392_ ;
	wire _w33391_ ;
	wire _w33390_ ;
	wire _w33389_ ;
	wire _w33388_ ;
	wire _w33387_ ;
	wire _w33386_ ;
	wire _w33385_ ;
	wire _w33384_ ;
	wire _w33383_ ;
	wire _w33382_ ;
	wire _w33381_ ;
	wire _w33380_ ;
	wire _w33379_ ;
	wire _w33378_ ;
	wire _w33377_ ;
	wire _w33376_ ;
	wire _w33375_ ;
	wire _w33374_ ;
	wire _w33373_ ;
	wire _w33372_ ;
	wire _w33371_ ;
	wire _w33370_ ;
	wire _w33369_ ;
	wire _w33368_ ;
	wire _w33367_ ;
	wire _w33366_ ;
	wire _w33365_ ;
	wire _w33364_ ;
	wire _w33363_ ;
	wire _w33362_ ;
	wire _w33361_ ;
	wire _w33360_ ;
	wire _w33359_ ;
	wire _w33358_ ;
	wire _w33357_ ;
	wire _w33356_ ;
	wire _w33355_ ;
	wire _w33354_ ;
	wire _w33353_ ;
	wire _w33352_ ;
	wire _w33351_ ;
	wire _w33350_ ;
	wire _w33349_ ;
	wire _w33348_ ;
	wire _w33347_ ;
	wire _w33346_ ;
	wire _w33345_ ;
	wire _w33344_ ;
	wire _w33343_ ;
	wire _w33342_ ;
	wire _w33341_ ;
	wire _w33340_ ;
	wire _w33339_ ;
	wire _w33338_ ;
	wire _w33337_ ;
	wire _w33336_ ;
	wire _w33335_ ;
	wire _w33334_ ;
	wire _w33333_ ;
	wire _w33332_ ;
	wire _w33331_ ;
	wire _w33330_ ;
	wire _w33329_ ;
	wire _w33328_ ;
	wire _w33327_ ;
	wire _w33326_ ;
	wire _w33325_ ;
	wire _w33324_ ;
	wire _w33323_ ;
	wire _w33322_ ;
	wire _w33321_ ;
	wire _w33320_ ;
	wire _w33319_ ;
	wire _w33318_ ;
	wire _w33317_ ;
	wire _w33316_ ;
	wire _w33315_ ;
	wire _w33314_ ;
	wire _w33313_ ;
	wire _w33312_ ;
	wire _w33311_ ;
	wire _w33310_ ;
	wire _w33309_ ;
	wire _w33308_ ;
	wire _w33307_ ;
	wire _w33306_ ;
	wire _w33305_ ;
	wire _w33304_ ;
	wire _w33303_ ;
	wire _w33302_ ;
	wire _w33301_ ;
	wire _w33300_ ;
	wire _w33299_ ;
	wire _w33298_ ;
	wire _w33297_ ;
	wire _w33296_ ;
	wire _w33295_ ;
	wire _w33294_ ;
	wire _w33293_ ;
	wire _w33292_ ;
	wire _w33291_ ;
	wire _w33290_ ;
	wire _w33289_ ;
	wire _w33288_ ;
	wire _w33287_ ;
	wire _w33286_ ;
	wire _w33285_ ;
	wire _w33284_ ;
	wire _w33283_ ;
	wire _w33282_ ;
	wire _w33281_ ;
	wire _w33280_ ;
	wire _w33279_ ;
	wire _w33278_ ;
	wire _w33277_ ;
	wire _w33276_ ;
	wire _w33275_ ;
	wire _w33274_ ;
	wire _w33273_ ;
	wire _w33272_ ;
	wire _w33271_ ;
	wire _w33270_ ;
	wire _w33269_ ;
	wire _w33268_ ;
	wire _w33267_ ;
	wire _w33266_ ;
	wire _w33265_ ;
	wire _w33264_ ;
	wire _w33263_ ;
	wire _w33262_ ;
	wire _w33261_ ;
	wire _w33260_ ;
	wire _w33259_ ;
	wire _w33258_ ;
	wire _w33257_ ;
	wire _w33256_ ;
	wire _w33255_ ;
	wire _w33254_ ;
	wire _w33253_ ;
	wire _w33252_ ;
	wire _w33251_ ;
	wire _w33250_ ;
	wire _w33249_ ;
	wire _w33248_ ;
	wire _w33247_ ;
	wire _w33246_ ;
	wire _w33245_ ;
	wire _w33244_ ;
	wire _w33243_ ;
	wire _w33242_ ;
	wire _w33241_ ;
	wire _w33240_ ;
	wire _w33239_ ;
	wire _w33238_ ;
	wire _w33237_ ;
	wire _w33236_ ;
	wire _w33235_ ;
	wire _w33234_ ;
	wire _w33233_ ;
	wire _w33232_ ;
	wire _w33231_ ;
	wire _w33230_ ;
	wire _w33229_ ;
	wire _w33228_ ;
	wire _w33227_ ;
	wire _w33226_ ;
	wire _w33225_ ;
	wire _w33224_ ;
	wire _w33223_ ;
	wire _w33222_ ;
	wire _w33221_ ;
	wire _w33220_ ;
	wire _w33219_ ;
	wire _w33218_ ;
	wire _w33217_ ;
	wire _w33216_ ;
	wire _w33215_ ;
	wire _w33214_ ;
	wire _w33213_ ;
	wire _w33212_ ;
	wire _w33211_ ;
	wire _w33210_ ;
	wire _w33209_ ;
	wire _w33208_ ;
	wire _w33207_ ;
	wire _w33206_ ;
	wire _w33205_ ;
	wire _w33204_ ;
	wire _w33203_ ;
	wire _w33202_ ;
	wire _w33201_ ;
	wire _w33200_ ;
	wire _w33199_ ;
	wire _w33198_ ;
	wire _w33197_ ;
	wire _w33196_ ;
	wire _w33195_ ;
	wire _w33194_ ;
	wire _w33193_ ;
	wire _w33192_ ;
	wire _w33191_ ;
	wire _w33190_ ;
	wire _w33189_ ;
	wire _w33188_ ;
	wire _w33187_ ;
	wire _w33186_ ;
	wire _w33185_ ;
	wire _w33184_ ;
	wire _w33183_ ;
	wire _w33182_ ;
	wire _w33181_ ;
	wire _w33180_ ;
	wire _w33179_ ;
	wire _w33178_ ;
	wire _w33177_ ;
	wire _w33176_ ;
	wire _w33175_ ;
	wire _w33174_ ;
	wire _w33173_ ;
	wire _w33172_ ;
	wire _w33171_ ;
	wire _w33170_ ;
	wire _w33169_ ;
	wire _w33168_ ;
	wire _w33167_ ;
	wire _w33166_ ;
	wire _w33165_ ;
	wire _w33164_ ;
	wire _w33163_ ;
	wire _w33162_ ;
	wire _w33161_ ;
	wire _w33160_ ;
	wire _w33159_ ;
	wire _w33158_ ;
	wire _w33157_ ;
	wire _w33156_ ;
	wire _w33155_ ;
	wire _w33154_ ;
	wire _w33153_ ;
	wire _w33152_ ;
	wire _w33151_ ;
	wire _w33150_ ;
	wire _w33149_ ;
	wire _w33148_ ;
	wire _w33147_ ;
	wire _w33146_ ;
	wire _w33145_ ;
	wire _w33144_ ;
	wire _w33143_ ;
	wire _w33142_ ;
	wire _w33141_ ;
	wire _w33140_ ;
	wire _w33139_ ;
	wire _w33138_ ;
	wire _w33137_ ;
	wire _w33136_ ;
	wire _w33135_ ;
	wire _w33134_ ;
	wire _w33133_ ;
	wire _w33132_ ;
	wire _w33131_ ;
	wire _w33130_ ;
	wire _w33129_ ;
	wire _w33128_ ;
	wire _w33127_ ;
	wire _w33126_ ;
	wire _w33125_ ;
	wire _w33124_ ;
	wire _w33123_ ;
	wire _w33122_ ;
	wire _w33121_ ;
	wire _w33120_ ;
	wire _w33119_ ;
	wire _w33118_ ;
	wire _w33117_ ;
	wire _w33116_ ;
	wire _w33115_ ;
	wire _w33114_ ;
	wire _w33113_ ;
	wire _w33112_ ;
	wire _w33111_ ;
	wire _w33110_ ;
	wire _w33109_ ;
	wire _w33108_ ;
	wire _w33107_ ;
	wire _w33106_ ;
	wire _w33105_ ;
	wire _w33104_ ;
	wire _w33103_ ;
	wire _w33102_ ;
	wire _w33101_ ;
	wire _w33100_ ;
	wire _w33099_ ;
	wire _w33098_ ;
	wire _w33097_ ;
	wire _w33096_ ;
	wire _w33095_ ;
	wire _w33094_ ;
	wire _w33093_ ;
	wire _w33092_ ;
	wire _w33091_ ;
	wire _w33090_ ;
	wire _w33089_ ;
	wire _w33088_ ;
	wire _w33087_ ;
	wire _w33086_ ;
	wire _w33085_ ;
	wire _w33084_ ;
	wire _w33083_ ;
	wire _w33082_ ;
	wire _w33081_ ;
	wire _w33080_ ;
	wire _w33079_ ;
	wire _w33078_ ;
	wire _w33077_ ;
	wire _w33076_ ;
	wire _w33075_ ;
	wire _w33074_ ;
	wire _w33073_ ;
	wire _w33072_ ;
	wire _w33071_ ;
	wire _w33070_ ;
	wire _w33069_ ;
	wire _w33068_ ;
	wire _w33067_ ;
	wire _w33066_ ;
	wire _w33065_ ;
	wire _w33064_ ;
	wire _w33063_ ;
	wire _w33062_ ;
	wire _w33061_ ;
	wire _w33060_ ;
	wire _w33059_ ;
	wire _w33058_ ;
	wire _w33057_ ;
	wire _w33056_ ;
	wire _w33055_ ;
	wire _w33054_ ;
	wire _w33053_ ;
	wire _w33052_ ;
	wire _w33051_ ;
	wire _w33050_ ;
	wire _w33049_ ;
	wire _w33048_ ;
	wire _w33047_ ;
	wire _w33046_ ;
	wire _w33045_ ;
	wire _w33044_ ;
	wire _w33043_ ;
	wire _w33042_ ;
	wire _w33041_ ;
	wire _w33040_ ;
	wire _w33039_ ;
	wire _w33038_ ;
	wire _w33037_ ;
	wire _w33036_ ;
	wire _w33035_ ;
	wire _w33034_ ;
	wire _w33033_ ;
	wire _w33032_ ;
	wire _w33031_ ;
	wire _w33030_ ;
	wire _w33029_ ;
	wire _w33028_ ;
	wire _w33027_ ;
	wire _w33026_ ;
	wire _w33025_ ;
	wire _w33024_ ;
	wire _w33023_ ;
	wire _w33022_ ;
	wire _w33021_ ;
	wire _w33020_ ;
	wire _w33019_ ;
	wire _w33018_ ;
	wire _w33017_ ;
	wire _w33016_ ;
	wire _w33015_ ;
	wire _w33014_ ;
	wire _w33013_ ;
	wire _w33012_ ;
	wire _w33011_ ;
	wire _w33010_ ;
	wire _w33009_ ;
	wire _w33008_ ;
	wire _w33007_ ;
	wire _w33006_ ;
	wire _w33005_ ;
	wire _w33004_ ;
	wire _w33003_ ;
	wire _w33002_ ;
	wire _w33001_ ;
	wire _w33000_ ;
	wire _w32999_ ;
	wire _w32998_ ;
	wire _w32997_ ;
	wire _w32996_ ;
	wire _w32995_ ;
	wire _w32994_ ;
	wire _w32993_ ;
	wire _w32992_ ;
	wire _w32991_ ;
	wire _w32990_ ;
	wire _w32989_ ;
	wire _w32988_ ;
	wire _w32987_ ;
	wire _w32986_ ;
	wire _w32985_ ;
	wire _w32984_ ;
	wire _w32983_ ;
	wire _w32982_ ;
	wire _w32981_ ;
	wire _w32980_ ;
	wire _w32979_ ;
	wire _w32978_ ;
	wire _w32977_ ;
	wire _w32976_ ;
	wire _w32975_ ;
	wire _w32974_ ;
	wire _w32973_ ;
	wire _w32972_ ;
	wire _w32971_ ;
	wire _w32970_ ;
	wire _w32969_ ;
	wire _w32968_ ;
	wire _w32967_ ;
	wire _w32966_ ;
	wire _w32965_ ;
	wire _w32964_ ;
	wire _w32963_ ;
	wire _w32962_ ;
	wire _w32961_ ;
	wire _w32960_ ;
	wire _w32959_ ;
	wire _w32958_ ;
	wire _w32957_ ;
	wire _w32956_ ;
	wire _w32955_ ;
	wire _w32954_ ;
	wire _w32953_ ;
	wire _w32952_ ;
	wire _w32951_ ;
	wire _w32950_ ;
	wire _w32949_ ;
	wire _w32948_ ;
	wire _w32947_ ;
	wire _w32946_ ;
	wire _w32945_ ;
	wire _w32944_ ;
	wire _w32943_ ;
	wire _w32942_ ;
	wire _w32941_ ;
	wire _w32940_ ;
	wire _w32939_ ;
	wire _w32938_ ;
	wire _w32937_ ;
	wire _w32936_ ;
	wire _w32935_ ;
	wire _w32934_ ;
	wire _w32933_ ;
	wire _w32932_ ;
	wire _w32931_ ;
	wire _w32930_ ;
	wire _w32929_ ;
	wire _w32928_ ;
	wire _w32927_ ;
	wire _w32926_ ;
	wire _w32925_ ;
	wire _w32924_ ;
	wire _w32923_ ;
	wire _w32922_ ;
	wire _w32921_ ;
	wire _w32920_ ;
	wire _w32919_ ;
	wire _w32918_ ;
	wire _w32917_ ;
	wire _w32916_ ;
	wire _w32915_ ;
	wire _w32914_ ;
	wire _w32913_ ;
	wire _w32912_ ;
	wire _w32911_ ;
	wire _w32910_ ;
	wire _w32909_ ;
	wire _w32908_ ;
	wire _w32907_ ;
	wire _w32906_ ;
	wire _w32905_ ;
	wire _w32904_ ;
	wire _w32903_ ;
	wire _w32902_ ;
	wire _w32901_ ;
	wire _w32900_ ;
	wire _w32899_ ;
	wire _w32898_ ;
	wire _w32897_ ;
	wire _w32896_ ;
	wire _w32895_ ;
	wire _w32894_ ;
	wire _w32893_ ;
	wire _w32892_ ;
	wire _w32891_ ;
	wire _w32890_ ;
	wire _w32889_ ;
	wire _w32888_ ;
	wire _w32887_ ;
	wire _w32886_ ;
	wire _w32885_ ;
	wire _w32884_ ;
	wire _w32883_ ;
	wire _w32882_ ;
	wire _w32881_ ;
	wire _w32880_ ;
	wire _w32879_ ;
	wire _w32878_ ;
	wire _w32877_ ;
	wire _w32876_ ;
	wire _w32875_ ;
	wire _w32874_ ;
	wire _w32873_ ;
	wire _w32872_ ;
	wire _w32871_ ;
	wire _w32870_ ;
	wire _w32869_ ;
	wire _w32868_ ;
	wire _w32867_ ;
	wire _w32866_ ;
	wire _w32865_ ;
	wire _w32864_ ;
	wire _w32863_ ;
	wire _w32862_ ;
	wire _w32861_ ;
	wire _w32860_ ;
	wire _w32859_ ;
	wire _w32858_ ;
	wire _w32857_ ;
	wire _w32856_ ;
	wire _w32855_ ;
	wire _w32854_ ;
	wire _w32853_ ;
	wire _w32852_ ;
	wire _w32851_ ;
	wire _w32850_ ;
	wire _w32849_ ;
	wire _w32848_ ;
	wire _w32847_ ;
	wire _w32846_ ;
	wire _w32845_ ;
	wire _w32844_ ;
	wire _w32843_ ;
	wire _w32842_ ;
	wire _w32841_ ;
	wire _w32840_ ;
	wire _w32839_ ;
	wire _w32838_ ;
	wire _w32837_ ;
	wire _w32836_ ;
	wire _w32835_ ;
	wire _w32834_ ;
	wire _w32833_ ;
	wire _w32832_ ;
	wire _w32831_ ;
	wire _w32830_ ;
	wire _w32829_ ;
	wire _w32828_ ;
	wire _w32827_ ;
	wire _w32826_ ;
	wire _w32825_ ;
	wire _w32824_ ;
	wire _w32823_ ;
	wire _w32822_ ;
	wire _w32821_ ;
	wire _w32820_ ;
	wire _w32819_ ;
	wire _w32818_ ;
	wire _w32817_ ;
	wire _w32816_ ;
	wire _w32815_ ;
	wire _w32814_ ;
	wire _w32813_ ;
	wire _w32812_ ;
	wire _w32811_ ;
	wire _w32810_ ;
	wire _w32809_ ;
	wire _w32808_ ;
	wire _w32807_ ;
	wire _w32806_ ;
	wire _w32805_ ;
	wire _w32804_ ;
	wire _w32803_ ;
	wire _w32802_ ;
	wire _w32801_ ;
	wire _w32800_ ;
	wire _w32799_ ;
	wire _w32798_ ;
	wire _w32797_ ;
	wire _w32796_ ;
	wire _w32795_ ;
	wire _w32794_ ;
	wire _w32793_ ;
	wire _w32792_ ;
	wire _w32791_ ;
	wire _w32790_ ;
	wire _w32789_ ;
	wire _w32788_ ;
	wire _w32787_ ;
	wire _w32786_ ;
	wire _w32785_ ;
	wire _w32784_ ;
	wire _w32783_ ;
	wire _w32782_ ;
	wire _w32781_ ;
	wire _w32780_ ;
	wire _w32779_ ;
	wire _w32778_ ;
	wire _w32777_ ;
	wire _w32776_ ;
	wire _w32775_ ;
	wire _w32774_ ;
	wire _w32773_ ;
	wire _w32772_ ;
	wire _w32771_ ;
	wire _w32770_ ;
	wire _w32769_ ;
	wire _w32768_ ;
	wire _w32767_ ;
	wire _w32766_ ;
	wire _w32765_ ;
	wire _w32764_ ;
	wire _w32763_ ;
	wire _w32762_ ;
	wire _w32761_ ;
	wire _w32760_ ;
	wire _w32759_ ;
	wire _w32758_ ;
	wire _w32757_ ;
	wire _w32756_ ;
	wire _w32755_ ;
	wire _w32754_ ;
	wire _w32753_ ;
	wire _w32752_ ;
	wire _w32751_ ;
	wire _w32750_ ;
	wire _w32749_ ;
	wire _w32748_ ;
	wire _w32747_ ;
	wire _w32746_ ;
	wire _w32745_ ;
	wire _w32744_ ;
	wire _w32743_ ;
	wire _w32742_ ;
	wire _w32741_ ;
	wire _w32740_ ;
	wire _w32739_ ;
	wire _w32738_ ;
	wire _w32737_ ;
	wire _w32736_ ;
	wire _w32735_ ;
	wire _w32734_ ;
	wire _w32733_ ;
	wire _w32732_ ;
	wire _w32731_ ;
	wire _w32730_ ;
	wire _w32729_ ;
	wire _w32728_ ;
	wire _w32727_ ;
	wire _w32726_ ;
	wire _w32725_ ;
	wire _w32724_ ;
	wire _w32723_ ;
	wire _w32722_ ;
	wire _w32721_ ;
	wire _w32720_ ;
	wire _w32719_ ;
	wire _w32718_ ;
	wire _w32717_ ;
	wire _w32716_ ;
	wire _w32715_ ;
	wire _w32714_ ;
	wire _w32713_ ;
	wire _w32712_ ;
	wire _w32711_ ;
	wire _w32710_ ;
	wire _w32709_ ;
	wire _w32708_ ;
	wire _w32707_ ;
	wire _w32706_ ;
	wire _w32705_ ;
	wire _w32704_ ;
	wire _w32703_ ;
	wire _w32702_ ;
	wire _w32701_ ;
	wire _w32700_ ;
	wire _w32699_ ;
	wire _w32698_ ;
	wire _w32697_ ;
	wire _w32696_ ;
	wire _w32695_ ;
	wire _w32694_ ;
	wire _w32693_ ;
	wire _w32692_ ;
	wire _w32691_ ;
	wire _w32690_ ;
	wire _w32689_ ;
	wire _w32688_ ;
	wire _w32687_ ;
	wire _w32686_ ;
	wire _w32685_ ;
	wire _w32684_ ;
	wire _w32683_ ;
	wire _w32682_ ;
	wire _w32681_ ;
	wire _w32680_ ;
	wire _w32679_ ;
	wire _w32678_ ;
	wire _w32677_ ;
	wire _w32676_ ;
	wire _w32675_ ;
	wire _w32674_ ;
	wire _w32673_ ;
	wire _w32672_ ;
	wire _w32671_ ;
	wire _w32670_ ;
	wire _w32669_ ;
	wire _w32668_ ;
	wire _w32667_ ;
	wire _w32666_ ;
	wire _w32665_ ;
	wire _w32664_ ;
	wire _w32663_ ;
	wire _w32662_ ;
	wire _w32661_ ;
	wire _w32660_ ;
	wire _w32659_ ;
	wire _w32658_ ;
	wire _w32657_ ;
	wire _w32656_ ;
	wire _w32655_ ;
	wire _w32654_ ;
	wire _w32653_ ;
	wire _w32652_ ;
	wire _w32651_ ;
	wire _w32650_ ;
	wire _w32649_ ;
	wire _w32648_ ;
	wire _w32647_ ;
	wire _w32646_ ;
	wire _w32645_ ;
	wire _w32644_ ;
	wire _w32643_ ;
	wire _w32642_ ;
	wire _w32641_ ;
	wire _w32640_ ;
	wire _w32639_ ;
	wire _w32638_ ;
	wire _w32637_ ;
	wire _w32636_ ;
	wire _w32635_ ;
	wire _w32634_ ;
	wire _w32633_ ;
	wire _w32632_ ;
	wire _w32631_ ;
	wire _w32630_ ;
	wire _w32629_ ;
	wire _w32628_ ;
	wire _w32627_ ;
	wire _w32626_ ;
	wire _w32625_ ;
	wire _w32624_ ;
	wire _w32623_ ;
	wire _w32622_ ;
	wire _w32621_ ;
	wire _w32620_ ;
	wire _w32619_ ;
	wire _w32618_ ;
	wire _w32617_ ;
	wire _w32616_ ;
	wire _w32615_ ;
	wire _w32614_ ;
	wire _w32613_ ;
	wire _w32612_ ;
	wire _w32611_ ;
	wire _w32610_ ;
	wire _w32609_ ;
	wire _w32608_ ;
	wire _w32607_ ;
	wire _w32606_ ;
	wire _w32605_ ;
	wire _w32604_ ;
	wire _w32603_ ;
	wire _w32602_ ;
	wire _w32601_ ;
	wire _w32600_ ;
	wire _w32599_ ;
	wire _w32598_ ;
	wire _w32597_ ;
	wire _w32596_ ;
	wire _w32595_ ;
	wire _w32594_ ;
	wire _w32593_ ;
	wire _w32592_ ;
	wire _w32591_ ;
	wire _w32590_ ;
	wire _w32589_ ;
	wire _w32588_ ;
	wire _w32587_ ;
	wire _w32586_ ;
	wire _w32585_ ;
	wire _w32584_ ;
	wire _w32583_ ;
	wire _w32582_ ;
	wire _w32581_ ;
	wire _w32580_ ;
	wire _w32579_ ;
	wire _w32578_ ;
	wire _w32577_ ;
	wire _w32576_ ;
	wire _w32575_ ;
	wire _w32574_ ;
	wire _w32573_ ;
	wire _w32572_ ;
	wire _w32571_ ;
	wire _w32570_ ;
	wire _w32569_ ;
	wire _w32568_ ;
	wire _w32567_ ;
	wire _w32566_ ;
	wire _w32565_ ;
	wire _w32564_ ;
	wire _w32563_ ;
	wire _w32562_ ;
	wire _w32561_ ;
	wire _w32560_ ;
	wire _w32559_ ;
	wire _w32558_ ;
	wire _w32557_ ;
	wire _w32556_ ;
	wire _w32555_ ;
	wire _w32554_ ;
	wire _w32553_ ;
	wire _w32552_ ;
	wire _w32551_ ;
	wire _w32550_ ;
	wire _w32549_ ;
	wire _w32548_ ;
	wire _w32547_ ;
	wire _w32546_ ;
	wire _w32545_ ;
	wire _w32544_ ;
	wire _w32543_ ;
	wire _w32542_ ;
	wire _w32541_ ;
	wire _w32540_ ;
	wire _w32539_ ;
	wire _w32538_ ;
	wire _w32537_ ;
	wire _w32536_ ;
	wire _w32535_ ;
	wire _w32534_ ;
	wire _w32533_ ;
	wire _w32532_ ;
	wire _w32531_ ;
	wire _w32530_ ;
	wire _w32529_ ;
	wire _w32528_ ;
	wire _w32527_ ;
	wire _w32526_ ;
	wire _w32525_ ;
	wire _w32524_ ;
	wire _w32523_ ;
	wire _w32522_ ;
	wire _w32521_ ;
	wire _w32520_ ;
	wire _w32519_ ;
	wire _w32518_ ;
	wire _w32517_ ;
	wire _w32516_ ;
	wire _w32515_ ;
	wire _w32514_ ;
	wire _w32513_ ;
	wire _w32512_ ;
	wire _w32511_ ;
	wire _w32510_ ;
	wire _w32509_ ;
	wire _w32508_ ;
	wire _w32507_ ;
	wire _w32506_ ;
	wire _w32505_ ;
	wire _w32504_ ;
	wire _w32503_ ;
	wire _w32502_ ;
	wire _w32501_ ;
	wire _w32500_ ;
	wire _w32499_ ;
	wire _w32498_ ;
	wire _w32497_ ;
	wire _w32496_ ;
	wire _w32495_ ;
	wire _w32494_ ;
	wire _w32493_ ;
	wire _w32492_ ;
	wire _w32491_ ;
	wire _w32490_ ;
	wire _w32489_ ;
	wire _w32488_ ;
	wire _w32487_ ;
	wire _w32486_ ;
	wire _w32485_ ;
	wire _w32484_ ;
	wire _w32483_ ;
	wire _w32482_ ;
	wire _w32481_ ;
	wire _w32480_ ;
	wire _w32479_ ;
	wire _w32478_ ;
	wire _w32477_ ;
	wire _w32476_ ;
	wire _w32475_ ;
	wire _w32474_ ;
	wire _w32473_ ;
	wire _w32472_ ;
	wire _w32471_ ;
	wire _w32470_ ;
	wire _w32469_ ;
	wire _w32468_ ;
	wire _w32467_ ;
	wire _w32466_ ;
	wire _w32465_ ;
	wire _w32464_ ;
	wire _w32463_ ;
	wire _w32462_ ;
	wire _w32461_ ;
	wire _w32460_ ;
	wire _w32459_ ;
	wire _w32458_ ;
	wire _w32457_ ;
	wire _w32456_ ;
	wire _w32455_ ;
	wire _w32454_ ;
	wire _w32453_ ;
	wire _w32452_ ;
	wire _w32451_ ;
	wire _w32450_ ;
	wire _w32449_ ;
	wire _w32448_ ;
	wire _w32447_ ;
	wire _w32446_ ;
	wire _w32445_ ;
	wire _w32444_ ;
	wire _w32443_ ;
	wire _w32442_ ;
	wire _w32441_ ;
	wire _w32440_ ;
	wire _w32439_ ;
	wire _w32438_ ;
	wire _w32437_ ;
	wire _w32436_ ;
	wire _w32435_ ;
	wire _w32434_ ;
	wire _w32433_ ;
	wire _w32432_ ;
	wire _w32431_ ;
	wire _w32430_ ;
	wire _w32429_ ;
	wire _w32428_ ;
	wire _w32427_ ;
	wire _w32426_ ;
	wire _w32425_ ;
	wire _w32424_ ;
	wire _w32423_ ;
	wire _w32422_ ;
	wire _w32421_ ;
	wire _w32420_ ;
	wire _w32419_ ;
	wire _w32418_ ;
	wire _w32417_ ;
	wire _w32416_ ;
	wire _w32415_ ;
	wire _w32414_ ;
	wire _w32413_ ;
	wire _w32412_ ;
	wire _w32411_ ;
	wire _w32410_ ;
	wire _w32409_ ;
	wire _w32408_ ;
	wire _w32407_ ;
	wire _w32406_ ;
	wire _w32405_ ;
	wire _w32404_ ;
	wire _w32403_ ;
	wire _w32402_ ;
	wire _w32401_ ;
	wire _w32400_ ;
	wire _w32399_ ;
	wire _w32398_ ;
	wire _w32397_ ;
	wire _w32396_ ;
	wire _w32395_ ;
	wire _w32394_ ;
	wire _w32393_ ;
	wire _w32392_ ;
	wire _w32391_ ;
	wire _w32390_ ;
	wire _w32389_ ;
	wire _w32388_ ;
	wire _w32387_ ;
	wire _w32386_ ;
	wire _w32385_ ;
	wire _w32384_ ;
	wire _w32383_ ;
	wire _w32382_ ;
	wire _w32381_ ;
	wire _w32380_ ;
	wire _w32379_ ;
	wire _w32378_ ;
	wire _w32377_ ;
	wire _w32376_ ;
	wire _w32375_ ;
	wire _w32374_ ;
	wire _w32373_ ;
	wire _w32372_ ;
	wire _w32371_ ;
	wire _w32370_ ;
	wire _w32369_ ;
	wire _w32368_ ;
	wire _w32367_ ;
	wire _w32366_ ;
	wire _w32365_ ;
	wire _w32364_ ;
	wire _w32363_ ;
	wire _w32362_ ;
	wire _w32361_ ;
	wire _w32360_ ;
	wire _w32359_ ;
	wire _w32358_ ;
	wire _w32357_ ;
	wire _w32356_ ;
	wire _w32355_ ;
	wire _w32354_ ;
	wire _w32353_ ;
	wire _w32352_ ;
	wire _w32351_ ;
	wire _w32350_ ;
	wire _w32349_ ;
	wire _w32348_ ;
	wire _w32347_ ;
	wire _w32346_ ;
	wire _w32345_ ;
	wire _w32344_ ;
	wire _w32343_ ;
	wire _w32342_ ;
	wire _w32341_ ;
	wire _w32340_ ;
	wire _w32339_ ;
	wire _w32338_ ;
	wire _w32337_ ;
	wire _w32336_ ;
	wire _w32335_ ;
	wire _w32334_ ;
	wire _w32333_ ;
	wire _w32332_ ;
	wire _w32331_ ;
	wire _w32330_ ;
	wire _w32329_ ;
	wire _w32328_ ;
	wire _w32327_ ;
	wire _w32326_ ;
	wire _w32325_ ;
	wire _w32324_ ;
	wire _w32323_ ;
	wire _w32322_ ;
	wire _w32321_ ;
	wire _w32320_ ;
	wire _w32319_ ;
	wire _w32318_ ;
	wire _w32317_ ;
	wire _w32316_ ;
	wire _w32315_ ;
	wire _w32314_ ;
	wire _w32313_ ;
	wire _w32312_ ;
	wire _w32311_ ;
	wire _w32310_ ;
	wire _w32309_ ;
	wire _w32308_ ;
	wire _w32307_ ;
	wire _w32306_ ;
	wire _w32305_ ;
	wire _w32304_ ;
	wire _w32303_ ;
	wire _w32302_ ;
	wire _w32301_ ;
	wire _w32300_ ;
	wire _w32299_ ;
	wire _w32298_ ;
	wire _w32297_ ;
	wire _w32296_ ;
	wire _w32295_ ;
	wire _w32294_ ;
	wire _w32293_ ;
	wire _w32292_ ;
	wire _w32291_ ;
	wire _w32290_ ;
	wire _w32289_ ;
	wire _w32288_ ;
	wire _w32287_ ;
	wire _w32286_ ;
	wire _w32285_ ;
	wire _w32284_ ;
	wire _w32283_ ;
	wire _w32282_ ;
	wire _w32281_ ;
	wire _w32280_ ;
	wire _w32279_ ;
	wire _w32278_ ;
	wire _w32277_ ;
	wire _w32276_ ;
	wire _w32275_ ;
	wire _w32274_ ;
	wire _w32273_ ;
	wire _w32272_ ;
	wire _w32271_ ;
	wire _w32270_ ;
	wire _w32269_ ;
	wire _w32268_ ;
	wire _w32267_ ;
	wire _w32266_ ;
	wire _w32265_ ;
	wire _w32264_ ;
	wire _w32263_ ;
	wire _w32262_ ;
	wire _w32261_ ;
	wire _w32260_ ;
	wire _w32259_ ;
	wire _w32258_ ;
	wire _w32257_ ;
	wire _w32256_ ;
	wire _w32255_ ;
	wire _w32254_ ;
	wire _w32253_ ;
	wire _w32252_ ;
	wire _w32251_ ;
	wire _w32250_ ;
	wire _w32249_ ;
	wire _w32248_ ;
	wire _w32247_ ;
	wire _w32246_ ;
	wire _w32245_ ;
	wire _w32244_ ;
	wire _w32243_ ;
	wire _w32242_ ;
	wire _w32241_ ;
	wire _w32240_ ;
	wire _w32239_ ;
	wire _w32238_ ;
	wire _w32237_ ;
	wire _w32236_ ;
	wire _w32235_ ;
	wire _w32234_ ;
	wire _w32233_ ;
	wire _w32232_ ;
	wire _w32231_ ;
	wire _w32230_ ;
	wire _w32229_ ;
	wire _w32228_ ;
	wire _w32227_ ;
	wire _w32226_ ;
	wire _w32225_ ;
	wire _w32224_ ;
	wire _w32223_ ;
	wire _w32222_ ;
	wire _w32221_ ;
	wire _w32220_ ;
	wire _w32219_ ;
	wire _w32218_ ;
	wire _w32217_ ;
	wire _w32216_ ;
	wire _w32215_ ;
	wire _w32214_ ;
	wire _w32213_ ;
	wire _w32212_ ;
	wire _w32211_ ;
	wire _w32210_ ;
	wire _w32209_ ;
	wire _w32208_ ;
	wire _w32207_ ;
	wire _w32206_ ;
	wire _w32205_ ;
	wire _w32204_ ;
	wire _w32203_ ;
	wire _w32202_ ;
	wire _w32201_ ;
	wire _w32200_ ;
	wire _w32199_ ;
	wire _w32198_ ;
	wire _w32197_ ;
	wire _w32196_ ;
	wire _w32195_ ;
	wire _w32194_ ;
	wire _w32193_ ;
	wire _w32192_ ;
	wire _w32191_ ;
	wire _w32190_ ;
	wire _w32189_ ;
	wire _w32188_ ;
	wire _w32187_ ;
	wire _w32186_ ;
	wire _w32185_ ;
	wire _w32184_ ;
	wire _w32183_ ;
	wire _w32182_ ;
	wire _w32181_ ;
	wire _w32180_ ;
	wire _w32179_ ;
	wire _w32178_ ;
	wire _w32177_ ;
	wire _w32176_ ;
	wire _w32175_ ;
	wire _w32174_ ;
	wire _w32173_ ;
	wire _w32172_ ;
	wire _w32171_ ;
	wire _w32170_ ;
	wire _w32169_ ;
	wire _w32168_ ;
	wire _w32167_ ;
	wire _w32166_ ;
	wire _w32165_ ;
	wire _w32164_ ;
	wire _w32163_ ;
	wire _w32162_ ;
	wire _w32161_ ;
	wire _w32160_ ;
	wire _w32159_ ;
	wire _w32158_ ;
	wire _w32157_ ;
	wire _w32156_ ;
	wire _w32155_ ;
	wire _w32154_ ;
	wire _w32153_ ;
	wire _w32152_ ;
	wire _w32151_ ;
	wire _w32150_ ;
	wire _w32149_ ;
	wire _w32148_ ;
	wire _w32147_ ;
	wire _w32146_ ;
	wire _w32145_ ;
	wire _w32144_ ;
	wire _w32143_ ;
	wire _w32142_ ;
	wire _w32141_ ;
	wire _w32140_ ;
	wire _w32139_ ;
	wire _w32138_ ;
	wire _w32137_ ;
	wire _w32136_ ;
	wire _w32135_ ;
	wire _w32134_ ;
	wire _w32133_ ;
	wire _w32132_ ;
	wire _w32131_ ;
	wire _w32130_ ;
	wire _w32129_ ;
	wire _w32128_ ;
	wire _w32127_ ;
	wire _w32126_ ;
	wire _w32125_ ;
	wire _w32124_ ;
	wire _w32123_ ;
	wire _w32122_ ;
	wire _w32121_ ;
	wire _w32120_ ;
	wire _w32119_ ;
	wire _w32118_ ;
	wire _w32117_ ;
	wire _w32116_ ;
	wire _w32115_ ;
	wire _w32114_ ;
	wire _w32113_ ;
	wire _w32112_ ;
	wire _w32111_ ;
	wire _w32110_ ;
	wire _w32109_ ;
	wire _w32108_ ;
	wire _w32107_ ;
	wire _w32106_ ;
	wire _w32105_ ;
	wire _w32104_ ;
	wire _w32103_ ;
	wire _w32102_ ;
	wire _w32101_ ;
	wire _w32100_ ;
	wire _w32099_ ;
	wire _w32098_ ;
	wire _w32097_ ;
	wire _w32096_ ;
	wire _w32095_ ;
	wire _w32094_ ;
	wire _w32093_ ;
	wire _w32092_ ;
	wire _w32091_ ;
	wire _w32090_ ;
	wire _w32089_ ;
	wire _w32088_ ;
	wire _w32087_ ;
	wire _w32086_ ;
	wire _w32085_ ;
	wire _w32084_ ;
	wire _w32083_ ;
	wire _w32082_ ;
	wire _w32081_ ;
	wire _w32080_ ;
	wire _w32079_ ;
	wire _w32078_ ;
	wire _w32077_ ;
	wire _w32076_ ;
	wire _w32075_ ;
	wire _w32074_ ;
	wire _w32073_ ;
	wire _w32072_ ;
	wire _w32071_ ;
	wire _w32070_ ;
	wire _w32069_ ;
	wire _w32068_ ;
	wire _w32067_ ;
	wire _w32066_ ;
	wire _w32065_ ;
	wire _w32064_ ;
	wire _w32063_ ;
	wire _w32062_ ;
	wire _w32061_ ;
	wire _w32060_ ;
	wire _w32059_ ;
	wire _w32058_ ;
	wire _w32057_ ;
	wire _w32056_ ;
	wire _w32055_ ;
	wire _w32054_ ;
	wire _w32053_ ;
	wire _w32052_ ;
	wire _w32051_ ;
	wire _w32050_ ;
	wire _w32049_ ;
	wire _w32048_ ;
	wire _w32047_ ;
	wire _w32046_ ;
	wire _w32045_ ;
	wire _w32044_ ;
	wire _w32043_ ;
	wire _w32042_ ;
	wire _w32041_ ;
	wire _w32040_ ;
	wire _w32039_ ;
	wire _w32038_ ;
	wire _w32037_ ;
	wire _w32036_ ;
	wire _w32035_ ;
	wire _w32034_ ;
	wire _w32033_ ;
	wire _w32032_ ;
	wire _w32031_ ;
	wire _w32030_ ;
	wire _w32029_ ;
	wire _w32028_ ;
	wire _w32027_ ;
	wire _w32026_ ;
	wire _w32025_ ;
	wire _w32024_ ;
	wire _w32023_ ;
	wire _w32022_ ;
	wire _w32021_ ;
	wire _w32020_ ;
	wire _w32019_ ;
	wire _w32018_ ;
	wire _w32017_ ;
	wire _w32016_ ;
	wire _w32015_ ;
	wire _w32014_ ;
	wire _w32013_ ;
	wire _w32012_ ;
	wire _w32011_ ;
	wire _w32010_ ;
	wire _w32009_ ;
	wire _w32008_ ;
	wire _w32007_ ;
	wire _w32006_ ;
	wire _w32005_ ;
	wire _w32004_ ;
	wire _w32003_ ;
	wire _w32002_ ;
	wire _w32001_ ;
	wire _w32000_ ;
	wire _w31999_ ;
	wire _w31998_ ;
	wire _w31997_ ;
	wire _w31996_ ;
	wire _w31995_ ;
	wire _w31994_ ;
	wire _w31993_ ;
	wire _w31992_ ;
	wire _w31991_ ;
	wire _w31990_ ;
	wire _w31989_ ;
	wire _w31988_ ;
	wire _w31987_ ;
	wire _w31986_ ;
	wire _w31985_ ;
	wire _w31984_ ;
	wire _w31983_ ;
	wire _w31982_ ;
	wire _w31981_ ;
	wire _w31980_ ;
	wire _w31979_ ;
	wire _w31978_ ;
	wire _w31977_ ;
	wire _w31976_ ;
	wire _w31975_ ;
	wire _w31974_ ;
	wire _w31973_ ;
	wire _w31972_ ;
	wire _w31971_ ;
	wire _w31970_ ;
	wire _w31969_ ;
	wire _w31968_ ;
	wire _w31967_ ;
	wire _w31966_ ;
	wire _w31965_ ;
	wire _w31964_ ;
	wire _w31963_ ;
	wire _w31962_ ;
	wire _w31961_ ;
	wire _w31960_ ;
	wire _w31959_ ;
	wire _w31958_ ;
	wire _w31957_ ;
	wire _w31956_ ;
	wire _w31955_ ;
	wire _w31954_ ;
	wire _w31953_ ;
	wire _w31952_ ;
	wire _w31951_ ;
	wire _w31950_ ;
	wire _w31949_ ;
	wire _w31948_ ;
	wire _w31947_ ;
	wire _w31946_ ;
	wire _w31945_ ;
	wire _w31944_ ;
	wire _w31943_ ;
	wire _w31942_ ;
	wire _w31941_ ;
	wire _w31940_ ;
	wire _w31939_ ;
	wire _w31938_ ;
	wire _w31937_ ;
	wire _w31936_ ;
	wire _w31935_ ;
	wire _w31934_ ;
	wire _w31933_ ;
	wire _w31932_ ;
	wire _w31931_ ;
	wire _w31930_ ;
	wire _w31929_ ;
	wire _w31928_ ;
	wire _w31927_ ;
	wire _w31926_ ;
	wire _w31925_ ;
	wire _w31924_ ;
	wire _w31923_ ;
	wire _w31922_ ;
	wire _w31921_ ;
	wire _w31920_ ;
	wire _w31919_ ;
	wire _w31918_ ;
	wire _w31917_ ;
	wire _w31916_ ;
	wire _w31915_ ;
	wire _w31914_ ;
	wire _w31913_ ;
	wire _w31912_ ;
	wire _w31911_ ;
	wire _w31910_ ;
	wire _w31909_ ;
	wire _w31908_ ;
	wire _w31907_ ;
	wire _w31906_ ;
	wire _w31905_ ;
	wire _w31904_ ;
	wire _w31903_ ;
	wire _w31902_ ;
	wire _w31901_ ;
	wire _w31900_ ;
	wire _w31899_ ;
	wire _w31898_ ;
	wire _w31897_ ;
	wire _w31896_ ;
	wire _w31895_ ;
	wire _w31894_ ;
	wire _w31893_ ;
	wire _w31892_ ;
	wire _w31891_ ;
	wire _w31890_ ;
	wire _w31889_ ;
	wire _w31888_ ;
	wire _w31887_ ;
	wire _w31886_ ;
	wire _w31885_ ;
	wire _w31884_ ;
	wire _w31883_ ;
	wire _w31882_ ;
	wire _w31881_ ;
	wire _w31880_ ;
	wire _w31879_ ;
	wire _w31878_ ;
	wire _w31877_ ;
	wire _w31876_ ;
	wire _w31875_ ;
	wire _w31874_ ;
	wire _w31873_ ;
	wire _w31872_ ;
	wire _w31871_ ;
	wire _w31870_ ;
	wire _w31869_ ;
	wire _w31868_ ;
	wire _w31867_ ;
	wire _w31866_ ;
	wire _w31865_ ;
	wire _w31864_ ;
	wire _w31863_ ;
	wire _w31862_ ;
	wire _w31861_ ;
	wire _w31860_ ;
	wire _w31859_ ;
	wire _w31858_ ;
	wire _w31857_ ;
	wire _w31856_ ;
	wire _w31855_ ;
	wire _w31854_ ;
	wire _w31853_ ;
	wire _w31852_ ;
	wire _w31851_ ;
	wire _w31850_ ;
	wire _w31849_ ;
	wire _w31848_ ;
	wire _w31847_ ;
	wire _w31846_ ;
	wire _w31845_ ;
	wire _w31844_ ;
	wire _w31843_ ;
	wire _w31842_ ;
	wire _w31841_ ;
	wire _w31840_ ;
	wire _w31839_ ;
	wire _w31838_ ;
	wire _w31837_ ;
	wire _w31836_ ;
	wire _w31835_ ;
	wire _w31834_ ;
	wire _w31833_ ;
	wire _w31832_ ;
	wire _w31831_ ;
	wire _w31830_ ;
	wire _w31829_ ;
	wire _w31828_ ;
	wire _w31827_ ;
	wire _w31826_ ;
	wire _w31825_ ;
	wire _w31824_ ;
	wire _w31823_ ;
	wire _w31822_ ;
	wire _w31821_ ;
	wire _w31820_ ;
	wire _w31819_ ;
	wire _w31818_ ;
	wire _w31817_ ;
	wire _w31816_ ;
	wire _w31815_ ;
	wire _w31814_ ;
	wire _w31813_ ;
	wire _w31812_ ;
	wire _w31811_ ;
	wire _w31810_ ;
	wire _w31809_ ;
	wire _w31808_ ;
	wire _w31807_ ;
	wire _w31806_ ;
	wire _w31805_ ;
	wire _w31804_ ;
	wire _w31803_ ;
	wire _w31802_ ;
	wire _w31801_ ;
	wire _w31800_ ;
	wire _w31799_ ;
	wire _w31798_ ;
	wire _w31797_ ;
	wire _w31796_ ;
	wire _w31795_ ;
	wire _w31794_ ;
	wire _w31793_ ;
	wire _w31792_ ;
	wire _w31791_ ;
	wire _w31790_ ;
	wire _w31789_ ;
	wire _w31788_ ;
	wire _w31787_ ;
	wire _w31786_ ;
	wire _w31785_ ;
	wire _w31784_ ;
	wire _w31783_ ;
	wire _w31782_ ;
	wire _w31781_ ;
	wire _w31780_ ;
	wire _w31779_ ;
	wire _w31778_ ;
	wire _w31777_ ;
	wire _w31776_ ;
	wire _w31775_ ;
	wire _w31774_ ;
	wire _w31773_ ;
	wire _w31772_ ;
	wire _w31771_ ;
	wire _w31770_ ;
	wire _w31769_ ;
	wire _w31768_ ;
	wire _w31767_ ;
	wire _w31766_ ;
	wire _w31765_ ;
	wire _w31764_ ;
	wire _w31763_ ;
	wire _w31762_ ;
	wire _w31761_ ;
	wire _w31760_ ;
	wire _w31759_ ;
	wire _w31758_ ;
	wire _w31757_ ;
	wire _w31756_ ;
	wire _w31755_ ;
	wire _w31754_ ;
	wire _w31753_ ;
	wire _w31752_ ;
	wire _w31751_ ;
	wire _w31750_ ;
	wire _w31749_ ;
	wire _w31748_ ;
	wire _w31747_ ;
	wire _w31746_ ;
	wire _w31745_ ;
	wire _w31744_ ;
	wire _w31743_ ;
	wire _w31742_ ;
	wire _w31741_ ;
	wire _w31740_ ;
	wire _w31739_ ;
	wire _w31738_ ;
	wire _w31737_ ;
	wire _w31736_ ;
	wire _w31735_ ;
	wire _w31734_ ;
	wire _w31733_ ;
	wire _w31732_ ;
	wire _w31731_ ;
	wire _w31730_ ;
	wire _w31729_ ;
	wire _w31728_ ;
	wire _w31727_ ;
	wire _w31726_ ;
	wire _w31725_ ;
	wire _w31724_ ;
	wire _w31723_ ;
	wire _w31722_ ;
	wire _w31721_ ;
	wire _w31720_ ;
	wire _w31719_ ;
	wire _w31718_ ;
	wire _w31717_ ;
	wire _w31716_ ;
	wire _w31715_ ;
	wire _w31714_ ;
	wire _w31713_ ;
	wire _w31712_ ;
	wire _w31711_ ;
	wire _w31710_ ;
	wire _w31709_ ;
	wire _w31708_ ;
	wire _w31707_ ;
	wire _w31706_ ;
	wire _w31705_ ;
	wire _w31704_ ;
	wire _w31703_ ;
	wire _w31702_ ;
	wire _w31701_ ;
	wire _w31700_ ;
	wire _w31699_ ;
	wire _w31698_ ;
	wire _w31697_ ;
	wire _w31696_ ;
	wire _w31695_ ;
	wire _w31694_ ;
	wire _w31693_ ;
	wire _w31692_ ;
	wire _w31691_ ;
	wire _w31690_ ;
	wire _w31689_ ;
	wire _w31688_ ;
	wire _w31687_ ;
	wire _w31686_ ;
	wire _w31685_ ;
	wire _w31684_ ;
	wire _w31683_ ;
	wire _w31682_ ;
	wire _w31681_ ;
	wire _w31680_ ;
	wire _w31679_ ;
	wire _w31678_ ;
	wire _w31677_ ;
	wire _w31676_ ;
	wire _w31675_ ;
	wire _w31674_ ;
	wire _w31673_ ;
	wire _w31672_ ;
	wire _w31671_ ;
	wire _w31670_ ;
	wire _w31669_ ;
	wire _w31668_ ;
	wire _w31667_ ;
	wire _w31666_ ;
	wire _w31665_ ;
	wire _w31664_ ;
	wire _w31663_ ;
	wire _w31662_ ;
	wire _w31661_ ;
	wire _w31660_ ;
	wire _w31659_ ;
	wire _w31658_ ;
	wire _w31657_ ;
	wire _w31656_ ;
	wire _w31655_ ;
	wire _w31654_ ;
	wire _w31653_ ;
	wire _w31652_ ;
	wire _w31651_ ;
	wire _w31650_ ;
	wire _w31649_ ;
	wire _w31648_ ;
	wire _w31647_ ;
	wire _w31646_ ;
	wire _w31645_ ;
	wire _w31644_ ;
	wire _w31643_ ;
	wire _w31642_ ;
	wire _w31641_ ;
	wire _w31640_ ;
	wire _w31639_ ;
	wire _w31638_ ;
	wire _w31637_ ;
	wire _w31636_ ;
	wire _w31635_ ;
	wire _w31634_ ;
	wire _w31633_ ;
	wire _w31632_ ;
	wire _w31631_ ;
	wire _w31630_ ;
	wire _w31629_ ;
	wire _w31628_ ;
	wire _w31627_ ;
	wire _w31626_ ;
	wire _w31625_ ;
	wire _w31624_ ;
	wire _w31623_ ;
	wire _w31622_ ;
	wire _w31621_ ;
	wire _w31620_ ;
	wire _w31619_ ;
	wire _w31618_ ;
	wire _w31617_ ;
	wire _w31616_ ;
	wire _w31615_ ;
	wire _w31614_ ;
	wire _w31613_ ;
	wire _w31612_ ;
	wire _w31611_ ;
	wire _w31610_ ;
	wire _w31609_ ;
	wire _w31608_ ;
	wire _w31607_ ;
	wire _w31606_ ;
	wire _w31605_ ;
	wire _w31604_ ;
	wire _w31603_ ;
	wire _w31602_ ;
	wire _w31601_ ;
	wire _w31600_ ;
	wire _w31599_ ;
	wire _w31598_ ;
	wire _w31597_ ;
	wire _w31596_ ;
	wire _w31595_ ;
	wire _w31594_ ;
	wire _w31593_ ;
	wire _w31592_ ;
	wire _w31591_ ;
	wire _w31590_ ;
	wire _w31589_ ;
	wire _w31588_ ;
	wire _w31587_ ;
	wire _w31586_ ;
	wire _w31585_ ;
	wire _w31584_ ;
	wire _w31583_ ;
	wire _w31582_ ;
	wire _w31581_ ;
	wire _w31580_ ;
	wire _w31579_ ;
	wire _w31578_ ;
	wire _w31577_ ;
	wire _w31576_ ;
	wire _w31575_ ;
	wire _w31574_ ;
	wire _w31573_ ;
	wire _w31572_ ;
	wire _w31571_ ;
	wire _w31570_ ;
	wire _w31569_ ;
	wire _w31568_ ;
	wire _w31567_ ;
	wire _w31566_ ;
	wire _w31565_ ;
	wire _w31564_ ;
	wire _w31563_ ;
	wire _w31562_ ;
	wire _w31561_ ;
	wire _w31560_ ;
	wire _w31559_ ;
	wire _w31558_ ;
	wire _w31557_ ;
	wire _w31556_ ;
	wire _w31555_ ;
	wire _w31554_ ;
	wire _w31553_ ;
	wire _w31552_ ;
	wire _w31551_ ;
	wire _w31550_ ;
	wire _w31549_ ;
	wire _w31548_ ;
	wire _w31547_ ;
	wire _w31546_ ;
	wire _w31545_ ;
	wire _w31544_ ;
	wire _w31543_ ;
	wire _w31542_ ;
	wire _w31541_ ;
	wire _w31540_ ;
	wire _w31539_ ;
	wire _w31538_ ;
	wire _w31537_ ;
	wire _w31536_ ;
	wire _w31535_ ;
	wire _w31534_ ;
	wire _w31533_ ;
	wire _w31532_ ;
	wire _w31531_ ;
	wire _w31530_ ;
	wire _w31529_ ;
	wire _w31528_ ;
	wire _w31527_ ;
	wire _w31526_ ;
	wire _w31525_ ;
	wire _w31524_ ;
	wire _w31523_ ;
	wire _w31522_ ;
	wire _w31521_ ;
	wire _w31520_ ;
	wire _w31519_ ;
	wire _w31518_ ;
	wire _w31517_ ;
	wire _w31516_ ;
	wire _w31515_ ;
	wire _w31514_ ;
	wire _w31513_ ;
	wire _w31512_ ;
	wire _w31511_ ;
	wire _w31510_ ;
	wire _w31509_ ;
	wire _w31508_ ;
	wire _w31507_ ;
	wire _w31506_ ;
	wire _w31505_ ;
	wire _w31504_ ;
	wire _w31503_ ;
	wire _w31502_ ;
	wire _w31501_ ;
	wire _w31500_ ;
	wire _w31499_ ;
	wire _w31498_ ;
	wire _w31497_ ;
	wire _w31496_ ;
	wire _w31495_ ;
	wire _w31494_ ;
	wire _w31493_ ;
	wire _w31492_ ;
	wire _w31491_ ;
	wire _w31490_ ;
	wire _w31489_ ;
	wire _w31488_ ;
	wire _w31487_ ;
	wire _w31486_ ;
	wire _w31485_ ;
	wire _w31484_ ;
	wire _w31483_ ;
	wire _w31482_ ;
	wire _w31481_ ;
	wire _w31480_ ;
	wire _w31479_ ;
	wire _w31478_ ;
	wire _w31477_ ;
	wire _w31476_ ;
	wire _w31475_ ;
	wire _w31474_ ;
	wire _w31473_ ;
	wire _w31472_ ;
	wire _w31471_ ;
	wire _w31470_ ;
	wire _w31469_ ;
	wire _w31468_ ;
	wire _w31467_ ;
	wire _w31466_ ;
	wire _w31465_ ;
	wire _w31464_ ;
	wire _w31463_ ;
	wire _w31462_ ;
	wire _w31461_ ;
	wire _w31460_ ;
	wire _w31459_ ;
	wire _w31458_ ;
	wire _w31457_ ;
	wire _w31456_ ;
	wire _w31455_ ;
	wire _w31454_ ;
	wire _w31453_ ;
	wire _w31452_ ;
	wire _w31451_ ;
	wire _w31450_ ;
	wire _w31449_ ;
	wire _w31448_ ;
	wire _w31447_ ;
	wire _w31446_ ;
	wire _w31445_ ;
	wire _w31444_ ;
	wire _w31443_ ;
	wire _w31442_ ;
	wire _w31441_ ;
	wire _w31440_ ;
	wire _w31439_ ;
	wire _w31438_ ;
	wire _w31437_ ;
	wire _w31436_ ;
	wire _w31435_ ;
	wire _w31434_ ;
	wire _w31433_ ;
	wire _w31432_ ;
	wire _w31431_ ;
	wire _w31430_ ;
	wire _w31429_ ;
	wire _w31428_ ;
	wire _w31427_ ;
	wire _w31426_ ;
	wire _w31425_ ;
	wire _w31424_ ;
	wire _w31423_ ;
	wire _w31422_ ;
	wire _w31421_ ;
	wire _w31420_ ;
	wire _w31419_ ;
	wire _w31418_ ;
	wire _w31417_ ;
	wire _w31416_ ;
	wire _w31415_ ;
	wire _w31414_ ;
	wire _w31413_ ;
	wire _w31412_ ;
	wire _w31411_ ;
	wire _w31410_ ;
	wire _w31409_ ;
	wire _w31408_ ;
	wire _w31407_ ;
	wire _w31406_ ;
	wire _w31405_ ;
	wire _w31404_ ;
	wire _w31403_ ;
	wire _w31402_ ;
	wire _w31401_ ;
	wire _w31400_ ;
	wire _w31399_ ;
	wire _w31398_ ;
	wire _w31397_ ;
	wire _w31396_ ;
	wire _w31395_ ;
	wire _w31394_ ;
	wire _w31393_ ;
	wire _w31392_ ;
	wire _w31391_ ;
	wire _w31390_ ;
	wire _w31389_ ;
	wire _w31388_ ;
	wire _w31387_ ;
	wire _w31386_ ;
	wire _w31385_ ;
	wire _w31384_ ;
	wire _w31383_ ;
	wire _w31382_ ;
	wire _w31381_ ;
	wire _w31380_ ;
	wire _w31379_ ;
	wire _w31378_ ;
	wire _w31377_ ;
	wire _w31376_ ;
	wire _w31375_ ;
	wire _w31374_ ;
	wire _w31373_ ;
	wire _w31372_ ;
	wire _w31371_ ;
	wire _w31370_ ;
	wire _w31369_ ;
	wire _w31368_ ;
	wire _w31367_ ;
	wire _w31366_ ;
	wire _w31365_ ;
	wire _w31364_ ;
	wire _w31363_ ;
	wire _w31362_ ;
	wire _w31361_ ;
	wire _w31360_ ;
	wire _w31359_ ;
	wire _w31358_ ;
	wire _w31357_ ;
	wire _w31356_ ;
	wire _w31355_ ;
	wire _w31354_ ;
	wire _w31353_ ;
	wire _w31352_ ;
	wire _w31351_ ;
	wire _w31350_ ;
	wire _w31349_ ;
	wire _w31348_ ;
	wire _w31347_ ;
	wire _w31346_ ;
	wire _w31345_ ;
	wire _w31344_ ;
	wire _w31343_ ;
	wire _w31342_ ;
	wire _w31341_ ;
	wire _w31340_ ;
	wire _w31339_ ;
	wire _w31338_ ;
	wire _w31337_ ;
	wire _w31336_ ;
	wire _w31335_ ;
	wire _w31334_ ;
	wire _w31333_ ;
	wire _w31332_ ;
	wire _w31331_ ;
	wire _w31330_ ;
	wire _w31329_ ;
	wire _w31328_ ;
	wire _w31327_ ;
	wire _w31326_ ;
	wire _w31325_ ;
	wire _w31324_ ;
	wire _w31323_ ;
	wire _w31322_ ;
	wire _w31321_ ;
	wire _w31320_ ;
	wire _w31319_ ;
	wire _w31318_ ;
	wire _w31317_ ;
	wire _w31316_ ;
	wire _w31315_ ;
	wire _w31314_ ;
	wire _w31313_ ;
	wire _w31312_ ;
	wire _w31311_ ;
	wire _w31310_ ;
	wire _w31309_ ;
	wire _w31308_ ;
	wire _w31307_ ;
	wire _w31306_ ;
	wire _w31305_ ;
	wire _w31304_ ;
	wire _w31303_ ;
	wire _w31302_ ;
	wire _w31301_ ;
	wire _w31300_ ;
	wire _w31299_ ;
	wire _w31298_ ;
	wire _w31297_ ;
	wire _w31296_ ;
	wire _w31295_ ;
	wire _w31294_ ;
	wire _w31293_ ;
	wire _w31292_ ;
	wire _w31291_ ;
	wire _w31290_ ;
	wire _w31289_ ;
	wire _w31288_ ;
	wire _w31287_ ;
	wire _w31286_ ;
	wire _w31285_ ;
	wire _w31284_ ;
	wire _w31283_ ;
	wire _w31282_ ;
	wire _w31281_ ;
	wire _w31280_ ;
	wire _w31279_ ;
	wire _w31278_ ;
	wire _w31277_ ;
	wire _w31276_ ;
	wire _w31275_ ;
	wire _w31274_ ;
	wire _w31273_ ;
	wire _w31272_ ;
	wire _w31271_ ;
	wire _w31270_ ;
	wire _w31269_ ;
	wire _w31268_ ;
	wire _w31267_ ;
	wire _w31266_ ;
	wire _w31265_ ;
	wire _w20784_ ;
	wire _w20783_ ;
	wire _w20782_ ;
	wire _w20781_ ;
	wire _w20780_ ;
	wire _w20779_ ;
	wire _w20778_ ;
	wire _w20777_ ;
	wire _w20776_ ;
	wire _w20775_ ;
	wire _w20774_ ;
	wire _w20773_ ;
	wire _w20772_ ;
	wire _w20771_ ;
	wire _w20770_ ;
	wire _w20769_ ;
	wire _w20768_ ;
	wire _w20767_ ;
	wire _w20766_ ;
	wire _w20765_ ;
	wire _w20764_ ;
	wire _w20763_ ;
	wire _w20762_ ;
	wire _w20761_ ;
	wire _w20760_ ;
	wire _w20759_ ;
	wire _w20758_ ;
	wire _w20757_ ;
	wire _w20756_ ;
	wire _w20755_ ;
	wire _w20754_ ;
	wire _w20753_ ;
	wire _w20752_ ;
	wire _w20751_ ;
	wire _w20750_ ;
	wire _w20749_ ;
	wire _w20748_ ;
	wire _w20747_ ;
	wire _w20746_ ;
	wire _w20745_ ;
	wire _w20744_ ;
	wire _w20743_ ;
	wire _w20742_ ;
	wire _w20741_ ;
	wire _w20740_ ;
	wire _w20739_ ;
	wire _w20738_ ;
	wire _w20737_ ;
	wire _w20736_ ;
	wire _w20735_ ;
	wire _w20734_ ;
	wire _w20733_ ;
	wire _w20732_ ;
	wire _w20731_ ;
	wire _w20730_ ;
	wire _w20729_ ;
	wire _w20728_ ;
	wire _w20727_ ;
	wire _w20726_ ;
	wire _w20725_ ;
	wire _w20724_ ;
	wire _w20723_ ;
	wire _w20722_ ;
	wire _w20721_ ;
	wire _w20720_ ;
	wire _w20719_ ;
	wire _w20718_ ;
	wire _w20717_ ;
	wire _w20716_ ;
	wire _w20715_ ;
	wire _w20714_ ;
	wire _w20713_ ;
	wire _w20712_ ;
	wire _w20711_ ;
	wire _w20710_ ;
	wire _w20709_ ;
	wire _w20708_ ;
	wire _w20707_ ;
	wire _w20706_ ;
	wire _w20705_ ;
	wire _w20704_ ;
	wire _w20703_ ;
	wire _w20702_ ;
	wire _w20701_ ;
	wire _w20700_ ;
	wire _w20699_ ;
	wire _w20698_ ;
	wire _w20697_ ;
	wire _w20696_ ;
	wire _w20695_ ;
	wire _w20694_ ;
	wire _w20693_ ;
	wire _w20692_ ;
	wire _w20691_ ;
	wire _w20690_ ;
	wire _w20689_ ;
	wire _w20688_ ;
	wire _w20687_ ;
	wire _w20686_ ;
	wire _w20685_ ;
	wire _w20684_ ;
	wire _w20683_ ;
	wire _w20682_ ;
	wire _w20681_ ;
	wire _w20680_ ;
	wire _w20679_ ;
	wire _w20678_ ;
	wire _w20677_ ;
	wire _w20676_ ;
	wire _w20675_ ;
	wire _w20674_ ;
	wire _w20673_ ;
	wire _w20672_ ;
	wire _w20671_ ;
	wire _w20670_ ;
	wire _w20669_ ;
	wire _w20668_ ;
	wire _w20667_ ;
	wire _w20666_ ;
	wire _w20665_ ;
	wire _w20664_ ;
	wire _w20663_ ;
	wire _w20662_ ;
	wire _w20661_ ;
	wire _w20660_ ;
	wire _w20659_ ;
	wire _w20658_ ;
	wire _w20657_ ;
	wire _w20656_ ;
	wire _w20655_ ;
	wire _w20654_ ;
	wire _w20653_ ;
	wire _w20652_ ;
	wire _w20651_ ;
	wire _w20650_ ;
	wire _w20649_ ;
	wire _w20648_ ;
	wire _w20647_ ;
	wire _w20646_ ;
	wire _w20645_ ;
	wire _w20644_ ;
	wire _w20643_ ;
	wire _w20642_ ;
	wire _w20641_ ;
	wire _w20640_ ;
	wire _w20639_ ;
	wire _w20638_ ;
	wire _w20637_ ;
	wire _w20636_ ;
	wire _w20635_ ;
	wire _w20634_ ;
	wire _w20633_ ;
	wire _w20632_ ;
	wire _w20631_ ;
	wire _w20630_ ;
	wire _w20629_ ;
	wire _w20628_ ;
	wire _w20627_ ;
	wire _w20626_ ;
	wire _w20625_ ;
	wire _w20624_ ;
	wire _w20623_ ;
	wire _w20622_ ;
	wire _w20621_ ;
	wire _w20620_ ;
	wire _w20619_ ;
	wire _w20618_ ;
	wire _w20617_ ;
	wire _w20616_ ;
	wire _w20615_ ;
	wire _w20614_ ;
	wire _w20613_ ;
	wire _w20612_ ;
	wire _w20611_ ;
	wire _w20610_ ;
	wire _w20609_ ;
	wire _w20608_ ;
	wire _w20607_ ;
	wire _w20606_ ;
	wire _w20605_ ;
	wire _w20604_ ;
	wire _w20603_ ;
	wire _w20602_ ;
	wire _w20601_ ;
	wire _w20600_ ;
	wire _w20599_ ;
	wire _w20598_ ;
	wire _w20597_ ;
	wire _w20596_ ;
	wire _w20595_ ;
	wire _w20594_ ;
	wire _w20593_ ;
	wire _w20592_ ;
	wire _w20591_ ;
	wire _w20590_ ;
	wire _w20589_ ;
	wire _w20588_ ;
	wire _w20587_ ;
	wire _w20586_ ;
	wire _w20585_ ;
	wire _w20584_ ;
	wire _w20583_ ;
	wire _w20582_ ;
	wire _w20581_ ;
	wire _w20580_ ;
	wire _w20579_ ;
	wire _w20578_ ;
	wire _w20577_ ;
	wire _w20576_ ;
	wire _w20575_ ;
	wire _w20574_ ;
	wire _w20573_ ;
	wire _w20572_ ;
	wire _w20571_ ;
	wire _w20570_ ;
	wire _w20569_ ;
	wire _w20568_ ;
	wire _w20567_ ;
	wire _w20566_ ;
	wire _w20565_ ;
	wire _w20564_ ;
	wire _w20563_ ;
	wire _w20562_ ;
	wire _w20561_ ;
	wire _w20560_ ;
	wire _w20559_ ;
	wire _w20558_ ;
	wire _w20557_ ;
	wire _w20556_ ;
	wire _w20555_ ;
	wire _w20554_ ;
	wire _w20553_ ;
	wire _w20552_ ;
	wire _w20551_ ;
	wire _w20550_ ;
	wire _w20549_ ;
	wire _w20548_ ;
	wire _w20547_ ;
	wire _w20546_ ;
	wire _w20545_ ;
	wire _w20544_ ;
	wire _w20543_ ;
	wire _w20542_ ;
	wire _w20541_ ;
	wire _w20540_ ;
	wire _w20539_ ;
	wire _w20538_ ;
	wire _w20537_ ;
	wire _w20536_ ;
	wire _w20535_ ;
	wire _w20534_ ;
	wire _w20533_ ;
	wire _w20532_ ;
	wire _w20531_ ;
	wire _w20530_ ;
	wire _w20529_ ;
	wire _w20528_ ;
	wire _w20527_ ;
	wire _w20526_ ;
	wire _w20525_ ;
	wire _w20524_ ;
	wire _w20523_ ;
	wire _w20522_ ;
	wire _w20521_ ;
	wire _w20520_ ;
	wire _w20519_ ;
	wire _w20518_ ;
	wire _w20517_ ;
	wire _w20516_ ;
	wire _w20515_ ;
	wire _w20514_ ;
	wire _w20513_ ;
	wire _w20512_ ;
	wire _w20511_ ;
	wire _w20510_ ;
	wire _w20509_ ;
	wire _w20508_ ;
	wire _w20507_ ;
	wire _w20506_ ;
	wire _w20505_ ;
	wire _w20504_ ;
	wire _w20503_ ;
	wire _w20502_ ;
	wire _w20501_ ;
	wire _w20500_ ;
	wire _w20499_ ;
	wire _w20498_ ;
	wire _w20497_ ;
	wire _w20496_ ;
	wire _w20495_ ;
	wire _w20494_ ;
	wire _w20493_ ;
	wire _w20492_ ;
	wire _w20491_ ;
	wire _w20490_ ;
	wire _w20489_ ;
	wire _w20488_ ;
	wire _w20487_ ;
	wire _w20486_ ;
	wire _w20485_ ;
	wire _w20484_ ;
	wire _w20483_ ;
	wire _w20482_ ;
	wire _w20481_ ;
	wire _w20480_ ;
	wire _w20479_ ;
	wire _w20478_ ;
	wire _w20477_ ;
	wire _w20476_ ;
	wire _w20475_ ;
	wire _w20474_ ;
	wire _w20473_ ;
	wire _w20472_ ;
	wire _w20471_ ;
	wire _w20470_ ;
	wire _w20469_ ;
	wire _w20468_ ;
	wire _w20467_ ;
	wire _w20466_ ;
	wire _w20465_ ;
	wire _w20464_ ;
	wire _w20463_ ;
	wire _w20462_ ;
	wire _w20461_ ;
	wire _w20460_ ;
	wire _w20459_ ;
	wire _w20458_ ;
	wire _w20457_ ;
	wire _w20456_ ;
	wire _w20455_ ;
	wire _w20454_ ;
	wire _w20453_ ;
	wire _w20452_ ;
	wire _w20451_ ;
	wire _w20450_ ;
	wire _w20449_ ;
	wire _w20448_ ;
	wire _w20447_ ;
	wire _w20446_ ;
	wire _w20445_ ;
	wire _w20444_ ;
	wire _w20443_ ;
	wire _w20442_ ;
	wire _w20441_ ;
	wire _w20440_ ;
	wire _w20439_ ;
	wire _w20438_ ;
	wire _w20437_ ;
	wire _w20436_ ;
	wire _w20435_ ;
	wire _w20434_ ;
	wire _w20433_ ;
	wire _w20432_ ;
	wire _w20431_ ;
	wire _w20430_ ;
	wire _w20429_ ;
	wire _w20428_ ;
	wire _w20427_ ;
	wire _w20426_ ;
	wire _w20425_ ;
	wire _w20424_ ;
	wire _w20423_ ;
	wire _w20422_ ;
	wire _w20421_ ;
	wire _w20420_ ;
	wire _w20419_ ;
	wire _w20418_ ;
	wire _w20417_ ;
	wire _w20416_ ;
	wire _w20415_ ;
	wire _w20414_ ;
	wire _w20413_ ;
	wire _w20412_ ;
	wire _w20411_ ;
	wire _w20410_ ;
	wire _w20409_ ;
	wire _w20408_ ;
	wire _w20407_ ;
	wire _w20406_ ;
	wire _w20405_ ;
	wire _w20404_ ;
	wire _w20403_ ;
	wire _w20402_ ;
	wire _w20401_ ;
	wire _w20400_ ;
	wire _w20399_ ;
	wire _w20398_ ;
	wire _w20397_ ;
	wire _w20396_ ;
	wire _w20395_ ;
	wire _w20394_ ;
	wire _w20393_ ;
	wire _w20392_ ;
	wire _w20391_ ;
	wire _w20390_ ;
	wire _w20389_ ;
	wire _w20388_ ;
	wire _w20387_ ;
	wire _w20386_ ;
	wire _w20385_ ;
	wire _w20384_ ;
	wire _w20383_ ;
	wire _w20382_ ;
	wire _w20381_ ;
	wire _w20380_ ;
	wire _w20379_ ;
	wire _w20378_ ;
	wire _w20377_ ;
	wire _w20376_ ;
	wire _w20375_ ;
	wire _w20374_ ;
	wire _w20373_ ;
	wire _w20372_ ;
	wire _w20371_ ;
	wire _w20370_ ;
	wire _w20369_ ;
	wire _w20368_ ;
	wire _w20367_ ;
	wire _w20366_ ;
	wire _w20365_ ;
	wire _w20364_ ;
	wire _w20363_ ;
	wire _w20362_ ;
	wire _w20361_ ;
	wire _w20360_ ;
	wire _w20359_ ;
	wire _w20358_ ;
	wire _w20357_ ;
	wire _w20356_ ;
	wire _w20355_ ;
	wire _w20354_ ;
	wire _w20353_ ;
	wire _w20352_ ;
	wire _w20351_ ;
	wire _w20350_ ;
	wire _w20349_ ;
	wire _w20348_ ;
	wire _w20347_ ;
	wire _w20346_ ;
	wire _w20345_ ;
	wire _w20344_ ;
	wire _w20343_ ;
	wire _w20342_ ;
	wire _w20341_ ;
	wire _w20340_ ;
	wire _w20339_ ;
	wire _w20338_ ;
	wire _w20337_ ;
	wire _w20336_ ;
	wire _w20335_ ;
	wire _w20334_ ;
	wire _w20333_ ;
	wire _w20332_ ;
	wire _w20331_ ;
	wire _w20330_ ;
	wire _w20329_ ;
	wire _w20328_ ;
	wire _w20327_ ;
	wire _w20326_ ;
	wire _w20325_ ;
	wire _w20324_ ;
	wire _w20323_ ;
	wire _w20322_ ;
	wire _w20321_ ;
	wire _w20320_ ;
	wire _w20319_ ;
	wire _w20318_ ;
	wire _w20317_ ;
	wire _w20316_ ;
	wire _w20315_ ;
	wire _w20314_ ;
	wire _w20313_ ;
	wire _w20312_ ;
	wire _w20311_ ;
	wire _w20310_ ;
	wire _w20309_ ;
	wire _w20308_ ;
	wire _w20307_ ;
	wire _w20306_ ;
	wire _w20305_ ;
	wire _w20304_ ;
	wire _w20303_ ;
	wire _w20302_ ;
	wire _w20301_ ;
	wire _w20300_ ;
	wire _w20299_ ;
	wire _w20298_ ;
	wire _w20297_ ;
	wire _w20296_ ;
	wire _w20295_ ;
	wire _w20294_ ;
	wire _w20293_ ;
	wire _w20292_ ;
	wire _w20291_ ;
	wire _w20290_ ;
	wire _w20289_ ;
	wire _w20288_ ;
	wire _w20287_ ;
	wire _w20286_ ;
	wire _w20285_ ;
	wire _w20284_ ;
	wire _w20283_ ;
	wire _w20282_ ;
	wire _w20281_ ;
	wire _w20280_ ;
	wire _w20279_ ;
	wire _w20278_ ;
	wire _w20277_ ;
	wire _w20276_ ;
	wire _w20275_ ;
	wire _w20274_ ;
	wire _w20273_ ;
	wire _w20272_ ;
	wire _w20271_ ;
	wire _w20270_ ;
	wire _w20269_ ;
	wire _w20268_ ;
	wire _w20267_ ;
	wire _w20266_ ;
	wire _w20265_ ;
	wire _w20264_ ;
	wire _w20263_ ;
	wire _w20262_ ;
	wire _w20261_ ;
	wire _w20260_ ;
	wire _w20259_ ;
	wire _w20258_ ;
	wire _w20257_ ;
	wire _w20256_ ;
	wire _w20255_ ;
	wire _w20254_ ;
	wire _w20253_ ;
	wire _w20252_ ;
	wire _w20251_ ;
	wire _w20250_ ;
	wire _w20249_ ;
	wire _w20248_ ;
	wire _w20247_ ;
	wire _w20246_ ;
	wire _w20245_ ;
	wire _w20244_ ;
	wire _w20243_ ;
	wire _w20242_ ;
	wire _w20241_ ;
	wire _w20240_ ;
	wire _w20239_ ;
	wire _w20238_ ;
	wire _w20237_ ;
	wire _w20236_ ;
	wire _w20235_ ;
	wire _w20234_ ;
	wire _w20233_ ;
	wire _w20232_ ;
	wire _w20231_ ;
	wire _w20230_ ;
	wire _w20229_ ;
	wire _w20228_ ;
	wire _w20227_ ;
	wire _w20226_ ;
	wire _w20225_ ;
	wire _w20224_ ;
	wire _w20223_ ;
	wire _w20222_ ;
	wire _w20221_ ;
	wire _w20220_ ;
	wire _w20219_ ;
	wire _w20218_ ;
	wire _w20217_ ;
	wire _w20216_ ;
	wire _w20215_ ;
	wire _w20214_ ;
	wire _w20213_ ;
	wire _w20212_ ;
	wire _w20211_ ;
	wire _w20210_ ;
	wire _w20209_ ;
	wire _w20208_ ;
	wire _w20207_ ;
	wire _w20206_ ;
	wire _w20205_ ;
	wire _w20204_ ;
	wire _w20203_ ;
	wire _w20202_ ;
	wire _w20201_ ;
	wire _w20200_ ;
	wire _w20199_ ;
	wire _w20198_ ;
	wire _w20197_ ;
	wire _w20196_ ;
	wire _w20195_ ;
	wire _w20194_ ;
	wire _w20193_ ;
	wire _w20192_ ;
	wire _w20191_ ;
	wire _w20190_ ;
	wire _w20189_ ;
	wire _w20188_ ;
	wire _w20187_ ;
	wire _w20186_ ;
	wire _w20185_ ;
	wire _w20184_ ;
	wire _w20183_ ;
	wire _w20182_ ;
	wire _w20181_ ;
	wire _w20180_ ;
	wire _w20179_ ;
	wire _w20178_ ;
	wire _w20177_ ;
	wire _w20176_ ;
	wire _w20175_ ;
	wire _w20174_ ;
	wire _w20173_ ;
	wire _w20172_ ;
	wire _w20171_ ;
	wire _w20170_ ;
	wire _w20169_ ;
	wire _w20168_ ;
	wire _w20167_ ;
	wire _w20166_ ;
	wire _w20165_ ;
	wire _w20164_ ;
	wire _w20163_ ;
	wire _w20162_ ;
	wire _w20161_ ;
	wire _w20160_ ;
	wire _w20159_ ;
	wire _w20158_ ;
	wire _w20157_ ;
	wire _w20156_ ;
	wire _w20155_ ;
	wire _w20154_ ;
	wire _w20153_ ;
	wire _w20152_ ;
	wire _w20151_ ;
	wire _w20150_ ;
	wire _w20149_ ;
	wire _w20148_ ;
	wire _w20147_ ;
	wire _w20146_ ;
	wire _w20145_ ;
	wire _w20144_ ;
	wire _w20143_ ;
	wire _w20142_ ;
	wire _w20141_ ;
	wire _w20140_ ;
	wire _w20139_ ;
	wire _w20138_ ;
	wire _w20137_ ;
	wire _w20136_ ;
	wire _w20135_ ;
	wire _w20134_ ;
	wire _w20133_ ;
	wire _w20132_ ;
	wire _w20131_ ;
	wire _w20130_ ;
	wire _w20129_ ;
	wire _w20128_ ;
	wire _w20127_ ;
	wire _w20126_ ;
	wire _w20125_ ;
	wire _w20124_ ;
	wire _w20123_ ;
	wire _w20122_ ;
	wire _w20121_ ;
	wire _w20120_ ;
	wire _w20119_ ;
	wire _w20118_ ;
	wire _w20117_ ;
	wire _w20116_ ;
	wire _w20115_ ;
	wire _w20114_ ;
	wire _w20113_ ;
	wire _w20112_ ;
	wire _w20111_ ;
	wire _w20110_ ;
	wire _w20109_ ;
	wire _w20108_ ;
	wire _w20107_ ;
	wire _w20106_ ;
	wire _w20105_ ;
	wire _w20104_ ;
	wire _w20103_ ;
	wire _w20102_ ;
	wire _w20101_ ;
	wire _w20100_ ;
	wire _w20099_ ;
	wire _w20098_ ;
	wire _w20097_ ;
	wire _w20096_ ;
	wire _w20095_ ;
	wire _w20094_ ;
	wire _w20093_ ;
	wire _w20092_ ;
	wire _w20091_ ;
	wire _w20090_ ;
	wire _w20089_ ;
	wire _w20088_ ;
	wire _w20087_ ;
	wire _w20086_ ;
	wire _w20085_ ;
	wire _w20084_ ;
	wire _w20083_ ;
	wire _w20082_ ;
	wire _w20081_ ;
	wire _w20080_ ;
	wire _w20079_ ;
	wire _w20078_ ;
	wire _w20077_ ;
	wire _w20076_ ;
	wire _w20075_ ;
	wire _w20074_ ;
	wire _w20073_ ;
	wire _w20072_ ;
	wire _w20071_ ;
	wire _w20070_ ;
	wire _w20069_ ;
	wire _w20068_ ;
	wire _w20067_ ;
	wire _w20066_ ;
	wire _w20065_ ;
	wire _w20064_ ;
	wire _w20063_ ;
	wire _w20062_ ;
	wire _w20061_ ;
	wire _w20060_ ;
	wire _w20059_ ;
	wire _w20058_ ;
	wire _w20057_ ;
	wire _w20056_ ;
	wire _w20055_ ;
	wire _w20054_ ;
	wire _w20053_ ;
	wire _w20052_ ;
	wire _w20051_ ;
	wire _w20050_ ;
	wire _w20049_ ;
	wire _w20048_ ;
	wire _w20047_ ;
	wire _w20046_ ;
	wire _w20045_ ;
	wire _w20044_ ;
	wire _w20043_ ;
	wire _w20042_ ;
	wire _w20041_ ;
	wire _w20040_ ;
	wire _w20039_ ;
	wire _w20038_ ;
	wire _w20037_ ;
	wire _w20036_ ;
	wire _w20035_ ;
	wire _w20034_ ;
	wire _w20033_ ;
	wire _w20032_ ;
	wire _w20031_ ;
	wire _w20030_ ;
	wire _w20029_ ;
	wire _w20028_ ;
	wire _w20027_ ;
	wire _w20026_ ;
	wire _w20025_ ;
	wire _w20024_ ;
	wire _w20023_ ;
	wire _w20022_ ;
	wire _w20021_ ;
	wire _w20020_ ;
	wire _w20019_ ;
	wire _w20018_ ;
	wire _w20017_ ;
	wire _w20016_ ;
	wire _w20015_ ;
	wire _w20014_ ;
	wire _w20013_ ;
	wire _w20012_ ;
	wire _w20011_ ;
	wire _w20010_ ;
	wire _w20009_ ;
	wire _w20008_ ;
	wire _w20007_ ;
	wire _w20006_ ;
	wire _w20005_ ;
	wire _w20004_ ;
	wire _w20003_ ;
	wire _w20002_ ;
	wire _w20001_ ;
	wire _w20000_ ;
	wire _w19999_ ;
	wire _w19998_ ;
	wire _w19997_ ;
	wire _w19996_ ;
	wire _w19995_ ;
	wire _w19994_ ;
	wire _w19993_ ;
	wire _w19992_ ;
	wire _w19991_ ;
	wire _w19990_ ;
	wire _w19989_ ;
	wire _w19988_ ;
	wire _w19987_ ;
	wire _w19986_ ;
	wire _w19985_ ;
	wire _w19984_ ;
	wire _w19983_ ;
	wire _w19982_ ;
	wire _w19981_ ;
	wire _w19980_ ;
	wire _w19979_ ;
	wire _w19978_ ;
	wire _w19977_ ;
	wire _w19976_ ;
	wire _w19975_ ;
	wire _w19974_ ;
	wire _w19973_ ;
	wire _w19972_ ;
	wire _w19971_ ;
	wire _w19970_ ;
	wire _w19969_ ;
	wire _w19968_ ;
	wire _w19967_ ;
	wire _w19966_ ;
	wire _w19965_ ;
	wire _w19964_ ;
	wire _w19963_ ;
	wire _w19962_ ;
	wire _w19961_ ;
	wire _w19960_ ;
	wire _w19959_ ;
	wire _w19958_ ;
	wire _w19957_ ;
	wire _w19956_ ;
	wire _w19955_ ;
	wire _w19954_ ;
	wire _w19953_ ;
	wire _w19952_ ;
	wire _w19951_ ;
	wire _w19950_ ;
	wire _w19949_ ;
	wire _w19948_ ;
	wire _w19947_ ;
	wire _w19946_ ;
	wire _w19945_ ;
	wire _w19944_ ;
	wire _w19943_ ;
	wire _w19942_ ;
	wire _w19941_ ;
	wire _w19940_ ;
	wire _w19939_ ;
	wire _w19938_ ;
	wire _w19937_ ;
	wire _w19936_ ;
	wire _w19935_ ;
	wire _w19934_ ;
	wire _w19933_ ;
	wire _w19932_ ;
	wire _w19931_ ;
	wire _w19930_ ;
	wire _w19929_ ;
	wire _w19928_ ;
	wire _w19927_ ;
	wire _w19926_ ;
	wire _w19925_ ;
	wire _w19924_ ;
	wire _w19923_ ;
	wire _w19922_ ;
	wire _w19921_ ;
	wire _w19920_ ;
	wire _w19919_ ;
	wire _w19918_ ;
	wire _w19917_ ;
	wire _w19916_ ;
	wire _w19915_ ;
	wire _w19914_ ;
	wire _w19913_ ;
	wire _w19912_ ;
	wire _w19911_ ;
	wire _w19910_ ;
	wire _w19909_ ;
	wire _w19908_ ;
	wire _w19907_ ;
	wire _w19906_ ;
	wire _w19905_ ;
	wire _w19904_ ;
	wire _w19903_ ;
	wire _w19902_ ;
	wire _w19901_ ;
	wire _w19900_ ;
	wire _w19899_ ;
	wire _w19898_ ;
	wire _w19897_ ;
	wire _w19896_ ;
	wire _w19895_ ;
	wire _w19894_ ;
	wire _w19893_ ;
	wire _w19892_ ;
	wire _w19891_ ;
	wire _w19890_ ;
	wire _w19889_ ;
	wire _w19888_ ;
	wire _w19887_ ;
	wire _w19886_ ;
	wire _w19885_ ;
	wire _w19884_ ;
	wire _w19883_ ;
	wire _w19882_ ;
	wire _w19881_ ;
	wire _w19880_ ;
	wire _w19879_ ;
	wire _w19878_ ;
	wire _w19877_ ;
	wire _w19876_ ;
	wire _w19875_ ;
	wire _w19874_ ;
	wire _w19873_ ;
	wire _w19872_ ;
	wire _w19871_ ;
	wire _w19870_ ;
	wire _w19869_ ;
	wire _w19868_ ;
	wire _w19867_ ;
	wire _w19866_ ;
	wire _w19865_ ;
	wire _w19864_ ;
	wire _w19863_ ;
	wire _w19862_ ;
	wire _w19861_ ;
	wire _w19860_ ;
	wire _w19859_ ;
	wire _w19858_ ;
	wire _w19857_ ;
	wire _w19856_ ;
	wire _w19855_ ;
	wire _w19854_ ;
	wire _w19853_ ;
	wire _w19852_ ;
	wire _w19851_ ;
	wire _w19850_ ;
	wire _w19849_ ;
	wire _w19848_ ;
	wire _w19847_ ;
	wire _w19846_ ;
	wire _w19845_ ;
	wire _w19844_ ;
	wire _w19843_ ;
	wire _w19842_ ;
	wire _w19841_ ;
	wire _w19840_ ;
	wire _w19839_ ;
	wire _w19838_ ;
	wire _w19837_ ;
	wire _w19836_ ;
	wire _w19835_ ;
	wire _w19834_ ;
	wire _w19833_ ;
	wire _w19832_ ;
	wire _w19831_ ;
	wire _w19830_ ;
	wire _w19829_ ;
	wire _w19828_ ;
	wire _w19827_ ;
	wire _w19826_ ;
	wire _w19825_ ;
	wire _w19824_ ;
	wire _w19823_ ;
	wire _w19822_ ;
	wire _w19821_ ;
	wire _w19820_ ;
	wire _w19819_ ;
	wire _w19818_ ;
	wire _w19817_ ;
	wire _w19816_ ;
	wire _w19815_ ;
	wire _w19814_ ;
	wire _w19813_ ;
	wire _w19812_ ;
	wire _w19811_ ;
	wire _w19810_ ;
	wire _w19809_ ;
	wire _w19808_ ;
	wire _w19807_ ;
	wire _w19806_ ;
	wire _w19805_ ;
	wire _w19804_ ;
	wire _w19803_ ;
	wire _w19802_ ;
	wire _w19801_ ;
	wire _w19800_ ;
	wire _w19799_ ;
	wire _w19798_ ;
	wire _w19797_ ;
	wire _w19796_ ;
	wire _w19795_ ;
	wire _w19794_ ;
	wire _w19793_ ;
	wire _w19792_ ;
	wire _w19791_ ;
	wire _w19790_ ;
	wire _w19789_ ;
	wire _w19788_ ;
	wire _w19787_ ;
	wire _w19786_ ;
	wire _w19785_ ;
	wire _w19784_ ;
	wire _w19783_ ;
	wire _w19782_ ;
	wire _w19781_ ;
	wire _w19780_ ;
	wire _w19779_ ;
	wire _w19778_ ;
	wire _w19777_ ;
	wire _w19776_ ;
	wire _w19775_ ;
	wire _w19774_ ;
	wire _w19773_ ;
	wire _w19772_ ;
	wire _w19771_ ;
	wire _w19770_ ;
	wire _w19769_ ;
	wire _w19768_ ;
	wire _w19767_ ;
	wire _w19766_ ;
	wire _w19765_ ;
	wire _w19764_ ;
	wire _w19763_ ;
	wire _w19762_ ;
	wire _w19761_ ;
	wire _w19760_ ;
	wire _w19759_ ;
	wire _w19758_ ;
	wire _w19757_ ;
	wire _w19756_ ;
	wire _w19755_ ;
	wire _w19754_ ;
	wire _w19753_ ;
	wire _w19752_ ;
	wire _w19751_ ;
	wire _w19750_ ;
	wire _w19749_ ;
	wire _w19748_ ;
	wire _w19747_ ;
	wire _w19746_ ;
	wire _w19745_ ;
	wire _w19744_ ;
	wire _w19743_ ;
	wire _w19742_ ;
	wire _w19741_ ;
	wire _w19740_ ;
	wire _w19739_ ;
	wire _w19738_ ;
	wire _w19737_ ;
	wire _w19736_ ;
	wire _w19735_ ;
	wire _w19734_ ;
	wire _w19733_ ;
	wire _w19732_ ;
	wire _w19731_ ;
	wire _w19730_ ;
	wire _w19729_ ;
	wire _w19728_ ;
	wire _w19727_ ;
	wire _w19726_ ;
	wire _w19725_ ;
	wire _w19724_ ;
	wire _w19723_ ;
	wire _w19722_ ;
	wire _w19721_ ;
	wire _w19720_ ;
	wire _w19719_ ;
	wire _w19718_ ;
	wire _w19717_ ;
	wire _w19716_ ;
	wire _w19715_ ;
	wire _w19714_ ;
	wire _w19713_ ;
	wire _w19712_ ;
	wire _w19711_ ;
	wire _w19710_ ;
	wire _w19709_ ;
	wire _w19708_ ;
	wire _w19707_ ;
	wire _w19706_ ;
	wire _w19705_ ;
	wire _w19704_ ;
	wire _w19703_ ;
	wire _w19702_ ;
	wire _w19701_ ;
	wire _w19700_ ;
	wire _w19699_ ;
	wire _w19698_ ;
	wire _w19697_ ;
	wire _w19696_ ;
	wire _w19695_ ;
	wire _w19694_ ;
	wire _w19693_ ;
	wire _w19692_ ;
	wire _w19691_ ;
	wire _w19690_ ;
	wire _w19689_ ;
	wire _w19688_ ;
	wire _w19687_ ;
	wire _w19686_ ;
	wire _w19685_ ;
	wire _w19684_ ;
	wire _w19683_ ;
	wire _w19682_ ;
	wire _w19681_ ;
	wire _w19680_ ;
	wire _w19679_ ;
	wire _w19678_ ;
	wire _w19677_ ;
	wire _w19676_ ;
	wire _w19675_ ;
	wire _w19674_ ;
	wire _w19673_ ;
	wire _w19672_ ;
	wire _w19671_ ;
	wire _w19670_ ;
	wire _w19669_ ;
	wire _w19668_ ;
	wire _w19667_ ;
	wire _w19666_ ;
	wire _w19665_ ;
	wire _w19664_ ;
	wire _w19663_ ;
	wire _w19662_ ;
	wire _w19661_ ;
	wire _w19660_ ;
	wire _w19659_ ;
	wire _w19658_ ;
	wire _w19657_ ;
	wire _w19656_ ;
	wire _w19655_ ;
	wire _w19654_ ;
	wire _w19653_ ;
	wire _w19652_ ;
	wire _w19651_ ;
	wire _w19650_ ;
	wire _w19649_ ;
	wire _w19648_ ;
	wire _w19647_ ;
	wire _w19646_ ;
	wire _w19645_ ;
	wire _w19644_ ;
	wire _w19643_ ;
	wire _w19642_ ;
	wire _w19641_ ;
	wire _w19640_ ;
	wire _w19639_ ;
	wire _w19638_ ;
	wire _w19637_ ;
	wire _w19636_ ;
	wire _w19635_ ;
	wire _w19634_ ;
	wire _w19633_ ;
	wire _w19632_ ;
	wire _w19631_ ;
	wire _w19630_ ;
	wire _w19629_ ;
	wire _w19628_ ;
	wire _w19627_ ;
	wire _w19626_ ;
	wire _w19625_ ;
	wire _w19624_ ;
	wire _w19623_ ;
	wire _w19622_ ;
	wire _w19621_ ;
	wire _w19620_ ;
	wire _w19619_ ;
	wire _w19618_ ;
	wire _w19617_ ;
	wire _w19616_ ;
	wire _w19615_ ;
	wire _w19614_ ;
	wire _w19613_ ;
	wire _w19612_ ;
	wire _w19611_ ;
	wire _w19610_ ;
	wire _w19609_ ;
	wire _w19608_ ;
	wire _w19607_ ;
	wire _w19606_ ;
	wire _w19605_ ;
	wire _w19604_ ;
	wire _w19603_ ;
	wire _w19602_ ;
	wire _w19601_ ;
	wire _w19600_ ;
	wire _w19599_ ;
	wire _w19598_ ;
	wire _w19597_ ;
	wire _w19596_ ;
	wire _w19595_ ;
	wire _w19594_ ;
	wire _w19593_ ;
	wire _w19592_ ;
	wire _w19591_ ;
	wire _w19590_ ;
	wire _w19589_ ;
	wire _w19588_ ;
	wire _w19587_ ;
	wire _w19586_ ;
	wire _w19585_ ;
	wire _w19584_ ;
	wire _w19583_ ;
	wire _w19582_ ;
	wire _w19581_ ;
	wire _w19580_ ;
	wire _w19579_ ;
	wire _w19578_ ;
	wire _w19577_ ;
	wire _w19576_ ;
	wire _w19575_ ;
	wire _w19574_ ;
	wire _w19573_ ;
	wire _w19572_ ;
	wire _w19571_ ;
	wire _w19570_ ;
	wire _w19569_ ;
	wire _w19568_ ;
	wire _w19567_ ;
	wire _w19566_ ;
	wire _w19565_ ;
	wire _w19564_ ;
	wire _w19563_ ;
	wire _w19562_ ;
	wire _w19561_ ;
	wire _w19560_ ;
	wire _w19559_ ;
	wire _w19558_ ;
	wire _w19557_ ;
	wire _w19556_ ;
	wire _w19555_ ;
	wire _w19554_ ;
	wire _w19553_ ;
	wire _w19552_ ;
	wire _w19551_ ;
	wire _w19550_ ;
	wire _w19549_ ;
	wire _w19548_ ;
	wire _w19547_ ;
	wire _w19546_ ;
	wire _w19545_ ;
	wire _w19544_ ;
	wire _w19543_ ;
	wire _w19542_ ;
	wire _w19541_ ;
	wire _w19540_ ;
	wire _w19539_ ;
	wire _w19538_ ;
	wire _w19537_ ;
	wire _w19536_ ;
	wire _w19535_ ;
	wire _w19534_ ;
	wire _w19533_ ;
	wire _w19532_ ;
	wire _w19531_ ;
	wire _w19530_ ;
	wire _w19529_ ;
	wire _w19528_ ;
	wire _w19527_ ;
	wire _w19526_ ;
	wire _w19525_ ;
	wire _w19524_ ;
	wire _w19523_ ;
	wire _w19522_ ;
	wire _w19521_ ;
	wire _w19520_ ;
	wire _w19519_ ;
	wire _w19518_ ;
	wire _w19517_ ;
	wire _w19516_ ;
	wire _w19515_ ;
	wire _w19514_ ;
	wire _w19513_ ;
	wire _w19512_ ;
	wire _w19511_ ;
	wire _w19510_ ;
	wire _w19509_ ;
	wire _w19508_ ;
	wire _w19507_ ;
	wire _w19506_ ;
	wire _w19505_ ;
	wire _w19504_ ;
	wire _w19503_ ;
	wire _w19502_ ;
	wire _w19501_ ;
	wire _w19500_ ;
	wire _w19499_ ;
	wire _w19498_ ;
	wire _w19497_ ;
	wire _w19496_ ;
	wire _w19495_ ;
	wire _w19494_ ;
	wire _w19493_ ;
	wire _w19492_ ;
	wire _w19491_ ;
	wire _w19490_ ;
	wire _w19489_ ;
	wire _w19488_ ;
	wire _w19487_ ;
	wire _w19486_ ;
	wire _w19485_ ;
	wire _w19484_ ;
	wire _w19483_ ;
	wire _w19482_ ;
	wire _w19481_ ;
	wire _w19480_ ;
	wire _w19479_ ;
	wire _w19478_ ;
	wire _w19477_ ;
	wire _w19476_ ;
	wire _w19475_ ;
	wire _w19474_ ;
	wire _w19473_ ;
	wire _w19472_ ;
	wire _w19471_ ;
	wire _w19470_ ;
	wire _w19469_ ;
	wire _w19468_ ;
	wire _w19467_ ;
	wire _w19466_ ;
	wire _w19465_ ;
	wire _w19464_ ;
	wire _w19463_ ;
	wire _w19462_ ;
	wire _w19461_ ;
	wire _w19460_ ;
	wire _w19459_ ;
	wire _w19458_ ;
	wire _w19457_ ;
	wire _w19456_ ;
	wire _w19455_ ;
	wire _w19454_ ;
	wire _w19453_ ;
	wire _w19452_ ;
	wire _w19451_ ;
	wire _w19450_ ;
	wire _w19449_ ;
	wire _w19448_ ;
	wire _w19447_ ;
	wire _w19446_ ;
	wire _w19445_ ;
	wire _w19444_ ;
	wire _w19443_ ;
	wire _w19442_ ;
	wire _w19441_ ;
	wire _w19440_ ;
	wire _w19439_ ;
	wire _w19438_ ;
	wire _w19437_ ;
	wire _w19436_ ;
	wire _w19435_ ;
	wire _w19434_ ;
	wire _w19433_ ;
	wire _w19432_ ;
	wire _w19431_ ;
	wire _w19430_ ;
	wire _w19429_ ;
	wire _w19428_ ;
	wire _w19427_ ;
	wire _w19426_ ;
	wire _w19425_ ;
	wire _w19424_ ;
	wire _w19423_ ;
	wire _w19422_ ;
	wire _w19421_ ;
	wire _w19420_ ;
	wire _w19419_ ;
	wire _w19418_ ;
	wire _w19417_ ;
	wire _w19416_ ;
	wire _w19415_ ;
	wire _w19414_ ;
	wire _w19413_ ;
	wire _w19412_ ;
	wire _w19411_ ;
	wire _w19410_ ;
	wire _w19409_ ;
	wire _w19408_ ;
	wire _w19407_ ;
	wire _w19406_ ;
	wire _w19405_ ;
	wire _w19404_ ;
	wire _w19403_ ;
	wire _w19402_ ;
	wire _w19401_ ;
	wire _w19400_ ;
	wire _w19399_ ;
	wire _w19398_ ;
	wire _w19397_ ;
	wire _w19396_ ;
	wire _w19395_ ;
	wire _w19394_ ;
	wire _w19393_ ;
	wire _w19392_ ;
	wire _w19391_ ;
	wire _w19390_ ;
	wire _w19389_ ;
	wire _w19388_ ;
	wire _w19387_ ;
	wire _w19386_ ;
	wire _w19385_ ;
	wire _w19384_ ;
	wire _w19383_ ;
	wire _w19382_ ;
	wire _w19381_ ;
	wire _w19380_ ;
	wire _w19379_ ;
	wire _w19378_ ;
	wire _w19377_ ;
	wire _w19376_ ;
	wire _w19375_ ;
	wire _w19374_ ;
	wire _w19373_ ;
	wire _w19372_ ;
	wire _w19371_ ;
	wire _w19370_ ;
	wire _w19369_ ;
	wire _w19368_ ;
	wire _w19367_ ;
	wire _w19366_ ;
	wire _w19365_ ;
	wire _w19364_ ;
	wire _w19363_ ;
	wire _w19362_ ;
	wire _w19361_ ;
	wire _w19360_ ;
	wire _w19359_ ;
	wire _w19358_ ;
	wire _w19357_ ;
	wire _w19356_ ;
	wire _w19355_ ;
	wire _w19354_ ;
	wire _w19353_ ;
	wire _w19352_ ;
	wire _w19351_ ;
	wire _w19350_ ;
	wire _w19349_ ;
	wire _w19348_ ;
	wire _w19347_ ;
	wire _w19346_ ;
	wire _w19345_ ;
	wire _w19344_ ;
	wire _w19343_ ;
	wire _w19342_ ;
	wire _w19341_ ;
	wire _w19340_ ;
	wire _w19339_ ;
	wire _w19338_ ;
	wire _w19337_ ;
	wire _w19336_ ;
	wire _w19335_ ;
	wire _w19334_ ;
	wire _w19333_ ;
	wire _w19332_ ;
	wire _w19331_ ;
	wire _w19330_ ;
	wire _w19329_ ;
	wire _w19328_ ;
	wire _w19327_ ;
	wire _w19326_ ;
	wire _w19325_ ;
	wire _w19324_ ;
	wire _w19323_ ;
	wire _w19322_ ;
	wire _w19321_ ;
	wire _w19320_ ;
	wire _w19319_ ;
	wire _w19318_ ;
	wire _w19317_ ;
	wire _w19316_ ;
	wire _w19315_ ;
	wire _w19314_ ;
	wire _w19313_ ;
	wire _w19312_ ;
	wire _w19311_ ;
	wire _w19310_ ;
	wire _w19309_ ;
	wire _w19308_ ;
	wire _w19307_ ;
	wire _w19306_ ;
	wire _w19305_ ;
	wire _w19304_ ;
	wire _w19303_ ;
	wire _w19302_ ;
	wire _w19301_ ;
	wire _w19300_ ;
	wire _w19299_ ;
	wire _w19298_ ;
	wire _w19297_ ;
	wire _w19296_ ;
	wire _w19295_ ;
	wire _w19294_ ;
	wire _w19293_ ;
	wire _w19292_ ;
	wire _w19291_ ;
	wire _w19290_ ;
	wire _w19289_ ;
	wire _w19288_ ;
	wire _w19287_ ;
	wire _w19286_ ;
	wire _w19285_ ;
	wire _w19284_ ;
	wire _w19283_ ;
	wire _w19282_ ;
	wire _w19281_ ;
	wire _w19280_ ;
	wire _w19279_ ;
	wire _w19278_ ;
	wire _w19277_ ;
	wire _w19276_ ;
	wire _w19275_ ;
	wire _w19274_ ;
	wire _w19273_ ;
	wire _w19272_ ;
	wire _w19271_ ;
	wire _w19270_ ;
	wire _w19269_ ;
	wire _w19268_ ;
	wire _w19267_ ;
	wire _w19266_ ;
	wire _w19265_ ;
	wire _w19264_ ;
	wire _w19263_ ;
	wire _w19262_ ;
	wire _w19261_ ;
	wire _w19260_ ;
	wire _w19259_ ;
	wire _w19258_ ;
	wire _w19257_ ;
	wire _w19256_ ;
	wire _w19255_ ;
	wire _w19254_ ;
	wire _w19253_ ;
	wire _w19252_ ;
	wire _w19251_ ;
	wire _w19250_ ;
	wire _w19249_ ;
	wire _w19248_ ;
	wire _w19247_ ;
	wire _w19246_ ;
	wire _w19245_ ;
	wire _w19244_ ;
	wire _w19243_ ;
	wire _w19242_ ;
	wire _w19241_ ;
	wire _w19240_ ;
	wire _w19239_ ;
	wire _w19238_ ;
	wire _w19237_ ;
	wire _w19236_ ;
	wire _w19235_ ;
	wire _w19234_ ;
	wire _w19233_ ;
	wire _w19232_ ;
	wire _w19231_ ;
	wire _w19230_ ;
	wire _w19229_ ;
	wire _w19228_ ;
	wire _w19227_ ;
	wire _w19226_ ;
	wire _w19225_ ;
	wire _w19224_ ;
	wire _w19223_ ;
	wire _w19222_ ;
	wire _w19221_ ;
	wire _w19220_ ;
	wire _w19219_ ;
	wire _w19218_ ;
	wire _w19217_ ;
	wire _w19216_ ;
	wire _w19215_ ;
	wire _w19214_ ;
	wire _w19213_ ;
	wire _w19212_ ;
	wire _w19211_ ;
	wire _w19210_ ;
	wire _w19209_ ;
	wire _w19208_ ;
	wire _w19207_ ;
	wire _w19206_ ;
	wire _w19205_ ;
	wire _w19204_ ;
	wire _w19203_ ;
	wire _w19202_ ;
	wire _w19201_ ;
	wire _w19200_ ;
	wire _w19199_ ;
	wire _w19198_ ;
	wire _w19197_ ;
	wire _w19196_ ;
	wire _w19195_ ;
	wire _w19194_ ;
	wire _w19193_ ;
	wire _w19192_ ;
	wire _w19191_ ;
	wire _w19190_ ;
	wire _w19189_ ;
	wire _w19188_ ;
	wire _w19187_ ;
	wire _w19186_ ;
	wire _w19185_ ;
	wire _w19184_ ;
	wire _w19183_ ;
	wire _w19182_ ;
	wire _w19181_ ;
	wire _w19180_ ;
	wire _w19179_ ;
	wire _w19178_ ;
	wire _w19177_ ;
	wire _w19176_ ;
	wire _w19175_ ;
	wire _w19174_ ;
	wire _w19173_ ;
	wire _w19172_ ;
	wire _w19171_ ;
	wire _w19170_ ;
	wire _w19169_ ;
	wire _w19168_ ;
	wire _w19167_ ;
	wire _w19166_ ;
	wire _w19165_ ;
	wire _w19164_ ;
	wire _w19163_ ;
	wire _w19162_ ;
	wire _w19161_ ;
	wire _w19160_ ;
	wire _w19159_ ;
	wire _w19158_ ;
	wire _w19157_ ;
	wire _w19156_ ;
	wire _w19155_ ;
	wire _w19154_ ;
	wire _w19153_ ;
	wire _w19152_ ;
	wire _w19151_ ;
	wire _w19150_ ;
	wire _w19149_ ;
	wire _w19148_ ;
	wire _w19147_ ;
	wire _w19146_ ;
	wire _w19145_ ;
	wire _w19144_ ;
	wire _w19143_ ;
	wire _w19142_ ;
	wire _w19141_ ;
	wire _w19140_ ;
	wire _w19139_ ;
	wire _w19138_ ;
	wire _w19137_ ;
	wire _w19136_ ;
	wire _w19135_ ;
	wire _w19134_ ;
	wire _w19133_ ;
	wire _w19132_ ;
	wire _w19131_ ;
	wire _w19130_ ;
	wire _w19129_ ;
	wire _w19128_ ;
	wire _w19127_ ;
	wire _w19126_ ;
	wire _w19125_ ;
	wire _w19124_ ;
	wire _w19123_ ;
	wire _w19122_ ;
	wire _w19121_ ;
	wire _w19120_ ;
	wire _w19119_ ;
	wire _w19118_ ;
	wire _w19117_ ;
	wire _w19116_ ;
	wire _w19115_ ;
	wire _w19114_ ;
	wire _w19113_ ;
	wire _w19112_ ;
	wire _w19111_ ;
	wire _w19110_ ;
	wire _w19109_ ;
	wire _w19108_ ;
	wire _w19107_ ;
	wire _w19106_ ;
	wire _w19105_ ;
	wire _w19104_ ;
	wire _w19103_ ;
	wire _w19102_ ;
	wire _w19101_ ;
	wire _w19100_ ;
	wire _w19099_ ;
	wire _w19098_ ;
	wire _w19097_ ;
	wire _w19096_ ;
	wire _w19095_ ;
	wire _w19094_ ;
	wire _w19093_ ;
	wire _w19092_ ;
	wire _w19091_ ;
	wire _w19090_ ;
	wire _w19089_ ;
	wire _w19088_ ;
	wire _w19087_ ;
	wire _w19086_ ;
	wire _w19085_ ;
	wire _w19084_ ;
	wire _w19083_ ;
	wire _w19082_ ;
	wire _w19081_ ;
	wire _w19080_ ;
	wire _w19079_ ;
	wire _w19078_ ;
	wire _w19077_ ;
	wire _w19076_ ;
	wire _w19075_ ;
	wire _w19074_ ;
	wire _w19073_ ;
	wire _w19072_ ;
	wire _w19071_ ;
	wire _w19070_ ;
	wire _w19069_ ;
	wire _w19068_ ;
	wire _w19067_ ;
	wire _w19066_ ;
	wire _w19065_ ;
	wire _w19064_ ;
	wire _w19063_ ;
	wire _w19062_ ;
	wire _w19061_ ;
	wire _w19060_ ;
	wire _w19059_ ;
	wire _w19058_ ;
	wire _w19057_ ;
	wire _w19056_ ;
	wire _w19055_ ;
	wire _w19054_ ;
	wire _w19053_ ;
	wire _w19052_ ;
	wire _w19051_ ;
	wire _w19050_ ;
	wire _w19049_ ;
	wire _w19048_ ;
	wire _w19047_ ;
	wire _w19046_ ;
	wire _w19045_ ;
	wire _w19044_ ;
	wire _w19043_ ;
	wire _w19042_ ;
	wire _w19041_ ;
	wire _w19040_ ;
	wire _w19039_ ;
	wire _w19038_ ;
	wire _w19037_ ;
	wire _w19036_ ;
	wire _w19035_ ;
	wire _w19034_ ;
	wire _w19033_ ;
	wire _w19032_ ;
	wire _w19031_ ;
	wire _w19030_ ;
	wire _w19029_ ;
	wire _w19028_ ;
	wire _w19027_ ;
	wire _w19026_ ;
	wire _w19025_ ;
	wire _w19024_ ;
	wire _w19023_ ;
	wire _w19022_ ;
	wire _w19021_ ;
	wire _w19020_ ;
	wire _w19019_ ;
	wire _w19018_ ;
	wire _w19017_ ;
	wire _w19016_ ;
	wire _w19015_ ;
	wire _w19014_ ;
	wire _w19013_ ;
	wire _w19012_ ;
	wire _w19011_ ;
	wire _w19010_ ;
	wire _w19009_ ;
	wire _w19008_ ;
	wire _w19007_ ;
	wire _w19006_ ;
	wire _w19005_ ;
	wire _w19004_ ;
	wire _w19003_ ;
	wire _w19002_ ;
	wire _w19001_ ;
	wire _w19000_ ;
	wire _w18999_ ;
	wire _w18998_ ;
	wire _w18997_ ;
	wire _w18996_ ;
	wire _w18995_ ;
	wire _w18994_ ;
	wire _w18993_ ;
	wire _w18992_ ;
	wire _w18991_ ;
	wire _w18990_ ;
	wire _w18989_ ;
	wire _w18988_ ;
	wire _w18987_ ;
	wire _w18986_ ;
	wire _w18985_ ;
	wire _w18984_ ;
	wire _w18983_ ;
	wire _w18982_ ;
	wire _w18981_ ;
	wire _w18980_ ;
	wire _w18979_ ;
	wire _w18978_ ;
	wire _w18977_ ;
	wire _w18976_ ;
	wire _w18975_ ;
	wire _w18974_ ;
	wire _w18973_ ;
	wire _w18972_ ;
	wire _w18971_ ;
	wire _w18970_ ;
	wire _w18969_ ;
	wire _w18968_ ;
	wire _w18967_ ;
	wire _w18966_ ;
	wire _w18965_ ;
	wire _w18964_ ;
	wire _w18963_ ;
	wire _w18962_ ;
	wire _w18961_ ;
	wire _w18960_ ;
	wire _w18959_ ;
	wire _w18958_ ;
	wire _w18957_ ;
	wire _w18956_ ;
	wire _w18955_ ;
	wire _w18954_ ;
	wire _w18953_ ;
	wire _w18952_ ;
	wire _w18951_ ;
	wire _w18950_ ;
	wire _w18949_ ;
	wire _w18948_ ;
	wire _w18947_ ;
	wire _w18946_ ;
	wire _w18945_ ;
	wire _w18944_ ;
	wire _w18943_ ;
	wire _w18942_ ;
	wire _w18941_ ;
	wire _w18940_ ;
	wire _w18939_ ;
	wire _w18938_ ;
	wire _w18937_ ;
	wire _w18936_ ;
	wire _w18935_ ;
	wire _w18934_ ;
	wire _w18933_ ;
	wire _w18932_ ;
	wire _w18931_ ;
	wire _w18930_ ;
	wire _w18929_ ;
	wire _w18928_ ;
	wire _w18927_ ;
	wire _w18926_ ;
	wire _w18925_ ;
	wire _w18924_ ;
	wire _w18923_ ;
	wire _w18922_ ;
	wire _w18921_ ;
	wire _w18920_ ;
	wire _w18919_ ;
	wire _w18918_ ;
	wire _w18917_ ;
	wire _w18916_ ;
	wire _w18915_ ;
	wire _w18914_ ;
	wire _w18913_ ;
	wire _w18912_ ;
	wire _w18911_ ;
	wire _w18910_ ;
	wire _w18909_ ;
	wire _w18908_ ;
	wire _w18907_ ;
	wire _w18906_ ;
	wire _w18905_ ;
	wire _w18904_ ;
	wire _w18903_ ;
	wire _w18902_ ;
	wire _w18901_ ;
	wire _w18900_ ;
	wire _w18899_ ;
	wire _w18898_ ;
	wire _w18897_ ;
	wire _w18896_ ;
	wire _w18895_ ;
	wire _w18894_ ;
	wire _w18893_ ;
	wire _w18892_ ;
	wire _w18891_ ;
	wire _w18890_ ;
	wire _w18889_ ;
	wire _w18888_ ;
	wire _w18887_ ;
	wire _w18886_ ;
	wire _w18885_ ;
	wire _w18884_ ;
	wire _w18883_ ;
	wire _w18882_ ;
	wire _w18881_ ;
	wire _w18880_ ;
	wire _w18879_ ;
	wire _w18878_ ;
	wire _w18877_ ;
	wire _w18876_ ;
	wire _w18875_ ;
	wire _w18874_ ;
	wire _w18873_ ;
	wire _w18872_ ;
	wire _w18871_ ;
	wire _w18870_ ;
	wire _w18869_ ;
	wire _w18868_ ;
	wire _w18867_ ;
	wire _w18866_ ;
	wire _w18865_ ;
	wire _w18864_ ;
	wire _w18863_ ;
	wire _w18862_ ;
	wire _w18861_ ;
	wire _w18860_ ;
	wire _w18859_ ;
	wire _w18858_ ;
	wire _w18857_ ;
	wire _w18856_ ;
	wire _w18855_ ;
	wire _w18854_ ;
	wire _w18853_ ;
	wire _w18852_ ;
	wire _w18851_ ;
	wire _w18850_ ;
	wire _w18849_ ;
	wire _w18848_ ;
	wire _w18847_ ;
	wire _w18846_ ;
	wire _w18845_ ;
	wire _w18844_ ;
	wire _w18843_ ;
	wire _w18842_ ;
	wire _w18841_ ;
	wire _w18840_ ;
	wire _w18839_ ;
	wire _w18838_ ;
	wire _w18837_ ;
	wire _w18836_ ;
	wire _w18835_ ;
	wire _w18834_ ;
	wire _w18833_ ;
	wire _w18832_ ;
	wire _w18831_ ;
	wire _w18830_ ;
	wire _w18829_ ;
	wire _w18828_ ;
	wire _w18827_ ;
	wire _w18826_ ;
	wire _w18825_ ;
	wire _w18824_ ;
	wire _w18823_ ;
	wire _w18822_ ;
	wire _w18821_ ;
	wire _w18820_ ;
	wire _w18819_ ;
	wire _w18818_ ;
	wire _w18817_ ;
	wire _w18816_ ;
	wire _w18815_ ;
	wire _w18814_ ;
	wire _w18813_ ;
	wire _w18812_ ;
	wire _w18811_ ;
	wire _w18810_ ;
	wire _w18809_ ;
	wire _w18808_ ;
	wire _w18807_ ;
	wire _w18806_ ;
	wire _w18805_ ;
	wire _w18804_ ;
	wire _w18803_ ;
	wire _w18802_ ;
	wire _w18801_ ;
	wire _w18800_ ;
	wire _w18799_ ;
	wire _w18798_ ;
	wire _w18797_ ;
	wire _w18796_ ;
	wire _w18795_ ;
	wire _w18794_ ;
	wire _w18793_ ;
	wire _w18792_ ;
	wire _w18791_ ;
	wire _w18790_ ;
	wire _w18789_ ;
	wire _w18788_ ;
	wire _w18787_ ;
	wire _w18786_ ;
	wire _w18785_ ;
	wire _w18784_ ;
	wire _w18783_ ;
	wire _w18782_ ;
	wire _w18781_ ;
	wire _w18780_ ;
	wire _w18779_ ;
	wire _w18778_ ;
	wire _w18777_ ;
	wire _w18776_ ;
	wire _w18775_ ;
	wire _w18774_ ;
	wire _w18773_ ;
	wire _w18772_ ;
	wire _w18771_ ;
	wire _w18770_ ;
	wire _w18769_ ;
	wire _w18768_ ;
	wire _w18767_ ;
	wire _w18766_ ;
	wire _w18765_ ;
	wire _w18764_ ;
	wire _w18763_ ;
	wire _w18762_ ;
	wire _w18761_ ;
	wire _w18760_ ;
	wire _w18759_ ;
	wire _w18758_ ;
	wire _w18757_ ;
	wire _w18756_ ;
	wire _w18755_ ;
	wire _w18754_ ;
	wire _w18753_ ;
	wire _w18752_ ;
	wire _w18751_ ;
	wire _w18750_ ;
	wire _w18749_ ;
	wire _w18748_ ;
	wire _w18747_ ;
	wire _w18746_ ;
	wire _w18745_ ;
	wire _w18744_ ;
	wire _w18743_ ;
	wire _w18742_ ;
	wire _w18741_ ;
	wire _w18740_ ;
	wire _w18739_ ;
	wire _w18738_ ;
	wire _w18737_ ;
	wire _w18736_ ;
	wire _w18735_ ;
	wire _w18734_ ;
	wire _w18733_ ;
	wire _w18732_ ;
	wire _w18731_ ;
	wire _w18730_ ;
	wire _w18729_ ;
	wire _w18728_ ;
	wire _w18727_ ;
	wire _w18726_ ;
	wire _w18725_ ;
	wire _w18724_ ;
	wire _w18723_ ;
	wire _w18722_ ;
	wire _w18721_ ;
	wire _w18720_ ;
	wire _w18719_ ;
	wire _w18718_ ;
	wire _w18717_ ;
	wire _w18716_ ;
	wire _w18715_ ;
	wire _w18714_ ;
	wire _w18713_ ;
	wire _w18712_ ;
	wire _w18711_ ;
	wire _w18710_ ;
	wire _w18709_ ;
	wire _w18708_ ;
	wire _w18707_ ;
	wire _w18706_ ;
	wire _w18705_ ;
	wire _w18704_ ;
	wire _w18703_ ;
	wire _w18702_ ;
	wire _w18701_ ;
	wire _w18700_ ;
	wire _w18699_ ;
	wire _w18698_ ;
	wire _w18697_ ;
	wire _w18696_ ;
	wire _w18695_ ;
	wire _w18694_ ;
	wire _w18693_ ;
	wire _w18692_ ;
	wire _w18691_ ;
	wire _w18690_ ;
	wire _w18689_ ;
	wire _w18688_ ;
	wire _w18687_ ;
	wire _w18686_ ;
	wire _w18685_ ;
	wire _w18684_ ;
	wire _w18683_ ;
	wire _w18682_ ;
	wire _w18681_ ;
	wire _w18680_ ;
	wire _w18679_ ;
	wire _w18678_ ;
	wire _w18677_ ;
	wire _w18676_ ;
	wire _w18675_ ;
	wire _w18674_ ;
	wire _w18673_ ;
	wire _w18672_ ;
	wire _w18671_ ;
	wire _w18670_ ;
	wire _w18669_ ;
	wire _w18668_ ;
	wire _w18667_ ;
	wire _w18666_ ;
	wire _w18665_ ;
	wire _w18664_ ;
	wire _w18663_ ;
	wire _w18662_ ;
	wire _w18661_ ;
	wire _w18660_ ;
	wire _w18659_ ;
	wire _w18658_ ;
	wire _w18657_ ;
	wire _w18656_ ;
	wire _w18655_ ;
	wire _w18654_ ;
	wire _w18653_ ;
	wire _w18652_ ;
	wire _w18651_ ;
	wire _w18650_ ;
	wire _w18649_ ;
	wire _w18648_ ;
	wire _w18647_ ;
	wire _w18646_ ;
	wire _w18645_ ;
	wire _w18644_ ;
	wire _w18643_ ;
	wire _w18642_ ;
	wire _w18641_ ;
	wire _w18640_ ;
	wire _w18639_ ;
	wire _w18638_ ;
	wire _w18637_ ;
	wire _w18636_ ;
	wire _w18635_ ;
	wire _w18634_ ;
	wire _w18633_ ;
	wire _w18632_ ;
	wire _w18631_ ;
	wire _w18630_ ;
	wire _w18629_ ;
	wire _w18628_ ;
	wire _w18627_ ;
	wire _w18626_ ;
	wire _w18625_ ;
	wire _w18624_ ;
	wire _w18623_ ;
	wire _w18622_ ;
	wire _w18621_ ;
	wire _w18620_ ;
	wire _w18619_ ;
	wire _w18618_ ;
	wire _w18617_ ;
	wire _w18616_ ;
	wire _w18615_ ;
	wire _w18614_ ;
	wire _w18613_ ;
	wire _w18612_ ;
	wire _w18611_ ;
	wire _w18610_ ;
	wire _w18609_ ;
	wire _w18608_ ;
	wire _w18607_ ;
	wire _w18606_ ;
	wire _w18605_ ;
	wire _w18604_ ;
	wire _w18603_ ;
	wire _w18602_ ;
	wire _w18601_ ;
	wire _w18600_ ;
	wire _w18599_ ;
	wire _w18598_ ;
	wire _w18597_ ;
	wire _w18596_ ;
	wire _w18595_ ;
	wire _w18594_ ;
	wire _w18593_ ;
	wire _w18592_ ;
	wire _w18591_ ;
	wire _w18590_ ;
	wire _w18589_ ;
	wire _w18588_ ;
	wire _w18587_ ;
	wire _w18586_ ;
	wire _w18585_ ;
	wire _w18584_ ;
	wire _w18583_ ;
	wire _w18582_ ;
	wire _w18581_ ;
	wire _w18580_ ;
	wire _w18579_ ;
	wire _w18578_ ;
	wire _w18577_ ;
	wire _w18576_ ;
	wire _w18575_ ;
	wire _w18574_ ;
	wire _w18573_ ;
	wire _w18572_ ;
	wire _w18571_ ;
	wire _w18570_ ;
	wire _w18569_ ;
	wire _w18568_ ;
	wire _w18567_ ;
	wire _w18566_ ;
	wire _w18565_ ;
	wire _w18564_ ;
	wire _w18563_ ;
	wire _w18562_ ;
	wire _w18561_ ;
	wire _w18560_ ;
	wire _w18559_ ;
	wire _w18558_ ;
	wire _w18557_ ;
	wire _w18556_ ;
	wire _w18555_ ;
	wire _w18554_ ;
	wire _w18553_ ;
	wire _w18552_ ;
	wire _w18551_ ;
	wire _w18550_ ;
	wire _w18549_ ;
	wire _w18548_ ;
	wire _w18547_ ;
	wire _w18546_ ;
	wire _w18545_ ;
	wire _w18544_ ;
	wire _w18543_ ;
	wire _w18542_ ;
	wire _w18541_ ;
	wire _w18540_ ;
	wire _w18539_ ;
	wire _w18538_ ;
	wire _w18537_ ;
	wire _w18536_ ;
	wire _w18535_ ;
	wire _w18534_ ;
	wire _w18533_ ;
	wire _w18532_ ;
	wire _w18531_ ;
	wire _w18530_ ;
	wire _w18529_ ;
	wire _w18528_ ;
	wire _w18527_ ;
	wire _w18526_ ;
	wire _w18525_ ;
	wire _w18524_ ;
	wire _w18523_ ;
	wire _w18522_ ;
	wire _w18521_ ;
	wire _w18520_ ;
	wire _w18519_ ;
	wire _w18518_ ;
	wire _w18517_ ;
	wire _w18516_ ;
	wire _w18515_ ;
	wire _w18514_ ;
	wire _w18513_ ;
	wire _w18512_ ;
	wire _w18511_ ;
	wire _w18510_ ;
	wire _w18509_ ;
	wire _w18508_ ;
	wire _w18507_ ;
	wire _w18506_ ;
	wire _w18505_ ;
	wire _w18504_ ;
	wire _w18503_ ;
	wire _w18502_ ;
	wire _w18501_ ;
	wire _w18500_ ;
	wire _w18499_ ;
	wire _w18498_ ;
	wire _w18497_ ;
	wire _w18496_ ;
	wire _w18495_ ;
	wire _w18494_ ;
	wire _w18493_ ;
	wire _w18492_ ;
	wire _w18491_ ;
	wire _w18490_ ;
	wire _w18489_ ;
	wire _w18488_ ;
	wire _w18487_ ;
	wire _w18486_ ;
	wire _w18485_ ;
	wire _w18484_ ;
	wire _w18483_ ;
	wire _w18482_ ;
	wire _w18481_ ;
	wire _w18480_ ;
	wire _w18479_ ;
	wire _w18478_ ;
	wire _w18477_ ;
	wire _w18476_ ;
	wire _w18475_ ;
	wire _w18474_ ;
	wire _w18473_ ;
	wire _w18472_ ;
	wire _w18471_ ;
	wire _w18470_ ;
	wire _w18469_ ;
	wire _w18468_ ;
	wire _w18467_ ;
	wire _w18466_ ;
	wire _w18465_ ;
	wire _w18464_ ;
	wire _w18463_ ;
	wire _w18462_ ;
	wire _w18461_ ;
	wire _w18460_ ;
	wire _w18459_ ;
	wire _w18458_ ;
	wire _w18457_ ;
	wire _w18456_ ;
	wire _w18455_ ;
	wire _w18454_ ;
	wire _w18453_ ;
	wire _w18452_ ;
	wire _w18451_ ;
	wire _w18450_ ;
	wire _w18449_ ;
	wire _w18448_ ;
	wire _w18447_ ;
	wire _w18446_ ;
	wire _w18445_ ;
	wire _w18444_ ;
	wire _w18443_ ;
	wire _w18442_ ;
	wire _w18441_ ;
	wire _w18440_ ;
	wire _w18439_ ;
	wire _w18438_ ;
	wire _w18437_ ;
	wire _w18436_ ;
	wire _w18435_ ;
	wire _w18434_ ;
	wire _w18433_ ;
	wire _w18432_ ;
	wire _w18431_ ;
	wire _w18430_ ;
	wire _w18429_ ;
	wire _w18428_ ;
	wire _w18427_ ;
	wire _w18426_ ;
	wire _w18425_ ;
	wire _w18424_ ;
	wire _w18423_ ;
	wire _w18422_ ;
	wire _w18421_ ;
	wire _w18420_ ;
	wire _w18419_ ;
	wire _w18418_ ;
	wire _w18417_ ;
	wire _w18416_ ;
	wire _w18415_ ;
	wire _w18414_ ;
	wire _w18413_ ;
	wire _w18412_ ;
	wire _w18411_ ;
	wire _w18410_ ;
	wire _w18409_ ;
	wire _w18408_ ;
	wire _w18407_ ;
	wire _w18406_ ;
	wire _w18405_ ;
	wire _w18404_ ;
	wire _w18403_ ;
	wire _w18402_ ;
	wire _w18401_ ;
	wire _w18400_ ;
	wire _w18399_ ;
	wire _w18398_ ;
	wire _w18397_ ;
	wire _w18396_ ;
	wire _w18395_ ;
	wire _w18394_ ;
	wire _w18393_ ;
	wire _w18392_ ;
	wire _w18391_ ;
	wire _w18390_ ;
	wire _w18389_ ;
	wire _w18388_ ;
	wire _w18387_ ;
	wire _w18386_ ;
	wire _w18385_ ;
	wire _w18384_ ;
	wire _w18383_ ;
	wire _w18382_ ;
	wire _w18381_ ;
	wire _w18380_ ;
	wire _w18379_ ;
	wire _w18378_ ;
	wire _w18377_ ;
	wire _w18376_ ;
	wire _w18375_ ;
	wire _w18374_ ;
	wire _w18373_ ;
	wire _w18372_ ;
	wire _w18371_ ;
	wire _w18370_ ;
	wire _w18369_ ;
	wire _w18368_ ;
	wire _w18367_ ;
	wire _w18366_ ;
	wire _w18365_ ;
	wire _w18364_ ;
	wire _w18363_ ;
	wire _w18362_ ;
	wire _w18361_ ;
	wire _w18360_ ;
	wire _w18359_ ;
	wire _w18358_ ;
	wire _w18357_ ;
	wire _w18356_ ;
	wire _w18355_ ;
	wire _w18354_ ;
	wire _w18353_ ;
	wire _w18352_ ;
	wire _w18351_ ;
	wire _w18350_ ;
	wire _w18349_ ;
	wire _w18348_ ;
	wire _w18347_ ;
	wire _w18346_ ;
	wire _w18345_ ;
	wire _w18344_ ;
	wire _w18343_ ;
	wire _w18342_ ;
	wire _w18341_ ;
	wire _w18340_ ;
	wire _w18339_ ;
	wire _w18338_ ;
	wire _w18337_ ;
	wire _w18336_ ;
	wire _w18335_ ;
	wire _w18334_ ;
	wire _w18333_ ;
	wire _w18332_ ;
	wire _w18331_ ;
	wire _w18330_ ;
	wire _w18329_ ;
	wire _w18328_ ;
	wire _w18327_ ;
	wire _w18326_ ;
	wire _w18325_ ;
	wire _w18324_ ;
	wire _w18323_ ;
	wire _w18322_ ;
	wire _w18321_ ;
	wire _w18320_ ;
	wire _w18319_ ;
	wire _w18318_ ;
	wire _w18317_ ;
	wire _w18316_ ;
	wire _w18315_ ;
	wire _w18314_ ;
	wire _w18313_ ;
	wire _w18312_ ;
	wire _w18311_ ;
	wire _w18310_ ;
	wire _w18309_ ;
	wire _w18308_ ;
	wire _w18307_ ;
	wire _w18306_ ;
	wire _w18305_ ;
	wire _w18304_ ;
	wire _w18303_ ;
	wire _w18302_ ;
	wire _w18301_ ;
	wire _w18300_ ;
	wire _w18299_ ;
	wire _w18298_ ;
	wire _w18297_ ;
	wire _w18296_ ;
	wire _w18295_ ;
	wire _w18294_ ;
	wire _w18293_ ;
	wire _w18292_ ;
	wire _w18291_ ;
	wire _w18290_ ;
	wire _w18289_ ;
	wire _w18288_ ;
	wire _w18287_ ;
	wire _w18286_ ;
	wire _w18285_ ;
	wire _w18284_ ;
	wire _w18283_ ;
	wire _w18282_ ;
	wire _w18281_ ;
	wire _w18280_ ;
	wire _w18279_ ;
	wire _w18278_ ;
	wire _w18277_ ;
	wire _w18276_ ;
	wire _w18275_ ;
	wire _w18274_ ;
	wire _w18273_ ;
	wire _w18272_ ;
	wire _w18271_ ;
	wire _w18270_ ;
	wire _w18269_ ;
	wire _w18268_ ;
	wire _w18267_ ;
	wire _w18266_ ;
	wire _w18265_ ;
	wire _w18264_ ;
	wire _w18263_ ;
	wire _w18262_ ;
	wire _w18261_ ;
	wire _w18260_ ;
	wire _w18259_ ;
	wire _w18258_ ;
	wire _w18257_ ;
	wire _w18256_ ;
	wire _w18255_ ;
	wire _w18254_ ;
	wire _w18253_ ;
	wire _w18252_ ;
	wire _w18251_ ;
	wire _w18250_ ;
	wire _w18249_ ;
	wire _w18248_ ;
	wire _w18247_ ;
	wire _w18246_ ;
	wire _w18245_ ;
	wire _w18244_ ;
	wire _w18243_ ;
	wire _w18242_ ;
	wire _w18241_ ;
	wire _w18240_ ;
	wire _w18239_ ;
	wire _w18238_ ;
	wire _w18237_ ;
	wire _w18236_ ;
	wire _w18235_ ;
	wire _w18234_ ;
	wire _w18233_ ;
	wire _w18232_ ;
	wire _w18231_ ;
	wire _w18230_ ;
	wire _w18229_ ;
	wire _w18228_ ;
	wire _w18227_ ;
	wire _w18226_ ;
	wire _w18225_ ;
	wire _w18224_ ;
	wire _w18223_ ;
	wire _w18222_ ;
	wire _w18221_ ;
	wire _w18220_ ;
	wire _w18219_ ;
	wire _w18218_ ;
	wire _w18217_ ;
	wire _w18216_ ;
	wire _w18215_ ;
	wire _w18214_ ;
	wire _w18213_ ;
	wire _w18212_ ;
	wire _w18211_ ;
	wire _w18210_ ;
	wire _w18209_ ;
	wire _w18208_ ;
	wire _w18207_ ;
	wire _w18206_ ;
	wire _w18205_ ;
	wire _w18204_ ;
	wire _w18203_ ;
	wire _w18202_ ;
	wire _w18201_ ;
	wire _w18200_ ;
	wire _w18199_ ;
	wire _w18198_ ;
	wire _w18197_ ;
	wire _w18196_ ;
	wire _w18195_ ;
	wire _w18194_ ;
	wire _w18193_ ;
	wire _w18192_ ;
	wire _w18191_ ;
	wire _w18190_ ;
	wire _w18189_ ;
	wire _w18188_ ;
	wire _w18187_ ;
	wire _w18186_ ;
	wire _w18185_ ;
	wire _w18184_ ;
	wire _w18183_ ;
	wire _w18182_ ;
	wire _w18181_ ;
	wire _w18180_ ;
	wire _w18179_ ;
	wire _w18178_ ;
	wire _w18177_ ;
	wire _w18176_ ;
	wire _w18175_ ;
	wire _w18174_ ;
	wire _w18173_ ;
	wire _w18172_ ;
	wire _w18171_ ;
	wire _w18170_ ;
	wire _w18169_ ;
	wire _w18168_ ;
	wire _w18167_ ;
	wire _w18166_ ;
	wire _w18165_ ;
	wire _w18164_ ;
	wire _w18163_ ;
	wire _w18162_ ;
	wire _w18161_ ;
	wire _w18160_ ;
	wire _w18159_ ;
	wire _w18158_ ;
	wire _w18157_ ;
	wire _w18156_ ;
	wire _w18155_ ;
	wire _w18154_ ;
	wire _w18153_ ;
	wire _w18152_ ;
	wire _w18151_ ;
	wire _w18150_ ;
	wire _w18149_ ;
	wire _w18148_ ;
	wire _w18147_ ;
	wire _w18146_ ;
	wire _w18145_ ;
	wire _w18144_ ;
	wire _w18143_ ;
	wire _w18142_ ;
	wire _w18141_ ;
	wire _w18140_ ;
	wire _w18139_ ;
	wire _w18138_ ;
	wire _w18137_ ;
	wire _w18136_ ;
	wire _w18135_ ;
	wire _w18134_ ;
	wire _w18133_ ;
	wire _w18132_ ;
	wire _w18131_ ;
	wire _w18130_ ;
	wire _w18129_ ;
	wire _w18128_ ;
	wire _w18127_ ;
	wire _w18126_ ;
	wire _w18125_ ;
	wire _w18124_ ;
	wire _w18123_ ;
	wire _w18122_ ;
	wire _w18121_ ;
	wire _w18120_ ;
	wire _w18119_ ;
	wire _w18118_ ;
	wire _w18117_ ;
	wire _w18116_ ;
	wire _w18115_ ;
	wire _w18114_ ;
	wire _w18113_ ;
	wire _w18112_ ;
	wire _w18111_ ;
	wire _w18110_ ;
	wire _w18109_ ;
	wire _w18108_ ;
	wire _w18107_ ;
	wire _w18106_ ;
	wire _w18105_ ;
	wire _w18104_ ;
	wire _w18103_ ;
	wire _w18102_ ;
	wire _w18101_ ;
	wire _w18100_ ;
	wire _w18099_ ;
	wire _w18098_ ;
	wire _w18097_ ;
	wire _w18096_ ;
	wire _w18095_ ;
	wire _w18094_ ;
	wire _w18093_ ;
	wire _w18092_ ;
	wire _w18091_ ;
	wire _w18090_ ;
	wire _w18089_ ;
	wire _w18088_ ;
	wire _w18087_ ;
	wire _w18086_ ;
	wire _w18085_ ;
	wire _w18084_ ;
	wire _w18083_ ;
	wire _w18082_ ;
	wire _w18081_ ;
	wire _w18080_ ;
	wire _w18079_ ;
	wire _w18078_ ;
	wire _w18077_ ;
	wire _w18076_ ;
	wire _w18075_ ;
	wire _w18074_ ;
	wire _w18073_ ;
	wire _w18072_ ;
	wire _w18071_ ;
	wire _w18070_ ;
	wire _w18069_ ;
	wire _w18068_ ;
	wire _w18067_ ;
	wire _w18066_ ;
	wire _w18065_ ;
	wire _w18064_ ;
	wire _w18063_ ;
	wire _w18062_ ;
	wire _w18061_ ;
	wire _w18060_ ;
	wire _w18059_ ;
	wire _w18058_ ;
	wire _w18057_ ;
	wire _w18056_ ;
	wire _w18055_ ;
	wire _w18054_ ;
	wire _w18053_ ;
	wire _w18052_ ;
	wire _w18051_ ;
	wire _w18050_ ;
	wire _w18049_ ;
	wire _w18048_ ;
	wire _w18047_ ;
	wire _w18046_ ;
	wire _w18045_ ;
	wire _w18044_ ;
	wire _w18043_ ;
	wire _w18042_ ;
	wire _w18041_ ;
	wire _w18040_ ;
	wire _w18039_ ;
	wire _w18038_ ;
	wire _w18037_ ;
	wire _w18036_ ;
	wire _w18035_ ;
	wire _w18034_ ;
	wire _w18033_ ;
	wire _w18032_ ;
	wire _w18031_ ;
	wire _w18030_ ;
	wire _w18029_ ;
	wire _w18028_ ;
	wire _w18027_ ;
	wire _w18026_ ;
	wire _w18025_ ;
	wire _w18024_ ;
	wire _w18023_ ;
	wire _w18022_ ;
	wire _w18021_ ;
	wire _w18020_ ;
	wire _w18019_ ;
	wire _w18018_ ;
	wire _w18017_ ;
	wire _w18016_ ;
	wire _w18015_ ;
	wire _w18014_ ;
	wire _w18013_ ;
	wire _w18012_ ;
	wire _w18011_ ;
	wire _w18010_ ;
	wire _w18009_ ;
	wire _w18008_ ;
	wire _w18007_ ;
	wire _w18006_ ;
	wire _w18005_ ;
	wire _w18004_ ;
	wire _w18003_ ;
	wire _w18002_ ;
	wire _w18001_ ;
	wire _w18000_ ;
	wire _w17999_ ;
	wire _w17998_ ;
	wire _w17997_ ;
	wire _w17996_ ;
	wire _w17995_ ;
	wire _w17994_ ;
	wire _w17993_ ;
	wire _w17992_ ;
	wire _w17991_ ;
	wire _w17990_ ;
	wire _w17989_ ;
	wire _w17988_ ;
	wire _w17987_ ;
	wire _w17986_ ;
	wire _w17985_ ;
	wire _w17984_ ;
	wire _w17983_ ;
	wire _w17982_ ;
	wire _w17981_ ;
	wire _w17980_ ;
	wire _w17979_ ;
	wire _w17978_ ;
	wire _w17977_ ;
	wire _w17976_ ;
	wire _w17975_ ;
	wire _w17974_ ;
	wire _w17973_ ;
	wire _w17972_ ;
	wire _w17971_ ;
	wire _w17970_ ;
	wire _w17969_ ;
	wire _w17968_ ;
	wire _w17967_ ;
	wire _w17966_ ;
	wire _w17965_ ;
	wire _w17964_ ;
	wire _w17963_ ;
	wire _w17962_ ;
	wire _w17961_ ;
	wire _w17960_ ;
	wire _w17959_ ;
	wire _w17958_ ;
	wire _w17957_ ;
	wire _w17956_ ;
	wire _w17955_ ;
	wire _w17954_ ;
	wire _w17953_ ;
	wire _w17952_ ;
	wire _w17951_ ;
	wire _w17950_ ;
	wire _w17949_ ;
	wire _w17948_ ;
	wire _w17947_ ;
	wire _w17946_ ;
	wire _w17945_ ;
	wire _w17944_ ;
	wire _w17943_ ;
	wire _w17942_ ;
	wire _w17941_ ;
	wire _w17940_ ;
	wire _w17939_ ;
	wire _w17938_ ;
	wire _w17937_ ;
	wire _w17936_ ;
	wire _w17935_ ;
	wire _w17934_ ;
	wire _w17933_ ;
	wire _w17932_ ;
	wire _w17931_ ;
	wire _w17930_ ;
	wire _w17929_ ;
	wire _w17928_ ;
	wire _w17927_ ;
	wire _w17926_ ;
	wire _w17925_ ;
	wire _w17924_ ;
	wire _w17923_ ;
	wire _w17922_ ;
	wire _w17921_ ;
	wire _w17920_ ;
	wire _w17919_ ;
	wire _w17918_ ;
	wire _w17917_ ;
	wire _w17916_ ;
	wire _w17915_ ;
	wire _w17914_ ;
	wire _w17913_ ;
	wire _w17912_ ;
	wire _w17911_ ;
	wire _w17910_ ;
	wire _w17909_ ;
	wire _w17908_ ;
	wire _w17907_ ;
	wire _w17906_ ;
	wire _w17905_ ;
	wire _w17904_ ;
	wire _w17903_ ;
	wire _w17902_ ;
	wire _w17901_ ;
	wire _w17900_ ;
	wire _w17899_ ;
	wire _w17898_ ;
	wire _w17897_ ;
	wire _w17896_ ;
	wire _w17895_ ;
	wire _w17894_ ;
	wire _w17893_ ;
	wire _w17892_ ;
	wire _w17891_ ;
	wire _w17890_ ;
	wire _w17889_ ;
	wire _w17888_ ;
	wire _w17887_ ;
	wire _w17886_ ;
	wire _w17885_ ;
	wire _w17884_ ;
	wire _w17883_ ;
	wire _w17882_ ;
	wire _w17881_ ;
	wire _w17880_ ;
	wire _w17879_ ;
	wire _w17878_ ;
	wire _w17877_ ;
	wire _w17876_ ;
	wire _w17875_ ;
	wire _w17874_ ;
	wire _w17873_ ;
	wire _w17872_ ;
	wire _w17871_ ;
	wire _w17870_ ;
	wire _w17869_ ;
	wire _w17868_ ;
	wire _w17867_ ;
	wire _w17866_ ;
	wire _w17865_ ;
	wire _w17864_ ;
	wire _w17863_ ;
	wire _w17862_ ;
	wire _w17861_ ;
	wire _w17860_ ;
	wire _w17859_ ;
	wire _w17858_ ;
	wire _w17857_ ;
	wire _w17856_ ;
	wire _w17855_ ;
	wire _w17854_ ;
	wire _w17853_ ;
	wire _w17852_ ;
	wire _w17851_ ;
	wire _w17850_ ;
	wire _w17849_ ;
	wire _w17848_ ;
	wire _w17847_ ;
	wire _w17846_ ;
	wire _w17845_ ;
	wire _w17844_ ;
	wire _w17843_ ;
	wire _w17842_ ;
	wire _w17841_ ;
	wire _w17840_ ;
	wire _w17839_ ;
	wire _w17838_ ;
	wire _w17837_ ;
	wire _w17836_ ;
	wire _w17835_ ;
	wire _w17834_ ;
	wire _w17833_ ;
	wire _w17832_ ;
	wire _w17831_ ;
	wire _w17830_ ;
	wire _w17829_ ;
	wire _w17828_ ;
	wire _w17827_ ;
	wire _w17826_ ;
	wire _w17825_ ;
	wire _w17824_ ;
	wire _w17823_ ;
	wire _w17822_ ;
	wire _w17821_ ;
	wire _w17820_ ;
	wire _w17819_ ;
	wire _w17818_ ;
	wire _w17817_ ;
	wire _w17816_ ;
	wire _w17815_ ;
	wire _w17814_ ;
	wire _w17813_ ;
	wire _w17812_ ;
	wire _w17811_ ;
	wire _w17810_ ;
	wire _w17809_ ;
	wire _w17808_ ;
	wire _w17807_ ;
	wire _w17806_ ;
	wire _w17805_ ;
	wire _w17804_ ;
	wire _w17803_ ;
	wire _w17802_ ;
	wire _w17801_ ;
	wire _w17800_ ;
	wire _w17799_ ;
	wire _w17798_ ;
	wire _w17797_ ;
	wire _w17796_ ;
	wire _w17795_ ;
	wire _w17794_ ;
	wire _w17793_ ;
	wire _w17792_ ;
	wire _w17791_ ;
	wire _w17790_ ;
	wire _w17789_ ;
	wire _w17788_ ;
	wire _w17787_ ;
	wire _w17786_ ;
	wire _w17785_ ;
	wire _w17784_ ;
	wire _w17783_ ;
	wire _w17782_ ;
	wire _w17781_ ;
	wire _w17780_ ;
	wire _w17779_ ;
	wire _w17778_ ;
	wire _w17777_ ;
	wire _w17776_ ;
	wire _w17775_ ;
	wire _w17774_ ;
	wire _w17773_ ;
	wire _w17772_ ;
	wire _w17771_ ;
	wire _w17770_ ;
	wire _w17769_ ;
	wire _w17768_ ;
	wire _w17767_ ;
	wire _w17766_ ;
	wire _w17765_ ;
	wire _w17764_ ;
	wire _w17763_ ;
	wire _w17762_ ;
	wire _w17761_ ;
	wire _w17760_ ;
	wire _w17759_ ;
	wire _w17758_ ;
	wire _w17757_ ;
	wire _w17756_ ;
	wire _w17755_ ;
	wire _w17754_ ;
	wire _w17753_ ;
	wire _w17752_ ;
	wire _w17751_ ;
	wire _w17750_ ;
	wire _w17749_ ;
	wire _w17748_ ;
	wire _w17747_ ;
	wire _w17746_ ;
	wire _w17745_ ;
	wire _w17744_ ;
	wire _w17743_ ;
	wire _w17742_ ;
	wire _w17741_ ;
	wire _w17740_ ;
	wire _w17739_ ;
	wire _w17738_ ;
	wire _w17737_ ;
	wire _w17736_ ;
	wire _w17735_ ;
	wire _w17734_ ;
	wire _w17733_ ;
	wire _w17732_ ;
	wire _w17731_ ;
	wire _w17730_ ;
	wire _w17729_ ;
	wire _w17728_ ;
	wire _w17727_ ;
	wire _w17726_ ;
	wire _w17725_ ;
	wire _w17724_ ;
	wire _w17723_ ;
	wire _w17722_ ;
	wire _w17721_ ;
	wire _w17720_ ;
	wire _w17719_ ;
	wire _w17718_ ;
	wire _w17717_ ;
	wire _w17716_ ;
	wire _w17715_ ;
	wire _w17714_ ;
	wire _w17713_ ;
	wire _w17712_ ;
	wire _w17711_ ;
	wire _w17710_ ;
	wire _w17709_ ;
	wire _w17708_ ;
	wire _w17707_ ;
	wire _w17706_ ;
	wire _w17705_ ;
	wire _w17704_ ;
	wire _w17703_ ;
	wire _w17702_ ;
	wire _w17701_ ;
	wire _w17700_ ;
	wire _w17699_ ;
	wire _w17698_ ;
	wire _w17697_ ;
	wire _w17696_ ;
	wire _w17695_ ;
	wire _w17694_ ;
	wire _w17693_ ;
	wire _w17692_ ;
	wire _w17691_ ;
	wire _w17690_ ;
	wire _w17689_ ;
	wire _w17688_ ;
	wire _w17687_ ;
	wire _w17686_ ;
	wire _w17685_ ;
	wire _w17684_ ;
	wire _w17683_ ;
	wire _w17682_ ;
	wire _w17681_ ;
	wire _w17680_ ;
	wire _w17679_ ;
	wire _w17678_ ;
	wire _w17677_ ;
	wire _w17676_ ;
	wire _w17675_ ;
	wire _w17674_ ;
	wire _w17673_ ;
	wire _w17672_ ;
	wire _w17671_ ;
	wire _w17670_ ;
	wire _w17669_ ;
	wire _w17668_ ;
	wire _w17667_ ;
	wire _w17666_ ;
	wire _w17665_ ;
	wire _w17664_ ;
	wire _w17663_ ;
	wire _w17662_ ;
	wire _w17661_ ;
	wire _w17660_ ;
	wire _w17659_ ;
	wire _w17658_ ;
	wire _w17657_ ;
	wire _w17656_ ;
	wire _w17655_ ;
	wire _w17654_ ;
	wire _w17653_ ;
	wire _w17652_ ;
	wire _w17651_ ;
	wire _w17650_ ;
	wire _w17649_ ;
	wire _w17648_ ;
	wire _w17647_ ;
	wire _w17646_ ;
	wire _w17645_ ;
	wire _w17644_ ;
	wire _w17643_ ;
	wire _w17642_ ;
	wire _w17641_ ;
	wire _w17640_ ;
	wire _w17639_ ;
	wire _w17638_ ;
	wire _w17637_ ;
	wire _w17636_ ;
	wire _w17635_ ;
	wire _w17634_ ;
	wire _w17633_ ;
	wire _w17632_ ;
	wire _w17631_ ;
	wire _w17630_ ;
	wire _w17629_ ;
	wire _w17628_ ;
	wire _w17627_ ;
	wire _w17626_ ;
	wire _w17625_ ;
	wire _w17624_ ;
	wire _w17623_ ;
	wire _w17622_ ;
	wire _w17621_ ;
	wire _w17620_ ;
	wire _w17619_ ;
	wire _w17618_ ;
	wire _w17617_ ;
	wire _w17616_ ;
	wire _w17615_ ;
	wire _w17614_ ;
	wire _w17613_ ;
	wire _w17612_ ;
	wire _w17611_ ;
	wire _w17610_ ;
	wire _w17609_ ;
	wire _w17608_ ;
	wire _w17607_ ;
	wire _w17606_ ;
	wire _w17605_ ;
	wire _w17604_ ;
	wire _w17603_ ;
	wire _w17602_ ;
	wire _w17601_ ;
	wire _w17600_ ;
	wire _w17599_ ;
	wire _w17598_ ;
	wire _w17597_ ;
	wire _w17596_ ;
	wire _w17595_ ;
	wire _w17594_ ;
	wire _w17593_ ;
	wire _w17592_ ;
	wire _w17591_ ;
	wire _w17590_ ;
	wire _w17589_ ;
	wire _w17588_ ;
	wire _w17587_ ;
	wire _w17586_ ;
	wire _w17585_ ;
	wire _w17584_ ;
	wire _w17583_ ;
	wire _w17582_ ;
	wire _w17581_ ;
	wire _w17580_ ;
	wire _w17579_ ;
	wire _w17578_ ;
	wire _w17577_ ;
	wire _w17576_ ;
	wire _w17575_ ;
	wire _w17574_ ;
	wire _w17573_ ;
	wire _w17572_ ;
	wire _w17571_ ;
	wire _w17570_ ;
	wire _w17569_ ;
	wire _w17568_ ;
	wire _w17567_ ;
	wire _w17566_ ;
	wire _w17565_ ;
	wire _w17564_ ;
	wire _w17563_ ;
	wire _w17562_ ;
	wire _w17561_ ;
	wire _w17560_ ;
	wire _w17559_ ;
	wire _w17558_ ;
	wire _w17557_ ;
	wire _w17556_ ;
	wire _w17555_ ;
	wire _w17554_ ;
	wire _w17553_ ;
	wire _w17552_ ;
	wire _w17551_ ;
	wire _w17550_ ;
	wire _w17549_ ;
	wire _w17548_ ;
	wire _w17547_ ;
	wire _w17546_ ;
	wire _w17545_ ;
	wire _w17544_ ;
	wire _w17543_ ;
	wire _w17542_ ;
	wire _w17541_ ;
	wire _w17540_ ;
	wire _w17539_ ;
	wire _w17538_ ;
	wire _w17537_ ;
	wire _w17536_ ;
	wire _w17535_ ;
	wire _w17534_ ;
	wire _w17533_ ;
	wire _w17532_ ;
	wire _w17531_ ;
	wire _w17530_ ;
	wire _w17529_ ;
	wire _w17528_ ;
	wire _w17527_ ;
	wire _w17526_ ;
	wire _w17525_ ;
	wire _w17524_ ;
	wire _w17523_ ;
	wire _w17522_ ;
	wire _w17521_ ;
	wire _w17520_ ;
	wire _w17519_ ;
	wire _w17518_ ;
	wire _w17517_ ;
	wire _w17516_ ;
	wire _w17515_ ;
	wire _w17514_ ;
	wire _w17513_ ;
	wire _w17512_ ;
	wire _w17511_ ;
	wire _w17510_ ;
	wire _w17509_ ;
	wire _w17508_ ;
	wire _w17507_ ;
	wire _w17506_ ;
	wire _w17505_ ;
	wire _w17504_ ;
	wire _w17503_ ;
	wire _w17502_ ;
	wire _w17501_ ;
	wire _w17500_ ;
	wire _w17499_ ;
	wire _w17498_ ;
	wire _w17497_ ;
	wire _w17496_ ;
	wire _w17495_ ;
	wire _w17494_ ;
	wire _w17493_ ;
	wire _w17492_ ;
	wire _w17491_ ;
	wire _w17490_ ;
	wire _w17489_ ;
	wire _w17488_ ;
	wire _w17487_ ;
	wire _w17486_ ;
	wire _w17485_ ;
	wire _w17484_ ;
	wire _w17483_ ;
	wire _w17482_ ;
	wire _w17481_ ;
	wire _w17480_ ;
	wire _w17479_ ;
	wire _w17478_ ;
	wire _w17477_ ;
	wire _w17476_ ;
	wire _w17475_ ;
	wire _w17474_ ;
	wire _w17473_ ;
	wire _w17472_ ;
	wire _w17471_ ;
	wire _w17470_ ;
	wire _w17469_ ;
	wire _w17468_ ;
	wire _w17467_ ;
	wire _w17466_ ;
	wire _w17465_ ;
	wire _w17464_ ;
	wire _w17463_ ;
	wire _w17462_ ;
	wire _w17461_ ;
	wire _w17460_ ;
	wire _w17459_ ;
	wire _w17458_ ;
	wire _w17457_ ;
	wire _w17456_ ;
	wire _w17455_ ;
	wire _w17454_ ;
	wire _w17453_ ;
	wire _w17452_ ;
	wire _w17451_ ;
	wire _w17450_ ;
	wire _w17449_ ;
	wire _w17448_ ;
	wire _w17447_ ;
	wire _w17446_ ;
	wire _w17445_ ;
	wire _w17444_ ;
	wire _w17443_ ;
	wire _w17442_ ;
	wire _w17441_ ;
	wire _w17440_ ;
	wire _w17439_ ;
	wire _w17438_ ;
	wire _w17437_ ;
	wire _w17436_ ;
	wire _w17435_ ;
	wire _w17434_ ;
	wire _w17433_ ;
	wire _w17432_ ;
	wire _w17431_ ;
	wire _w17430_ ;
	wire _w17429_ ;
	wire _w17428_ ;
	wire _w17427_ ;
	wire _w17426_ ;
	wire _w17425_ ;
	wire _w17424_ ;
	wire _w17423_ ;
	wire _w17422_ ;
	wire _w17421_ ;
	wire _w17420_ ;
	wire _w17419_ ;
	wire _w17418_ ;
	wire _w17417_ ;
	wire _w17416_ ;
	wire _w17415_ ;
	wire _w17414_ ;
	wire _w17413_ ;
	wire _w17412_ ;
	wire _w17411_ ;
	wire _w17410_ ;
	wire _w17409_ ;
	wire _w17408_ ;
	wire _w17407_ ;
	wire _w17406_ ;
	wire _w17405_ ;
	wire _w17404_ ;
	wire _w17403_ ;
	wire _w17402_ ;
	wire _w17401_ ;
	wire _w17400_ ;
	wire _w17399_ ;
	wire _w17398_ ;
	wire _w17397_ ;
	wire _w17396_ ;
	wire _w17395_ ;
	wire _w17394_ ;
	wire _w17393_ ;
	wire _w17392_ ;
	wire _w17391_ ;
	wire _w17390_ ;
	wire _w17389_ ;
	wire _w17388_ ;
	wire _w17387_ ;
	wire _w17386_ ;
	wire _w17385_ ;
	wire _w17384_ ;
	wire _w17383_ ;
	wire _w17382_ ;
	wire _w17381_ ;
	wire _w17380_ ;
	wire _w17379_ ;
	wire _w17378_ ;
	wire _w17377_ ;
	wire _w17376_ ;
	wire _w17375_ ;
	wire _w17374_ ;
	wire _w17373_ ;
	wire _w17372_ ;
	wire _w17371_ ;
	wire _w17370_ ;
	wire _w17369_ ;
	wire _w17368_ ;
	wire _w17367_ ;
	wire _w17366_ ;
	wire _w17365_ ;
	wire _w17364_ ;
	wire _w17363_ ;
	wire _w17362_ ;
	wire _w17361_ ;
	wire _w17360_ ;
	wire _w17359_ ;
	wire _w17358_ ;
	wire _w17357_ ;
	wire _w17356_ ;
	wire _w17355_ ;
	wire _w17354_ ;
	wire _w17353_ ;
	wire _w17352_ ;
	wire _w17351_ ;
	wire _w17350_ ;
	wire _w17349_ ;
	wire _w17348_ ;
	wire _w17347_ ;
	wire _w17346_ ;
	wire _w17345_ ;
	wire _w17344_ ;
	wire _w17343_ ;
	wire _w17342_ ;
	wire _w17341_ ;
	wire _w17340_ ;
	wire _w17339_ ;
	wire _w17338_ ;
	wire _w17337_ ;
	wire _w17336_ ;
	wire _w17335_ ;
	wire _w17334_ ;
	wire _w17333_ ;
	wire _w17332_ ;
	wire _w17331_ ;
	wire _w17330_ ;
	wire _w17329_ ;
	wire _w17328_ ;
	wire _w17327_ ;
	wire _w17326_ ;
	wire _w17325_ ;
	wire _w17324_ ;
	wire _w17323_ ;
	wire _w17322_ ;
	wire _w17321_ ;
	wire _w17320_ ;
	wire _w17319_ ;
	wire _w17318_ ;
	wire _w17317_ ;
	wire _w17316_ ;
	wire _w17315_ ;
	wire _w17314_ ;
	wire _w17313_ ;
	wire _w17312_ ;
	wire _w17311_ ;
	wire _w17310_ ;
	wire _w17309_ ;
	wire _w17308_ ;
	wire _w17307_ ;
	wire _w17306_ ;
	wire _w17305_ ;
	wire _w17304_ ;
	wire _w17303_ ;
	wire _w17302_ ;
	wire _w17301_ ;
	wire _w17300_ ;
	wire _w17299_ ;
	wire _w17298_ ;
	wire _w17297_ ;
	wire _w17296_ ;
	wire _w17295_ ;
	wire _w17294_ ;
	wire _w17293_ ;
	wire _w17292_ ;
	wire _w17291_ ;
	wire _w17290_ ;
	wire _w17289_ ;
	wire _w17288_ ;
	wire _w17287_ ;
	wire _w17286_ ;
	wire _w17285_ ;
	wire _w17284_ ;
	wire _w17283_ ;
	wire _w17282_ ;
	wire _w17281_ ;
	wire _w17280_ ;
	wire _w17279_ ;
	wire _w17278_ ;
	wire _w17277_ ;
	wire _w17276_ ;
	wire _w17275_ ;
	wire _w17274_ ;
	wire _w17273_ ;
	wire _w17272_ ;
	wire _w17271_ ;
	wire _w17270_ ;
	wire _w17269_ ;
	wire _w17268_ ;
	wire _w17267_ ;
	wire _w17266_ ;
	wire _w17265_ ;
	wire _w17264_ ;
	wire _w17263_ ;
	wire _w17262_ ;
	wire _w17261_ ;
	wire _w17260_ ;
	wire _w17259_ ;
	wire _w17258_ ;
	wire _w17257_ ;
	wire _w17256_ ;
	wire _w17255_ ;
	wire _w17254_ ;
	wire _w17253_ ;
	wire _w17252_ ;
	wire _w17251_ ;
	wire _w17250_ ;
	wire _w17249_ ;
	wire _w17248_ ;
	wire _w17247_ ;
	wire _w17246_ ;
	wire _w17245_ ;
	wire _w17244_ ;
	wire _w17243_ ;
	wire _w17242_ ;
	wire _w17241_ ;
	wire _w17240_ ;
	wire _w17239_ ;
	wire _w17238_ ;
	wire _w17237_ ;
	wire _w17236_ ;
	wire _w17235_ ;
	wire _w17234_ ;
	wire _w17233_ ;
	wire _w17232_ ;
	wire _w17231_ ;
	wire _w17230_ ;
	wire _w17229_ ;
	wire _w17228_ ;
	wire _w17227_ ;
	wire _w17226_ ;
	wire _w17225_ ;
	wire _w17224_ ;
	wire _w17223_ ;
	wire _w17222_ ;
	wire _w17221_ ;
	wire _w17220_ ;
	wire _w17219_ ;
	wire _w17218_ ;
	wire _w17217_ ;
	wire _w17216_ ;
	wire _w17215_ ;
	wire _w17214_ ;
	wire _w17213_ ;
	wire _w17212_ ;
	wire _w17211_ ;
	wire _w17210_ ;
	wire _w17209_ ;
	wire _w17208_ ;
	wire _w17207_ ;
	wire _w17206_ ;
	wire _w17205_ ;
	wire _w17204_ ;
	wire _w17203_ ;
	wire _w17202_ ;
	wire _w17201_ ;
	wire _w17200_ ;
	wire _w17199_ ;
	wire _w17198_ ;
	wire _w17197_ ;
	wire _w17196_ ;
	wire _w17195_ ;
	wire _w17194_ ;
	wire _w17193_ ;
	wire _w17192_ ;
	wire _w17191_ ;
	wire _w17190_ ;
	wire _w17189_ ;
	wire _w17188_ ;
	wire _w17187_ ;
	wire _w17186_ ;
	wire _w17185_ ;
	wire _w17184_ ;
	wire _w17183_ ;
	wire _w17182_ ;
	wire _w17181_ ;
	wire _w17180_ ;
	wire _w17179_ ;
	wire _w17178_ ;
	wire _w17177_ ;
	wire _w17176_ ;
	wire _w17175_ ;
	wire _w17174_ ;
	wire _w17173_ ;
	wire _w17172_ ;
	wire _w17171_ ;
	wire _w17170_ ;
	wire _w17169_ ;
	wire _w17168_ ;
	wire _w17167_ ;
	wire _w17166_ ;
	wire _w17165_ ;
	wire _w17164_ ;
	wire _w17163_ ;
	wire _w17162_ ;
	wire _w17161_ ;
	wire _w17160_ ;
	wire _w17159_ ;
	wire _w17158_ ;
	wire _w17157_ ;
	wire _w17156_ ;
	wire _w17155_ ;
	wire _w17154_ ;
	wire _w17153_ ;
	wire _w17152_ ;
	wire _w17151_ ;
	wire _w17150_ ;
	wire _w17149_ ;
	wire _w17148_ ;
	wire _w17147_ ;
	wire _w17146_ ;
	wire _w17145_ ;
	wire _w17144_ ;
	wire _w17143_ ;
	wire _w17142_ ;
	wire _w17141_ ;
	wire _w17140_ ;
	wire _w17139_ ;
	wire _w17138_ ;
	wire _w17137_ ;
	wire _w17136_ ;
	wire _w17135_ ;
	wire _w17134_ ;
	wire _w17133_ ;
	wire _w17132_ ;
	wire _w17131_ ;
	wire _w17130_ ;
	wire _w17129_ ;
	wire _w17128_ ;
	wire _w17127_ ;
	wire _w17126_ ;
	wire _w17125_ ;
	wire _w17124_ ;
	wire _w17123_ ;
	wire _w17122_ ;
	wire _w17121_ ;
	wire _w17120_ ;
	wire _w17119_ ;
	wire _w17118_ ;
	wire _w17117_ ;
	wire _w17116_ ;
	wire _w17115_ ;
	wire _w17114_ ;
	wire _w17113_ ;
	wire _w17112_ ;
	wire _w17111_ ;
	wire _w17110_ ;
	wire _w17109_ ;
	wire _w17108_ ;
	wire _w17107_ ;
	wire _w17106_ ;
	wire _w17105_ ;
	wire _w17104_ ;
	wire _w17103_ ;
	wire _w17102_ ;
	wire _w17101_ ;
	wire _w17100_ ;
	wire _w17099_ ;
	wire _w17098_ ;
	wire _w17097_ ;
	wire _w17096_ ;
	wire _w17095_ ;
	wire _w17094_ ;
	wire _w17093_ ;
	wire _w17092_ ;
	wire _w17091_ ;
	wire _w17090_ ;
	wire _w17089_ ;
	wire _w17088_ ;
	wire _w17087_ ;
	wire _w17086_ ;
	wire _w17085_ ;
	wire _w17084_ ;
	wire _w17083_ ;
	wire _w17082_ ;
	wire _w17081_ ;
	wire _w17080_ ;
	wire _w17079_ ;
	wire _w17078_ ;
	wire _w17077_ ;
	wire _w17076_ ;
	wire _w17075_ ;
	wire _w17074_ ;
	wire _w17073_ ;
	wire _w17072_ ;
	wire _w17071_ ;
	wire _w17070_ ;
	wire _w17069_ ;
	wire _w17068_ ;
	wire _w17067_ ;
	wire _w17066_ ;
	wire _w17065_ ;
	wire _w17064_ ;
	wire _w17063_ ;
	wire _w17062_ ;
	wire _w17061_ ;
	wire _w17060_ ;
	wire _w17059_ ;
	wire _w17058_ ;
	wire _w17057_ ;
	wire _w17056_ ;
	wire _w17055_ ;
	wire _w17054_ ;
	wire _w17053_ ;
	wire _w17052_ ;
	wire _w17051_ ;
	wire _w17050_ ;
	wire _w17049_ ;
	wire _w17048_ ;
	wire _w17047_ ;
	wire _w17046_ ;
	wire _w17045_ ;
	wire _w17044_ ;
	wire _w17043_ ;
	wire _w17042_ ;
	wire _w17041_ ;
	wire _w17040_ ;
	wire _w17039_ ;
	wire _w17038_ ;
	wire _w17037_ ;
	wire _w17036_ ;
	wire _w17035_ ;
	wire _w17034_ ;
	wire _w17033_ ;
	wire _w17032_ ;
	wire _w17031_ ;
	wire _w17030_ ;
	wire _w17029_ ;
	wire _w17028_ ;
	wire _w17027_ ;
	wire _w17026_ ;
	wire _w17025_ ;
	wire _w17024_ ;
	wire _w17023_ ;
	wire _w17022_ ;
	wire _w17021_ ;
	wire _w17020_ ;
	wire _w17019_ ;
	wire _w17018_ ;
	wire _w17017_ ;
	wire _w17016_ ;
	wire _w17015_ ;
	wire _w17014_ ;
	wire _w17013_ ;
	wire _w17012_ ;
	wire _w17011_ ;
	wire _w17010_ ;
	wire _w17009_ ;
	wire _w17008_ ;
	wire _w17007_ ;
	wire _w17006_ ;
	wire _w17005_ ;
	wire _w17004_ ;
	wire _w17003_ ;
	wire _w17002_ ;
	wire _w17001_ ;
	wire _w17000_ ;
	wire _w16999_ ;
	wire _w16998_ ;
	wire _w16997_ ;
	wire _w16996_ ;
	wire _w16995_ ;
	wire _w16994_ ;
	wire _w16993_ ;
	wire _w16992_ ;
	wire _w16991_ ;
	wire _w16990_ ;
	wire _w16989_ ;
	wire _w16988_ ;
	wire _w16987_ ;
	wire _w16986_ ;
	wire _w16985_ ;
	wire _w16984_ ;
	wire _w16983_ ;
	wire _w16982_ ;
	wire _w16981_ ;
	wire _w16980_ ;
	wire _w16979_ ;
	wire _w16978_ ;
	wire _w16977_ ;
	wire _w16976_ ;
	wire _w16975_ ;
	wire _w16974_ ;
	wire _w16973_ ;
	wire _w16972_ ;
	wire _w16971_ ;
	wire _w16970_ ;
	wire _w16969_ ;
	wire _w16968_ ;
	wire _w16967_ ;
	wire _w16966_ ;
	wire _w16965_ ;
	wire _w16964_ ;
	wire _w16963_ ;
	wire _w16962_ ;
	wire _w16961_ ;
	wire _w16960_ ;
	wire _w16959_ ;
	wire _w16958_ ;
	wire _w16957_ ;
	wire _w16956_ ;
	wire _w16955_ ;
	wire _w16954_ ;
	wire _w16953_ ;
	wire _w16952_ ;
	wire _w16951_ ;
	wire _w16950_ ;
	wire _w16949_ ;
	wire _w16948_ ;
	wire _w16947_ ;
	wire _w16946_ ;
	wire _w16945_ ;
	wire _w16944_ ;
	wire _w16943_ ;
	wire _w16942_ ;
	wire _w16941_ ;
	wire _w16940_ ;
	wire _w16939_ ;
	wire _w16938_ ;
	wire _w16937_ ;
	wire _w16936_ ;
	wire _w16935_ ;
	wire _w16934_ ;
	wire _w16933_ ;
	wire _w16932_ ;
	wire _w16931_ ;
	wire _w16930_ ;
	wire _w16929_ ;
	wire _w16928_ ;
	wire _w16927_ ;
	wire _w16926_ ;
	wire _w16925_ ;
	wire _w16924_ ;
	wire _w16923_ ;
	wire _w16922_ ;
	wire _w16921_ ;
	wire _w16920_ ;
	wire _w16919_ ;
	wire _w16918_ ;
	wire _w16917_ ;
	wire _w16916_ ;
	wire _w16915_ ;
	wire _w16914_ ;
	wire _w16913_ ;
	wire _w16912_ ;
	wire _w16911_ ;
	wire _w16910_ ;
	wire _w16909_ ;
	wire _w16908_ ;
	wire _w16907_ ;
	wire _w16906_ ;
	wire _w16905_ ;
	wire _w16904_ ;
	wire _w16903_ ;
	wire _w16902_ ;
	wire _w16901_ ;
	wire _w16900_ ;
	wire _w16899_ ;
	wire _w16898_ ;
	wire _w16897_ ;
	wire _w16896_ ;
	wire _w16895_ ;
	wire _w16894_ ;
	wire _w16893_ ;
	wire _w16892_ ;
	wire _w16891_ ;
	wire _w16890_ ;
	wire _w16889_ ;
	wire _w16888_ ;
	wire _w16887_ ;
	wire _w16886_ ;
	wire _w16885_ ;
	wire _w16884_ ;
	wire _w16883_ ;
	wire _w16882_ ;
	wire _w16881_ ;
	wire _w16880_ ;
	wire _w16879_ ;
	wire _w16878_ ;
	wire _w16877_ ;
	wire _w16876_ ;
	wire _w16875_ ;
	wire _w16874_ ;
	wire _w16873_ ;
	wire _w16872_ ;
	wire _w16871_ ;
	wire _w16870_ ;
	wire _w16869_ ;
	wire _w16868_ ;
	wire _w16867_ ;
	wire _w16866_ ;
	wire _w16865_ ;
	wire _w16864_ ;
	wire _w16863_ ;
	wire _w16862_ ;
	wire _w16861_ ;
	wire _w16860_ ;
	wire _w16859_ ;
	wire _w16858_ ;
	wire _w16857_ ;
	wire _w16856_ ;
	wire _w16855_ ;
	wire _w16854_ ;
	wire _w16853_ ;
	wire _w16852_ ;
	wire _w16851_ ;
	wire _w16850_ ;
	wire _w16849_ ;
	wire _w16848_ ;
	wire _w16847_ ;
	wire _w16846_ ;
	wire _w16845_ ;
	wire _w16844_ ;
	wire _w16843_ ;
	wire _w16842_ ;
	wire _w16841_ ;
	wire _w16840_ ;
	wire _w16839_ ;
	wire _w16838_ ;
	wire _w16837_ ;
	wire _w16836_ ;
	wire _w16835_ ;
	wire _w16834_ ;
	wire _w16833_ ;
	wire _w16832_ ;
	wire _w16831_ ;
	wire _w16830_ ;
	wire _w16829_ ;
	wire _w16828_ ;
	wire _w16827_ ;
	wire _w16826_ ;
	wire _w16825_ ;
	wire _w16824_ ;
	wire _w16823_ ;
	wire _w16822_ ;
	wire _w16821_ ;
	wire _w16820_ ;
	wire _w16819_ ;
	wire _w16818_ ;
	wire _w16817_ ;
	wire _w16816_ ;
	wire _w16815_ ;
	wire _w16814_ ;
	wire _w16813_ ;
	wire _w16812_ ;
	wire _w16811_ ;
	wire _w16810_ ;
	wire _w16809_ ;
	wire _w16808_ ;
	wire _w16807_ ;
	wire _w16806_ ;
	wire _w16805_ ;
	wire _w16804_ ;
	wire _w16803_ ;
	wire _w16802_ ;
	wire _w16801_ ;
	wire _w16800_ ;
	wire _w16799_ ;
	wire _w16798_ ;
	wire _w16797_ ;
	wire _w16796_ ;
	wire _w16795_ ;
	wire _w16794_ ;
	wire _w16793_ ;
	wire _w16792_ ;
	wire _w16791_ ;
	wire _w16790_ ;
	wire _w16789_ ;
	wire _w16788_ ;
	wire _w16787_ ;
	wire _w16786_ ;
	wire _w16785_ ;
	wire _w16784_ ;
	wire _w16783_ ;
	wire _w16782_ ;
	wire _w16781_ ;
	wire _w16780_ ;
	wire _w16779_ ;
	wire _w16778_ ;
	wire _w16777_ ;
	wire _w16776_ ;
	wire _w16775_ ;
	wire _w16774_ ;
	wire _w16773_ ;
	wire _w16772_ ;
	wire _w16771_ ;
	wire _w16770_ ;
	wire _w16769_ ;
	wire _w16768_ ;
	wire _w16767_ ;
	wire _w16766_ ;
	wire _w16765_ ;
	wire _w16764_ ;
	wire _w16763_ ;
	wire _w16762_ ;
	wire _w16761_ ;
	wire _w16760_ ;
	wire _w16759_ ;
	wire _w16758_ ;
	wire _w16757_ ;
	wire _w16756_ ;
	wire _w16755_ ;
	wire _w16754_ ;
	wire _w16753_ ;
	wire _w16752_ ;
	wire _w16751_ ;
	wire _w16750_ ;
	wire _w16749_ ;
	wire _w16748_ ;
	wire _w16747_ ;
	wire _w16746_ ;
	wire _w16745_ ;
	wire _w16744_ ;
	wire _w16743_ ;
	wire _w16742_ ;
	wire _w16741_ ;
	wire _w16740_ ;
	wire _w16739_ ;
	wire _w16738_ ;
	wire _w16737_ ;
	wire _w16736_ ;
	wire _w16735_ ;
	wire _w16734_ ;
	wire _w16733_ ;
	wire _w16732_ ;
	wire _w16731_ ;
	wire _w16730_ ;
	wire _w16729_ ;
	wire _w16728_ ;
	wire _w16727_ ;
	wire _w16726_ ;
	wire _w16725_ ;
	wire _w16724_ ;
	wire _w16723_ ;
	wire _w16722_ ;
	wire _w16721_ ;
	wire _w16720_ ;
	wire _w16719_ ;
	wire _w16718_ ;
	wire _w16717_ ;
	wire _w16716_ ;
	wire _w16715_ ;
	wire _w16714_ ;
	wire _w16713_ ;
	wire _w16712_ ;
	wire _w16711_ ;
	wire _w16710_ ;
	wire _w16709_ ;
	wire _w16708_ ;
	wire _w16707_ ;
	wire _w16706_ ;
	wire _w16705_ ;
	wire _w16704_ ;
	wire _w16703_ ;
	wire _w16702_ ;
	wire _w16701_ ;
	wire _w16700_ ;
	wire _w16699_ ;
	wire _w16698_ ;
	wire _w16697_ ;
	wire _w16696_ ;
	wire _w16695_ ;
	wire _w16694_ ;
	wire _w16693_ ;
	wire _w16692_ ;
	wire _w16691_ ;
	wire _w16690_ ;
	wire _w16689_ ;
	wire _w16688_ ;
	wire _w16687_ ;
	wire _w16686_ ;
	wire _w16685_ ;
	wire _w16684_ ;
	wire _w16683_ ;
	wire _w16682_ ;
	wire _w16681_ ;
	wire _w16680_ ;
	wire _w16679_ ;
	wire _w16678_ ;
	wire _w16677_ ;
	wire _w16676_ ;
	wire _w16675_ ;
	wire _w16674_ ;
	wire _w16673_ ;
	wire _w16672_ ;
	wire _w16671_ ;
	wire _w16670_ ;
	wire _w16669_ ;
	wire _w16668_ ;
	wire _w16667_ ;
	wire _w16666_ ;
	wire _w16665_ ;
	wire _w16664_ ;
	wire _w16663_ ;
	wire _w16662_ ;
	wire _w16661_ ;
	wire _w16660_ ;
	wire _w16659_ ;
	wire _w16658_ ;
	wire _w16657_ ;
	wire _w16656_ ;
	wire _w16655_ ;
	wire _w16654_ ;
	wire _w16653_ ;
	wire _w16652_ ;
	wire _w16651_ ;
	wire _w16650_ ;
	wire _w16649_ ;
	wire _w16648_ ;
	wire _w16647_ ;
	wire _w16646_ ;
	wire _w16645_ ;
	wire _w16644_ ;
	wire _w16643_ ;
	wire _w16642_ ;
	wire _w16641_ ;
	wire _w16640_ ;
	wire _w16639_ ;
	wire _w16638_ ;
	wire _w16637_ ;
	wire _w16636_ ;
	wire _w16635_ ;
	wire _w16634_ ;
	wire _w16633_ ;
	wire _w16632_ ;
	wire _w16631_ ;
	wire _w16630_ ;
	wire _w16629_ ;
	wire _w16628_ ;
	wire _w16627_ ;
	wire _w16626_ ;
	wire _w16625_ ;
	wire _w16624_ ;
	wire _w16623_ ;
	wire _w16622_ ;
	wire _w16621_ ;
	wire _w16620_ ;
	wire _w16619_ ;
	wire _w16618_ ;
	wire _w16617_ ;
	wire _w16616_ ;
	wire _w16615_ ;
	wire _w16614_ ;
	wire _w16613_ ;
	wire _w16612_ ;
	wire _w16611_ ;
	wire _w16610_ ;
	wire _w16609_ ;
	wire _w16608_ ;
	wire _w16607_ ;
	wire _w16606_ ;
	wire _w16605_ ;
	wire _w16604_ ;
	wire _w16603_ ;
	wire _w16602_ ;
	wire _w16601_ ;
	wire _w16600_ ;
	wire _w16599_ ;
	wire _w16598_ ;
	wire _w16597_ ;
	wire _w16596_ ;
	wire _w16595_ ;
	wire _w16594_ ;
	wire _w16593_ ;
	wire _w16592_ ;
	wire _w16591_ ;
	wire _w16590_ ;
	wire _w16589_ ;
	wire _w16588_ ;
	wire _w16587_ ;
	wire _w16586_ ;
	wire _w16585_ ;
	wire _w16584_ ;
	wire _w16583_ ;
	wire _w16582_ ;
	wire _w16581_ ;
	wire _w16580_ ;
	wire _w16579_ ;
	wire _w16578_ ;
	wire _w16577_ ;
	wire _w16576_ ;
	wire _w16575_ ;
	wire _w16574_ ;
	wire _w16573_ ;
	wire _w16572_ ;
	wire _w16571_ ;
	wire _w16570_ ;
	wire _w16569_ ;
	wire _w16568_ ;
	wire _w16567_ ;
	wire _w16566_ ;
	wire _w16565_ ;
	wire _w16564_ ;
	wire _w16563_ ;
	wire _w16562_ ;
	wire _w16561_ ;
	wire _w16560_ ;
	wire _w16559_ ;
	wire _w16558_ ;
	wire _w16557_ ;
	wire _w16556_ ;
	wire _w16555_ ;
	wire _w16554_ ;
	wire _w16553_ ;
	wire _w16552_ ;
	wire _w16551_ ;
	wire _w16550_ ;
	wire _w16549_ ;
	wire _w16548_ ;
	wire _w16547_ ;
	wire _w16546_ ;
	wire _w16545_ ;
	wire _w16544_ ;
	wire _w16543_ ;
	wire _w16542_ ;
	wire _w16541_ ;
	wire _w16540_ ;
	wire _w16539_ ;
	wire _w16538_ ;
	wire _w16537_ ;
	wire _w16536_ ;
	wire _w16535_ ;
	wire _w16534_ ;
	wire _w16533_ ;
	wire _w16532_ ;
	wire _w16531_ ;
	wire _w16530_ ;
	wire _w16529_ ;
	wire _w16528_ ;
	wire _w16527_ ;
	wire _w16526_ ;
	wire _w16525_ ;
	wire _w16524_ ;
	wire _w16523_ ;
	wire _w16522_ ;
	wire _w16521_ ;
	wire _w16520_ ;
	wire _w16519_ ;
	wire _w16518_ ;
	wire _w16517_ ;
	wire _w16516_ ;
	wire _w16515_ ;
	wire _w16514_ ;
	wire _w16513_ ;
	wire _w16512_ ;
	wire _w16511_ ;
	wire _w16510_ ;
	wire _w16509_ ;
	wire _w16508_ ;
	wire _w16507_ ;
	wire _w16506_ ;
	wire _w16505_ ;
	wire _w16504_ ;
	wire _w16503_ ;
	wire _w16502_ ;
	wire _w16501_ ;
	wire _w16500_ ;
	wire _w16499_ ;
	wire _w16498_ ;
	wire _w16497_ ;
	wire _w16496_ ;
	wire _w16495_ ;
	wire _w16494_ ;
	wire _w16493_ ;
	wire _w16492_ ;
	wire _w16491_ ;
	wire _w16490_ ;
	wire _w16489_ ;
	wire _w16488_ ;
	wire _w16487_ ;
	wire _w16486_ ;
	wire _w16485_ ;
	wire _w16484_ ;
	wire _w16483_ ;
	wire _w16482_ ;
	wire _w16481_ ;
	wire _w16480_ ;
	wire _w16479_ ;
	wire _w16478_ ;
	wire _w16477_ ;
	wire _w16476_ ;
	wire _w16475_ ;
	wire _w16474_ ;
	wire _w16473_ ;
	wire _w16472_ ;
	wire _w16471_ ;
	wire _w16470_ ;
	wire _w16469_ ;
	wire _w16468_ ;
	wire _w16467_ ;
	wire _w16466_ ;
	wire _w16465_ ;
	wire _w16464_ ;
	wire _w16463_ ;
	wire _w16462_ ;
	wire _w16461_ ;
	wire _w16460_ ;
	wire _w16459_ ;
	wire _w16458_ ;
	wire _w16457_ ;
	wire _w16456_ ;
	wire _w16455_ ;
	wire _w16454_ ;
	wire _w16453_ ;
	wire _w16452_ ;
	wire _w16451_ ;
	wire _w16450_ ;
	wire _w16449_ ;
	wire _w16448_ ;
	wire _w16447_ ;
	wire _w16446_ ;
	wire _w16445_ ;
	wire _w16444_ ;
	wire _w16443_ ;
	wire _w16442_ ;
	wire _w16441_ ;
	wire _w16440_ ;
	wire _w16439_ ;
	wire _w16438_ ;
	wire _w16437_ ;
	wire _w16436_ ;
	wire _w16435_ ;
	wire _w16434_ ;
	wire _w16433_ ;
	wire _w16432_ ;
	wire _w16431_ ;
	wire _w16430_ ;
	wire _w16429_ ;
	wire _w16428_ ;
	wire _w16427_ ;
	wire _w16426_ ;
	wire _w16425_ ;
	wire _w16424_ ;
	wire _w16423_ ;
	wire _w16422_ ;
	wire _w16421_ ;
	wire _w16420_ ;
	wire _w16419_ ;
	wire _w16418_ ;
	wire _w16417_ ;
	wire _w16416_ ;
	wire _w16415_ ;
	wire _w16414_ ;
	wire _w16413_ ;
	wire _w16412_ ;
	wire _w16411_ ;
	wire _w16410_ ;
	wire _w16409_ ;
	wire _w16408_ ;
	wire _w16407_ ;
	wire _w16406_ ;
	wire _w16405_ ;
	wire _w16404_ ;
	wire _w16403_ ;
	wire _w16402_ ;
	wire _w16401_ ;
	wire _w16400_ ;
	wire _w16399_ ;
	wire _w16398_ ;
	wire _w16397_ ;
	wire _w16396_ ;
	wire _w16395_ ;
	wire _w16394_ ;
	wire _w16393_ ;
	wire _w16392_ ;
	wire _w16391_ ;
	wire _w16390_ ;
	wire _w16389_ ;
	wire _w16388_ ;
	wire _w16387_ ;
	wire _w16386_ ;
	wire _w16385_ ;
	wire _w16384_ ;
	wire _w16383_ ;
	wire _w16382_ ;
	wire _w16381_ ;
	wire _w16380_ ;
	wire _w16379_ ;
	wire _w16378_ ;
	wire _w16377_ ;
	wire _w16376_ ;
	wire _w16375_ ;
	wire _w16374_ ;
	wire _w16373_ ;
	wire _w16372_ ;
	wire _w16371_ ;
	wire _w16370_ ;
	wire _w16369_ ;
	wire _w16368_ ;
	wire _w16367_ ;
	wire _w16366_ ;
	wire _w16365_ ;
	wire _w16364_ ;
	wire _w16363_ ;
	wire _w16362_ ;
	wire _w16361_ ;
	wire _w16360_ ;
	wire _w16359_ ;
	wire _w16358_ ;
	wire _w16357_ ;
	wire _w16356_ ;
	wire _w16355_ ;
	wire _w16354_ ;
	wire _w16353_ ;
	wire _w16352_ ;
	wire _w16351_ ;
	wire _w16350_ ;
	wire _w16349_ ;
	wire _w16348_ ;
	wire _w16347_ ;
	wire _w16346_ ;
	wire _w16345_ ;
	wire _w16344_ ;
	wire _w16343_ ;
	wire _w16342_ ;
	wire _w16341_ ;
	wire _w16340_ ;
	wire _w16339_ ;
	wire _w16338_ ;
	wire _w16337_ ;
	wire _w16336_ ;
	wire _w16335_ ;
	wire _w16334_ ;
	wire _w16333_ ;
	wire _w16332_ ;
	wire _w16331_ ;
	wire _w16330_ ;
	wire _w16329_ ;
	wire _w16328_ ;
	wire _w16327_ ;
	wire _w16326_ ;
	wire _w16325_ ;
	wire _w16324_ ;
	wire _w16323_ ;
	wire _w16322_ ;
	wire _w16321_ ;
	wire _w16320_ ;
	wire _w16319_ ;
	wire _w16318_ ;
	wire _w16317_ ;
	wire _w16316_ ;
	wire _w16315_ ;
	wire _w16314_ ;
	wire _w16313_ ;
	wire _w16312_ ;
	wire _w16311_ ;
	wire _w16310_ ;
	wire _w16309_ ;
	wire _w16308_ ;
	wire _w16307_ ;
	wire _w16306_ ;
	wire _w16305_ ;
	wire _w16304_ ;
	wire _w16303_ ;
	wire _w16302_ ;
	wire _w16301_ ;
	wire _w16300_ ;
	wire _w16299_ ;
	wire _w16298_ ;
	wire _w16297_ ;
	wire _w16296_ ;
	wire _w16295_ ;
	wire _w16294_ ;
	wire _w16293_ ;
	wire _w16292_ ;
	wire _w16291_ ;
	wire _w16290_ ;
	wire _w16289_ ;
	wire _w16288_ ;
	wire _w16287_ ;
	wire _w16286_ ;
	wire _w16285_ ;
	wire _w16284_ ;
	wire _w16283_ ;
	wire _w16282_ ;
	wire _w16281_ ;
	wire _w16280_ ;
	wire _w16279_ ;
	wire _w16278_ ;
	wire _w16277_ ;
	wire _w16276_ ;
	wire _w16275_ ;
	wire _w16274_ ;
	wire _w16273_ ;
	wire _w16272_ ;
	wire _w16271_ ;
	wire _w16270_ ;
	wire _w16269_ ;
	wire _w16268_ ;
	wire _w16267_ ;
	wire _w16266_ ;
	wire _w16265_ ;
	wire _w16264_ ;
	wire _w16263_ ;
	wire _w16262_ ;
	wire _w16261_ ;
	wire _w16260_ ;
	wire _w16259_ ;
	wire _w16258_ ;
	wire _w16257_ ;
	wire _w16256_ ;
	wire _w16255_ ;
	wire _w16254_ ;
	wire _w16253_ ;
	wire _w16252_ ;
	wire _w16251_ ;
	wire _w16250_ ;
	wire _w16249_ ;
	wire _w16248_ ;
	wire _w16247_ ;
	wire _w16246_ ;
	wire _w16245_ ;
	wire _w16244_ ;
	wire _w16243_ ;
	wire _w16242_ ;
	wire _w16241_ ;
	wire _w16240_ ;
	wire _w16239_ ;
	wire _w16238_ ;
	wire _w16237_ ;
	wire _w16236_ ;
	wire _w16235_ ;
	wire _w16234_ ;
	wire _w16233_ ;
	wire _w16232_ ;
	wire _w16231_ ;
	wire _w16230_ ;
	wire _w16229_ ;
	wire _w16228_ ;
	wire _w16227_ ;
	wire _w16226_ ;
	wire _w16225_ ;
	wire _w16224_ ;
	wire _w16223_ ;
	wire _w16222_ ;
	wire _w16221_ ;
	wire _w16220_ ;
	wire _w16219_ ;
	wire _w16218_ ;
	wire _w16217_ ;
	wire _w16216_ ;
	wire _w16215_ ;
	wire _w16214_ ;
	wire _w16213_ ;
	wire _w16212_ ;
	wire _w16211_ ;
	wire _w16210_ ;
	wire _w16209_ ;
	wire _w16208_ ;
	wire _w16207_ ;
	wire _w16206_ ;
	wire _w16205_ ;
	wire _w16204_ ;
	wire _w16203_ ;
	wire _w16202_ ;
	wire _w16201_ ;
	wire _w16200_ ;
	wire _w16199_ ;
	wire _w16198_ ;
	wire _w16197_ ;
	wire _w16196_ ;
	wire _w16195_ ;
	wire _w16194_ ;
	wire _w16193_ ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10638_ ;
	wire _w10637_ ;
	wire _w10636_ ;
	wire _w10635_ ;
	wire _w10634_ ;
	wire _w10633_ ;
	wire _w10632_ ;
	wire _w10631_ ;
	wire _w10630_ ;
	wire _w10629_ ;
	wire _w10628_ ;
	wire _w10627_ ;
	wire _w10626_ ;
	wire _w10625_ ;
	wire _w10624_ ;
	wire _w10623_ ;
	wire _w10622_ ;
	wire _w10621_ ;
	wire _w10620_ ;
	wire _w10619_ ;
	wire _w10618_ ;
	wire _w10617_ ;
	wire _w10616_ ;
	wire _w10615_ ;
	wire _w10614_ ;
	wire _w10613_ ;
	wire _w10612_ ;
	wire _w10611_ ;
	wire _w10610_ ;
	wire _w10609_ ;
	wire _w10608_ ;
	wire _w10607_ ;
	wire _w10606_ ;
	wire _w10605_ ;
	wire _w10604_ ;
	wire _w10603_ ;
	wire _w10602_ ;
	wire _w10601_ ;
	wire _w10600_ ;
	wire _w10599_ ;
	wire _w10598_ ;
	wire _w10597_ ;
	wire _w10596_ ;
	wire _w10595_ ;
	wire _w10594_ ;
	wire _w10593_ ;
	wire _w10592_ ;
	wire _w10591_ ;
	wire _w10590_ ;
	wire _w10589_ ;
	wire _w10588_ ;
	wire _w10587_ ;
	wire _w10586_ ;
	wire _w10585_ ;
	wire _w10584_ ;
	wire _w10583_ ;
	wire _w10582_ ;
	wire _w10581_ ;
	wire _w10580_ ;
	wire _w10579_ ;
	wire _w10578_ ;
	wire _w10577_ ;
	wire _w10576_ ;
	wire _w10575_ ;
	wire _w10574_ ;
	wire _w10573_ ;
	wire _w10572_ ;
	wire _w10571_ ;
	wire _w10540_ ;
	wire _w10539_ ;
	wire _w10538_ ;
	wire _w10537_ ;
	wire _w10536_ ;
	wire _w10535_ ;
	wire _w10534_ ;
	wire _w10533_ ;
	wire _w10532_ ;
	wire _w10531_ ;
	wire _w10530_ ;
	wire _w10529_ ;
	wire _w10528_ ;
	wire _w10527_ ;
	wire _w10526_ ;
	wire _w10525_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w11053_ ;
	wire _w11054_ ;
	wire _w11055_ ;
	wire _w11056_ ;
	wire _w11057_ ;
	wire _w11058_ ;
	wire _w11059_ ;
	wire _w11060_ ;
	wire _w11061_ ;
	wire _w11062_ ;
	wire _w11063_ ;
	wire _w11064_ ;
	wire _w11065_ ;
	wire _w11066_ ;
	wire _w11067_ ;
	wire _w11068_ ;
	wire _w11069_ ;
	wire _w11070_ ;
	wire _w11071_ ;
	wire _w11072_ ;
	wire _w11073_ ;
	wire _w11074_ ;
	wire _w11075_ ;
	wire _w11076_ ;
	wire _w11077_ ;
	wire _w11078_ ;
	wire _w11079_ ;
	wire _w11080_ ;
	wire _w11081_ ;
	wire _w11082_ ;
	wire _w11083_ ;
	wire _w11084_ ;
	wire _w11085_ ;
	wire _w11086_ ;
	wire _w11087_ ;
	wire _w11088_ ;
	wire _w11089_ ;
	wire _w11090_ ;
	wire _w11091_ ;
	wire _w11092_ ;
	wire _w11093_ ;
	wire _w11094_ ;
	wire _w11095_ ;
	wire _w11096_ ;
	wire _w11097_ ;
	wire _w11098_ ;
	wire _w11099_ ;
	wire _w11100_ ;
	wire _w11101_ ;
	wire _w11102_ ;
	wire _w11103_ ;
	wire _w11104_ ;
	wire _w11105_ ;
	wire _w11106_ ;
	wire _w11107_ ;
	wire _w11108_ ;
	wire _w11109_ ;
	wire _w11110_ ;
	wire _w11111_ ;
	wire _w11112_ ;
	wire _w11113_ ;
	wire _w11114_ ;
	wire _w11115_ ;
	wire _w11116_ ;
	wire _w11117_ ;
	wire _w11118_ ;
	wire _w11119_ ;
	wire _w11120_ ;
	wire _w11121_ ;
	wire _w11122_ ;
	wire _w11123_ ;
	wire _w11124_ ;
	wire _w11125_ ;
	wire _w11126_ ;
	wire _w11127_ ;
	wire _w11128_ ;
	wire _w11129_ ;
	wire _w11130_ ;
	wire _w11131_ ;
	wire _w11132_ ;
	wire _w11133_ ;
	wire _w11134_ ;
	wire _w11135_ ;
	wire _w11136_ ;
	wire _w11137_ ;
	wire _w11138_ ;
	wire _w11139_ ;
	wire _w11140_ ;
	wire _w11141_ ;
	wire _w11142_ ;
	wire _w11143_ ;
	wire _w11144_ ;
	wire _w11145_ ;
	wire _w11146_ ;
	wire _w11147_ ;
	wire _w11148_ ;
	wire _w11149_ ;
	wire _w11150_ ;
	wire _w11151_ ;
	wire _w11152_ ;
	wire _w11153_ ;
	wire _w11154_ ;
	wire _w11155_ ;
	wire _w11156_ ;
	wire _w11157_ ;
	wire _w11158_ ;
	wire _w11159_ ;
	wire _w11160_ ;
	wire _w11161_ ;
	wire _w11162_ ;
	wire _w11163_ ;
	wire _w11164_ ;
	wire _w11165_ ;
	wire _w11166_ ;
	wire _w11167_ ;
	wire _w11168_ ;
	wire _w11169_ ;
	wire _w11170_ ;
	wire _w11171_ ;
	wire _w11172_ ;
	wire _w11173_ ;
	wire _w11174_ ;
	wire _w11175_ ;
	wire _w11176_ ;
	wire _w11177_ ;
	wire _w11178_ ;
	wire _w11179_ ;
	wire _w11180_ ;
	wire _w11181_ ;
	wire _w11182_ ;
	wire _w11183_ ;
	wire _w11184_ ;
	wire _w11185_ ;
	wire _w11186_ ;
	wire _w11187_ ;
	wire _w11188_ ;
	wire _w11189_ ;
	wire _w11190_ ;
	wire _w11191_ ;
	wire _w11192_ ;
	wire _w11193_ ;
	wire _w11194_ ;
	wire _w11195_ ;
	wire _w11196_ ;
	wire _w11197_ ;
	wire _w11198_ ;
	wire _w11199_ ;
	wire _w11200_ ;
	wire _w11201_ ;
	wire _w11202_ ;
	wire _w11203_ ;
	wire _w11204_ ;
	wire _w11205_ ;
	wire _w11206_ ;
	wire _w11207_ ;
	wire _w11208_ ;
	wire _w11209_ ;
	wire _w11210_ ;
	wire _w11211_ ;
	wire _w11212_ ;
	wire _w11213_ ;
	wire _w11214_ ;
	wire _w11215_ ;
	wire _w11216_ ;
	wire _w11217_ ;
	wire _w11218_ ;
	wire _w11219_ ;
	wire _w11220_ ;
	wire _w11221_ ;
	wire _w11222_ ;
	wire _w11223_ ;
	wire _w11224_ ;
	wire _w11225_ ;
	wire _w11226_ ;
	wire _w11227_ ;
	wire _w11228_ ;
	wire _w11229_ ;
	wire _w11230_ ;
	wire _w11231_ ;
	wire _w11232_ ;
	wire _w11233_ ;
	wire _w11234_ ;
	wire _w11235_ ;
	wire _w11236_ ;
	wire _w11237_ ;
	wire _w11238_ ;
	wire _w11239_ ;
	wire _w11240_ ;
	wire _w11241_ ;
	wire _w11242_ ;
	wire _w11243_ ;
	wire _w11244_ ;
	wire _w11245_ ;
	wire _w11246_ ;
	wire _w11247_ ;
	wire _w11248_ ;
	wire _w11249_ ;
	wire _w11250_ ;
	wire _w11251_ ;
	wire _w11252_ ;
	wire _w11253_ ;
	wire _w11254_ ;
	wire _w11255_ ;
	wire _w11256_ ;
	wire _w11257_ ;
	wire _w11258_ ;
	wire _w11259_ ;
	wire _w11260_ ;
	wire _w11261_ ;
	wire _w11262_ ;
	wire _w11263_ ;
	wire _w11264_ ;
	wire _w11265_ ;
	wire _w11266_ ;
	wire _w11267_ ;
	wire _w11268_ ;
	wire _w11269_ ;
	wire _w11270_ ;
	wire _w11271_ ;
	wire _w11272_ ;
	wire _w11273_ ;
	wire _w11274_ ;
	wire _w11275_ ;
	wire _w11276_ ;
	wire _w11277_ ;
	wire _w11278_ ;
	wire _w11279_ ;
	wire _w11280_ ;
	wire _w11281_ ;
	wire _w11282_ ;
	wire _w11283_ ;
	wire _w11284_ ;
	wire _w11285_ ;
	wire _w11286_ ;
	wire _w11287_ ;
	wire _w11288_ ;
	wire _w11289_ ;
	wire _w11290_ ;
	wire _w11291_ ;
	wire _w11292_ ;
	wire _w11293_ ;
	wire _w11294_ ;
	wire _w11295_ ;
	wire _w11296_ ;
	wire _w11297_ ;
	wire _w11298_ ;
	wire _w11299_ ;
	wire _w11300_ ;
	wire _w11301_ ;
	wire _w11302_ ;
	wire _w11303_ ;
	wire _w11304_ ;
	wire _w11305_ ;
	wire _w11306_ ;
	wire _w11307_ ;
	wire _w11308_ ;
	wire _w11309_ ;
	wire _w11310_ ;
	wire _w11311_ ;
	wire _w11312_ ;
	wire _w11313_ ;
	wire _w11314_ ;
	wire _w11315_ ;
	wire _w11316_ ;
	wire _w11317_ ;
	wire _w11318_ ;
	wire _w11319_ ;
	wire _w11320_ ;
	wire _w11321_ ;
	wire _w11322_ ;
	wire _w11323_ ;
	wire _w11324_ ;
	wire _w11325_ ;
	wire _w11326_ ;
	wire _w11327_ ;
	wire _w11328_ ;
	wire _w11329_ ;
	wire _w11330_ ;
	wire _w11331_ ;
	wire _w11332_ ;
	wire _w11333_ ;
	wire _w11334_ ;
	wire _w11335_ ;
	wire _w11336_ ;
	wire _w11337_ ;
	wire _w11338_ ;
	wire _w11339_ ;
	wire _w11340_ ;
	wire _w11341_ ;
	wire _w11342_ ;
	wire _w11343_ ;
	wire _w11344_ ;
	wire _w11345_ ;
	wire _w11346_ ;
	wire _w11347_ ;
	wire _w11348_ ;
	wire _w11349_ ;
	wire _w11350_ ;
	wire _w11351_ ;
	wire _w11352_ ;
	wire _w11353_ ;
	wire _w11354_ ;
	wire _w11355_ ;
	wire _w11356_ ;
	wire _w11357_ ;
	wire _w11358_ ;
	wire _w11359_ ;
	wire _w11360_ ;
	wire _w11361_ ;
	wire _w11362_ ;
	wire _w11363_ ;
	wire _w11364_ ;
	wire _w11365_ ;
	wire _w11366_ ;
	wire _w11367_ ;
	wire _w11368_ ;
	wire _w11369_ ;
	wire _w11370_ ;
	wire _w11371_ ;
	wire _w11372_ ;
	wire _w11373_ ;
	wire _w11374_ ;
	wire _w11375_ ;
	wire _w11376_ ;
	wire _w11377_ ;
	wire _w11378_ ;
	wire _w11379_ ;
	wire _w11380_ ;
	wire _w11381_ ;
	wire _w11382_ ;
	wire _w11383_ ;
	wire _w11384_ ;
	wire _w11385_ ;
	wire _w11386_ ;
	wire _w11387_ ;
	wire _w11388_ ;
	wire _w11389_ ;
	wire _w11390_ ;
	wire _w11391_ ;
	wire _w11392_ ;
	wire _w11393_ ;
	wire _w11394_ ;
	wire _w11395_ ;
	wire _w11396_ ;
	wire _w11397_ ;
	wire _w11398_ ;
	wire _w11399_ ;
	wire _w11400_ ;
	wire _w11401_ ;
	wire _w11402_ ;
	wire _w11403_ ;
	wire _w11404_ ;
	wire _w11405_ ;
	wire _w11406_ ;
	wire _w11407_ ;
	wire _w11408_ ;
	wire _w11409_ ;
	wire _w11410_ ;
	wire _w11411_ ;
	wire _w11412_ ;
	wire _w11413_ ;
	wire _w11414_ ;
	wire _w11415_ ;
	wire _w11416_ ;
	wire _w11417_ ;
	wire _w11418_ ;
	wire _w11419_ ;
	wire _w11420_ ;
	wire _w11421_ ;
	wire _w11422_ ;
	wire _w11423_ ;
	wire _w11424_ ;
	wire _w11425_ ;
	wire _w11426_ ;
	wire _w11427_ ;
	wire _w11428_ ;
	wire _w11429_ ;
	wire _w11430_ ;
	wire _w11431_ ;
	wire _w11432_ ;
	wire _w11433_ ;
	wire _w11434_ ;
	wire _w11435_ ;
	wire _w11436_ ;
	wire _w11437_ ;
	wire _w11438_ ;
	wire _w11439_ ;
	wire _w11440_ ;
	wire _w11441_ ;
	wire _w11442_ ;
	wire _w11443_ ;
	wire _w11444_ ;
	wire _w11445_ ;
	wire _w11446_ ;
	wire _w11447_ ;
	wire _w11448_ ;
	wire _w11449_ ;
	wire _w11450_ ;
	wire _w11451_ ;
	wire _w11452_ ;
	wire _w11453_ ;
	wire _w11454_ ;
	wire _w11455_ ;
	wire _w11456_ ;
	wire _w11457_ ;
	wire _w11458_ ;
	wire _w11459_ ;
	wire _w11460_ ;
	wire _w11461_ ;
	wire _w11462_ ;
	wire _w11463_ ;
	wire _w11464_ ;
	wire _w11465_ ;
	wire _w11466_ ;
	wire _w11467_ ;
	wire _w11468_ ;
	wire _w11469_ ;
	wire _w11470_ ;
	wire _w11471_ ;
	wire _w11472_ ;
	wire _w11473_ ;
	wire _w11474_ ;
	wire _w11475_ ;
	wire _w11476_ ;
	wire _w11477_ ;
	wire _w11478_ ;
	wire _w11479_ ;
	wire _w11480_ ;
	wire _w11481_ ;
	wire _w11482_ ;
	wire _w11483_ ;
	wire _w11484_ ;
	wire _w11485_ ;
	wire _w11486_ ;
	wire _w11487_ ;
	wire _w11488_ ;
	wire _w11489_ ;
	wire _w11490_ ;
	wire _w11491_ ;
	wire _w11492_ ;
	wire _w11493_ ;
	wire _w11494_ ;
	wire _w11495_ ;
	wire _w11496_ ;
	wire _w11497_ ;
	wire _w11498_ ;
	wire _w11499_ ;
	wire _w11500_ ;
	wire _w11501_ ;
	wire _w11502_ ;
	wire _w11503_ ;
	wire _w11504_ ;
	wire _w11505_ ;
	wire _w11506_ ;
	wire _w11507_ ;
	wire _w11508_ ;
	wire _w11509_ ;
	wire _w11510_ ;
	wire _w11511_ ;
	wire _w11512_ ;
	wire _w11513_ ;
	wire _w11514_ ;
	wire _w11515_ ;
	wire _w11516_ ;
	wire _w11517_ ;
	wire _w11518_ ;
	wire _w11519_ ;
	wire _w11520_ ;
	wire _w11521_ ;
	wire _w11522_ ;
	wire _w11523_ ;
	wire _w11524_ ;
	wire _w11525_ ;
	wire _w11526_ ;
	wire _w11527_ ;
	wire _w11528_ ;
	wire _w11529_ ;
	wire _w11530_ ;
	wire _w11531_ ;
	wire _w11532_ ;
	wire _w11533_ ;
	wire _w11534_ ;
	wire _w11535_ ;
	wire _w11536_ ;
	wire _w11537_ ;
	wire _w11538_ ;
	wire _w11539_ ;
	wire _w11540_ ;
	wire _w11541_ ;
	wire _w11542_ ;
	wire _w11543_ ;
	wire _w11544_ ;
	wire _w11545_ ;
	wire _w11546_ ;
	wire _w11547_ ;
	wire _w11548_ ;
	wire _w11549_ ;
	wire _w11550_ ;
	wire _w11551_ ;
	wire _w11552_ ;
	wire _w11553_ ;
	wire _w11554_ ;
	wire _w11555_ ;
	wire _w11556_ ;
	wire _w11557_ ;
	wire _w11558_ ;
	wire _w11559_ ;
	wire _w11560_ ;
	wire _w11561_ ;
	wire _w11562_ ;
	wire _w11563_ ;
	wire _w11564_ ;
	wire _w11565_ ;
	wire _w11566_ ;
	wire _w11567_ ;
	wire _w11568_ ;
	wire _w11569_ ;
	wire _w11570_ ;
	wire _w11571_ ;
	wire _w11572_ ;
	wire _w11573_ ;
	wire _w11574_ ;
	wire _w11575_ ;
	wire _w11576_ ;
	wire _w11577_ ;
	wire _w11578_ ;
	wire _w11579_ ;
	wire _w11580_ ;
	wire _w11581_ ;
	wire _w11582_ ;
	wire _w11583_ ;
	wire _w11584_ ;
	wire _w11585_ ;
	wire _w11586_ ;
	wire _w11587_ ;
	wire _w11588_ ;
	wire _w11589_ ;
	wire _w11590_ ;
	wire _w11591_ ;
	wire _w11592_ ;
	wire _w11593_ ;
	wire _w11594_ ;
	wire _w11595_ ;
	wire _w11596_ ;
	wire _w11597_ ;
	wire _w11598_ ;
	wire _w11599_ ;
	wire _w11600_ ;
	wire _w11601_ ;
	wire _w11602_ ;
	wire _w11603_ ;
	wire _w11604_ ;
	wire _w11605_ ;
	wire _w11606_ ;
	wire _w11607_ ;
	wire _w11608_ ;
	wire _w11609_ ;
	wire _w11610_ ;
	wire _w11611_ ;
	wire _w11612_ ;
	wire _w11613_ ;
	wire _w11614_ ;
	wire _w11615_ ;
	wire _w11616_ ;
	wire _w11617_ ;
	wire _w11618_ ;
	wire _w11619_ ;
	wire _w11620_ ;
	wire _w12869_ ;
	wire _w12870_ ;
	wire _w12871_ ;
	wire _w12872_ ;
	wire _w12873_ ;
	wire _w12874_ ;
	wire _w12875_ ;
	wire _w12876_ ;
	wire _w12877_ ;
	wire _w12878_ ;
	wire _w12879_ ;
	wire _w12880_ ;
	wire _w12881_ ;
	wire _w12882_ ;
	wire _w12883_ ;
	wire _w12884_ ;
	wire _w12885_ ;
	wire _w12886_ ;
	wire _w12887_ ;
	wire _w12888_ ;
	wire _w12889_ ;
	wire _w12890_ ;
	wire _w12891_ ;
	wire _w12892_ ;
	wire _w12893_ ;
	wire _w12894_ ;
	wire _w12895_ ;
	wire _w12896_ ;
	wire _w12897_ ;
	wire _w12898_ ;
	wire _w12899_ ;
	wire _w12900_ ;
	wire _w12901_ ;
	wire _w12902_ ;
	wire _w12903_ ;
	wire _w12904_ ;
	wire _w12905_ ;
	wire _w12906_ ;
	wire _w12907_ ;
	wire _w12908_ ;
	wire _w12909_ ;
	wire _w12910_ ;
	wire _w12911_ ;
	wire _w12912_ ;
	wire _w12913_ ;
	wire _w12914_ ;
	wire _w12915_ ;
	wire _w12916_ ;
	wire _w12917_ ;
	wire _w12918_ ;
	wire _w12919_ ;
	wire _w12920_ ;
	wire _w12921_ ;
	wire _w12922_ ;
	wire _w12923_ ;
	wire _w12924_ ;
	wire _w12925_ ;
	wire _w12926_ ;
	wire _w12927_ ;
	wire _w12928_ ;
	wire _w12929_ ;
	wire _w12930_ ;
	wire _w12931_ ;
	wire _w12932_ ;
	wire _w12933_ ;
	wire _w12934_ ;
	wire _w12935_ ;
	wire _w12936_ ;
	wire _w12937_ ;
	wire _w12938_ ;
	wire _w12939_ ;
	wire _w12940_ ;
	wire _w12941_ ;
	wire _w12942_ ;
	wire _w12943_ ;
	wire _w12944_ ;
	wire _w12945_ ;
	wire _w12946_ ;
	wire _w12947_ ;
	wire _w12948_ ;
	wire _w12949_ ;
	wire _w12950_ ;
	wire _w12951_ ;
	wire _w12952_ ;
	wire _w12953_ ;
	wire _w12954_ ;
	wire _w12955_ ;
	wire _w12956_ ;
	wire _w12957_ ;
	wire _w12958_ ;
	wire _w12959_ ;
	wire _w12960_ ;
	wire _w12961_ ;
	wire _w12962_ ;
	wire _w12963_ ;
	wire _w12964_ ;
	wire _w12965_ ;
	wire _w12966_ ;
	wire _w12967_ ;
	wire _w12968_ ;
	wire _w12969_ ;
	wire _w12970_ ;
	wire _w12971_ ;
	wire _w12972_ ;
	wire _w12973_ ;
	wire _w12974_ ;
	wire _w12975_ ;
	wire _w12976_ ;
	wire _w12977_ ;
	wire _w12978_ ;
	wire _w12979_ ;
	wire _w12980_ ;
	wire _w12981_ ;
	wire _w12982_ ;
	wire _w12983_ ;
	wire _w12984_ ;
	wire _w12985_ ;
	wire _w12986_ ;
	wire _w12987_ ;
	wire _w12988_ ;
	wire _w12989_ ;
	wire _w12990_ ;
	wire _w12991_ ;
	wire _w12992_ ;
	wire _w12993_ ;
	wire _w12994_ ;
	wire _w12995_ ;
	wire _w12996_ ;
	wire _w12997_ ;
	wire _w12998_ ;
	wire _w12999_ ;
	wire _w13000_ ;
	wire _w13001_ ;
	wire _w13002_ ;
	wire _w13003_ ;
	wire _w13004_ ;
	wire _w13005_ ;
	wire _w13006_ ;
	wire _w13007_ ;
	wire _w13008_ ;
	wire _w13009_ ;
	wire _w13010_ ;
	wire _w13011_ ;
	wire _w13012_ ;
	wire _w13013_ ;
	wire _w13014_ ;
	wire _w13015_ ;
	wire _w13016_ ;
	wire _w13017_ ;
	wire _w13018_ ;
	wire _w13019_ ;
	wire _w13020_ ;
	wire _w13021_ ;
	wire _w13022_ ;
	wire _w13023_ ;
	wire _w13024_ ;
	wire _w13025_ ;
	wire _w13026_ ;
	wire _w13027_ ;
	wire _w13028_ ;
	wire _w13029_ ;
	wire _w13030_ ;
	wire _w13031_ ;
	wire _w13032_ ;
	wire _w13033_ ;
	wire _w13034_ ;
	wire _w13035_ ;
	wire _w13036_ ;
	wire _w13037_ ;
	wire _w13038_ ;
	wire _w13039_ ;
	wire _w13040_ ;
	wire _w13041_ ;
	wire _w13042_ ;
	wire _w13043_ ;
	wire _w13044_ ;
	wire _w13045_ ;
	wire _w13046_ ;
	wire _w13047_ ;
	wire _w13048_ ;
	wire _w13049_ ;
	wire _w13050_ ;
	wire _w13051_ ;
	wire _w13052_ ;
	wire _w13053_ ;
	wire _w13054_ ;
	wire _w13055_ ;
	wire _w13056_ ;
	wire _w13057_ ;
	wire _w13058_ ;
	wire _w13059_ ;
	wire _w13060_ ;
	wire _w13061_ ;
	wire _w13062_ ;
	wire _w13063_ ;
	wire _w13064_ ;
	wire _w13065_ ;
	wire _w13066_ ;
	wire _w13067_ ;
	wire _w13068_ ;
	wire _w13069_ ;
	wire _w13070_ ;
	wire _w13071_ ;
	wire _w13072_ ;
	wire _w13073_ ;
	wire _w13074_ ;
	wire _w13075_ ;
	wire _w13076_ ;
	wire _w13077_ ;
	wire _w13078_ ;
	wire _w13079_ ;
	wire _w13080_ ;
	wire _w13081_ ;
	wire _w13082_ ;
	wire _w13083_ ;
	wire _w13084_ ;
	wire _w13085_ ;
	wire _w13086_ ;
	wire _w13087_ ;
	wire _w13088_ ;
	wire _w13089_ ;
	wire _w13090_ ;
	wire _w13091_ ;
	wire _w13092_ ;
	wire _w13093_ ;
	wire _w13094_ ;
	wire _w13095_ ;
	wire _w13096_ ;
	wire _w13097_ ;
	wire _w13098_ ;
	wire _w13099_ ;
	wire _w13100_ ;
	wire _w13101_ ;
	wire _w13102_ ;
	wire _w13103_ ;
	wire _w13104_ ;
	wire _w13105_ ;
	wire _w13106_ ;
	wire _w13107_ ;
	wire _w13108_ ;
	wire _w13109_ ;
	wire _w13110_ ;
	wire _w13111_ ;
	wire _w13112_ ;
	wire _w13113_ ;
	wire _w13114_ ;
	wire _w13115_ ;
	wire _w13116_ ;
	wire _w13117_ ;
	wire _w13118_ ;
	wire _w13119_ ;
	wire _w13120_ ;
	wire _w13121_ ;
	wire _w13122_ ;
	wire _w13123_ ;
	wire _w13124_ ;
	wire _w13125_ ;
	wire _w13126_ ;
	wire _w13127_ ;
	wire _w13128_ ;
	wire _w13129_ ;
	wire _w13130_ ;
	wire _w13131_ ;
	wire _w13132_ ;
	wire _w13133_ ;
	wire _w13134_ ;
	wire _w13135_ ;
	wire _w13136_ ;
	wire _w13137_ ;
	wire _w13138_ ;
	wire _w13139_ ;
	wire _w13140_ ;
	wire _w13141_ ;
	wire _w13142_ ;
	wire _w13143_ ;
	wire _w13144_ ;
	wire _w13145_ ;
	wire _w13146_ ;
	wire _w13147_ ;
	wire _w13148_ ;
	wire _w13149_ ;
	wire _w13150_ ;
	wire _w13151_ ;
	wire _w13152_ ;
	wire _w13153_ ;
	wire _w13154_ ;
	wire _w13155_ ;
	wire _w13156_ ;
	wire _w13157_ ;
	wire _w13158_ ;
	wire _w13159_ ;
	wire _w13160_ ;
	wire _w13161_ ;
	wire _w13162_ ;
	wire _w13163_ ;
	wire _w13164_ ;
	wire _w13165_ ;
	wire _w13166_ ;
	wire _w13167_ ;
	wire _w13168_ ;
	wire _w13169_ ;
	wire _w13170_ ;
	wire _w13171_ ;
	wire _w13172_ ;
	wire _w13173_ ;
	wire _w13174_ ;
	wire _w13175_ ;
	wire _w13176_ ;
	wire _w13177_ ;
	wire _w13178_ ;
	wire _w13179_ ;
	wire _w13180_ ;
	wire _w13181_ ;
	wire _w13182_ ;
	wire _w13183_ ;
	wire _w13184_ ;
	wire _w13185_ ;
	wire _w13186_ ;
	wire _w13187_ ;
	wire _w13188_ ;
	wire _w13189_ ;
	wire _w13190_ ;
	wire _w13191_ ;
	wire _w13192_ ;
	wire _w13193_ ;
	wire _w13194_ ;
	wire _w13195_ ;
	wire _w13196_ ;
	wire _w13197_ ;
	wire _w13198_ ;
	wire _w13199_ ;
	wire _w13200_ ;
	wire _w13201_ ;
	wire _w13202_ ;
	wire _w13203_ ;
	wire _w13204_ ;
	wire _w13205_ ;
	wire _w13206_ ;
	wire _w13207_ ;
	wire _w13208_ ;
	wire _w13209_ ;
	wire _w13210_ ;
	wire _w13211_ ;
	wire _w13212_ ;
	wire _w13213_ ;
	wire _w13214_ ;
	wire _w13215_ ;
	wire _w13216_ ;
	wire _w13217_ ;
	wire _w13218_ ;
	wire _w13219_ ;
	wire _w13220_ ;
	wire _w13221_ ;
	wire _w13222_ ;
	wire _w13223_ ;
	wire _w13224_ ;
	wire _w13225_ ;
	wire _w13226_ ;
	wire _w13227_ ;
	wire _w13228_ ;
	wire _w13229_ ;
	wire _w13230_ ;
	wire _w13231_ ;
	wire _w13232_ ;
	wire _w13233_ ;
	wire _w13234_ ;
	wire _w13235_ ;
	wire _w13236_ ;
	wire _w13237_ ;
	wire _w13238_ ;
	wire _w13239_ ;
	wire _w13240_ ;
	wire _w13241_ ;
	wire _w13242_ ;
	wire _w13243_ ;
	wire _w13244_ ;
	wire _w13245_ ;
	wire _w13246_ ;
	wire _w13247_ ;
	wire _w13248_ ;
	wire _w13249_ ;
	wire _w13250_ ;
	wire _w13251_ ;
	wire _w13252_ ;
	wire _w13253_ ;
	wire _w13254_ ;
	wire _w13255_ ;
	wire _w13256_ ;
	wire _w13257_ ;
	wire _w13258_ ;
	wire _w13259_ ;
	wire _w13260_ ;
	wire _w13261_ ;
	wire _w13262_ ;
	wire _w13263_ ;
	wire _w13264_ ;
	wire _w13265_ ;
	wire _w13266_ ;
	wire _w13267_ ;
	wire _w13268_ ;
	wire _w13269_ ;
	wire _w13270_ ;
	wire _w13271_ ;
	wire _w13272_ ;
	wire _w13273_ ;
	wire _w13274_ ;
	wire _w13275_ ;
	wire _w13276_ ;
	wire _w13277_ ;
	wire _w13278_ ;
	wire _w13279_ ;
	wire _w13280_ ;
	wire _w13281_ ;
	wire _w13282_ ;
	wire _w13283_ ;
	wire _w13284_ ;
	wire _w13285_ ;
	wire _w13286_ ;
	wire _w13287_ ;
	wire _w13288_ ;
	wire _w13289_ ;
	wire _w13290_ ;
	wire _w13291_ ;
	wire _w13292_ ;
	wire _w13293_ ;
	wire _w13294_ ;
	wire _w13295_ ;
	wire _w13296_ ;
	wire _w13297_ ;
	wire _w13298_ ;
	wire _w13299_ ;
	wire _w13300_ ;
	wire _w13301_ ;
	wire _w13302_ ;
	wire _w13303_ ;
	wire _w13304_ ;
	wire _w13305_ ;
	wire _w13306_ ;
	wire _w13307_ ;
	wire _w13308_ ;
	wire _w13309_ ;
	wire _w13310_ ;
	wire _w13311_ ;
	wire _w13312_ ;
	wire _w13313_ ;
	wire _w13314_ ;
	wire _w13315_ ;
	wire _w13316_ ;
	wire _w13317_ ;
	wire _w13318_ ;
	wire _w13319_ ;
	wire _w13320_ ;
	wire _w13321_ ;
	wire _w13322_ ;
	wire _w13323_ ;
	wire _w13324_ ;
	wire _w13325_ ;
	wire _w13326_ ;
	wire _w13327_ ;
	wire _w13328_ ;
	wire _w13329_ ;
	wire _w13330_ ;
	wire _w13331_ ;
	wire _w13332_ ;
	wire _w13333_ ;
	wire _w13334_ ;
	wire _w13335_ ;
	wire _w13336_ ;
	wire _w13337_ ;
	wire _w13338_ ;
	wire _w13339_ ;
	wire _w13340_ ;
	wire _w13341_ ;
	wire _w13342_ ;
	wire _w13343_ ;
	wire _w13344_ ;
	wire _w13345_ ;
	wire _w13346_ ;
	wire _w13347_ ;
	wire _w13348_ ;
	wire _w13349_ ;
	wire _w13350_ ;
	wire _w13351_ ;
	wire _w13352_ ;
	wire _w13353_ ;
	wire _w13354_ ;
	wire _w13355_ ;
	wire _w13356_ ;
	wire _w13357_ ;
	wire _w13358_ ;
	wire _w13359_ ;
	wire _w13360_ ;
	wire _w13361_ ;
	wire _w13362_ ;
	wire _w13363_ ;
	wire _w13364_ ;
	wire _w13365_ ;
	wire _w13366_ ;
	wire _w13367_ ;
	wire _w13368_ ;
	wire _w13369_ ;
	wire _w13370_ ;
	wire _w13371_ ;
	wire _w13372_ ;
	wire _w13373_ ;
	wire _w13374_ ;
	wire _w13375_ ;
	wire _w13376_ ;
	wire _w13377_ ;
	wire _w13378_ ;
	wire _w13379_ ;
	wire _w13380_ ;
	wire _w13381_ ;
	wire _w13382_ ;
	wire _w13383_ ;
	wire _w13384_ ;
	wire _w13385_ ;
	wire _w13386_ ;
	wire _w13387_ ;
	wire _w13388_ ;
	wire _w13389_ ;
	wire _w13390_ ;
	wire _w13391_ ;
	wire _w13392_ ;
	wire _w13393_ ;
	wire _w13394_ ;
	wire _w13395_ ;
	wire _w13396_ ;
	wire _w13397_ ;
	wire _w13398_ ;
	wire _w13399_ ;
	wire _w13400_ ;
	wire _w13401_ ;
	wire _w13402_ ;
	wire _w13403_ ;
	wire _w13404_ ;
	wire _w13405_ ;
	wire _w13406_ ;
	wire _w13407_ ;
	wire _w13408_ ;
	wire _w13409_ ;
	wire _w13410_ ;
	wire _w13411_ ;
	wire _w13412_ ;
	wire _w13413_ ;
	wire _w13414_ ;
	wire _w13415_ ;
	wire _w13416_ ;
	wire _w13417_ ;
	wire _w13418_ ;
	wire _w13419_ ;
	wire _w13420_ ;
	wire _w13421_ ;
	wire _w13422_ ;
	wire _w13423_ ;
	wire _w13424_ ;
	wire _w13425_ ;
	wire _w13426_ ;
	wire _w13427_ ;
	wire _w13428_ ;
	wire _w13429_ ;
	wire _w13430_ ;
	wire _w13431_ ;
	wire _w13432_ ;
	wire _w13433_ ;
	wire _w13434_ ;
	wire _w13435_ ;
	wire _w13436_ ;
	wire _w13437_ ;
	wire _w13438_ ;
	wire _w13439_ ;
	wire _w13440_ ;
	wire _w13441_ ;
	wire _w13442_ ;
	wire _w13443_ ;
	wire _w13444_ ;
	wire _w13445_ ;
	wire _w13446_ ;
	wire _w13447_ ;
	wire _w13448_ ;
	wire _w13449_ ;
	wire _w13450_ ;
	wire _w13451_ ;
	wire _w13452_ ;
	wire _w13453_ ;
	wire _w13454_ ;
	wire _w13455_ ;
	wire _w13456_ ;
	wire _w13457_ ;
	wire _w13458_ ;
	wire _w13459_ ;
	wire _w13460_ ;
	wire _w13461_ ;
	wire _w13462_ ;
	wire _w13463_ ;
	wire _w13464_ ;
	wire _w13465_ ;
	wire _w13466_ ;
	wire _w13467_ ;
	wire _w13468_ ;
	wire _w13469_ ;
	wire _w13470_ ;
	wire _w13471_ ;
	wire _w13472_ ;
	wire _w13473_ ;
	wire _w13474_ ;
	wire _w13475_ ;
	wire _w13476_ ;
	wire _w13477_ ;
	wire _w13478_ ;
	wire _w13479_ ;
	wire _w13480_ ;
	wire _w13481_ ;
	wire _w13482_ ;
	wire _w13483_ ;
	wire _w13484_ ;
	wire _w13485_ ;
	wire _w13486_ ;
	wire _w13487_ ;
	wire _w13488_ ;
	wire _w13489_ ;
	wire _w13490_ ;
	wire _w13491_ ;
	wire _w13492_ ;
	wire _w13493_ ;
	wire _w13494_ ;
	wire _w13495_ ;
	wire _w13496_ ;
	wire _w13497_ ;
	wire _w13498_ ;
	wire _w13499_ ;
	wire _w13500_ ;
	wire _w13501_ ;
	wire _w13502_ ;
	wire _w13503_ ;
	wire _w13504_ ;
	wire _w13505_ ;
	wire _w13506_ ;
	wire _w13507_ ;
	wire _w13508_ ;
	wire _w13509_ ;
	wire _w13510_ ;
	wire _w13511_ ;
	wire _w13512_ ;
	wire _w13513_ ;
	wire _w13514_ ;
	wire _w13515_ ;
	wire _w13516_ ;
	wire _w13517_ ;
	wire _w13518_ ;
	wire _w13519_ ;
	wire _w13520_ ;
	wire _w13521_ ;
	wire _w13522_ ;
	wire _w13523_ ;
	wire _w13524_ ;
	wire _w13525_ ;
	wire _w13526_ ;
	wire _w13527_ ;
	wire _w13528_ ;
	wire _w13529_ ;
	wire _w13530_ ;
	wire _w13531_ ;
	wire _w13532_ ;
	wire _w13533_ ;
	wire _w13534_ ;
	wire _w13535_ ;
	wire _w13536_ ;
	wire _w13537_ ;
	wire _w13538_ ;
	wire _w13539_ ;
	wire _w13540_ ;
	wire _w13541_ ;
	wire _w13542_ ;
	wire _w13543_ ;
	wire _w13544_ ;
	wire _w13545_ ;
	wire _w13546_ ;
	wire _w13547_ ;
	wire _w13548_ ;
	wire _w13549_ ;
	wire _w13550_ ;
	wire _w13551_ ;
	wire _w13552_ ;
	wire _w13553_ ;
	wire _w13554_ ;
	wire _w13555_ ;
	wire _w13556_ ;
	wire _w13557_ ;
	wire _w13558_ ;
	wire _w13559_ ;
	wire _w13560_ ;
	wire _w13561_ ;
	wire _w13562_ ;
	wire _w13563_ ;
	wire _w13564_ ;
	wire _w13565_ ;
	wire _w13566_ ;
	wire _w13567_ ;
	wire _w13568_ ;
	wire _w13569_ ;
	wire _w13570_ ;
	wire _w13571_ ;
	wire _w13572_ ;
	wire _w13573_ ;
	wire _w13574_ ;
	wire _w13575_ ;
	wire _w13576_ ;
	wire _w13577_ ;
	wire _w13578_ ;
	wire _w13579_ ;
	wire _w13580_ ;
	wire _w13581_ ;
	wire _w13582_ ;
	wire _w13583_ ;
	wire _w13584_ ;
	wire _w13585_ ;
	wire _w13586_ ;
	wire _w13587_ ;
	wire _w13588_ ;
	wire _w13589_ ;
	wire _w13590_ ;
	wire _w13591_ ;
	wire _w13592_ ;
	wire _w13593_ ;
	wire _w13594_ ;
	wire _w13595_ ;
	wire _w13596_ ;
	wire _w13597_ ;
	wire _w13598_ ;
	wire _w13599_ ;
	wire _w13600_ ;
	wire _w13601_ ;
	wire _w13602_ ;
	wire _w13603_ ;
	wire _w13604_ ;
	wire _w13605_ ;
	wire _w13606_ ;
	wire _w13607_ ;
	wire _w13608_ ;
	wire _w13609_ ;
	wire _w13610_ ;
	wire _w13611_ ;
	wire _w13612_ ;
	wire _w13613_ ;
	wire _w13614_ ;
	wire _w13615_ ;
	wire _w13616_ ;
	wire _w13617_ ;
	wire _w13618_ ;
	wire _w13619_ ;
	wire _w13620_ ;
	wire _w13621_ ;
	wire _w13622_ ;
	wire _w13623_ ;
	wire _w13624_ ;
	wire _w13625_ ;
	wire _w13626_ ;
	wire _w13627_ ;
	wire _w13628_ ;
	wire _w13629_ ;
	wire _w13630_ ;
	wire _w13631_ ;
	wire _w13632_ ;
	wire _w13633_ ;
	wire _w13634_ ;
	wire _w13635_ ;
	wire _w13636_ ;
	wire _w13637_ ;
	wire _w13638_ ;
	wire _w13639_ ;
	wire _w13640_ ;
	wire _w13641_ ;
	wire _w13642_ ;
	wire _w13643_ ;
	wire _w13644_ ;
	wire _w13645_ ;
	wire _w13646_ ;
	wire _w13647_ ;
	wire _w13648_ ;
	wire _w13649_ ;
	wire _w13650_ ;
	wire _w13651_ ;
	wire _w13652_ ;
	wire _w13653_ ;
	wire _w13654_ ;
	wire _w13655_ ;
	wire _w13656_ ;
	wire _w13657_ ;
	wire _w13658_ ;
	wire _w13659_ ;
	wire _w13660_ ;
	wire _w13661_ ;
	wire _w13662_ ;
	wire _w13663_ ;
	wire _w13664_ ;
	wire _w13665_ ;
	wire _w13666_ ;
	wire _w13667_ ;
	wire _w13668_ ;
	wire _w13669_ ;
	wire _w13670_ ;
	wire _w13671_ ;
	wire _w13672_ ;
	wire _w13673_ ;
	wire _w13674_ ;
	wire _w13675_ ;
	wire _w13676_ ;
	wire _w13677_ ;
	wire _w13678_ ;
	wire _w13679_ ;
	wire _w13680_ ;
	wire _w13681_ ;
	wire _w13682_ ;
	wire _w13683_ ;
	wire _w13684_ ;
	wire _w13685_ ;
	wire _w13686_ ;
	wire _w13687_ ;
	wire _w13688_ ;
	wire _w13689_ ;
	wire _w13690_ ;
	wire _w13691_ ;
	wire _w13692_ ;
	wire _w13693_ ;
	wire _w13694_ ;
	wire _w13695_ ;
	wire _w13696_ ;
	wire _w13697_ ;
	wire _w13698_ ;
	wire _w13699_ ;
	wire _w13700_ ;
	wire _w13701_ ;
	wire _w13702_ ;
	wire _w13703_ ;
	wire _w13704_ ;
	wire _w13705_ ;
	wire _w13706_ ;
	wire _w13707_ ;
	wire _w13708_ ;
	wire _w13709_ ;
	wire _w13710_ ;
	wire _w13711_ ;
	wire _w13712_ ;
	wire _w13713_ ;
	wire _w13714_ ;
	wire _w13715_ ;
	wire _w13716_ ;
	wire _w13717_ ;
	wire _w13718_ ;
	wire _w13719_ ;
	wire _w13720_ ;
	wire _w13721_ ;
	wire _w13722_ ;
	wire _w13723_ ;
	wire _w13724_ ;
	wire _w13725_ ;
	wire _w13726_ ;
	wire _w13727_ ;
	wire _w13728_ ;
	wire _w13729_ ;
	wire _w13730_ ;
	wire _w13731_ ;
	wire _w13732_ ;
	wire _w13733_ ;
	wire _w13734_ ;
	wire _w13735_ ;
	wire _w13736_ ;
	wire _w13737_ ;
	wire _w13738_ ;
	wire _w13739_ ;
	wire _w13740_ ;
	wire _w13741_ ;
	wire _w13742_ ;
	wire _w13743_ ;
	wire _w13744_ ;
	wire _w13745_ ;
	wire _w13746_ ;
	wire _w13747_ ;
	wire _w13748_ ;
	wire _w13749_ ;
	wire _w13750_ ;
	wire _w13751_ ;
	wire _w13752_ ;
	wire _w13753_ ;
	wire _w13754_ ;
	wire _w13755_ ;
	wire _w13756_ ;
	wire _w13757_ ;
	wire _w13758_ ;
	wire _w13759_ ;
	wire _w13760_ ;
	wire _w13761_ ;
	wire _w13762_ ;
	wire _w13763_ ;
	wire _w13764_ ;
	wire _w13765_ ;
	wire _w13766_ ;
	wire _w13767_ ;
	wire _w13768_ ;
	wire _w13769_ ;
	wire _w13770_ ;
	wire _w13771_ ;
	wire _w13772_ ;
	wire _w13773_ ;
	wire _w13774_ ;
	wire _w13775_ ;
	wire _w13776_ ;
	wire _w13777_ ;
	wire _w13778_ ;
	wire _w13779_ ;
	wire _w13780_ ;
	wire _w13781_ ;
	wire _w13782_ ;
	wire _w13783_ ;
	wire _w13784_ ;
	wire _w13785_ ;
	wire _w13786_ ;
	wire _w13787_ ;
	wire _w13788_ ;
	wire _w13789_ ;
	wire _w13790_ ;
	wire _w13791_ ;
	wire _w13792_ ;
	wire _w13793_ ;
	wire _w13794_ ;
	wire _w13795_ ;
	wire _w13796_ ;
	wire _w13797_ ;
	wire _w13798_ ;
	wire _w13799_ ;
	wire _w13800_ ;
	wire _w13801_ ;
	wire _w13802_ ;
	wire _w13803_ ;
	wire _w13804_ ;
	wire _w13805_ ;
	wire _w13806_ ;
	wire _w13807_ ;
	wire _w13808_ ;
	wire _w13809_ ;
	wire _w13810_ ;
	wire _w13811_ ;
	wire _w13812_ ;
	wire _w13813_ ;
	wire _w13814_ ;
	wire _w13815_ ;
	wire _w13816_ ;
	wire _w13817_ ;
	wire _w13818_ ;
	wire _w13819_ ;
	wire _w13820_ ;
	wire _w13821_ ;
	wire _w13822_ ;
	wire _w13823_ ;
	wire _w13824_ ;
	wire _w13825_ ;
	wire _w13826_ ;
	wire _w13827_ ;
	wire _w13828_ ;
	wire _w13829_ ;
	wire _w13830_ ;
	wire _w13831_ ;
	wire _w13832_ ;
	wire _w13833_ ;
	wire _w13834_ ;
	wire _w13835_ ;
	wire _w13836_ ;
	wire _w13837_ ;
	wire _w13838_ ;
	wire _w13839_ ;
	wire _w13840_ ;
	wire _w13841_ ;
	wire _w13842_ ;
	wire _w13843_ ;
	wire _w13844_ ;
	wire _w13845_ ;
	wire _w13846_ ;
	wire _w13847_ ;
	wire _w13848_ ;
	wire _w13849_ ;
	wire _w13850_ ;
	wire _w13851_ ;
	wire _w13852_ ;
	wire _w13853_ ;
	wire _w13854_ ;
	wire _w13855_ ;
	wire _w13856_ ;
	wire _w13857_ ;
	wire _w13858_ ;
	wire _w13859_ ;
	wire _w13860_ ;
	wire _w13861_ ;
	wire _w13862_ ;
	wire _w13863_ ;
	wire _w13864_ ;
	wire _w13865_ ;
	wire _w13866_ ;
	wire _w13867_ ;
	wire _w13868_ ;
	wire _w13869_ ;
	wire _w13870_ ;
	wire _w13871_ ;
	wire _w13872_ ;
	wire _w13873_ ;
	wire _w13874_ ;
	wire _w13875_ ;
	wire _w13876_ ;
	wire _w13877_ ;
	wire _w13878_ ;
	wire _w13879_ ;
	wire _w13880_ ;
	wire _w13881_ ;
	wire _w13882_ ;
	wire _w13883_ ;
	wire _w13884_ ;
	wire _w13885_ ;
	wire _w13886_ ;
	wire _w13887_ ;
	wire _w13888_ ;
	wire _w13889_ ;
	wire _w13890_ ;
	wire _w13891_ ;
	wire _w13892_ ;
	wire _w13893_ ;
	wire _w13894_ ;
	wire _w13895_ ;
	wire _w13896_ ;
	wire _w13897_ ;
	wire _w13898_ ;
	wire _w13899_ ;
	wire _w13900_ ;
	wire _w13901_ ;
	wire _w13902_ ;
	wire _w13903_ ;
	wire _w13904_ ;
	wire _w13905_ ;
	wire _w13906_ ;
	wire _w13907_ ;
	wire _w13908_ ;
	wire _w13909_ ;
	wire _w13910_ ;
	wire _w13911_ ;
	wire _w13912_ ;
	wire _w13913_ ;
	wire _w13914_ ;
	wire _w13915_ ;
	wire _w13916_ ;
	wire _w13917_ ;
	wire _w13918_ ;
	wire _w13919_ ;
	wire _w13920_ ;
	wire _w13921_ ;
	wire _w13922_ ;
	wire _w13923_ ;
	wire _w13924_ ;
	wire _w13925_ ;
	wire _w13926_ ;
	wire _w13927_ ;
	wire _w13928_ ;
	wire _w13929_ ;
	wire _w13930_ ;
	wire _w13931_ ;
	wire _w13932_ ;
	wire _w13933_ ;
	wire _w13934_ ;
	wire _w13935_ ;
	wire _w13936_ ;
	wire _w13937_ ;
	wire _w13938_ ;
	wire _w13939_ ;
	wire _w13940_ ;
	wire _w13941_ ;
	wire _w13942_ ;
	wire _w13943_ ;
	wire _w13944_ ;
	wire _w13945_ ;
	wire _w13946_ ;
	wire _w13947_ ;
	wire _w13948_ ;
	wire _w13949_ ;
	wire _w13950_ ;
	wire _w13951_ ;
	wire _w13952_ ;
	wire _w13953_ ;
	wire _w13954_ ;
	wire _w13955_ ;
	wire _w13956_ ;
	wire _w13957_ ;
	wire _w13958_ ;
	wire _w13959_ ;
	wire _w13960_ ;
	wire _w13961_ ;
	wire _w13962_ ;
	wire _w13963_ ;
	wire _w13964_ ;
	wire _w13965_ ;
	wire _w13966_ ;
	wire _w13967_ ;
	wire _w13968_ ;
	wire _w13969_ ;
	wire _w13970_ ;
	wire _w13971_ ;
	wire _w13972_ ;
	wire _w13973_ ;
	wire _w13974_ ;
	wire _w13975_ ;
	wire _w13976_ ;
	wire _w13977_ ;
	wire _w13978_ ;
	wire _w13979_ ;
	wire _w13980_ ;
	wire _w13981_ ;
	wire _w13982_ ;
	wire _w13983_ ;
	wire _w13984_ ;
	wire _w13985_ ;
	wire _w13986_ ;
	wire _w13987_ ;
	wire _w13988_ ;
	wire _w13989_ ;
	wire _w13990_ ;
	wire _w13991_ ;
	wire _w13992_ ;
	wire _w13993_ ;
	wire _w13994_ ;
	wire _w13995_ ;
	wire _w13996_ ;
	wire _w13997_ ;
	wire _w13998_ ;
	wire _w13999_ ;
	wire _w14000_ ;
	wire _w14001_ ;
	wire _w14002_ ;
	wire _w14003_ ;
	wire _w14004_ ;
	wire _w14005_ ;
	wire _w14006_ ;
	wire _w14007_ ;
	wire _w14008_ ;
	wire _w14009_ ;
	wire _w14010_ ;
	wire _w14011_ ;
	wire _w14012_ ;
	wire _w14013_ ;
	wire _w14014_ ;
	wire _w14015_ ;
	wire _w14016_ ;
	wire _w14017_ ;
	wire _w14018_ ;
	wire _w14019_ ;
	wire _w14020_ ;
	wire _w14021_ ;
	wire _w14022_ ;
	wire _w14023_ ;
	wire _w14024_ ;
	wire _w14025_ ;
	wire _w14026_ ;
	wire _w14027_ ;
	wire _w14028_ ;
	wire _w14029_ ;
	wire _w14030_ ;
	wire _w14031_ ;
	wire _w14032_ ;
	wire _w14033_ ;
	wire _w14034_ ;
	wire _w14035_ ;
	wire _w14036_ ;
	wire _w14037_ ;
	wire _w14038_ ;
	wire _w14039_ ;
	wire _w14040_ ;
	wire _w14041_ ;
	wire _w14042_ ;
	wire _w14043_ ;
	wire _w14044_ ;
	wire _w14045_ ;
	wire _w14046_ ;
	wire _w14047_ ;
	wire _w14048_ ;
	wire _w14049_ ;
	wire _w14050_ ;
	wire _w14051_ ;
	wire _w14052_ ;
	wire _w14053_ ;
	wire _w14054_ ;
	wire _w14055_ ;
	wire _w14056_ ;
	wire _w14057_ ;
	wire _w14058_ ;
	wire _w14059_ ;
	wire _w14060_ ;
	wire _w14061_ ;
	wire _w14062_ ;
	wire _w14063_ ;
	wire _w14064_ ;
	wire _w14065_ ;
	wire _w14066_ ;
	wire _w14067_ ;
	wire _w14068_ ;
	wire _w14069_ ;
	wire _w14070_ ;
	wire _w14071_ ;
	wire _w14072_ ;
	wire _w14073_ ;
	wire _w14074_ ;
	wire _w14075_ ;
	wire _w14076_ ;
	wire _w14077_ ;
	wire _w14078_ ;
	wire _w14079_ ;
	wire _w14080_ ;
	wire _w14081_ ;
	wire _w14082_ ;
	wire _w14083_ ;
	wire _w14084_ ;
	wire _w14085_ ;
	wire _w14086_ ;
	wire _w14087_ ;
	wire _w14088_ ;
	wire _w14089_ ;
	wire _w14090_ ;
	wire _w14091_ ;
	wire _w14092_ ;
	wire _w14093_ ;
	wire _w14094_ ;
	wire _w14095_ ;
	wire _w14096_ ;
	wire _w14097_ ;
	wire _w14098_ ;
	wire _w14099_ ;
	wire _w14100_ ;
	wire _w14101_ ;
	wire _w14102_ ;
	wire _w14103_ ;
	wire _w14104_ ;
	wire _w14105_ ;
	wire _w14106_ ;
	wire _w14107_ ;
	wire _w14108_ ;
	wire _w14109_ ;
	wire _w14110_ ;
	wire _w14111_ ;
	wire _w14112_ ;
	wire _w14113_ ;
	wire _w14114_ ;
	wire _w14115_ ;
	wire _w14116_ ;
	wire _w14117_ ;
	wire _w14118_ ;
	wire _w14119_ ;
	wire _w14120_ ;
	wire _w14121_ ;
	wire _w14122_ ;
	wire _w14123_ ;
	wire _w14124_ ;
	wire _w14125_ ;
	wire _w14126_ ;
	wire _w14127_ ;
	wire _w14128_ ;
	wire _w14129_ ;
	wire _w14130_ ;
	wire _w14131_ ;
	wire _w14132_ ;
	wire _w14133_ ;
	wire _w14134_ ;
	wire _w14135_ ;
	wire _w14136_ ;
	wire _w14137_ ;
	wire _w14138_ ;
	wire _w14139_ ;
	wire _w14140_ ;
	wire _w14141_ ;
	wire _w14142_ ;
	wire _w14143_ ;
	wire _w14144_ ;
	wire _w14145_ ;
	wire _w14146_ ;
	wire _w14147_ ;
	wire _w14148_ ;
	wire _w14149_ ;
	wire _w14150_ ;
	wire _w14151_ ;
	wire _w14152_ ;
	wire _w14153_ ;
	wire _w14154_ ;
	wire _w14155_ ;
	wire _w14156_ ;
	wire _w14157_ ;
	wire _w14158_ ;
	wire _w14159_ ;
	wire _w14160_ ;
	wire _w14161_ ;
	wire _w14162_ ;
	wire _w14163_ ;
	wire _w14164_ ;
	wire _w14165_ ;
	wire _w14166_ ;
	wire _w14167_ ;
	wire _w14168_ ;
	wire _w14169_ ;
	wire _w14170_ ;
	wire _w14171_ ;
	wire _w14172_ ;
	wire _w14173_ ;
	wire _w14174_ ;
	wire _w14175_ ;
	wire _w14176_ ;
	wire _w14177_ ;
	wire _w14178_ ;
	wire _w14179_ ;
	wire _w14180_ ;
	wire _w14181_ ;
	wire _w14182_ ;
	wire _w14183_ ;
	wire _w14184_ ;
	wire _w14185_ ;
	wire _w14186_ ;
	wire _w14187_ ;
	wire _w14188_ ;
	wire _w14189_ ;
	wire _w14190_ ;
	wire _w14191_ ;
	wire _w14192_ ;
	wire _w14193_ ;
	wire _w14194_ ;
	wire _w14195_ ;
	wire _w14196_ ;
	wire _w14197_ ;
	wire _w14198_ ;
	wire _w14199_ ;
	wire _w14200_ ;
	wire _w14201_ ;
	wire _w14202_ ;
	wire _w14203_ ;
	wire _w14204_ ;
	wire _w14205_ ;
	wire _w14206_ ;
	wire _w14207_ ;
	wire _w14208_ ;
	wire _w14209_ ;
	wire _w14210_ ;
	wire _w14211_ ;
	wire _w14212_ ;
	wire _w14213_ ;
	wire _w14214_ ;
	wire _w14215_ ;
	wire _w14216_ ;
	wire _w14217_ ;
	wire _w14218_ ;
	wire _w14219_ ;
	wire _w14220_ ;
	wire _w14221_ ;
	wire _w14222_ ;
	wire _w14223_ ;
	wire _w14224_ ;
	wire _w14225_ ;
	wire _w14226_ ;
	wire _w14227_ ;
	wire _w14228_ ;
	wire _w14229_ ;
	wire _w14230_ ;
	wire _w14231_ ;
	wire _w14232_ ;
	wire _w14233_ ;
	wire _w14234_ ;
	wire _w14235_ ;
	wire _w14236_ ;
	wire _w14237_ ;
	wire _w14238_ ;
	wire _w14239_ ;
	wire _w14240_ ;
	wire _w14241_ ;
	wire _w14242_ ;
	wire _w14243_ ;
	wire _w14244_ ;
	wire _w14245_ ;
	wire _w14246_ ;
	wire _w14247_ ;
	wire _w14248_ ;
	wire _w14249_ ;
	wire _w14250_ ;
	wire _w14251_ ;
	wire _w14252_ ;
	wire _w14253_ ;
	wire _w14254_ ;
	wire _w14255_ ;
	wire _w14256_ ;
	wire _w14257_ ;
	wire _w14258_ ;
	wire _w14259_ ;
	wire _w14260_ ;
	wire _w14261_ ;
	wire _w14262_ ;
	wire _w14263_ ;
	wire _w14264_ ;
	wire _w14265_ ;
	wire _w14266_ ;
	wire _w14267_ ;
	wire _w14268_ ;
	wire _w14269_ ;
	wire _w14270_ ;
	wire _w14271_ ;
	wire _w14272_ ;
	wire _w14273_ ;
	wire _w14274_ ;
	wire _w14275_ ;
	wire _w14276_ ;
	wire _w14277_ ;
	wire _w14278_ ;
	wire _w14279_ ;
	wire _w14280_ ;
	wire _w14281_ ;
	wire _w14282_ ;
	wire _w14283_ ;
	wire _w14284_ ;
	wire _w14285_ ;
	wire _w14286_ ;
	wire _w14287_ ;
	wire _w14288_ ;
	wire _w14289_ ;
	wire _w14290_ ;
	wire _w14291_ ;
	wire _w14292_ ;
	wire _w14293_ ;
	wire _w14294_ ;
	wire _w14295_ ;
	wire _w14296_ ;
	wire _w14297_ ;
	wire _w14298_ ;
	wire _w14299_ ;
	wire _w14300_ ;
	wire _w14301_ ;
	wire _w14302_ ;
	wire _w14303_ ;
	wire _w14304_ ;
	wire _w14305_ ;
	wire _w14306_ ;
	wire _w14307_ ;
	wire _w14308_ ;
	wire _w14309_ ;
	wire _w14310_ ;
	wire _w14311_ ;
	wire _w14312_ ;
	wire _w14313_ ;
	wire _w14314_ ;
	wire _w14315_ ;
	wire _w14316_ ;
	wire _w14317_ ;
	wire _w14318_ ;
	wire _w14319_ ;
	wire _w14320_ ;
	wire _w14321_ ;
	wire _w14322_ ;
	wire _w14323_ ;
	wire _w14324_ ;
	wire _w14325_ ;
	wire _w14326_ ;
	wire _w14327_ ;
	wire _w14328_ ;
	wire _w14329_ ;
	wire _w14330_ ;
	wire _w14331_ ;
	wire _w14332_ ;
	wire _w14333_ ;
	wire _w14334_ ;
	wire _w14335_ ;
	wire _w14336_ ;
	wire _w14337_ ;
	wire _w14338_ ;
	wire _w14339_ ;
	wire _w14340_ ;
	wire _w14341_ ;
	wire _w14342_ ;
	wire _w14343_ ;
	wire _w14344_ ;
	wire _w14345_ ;
	wire _w14346_ ;
	wire _w14347_ ;
	wire _w14348_ ;
	wire _w14349_ ;
	wire _w14350_ ;
	wire _w14351_ ;
	wire _w14352_ ;
	wire _w14353_ ;
	wire _w14354_ ;
	wire _w14355_ ;
	wire _w14356_ ;
	wire _w14357_ ;
	wire _w14358_ ;
	wire _w14359_ ;
	wire _w14360_ ;
	wire _w14361_ ;
	wire _w14362_ ;
	wire _w14363_ ;
	wire _w14364_ ;
	wire _w14365_ ;
	wire _w14366_ ;
	wire _w14367_ ;
	wire _w14368_ ;
	wire _w14369_ ;
	wire _w14370_ ;
	wire _w14371_ ;
	wire _w14372_ ;
	wire _w14373_ ;
	wire _w14374_ ;
	wire _w14375_ ;
	wire _w14376_ ;
	wire _w14377_ ;
	wire _w14378_ ;
	wire _w14379_ ;
	wire _w14380_ ;
	wire _w14381_ ;
	wire _w14382_ ;
	wire _w14383_ ;
	wire _w14384_ ;
	wire _w14385_ ;
	wire _w14386_ ;
	wire _w14387_ ;
	wire _w14388_ ;
	wire _w14389_ ;
	wire _w14390_ ;
	wire _w14391_ ;
	wire _w14392_ ;
	wire _w14393_ ;
	wire _w14394_ ;
	wire _w14395_ ;
	wire _w14396_ ;
	wire _w14397_ ;
	wire _w14398_ ;
	wire _w14399_ ;
	wire _w14400_ ;
	wire _w14401_ ;
	wire _w14402_ ;
	wire _w14403_ ;
	wire _w14404_ ;
	wire _w14405_ ;
	wire _w14406_ ;
	wire _w14407_ ;
	wire _w14408_ ;
	wire _w14409_ ;
	wire _w14410_ ;
	wire _w14411_ ;
	wire _w14412_ ;
	wire _w14413_ ;
	wire _w14414_ ;
	wire _w14415_ ;
	wire _w14416_ ;
	wire _w14417_ ;
	wire _w14418_ ;
	wire _w14419_ ;
	wire _w14420_ ;
	wire _w14421_ ;
	wire _w14422_ ;
	wire _w14423_ ;
	wire _w14424_ ;
	wire _w14425_ ;
	wire _w14426_ ;
	wire _w14427_ ;
	wire _w14428_ ;
	wire _w14429_ ;
	wire _w14430_ ;
	wire _w14431_ ;
	wire _w14432_ ;
	wire _w14433_ ;
	wire _w14434_ ;
	wire _w14435_ ;
	wire _w14436_ ;
	wire _w14437_ ;
	wire _w14438_ ;
	wire _w14439_ ;
	wire _w14440_ ;
	wire _w14441_ ;
	wire _w14442_ ;
	wire _w14443_ ;
	wire _w14444_ ;
	wire _w14445_ ;
	wire _w14446_ ;
	wire _w14447_ ;
	wire _w14448_ ;
	wire _w14449_ ;
	wire _w14450_ ;
	wire _w14451_ ;
	wire _w14452_ ;
	wire _w14453_ ;
	wire _w14454_ ;
	wire _w14455_ ;
	wire _w14456_ ;
	wire _w14457_ ;
	wire _w14458_ ;
	wire _w14459_ ;
	wire _w14460_ ;
	wire _w14461_ ;
	wire _w14462_ ;
	wire _w14463_ ;
	wire _w14464_ ;
	wire _w14465_ ;
	wire _w14466_ ;
	wire _w14467_ ;
	wire _w14468_ ;
	wire _w14469_ ;
	wire _w14470_ ;
	wire _w14471_ ;
	wire _w14472_ ;
	wire _w14473_ ;
	wire _w14474_ ;
	wire _w14475_ ;
	wire _w14476_ ;
	wire _w14477_ ;
	wire _w14478_ ;
	wire _w14479_ ;
	wire _w14480_ ;
	wire _w14481_ ;
	wire _w14482_ ;
	wire _w14483_ ;
	wire _w14484_ ;
	wire _w14485_ ;
	wire _w14486_ ;
	wire _w14487_ ;
	wire _w14488_ ;
	wire _w14489_ ;
	wire _w14490_ ;
	wire _w14491_ ;
	wire _w14492_ ;
	wire _w14493_ ;
	wire _w14494_ ;
	wire _w14495_ ;
	wire _w14496_ ;
	wire _w14497_ ;
	wire _w14498_ ;
	wire _w14499_ ;
	wire _w14500_ ;
	wire _w14501_ ;
	wire _w14502_ ;
	wire _w14503_ ;
	wire _w14504_ ;
	wire _w14505_ ;
	wire _w14506_ ;
	wire _w14507_ ;
	wire _w14508_ ;
	wire _w14509_ ;
	wire _w14510_ ;
	wire _w14511_ ;
	wire _w14512_ ;
	wire _w14513_ ;
	wire _w14514_ ;
	wire _w14515_ ;
	wire _w14516_ ;
	wire _w14517_ ;
	wire _w14518_ ;
	wire _w14519_ ;
	wire _w14520_ ;
	wire _w14521_ ;
	wire _w14522_ ;
	wire _w14523_ ;
	wire _w14524_ ;
	wire _w14525_ ;
	wire _w14526_ ;
	wire _w14527_ ;
	wire _w14528_ ;
	wire _w14529_ ;
	wire _w14530_ ;
	wire _w14531_ ;
	wire _w14532_ ;
	wire _w14533_ ;
	wire _w14534_ ;
	wire _w14535_ ;
	wire _w14536_ ;
	wire _w14537_ ;
	wire _w14538_ ;
	wire _w14539_ ;
	wire _w14540_ ;
	wire _w14541_ ;
	wire _w14542_ ;
	wire _w14543_ ;
	wire _w14544_ ;
	wire _w14545_ ;
	wire _w14546_ ;
	wire _w14547_ ;
	wire _w14548_ ;
	wire _w14549_ ;
	wire _w14550_ ;
	wire _w14551_ ;
	wire _w14552_ ;
	wire _w14553_ ;
	wire _w14554_ ;
	wire _w14555_ ;
	wire _w14556_ ;
	wire _w14557_ ;
	wire _w14558_ ;
	wire _w14559_ ;
	wire _w14560_ ;
	wire _w14561_ ;
	wire _w14562_ ;
	wire _w14563_ ;
	wire _w14564_ ;
	wire _w14565_ ;
	wire _w14566_ ;
	wire _w14567_ ;
	wire _w14568_ ;
	wire _w14569_ ;
	wire _w14570_ ;
	wire _w14571_ ;
	wire _w14572_ ;
	wire _w14573_ ;
	wire _w14574_ ;
	wire _w14575_ ;
	wire _w14576_ ;
	wire _w14577_ ;
	wire _w14578_ ;
	wire _w14579_ ;
	wire _w14580_ ;
	wire _w14581_ ;
	wire _w14582_ ;
	wire _w14583_ ;
	wire _w14584_ ;
	wire _w14585_ ;
	wire _w14586_ ;
	wire _w14587_ ;
	wire _w14588_ ;
	wire _w14589_ ;
	wire _w14590_ ;
	wire _w14591_ ;
	wire _w14592_ ;
	wire _w14593_ ;
	wire _w14594_ ;
	wire _w14595_ ;
	wire _w14596_ ;
	wire _w14597_ ;
	wire _w14598_ ;
	wire _w14599_ ;
	wire _w14600_ ;
	wire _w14601_ ;
	wire _w14602_ ;
	wire _w14603_ ;
	wire _w14604_ ;
	wire _w14605_ ;
	wire _w14606_ ;
	wire _w14607_ ;
	wire _w14608_ ;
	wire _w14609_ ;
	wire _w14610_ ;
	wire _w14611_ ;
	wire _w14612_ ;
	wire _w14613_ ;
	wire _w14614_ ;
	wire _w14615_ ;
	wire _w14616_ ;
	wire _w14617_ ;
	wire _w14618_ ;
	wire _w14619_ ;
	wire _w14620_ ;
	wire _w14621_ ;
	wire _w14622_ ;
	wire _w14623_ ;
	wire _w14624_ ;
	wire _w14625_ ;
	wire _w14626_ ;
	wire _w14627_ ;
	wire _w14628_ ;
	wire _w14629_ ;
	wire _w14630_ ;
	wire _w14631_ ;
	wire _w14632_ ;
	wire _w14633_ ;
	wire _w14634_ ;
	wire _w14635_ ;
	wire _w14636_ ;
	wire _w14637_ ;
	wire _w14638_ ;
	wire _w14639_ ;
	wire _w14640_ ;
	wire _w14641_ ;
	wire _w14642_ ;
	wire _w14643_ ;
	wire _w14644_ ;
	wire _w14645_ ;
	wire _w14646_ ;
	wire _w14647_ ;
	wire _w14648_ ;
	wire _w14649_ ;
	wire _w14650_ ;
	wire _w14651_ ;
	wire _w14652_ ;
	wire _w14653_ ;
	wire _w14654_ ;
	wire _w14655_ ;
	wire _w14656_ ;
	wire _w14657_ ;
	wire _w14658_ ;
	wire _w14659_ ;
	wire _w14660_ ;
	wire _w14661_ ;
	wire _w14662_ ;
	wire _w14663_ ;
	wire _w14664_ ;
	wire _w14665_ ;
	wire _w14666_ ;
	wire _w14667_ ;
	wire _w14668_ ;
	wire _w14669_ ;
	wire _w14670_ ;
	wire _w14671_ ;
	wire _w14672_ ;
	wire _w14673_ ;
	wire _w14674_ ;
	wire _w14675_ ;
	wire _w14676_ ;
	wire _w14677_ ;
	wire _w14678_ ;
	wire _w14679_ ;
	wire _w14680_ ;
	wire _w14681_ ;
	wire _w14682_ ;
	wire _w14683_ ;
	wire _w14684_ ;
	wire _w14685_ ;
	wire _w14686_ ;
	wire _w14687_ ;
	wire _w14688_ ;
	wire _w14689_ ;
	wire _w14690_ ;
	wire _w14691_ ;
	wire _w14692_ ;
	wire _w14693_ ;
	wire _w14694_ ;
	wire _w14695_ ;
	wire _w14696_ ;
	wire _w14697_ ;
	wire _w14698_ ;
	wire _w14699_ ;
	wire _w14700_ ;
	wire _w14701_ ;
	wire _w14702_ ;
	wire _w14703_ ;
	wire _w14704_ ;
	wire _w14705_ ;
	wire _w14706_ ;
	wire _w14707_ ;
	wire _w14708_ ;
	wire _w14709_ ;
	wire _w14710_ ;
	wire _w14711_ ;
	wire _w14712_ ;
	wire _w14713_ ;
	wire _w14714_ ;
	wire _w14715_ ;
	wire _w14716_ ;
	wire _w14717_ ;
	wire _w14718_ ;
	wire _w14719_ ;
	wire _w14720_ ;
	wire _w14721_ ;
	wire _w14722_ ;
	wire _w14723_ ;
	wire _w14724_ ;
	wire _w14725_ ;
	wire _w14726_ ;
	wire _w14727_ ;
	wire _w14728_ ;
	wire _w14729_ ;
	wire _w14730_ ;
	wire _w14731_ ;
	wire _w14732_ ;
	wire _w14733_ ;
	wire _w14734_ ;
	wire _w14735_ ;
	wire _w14736_ ;
	wire _w14737_ ;
	wire _w14738_ ;
	wire _w14739_ ;
	wire _w14740_ ;
	wire _w14741_ ;
	wire _w14742_ ;
	wire _w14743_ ;
	wire _w14744_ ;
	wire _w14745_ ;
	wire _w14746_ ;
	wire _w14747_ ;
	wire _w14748_ ;
	wire _w14749_ ;
	wire _w14750_ ;
	wire _w14751_ ;
	wire _w14752_ ;
	wire _w14753_ ;
	wire _w14754_ ;
	wire _w14755_ ;
	wire _w14756_ ;
	wire _w14757_ ;
	wire _w14758_ ;
	wire _w14759_ ;
	wire _w14760_ ;
	wire _w14761_ ;
	wire _w14762_ ;
	wire _w14763_ ;
	wire _w14764_ ;
	wire _w14765_ ;
	wire _w14766_ ;
	wire _w14767_ ;
	wire _w14768_ ;
	wire _w14769_ ;
	wire _w14770_ ;
	wire _w14771_ ;
	wire _w14772_ ;
	wire _w14773_ ;
	wire _w14774_ ;
	wire _w14775_ ;
	wire _w14776_ ;
	wire _w14777_ ;
	wire _w14778_ ;
	wire _w14779_ ;
	wire _w14780_ ;
	wire _w14781_ ;
	wire _w14782_ ;
	wire _w14783_ ;
	wire _w14784_ ;
	wire _w14785_ ;
	wire _w14786_ ;
	wire _w14787_ ;
	wire _w14788_ ;
	wire _w14789_ ;
	wire _w14790_ ;
	wire _w14791_ ;
	wire _w14792_ ;
	wire _w14793_ ;
	wire _w14794_ ;
	wire _w14795_ ;
	wire _w14796_ ;
	wire _w14797_ ;
	wire _w14798_ ;
	wire _w14799_ ;
	wire _w14800_ ;
	wire _w14801_ ;
	wire _w14802_ ;
	wire _w14803_ ;
	wire _w14804_ ;
	wire _w14805_ ;
	wire _w14806_ ;
	wire _w14807_ ;
	wire _w14808_ ;
	wire _w14809_ ;
	wire _w14810_ ;
	wire _w14811_ ;
	wire _w14812_ ;
	wire _w14813_ ;
	wire _w14814_ ;
	wire _w14815_ ;
	wire _w14816_ ;
	wire _w14817_ ;
	wire _w14818_ ;
	wire _w14819_ ;
	wire _w14820_ ;
	wire _w14821_ ;
	wire _w14822_ ;
	wire _w14823_ ;
	wire _w14824_ ;
	wire _w14825_ ;
	wire _w14826_ ;
	wire _w14827_ ;
	wire _w14828_ ;
	wire _w14829_ ;
	wire _w14830_ ;
	wire _w14831_ ;
	wire _w14832_ ;
	wire _w14833_ ;
	wire _w14834_ ;
	wire _w14835_ ;
	wire _w14836_ ;
	wire _w14837_ ;
	wire _w14838_ ;
	wire _w14839_ ;
	wire _w14840_ ;
	wire _w14841_ ;
	wire _w14842_ ;
	wire _w14843_ ;
	wire _w14844_ ;
	wire _w14845_ ;
	wire _w14846_ ;
	wire _w14847_ ;
	wire _w14848_ ;
	wire _w14849_ ;
	wire _w14850_ ;
	wire _w14851_ ;
	wire _w14852_ ;
	wire _w14853_ ;
	wire _w14854_ ;
	wire _w14855_ ;
	wire _w14856_ ;
	wire _w14857_ ;
	wire _w14858_ ;
	wire _w14859_ ;
	wire _w14860_ ;
	wire _w14861_ ;
	wire _w14862_ ;
	wire _w14863_ ;
	wire _w14864_ ;
	wire _w14865_ ;
	wire _w14866_ ;
	wire _w14867_ ;
	wire _w14868_ ;
	wire _w14869_ ;
	wire _w14870_ ;
	wire _w14871_ ;
	wire _w14872_ ;
	wire _w14873_ ;
	wire _w14874_ ;
	wire _w14875_ ;
	wire _w14876_ ;
	wire _w14877_ ;
	wire _w14878_ ;
	wire _w14879_ ;
	wire _w14880_ ;
	wire _w14881_ ;
	wire _w14882_ ;
	wire _w14883_ ;
	wire _w14884_ ;
	wire _w14885_ ;
	wire _w14886_ ;
	wire _w14887_ ;
	wire _w14888_ ;
	wire _w14889_ ;
	wire _w14890_ ;
	wire _w14891_ ;
	wire _w14892_ ;
	wire _w14893_ ;
	wire _w14894_ ;
	wire _w14895_ ;
	wire _w14896_ ;
	wire _w14897_ ;
	wire _w14898_ ;
	wire _w14899_ ;
	wire _w14900_ ;
	wire _w14901_ ;
	wire _w14902_ ;
	wire _w14903_ ;
	wire _w14904_ ;
	wire _w14905_ ;
	wire _w14906_ ;
	wire _w14907_ ;
	wire _w14908_ ;
	wire _w14909_ ;
	wire _w14910_ ;
	wire _w14911_ ;
	wire _w14912_ ;
	wire _w14913_ ;
	wire _w14914_ ;
	wire _w14915_ ;
	wire _w14916_ ;
	wire _w14917_ ;
	wire _w14918_ ;
	wire _w14919_ ;
	wire _w14920_ ;
	wire _w14921_ ;
	wire _w14922_ ;
	wire _w14923_ ;
	wire _w14924_ ;
	wire _w14925_ ;
	wire _w14926_ ;
	wire _w14927_ ;
	wire _w14928_ ;
	wire _w14929_ ;
	wire _w14930_ ;
	wire _w14931_ ;
	wire _w14932_ ;
	wire _w14933_ ;
	wire _w14934_ ;
	wire _w14935_ ;
	wire _w14936_ ;
	wire _w14937_ ;
	wire _w14938_ ;
	wire _w14939_ ;
	wire _w14940_ ;
	wire _w14941_ ;
	wire _w14942_ ;
	wire _w14943_ ;
	wire _w14944_ ;
	wire _w14945_ ;
	wire _w14946_ ;
	wire _w14947_ ;
	wire _w14948_ ;
	wire _w14949_ ;
	wire _w14950_ ;
	wire _w14951_ ;
	wire _w14952_ ;
	wire _w14953_ ;
	wire _w14954_ ;
	wire _w14955_ ;
	wire _w14956_ ;
	wire _w14957_ ;
	wire _w14958_ ;
	wire _w14959_ ;
	wire _w14960_ ;
	wire _w14961_ ;
	wire _w14962_ ;
	wire _w14963_ ;
	wire _w14964_ ;
	wire _w14965_ ;
	wire _w14966_ ;
	wire _w14967_ ;
	wire _w14968_ ;
	wire _w14969_ ;
	wire _w14970_ ;
	wire _w14971_ ;
	wire _w14972_ ;
	wire _w14973_ ;
	wire _w14974_ ;
	wire _w14975_ ;
	wire _w14976_ ;
	wire _w14977_ ;
	wire _w14978_ ;
	wire _w14979_ ;
	wire _w14980_ ;
	wire _w14981_ ;
	wire _w14982_ ;
	wire _w14983_ ;
	wire _w14984_ ;
	wire _w14985_ ;
	wire _w14986_ ;
	wire _w14987_ ;
	wire _w14988_ ;
	wire _w14989_ ;
	wire _w14990_ ;
	wire _w14991_ ;
	wire _w14992_ ;
	wire _w14993_ ;
	wire _w14994_ ;
	wire _w14995_ ;
	wire _w14996_ ;
	wire _w14997_ ;
	wire _w14998_ ;
	wire _w14999_ ;
	wire _w15000_ ;
	wire _w15001_ ;
	wire _w15002_ ;
	wire _w15003_ ;
	wire _w15004_ ;
	wire _w15005_ ;
	wire _w15006_ ;
	wire _w15007_ ;
	wire _w15008_ ;
	wire _w15009_ ;
	wire _w15010_ ;
	wire _w15011_ ;
	wire _w15012_ ;
	wire _w15013_ ;
	wire _w15014_ ;
	wire _w15015_ ;
	wire _w15016_ ;
	wire _w15017_ ;
	wire _w15018_ ;
	wire _w15019_ ;
	wire _w15020_ ;
	wire _w15021_ ;
	wire _w15022_ ;
	wire _w15023_ ;
	wire _w15024_ ;
	wire _w15025_ ;
	wire _w15026_ ;
	wire _w15027_ ;
	wire _w15028_ ;
	wire _w15029_ ;
	wire _w15030_ ;
	wire _w15031_ ;
	wire _w15032_ ;
	wire _w15033_ ;
	wire _w15034_ ;
	wire _w15035_ ;
	wire _w15036_ ;
	wire _w15037_ ;
	wire _w15038_ ;
	wire _w15039_ ;
	wire _w15040_ ;
	wire _w15041_ ;
	wire _w15042_ ;
	wire _w15043_ ;
	wire _w15044_ ;
	wire _w15045_ ;
	wire _w15046_ ;
	wire _w15047_ ;
	wire _w15048_ ;
	wire _w15049_ ;
	wire _w15050_ ;
	wire _w15051_ ;
	wire _w15052_ ;
	wire _w15053_ ;
	wire _w15054_ ;
	wire _w15055_ ;
	wire _w15056_ ;
	wire _w15057_ ;
	wire _w15058_ ;
	wire _w15059_ ;
	wire _w15060_ ;
	wire _w15061_ ;
	wire _w15062_ ;
	wire _w15063_ ;
	wire _w15064_ ;
	wire _w15065_ ;
	wire _w15066_ ;
	wire _w15067_ ;
	wire _w15068_ ;
	wire _w15069_ ;
	wire _w15070_ ;
	wire _w15071_ ;
	wire _w15072_ ;
	wire _w15073_ ;
	wire _w15074_ ;
	wire _w15075_ ;
	wire _w15076_ ;
	wire _w15077_ ;
	wire _w15078_ ;
	wire _w15079_ ;
	wire _w15080_ ;
	wire _w15081_ ;
	wire _w15082_ ;
	wire _w15083_ ;
	wire _w15084_ ;
	wire _w15085_ ;
	wire _w15086_ ;
	wire _w15087_ ;
	wire _w15088_ ;
	wire _w15089_ ;
	wire _w15090_ ;
	wire _w15091_ ;
	wire _w15092_ ;
	wire _w15093_ ;
	wire _w15094_ ;
	wire _w15095_ ;
	wire _w15096_ ;
	wire _w15097_ ;
	wire _w15098_ ;
	wire _w15099_ ;
	wire _w15100_ ;
	wire _w15101_ ;
	wire _w15102_ ;
	wire _w15103_ ;
	wire _w15104_ ;
	wire _w15105_ ;
	wire _w15106_ ;
	wire _w15107_ ;
	wire _w15108_ ;
	wire _w15109_ ;
	wire _w15110_ ;
	wire _w15111_ ;
	wire _w15112_ ;
	wire _w15113_ ;
	wire _w15114_ ;
	wire _w15115_ ;
	wire _w15116_ ;
	wire _w15117_ ;
	wire _w15118_ ;
	wire _w15119_ ;
	wire _w15120_ ;
	wire _w15121_ ;
	wire _w15122_ ;
	wire _w15123_ ;
	wire _w15124_ ;
	wire _w15125_ ;
	wire _w15126_ ;
	wire _w15127_ ;
	wire _w15128_ ;
	wire _w15129_ ;
	wire _w15130_ ;
	wire _w15131_ ;
	wire _w15132_ ;
	wire _w15133_ ;
	wire _w15134_ ;
	wire _w15135_ ;
	wire _w15136_ ;
	wire _w15137_ ;
	wire _w15138_ ;
	wire _w15139_ ;
	wire _w15140_ ;
	wire _w15141_ ;
	wire _w15142_ ;
	wire _w15143_ ;
	wire _w15144_ ;
	wire _w15145_ ;
	wire _w15146_ ;
	wire _w15147_ ;
	wire _w15148_ ;
	wire _w15149_ ;
	wire _w15150_ ;
	wire _w15151_ ;
	wire _w15152_ ;
	wire _w15153_ ;
	wire _w15154_ ;
	wire _w15155_ ;
	wire _w15156_ ;
	wire _w15157_ ;
	wire _w15158_ ;
	wire _w15159_ ;
	wire _w15160_ ;
	wire _w15161_ ;
	wire _w15162_ ;
	wire _w15163_ ;
	wire _w15164_ ;
	wire _w15165_ ;
	wire _w15166_ ;
	wire _w15167_ ;
	wire _w15168_ ;
	wire _w15169_ ;
	wire _w15170_ ;
	wire _w15171_ ;
	wire _w15172_ ;
	wire _w15173_ ;
	wire _w15174_ ;
	wire _w15175_ ;
	wire _w15176_ ;
	wire _w15177_ ;
	wire _w15178_ ;
	wire _w15179_ ;
	wire _w15180_ ;
	wire _w15181_ ;
	wire _w15182_ ;
	wire _w15183_ ;
	wire _w15184_ ;
	wire _w15185_ ;
	wire _w15186_ ;
	wire _w15187_ ;
	wire _w15188_ ;
	wire _w15189_ ;
	wire _w15190_ ;
	wire _w15191_ ;
	wire _w15192_ ;
	wire _w15193_ ;
	wire _w15194_ ;
	wire _w15195_ ;
	wire _w15196_ ;
	wire _w15197_ ;
	wire _w15198_ ;
	wire _w15199_ ;
	wire _w15200_ ;
	wire _w15201_ ;
	wire _w15202_ ;
	wire _w15203_ ;
	wire _w15204_ ;
	wire _w15205_ ;
	wire _w15206_ ;
	wire _w15207_ ;
	wire _w15208_ ;
	wire _w15209_ ;
	wire _w15210_ ;
	wire _w15211_ ;
	wire _w15212_ ;
	wire _w15213_ ;
	wire _w15214_ ;
	wire _w15215_ ;
	wire _w15216_ ;
	wire _w15217_ ;
	wire _w15218_ ;
	wire _w15219_ ;
	wire _w15220_ ;
	wire _w15221_ ;
	wire _w15222_ ;
	wire _w15223_ ;
	wire _w15224_ ;
	wire _w15225_ ;
	wire _w15226_ ;
	wire _w15227_ ;
	wire _w15228_ ;
	wire _w15229_ ;
	wire _w15230_ ;
	wire _w15231_ ;
	wire _w15232_ ;
	wire _w15233_ ;
	wire _w15234_ ;
	wire _w15235_ ;
	wire _w15236_ ;
	wire _w15237_ ;
	wire _w15238_ ;
	wire _w15239_ ;
	wire _w15240_ ;
	wire _w15241_ ;
	wire _w15242_ ;
	wire _w15243_ ;
	wire _w15244_ ;
	wire _w15245_ ;
	wire _w15246_ ;
	wire _w15247_ ;
	wire _w15248_ ;
	wire _w15249_ ;
	wire _w15250_ ;
	wire _w15251_ ;
	wire _w15252_ ;
	wire _w15253_ ;
	wire _w15254_ ;
	wire _w15255_ ;
	wire _w15256_ ;
	wire _w15257_ ;
	wire _w15258_ ;
	wire _w15259_ ;
	wire _w15260_ ;
	wire _w15261_ ;
	wire _w15262_ ;
	wire _w15263_ ;
	wire _w15264_ ;
	wire _w15265_ ;
	wire _w15266_ ;
	wire _w15267_ ;
	wire _w15268_ ;
	wire _w15269_ ;
	wire _w15270_ ;
	wire _w15271_ ;
	wire _w15272_ ;
	wire _w15273_ ;
	wire _w15274_ ;
	wire _w15275_ ;
	wire _w15276_ ;
	wire _w15277_ ;
	wire _w15278_ ;
	wire _w15279_ ;
	wire _w15280_ ;
	wire _w15281_ ;
	wire _w15282_ ;
	wire _w15283_ ;
	wire _w15284_ ;
	wire _w15285_ ;
	wire _w15286_ ;
	wire _w15287_ ;
	wire _w15288_ ;
	wire _w15289_ ;
	wire _w15290_ ;
	wire _w15291_ ;
	wire _w15292_ ;
	wire _w15293_ ;
	wire _w15294_ ;
	wire _w15295_ ;
	wire _w15296_ ;
	wire _w15297_ ;
	wire _w15298_ ;
	wire _w15299_ ;
	wire _w15300_ ;
	wire _w15301_ ;
	wire _w15302_ ;
	wire _w15303_ ;
	wire _w15304_ ;
	wire _w15305_ ;
	wire _w15306_ ;
	wire _w15307_ ;
	wire _w15308_ ;
	wire _w15309_ ;
	wire _w15310_ ;
	wire _w15311_ ;
	wire _w15312_ ;
	wire _w15313_ ;
	wire _w15314_ ;
	wire _w15315_ ;
	wire _w15316_ ;
	wire _w15317_ ;
	wire _w15318_ ;
	wire _w15319_ ;
	wire _w15320_ ;
	wire _w15321_ ;
	wire _w15322_ ;
	wire _w15323_ ;
	wire _w15324_ ;
	wire _w15325_ ;
	wire _w15326_ ;
	wire _w15327_ ;
	wire _w15328_ ;
	wire _w15329_ ;
	wire _w15330_ ;
	wire _w15331_ ;
	wire _w15332_ ;
	wire _w15333_ ;
	wire _w15334_ ;
	wire _w15335_ ;
	wire _w15336_ ;
	wire _w15337_ ;
	wire _w15338_ ;
	wire _w15339_ ;
	wire _w15340_ ;
	wire _w15341_ ;
	wire _w15342_ ;
	wire _w15343_ ;
	wire _w15344_ ;
	wire _w15345_ ;
	wire _w15346_ ;
	wire _w15347_ ;
	wire _w15348_ ;
	wire _w15349_ ;
	wire _w15350_ ;
	wire _w15351_ ;
	wire _w15352_ ;
	wire _w15353_ ;
	wire _w15354_ ;
	wire _w15355_ ;
	wire _w15356_ ;
	wire _w15357_ ;
	wire _w15358_ ;
	wire _w15359_ ;
	wire _w15360_ ;
	wire _w15361_ ;
	wire _w15362_ ;
	wire _w15363_ ;
	wire _w15364_ ;
	wire _w15365_ ;
	wire _w15366_ ;
	wire _w15367_ ;
	wire _w15368_ ;
	wire _w15369_ ;
	wire _w15370_ ;
	wire _w15371_ ;
	wire _w15372_ ;
	wire _w15373_ ;
	wire _w15374_ ;
	wire _w15375_ ;
	wire _w15376_ ;
	wire _w15377_ ;
	wire _w15378_ ;
	wire _w15379_ ;
	wire _w15380_ ;
	wire _w15381_ ;
	wire _w15382_ ;
	wire _w15383_ ;
	wire _w15384_ ;
	wire _w15385_ ;
	wire _w15386_ ;
	wire _w15387_ ;
	wire _w15388_ ;
	wire _w15389_ ;
	wire _w15390_ ;
	wire _w15391_ ;
	wire _w15392_ ;
	wire _w15393_ ;
	wire _w15394_ ;
	wire _w15395_ ;
	wire _w15396_ ;
	wire _w15397_ ;
	wire _w15398_ ;
	wire _w15399_ ;
	wire _w15400_ ;
	wire _w15401_ ;
	wire _w15402_ ;
	wire _w15403_ ;
	wire _w15404_ ;
	wire _w15405_ ;
	wire _w15406_ ;
	wire _w15407_ ;
	wire _w15408_ ;
	wire _w15409_ ;
	wire _w15410_ ;
	wire _w15411_ ;
	wire _w15412_ ;
	wire _w15413_ ;
	wire _w15414_ ;
	wire _w15415_ ;
	wire _w15416_ ;
	wire _w15417_ ;
	wire _w15418_ ;
	wire _w15419_ ;
	wire _w15420_ ;
	wire _w15421_ ;
	wire _w15422_ ;
	wire _w15423_ ;
	wire _w15424_ ;
	wire _w15425_ ;
	wire _w15426_ ;
	wire _w15427_ ;
	wire _w15428_ ;
	wire _w15429_ ;
	wire _w15430_ ;
	wire _w15431_ ;
	wire _w15432_ ;
	wire _w15433_ ;
	wire _w15434_ ;
	wire _w15435_ ;
	wire _w15436_ ;
	wire _w15437_ ;
	wire _w15438_ ;
	wire _w15439_ ;
	wire _w15440_ ;
	wire _w15441_ ;
	wire _w15442_ ;
	wire _w15443_ ;
	wire _w15444_ ;
	wire _w15445_ ;
	wire _w15446_ ;
	wire _w15447_ ;
	wire _w15448_ ;
	wire _w15449_ ;
	wire _w15450_ ;
	wire _w15451_ ;
	wire _w15452_ ;
	wire _w15453_ ;
	wire _w15454_ ;
	wire _w15455_ ;
	wire _w15456_ ;
	wire _w15457_ ;
	wire _w15458_ ;
	wire _w15459_ ;
	wire _w15460_ ;
	wire _w15461_ ;
	wire _w15462_ ;
	wire _w15463_ ;
	wire _w15464_ ;
	wire _w15465_ ;
	wire _w15466_ ;
	wire _w15467_ ;
	wire _w15468_ ;
	wire _w15469_ ;
	wire _w15470_ ;
	wire _w15471_ ;
	wire _w15472_ ;
	wire _w15473_ ;
	wire _w15474_ ;
	wire _w15475_ ;
	wire _w15476_ ;
	wire _w15477_ ;
	wire _w15478_ ;
	wire _w15479_ ;
	wire _w15480_ ;
	wire _w15481_ ;
	wire _w15482_ ;
	wire _w15483_ ;
	wire _w15484_ ;
	wire _w15485_ ;
	wire _w15486_ ;
	wire _w15487_ ;
	wire _w15488_ ;
	wire _w15489_ ;
	wire _w15490_ ;
	wire _w15491_ ;
	wire _w15492_ ;
	wire _w15493_ ;
	wire _w15494_ ;
	wire _w15495_ ;
	wire _w15496_ ;
	wire _w15497_ ;
	wire _w15498_ ;
	wire _w15499_ ;
	wire _w15500_ ;
	wire _w15501_ ;
	wire _w15502_ ;
	wire _w15503_ ;
	wire _w15504_ ;
	wire _w15505_ ;
	wire _w15506_ ;
	wire _w15507_ ;
	wire _w15508_ ;
	wire _w15509_ ;
	wire _w15510_ ;
	wire _w15511_ ;
	wire _w15512_ ;
	wire _w15513_ ;
	wire _w15514_ ;
	wire _w15515_ ;
	wire _w15516_ ;
	wire _w15517_ ;
	wire _w15518_ ;
	wire _w15519_ ;
	wire _w15520_ ;
	wire _w15521_ ;
	wire _w15522_ ;
	wire _w15523_ ;
	wire _w15524_ ;
	wire _w15525_ ;
	wire _w15526_ ;
	wire _w15527_ ;
	wire _w15528_ ;
	wire _w15529_ ;
	wire _w15530_ ;
	wire _w15531_ ;
	wire _w15532_ ;
	wire _w15533_ ;
	wire _w15534_ ;
	wire _w15535_ ;
	wire _w15536_ ;
	wire _w15537_ ;
	wire _w15538_ ;
	wire _w15539_ ;
	wire _w15540_ ;
	wire _w15541_ ;
	wire _w15542_ ;
	wire _w15543_ ;
	wire _w15544_ ;
	wire _w15545_ ;
	wire _w15546_ ;
	wire _w15547_ ;
	wire _w15548_ ;
	wire _w15549_ ;
	wire _w15550_ ;
	wire _w15551_ ;
	wire _w15552_ ;
	wire _w15553_ ;
	wire _w15554_ ;
	wire _w15555_ ;
	wire _w15556_ ;
	wire _w15557_ ;
	wire _w15558_ ;
	wire _w15559_ ;
	wire _w15560_ ;
	wire _w15561_ ;
	wire _w15562_ ;
	wire _w15563_ ;
	wire _w15564_ ;
	wire _w15565_ ;
	wire _w15566_ ;
	wire _w15567_ ;
	wire _w15568_ ;
	wire _w15569_ ;
	wire _w15570_ ;
	wire _w15571_ ;
	wire _w15572_ ;
	wire _w15573_ ;
	wire _w15574_ ;
	wire _w15575_ ;
	wire _w15576_ ;
	wire _w15577_ ;
	wire _w15578_ ;
	wire _w15579_ ;
	wire _w15580_ ;
	wire _w15581_ ;
	wire _w15582_ ;
	wire _w15583_ ;
	wire _w15584_ ;
	wire _w15585_ ;
	wire _w15586_ ;
	wire _w15587_ ;
	wire _w15588_ ;
	wire _w15589_ ;
	wire _w15590_ ;
	wire _w15591_ ;
	wire _w15592_ ;
	wire _w15593_ ;
	wire _w15594_ ;
	wire _w15595_ ;
	wire _w15596_ ;
	wire _w15597_ ;
	wire _w15598_ ;
	wire _w20785_ ;
	wire _w20786_ ;
	wire _w20787_ ;
	wire _w20788_ ;
	wire _w20789_ ;
	wire _w20790_ ;
	wire _w20791_ ;
	wire _w20792_ ;
	wire _w20793_ ;
	wire _w20794_ ;
	wire _w20795_ ;
	wire _w20796_ ;
	wire _w20797_ ;
	wire _w20798_ ;
	wire _w20799_ ;
	wire _w20800_ ;
	wire _w20801_ ;
	wire _w20802_ ;
	wire _w20803_ ;
	wire _w20804_ ;
	wire _w20805_ ;
	wire _w20806_ ;
	wire _w20807_ ;
	wire _w20808_ ;
	wire _w20809_ ;
	wire _w20810_ ;
	wire _w20811_ ;
	wire _w20812_ ;
	wire _w20813_ ;
	wire _w20814_ ;
	wire _w20815_ ;
	wire _w20816_ ;
	wire _w20817_ ;
	wire _w20818_ ;
	wire _w20819_ ;
	wire _w20820_ ;
	wire _w20821_ ;
	wire _w20822_ ;
	wire _w20823_ ;
	wire _w20824_ ;
	wire _w20825_ ;
	wire _w20826_ ;
	wire _w20827_ ;
	wire _w20828_ ;
	wire _w20829_ ;
	wire _w20830_ ;
	wire _w20831_ ;
	wire _w20832_ ;
	wire _w20833_ ;
	wire _w20834_ ;
	wire _w20835_ ;
	wire _w20836_ ;
	wire _w20837_ ;
	wire _w20838_ ;
	wire _w20839_ ;
	wire _w20840_ ;
	wire _w20841_ ;
	wire _w20842_ ;
	wire _w20843_ ;
	wire _w20844_ ;
	wire _w20845_ ;
	wire _w20846_ ;
	wire _w20847_ ;
	wire _w20848_ ;
	wire _w20849_ ;
	wire _w20850_ ;
	wire _w20851_ ;
	wire _w20852_ ;
	wire _w20853_ ;
	wire _w20854_ ;
	wire _w20855_ ;
	wire _w20856_ ;
	wire _w20857_ ;
	wire _w20858_ ;
	wire _w20859_ ;
	wire _w20860_ ;
	wire _w20861_ ;
	wire _w20862_ ;
	wire _w20863_ ;
	wire _w20864_ ;
	wire _w20865_ ;
	wire _w20866_ ;
	wire _w20867_ ;
	wire _w20868_ ;
	wire _w20869_ ;
	wire _w20870_ ;
	wire _w20871_ ;
	wire _w20872_ ;
	wire _w20873_ ;
	wire _w20874_ ;
	wire _w20875_ ;
	wire _w20876_ ;
	wire _w20877_ ;
	wire _w20878_ ;
	wire _w20879_ ;
	wire _w20880_ ;
	wire _w20881_ ;
	wire _w20882_ ;
	wire _w20883_ ;
	wire _w20884_ ;
	wire _w20885_ ;
	wire _w20886_ ;
	wire _w20887_ ;
	wire _w20888_ ;
	wire _w20889_ ;
	wire _w20890_ ;
	wire _w20891_ ;
	wire _w20892_ ;
	wire _w20893_ ;
	wire _w20894_ ;
	wire _w20895_ ;
	wire _w20896_ ;
	wire _w20897_ ;
	wire _w20898_ ;
	wire _w20899_ ;
	wire _w20900_ ;
	wire _w20901_ ;
	wire _w20902_ ;
	wire _w20903_ ;
	wire _w20904_ ;
	wire _w20905_ ;
	wire _w20906_ ;
	wire _w20907_ ;
	wire _w20908_ ;
	wire _w20909_ ;
	wire _w20910_ ;
	wire _w20911_ ;
	wire _w20912_ ;
	wire _w20913_ ;
	wire _w20914_ ;
	wire _w20915_ ;
	wire _w20916_ ;
	wire _w20917_ ;
	wire _w20918_ ;
	wire _w20919_ ;
	wire _w20920_ ;
	wire _w20921_ ;
	wire _w20922_ ;
	wire _w20923_ ;
	wire _w20924_ ;
	wire _w20925_ ;
	wire _w20926_ ;
	wire _w20927_ ;
	wire _w20928_ ;
	wire _w20929_ ;
	wire _w20930_ ;
	wire _w20931_ ;
	wire _w20932_ ;
	wire _w20933_ ;
	wire _w20934_ ;
	wire _w20935_ ;
	wire _w20936_ ;
	wire _w20937_ ;
	wire _w20938_ ;
	wire _w20939_ ;
	wire _w20940_ ;
	wire _w20941_ ;
	wire _w20942_ ;
	wire _w20943_ ;
	wire _w20944_ ;
	wire _w20945_ ;
	wire _w20946_ ;
	wire _w20947_ ;
	wire _w20948_ ;
	wire _w20949_ ;
	wire _w20950_ ;
	wire _w20951_ ;
	wire _w20952_ ;
	wire _w20953_ ;
	wire _w20954_ ;
	wire _w20955_ ;
	wire _w20956_ ;
	wire _w20957_ ;
	wire _w20958_ ;
	wire _w20959_ ;
	wire _w20960_ ;
	wire _w20961_ ;
	wire _w20962_ ;
	wire _w20963_ ;
	wire _w20964_ ;
	wire _w20965_ ;
	wire _w20966_ ;
	wire _w20967_ ;
	wire _w20968_ ;
	wire _w20969_ ;
	wire _w20970_ ;
	wire _w20971_ ;
	wire _w20972_ ;
	wire _w20973_ ;
	wire _w20974_ ;
	wire _w20975_ ;
	wire _w20976_ ;
	wire _w20977_ ;
	wire _w20978_ ;
	wire _w20979_ ;
	wire _w20980_ ;
	wire _w20981_ ;
	wire _w20982_ ;
	wire _w20983_ ;
	wire _w20984_ ;
	wire _w20985_ ;
	wire _w20986_ ;
	wire _w20987_ ;
	wire _w20988_ ;
	wire _w20989_ ;
	wire _w20990_ ;
	wire _w20991_ ;
	wire _w20992_ ;
	wire _w20993_ ;
	wire _w20994_ ;
	wire _w20995_ ;
	wire _w20996_ ;
	wire _w20997_ ;
	wire _w20998_ ;
	wire _w20999_ ;
	wire _w21000_ ;
	wire _w21001_ ;
	wire _w21002_ ;
	wire _w21003_ ;
	wire _w21004_ ;
	wire _w21005_ ;
	wire _w21006_ ;
	wire _w21007_ ;
	wire _w21008_ ;
	wire _w21009_ ;
	wire _w21010_ ;
	wire _w21011_ ;
	wire _w21012_ ;
	wire _w21013_ ;
	wire _w21014_ ;
	wire _w21015_ ;
	wire _w21016_ ;
	wire _w21017_ ;
	wire _w21018_ ;
	wire _w21019_ ;
	wire _w21020_ ;
	wire _w21021_ ;
	wire _w21022_ ;
	wire _w21023_ ;
	wire _w21024_ ;
	wire _w21025_ ;
	wire _w21026_ ;
	wire _w21027_ ;
	wire _w21028_ ;
	wire _w21029_ ;
	wire _w21030_ ;
	wire _w21031_ ;
	wire _w21032_ ;
	wire _w21033_ ;
	wire _w21034_ ;
	wire _w21035_ ;
	wire _w21036_ ;
	wire _w21037_ ;
	wire _w21038_ ;
	wire _w21039_ ;
	wire _w21040_ ;
	wire _w21041_ ;
	wire _w21042_ ;
	wire _w21043_ ;
	wire _w21044_ ;
	wire _w21045_ ;
	wire _w21046_ ;
	wire _w21047_ ;
	wire _w21048_ ;
	wire _w21049_ ;
	wire _w21050_ ;
	wire _w21051_ ;
	wire _w21052_ ;
	wire _w21053_ ;
	wire _w21054_ ;
	wire _w21055_ ;
	wire _w21056_ ;
	wire _w21057_ ;
	wire _w21058_ ;
	wire _w21059_ ;
	wire _w21060_ ;
	wire _w21061_ ;
	wire _w21062_ ;
	wire _w21063_ ;
	wire _w21064_ ;
	wire _w21065_ ;
	wire _w21066_ ;
	wire _w21067_ ;
	wire _w21068_ ;
	wire _w21069_ ;
	wire _w21070_ ;
	wire _w21071_ ;
	wire _w21072_ ;
	wire _w21073_ ;
	wire _w21074_ ;
	wire _w21075_ ;
	wire _w21076_ ;
	wire _w21077_ ;
	wire _w21078_ ;
	wire _w21079_ ;
	wire _w21080_ ;
	wire _w21081_ ;
	wire _w21082_ ;
	wire _w21083_ ;
	wire _w21084_ ;
	wire _w21085_ ;
	wire _w21086_ ;
	wire _w21087_ ;
	wire _w21088_ ;
	wire _w21089_ ;
	wire _w21090_ ;
	wire _w21091_ ;
	wire _w21092_ ;
	wire _w21093_ ;
	wire _w21094_ ;
	wire _w21095_ ;
	wire _w21096_ ;
	wire _w21097_ ;
	wire _w21098_ ;
	wire _w21099_ ;
	wire _w21100_ ;
	wire _w21101_ ;
	wire _w21102_ ;
	wire _w21103_ ;
	wire _w21104_ ;
	wire _w21105_ ;
	wire _w21106_ ;
	wire _w21107_ ;
	wire _w21108_ ;
	wire _w21109_ ;
	wire _w21110_ ;
	wire _w21111_ ;
	wire _w21112_ ;
	wire _w21113_ ;
	wire _w21114_ ;
	wire _w21115_ ;
	wire _w21116_ ;
	wire _w21117_ ;
	wire _w21118_ ;
	wire _w21119_ ;
	wire _w21120_ ;
	wire _w21121_ ;
	wire _w21122_ ;
	wire _w21123_ ;
	wire _w21124_ ;
	wire _w21125_ ;
	wire _w21126_ ;
	wire _w21127_ ;
	wire _w21128_ ;
	wire _w21129_ ;
	wire _w21130_ ;
	wire _w21131_ ;
	wire _w21132_ ;
	wire _w21133_ ;
	wire _w21134_ ;
	wire _w21135_ ;
	wire _w21136_ ;
	wire _w21137_ ;
	wire _w21138_ ;
	wire _w21139_ ;
	wire _w21140_ ;
	wire _w21141_ ;
	wire _w21142_ ;
	wire _w21143_ ;
	wire _w21144_ ;
	wire _w21145_ ;
	wire _w21146_ ;
	wire _w21147_ ;
	wire _w21148_ ;
	wire _w21149_ ;
	wire _w21150_ ;
	wire _w21151_ ;
	wire _w21152_ ;
	wire _w21153_ ;
	wire _w21154_ ;
	wire _w21155_ ;
	wire _w21156_ ;
	wire _w21157_ ;
	wire _w21158_ ;
	wire _w21159_ ;
	wire _w21160_ ;
	wire _w21161_ ;
	wire _w21162_ ;
	wire _w21163_ ;
	wire _w21164_ ;
	wire _w21165_ ;
	wire _w21166_ ;
	wire _w21167_ ;
	wire _w21168_ ;
	wire _w21169_ ;
	wire _w21170_ ;
	wire _w21171_ ;
	wire _w21172_ ;
	wire _w21173_ ;
	wire _w21174_ ;
	wire _w21175_ ;
	wire _w21176_ ;
	wire _w21177_ ;
	wire _w21178_ ;
	wire _w21179_ ;
	wire _w21180_ ;
	wire _w21181_ ;
	wire _w21182_ ;
	wire _w21183_ ;
	wire _w21184_ ;
	wire _w21185_ ;
	wire _w21186_ ;
	wire _w21187_ ;
	wire _w21188_ ;
	wire _w21189_ ;
	wire _w21190_ ;
	wire _w21191_ ;
	wire _w21192_ ;
	wire _w21193_ ;
	wire _w21194_ ;
	wire _w21195_ ;
	wire _w21196_ ;
	wire _w21197_ ;
	wire _w21198_ ;
	wire _w21199_ ;
	wire _w21200_ ;
	wire _w21201_ ;
	wire _w21202_ ;
	wire _w21203_ ;
	wire _w21204_ ;
	wire _w21205_ ;
	wire _w21206_ ;
	wire _w21207_ ;
	wire _w21208_ ;
	wire _w21209_ ;
	wire _w21210_ ;
	wire _w21211_ ;
	wire _w21212_ ;
	wire _w21213_ ;
	wire _w21214_ ;
	wire _w21215_ ;
	wire _w21216_ ;
	wire _w21217_ ;
	wire _w21218_ ;
	wire _w21219_ ;
	wire _w21220_ ;
	wire _w21221_ ;
	wire _w21222_ ;
	wire _w21223_ ;
	wire _w21224_ ;
	wire _w21225_ ;
	wire _w21226_ ;
	wire _w21227_ ;
	wire _w21228_ ;
	wire _w21229_ ;
	wire _w21230_ ;
	wire _w21231_ ;
	wire _w21232_ ;
	wire _w21233_ ;
	wire _w21234_ ;
	wire _w21235_ ;
	wire _w21236_ ;
	wire _w21237_ ;
	wire _w21238_ ;
	wire _w21239_ ;
	wire _w21240_ ;
	wire _w21241_ ;
	wire _w21242_ ;
	wire _w21243_ ;
	wire _w21244_ ;
	wire _w21245_ ;
	wire _w21246_ ;
	wire _w21247_ ;
	wire _w21248_ ;
	wire _w21249_ ;
	wire _w21250_ ;
	wire _w21251_ ;
	wire _w21252_ ;
	wire _w21253_ ;
	wire _w21254_ ;
	wire _w21255_ ;
	wire _w21256_ ;
	wire _w21257_ ;
	wire _w21258_ ;
	wire _w21259_ ;
	wire _w21260_ ;
	wire _w21261_ ;
	wire _w21262_ ;
	wire _w21263_ ;
	wire _w21264_ ;
	wire _w21265_ ;
	wire _w21266_ ;
	wire _w21267_ ;
	wire _w21268_ ;
	wire _w21269_ ;
	wire _w21270_ ;
	wire _w21271_ ;
	wire _w21272_ ;
	wire _w21273_ ;
	wire _w21274_ ;
	wire _w21275_ ;
	wire _w21276_ ;
	wire _w21277_ ;
	wire _w21278_ ;
	wire _w21279_ ;
	wire _w21280_ ;
	wire _w21281_ ;
	wire _w21282_ ;
	wire _w21283_ ;
	wire _w21284_ ;
	wire _w21285_ ;
	wire _w21286_ ;
	wire _w21287_ ;
	wire _w21288_ ;
	wire _w21289_ ;
	wire _w21290_ ;
	wire _w21291_ ;
	wire _w21292_ ;
	wire _w21293_ ;
	wire _w21294_ ;
	wire _w21295_ ;
	wire _w21296_ ;
	wire _w21297_ ;
	wire _w21298_ ;
	wire _w21299_ ;
	wire _w21300_ ;
	wire _w21301_ ;
	wire _w21302_ ;
	wire _w21303_ ;
	wire _w21304_ ;
	wire _w21305_ ;
	wire _w21306_ ;
	wire _w21307_ ;
	wire _w21308_ ;
	wire _w21309_ ;
	wire _w21310_ ;
	wire _w21311_ ;
	wire _w21312_ ;
	wire _w21313_ ;
	wire _w21314_ ;
	wire _w21315_ ;
	wire _w21316_ ;
	wire _w21317_ ;
	wire _w21318_ ;
	wire _w21319_ ;
	wire _w21320_ ;
	wire _w21321_ ;
	wire _w21322_ ;
	wire _w21323_ ;
	wire _w21324_ ;
	wire _w21325_ ;
	wire _w21326_ ;
	wire _w21327_ ;
	wire _w21328_ ;
	wire _w21329_ ;
	wire _w21330_ ;
	wire _w21331_ ;
	wire _w21332_ ;
	wire _w21333_ ;
	wire _w21334_ ;
	wire _w21335_ ;
	wire _w21336_ ;
	wire _w21337_ ;
	wire _w21338_ ;
	wire _w21339_ ;
	wire _w21340_ ;
	wire _w21341_ ;
	wire _w21342_ ;
	wire _w21343_ ;
	wire _w21344_ ;
	wire _w21345_ ;
	wire _w21346_ ;
	wire _w21347_ ;
	wire _w21348_ ;
	wire _w21349_ ;
	wire _w21350_ ;
	wire _w21351_ ;
	wire _w21352_ ;
	wire _w21353_ ;
	wire _w21354_ ;
	wire _w21355_ ;
	wire _w21356_ ;
	wire _w21357_ ;
	wire _w21358_ ;
	wire _w21359_ ;
	wire _w21360_ ;
	wire _w21361_ ;
	wire _w21362_ ;
	wire _w21363_ ;
	wire _w21364_ ;
	wire _w21365_ ;
	wire _w21366_ ;
	wire _w21367_ ;
	wire _w21368_ ;
	wire _w21369_ ;
	wire _w21370_ ;
	wire _w21371_ ;
	wire _w21372_ ;
	wire _w21373_ ;
	wire _w21374_ ;
	wire _w21375_ ;
	wire _w21376_ ;
	wire _w21377_ ;
	wire _w21378_ ;
	wire _w21379_ ;
	wire _w21380_ ;
	wire _w21381_ ;
	wire _w21382_ ;
	wire _w21383_ ;
	wire _w21384_ ;
	wire _w21385_ ;
	wire _w21386_ ;
	wire _w21387_ ;
	wire _w21388_ ;
	wire _w21389_ ;
	wire _w21390_ ;
	wire _w21391_ ;
	wire _w21392_ ;
	wire _w21393_ ;
	wire _w21394_ ;
	wire _w21395_ ;
	wire _w21396_ ;
	wire _w21397_ ;
	wire _w21398_ ;
	wire _w21399_ ;
	wire _w21400_ ;
	wire _w21401_ ;
	wire _w21402_ ;
	wire _w21403_ ;
	wire _w21404_ ;
	wire _w21405_ ;
	wire _w21406_ ;
	wire _w21407_ ;
	wire _w21408_ ;
	wire _w21409_ ;
	wire _w21410_ ;
	wire _w21411_ ;
	wire _w21412_ ;
	wire _w21413_ ;
	wire _w21414_ ;
	wire _w21415_ ;
	wire _w21416_ ;
	wire _w21417_ ;
	wire _w21418_ ;
	wire _w21419_ ;
	wire _w21420_ ;
	wire _w21421_ ;
	wire _w21422_ ;
	wire _w21423_ ;
	wire _w21424_ ;
	wire _w21425_ ;
	wire _w21426_ ;
	wire _w21427_ ;
	wire _w21428_ ;
	wire _w21429_ ;
	wire _w21430_ ;
	wire _w21431_ ;
	wire _w21432_ ;
	wire _w21433_ ;
	wire _w21434_ ;
	wire _w21435_ ;
	wire _w21436_ ;
	wire _w21437_ ;
	wire _w21438_ ;
	wire _w21439_ ;
	wire _w21440_ ;
	wire _w21441_ ;
	wire _w21442_ ;
	wire _w21443_ ;
	wire _w21444_ ;
	wire _w21445_ ;
	wire _w21446_ ;
	wire _w21447_ ;
	wire _w21448_ ;
	wire _w21449_ ;
	wire _w21450_ ;
	wire _w21451_ ;
	wire _w21452_ ;
	wire _w21453_ ;
	wire _w21454_ ;
	wire _w21455_ ;
	wire _w21456_ ;
	wire _w21457_ ;
	wire _w21458_ ;
	wire _w21459_ ;
	wire _w21460_ ;
	wire _w21461_ ;
	wire _w21462_ ;
	wire _w21463_ ;
	wire _w21464_ ;
	wire _w21465_ ;
	wire _w21466_ ;
	wire _w21467_ ;
	wire _w21468_ ;
	wire _w21469_ ;
	wire _w21470_ ;
	wire _w21471_ ;
	wire _w21472_ ;
	wire _w21473_ ;
	wire _w21474_ ;
	wire _w21475_ ;
	wire _w21476_ ;
	wire _w21477_ ;
	wire _w21478_ ;
	wire _w21479_ ;
	wire _w21480_ ;
	wire _w21481_ ;
	wire _w21482_ ;
	wire _w21483_ ;
	wire _w21484_ ;
	wire _w21485_ ;
	wire _w21486_ ;
	wire _w21487_ ;
	wire _w21488_ ;
	wire _w21489_ ;
	wire _w21490_ ;
	wire _w21491_ ;
	wire _w21492_ ;
	wire _w21493_ ;
	wire _w21494_ ;
	wire _w21495_ ;
	wire _w21496_ ;
	wire _w21497_ ;
	wire _w21498_ ;
	wire _w21499_ ;
	wire _w21500_ ;
	wire _w21501_ ;
	wire _w21502_ ;
	wire _w21503_ ;
	wire _w21504_ ;
	wire _w21505_ ;
	wire _w21506_ ;
	wire _w21507_ ;
	wire _w21508_ ;
	wire _w21509_ ;
	wire _w21510_ ;
	wire _w21511_ ;
	wire _w21512_ ;
	wire _w21513_ ;
	wire _w21514_ ;
	wire _w21515_ ;
	wire _w21516_ ;
	wire _w21517_ ;
	wire _w21518_ ;
	wire _w21519_ ;
	wire _w21520_ ;
	wire _w21521_ ;
	wire _w21522_ ;
	wire _w21523_ ;
	wire _w21524_ ;
	wire _w21525_ ;
	wire _w21526_ ;
	wire _w21527_ ;
	wire _w21528_ ;
	wire _w21529_ ;
	wire _w21530_ ;
	wire _w21531_ ;
	wire _w21532_ ;
	wire _w21533_ ;
	wire _w21534_ ;
	wire _w21535_ ;
	wire _w21536_ ;
	wire _w21537_ ;
	wire _w21538_ ;
	wire _w21539_ ;
	wire _w21540_ ;
	wire _w21541_ ;
	wire _w21542_ ;
	wire _w21543_ ;
	wire _w21544_ ;
	wire _w21545_ ;
	wire _w21546_ ;
	wire _w21547_ ;
	wire _w21548_ ;
	wire _w21549_ ;
	wire _w21550_ ;
	wire _w21551_ ;
	wire _w21552_ ;
	wire _w21553_ ;
	wire _w21554_ ;
	wire _w21555_ ;
	wire _w21556_ ;
	wire _w21557_ ;
	wire _w21558_ ;
	wire _w21559_ ;
	wire _w21560_ ;
	wire _w21561_ ;
	wire _w21562_ ;
	wire _w21563_ ;
	wire _w21564_ ;
	wire _w21565_ ;
	wire _w21566_ ;
	wire _w21567_ ;
	wire _w21568_ ;
	wire _w21569_ ;
	wire _w21570_ ;
	wire _w21571_ ;
	wire _w21572_ ;
	wire _w21573_ ;
	wire _w21574_ ;
	wire _w21575_ ;
	wire _w21576_ ;
	wire _w21577_ ;
	wire _w21578_ ;
	wire _w21579_ ;
	wire _w21580_ ;
	wire _w21581_ ;
	wire _w21582_ ;
	wire _w21583_ ;
	wire _w21584_ ;
	wire _w21585_ ;
	wire _w21586_ ;
	wire _w21587_ ;
	wire _w21588_ ;
	wire _w21589_ ;
	wire _w21590_ ;
	wire _w21591_ ;
	wire _w21592_ ;
	wire _w21593_ ;
	wire _w21594_ ;
	wire _w21595_ ;
	wire _w21596_ ;
	wire _w21597_ ;
	wire _w21598_ ;
	wire _w21599_ ;
	wire _w21600_ ;
	wire _w21601_ ;
	wire _w21602_ ;
	wire _w21603_ ;
	wire _w21604_ ;
	wire _w21605_ ;
	wire _w21606_ ;
	wire _w21607_ ;
	wire _w21608_ ;
	wire _w21609_ ;
	wire _w21610_ ;
	wire _w21611_ ;
	wire _w21612_ ;
	wire _w21613_ ;
	wire _w21614_ ;
	wire _w21615_ ;
	wire _w21616_ ;
	wire _w21617_ ;
	wire _w21618_ ;
	wire _w21619_ ;
	wire _w21620_ ;
	wire _w21621_ ;
	wire _w21622_ ;
	wire _w21623_ ;
	wire _w21624_ ;
	wire _w21625_ ;
	wire _w21626_ ;
	wire _w21627_ ;
	wire _w21628_ ;
	wire _w21629_ ;
	wire _w21630_ ;
	wire _w21631_ ;
	wire _w21632_ ;
	wire _w21633_ ;
	wire _w21634_ ;
	wire _w21635_ ;
	wire _w21636_ ;
	wire _w21637_ ;
	wire _w21638_ ;
	wire _w21639_ ;
	wire _w21640_ ;
	wire _w21641_ ;
	wire _w21642_ ;
	wire _w21643_ ;
	wire _w21644_ ;
	wire _w21645_ ;
	wire _w21646_ ;
	wire _w21647_ ;
	wire _w21648_ ;
	wire _w21649_ ;
	wire _w21650_ ;
	wire _w21651_ ;
	wire _w21652_ ;
	wire _w21653_ ;
	wire _w21654_ ;
	wire _w21655_ ;
	wire _w21656_ ;
	wire _w21657_ ;
	wire _w21658_ ;
	wire _w21659_ ;
	wire _w21660_ ;
	wire _w21661_ ;
	wire _w21662_ ;
	wire _w21663_ ;
	wire _w21664_ ;
	wire _w21665_ ;
	wire _w21666_ ;
	wire _w21667_ ;
	wire _w21668_ ;
	wire _w21669_ ;
	wire _w21670_ ;
	wire _w21671_ ;
	wire _w21672_ ;
	wire _w21673_ ;
	wire _w21674_ ;
	wire _w21675_ ;
	wire _w21676_ ;
	wire _w21677_ ;
	wire _w21678_ ;
	wire _w21679_ ;
	wire _w21680_ ;
	wire _w21681_ ;
	wire _w21682_ ;
	wire _w21683_ ;
	wire _w21684_ ;
	wire _w21685_ ;
	wire _w21686_ ;
	wire _w21687_ ;
	wire _w21688_ ;
	wire _w21689_ ;
	wire _w21690_ ;
	wire _w21691_ ;
	wire _w21692_ ;
	wire _w21693_ ;
	wire _w21694_ ;
	wire _w21695_ ;
	wire _w21696_ ;
	wire _w21697_ ;
	wire _w21698_ ;
	wire _w21699_ ;
	wire _w21700_ ;
	wire _w21701_ ;
	wire _w21702_ ;
	wire _w21703_ ;
	wire _w21704_ ;
	wire _w21705_ ;
	wire _w21706_ ;
	wire _w21707_ ;
	wire _w21708_ ;
	wire _w21709_ ;
	wire _w21710_ ;
	wire _w21711_ ;
	wire _w21712_ ;
	wire _w21713_ ;
	wire _w21714_ ;
	wire _w21715_ ;
	wire _w21716_ ;
	wire _w21717_ ;
	wire _w21718_ ;
	wire _w21719_ ;
	wire _w21720_ ;
	wire _w21721_ ;
	wire _w21722_ ;
	wire _w21723_ ;
	wire _w21724_ ;
	wire _w21725_ ;
	wire _w21726_ ;
	wire _w21727_ ;
	wire _w21728_ ;
	wire _w21729_ ;
	wire _w21730_ ;
	wire _w21731_ ;
	wire _w21732_ ;
	wire _w21733_ ;
	wire _w21734_ ;
	wire _w21735_ ;
	wire _w21736_ ;
	wire _w21737_ ;
	wire _w21738_ ;
	wire _w21739_ ;
	wire _w21740_ ;
	wire _w21741_ ;
	wire _w21742_ ;
	wire _w21743_ ;
	wire _w21744_ ;
	wire _w21745_ ;
	wire _w21746_ ;
	wire _w21747_ ;
	wire _w21748_ ;
	wire _w21749_ ;
	wire _w21750_ ;
	wire _w21751_ ;
	wire _w21752_ ;
	wire _w21753_ ;
	wire _w21754_ ;
	wire _w21755_ ;
	wire _w21756_ ;
	wire _w21757_ ;
	wire _w21758_ ;
	wire _w21759_ ;
	wire _w21760_ ;
	wire _w21761_ ;
	wire _w21762_ ;
	wire _w21763_ ;
	wire _w21764_ ;
	wire _w21765_ ;
	wire _w21766_ ;
	wire _w21767_ ;
	wire _w21768_ ;
	wire _w21769_ ;
	wire _w21770_ ;
	wire _w21771_ ;
	wire _w21772_ ;
	wire _w21773_ ;
	wire _w21774_ ;
	wire _w21775_ ;
	wire _w21776_ ;
	wire _w21777_ ;
	wire _w21778_ ;
	wire _w21779_ ;
	wire _w21780_ ;
	wire _w21781_ ;
	wire _w21782_ ;
	wire _w21783_ ;
	wire _w21784_ ;
	wire _w21785_ ;
	wire _w21786_ ;
	wire _w21787_ ;
	wire _w21788_ ;
	wire _w21789_ ;
	wire _w21790_ ;
	wire _w21791_ ;
	wire _w21792_ ;
	wire _w21793_ ;
	wire _w21794_ ;
	wire _w21795_ ;
	wire _w21796_ ;
	wire _w21797_ ;
	wire _w21798_ ;
	wire _w21799_ ;
	wire _w21800_ ;
	wire _w21801_ ;
	wire _w21802_ ;
	wire _w21803_ ;
	wire _w21804_ ;
	wire _w21805_ ;
	wire _w21806_ ;
	wire _w21807_ ;
	wire _w21808_ ;
	wire _w21809_ ;
	wire _w21810_ ;
	wire _w21811_ ;
	wire _w21812_ ;
	wire _w21813_ ;
	wire _w21814_ ;
	wire _w21815_ ;
	wire _w21816_ ;
	wire _w21817_ ;
	wire _w21818_ ;
	wire _w21819_ ;
	wire _w21820_ ;
	wire _w21821_ ;
	wire _w21822_ ;
	wire _w21823_ ;
	wire _w21824_ ;
	wire _w21825_ ;
	wire _w21826_ ;
	wire _w21827_ ;
	wire _w21828_ ;
	wire _w21829_ ;
	wire _w21830_ ;
	wire _w21831_ ;
	wire _w21832_ ;
	wire _w21833_ ;
	wire _w21834_ ;
	wire _w21835_ ;
	wire _w21836_ ;
	wire _w21837_ ;
	wire _w21838_ ;
	wire _w21839_ ;
	wire _w21840_ ;
	wire _w21841_ ;
	wire _w21842_ ;
	wire _w21843_ ;
	wire _w21844_ ;
	wire _w21845_ ;
	wire _w21846_ ;
	wire _w21847_ ;
	wire _w21848_ ;
	wire _w21849_ ;
	wire _w21850_ ;
	wire _w21851_ ;
	wire _w21852_ ;
	wire _w21853_ ;
	wire _w21854_ ;
	wire _w21855_ ;
	wire _w21856_ ;
	wire _w21857_ ;
	wire _w21858_ ;
	wire _w21859_ ;
	wire _w21860_ ;
	wire _w21861_ ;
	wire _w21862_ ;
	wire _w21863_ ;
	wire _w21864_ ;
	wire _w21865_ ;
	wire _w21866_ ;
	wire _w21867_ ;
	wire _w21868_ ;
	wire _w21869_ ;
	wire _w21870_ ;
	wire _w21871_ ;
	wire _w21872_ ;
	wire _w21873_ ;
	wire _w21874_ ;
	wire _w21875_ ;
	wire _w21876_ ;
	wire _w21877_ ;
	wire _w21878_ ;
	wire _w21879_ ;
	wire _w21880_ ;
	wire _w21881_ ;
	wire _w21882_ ;
	wire _w21883_ ;
	wire _w21884_ ;
	wire _w21885_ ;
	wire _w21886_ ;
	wire _w21887_ ;
	wire _w21888_ ;
	wire _w21889_ ;
	wire _w21890_ ;
	wire _w21891_ ;
	wire _w21892_ ;
	wire _w21893_ ;
	wire _w21894_ ;
	wire _w21895_ ;
	wire _w21896_ ;
	wire _w21897_ ;
	wire _w21898_ ;
	wire _w21899_ ;
	wire _w21900_ ;
	wire _w21901_ ;
	wire _w21902_ ;
	wire _w21903_ ;
	wire _w21904_ ;
	wire _w21905_ ;
	wire _w21906_ ;
	wire _w21907_ ;
	wire _w21908_ ;
	wire _w21909_ ;
	wire _w21910_ ;
	wire _w21911_ ;
	wire _w21912_ ;
	wire _w21913_ ;
	wire _w21914_ ;
	wire _w21915_ ;
	wire _w21916_ ;
	wire _w21917_ ;
	wire _w21918_ ;
	wire _w21919_ ;
	wire _w21920_ ;
	wire _w21921_ ;
	wire _w21922_ ;
	wire _w21923_ ;
	wire _w21924_ ;
	wire _w21925_ ;
	wire _w21926_ ;
	wire _w21927_ ;
	wire _w21928_ ;
	wire _w21929_ ;
	wire _w21930_ ;
	wire _w21931_ ;
	wire _w21932_ ;
	wire _w21933_ ;
	wire _w21934_ ;
	wire _w21935_ ;
	wire _w21936_ ;
	wire _w21937_ ;
	wire _w21938_ ;
	wire _w21939_ ;
	wire _w21940_ ;
	wire _w21941_ ;
	wire _w21942_ ;
	wire _w21943_ ;
	wire _w21944_ ;
	wire _w21945_ ;
	wire _w21946_ ;
	wire _w21947_ ;
	wire _w21948_ ;
	wire _w21949_ ;
	wire _w21950_ ;
	wire _w21951_ ;
	wire _w21952_ ;
	wire _w21953_ ;
	wire _w21954_ ;
	wire _w21955_ ;
	wire _w21956_ ;
	wire _w21957_ ;
	wire _w21958_ ;
	wire _w21959_ ;
	wire _w21960_ ;
	wire _w21961_ ;
	wire _w21962_ ;
	wire _w21963_ ;
	wire _w21964_ ;
	wire _w21965_ ;
	wire _w21966_ ;
	wire _w21967_ ;
	wire _w21968_ ;
	wire _w21969_ ;
	wire _w21970_ ;
	wire _w21971_ ;
	wire _w21972_ ;
	wire _w21973_ ;
	wire _w21974_ ;
	wire _w21975_ ;
	wire _w21976_ ;
	wire _w21977_ ;
	wire _w21978_ ;
	wire _w21979_ ;
	wire _w21980_ ;
	wire _w21981_ ;
	wire _w21982_ ;
	wire _w21983_ ;
	wire _w21984_ ;
	wire _w21985_ ;
	wire _w21986_ ;
	wire _w21987_ ;
	wire _w21988_ ;
	wire _w21989_ ;
	wire _w21990_ ;
	wire _w21991_ ;
	wire _w21992_ ;
	wire _w21993_ ;
	wire _w21994_ ;
	wire _w21995_ ;
	wire _w21996_ ;
	wire _w21997_ ;
	wire _w21998_ ;
	wire _w21999_ ;
	wire _w22000_ ;
	wire _w22001_ ;
	wire _w22002_ ;
	wire _w22003_ ;
	wire _w22004_ ;
	wire _w22005_ ;
	wire _w22006_ ;
	wire _w22007_ ;
	wire _w22008_ ;
	wire _w22009_ ;
	wire _w22010_ ;
	wire _w22011_ ;
	wire _w22012_ ;
	wire _w22013_ ;
	wire _w22014_ ;
	wire _w22015_ ;
	wire _w22016_ ;
	wire _w22017_ ;
	wire _w22018_ ;
	wire _w22019_ ;
	wire _w22020_ ;
	wire _w22021_ ;
	wire _w22022_ ;
	wire _w22023_ ;
	wire _w22024_ ;
	wire _w22025_ ;
	wire _w22026_ ;
	wire _w22027_ ;
	wire _w22028_ ;
	wire _w22029_ ;
	wire _w22030_ ;
	wire _w22031_ ;
	wire _w22032_ ;
	wire _w22033_ ;
	wire _w22034_ ;
	wire _w22035_ ;
	wire _w22036_ ;
	wire _w22037_ ;
	wire _w22038_ ;
	wire _w22039_ ;
	wire _w22040_ ;
	wire _w22041_ ;
	wire _w22042_ ;
	wire _w22043_ ;
	wire _w22044_ ;
	wire _w22045_ ;
	wire _w22046_ ;
	wire _w22047_ ;
	wire _w22048_ ;
	wire _w22049_ ;
	wire _w22050_ ;
	wire _w22051_ ;
	wire _w22052_ ;
	wire _w22053_ ;
	wire _w22054_ ;
	wire _w22055_ ;
	wire _w22056_ ;
	wire _w22057_ ;
	wire _w22058_ ;
	wire _w22059_ ;
	wire _w22060_ ;
	wire _w22061_ ;
	wire _w22062_ ;
	wire _w22063_ ;
	wire _w22064_ ;
	wire _w22065_ ;
	wire _w22066_ ;
	wire _w22067_ ;
	wire _w22068_ ;
	wire _w22069_ ;
	wire _w22070_ ;
	wire _w22071_ ;
	wire _w22072_ ;
	wire _w22073_ ;
	wire _w22074_ ;
	wire _w22075_ ;
	wire _w22076_ ;
	wire _w22077_ ;
	wire _w22078_ ;
	wire _w22079_ ;
	wire _w22080_ ;
	wire _w22081_ ;
	wire _w22082_ ;
	wire _w22083_ ;
	wire _w22084_ ;
	wire _w22085_ ;
	wire _w22086_ ;
	wire _w22087_ ;
	wire _w22088_ ;
	wire _w22089_ ;
	wire _w22090_ ;
	wire _w22091_ ;
	wire _w22092_ ;
	wire _w22093_ ;
	wire _w22094_ ;
	wire _w22095_ ;
	wire _w22096_ ;
	wire _w22097_ ;
	wire _w22098_ ;
	wire _w22099_ ;
	wire _w22100_ ;
	wire _w22101_ ;
	wire _w22102_ ;
	wire _w22103_ ;
	wire _w22104_ ;
	wire _w22105_ ;
	wire _w22106_ ;
	wire _w22107_ ;
	wire _w22108_ ;
	wire _w22109_ ;
	wire _w22110_ ;
	wire _w22111_ ;
	wire _w22112_ ;
	wire _w22113_ ;
	wire _w22114_ ;
	wire _w22115_ ;
	wire _w22116_ ;
	wire _w22117_ ;
	wire _w22118_ ;
	wire _w22119_ ;
	wire _w22120_ ;
	wire _w22121_ ;
	wire _w22122_ ;
	wire _w22123_ ;
	wire _w22124_ ;
	wire _w22125_ ;
	wire _w22126_ ;
	wire _w22127_ ;
	wire _w22128_ ;
	wire _w22129_ ;
	wire _w22130_ ;
	wire _w22131_ ;
	wire _w22132_ ;
	wire _w22133_ ;
	wire _w22134_ ;
	wire _w22135_ ;
	wire _w22136_ ;
	wire _w22137_ ;
	wire _w22138_ ;
	wire _w22139_ ;
	wire _w22140_ ;
	wire _w22141_ ;
	wire _w22142_ ;
	wire _w22143_ ;
	wire _w22144_ ;
	wire _w22145_ ;
	wire _w22146_ ;
	wire _w22147_ ;
	wire _w22148_ ;
	wire _w22149_ ;
	wire _w22150_ ;
	wire _w22151_ ;
	wire _w22152_ ;
	wire _w22153_ ;
	wire _w22154_ ;
	wire _w22155_ ;
	wire _w22156_ ;
	wire _w22157_ ;
	wire _w22158_ ;
	wire _w22159_ ;
	wire _w22160_ ;
	wire _w22161_ ;
	wire _w22162_ ;
	wire _w22163_ ;
	wire _w22164_ ;
	wire _w22165_ ;
	wire _w22166_ ;
	wire _w22167_ ;
	wire _w22168_ ;
	wire _w22169_ ;
	wire _w22170_ ;
	wire _w22171_ ;
	wire _w22172_ ;
	wire _w22173_ ;
	wire _w22174_ ;
	wire _w22175_ ;
	wire _w22176_ ;
	wire _w22177_ ;
	wire _w22178_ ;
	wire _w22179_ ;
	wire _w22180_ ;
	wire _w22181_ ;
	wire _w22182_ ;
	wire _w22183_ ;
	wire _w22184_ ;
	wire _w22185_ ;
	wire _w22186_ ;
	wire _w22187_ ;
	wire _w22188_ ;
	wire _w22189_ ;
	wire _w22190_ ;
	wire _w22191_ ;
	wire _w22192_ ;
	wire _w22193_ ;
	wire _w22194_ ;
	wire _w22195_ ;
	wire _w22196_ ;
	wire _w22197_ ;
	wire _w22198_ ;
	wire _w22199_ ;
	wire _w22200_ ;
	wire _w22201_ ;
	wire _w22202_ ;
	wire _w22203_ ;
	wire _w22204_ ;
	wire _w22205_ ;
	wire _w22206_ ;
	wire _w22207_ ;
	wire _w22208_ ;
	wire _w22209_ ;
	wire _w22210_ ;
	wire _w22211_ ;
	wire _w22212_ ;
	wire _w22213_ ;
	wire _w22214_ ;
	wire _w22215_ ;
	wire _w22216_ ;
	wire _w22217_ ;
	wire _w22218_ ;
	wire _w22219_ ;
	wire _w22220_ ;
	wire _w22221_ ;
	wire _w22222_ ;
	wire _w22223_ ;
	wire _w22224_ ;
	wire _w22225_ ;
	wire _w22226_ ;
	wire _w22227_ ;
	wire _w22228_ ;
	wire _w22229_ ;
	wire _w22230_ ;
	wire _w22231_ ;
	wire _w22232_ ;
	wire _w22233_ ;
	wire _w22234_ ;
	wire _w22235_ ;
	wire _w22236_ ;
	wire _w22237_ ;
	wire _w22238_ ;
	wire _w22239_ ;
	wire _w22240_ ;
	wire _w22241_ ;
	wire _w22242_ ;
	wire _w22243_ ;
	wire _w22244_ ;
	wire _w22245_ ;
	wire _w22246_ ;
	wire _w22247_ ;
	wire _w22248_ ;
	wire _w22249_ ;
	wire _w22250_ ;
	wire _w22251_ ;
	wire _w22252_ ;
	wire _w22253_ ;
	wire _w22254_ ;
	wire _w22255_ ;
	wire _w22256_ ;
	wire _w22257_ ;
	wire _w22258_ ;
	wire _w22259_ ;
	wire _w22260_ ;
	wire _w22261_ ;
	wire _w22262_ ;
	wire _w22263_ ;
	wire _w22264_ ;
	wire _w22265_ ;
	wire _w22266_ ;
	wire _w22267_ ;
	wire _w22268_ ;
	wire _w22269_ ;
	wire _w22270_ ;
	wire _w22271_ ;
	wire _w22272_ ;
	wire _w22273_ ;
	wire _w22274_ ;
	wire _w22275_ ;
	wire _w22276_ ;
	wire _w22277_ ;
	wire _w22278_ ;
	wire _w22279_ ;
	wire _w22280_ ;
	wire _w22281_ ;
	wire _w22282_ ;
	wire _w22283_ ;
	wire _w22284_ ;
	wire _w22285_ ;
	wire _w22286_ ;
	wire _w22287_ ;
	wire _w22288_ ;
	wire _w22289_ ;
	wire _w22290_ ;
	wire _w22291_ ;
	wire _w22292_ ;
	wire _w22293_ ;
	wire _w22294_ ;
	wire _w22295_ ;
	wire _w22296_ ;
	wire _w22297_ ;
	wire _w22298_ ;
	wire _w22299_ ;
	wire _w22300_ ;
	wire _w22301_ ;
	wire _w22302_ ;
	wire _w22303_ ;
	wire _w22304_ ;
	wire _w22305_ ;
	wire _w22306_ ;
	wire _w22307_ ;
	wire _w22308_ ;
	wire _w22309_ ;
	wire _w22310_ ;
	wire _w22311_ ;
	wire _w22312_ ;
	wire _w22313_ ;
	wire _w22314_ ;
	wire _w22315_ ;
	wire _w22316_ ;
	wire _w22317_ ;
	wire _w22318_ ;
	wire _w22319_ ;
	wire _w22320_ ;
	wire _w22321_ ;
	wire _w22322_ ;
	wire _w22323_ ;
	wire _w22324_ ;
	wire _w22325_ ;
	wire _w22326_ ;
	wire _w22327_ ;
	wire _w22328_ ;
	wire _w22329_ ;
	wire _w22330_ ;
	wire _w22331_ ;
	wire _w22332_ ;
	wire _w22333_ ;
	wire _w22334_ ;
	wire _w22335_ ;
	wire _w22336_ ;
	wire _w22337_ ;
	wire _w22338_ ;
	wire _w22339_ ;
	wire _w22340_ ;
	wire _w22341_ ;
	wire _w22342_ ;
	wire _w22343_ ;
	wire _w22344_ ;
	wire _w22345_ ;
	wire _w22346_ ;
	wire _w22347_ ;
	wire _w22348_ ;
	wire _w22349_ ;
	wire _w22350_ ;
	wire _w22351_ ;
	wire _w22352_ ;
	wire _w22353_ ;
	wire _w22354_ ;
	wire _w22355_ ;
	wire _w22356_ ;
	wire _w22357_ ;
	wire _w22358_ ;
	wire _w22359_ ;
	wire _w22360_ ;
	wire _w22361_ ;
	wire _w22362_ ;
	wire _w22363_ ;
	wire _w22364_ ;
	wire _w22365_ ;
	wire _w22366_ ;
	wire _w22367_ ;
	wire _w22368_ ;
	wire _w22369_ ;
	wire _w22370_ ;
	wire _w22371_ ;
	wire _w22372_ ;
	wire _w22373_ ;
	wire _w22374_ ;
	wire _w22375_ ;
	wire _w22376_ ;
	wire _w22377_ ;
	wire _w22378_ ;
	wire _w22379_ ;
	wire _w22380_ ;
	wire _w22381_ ;
	wire _w22382_ ;
	wire _w22383_ ;
	wire _w22384_ ;
	wire _w22385_ ;
	wire _w22386_ ;
	wire _w22387_ ;
	wire _w22388_ ;
	wire _w22389_ ;
	wire _w22390_ ;
	wire _w22391_ ;
	wire _w22392_ ;
	wire _w22393_ ;
	wire _w22394_ ;
	wire _w22395_ ;
	wire _w22396_ ;
	wire _w22397_ ;
	wire _w22398_ ;
	wire _w22399_ ;
	wire _w22400_ ;
	wire _w22401_ ;
	wire _w22402_ ;
	wire _w22403_ ;
	wire _w22404_ ;
	wire _w22405_ ;
	wire _w22406_ ;
	wire _w22407_ ;
	wire _w22408_ ;
	wire _w22409_ ;
	wire _w22410_ ;
	wire _w22411_ ;
	wire _w22412_ ;
	wire _w22413_ ;
	wire _w22414_ ;
	wire _w22415_ ;
	wire _w22416_ ;
	wire _w22417_ ;
	wire _w22418_ ;
	wire _w22419_ ;
	wire _w22420_ ;
	wire _w22421_ ;
	wire _w22422_ ;
	wire _w22423_ ;
	wire _w22424_ ;
	wire _w22425_ ;
	wire _w22426_ ;
	wire _w22427_ ;
	wire _w22428_ ;
	wire _w22429_ ;
	wire _w22430_ ;
	wire _w22431_ ;
	wire _w22432_ ;
	wire _w22433_ ;
	wire _w22434_ ;
	wire _w22435_ ;
	wire _w22436_ ;
	wire _w22437_ ;
	wire _w22438_ ;
	wire _w22439_ ;
	wire _w22440_ ;
	wire _w22441_ ;
	wire _w22442_ ;
	wire _w22443_ ;
	wire _w22444_ ;
	wire _w22445_ ;
	wire _w22446_ ;
	wire _w22447_ ;
	wire _w22448_ ;
	wire _w22449_ ;
	wire _w22450_ ;
	wire _w22451_ ;
	wire _w22452_ ;
	wire _w22453_ ;
	wire _w22454_ ;
	wire _w22455_ ;
	wire _w22456_ ;
	wire _w22457_ ;
	wire _w22458_ ;
	wire _w22459_ ;
	wire _w22460_ ;
	wire _w22461_ ;
	wire _w22462_ ;
	wire _w22463_ ;
	wire _w22464_ ;
	wire _w22465_ ;
	wire _w22466_ ;
	wire _w22467_ ;
	wire _w22468_ ;
	wire _w22469_ ;
	wire _w22470_ ;
	wire _w22471_ ;
	wire _w22472_ ;
	wire _w22473_ ;
	wire _w22474_ ;
	wire _w22475_ ;
	wire _w22476_ ;
	wire _w22477_ ;
	wire _w22478_ ;
	wire _w22479_ ;
	wire _w22480_ ;
	wire _w22481_ ;
	wire _w22482_ ;
	wire _w22483_ ;
	wire _w22484_ ;
	wire _w22485_ ;
	wire _w22486_ ;
	wire _w22487_ ;
	wire _w22488_ ;
	wire _w22489_ ;
	wire _w22490_ ;
	wire _w22491_ ;
	wire _w22492_ ;
	wire _w22493_ ;
	wire _w22494_ ;
	wire _w22495_ ;
	wire _w22496_ ;
	wire _w22497_ ;
	wire _w22498_ ;
	wire _w22499_ ;
	wire _w22500_ ;
	wire _w22501_ ;
	wire _w22502_ ;
	wire _w22503_ ;
	wire _w22504_ ;
	wire _w22505_ ;
	wire _w22506_ ;
	wire _w22507_ ;
	wire _w22508_ ;
	wire _w22509_ ;
	wire _w22510_ ;
	wire _w22511_ ;
	wire _w22512_ ;
	wire _w22513_ ;
	wire _w22514_ ;
	wire _w22515_ ;
	wire _w22516_ ;
	wire _w22517_ ;
	wire _w22518_ ;
	wire _w22519_ ;
	wire _w22520_ ;
	wire _w22521_ ;
	wire _w22522_ ;
	wire _w22523_ ;
	wire _w22524_ ;
	wire _w22525_ ;
	wire _w22526_ ;
	wire _w22527_ ;
	wire _w22528_ ;
	wire _w22529_ ;
	wire _w22530_ ;
	wire _w22531_ ;
	wire _w22532_ ;
	wire _w22533_ ;
	wire _w22534_ ;
	wire _w22535_ ;
	wire _w22536_ ;
	wire _w22537_ ;
	wire _w22538_ ;
	wire _w22539_ ;
	wire _w22540_ ;
	wire _w22541_ ;
	wire _w22542_ ;
	wire _w22543_ ;
	wire _w22544_ ;
	wire _w22545_ ;
	wire _w22546_ ;
	wire _w22547_ ;
	wire _w22548_ ;
	wire _w22549_ ;
	wire _w22550_ ;
	wire _w22551_ ;
	wire _w22552_ ;
	wire _w22553_ ;
	wire _w22554_ ;
	wire _w22555_ ;
	wire _w22556_ ;
	wire _w22557_ ;
	wire _w22558_ ;
	wire _w22559_ ;
	wire _w22560_ ;
	wire _w22561_ ;
	wire _w22562_ ;
	wire _w22563_ ;
	wire _w22564_ ;
	wire _w22565_ ;
	wire _w22566_ ;
	wire _w22567_ ;
	wire _w22568_ ;
	wire _w22569_ ;
	wire _w22570_ ;
	wire _w22571_ ;
	wire _w22572_ ;
	wire _w22573_ ;
	wire _w22574_ ;
	wire _w22575_ ;
	wire _w22576_ ;
	wire _w22577_ ;
	wire _w22578_ ;
	wire _w22579_ ;
	wire _w22580_ ;
	wire _w22581_ ;
	wire _w22582_ ;
	wire _w22583_ ;
	wire _w22584_ ;
	wire _w22585_ ;
	wire _w22586_ ;
	wire _w22587_ ;
	wire _w22588_ ;
	wire _w22589_ ;
	wire _w22590_ ;
	wire _w22591_ ;
	wire _w22592_ ;
	wire _w22593_ ;
	wire _w22594_ ;
	wire _w22595_ ;
	wire _w22596_ ;
	wire _w22597_ ;
	wire _w22598_ ;
	wire _w22599_ ;
	wire _w22600_ ;
	wire _w22601_ ;
	wire _w22602_ ;
	wire _w22603_ ;
	wire _w22604_ ;
	wire _w22605_ ;
	wire _w22606_ ;
	wire _w22607_ ;
	wire _w22608_ ;
	wire _w22609_ ;
	wire _w22610_ ;
	wire _w22611_ ;
	wire _w22612_ ;
	wire _w22613_ ;
	wire _w22614_ ;
	wire _w22615_ ;
	wire _w22616_ ;
	wire _w22617_ ;
	wire _w22618_ ;
	wire _w22619_ ;
	wire _w22620_ ;
	wire _w22621_ ;
	wire _w22622_ ;
	wire _w22623_ ;
	wire _w22624_ ;
	wire _w22625_ ;
	wire _w22626_ ;
	wire _w22627_ ;
	wire _w22628_ ;
	wire _w22629_ ;
	wire _w22630_ ;
	wire _w22631_ ;
	wire _w22632_ ;
	wire _w22633_ ;
	wire _w22634_ ;
	wire _w22635_ ;
	wire _w22636_ ;
	wire _w22637_ ;
	wire _w22638_ ;
	wire _w22639_ ;
	wire _w22640_ ;
	wire _w22641_ ;
	wire _w22642_ ;
	wire _w22643_ ;
	wire _w22644_ ;
	wire _w22645_ ;
	wire _w22646_ ;
	wire _w22647_ ;
	wire _w22648_ ;
	wire _w22649_ ;
	wire _w22650_ ;
	wire _w22651_ ;
	wire _w22652_ ;
	wire _w22653_ ;
	wire _w22654_ ;
	wire _w22655_ ;
	wire _w22656_ ;
	wire _w22657_ ;
	wire _w22658_ ;
	wire _w22659_ ;
	wire _w22660_ ;
	wire _w22661_ ;
	wire _w22662_ ;
	wire _w22663_ ;
	wire _w22664_ ;
	wire _w22665_ ;
	wire _w22666_ ;
	wire _w22667_ ;
	wire _w22668_ ;
	wire _w22669_ ;
	wire _w22670_ ;
	wire _w22671_ ;
	wire _w22672_ ;
	wire _w22673_ ;
	wire _w22674_ ;
	wire _w22675_ ;
	wire _w22676_ ;
	wire _w22677_ ;
	wire _w22678_ ;
	wire _w22679_ ;
	wire _w22680_ ;
	wire _w22681_ ;
	wire _w22682_ ;
	wire _w22683_ ;
	wire _w22684_ ;
	wire _w22685_ ;
	wire _w22686_ ;
	wire _w22687_ ;
	wire _w22688_ ;
	wire _w22689_ ;
	wire _w22690_ ;
	wire _w22691_ ;
	wire _w22692_ ;
	wire _w22693_ ;
	wire _w22694_ ;
	wire _w22695_ ;
	wire _w22696_ ;
	wire _w22697_ ;
	wire _w22698_ ;
	wire _w22699_ ;
	wire _w22700_ ;
	wire _w22701_ ;
	wire _w22702_ ;
	wire _w22703_ ;
	wire _w22704_ ;
	wire _w22705_ ;
	wire _w22706_ ;
	wire _w22707_ ;
	wire _w22708_ ;
	wire _w22709_ ;
	wire _w22710_ ;
	wire _w22711_ ;
	wire _w22712_ ;
	wire _w22713_ ;
	wire _w22714_ ;
	wire _w22715_ ;
	wire _w22716_ ;
	wire _w22717_ ;
	wire _w22718_ ;
	wire _w22719_ ;
	wire _w22720_ ;
	wire _w22721_ ;
	wire _w22722_ ;
	wire _w22723_ ;
	wire _w22724_ ;
	wire _w22725_ ;
	wire _w22726_ ;
	wire _w22727_ ;
	wire _w22728_ ;
	wire _w22729_ ;
	wire _w22730_ ;
	wire _w22731_ ;
	wire _w22732_ ;
	wire _w22733_ ;
	wire _w22734_ ;
	wire _w22735_ ;
	wire _w22736_ ;
	wire _w22737_ ;
	wire _w22738_ ;
	wire _w22739_ ;
	wire _w22740_ ;
	wire _w22741_ ;
	wire _w22742_ ;
	wire _w22743_ ;
	wire _w22744_ ;
	wire _w22745_ ;
	wire _w22746_ ;
	wire _w22747_ ;
	wire _w22748_ ;
	wire _w22749_ ;
	wire _w22750_ ;
	wire _w22751_ ;
	wire _w22752_ ;
	wire _w22753_ ;
	wire _w22754_ ;
	wire _w22755_ ;
	wire _w22756_ ;
	wire _w22757_ ;
	wire _w22758_ ;
	wire _w22759_ ;
	wire _w22760_ ;
	wire _w22761_ ;
	wire _w22762_ ;
	wire _w22763_ ;
	wire _w22764_ ;
	wire _w22765_ ;
	wire _w22766_ ;
	wire _w22767_ ;
	wire _w22768_ ;
	wire _w22769_ ;
	wire _w22770_ ;
	wire _w22771_ ;
	wire _w22772_ ;
	wire _w22773_ ;
	wire _w22774_ ;
	wire _w22775_ ;
	wire _w22776_ ;
	wire _w22777_ ;
	wire _w22778_ ;
	wire _w22779_ ;
	wire _w22780_ ;
	wire _w22781_ ;
	wire _w22782_ ;
	wire _w22783_ ;
	wire _w22784_ ;
	wire _w22785_ ;
	wire _w22786_ ;
	wire _w22787_ ;
	wire _w22788_ ;
	wire _w22789_ ;
	wire _w22790_ ;
	wire _w22791_ ;
	wire _w22792_ ;
	wire _w22793_ ;
	wire _w22794_ ;
	wire _w22795_ ;
	wire _w22796_ ;
	wire _w22797_ ;
	wire _w22798_ ;
	wire _w22799_ ;
	wire _w22800_ ;
	wire _w22801_ ;
	wire _w22802_ ;
	wire _w22803_ ;
	wire _w22804_ ;
	wire _w22805_ ;
	wire _w22806_ ;
	wire _w22807_ ;
	wire _w22808_ ;
	wire _w22809_ ;
	wire _w22810_ ;
	wire _w22811_ ;
	wire _w22812_ ;
	wire _w22813_ ;
	wire _w22814_ ;
	wire _w22815_ ;
	wire _w22816_ ;
	wire _w22817_ ;
	wire _w22818_ ;
	wire _w22819_ ;
	wire _w22820_ ;
	wire _w22821_ ;
	wire _w22822_ ;
	wire _w22823_ ;
	wire _w22824_ ;
	wire _w22825_ ;
	wire _w22826_ ;
	wire _w22827_ ;
	wire _w22828_ ;
	wire _w22829_ ;
	wire _w22830_ ;
	wire _w22831_ ;
	wire _w22832_ ;
	wire _w22833_ ;
	wire _w22834_ ;
	wire _w22835_ ;
	wire _w22836_ ;
	wire _w22837_ ;
	wire _w22838_ ;
	wire _w22839_ ;
	wire _w22840_ ;
	wire _w22841_ ;
	wire _w22842_ ;
	wire _w22843_ ;
	wire _w22844_ ;
	wire _w22845_ ;
	wire _w22846_ ;
	wire _w22847_ ;
	wire _w22848_ ;
	wire _w22849_ ;
	wire _w22850_ ;
	wire _w22851_ ;
	wire _w22852_ ;
	wire _w22853_ ;
	wire _w22854_ ;
	wire _w22855_ ;
	wire _w22856_ ;
	wire _w22857_ ;
	wire _w22858_ ;
	wire _w22859_ ;
	wire _w22860_ ;
	wire _w22861_ ;
	wire _w22862_ ;
	wire _w22863_ ;
	wire _w22864_ ;
	wire _w22865_ ;
	wire _w22866_ ;
	wire _w22867_ ;
	wire _w22868_ ;
	wire _w22869_ ;
	wire _w22870_ ;
	wire _w22871_ ;
	wire _w22872_ ;
	wire _w22873_ ;
	wire _w22874_ ;
	wire _w22875_ ;
	wire _w22876_ ;
	wire _w22877_ ;
	wire _w22878_ ;
	wire _w22879_ ;
	wire _w22880_ ;
	wire _w22881_ ;
	wire _w22882_ ;
	wire _w22883_ ;
	wire _w22884_ ;
	wire _w22885_ ;
	wire _w22886_ ;
	wire _w22887_ ;
	wire _w22888_ ;
	wire _w22889_ ;
	wire _w22890_ ;
	wire _w22891_ ;
	wire _w22892_ ;
	wire _w22893_ ;
	wire _w22894_ ;
	wire _w22895_ ;
	wire _w22896_ ;
	wire _w22897_ ;
	wire _w22898_ ;
	wire _w22899_ ;
	wire _w22900_ ;
	wire _w22901_ ;
	wire _w22902_ ;
	wire _w22903_ ;
	wire _w22904_ ;
	wire _w22905_ ;
	wire _w22906_ ;
	wire _w22907_ ;
	wire _w22908_ ;
	wire _w22909_ ;
	wire _w22910_ ;
	wire _w22911_ ;
	wire _w22912_ ;
	wire _w22913_ ;
	wire _w22914_ ;
	wire _w22915_ ;
	wire _w22916_ ;
	wire _w22917_ ;
	wire _w22918_ ;
	wire _w22919_ ;
	wire _w22920_ ;
	wire _w22921_ ;
	wire _w22922_ ;
	wire _w22923_ ;
	wire _w22924_ ;
	wire _w22925_ ;
	wire _w22926_ ;
	wire _w22927_ ;
	wire _w22928_ ;
	wire _w22929_ ;
	wire _w22930_ ;
	wire _w22931_ ;
	wire _w22932_ ;
	wire _w22933_ ;
	wire _w22934_ ;
	wire _w22935_ ;
	wire _w22936_ ;
	wire _w22937_ ;
	wire _w22938_ ;
	wire _w22939_ ;
	wire _w22940_ ;
	wire _w22941_ ;
	wire _w22942_ ;
	wire _w22943_ ;
	wire _w22944_ ;
	wire _w22945_ ;
	wire _w22946_ ;
	wire _w22947_ ;
	wire _w22948_ ;
	wire _w22949_ ;
	wire _w22950_ ;
	wire _w22951_ ;
	wire _w22952_ ;
	wire _w22953_ ;
	wire _w22954_ ;
	wire _w22955_ ;
	wire _w22956_ ;
	wire _w22957_ ;
	wire _w22958_ ;
	wire _w22959_ ;
	wire _w22960_ ;
	wire _w22961_ ;
	wire _w22962_ ;
	wire _w22963_ ;
	wire _w22964_ ;
	wire _w22965_ ;
	wire _w22966_ ;
	wire _w22967_ ;
	wire _w22968_ ;
	wire _w22969_ ;
	wire _w22970_ ;
	wire _w22971_ ;
	wire _w22972_ ;
	wire _w22973_ ;
	wire _w22974_ ;
	wire _w22975_ ;
	wire _w22976_ ;
	wire _w22977_ ;
	wire _w22978_ ;
	wire _w22979_ ;
	wire _w22980_ ;
	wire _w22981_ ;
	wire _w22982_ ;
	wire _w22983_ ;
	wire _w22984_ ;
	wire _w22985_ ;
	wire _w22986_ ;
	wire _w22987_ ;
	wire _w22988_ ;
	wire _w22989_ ;
	wire _w22990_ ;
	wire _w22991_ ;
	wire _w22992_ ;
	wire _w22993_ ;
	wire _w22994_ ;
	wire _w22995_ ;
	wire _w22996_ ;
	wire _w22997_ ;
	wire _w22998_ ;
	wire _w22999_ ;
	wire _w23000_ ;
	wire _w23001_ ;
	wire _w23002_ ;
	wire _w23003_ ;
	wire _w23004_ ;
	wire _w23005_ ;
	wire _w23006_ ;
	wire _w23007_ ;
	wire _w23008_ ;
	wire _w23009_ ;
	wire _w23010_ ;
	wire _w23011_ ;
	wire _w23012_ ;
	wire _w23013_ ;
	wire _w23014_ ;
	wire _w23015_ ;
	wire _w23016_ ;
	wire _w23017_ ;
	wire _w23018_ ;
	wire _w23019_ ;
	wire _w23020_ ;
	wire _w23021_ ;
	wire _w23022_ ;
	wire _w23023_ ;
	wire _w23024_ ;
	wire _w23025_ ;
	wire _w23026_ ;
	wire _w23027_ ;
	wire _w23028_ ;
	wire _w23029_ ;
	wire _w23030_ ;
	wire _w23031_ ;
	wire _w23032_ ;
	wire _w23033_ ;
	wire _w23034_ ;
	wire _w23035_ ;
	wire _w23036_ ;
	wire _w23037_ ;
	wire _w23038_ ;
	wire _w23039_ ;
	wire _w23040_ ;
	wire _w23041_ ;
	wire _w23042_ ;
	wire _w23043_ ;
	wire _w23044_ ;
	wire _w23045_ ;
	wire _w23046_ ;
	wire _w23047_ ;
	wire _w23048_ ;
	wire _w23049_ ;
	wire _w23050_ ;
	wire _w23051_ ;
	wire _w23052_ ;
	wire _w23053_ ;
	wire _w23054_ ;
	wire _w23055_ ;
	wire _w23056_ ;
	wire _w23057_ ;
	wire _w23058_ ;
	wire _w23059_ ;
	wire _w23060_ ;
	wire _w23061_ ;
	wire _w23062_ ;
	wire _w23063_ ;
	wire _w23064_ ;
	wire _w23065_ ;
	wire _w23066_ ;
	wire _w23067_ ;
	wire _w23068_ ;
	wire _w23069_ ;
	wire _w23070_ ;
	wire _w23071_ ;
	wire _w23072_ ;
	wire _w23073_ ;
	wire _w23074_ ;
	wire _w23075_ ;
	wire _w23076_ ;
	wire _w23077_ ;
	wire _w23078_ ;
	wire _w23079_ ;
	wire _w23080_ ;
	wire _w23081_ ;
	wire _w23082_ ;
	wire _w23083_ ;
	wire _w23084_ ;
	wire _w23085_ ;
	wire _w23086_ ;
	wire _w23087_ ;
	wire _w23088_ ;
	wire _w23089_ ;
	wire _w23090_ ;
	wire _w23091_ ;
	wire _w23092_ ;
	wire _w23093_ ;
	wire _w23094_ ;
	wire _w23095_ ;
	wire _w23096_ ;
	wire _w23097_ ;
	wire _w23098_ ;
	wire _w23099_ ;
	wire _w23100_ ;
	wire _w23101_ ;
	wire _w23102_ ;
	wire _w23103_ ;
	wire _w23104_ ;
	wire _w23105_ ;
	wire _w23106_ ;
	wire _w23107_ ;
	wire _w23108_ ;
	wire _w23109_ ;
	wire _w23110_ ;
	wire _w23111_ ;
	wire _w23112_ ;
	wire _w23113_ ;
	wire _w23114_ ;
	wire _w23115_ ;
	wire _w23116_ ;
	wire _w23117_ ;
	wire _w23118_ ;
	wire _w23119_ ;
	wire _w23120_ ;
	wire _w23121_ ;
	wire _w23122_ ;
	wire _w23123_ ;
	wire _w23124_ ;
	wire _w23125_ ;
	wire _w23126_ ;
	wire _w23127_ ;
	wire _w23128_ ;
	wire _w23129_ ;
	wire _w23130_ ;
	wire _w23131_ ;
	wire _w23132_ ;
	wire _w23133_ ;
	wire _w23134_ ;
	wire _w23135_ ;
	wire _w23136_ ;
	wire _w23137_ ;
	wire _w23138_ ;
	wire _w23139_ ;
	wire _w23140_ ;
	wire _w23141_ ;
	wire _w23142_ ;
	wire _w23143_ ;
	wire _w23144_ ;
	wire _w23145_ ;
	wire _w23146_ ;
	wire _w23147_ ;
	wire _w23148_ ;
	wire _w23149_ ;
	wire _w23150_ ;
	wire _w23151_ ;
	wire _w23152_ ;
	wire _w23153_ ;
	wire _w23154_ ;
	wire _w23155_ ;
	wire _w23156_ ;
	wire _w23157_ ;
	wire _w23158_ ;
	wire _w23159_ ;
	wire _w23160_ ;
	wire _w23161_ ;
	wire _w23162_ ;
	wire _w23163_ ;
	wire _w23164_ ;
	wire _w23165_ ;
	wire _w23166_ ;
	wire _w23167_ ;
	wire _w23168_ ;
	wire _w23169_ ;
	wire _w23170_ ;
	wire _w23171_ ;
	wire _w23172_ ;
	wire _w23173_ ;
	wire _w23174_ ;
	wire _w23175_ ;
	wire _w23176_ ;
	wire _w23177_ ;
	wire _w23178_ ;
	wire _w23179_ ;
	wire _w23180_ ;
	wire _w23181_ ;
	wire _w23182_ ;
	wire _w23183_ ;
	wire _w23184_ ;
	wire _w23185_ ;
	wire _w23186_ ;
	wire _w23187_ ;
	wire _w23188_ ;
	wire _w23189_ ;
	wire _w23190_ ;
	wire _w23191_ ;
	wire _w23192_ ;
	wire _w23193_ ;
	wire _w23194_ ;
	wire _w23195_ ;
	wire _w23196_ ;
	wire _w23197_ ;
	wire _w23198_ ;
	wire _w23199_ ;
	wire _w23200_ ;
	wire _w23201_ ;
	wire _w23202_ ;
	wire _w23203_ ;
	wire _w23204_ ;
	wire _w23205_ ;
	wire _w23206_ ;
	wire _w23207_ ;
	wire _w23208_ ;
	wire _w23209_ ;
	wire _w23210_ ;
	wire _w23211_ ;
	wire _w23212_ ;
	wire _w23213_ ;
	wire _w23214_ ;
	wire _w23215_ ;
	wire _w23216_ ;
	wire _w23217_ ;
	wire _w23218_ ;
	wire _w23219_ ;
	wire _w23220_ ;
	wire _w23221_ ;
	wire _w23222_ ;
	wire _w23223_ ;
	wire _w23224_ ;
	wire _w23225_ ;
	wire _w23226_ ;
	wire _w23227_ ;
	wire _w23228_ ;
	wire _w23229_ ;
	wire _w23230_ ;
	wire _w23231_ ;
	wire _w23232_ ;
	wire _w23233_ ;
	wire _w23234_ ;
	wire _w23235_ ;
	wire _w23236_ ;
	wire _w23237_ ;
	wire _w23238_ ;
	wire _w23239_ ;
	wire _w23240_ ;
	wire _w23241_ ;
	wire _w23242_ ;
	wire _w23243_ ;
	wire _w23244_ ;
	wire _w23245_ ;
	wire _w23246_ ;
	wire _w23247_ ;
	wire _w23248_ ;
	wire _w23249_ ;
	wire _w23250_ ;
	wire _w23251_ ;
	wire _w23252_ ;
	wire _w23253_ ;
	wire _w23254_ ;
	wire _w23255_ ;
	wire _w23256_ ;
	wire _w23257_ ;
	wire _w23258_ ;
	wire _w23259_ ;
	wire _w23260_ ;
	wire _w23261_ ;
	wire _w23262_ ;
	wire _w23263_ ;
	wire _w23264_ ;
	wire _w23265_ ;
	wire _w23266_ ;
	wire _w23267_ ;
	wire _w23268_ ;
	wire _w23269_ ;
	wire _w23270_ ;
	wire _w23271_ ;
	wire _w23272_ ;
	wire _w23273_ ;
	wire _w23274_ ;
	wire _w23275_ ;
	wire _w23276_ ;
	wire _w23277_ ;
	wire _w23278_ ;
	wire _w23279_ ;
	wire _w23280_ ;
	wire _w23281_ ;
	wire _w23282_ ;
	wire _w23283_ ;
	wire _w23284_ ;
	wire _w23285_ ;
	wire _w23286_ ;
	wire _w23287_ ;
	wire _w23288_ ;
	wire _w23289_ ;
	wire _w23290_ ;
	wire _w23291_ ;
	wire _w23292_ ;
	wire _w23293_ ;
	wire _w23294_ ;
	wire _w23295_ ;
	wire _w23296_ ;
	wire _w23297_ ;
	wire _w23298_ ;
	wire _w23299_ ;
	wire _w23300_ ;
	wire _w23301_ ;
	wire _w23302_ ;
	wire _w23303_ ;
	wire _w23304_ ;
	wire _w23305_ ;
	wire _w23306_ ;
	wire _w23307_ ;
	wire _w23308_ ;
	wire _w23309_ ;
	wire _w23310_ ;
	wire _w23311_ ;
	wire _w23312_ ;
	wire _w23313_ ;
	wire _w23314_ ;
	wire _w23315_ ;
	wire _w23316_ ;
	wire _w23317_ ;
	wire _w23318_ ;
	wire _w23319_ ;
	wire _w23320_ ;
	wire _w23321_ ;
	wire _w23322_ ;
	wire _w23323_ ;
	wire _w23324_ ;
	wire _w23325_ ;
	wire _w23326_ ;
	wire _w23327_ ;
	wire _w23328_ ;
	wire _w23329_ ;
	wire _w23330_ ;
	wire _w23331_ ;
	wire _w23332_ ;
	wire _w23333_ ;
	wire _w23334_ ;
	wire _w23335_ ;
	wire _w23336_ ;
	wire _w23337_ ;
	wire _w23338_ ;
	wire _w23339_ ;
	wire _w23340_ ;
	wire _w23341_ ;
	wire _w23342_ ;
	wire _w23343_ ;
	wire _w23344_ ;
	wire _w23345_ ;
	wire _w23346_ ;
	wire _w23347_ ;
	wire _w23348_ ;
	wire _w23349_ ;
	wire _w23350_ ;
	wire _w23351_ ;
	wire _w23352_ ;
	wire _w23353_ ;
	wire _w23354_ ;
	wire _w23355_ ;
	wire _w23356_ ;
	wire _w23357_ ;
	wire _w23358_ ;
	wire _w23359_ ;
	wire _w23360_ ;
	wire _w23361_ ;
	wire _w23362_ ;
	wire _w23363_ ;
	wire _w23364_ ;
	wire _w23365_ ;
	wire _w23366_ ;
	wire _w23367_ ;
	wire _w23368_ ;
	wire _w23369_ ;
	wire _w23370_ ;
	wire _w23371_ ;
	wire _w23372_ ;
	wire _w23373_ ;
	wire _w23374_ ;
	wire _w23375_ ;
	wire _w23376_ ;
	wire _w23377_ ;
	wire _w23378_ ;
	wire _w23379_ ;
	wire _w23380_ ;
	wire _w23381_ ;
	wire _w23382_ ;
	wire _w23383_ ;
	wire _w23384_ ;
	wire _w23385_ ;
	wire _w23386_ ;
	wire _w23387_ ;
	wire _w23388_ ;
	wire _w23389_ ;
	wire _w23390_ ;
	wire _w23391_ ;
	wire _w23392_ ;
	wire _w23393_ ;
	wire _w23394_ ;
	wire _w23395_ ;
	wire _w23396_ ;
	wire _w23397_ ;
	wire _w23398_ ;
	wire _w23399_ ;
	wire _w23400_ ;
	wire _w23401_ ;
	wire _w23402_ ;
	wire _w23403_ ;
	wire _w23404_ ;
	wire _w23405_ ;
	wire _w23406_ ;
	wire _w23407_ ;
	wire _w23408_ ;
	wire _w23409_ ;
	wire _w23410_ ;
	wire _w23411_ ;
	wire _w23412_ ;
	wire _w23413_ ;
	wire _w23414_ ;
	wire _w23415_ ;
	wire _w23416_ ;
	wire _w23417_ ;
	wire _w23418_ ;
	wire _w23419_ ;
	wire _w23420_ ;
	wire _w23421_ ;
	wire _w23422_ ;
	wire _w23423_ ;
	wire _w23424_ ;
	wire _w23425_ ;
	wire _w23426_ ;
	wire _w23427_ ;
	wire _w23428_ ;
	wire _w23429_ ;
	wire _w23430_ ;
	wire _w23431_ ;
	wire _w23432_ ;
	wire _w23433_ ;
	wire _w23434_ ;
	wire _w23435_ ;
	wire _w23436_ ;
	wire _w23437_ ;
	wire _w23438_ ;
	wire _w23439_ ;
	wire _w23440_ ;
	wire _w23441_ ;
	wire _w23442_ ;
	wire _w23443_ ;
	wire _w23444_ ;
	wire _w23445_ ;
	wire _w23446_ ;
	wire _w23447_ ;
	wire _w23448_ ;
	wire _w23449_ ;
	wire _w23450_ ;
	wire _w23451_ ;
	wire _w23452_ ;
	wire _w23453_ ;
	wire _w23454_ ;
	wire _w23455_ ;
	wire _w23456_ ;
	wire _w23457_ ;
	wire _w23458_ ;
	wire _w23459_ ;
	wire _w23460_ ;
	wire _w23461_ ;
	wire _w23462_ ;
	wire _w23463_ ;
	wire _w23464_ ;
	wire _w23465_ ;
	wire _w23466_ ;
	wire _w23467_ ;
	wire _w23468_ ;
	wire _w23469_ ;
	wire _w23470_ ;
	wire _w23471_ ;
	wire _w23472_ ;
	wire _w23473_ ;
	wire _w23474_ ;
	wire _w23475_ ;
	wire _w23476_ ;
	wire _w23477_ ;
	wire _w23478_ ;
	wire _w23479_ ;
	wire _w23480_ ;
	wire _w23481_ ;
	wire _w23482_ ;
	wire _w23483_ ;
	wire _w23484_ ;
	wire _w23485_ ;
	wire _w23486_ ;
	wire _w23487_ ;
	wire _w23488_ ;
	wire _w23489_ ;
	wire _w23490_ ;
	wire _w23491_ ;
	wire _w23492_ ;
	wire _w23493_ ;
	wire _w23494_ ;
	wire _w23495_ ;
	wire _w23496_ ;
	wire _w23497_ ;
	wire _w23498_ ;
	wire _w23499_ ;
	wire _w23500_ ;
	wire _w23501_ ;
	wire _w23502_ ;
	wire _w23503_ ;
	wire _w23504_ ;
	wire _w23505_ ;
	wire _w23506_ ;
	wire _w23507_ ;
	wire _w23508_ ;
	wire _w23509_ ;
	wire _w23510_ ;
	wire _w23511_ ;
	wire _w23512_ ;
	wire _w23513_ ;
	wire _w23514_ ;
	wire _w23515_ ;
	wire _w23516_ ;
	wire _w23517_ ;
	wire _w23518_ ;
	wire _w23519_ ;
	wire _w23520_ ;
	wire _w23521_ ;
	wire _w23522_ ;
	wire _w23523_ ;
	wire _w23524_ ;
	wire _w23525_ ;
	wire _w23526_ ;
	wire _w23527_ ;
	wire _w23528_ ;
	wire _w23529_ ;
	wire _w23530_ ;
	wire _w23531_ ;
	wire _w23532_ ;
	wire _w23533_ ;
	wire _w23534_ ;
	wire _w23535_ ;
	wire _w23536_ ;
	wire _w23537_ ;
	wire _w23538_ ;
	wire _w23539_ ;
	wire _w23540_ ;
	wire _w23541_ ;
	wire _w23542_ ;
	wire _w23543_ ;
	wire _w23544_ ;
	wire _w23545_ ;
	wire _w23546_ ;
	wire _w23547_ ;
	wire _w23548_ ;
	wire _w23549_ ;
	wire _w23550_ ;
	wire _w23551_ ;
	wire _w23552_ ;
	wire _w23553_ ;
	wire _w23554_ ;
	wire _w23555_ ;
	wire _w23556_ ;
	wire _w23557_ ;
	wire _w23558_ ;
	wire _w23559_ ;
	wire _w23560_ ;
	wire _w23561_ ;
	wire _w23562_ ;
	wire _w23563_ ;
	wire _w23564_ ;
	wire _w23565_ ;
	wire _w23566_ ;
	wire _w23567_ ;
	wire _w23568_ ;
	wire _w23569_ ;
	wire _w23570_ ;
	wire _w23571_ ;
	wire _w23572_ ;
	wire _w23573_ ;
	wire _w23574_ ;
	wire _w23575_ ;
	wire _w23576_ ;
	wire _w23577_ ;
	wire _w23578_ ;
	wire _w23579_ ;
	wire _w23580_ ;
	wire _w23581_ ;
	wire _w23582_ ;
	wire _w23583_ ;
	wire _w23584_ ;
	wire _w23585_ ;
	wire _w23586_ ;
	wire _w23587_ ;
	wire _w23588_ ;
	wire _w23589_ ;
	wire _w23590_ ;
	wire _w23591_ ;
	wire _w23592_ ;
	wire _w23593_ ;
	wire _w23594_ ;
	wire _w23595_ ;
	wire _w23596_ ;
	wire _w23597_ ;
	wire _w23598_ ;
	wire _w23599_ ;
	wire _w23600_ ;
	wire _w23601_ ;
	wire _w23602_ ;
	wire _w23603_ ;
	wire _w23604_ ;
	wire _w23605_ ;
	wire _w23606_ ;
	wire _w23607_ ;
	wire _w23608_ ;
	wire _w23609_ ;
	wire _w23610_ ;
	wire _w23611_ ;
	wire _w23612_ ;
	wire _w23613_ ;
	wire _w23614_ ;
	wire _w23615_ ;
	wire _w23616_ ;
	wire _w23617_ ;
	wire _w23618_ ;
	wire _w23619_ ;
	wire _w23620_ ;
	wire _w23621_ ;
	wire _w23622_ ;
	wire _w23623_ ;
	wire _w23624_ ;
	wire _w23625_ ;
	wire _w23626_ ;
	wire _w23627_ ;
	wire _w23628_ ;
	wire _w23629_ ;
	wire _w23630_ ;
	wire _w23631_ ;
	wire _w23632_ ;
	wire _w23633_ ;
	wire _w23634_ ;
	wire _w23635_ ;
	wire _w23636_ ;
	wire _w23637_ ;
	wire _w23638_ ;
	wire _w23639_ ;
	wire _w23640_ ;
	wire _w23641_ ;
	wire _w23642_ ;
	wire _w23643_ ;
	wire _w23644_ ;
	wire _w23645_ ;
	wire _w23646_ ;
	wire _w23647_ ;
	wire _w23648_ ;
	wire _w23649_ ;
	wire _w23650_ ;
	wire _w23651_ ;
	wire _w23652_ ;
	wire _w23653_ ;
	wire _w23654_ ;
	wire _w23655_ ;
	wire _w23656_ ;
	wire _w23657_ ;
	wire _w23658_ ;
	wire _w23659_ ;
	wire _w23660_ ;
	wire _w23661_ ;
	wire _w23662_ ;
	wire _w23663_ ;
	wire _w23664_ ;
	wire _w23665_ ;
	wire _w23666_ ;
	wire _w23667_ ;
	wire _w23668_ ;
	wire _w23669_ ;
	wire _w23670_ ;
	wire _w23671_ ;
	wire _w23672_ ;
	wire _w23673_ ;
	wire _w23674_ ;
	wire _w23675_ ;
	wire _w23676_ ;
	wire _w23677_ ;
	wire _w23678_ ;
	wire _w23679_ ;
	wire _w23680_ ;
	wire _w23681_ ;
	wire _w23682_ ;
	wire _w23683_ ;
	wire _w23684_ ;
	wire _w23685_ ;
	wire _w23686_ ;
	wire _w23687_ ;
	wire _w23688_ ;
	wire _w23689_ ;
	wire _w23690_ ;
	wire _w23691_ ;
	wire _w23692_ ;
	wire _w23693_ ;
	wire _w23694_ ;
	wire _w23695_ ;
	wire _w23696_ ;
	wire _w23697_ ;
	wire _w23698_ ;
	wire _w23699_ ;
	wire _w23700_ ;
	wire _w23701_ ;
	wire _w23702_ ;
	wire _w23703_ ;
	wire _w23704_ ;
	wire _w23705_ ;
	wire _w23706_ ;
	wire _w23707_ ;
	wire _w23708_ ;
	wire _w23709_ ;
	wire _w23710_ ;
	wire _w23711_ ;
	wire _w23712_ ;
	wire _w23713_ ;
	wire _w23714_ ;
	wire _w23715_ ;
	wire _w23716_ ;
	wire _w23717_ ;
	wire _w23718_ ;
	wire _w23719_ ;
	wire _w23720_ ;
	wire _w23721_ ;
	wire _w23722_ ;
	wire _w23723_ ;
	wire _w23724_ ;
	wire _w23725_ ;
	wire _w23726_ ;
	wire _w23727_ ;
	wire _w23728_ ;
	wire _w23729_ ;
	wire _w23730_ ;
	wire _w23731_ ;
	wire _w23732_ ;
	wire _w23733_ ;
	wire _w23734_ ;
	wire _w23735_ ;
	wire _w23736_ ;
	wire _w23737_ ;
	wire _w23738_ ;
	wire _w23739_ ;
	wire _w23740_ ;
	wire _w23741_ ;
	wire _w23742_ ;
	wire _w23743_ ;
	wire _w23744_ ;
	wire _w23745_ ;
	wire _w23746_ ;
	wire _w23747_ ;
	wire _w23748_ ;
	wire _w23749_ ;
	wire _w23750_ ;
	wire _w23751_ ;
	wire _w23752_ ;
	wire _w23753_ ;
	wire _w23754_ ;
	wire _w23755_ ;
	wire _w23756_ ;
	wire _w23757_ ;
	wire _w23758_ ;
	wire _w23759_ ;
	wire _w23760_ ;
	wire _w23761_ ;
	wire _w23762_ ;
	wire _w23763_ ;
	wire _w23764_ ;
	wire _w23765_ ;
	wire _w23766_ ;
	wire _w23767_ ;
	wire _w23768_ ;
	wire _w23769_ ;
	wire _w23770_ ;
	wire _w23771_ ;
	wire _w23772_ ;
	wire _w23773_ ;
	wire _w23774_ ;
	wire _w23775_ ;
	wire _w23776_ ;
	wire _w23777_ ;
	wire _w23778_ ;
	wire _w23779_ ;
	wire _w23780_ ;
	wire _w23781_ ;
	wire _w23782_ ;
	wire _w23783_ ;
	wire _w23784_ ;
	wire _w23785_ ;
	wire _w23786_ ;
	wire _w23787_ ;
	wire _w23788_ ;
	wire _w23789_ ;
	wire _w23790_ ;
	wire _w23791_ ;
	wire _w23792_ ;
	wire _w23793_ ;
	wire _w23794_ ;
	wire _w23795_ ;
	wire _w23796_ ;
	wire _w23797_ ;
	wire _w23798_ ;
	wire _w23799_ ;
	wire _w23800_ ;
	wire _w23801_ ;
	wire _w23802_ ;
	wire _w23803_ ;
	wire _w23804_ ;
	wire _w23805_ ;
	wire _w23806_ ;
	wire _w23807_ ;
	wire _w23808_ ;
	wire _w23809_ ;
	wire _w23810_ ;
	wire _w23811_ ;
	wire _w23812_ ;
	wire _w23813_ ;
	wire _w23814_ ;
	wire _w23815_ ;
	wire _w23816_ ;
	wire _w23817_ ;
	wire _w23818_ ;
	wire _w23819_ ;
	wire _w23820_ ;
	wire _w23821_ ;
	wire _w23822_ ;
	wire _w23823_ ;
	wire _w23824_ ;
	wire _w23825_ ;
	wire _w23826_ ;
	wire _w23827_ ;
	wire _w23828_ ;
	wire _w23829_ ;
	wire _w23830_ ;
	wire _w23831_ ;
	wire _w23832_ ;
	wire _w23833_ ;
	wire _w23834_ ;
	wire _w23835_ ;
	wire _w23836_ ;
	wire _w23837_ ;
	wire _w23838_ ;
	wire _w23839_ ;
	wire _w23840_ ;
	wire _w23841_ ;
	wire _w23842_ ;
	wire _w23843_ ;
	wire _w23844_ ;
	wire _w23845_ ;
	wire _w23846_ ;
	wire _w23847_ ;
	wire _w23848_ ;
	wire _w23849_ ;
	wire _w23850_ ;
	wire _w23851_ ;
	wire _w23852_ ;
	wire _w23853_ ;
	wire _w23854_ ;
	wire _w23855_ ;
	wire _w23856_ ;
	wire _w23857_ ;
	wire _w23858_ ;
	wire _w23859_ ;
	wire _w23860_ ;
	wire _w23861_ ;
	wire _w23862_ ;
	wire _w23863_ ;
	wire _w23864_ ;
	wire _w23865_ ;
	wire _w23866_ ;
	wire _w23867_ ;
	wire _w23868_ ;
	wire _w23869_ ;
	wire _w23870_ ;
	wire _w23871_ ;
	wire _w23872_ ;
	wire _w23873_ ;
	wire _w23874_ ;
	wire _w23875_ ;
	wire _w23876_ ;
	wire _w23877_ ;
	wire _w23878_ ;
	wire _w23879_ ;
	wire _w23880_ ;
	wire _w23881_ ;
	wire _w23882_ ;
	wire _w23883_ ;
	wire _w23884_ ;
	wire _w23885_ ;
	wire _w23886_ ;
	wire _w23887_ ;
	wire _w23888_ ;
	wire _w23889_ ;
	wire _w23890_ ;
	wire _w23891_ ;
	wire _w23892_ ;
	wire _w23893_ ;
	wire _w23894_ ;
	wire _w23895_ ;
	wire _w23896_ ;
	wire _w23897_ ;
	wire _w23898_ ;
	wire _w23899_ ;
	wire _w23900_ ;
	wire _w23901_ ;
	wire _w23902_ ;
	wire _w23903_ ;
	wire _w23904_ ;
	wire _w23905_ ;
	wire _w23906_ ;
	wire _w23907_ ;
	wire _w23908_ ;
	wire _w23909_ ;
	wire _w23910_ ;
	wire _w23911_ ;
	wire _w23912_ ;
	wire _w23913_ ;
	wire _w23914_ ;
	wire _w23915_ ;
	wire _w23916_ ;
	wire _w23917_ ;
	wire _w23918_ ;
	wire _w23919_ ;
	wire _w23920_ ;
	wire _w23921_ ;
	wire _w23922_ ;
	wire _w23923_ ;
	wire _w23924_ ;
	wire _w23925_ ;
	wire _w23926_ ;
	wire _w23927_ ;
	wire _w23928_ ;
	wire _w23929_ ;
	wire _w23930_ ;
	wire _w23931_ ;
	wire _w23932_ ;
	wire _w23933_ ;
	wire _w23934_ ;
	wire _w23935_ ;
	wire _w23936_ ;
	wire _w23937_ ;
	wire _w23938_ ;
	wire _w23939_ ;
	wire _w23940_ ;
	wire _w23941_ ;
	wire _w23942_ ;
	wire _w23943_ ;
	wire _w23944_ ;
	wire _w23945_ ;
	wire _w23946_ ;
	wire _w23947_ ;
	wire _w23948_ ;
	wire _w23949_ ;
	wire _w23950_ ;
	wire _w23951_ ;
	wire _w23952_ ;
	wire _w23953_ ;
	wire _w23954_ ;
	wire _w23955_ ;
	wire _w23956_ ;
	wire _w23957_ ;
	wire _w23958_ ;
	wire _w23959_ ;
	wire _w23960_ ;
	wire _w23961_ ;
	wire _w23962_ ;
	wire _w23963_ ;
	wire _w23964_ ;
	wire _w23965_ ;
	wire _w23966_ ;
	wire _w23967_ ;
	wire _w23968_ ;
	wire _w23969_ ;
	wire _w23970_ ;
	wire _w23971_ ;
	wire _w23972_ ;
	wire _w23973_ ;
	wire _w23974_ ;
	wire _w23975_ ;
	wire _w23976_ ;
	wire _w23977_ ;
	wire _w23978_ ;
	wire _w23979_ ;
	wire _w23980_ ;
	wire _w23981_ ;
	wire _w23982_ ;
	wire _w23983_ ;
	wire _w23984_ ;
	wire _w23985_ ;
	wire _w23986_ ;
	wire _w23987_ ;
	wire _w23988_ ;
	wire _w23989_ ;
	wire _w23990_ ;
	wire _w23991_ ;
	wire _w23992_ ;
	wire _w23993_ ;
	wire _w23994_ ;
	wire _w23995_ ;
	wire _w23996_ ;
	wire _w23997_ ;
	wire _w23998_ ;
	wire _w23999_ ;
	wire _w24000_ ;
	wire _w24001_ ;
	wire _w24002_ ;
	wire _w24003_ ;
	wire _w24004_ ;
	wire _w24005_ ;
	wire _w24006_ ;
	wire _w24007_ ;
	wire _w24008_ ;
	wire _w24009_ ;
	wire _w24010_ ;
	wire _w24011_ ;
	wire _w24012_ ;
	wire _w24013_ ;
	wire _w24014_ ;
	wire _w24015_ ;
	wire _w24016_ ;
	wire _w24017_ ;
	wire _w24018_ ;
	wire _w24019_ ;
	wire _w24020_ ;
	wire _w24021_ ;
	wire _w24022_ ;
	wire _w24023_ ;
	wire _w24024_ ;
	wire _w24025_ ;
	wire _w24026_ ;
	wire _w24027_ ;
	wire _w24028_ ;
	wire _w24029_ ;
	wire _w24030_ ;
	wire _w24031_ ;
	wire _w24032_ ;
	wire _w24033_ ;
	wire _w24034_ ;
	wire _w24035_ ;
	wire _w24036_ ;
	wire _w24037_ ;
	wire _w24038_ ;
	wire _w24039_ ;
	wire _w24040_ ;
	wire _w24041_ ;
	wire _w24042_ ;
	wire _w24043_ ;
	wire _w24044_ ;
	wire _w24045_ ;
	wire _w24046_ ;
	wire _w24047_ ;
	wire _w24048_ ;
	wire _w24049_ ;
	wire _w24050_ ;
	wire _w24051_ ;
	wire _w24052_ ;
	wire _w24053_ ;
	wire _w24054_ ;
	wire _w24055_ ;
	wire _w24056_ ;
	wire _w24057_ ;
	wire _w24058_ ;
	wire _w24059_ ;
	wire _w24060_ ;
	wire _w24061_ ;
	wire _w24062_ ;
	wire _w24063_ ;
	wire _w24064_ ;
	wire _w24065_ ;
	wire _w24066_ ;
	wire _w24067_ ;
	wire _w24068_ ;
	wire _w24069_ ;
	wire _w24070_ ;
	wire _w24071_ ;
	wire _w24072_ ;
	wire _w24073_ ;
	wire _w24074_ ;
	wire _w24075_ ;
	wire _w24076_ ;
	wire _w24077_ ;
	wire _w24078_ ;
	wire _w24079_ ;
	wire _w24080_ ;
	wire _w24081_ ;
	wire _w24082_ ;
	wire _w24083_ ;
	wire _w24084_ ;
	wire _w24085_ ;
	wire _w24086_ ;
	wire _w24087_ ;
	wire _w24088_ ;
	wire _w24089_ ;
	wire _w24090_ ;
	wire _w24091_ ;
	wire _w24092_ ;
	wire _w24093_ ;
	wire _w24094_ ;
	wire _w24095_ ;
	wire _w24096_ ;
	wire _w24097_ ;
	wire _w24098_ ;
	wire _w24099_ ;
	wire _w24100_ ;
	wire _w24101_ ;
	wire _w24102_ ;
	wire _w24103_ ;
	wire _w24104_ ;
	wire _w24105_ ;
	wire _w24106_ ;
	wire _w24107_ ;
	wire _w24108_ ;
	wire _w24109_ ;
	wire _w24110_ ;
	wire _w24111_ ;
	wire _w24112_ ;
	wire _w24113_ ;
	wire _w24114_ ;
	wire _w24115_ ;
	wire _w24116_ ;
	wire _w24117_ ;
	wire _w24118_ ;
	wire _w24119_ ;
	wire _w24120_ ;
	wire _w24121_ ;
	wire _w24122_ ;
	wire _w24123_ ;
	wire _w24124_ ;
	wire _w24125_ ;
	wire _w24126_ ;
	wire _w24127_ ;
	wire _w24128_ ;
	wire _w24129_ ;
	wire _w24130_ ;
	wire _w24131_ ;
	wire _w24132_ ;
	wire _w24133_ ;
	wire _w24134_ ;
	wire _w24135_ ;
	wire _w24136_ ;
	wire _w24137_ ;
	wire _w24138_ ;
	wire _w24139_ ;
	wire _w24140_ ;
	wire _w24141_ ;
	wire _w24142_ ;
	wire _w24143_ ;
	wire _w24144_ ;
	wire _w24145_ ;
	wire _w24146_ ;
	wire _w24147_ ;
	wire _w24148_ ;
	wire _w24149_ ;
	wire _w24150_ ;
	wire _w24151_ ;
	wire _w24152_ ;
	wire _w24153_ ;
	wire _w24154_ ;
	wire _w24155_ ;
	wire _w24156_ ;
	wire _w24157_ ;
	wire _w24158_ ;
	wire _w24159_ ;
	wire _w24160_ ;
	wire _w24161_ ;
	wire _w24162_ ;
	wire _w24163_ ;
	wire _w24164_ ;
	wire _w24165_ ;
	wire _w24166_ ;
	wire _w24167_ ;
	wire _w24168_ ;
	wire _w24169_ ;
	wire _w24170_ ;
	wire _w24171_ ;
	wire _w24172_ ;
	wire _w24173_ ;
	wire _w24174_ ;
	wire _w24175_ ;
	wire _w24176_ ;
	wire _w24177_ ;
	wire _w24178_ ;
	wire _w24179_ ;
	wire _w24180_ ;
	wire _w24181_ ;
	wire _w24182_ ;
	wire _w24183_ ;
	wire _w24184_ ;
	wire _w24185_ ;
	wire _w24186_ ;
	wire _w24187_ ;
	wire _w24188_ ;
	wire _w24189_ ;
	wire _w24190_ ;
	wire _w24191_ ;
	wire _w24192_ ;
	wire _w24193_ ;
	wire _w24194_ ;
	wire _w24195_ ;
	wire _w24196_ ;
	wire _w24197_ ;
	wire _w24198_ ;
	wire _w24199_ ;
	wire _w24200_ ;
	wire _w24201_ ;
	wire _w24202_ ;
	wire _w24203_ ;
	wire _w24204_ ;
	wire _w24205_ ;
	wire _w24206_ ;
	wire _w24207_ ;
	wire _w24208_ ;
	wire _w24209_ ;
	wire _w24210_ ;
	wire _w24211_ ;
	wire _w24212_ ;
	wire _w24213_ ;
	wire _w24214_ ;
	wire _w24215_ ;
	wire _w24216_ ;
	wire _w24217_ ;
	wire _w24218_ ;
	wire _w24219_ ;
	wire _w24220_ ;
	wire _w24221_ ;
	wire _w24222_ ;
	wire _w24223_ ;
	wire _w24224_ ;
	wire _w24225_ ;
	wire _w24226_ ;
	wire _w24227_ ;
	wire _w24228_ ;
	wire _w24229_ ;
	wire _w24230_ ;
	wire _w24231_ ;
	wire _w24232_ ;
	wire _w24233_ ;
	wire _w24234_ ;
	wire _w24235_ ;
	wire _w24236_ ;
	wire _w24237_ ;
	wire _w24238_ ;
	wire _w24239_ ;
	wire _w24240_ ;
	wire _w24241_ ;
	wire _w24242_ ;
	wire _w24243_ ;
	wire _w24244_ ;
	wire _w24245_ ;
	wire _w24246_ ;
	wire _w24247_ ;
	wire _w24248_ ;
	wire _w24249_ ;
	wire _w24250_ ;
	wire _w24251_ ;
	wire _w24252_ ;
	wire _w24253_ ;
	wire _w24254_ ;
	wire _w24255_ ;
	wire _w24256_ ;
	wire _w24257_ ;
	wire _w24258_ ;
	wire _w24259_ ;
	wire _w24260_ ;
	wire _w24261_ ;
	wire _w24262_ ;
	wire _w24263_ ;
	wire _w24264_ ;
	wire _w24265_ ;
	wire _w24266_ ;
	wire _w24267_ ;
	wire _w24268_ ;
	wire _w24269_ ;
	wire _w24270_ ;
	wire _w24271_ ;
	wire _w24272_ ;
	wire _w24273_ ;
	wire _w24274_ ;
	wire _w24275_ ;
	wire _w24276_ ;
	wire _w24277_ ;
	wire _w24278_ ;
	wire _w24279_ ;
	wire _w24280_ ;
	wire _w24281_ ;
	wire _w24282_ ;
	wire _w24283_ ;
	wire _w24284_ ;
	wire _w24285_ ;
	wire _w24286_ ;
	wire _w24287_ ;
	wire _w24288_ ;
	wire _w24289_ ;
	wire _w24290_ ;
	wire _w24291_ ;
	wire _w24292_ ;
	wire _w24293_ ;
	wire _w24294_ ;
	wire _w24295_ ;
	wire _w24296_ ;
	wire _w24297_ ;
	wire _w24298_ ;
	wire _w24299_ ;
	wire _w24300_ ;
	wire _w24301_ ;
	wire _w24302_ ;
	wire _w24303_ ;
	wire _w24304_ ;
	wire _w24305_ ;
	wire _w24306_ ;
	wire _w24307_ ;
	wire _w24308_ ;
	wire _w24309_ ;
	wire _w24310_ ;
	wire _w24311_ ;
	wire _w24312_ ;
	wire _w24313_ ;
	wire _w24314_ ;
	wire _w24315_ ;
	wire _w24316_ ;
	wire _w24317_ ;
	wire _w24318_ ;
	wire _w24319_ ;
	wire _w24320_ ;
	wire _w24321_ ;
	wire _w24322_ ;
	wire _w24323_ ;
	wire _w24324_ ;
	wire _w24325_ ;
	wire _w24326_ ;
	wire _w24327_ ;
	wire _w24328_ ;
	wire _w24329_ ;
	wire _w24330_ ;
	wire _w24331_ ;
	wire _w24332_ ;
	wire _w24333_ ;
	wire _w24334_ ;
	wire _w24335_ ;
	wire _w24336_ ;
	wire _w24337_ ;
	wire _w24338_ ;
	wire _w24339_ ;
	wire _w24340_ ;
	wire _w24341_ ;
	wire _w24342_ ;
	wire _w24343_ ;
	wire _w24344_ ;
	wire _w24345_ ;
	wire _w24346_ ;
	wire _w24347_ ;
	wire _w24348_ ;
	wire _w24349_ ;
	wire _w24350_ ;
	wire _w24351_ ;
	wire _w24352_ ;
	wire _w24353_ ;
	wire _w24354_ ;
	wire _w24355_ ;
	wire _w24356_ ;
	wire _w24357_ ;
	wire _w24358_ ;
	wire _w24359_ ;
	wire _w24360_ ;
	wire _w24361_ ;
	wire _w24362_ ;
	wire _w24363_ ;
	wire _w24364_ ;
	wire _w24365_ ;
	wire _w24366_ ;
	wire _w24367_ ;
	wire _w24368_ ;
	wire _w24369_ ;
	wire _w24370_ ;
	wire _w24371_ ;
	wire _w24372_ ;
	wire _w24373_ ;
	wire _w24374_ ;
	wire _w24375_ ;
	wire _w24376_ ;
	wire _w24377_ ;
	wire _w24378_ ;
	wire _w24379_ ;
	wire _w24380_ ;
	wire _w24381_ ;
	wire _w24382_ ;
	wire _w24383_ ;
	wire _w24384_ ;
	wire _w24385_ ;
	wire _w24386_ ;
	wire _w24387_ ;
	wire _w24388_ ;
	wire _w24389_ ;
	wire _w24390_ ;
	wire _w24391_ ;
	wire _w24392_ ;
	wire _w24393_ ;
	wire _w24394_ ;
	wire _w24395_ ;
	wire _w24396_ ;
	wire _w24397_ ;
	wire _w24398_ ;
	wire _w24399_ ;
	wire _w24400_ ;
	wire _w24401_ ;
	wire _w24402_ ;
	wire _w24403_ ;
	wire _w24404_ ;
	wire _w24405_ ;
	wire _w24406_ ;
	wire _w24407_ ;
	wire _w24408_ ;
	wire _w24409_ ;
	wire _w24410_ ;
	wire _w24411_ ;
	wire _w24412_ ;
	wire _w24413_ ;
	wire _w24414_ ;
	wire _w24415_ ;
	wire _w24416_ ;
	wire _w24417_ ;
	wire _w24418_ ;
	wire _w24419_ ;
	wire _w24420_ ;
	wire _w24421_ ;
	wire _w24422_ ;
	wire _w24423_ ;
	wire _w24424_ ;
	wire _w24425_ ;
	wire _w24426_ ;
	wire _w24427_ ;
	wire _w24428_ ;
	wire _w24429_ ;
	wire _w24430_ ;
	wire _w24431_ ;
	wire _w24432_ ;
	wire _w24433_ ;
	wire _w24434_ ;
	wire _w24435_ ;
	wire _w24436_ ;
	wire _w24437_ ;
	wire _w24438_ ;
	wire _w24439_ ;
	wire _w24440_ ;
	wire _w24441_ ;
	wire _w24442_ ;
	wire _w24443_ ;
	wire _w24444_ ;
	wire _w24445_ ;
	wire _w24446_ ;
	wire _w24447_ ;
	wire _w24448_ ;
	wire _w24449_ ;
	wire _w24450_ ;
	wire _w24451_ ;
	wire _w24452_ ;
	wire _w24453_ ;
	wire _w24454_ ;
	wire _w24455_ ;
	wire _w24456_ ;
	wire _w24457_ ;
	wire _w24458_ ;
	wire _w24459_ ;
	wire _w24460_ ;
	wire _w24461_ ;
	wire _w24462_ ;
	wire _w24463_ ;
	wire _w24464_ ;
	wire _w24465_ ;
	wire _w24466_ ;
	wire _w24467_ ;
	wire _w24468_ ;
	wire _w24469_ ;
	wire _w24470_ ;
	wire _w24471_ ;
	wire _w24472_ ;
	wire _w24473_ ;
	wire _w24474_ ;
	wire _w24475_ ;
	wire _w24476_ ;
	wire _w24477_ ;
	wire _w24478_ ;
	wire _w24479_ ;
	wire _w24480_ ;
	wire _w24481_ ;
	wire _w24482_ ;
	wire _w24483_ ;
	wire _w24484_ ;
	wire _w24485_ ;
	wire _w24486_ ;
	wire _w24487_ ;
	wire _w24488_ ;
	wire _w24489_ ;
	wire _w24490_ ;
	wire _w24491_ ;
	wire _w24492_ ;
	wire _w24493_ ;
	wire _w24494_ ;
	wire _w24495_ ;
	wire _w24496_ ;
	wire _w24497_ ;
	wire _w24498_ ;
	wire _w24499_ ;
	wire _w24500_ ;
	wire _w24501_ ;
	wire _w24502_ ;
	wire _w24503_ ;
	wire _w24504_ ;
	wire _w24505_ ;
	wire _w24506_ ;
	wire _w24507_ ;
	wire _w24508_ ;
	wire _w24509_ ;
	wire _w24510_ ;
	wire _w24511_ ;
	wire _w24512_ ;
	wire _w24513_ ;
	wire _w24514_ ;
	wire _w24515_ ;
	wire _w24516_ ;
	wire _w24517_ ;
	wire _w24518_ ;
	wire _w24519_ ;
	wire _w24520_ ;
	wire _w24521_ ;
	wire _w24522_ ;
	wire _w24523_ ;
	wire _w24524_ ;
	wire _w24525_ ;
	wire _w24526_ ;
	wire _w24527_ ;
	wire _w24528_ ;
	wire _w24529_ ;
	wire _w24530_ ;
	wire _w24531_ ;
	wire _w24532_ ;
	wire _w24533_ ;
	wire _w24534_ ;
	wire _w24535_ ;
	wire _w24536_ ;
	wire _w24537_ ;
	wire _w24538_ ;
	wire _w24539_ ;
	wire _w24540_ ;
	wire _w24541_ ;
	wire _w24542_ ;
	wire _w24543_ ;
	wire _w24544_ ;
	wire _w24545_ ;
	wire _w24546_ ;
	wire _w24547_ ;
	wire _w24548_ ;
	wire _w24549_ ;
	wire _w24550_ ;
	wire _w24551_ ;
	wire _w24552_ ;
	wire _w24553_ ;
	wire _w24554_ ;
	wire _w24555_ ;
	wire _w24556_ ;
	wire _w24557_ ;
	wire _w24558_ ;
	wire _w24559_ ;
	wire _w24560_ ;
	wire _w24561_ ;
	wire _w24562_ ;
	wire _w24563_ ;
	wire _w24564_ ;
	wire _w24565_ ;
	wire _w24566_ ;
	wire _w24567_ ;
	wire _w24568_ ;
	wire _w24569_ ;
	wire _w24570_ ;
	wire _w24571_ ;
	wire _w24572_ ;
	wire _w24573_ ;
	wire _w24574_ ;
	wire _w24575_ ;
	wire _w24576_ ;
	wire _w24577_ ;
	wire _w24578_ ;
	wire _w24579_ ;
	wire _w24580_ ;
	wire _w24581_ ;
	wire _w24582_ ;
	wire _w24583_ ;
	wire _w24584_ ;
	wire _w24585_ ;
	wire _w24586_ ;
	wire _w24587_ ;
	wire _w24588_ ;
	wire _w24589_ ;
	wire _w24590_ ;
	wire _w24591_ ;
	wire _w24592_ ;
	wire _w24593_ ;
	wire _w24594_ ;
	wire _w24595_ ;
	wire _w24596_ ;
	wire _w24597_ ;
	wire _w24598_ ;
	wire _w24599_ ;
	wire _w24600_ ;
	wire _w24601_ ;
	wire _w24602_ ;
	wire _w24603_ ;
	wire _w24604_ ;
	wire _w24605_ ;
	wire _w24606_ ;
	wire _w24607_ ;
	wire _w24608_ ;
	wire _w24609_ ;
	wire _w24610_ ;
	wire _w24611_ ;
	wire _w24612_ ;
	wire _w24613_ ;
	wire _w24614_ ;
	wire _w24615_ ;
	wire _w24616_ ;
	wire _w24617_ ;
	wire _w24618_ ;
	wire _w24619_ ;
	wire _w24620_ ;
	wire _w24621_ ;
	wire _w24622_ ;
	wire _w24623_ ;
	wire _w24624_ ;
	wire _w24625_ ;
	wire _w24626_ ;
	wire _w24627_ ;
	wire _w24628_ ;
	wire _w24629_ ;
	wire _w24630_ ;
	wire _w24631_ ;
	wire _w24632_ ;
	wire _w24633_ ;
	wire _w24634_ ;
	wire _w24635_ ;
	wire _w24636_ ;
	wire _w24637_ ;
	wire _w24638_ ;
	wire _w24639_ ;
	wire _w24640_ ;
	wire _w24641_ ;
	wire _w24642_ ;
	wire _w24643_ ;
	wire _w24644_ ;
	wire _w24645_ ;
	wire _w24646_ ;
	wire _w24647_ ;
	wire _w24648_ ;
	wire _w24649_ ;
	wire _w24650_ ;
	wire _w24651_ ;
	wire _w24652_ ;
	wire _w24653_ ;
	wire _w24654_ ;
	wire _w24655_ ;
	wire _w24656_ ;
	wire _w24657_ ;
	wire _w24658_ ;
	wire _w24659_ ;
	wire _w24660_ ;
	wire _w24661_ ;
	wire _w24662_ ;
	wire _w24663_ ;
	wire _w24664_ ;
	wire _w24665_ ;
	wire _w24666_ ;
	wire _w24667_ ;
	wire _w24668_ ;
	wire _w24669_ ;
	wire _w24670_ ;
	wire _w24671_ ;
	wire _w24672_ ;
	wire _w24673_ ;
	wire _w24674_ ;
	wire _w24675_ ;
	wire _w24676_ ;
	wire _w24677_ ;
	wire _w24678_ ;
	wire _w24679_ ;
	wire _w24680_ ;
	wire _w24681_ ;
	wire _w24682_ ;
	wire _w24683_ ;
	wire _w24684_ ;
	wire _w24685_ ;
	wire _w24686_ ;
	wire _w24687_ ;
	wire _w24688_ ;
	wire _w24689_ ;
	wire _w24690_ ;
	wire _w24691_ ;
	wire _w24692_ ;
	wire _w24693_ ;
	wire _w24694_ ;
	wire _w24695_ ;
	wire _w24696_ ;
	wire _w24697_ ;
	wire _w24698_ ;
	wire _w24699_ ;
	wire _w24700_ ;
	wire _w24701_ ;
	wire _w24702_ ;
	wire _w24703_ ;
	wire _w24704_ ;
	wire _w24705_ ;
	wire _w24706_ ;
	wire _w24707_ ;
	wire _w24708_ ;
	wire _w24709_ ;
	wire _w24710_ ;
	wire _w24711_ ;
	wire _w24712_ ;
	wire _w24713_ ;
	wire _w24714_ ;
	wire _w24715_ ;
	wire _w24716_ ;
	wire _w24717_ ;
	wire _w24718_ ;
	wire _w24719_ ;
	wire _w24720_ ;
	wire _w24721_ ;
	wire _w24722_ ;
	wire _w24723_ ;
	wire _w24724_ ;
	wire _w24725_ ;
	wire _w24726_ ;
	wire _w24727_ ;
	wire _w24728_ ;
	wire _w24729_ ;
	wire _w24730_ ;
	wire _w24731_ ;
	wire _w24732_ ;
	wire _w24733_ ;
	wire _w24734_ ;
	wire _w24735_ ;
	wire _w24736_ ;
	wire _w24737_ ;
	wire _w24738_ ;
	wire _w24739_ ;
	wire _w24740_ ;
	wire _w24741_ ;
	wire _w24742_ ;
	wire _w24743_ ;
	wire _w24744_ ;
	wire _w24745_ ;
	wire _w24746_ ;
	wire _w24747_ ;
	wire _w24748_ ;
	wire _w24749_ ;
	wire _w24750_ ;
	wire _w24751_ ;
	wire _w24752_ ;
	wire _w24753_ ;
	wire _w24754_ ;
	wire _w24755_ ;
	wire _w24756_ ;
	wire _w24757_ ;
	wire _w24758_ ;
	wire _w24759_ ;
	wire _w24760_ ;
	wire _w24761_ ;
	wire _w24762_ ;
	wire _w24763_ ;
	wire _w24764_ ;
	wire _w24765_ ;
	wire _w24766_ ;
	wire _w24767_ ;
	wire _w24768_ ;
	wire _w24769_ ;
	wire _w24770_ ;
	wire _w24771_ ;
	wire _w24772_ ;
	wire _w24773_ ;
	wire _w24774_ ;
	wire _w24775_ ;
	wire _w24776_ ;
	wire _w24777_ ;
	wire _w24778_ ;
	wire _w24779_ ;
	wire _w24780_ ;
	wire _w24781_ ;
	wire _w24782_ ;
	wire _w24783_ ;
	wire _w24784_ ;
	wire _w24785_ ;
	wire _w24786_ ;
	wire _w24787_ ;
	wire _w24788_ ;
	wire _w24789_ ;
	wire _w24790_ ;
	wire _w24791_ ;
	wire _w24792_ ;
	wire _w24793_ ;
	wire _w24794_ ;
	wire _w24795_ ;
	wire _w24796_ ;
	wire _w24797_ ;
	wire _w24798_ ;
	wire _w24799_ ;
	wire _w24800_ ;
	wire _w24801_ ;
	wire _w24802_ ;
	wire _w24803_ ;
	wire _w24804_ ;
	wire _w24805_ ;
	wire _w24806_ ;
	wire _w24807_ ;
	wire _w24808_ ;
	wire _w24809_ ;
	wire _w24810_ ;
	wire _w24811_ ;
	wire _w24812_ ;
	wire _w24813_ ;
	wire _w24814_ ;
	wire _w24815_ ;
	wire _w24816_ ;
	wire _w24817_ ;
	wire _w24818_ ;
	wire _w24819_ ;
	wire _w24820_ ;
	wire _w24821_ ;
	wire _w24822_ ;
	wire _w24823_ ;
	wire _w24824_ ;
	wire _w24825_ ;
	wire _w24826_ ;
	wire _w24827_ ;
	wire _w24828_ ;
	wire _w24829_ ;
	wire _w24830_ ;
	wire _w24831_ ;
	wire _w24832_ ;
	wire _w24833_ ;
	wire _w24834_ ;
	wire _w24835_ ;
	wire _w24836_ ;
	wire _w24837_ ;
	wire _w24838_ ;
	wire _w24839_ ;
	wire _w24840_ ;
	wire _w24841_ ;
	wire _w24842_ ;
	wire _w24843_ ;
	wire _w24844_ ;
	wire _w24845_ ;
	wire _w24846_ ;
	wire _w24847_ ;
	wire _w24848_ ;
	wire _w24849_ ;
	wire _w24850_ ;
	wire _w24851_ ;
	wire _w24852_ ;
	wire _w24853_ ;
	wire _w24854_ ;
	wire _w24855_ ;
	wire _w24856_ ;
	wire _w24857_ ;
	wire _w24858_ ;
	wire _w24859_ ;
	wire _w24860_ ;
	wire _w24861_ ;
	wire _w24862_ ;
	wire _w24863_ ;
	wire _w24864_ ;
	wire _w24865_ ;
	wire _w24866_ ;
	wire _w24867_ ;
	wire _w24868_ ;
	wire _w24869_ ;
	wire _w24870_ ;
	wire _w24871_ ;
	wire _w24872_ ;
	wire _w24873_ ;
	wire _w24874_ ;
	wire _w24875_ ;
	wire _w24876_ ;
	wire _w24877_ ;
	wire _w24878_ ;
	wire _w24879_ ;
	wire _w24880_ ;
	wire _w24881_ ;
	wire _w24882_ ;
	wire _w24883_ ;
	wire _w24884_ ;
	wire _w24885_ ;
	wire _w24886_ ;
	wire _w24887_ ;
	wire _w24888_ ;
	wire _w24889_ ;
	wire _w24890_ ;
	wire _w24891_ ;
	wire _w24892_ ;
	wire _w24893_ ;
	wire _w24894_ ;
	wire _w24895_ ;
	wire _w24896_ ;
	wire _w24897_ ;
	wire _w24898_ ;
	wire _w24899_ ;
	wire _w24900_ ;
	wire _w24901_ ;
	wire _w24902_ ;
	wire _w24903_ ;
	wire _w24904_ ;
	wire _w24905_ ;
	wire _w24906_ ;
	wire _w24907_ ;
	wire _w24908_ ;
	wire _w24909_ ;
	wire _w24910_ ;
	wire _w24911_ ;
	wire _w24912_ ;
	wire _w24913_ ;
	wire _w24914_ ;
	wire _w24915_ ;
	wire _w24916_ ;
	wire _w24917_ ;
	wire _w24918_ ;
	wire _w24919_ ;
	wire _w24920_ ;
	wire _w24921_ ;
	wire _w24922_ ;
	wire _w24923_ ;
	wire _w24924_ ;
	wire _w24925_ ;
	wire _w24926_ ;
	wire _w24927_ ;
	wire _w24928_ ;
	wire _w24929_ ;
	wire _w24930_ ;
	wire _w24931_ ;
	wire _w24932_ ;
	wire _w24933_ ;
	wire _w24934_ ;
	wire _w24935_ ;
	wire _w24936_ ;
	wire _w24937_ ;
	wire _w24938_ ;
	wire _w24939_ ;
	wire _w24940_ ;
	wire _w24941_ ;
	wire _w24942_ ;
	wire _w24943_ ;
	wire _w24944_ ;
	wire _w24945_ ;
	wire _w24946_ ;
	wire _w24947_ ;
	wire _w24948_ ;
	wire _w24949_ ;
	wire _w24950_ ;
	wire _w24951_ ;
	wire _w24952_ ;
	wire _w24953_ ;
	wire _w24954_ ;
	wire _w24955_ ;
	wire _w24956_ ;
	wire _w24957_ ;
	wire _w24958_ ;
	wire _w24959_ ;
	wire _w24960_ ;
	wire _w24961_ ;
	wire _w24962_ ;
	wire _w24963_ ;
	wire _w24964_ ;
	wire _w24965_ ;
	wire _w24966_ ;
	wire _w24967_ ;
	wire _w24968_ ;
	wire _w24969_ ;
	wire _w24970_ ;
	wire _w24971_ ;
	wire _w24972_ ;
	wire _w24973_ ;
	wire _w24974_ ;
	wire _w24975_ ;
	wire _w24976_ ;
	wire _w24977_ ;
	wire _w24978_ ;
	wire _w24979_ ;
	wire _w24980_ ;
	wire _w24981_ ;
	wire _w24982_ ;
	wire _w24983_ ;
	wire _w24984_ ;
	wire _w24985_ ;
	wire _w24986_ ;
	wire _w24987_ ;
	wire _w24988_ ;
	wire _w24989_ ;
	wire _w24990_ ;
	wire _w24991_ ;
	wire _w24992_ ;
	wire _w24993_ ;
	wire _w24994_ ;
	wire _w24995_ ;
	wire _w24996_ ;
	wire _w24997_ ;
	wire _w24998_ ;
	wire _w24999_ ;
	wire _w25000_ ;
	wire _w25001_ ;
	wire _w25002_ ;
	wire _w25003_ ;
	wire _w25004_ ;
	wire _w25005_ ;
	wire _w25006_ ;
	wire _w25007_ ;
	wire _w25008_ ;
	wire _w25009_ ;
	wire _w25010_ ;
	wire _w25011_ ;
	wire _w25012_ ;
	wire _w25013_ ;
	wire _w25014_ ;
	wire _w25015_ ;
	wire _w25016_ ;
	wire _w25017_ ;
	wire _w25018_ ;
	wire _w25019_ ;
	wire _w25020_ ;
	wire _w25021_ ;
	wire _w25022_ ;
	wire _w25023_ ;
	wire _w25024_ ;
	wire _w25025_ ;
	wire _w25026_ ;
	wire _w25027_ ;
	wire _w25028_ ;
	wire _w25029_ ;
	wire _w25030_ ;
	wire _w25031_ ;
	wire _w25032_ ;
	wire _w25033_ ;
	wire _w25034_ ;
	wire _w25035_ ;
	wire _w25036_ ;
	wire _w25037_ ;
	wire _w25038_ ;
	wire _w25039_ ;
	wire _w25040_ ;
	wire _w25041_ ;
	wire _w25042_ ;
	wire _w25043_ ;
	wire _w25044_ ;
	wire _w25045_ ;
	wire _w25046_ ;
	wire _w25047_ ;
	wire _w25048_ ;
	wire _w25049_ ;
	wire _w25050_ ;
	wire _w25051_ ;
	wire _w25052_ ;
	wire _w25053_ ;
	wire _w25054_ ;
	wire _w25055_ ;
	wire _w25056_ ;
	wire _w25057_ ;
	wire _w25058_ ;
	wire _w25059_ ;
	wire _w25060_ ;
	wire _w25061_ ;
	wire _w25062_ ;
	wire _w25063_ ;
	wire _w25064_ ;
	wire _w25065_ ;
	wire _w25066_ ;
	wire _w25067_ ;
	wire _w25068_ ;
	wire _w25069_ ;
	wire _w25070_ ;
	wire _w25071_ ;
	wire _w25072_ ;
	wire _w25073_ ;
	wire _w25074_ ;
	wire _w25075_ ;
	wire _w25076_ ;
	wire _w25077_ ;
	wire _w25078_ ;
	wire _w25079_ ;
	wire _w25080_ ;
	wire _w25081_ ;
	wire _w25082_ ;
	wire _w25083_ ;
	wire _w25084_ ;
	wire _w25085_ ;
	wire _w25086_ ;
	wire _w25087_ ;
	wire _w25088_ ;
	wire _w25089_ ;
	wire _w25090_ ;
	wire _w25091_ ;
	wire _w25092_ ;
	wire _w25093_ ;
	wire _w25094_ ;
	wire _w25095_ ;
	wire _w25096_ ;
	wire _w25097_ ;
	wire _w25098_ ;
	wire _w25099_ ;
	wire _w25100_ ;
	wire _w25101_ ;
	wire _w25102_ ;
	wire _w25103_ ;
	wire _w25104_ ;
	wire _w25105_ ;
	wire _w25106_ ;
	wire _w25107_ ;
	wire _w25108_ ;
	wire _w25109_ ;
	wire _w25110_ ;
	wire _w25111_ ;
	wire _w25112_ ;
	wire _w25113_ ;
	wire _w25114_ ;
	wire _w25115_ ;
	wire _w25116_ ;
	wire _w25117_ ;
	wire _w25118_ ;
	wire _w25119_ ;
	wire _w25120_ ;
	wire _w25121_ ;
	wire _w25122_ ;
	wire _w25123_ ;
	wire _w25124_ ;
	wire _w25125_ ;
	wire _w25126_ ;
	wire _w25127_ ;
	wire _w25128_ ;
	wire _w25129_ ;
	wire _w25130_ ;
	wire _w25131_ ;
	wire _w25132_ ;
	wire _w25133_ ;
	wire _w25134_ ;
	wire _w25135_ ;
	wire _w25136_ ;
	wire _w25137_ ;
	wire _w25138_ ;
	wire _w25139_ ;
	wire _w25140_ ;
	wire _w25141_ ;
	wire _w25142_ ;
	wire _w25143_ ;
	wire _w25144_ ;
	wire _w25145_ ;
	wire _w25146_ ;
	wire _w25147_ ;
	wire _w25148_ ;
	wire _w25149_ ;
	wire _w25150_ ;
	wire _w25151_ ;
	wire _w25152_ ;
	wire _w25153_ ;
	wire _w25154_ ;
	wire _w25155_ ;
	wire _w25156_ ;
	wire _w25157_ ;
	wire _w25158_ ;
	wire _w25159_ ;
	wire _w25160_ ;
	wire _w25161_ ;
	wire _w25162_ ;
	wire _w25163_ ;
	wire _w25164_ ;
	wire _w25165_ ;
	wire _w25166_ ;
	wire _w25167_ ;
	wire _w25168_ ;
	wire _w25169_ ;
	wire _w25170_ ;
	wire _w25171_ ;
	wire _w25172_ ;
	wire _w25173_ ;
	wire _w25174_ ;
	wire _w25175_ ;
	wire _w25176_ ;
	wire _w25177_ ;
	wire _w25178_ ;
	wire _w25179_ ;
	wire _w25180_ ;
	wire _w25181_ ;
	wire _w25182_ ;
	wire _w25183_ ;
	wire _w25184_ ;
	wire _w25185_ ;
	wire _w25186_ ;
	wire _w25187_ ;
	wire _w25188_ ;
	wire _w25189_ ;
	wire _w25190_ ;
	wire _w25191_ ;
	wire _w25192_ ;
	wire _w25193_ ;
	wire _w25194_ ;
	wire _w25195_ ;
	wire _w25196_ ;
	wire _w25197_ ;
	wire _w25198_ ;
	wire _w25199_ ;
	wire _w25200_ ;
	wire _w25201_ ;
	wire _w25202_ ;
	wire _w25203_ ;
	wire _w25204_ ;
	wire _w25205_ ;
	wire _w25206_ ;
	wire _w25207_ ;
	wire _w25208_ ;
	wire _w25209_ ;
	wire _w25210_ ;
	wire _w25211_ ;
	wire _w25212_ ;
	wire _w25213_ ;
	wire _w25214_ ;
	wire _w25215_ ;
	wire _w25216_ ;
	wire _w25217_ ;
	wire _w25218_ ;
	wire _w25219_ ;
	wire _w25220_ ;
	wire _w25221_ ;
	wire _w25222_ ;
	wire _w25223_ ;
	wire _w25224_ ;
	wire _w25225_ ;
	wire _w25226_ ;
	wire _w25227_ ;
	wire _w25228_ ;
	wire _w25229_ ;
	wire _w25230_ ;
	wire _w25231_ ;
	wire _w25232_ ;
	wire _w25233_ ;
	wire _w25234_ ;
	wire _w25235_ ;
	wire _w25236_ ;
	wire _w25237_ ;
	wire _w25238_ ;
	wire _w25239_ ;
	wire _w25240_ ;
	wire _w25241_ ;
	wire _w25242_ ;
	wire _w25243_ ;
	wire _w25244_ ;
	wire _w25245_ ;
	wire _w25246_ ;
	wire _w25247_ ;
	wire _w25248_ ;
	wire _w25249_ ;
	wire _w25250_ ;
	wire _w25251_ ;
	wire _w25252_ ;
	wire _w25253_ ;
	wire _w25254_ ;
	wire _w25255_ ;
	wire _w25256_ ;
	wire _w25257_ ;
	wire _w25258_ ;
	wire _w25259_ ;
	wire _w25260_ ;
	wire _w25261_ ;
	wire _w25262_ ;
	wire _w25263_ ;
	wire _w25264_ ;
	wire _w25265_ ;
	wire _w25266_ ;
	wire _w25267_ ;
	wire _w25268_ ;
	wire _w25269_ ;
	wire _w25270_ ;
	wire _w25271_ ;
	wire _w25272_ ;
	wire _w25273_ ;
	wire _w25274_ ;
	wire _w25275_ ;
	wire _w25276_ ;
	wire _w25277_ ;
	wire _w25278_ ;
	wire _w25279_ ;
	wire _w25280_ ;
	wire _w25281_ ;
	wire _w25282_ ;
	wire _w25283_ ;
	wire _w25284_ ;
	wire _w25285_ ;
	wire _w25286_ ;
	wire _w25287_ ;
	wire _w25288_ ;
	wire _w25289_ ;
	wire _w25290_ ;
	wire _w25291_ ;
	wire _w25292_ ;
	wire _w25293_ ;
	wire _w25294_ ;
	wire _w25295_ ;
	wire _w25296_ ;
	wire _w25297_ ;
	wire _w25298_ ;
	wire _w25299_ ;
	wire _w25300_ ;
	wire _w25301_ ;
	wire _w25302_ ;
	wire _w25303_ ;
	wire _w25304_ ;
	wire _w25305_ ;
	wire _w25306_ ;
	wire _w25307_ ;
	wire _w25308_ ;
	wire _w25309_ ;
	wire _w25310_ ;
	wire _w25311_ ;
	wire _w25312_ ;
	wire _w25313_ ;
	wire _w25314_ ;
	wire _w25315_ ;
	wire _w25316_ ;
	wire _w25317_ ;
	wire _w25318_ ;
	wire _w25319_ ;
	wire _w25320_ ;
	wire _w25321_ ;
	wire _w25322_ ;
	wire _w25323_ ;
	wire _w25324_ ;
	wire _w25325_ ;
	wire _w25326_ ;
	wire _w25327_ ;
	wire _w25328_ ;
	wire _w25329_ ;
	wire _w25330_ ;
	wire _w25331_ ;
	wire _w25332_ ;
	wire _w25333_ ;
	wire _w25334_ ;
	wire _w25335_ ;
	wire _w25336_ ;
	wire _w25337_ ;
	wire _w25338_ ;
	wire _w25339_ ;
	wire _w25340_ ;
	wire _w25341_ ;
	wire _w25342_ ;
	wire _w25343_ ;
	wire _w25344_ ;
	wire _w25345_ ;
	wire _w25346_ ;
	wire _w25347_ ;
	wire _w25348_ ;
	wire _w25349_ ;
	wire _w25350_ ;
	wire _w25351_ ;
	wire _w25352_ ;
	wire _w25353_ ;
	wire _w25354_ ;
	wire _w25355_ ;
	wire _w25356_ ;
	wire _w25357_ ;
	wire _w25358_ ;
	wire _w25359_ ;
	wire _w25360_ ;
	wire _w25361_ ;
	wire _w25362_ ;
	wire _w25363_ ;
	wire _w25364_ ;
	wire _w25365_ ;
	wire _w25366_ ;
	wire _w25367_ ;
	wire _w25368_ ;
	wire _w25369_ ;
	wire _w25370_ ;
	wire _w25371_ ;
	wire _w25372_ ;
	wire _w25373_ ;
	wire _w25374_ ;
	wire _w25375_ ;
	wire _w25376_ ;
	wire _w25377_ ;
	wire _w25378_ ;
	wire _w25379_ ;
	wire _w25380_ ;
	wire _w25381_ ;
	wire _w25382_ ;
	wire _w25383_ ;
	wire _w25384_ ;
	wire _w25385_ ;
	wire _w25386_ ;
	wire _w25387_ ;
	wire _w25388_ ;
	wire _w25389_ ;
	wire _w25390_ ;
	wire _w25391_ ;
	wire _w25392_ ;
	wire _w25393_ ;
	wire _w25394_ ;
	wire _w25395_ ;
	wire _w25396_ ;
	wire _w25397_ ;
	wire _w25398_ ;
	wire _w25399_ ;
	wire _w25400_ ;
	wire _w25401_ ;
	wire _w25402_ ;
	wire _w25403_ ;
	wire _w25404_ ;
	wire _w25405_ ;
	wire _w25406_ ;
	wire _w25407_ ;
	wire _w25408_ ;
	wire _w25409_ ;
	wire _w25410_ ;
	wire _w25411_ ;
	wire _w25412_ ;
	wire _w25413_ ;
	wire _w25414_ ;
	wire _w25415_ ;
	wire _w25416_ ;
	wire _w25417_ ;
	wire _w25418_ ;
	wire _w25419_ ;
	wire _w25420_ ;
	wire _w25421_ ;
	wire _w25422_ ;
	wire _w25423_ ;
	wire _w25424_ ;
	wire _w25425_ ;
	wire _w25426_ ;
	wire _w25427_ ;
	wire _w25428_ ;
	wire _w25429_ ;
	wire _w25430_ ;
	wire _w25431_ ;
	wire _w25432_ ;
	wire _w25433_ ;
	wire _w25434_ ;
	wire _w25435_ ;
	wire _w25436_ ;
	wire _w25437_ ;
	wire _w25438_ ;
	wire _w25439_ ;
	wire _w25440_ ;
	wire _w25441_ ;
	wire _w25442_ ;
	wire _w25443_ ;
	wire _w25444_ ;
	wire _w25445_ ;
	wire _w25446_ ;
	wire _w25447_ ;
	wire _w25448_ ;
	wire _w25449_ ;
	wire _w25450_ ;
	wire _w25451_ ;
	wire _w25452_ ;
	wire _w25453_ ;
	wire _w25454_ ;
	wire _w25455_ ;
	wire _w25456_ ;
	wire _w25457_ ;
	wire _w25458_ ;
	wire _w25459_ ;
	wire _w25460_ ;
	wire _w25461_ ;
	wire _w25462_ ;
	wire _w25463_ ;
	wire _w25464_ ;
	wire _w25465_ ;
	wire _w25466_ ;
	wire _w25467_ ;
	wire _w25468_ ;
	wire _w25469_ ;
	wire _w25470_ ;
	wire _w25471_ ;
	wire _w25472_ ;
	wire _w25473_ ;
	wire _w25474_ ;
	wire _w25475_ ;
	wire _w25476_ ;
	wire _w25477_ ;
	wire _w25478_ ;
	wire _w25479_ ;
	wire _w25480_ ;
	wire _w25481_ ;
	wire _w25482_ ;
	wire _w25483_ ;
	wire _w25484_ ;
	wire _w25485_ ;
	wire _w25486_ ;
	wire _w25487_ ;
	wire _w25488_ ;
	wire _w25489_ ;
	wire _w25490_ ;
	wire _w25491_ ;
	wire _w25492_ ;
	wire _w25493_ ;
	wire _w25494_ ;
	wire _w25495_ ;
	wire _w25496_ ;
	wire _w25497_ ;
	wire _w25498_ ;
	wire _w25499_ ;
	wire _w25500_ ;
	wire _w25501_ ;
	wire _w25502_ ;
	wire _w25503_ ;
	wire _w25504_ ;
	wire _w25505_ ;
	wire _w25506_ ;
	wire _w25507_ ;
	wire _w25508_ ;
	wire _w25509_ ;
	wire _w25510_ ;
	wire _w25511_ ;
	wire _w25512_ ;
	wire _w25513_ ;
	wire _w25514_ ;
	wire _w25515_ ;
	wire _w25516_ ;
	wire _w25517_ ;
	wire _w25518_ ;
	wire _w25519_ ;
	wire _w25520_ ;
	wire _w25521_ ;
	wire _w25522_ ;
	wire _w25523_ ;
	wire _w25524_ ;
	wire _w25525_ ;
	wire _w25526_ ;
	wire _w25527_ ;
	wire _w25528_ ;
	wire _w25529_ ;
	wire _w25530_ ;
	wire _w25531_ ;
	wire _w25532_ ;
	wire _w25533_ ;
	wire _w25534_ ;
	wire _w25535_ ;
	wire _w25536_ ;
	wire _w25537_ ;
	wire _w25538_ ;
	wire _w25539_ ;
	wire _w25540_ ;
	wire _w25541_ ;
	wire _w25542_ ;
	wire _w25543_ ;
	wire _w25544_ ;
	wire _w25545_ ;
	wire _w25546_ ;
	wire _w25547_ ;
	wire _w25548_ ;
	wire _w25549_ ;
	wire _w25550_ ;
	wire _w25551_ ;
	wire _w25552_ ;
	wire _w25553_ ;
	wire _w25554_ ;
	wire _w25555_ ;
	wire _w25556_ ;
	wire _w25557_ ;
	wire _w25558_ ;
	wire _w25559_ ;
	wire _w25560_ ;
	wire _w25561_ ;
	wire _w25562_ ;
	wire _w25563_ ;
	wire _w25564_ ;
	wire _w25565_ ;
	wire _w25566_ ;
	wire _w25567_ ;
	wire _w25568_ ;
	wire _w25569_ ;
	wire _w25570_ ;
	wire _w25571_ ;
	wire _w25572_ ;
	wire _w25573_ ;
	wire _w25574_ ;
	wire _w25575_ ;
	wire _w25576_ ;
	wire _w25577_ ;
	wire _w25578_ ;
	wire _w25579_ ;
	wire _w25580_ ;
	wire _w25581_ ;
	wire _w25582_ ;
	wire _w25583_ ;
	wire _w25584_ ;
	wire _w25585_ ;
	wire _w25586_ ;
	wire _w25587_ ;
	wire _w25588_ ;
	wire _w25589_ ;
	wire _w25590_ ;
	wire _w25591_ ;
	wire _w25592_ ;
	wire _w25593_ ;
	wire _w25594_ ;
	wire _w25595_ ;
	wire _w25596_ ;
	wire _w25597_ ;
	wire _w25598_ ;
	wire _w25599_ ;
	wire _w25600_ ;
	wire _w25601_ ;
	wire _w25602_ ;
	wire _w25603_ ;
	wire _w25604_ ;
	wire _w25605_ ;
	wire _w25606_ ;
	wire _w25607_ ;
	wire _w25608_ ;
	wire _w25609_ ;
	wire _w25610_ ;
	wire _w25611_ ;
	wire _w25612_ ;
	wire _w25613_ ;
	wire _w25614_ ;
	wire _w25615_ ;
	wire _w25616_ ;
	wire _w25617_ ;
	wire _w25618_ ;
	wire _w25619_ ;
	wire _w25620_ ;
	wire _w25621_ ;
	wire _w25622_ ;
	wire _w25623_ ;
	wire _w25624_ ;
	wire _w25625_ ;
	wire _w25626_ ;
	wire _w25627_ ;
	wire _w25628_ ;
	wire _w25629_ ;
	wire _w25630_ ;
	wire _w25631_ ;
	wire _w25632_ ;
	wire _w25633_ ;
	wire _w25634_ ;
	wire _w25635_ ;
	wire _w25636_ ;
	wire _w25637_ ;
	wire _w25638_ ;
	wire _w25639_ ;
	wire _w25640_ ;
	wire _w25641_ ;
	wire _w25642_ ;
	wire _w25643_ ;
	wire _w25644_ ;
	wire _w25645_ ;
	wire _w25646_ ;
	wire _w25647_ ;
	wire _w25648_ ;
	wire _w25649_ ;
	wire _w25650_ ;
	wire _w25651_ ;
	wire _w25652_ ;
	wire _w25653_ ;
	wire _w25654_ ;
	wire _w25655_ ;
	wire _w25656_ ;
	wire _w25657_ ;
	wire _w25658_ ;
	wire _w25659_ ;
	wire _w25660_ ;
	wire _w25661_ ;
	wire _w25662_ ;
	wire _w25663_ ;
	wire _w25664_ ;
	wire _w25665_ ;
	wire _w25666_ ;
	wire _w25667_ ;
	wire _w25668_ ;
	wire _w25669_ ;
	wire _w25670_ ;
	wire _w25671_ ;
	wire _w25672_ ;
	wire _w25673_ ;
	wire _w25674_ ;
	wire _w25675_ ;
	wire _w25676_ ;
	wire _w25677_ ;
	wire _w25678_ ;
	wire _w25679_ ;
	wire _w25680_ ;
	wire _w25681_ ;
	wire _w25682_ ;
	wire _w25683_ ;
	wire _w25684_ ;
	wire _w25685_ ;
	wire _w25686_ ;
	wire _w25687_ ;
	wire _w25688_ ;
	wire _w25689_ ;
	wire _w25690_ ;
	wire _w25691_ ;
	wire _w25692_ ;
	wire _w25693_ ;
	wire _w25694_ ;
	wire _w25695_ ;
	wire _w25696_ ;
	wire _w25697_ ;
	wire _w25698_ ;
	wire _w25699_ ;
	wire _w25700_ ;
	wire _w25701_ ;
	wire _w25702_ ;
	wire _w25703_ ;
	wire _w25704_ ;
	wire _w25705_ ;
	wire _w25706_ ;
	wire _w25707_ ;
	wire _w25708_ ;
	wire _w25709_ ;
	wire _w25710_ ;
	wire _w25711_ ;
	wire _w25712_ ;
	wire _w25713_ ;
	wire _w25714_ ;
	wire _w25715_ ;
	wire _w25716_ ;
	wire _w25717_ ;
	wire _w25718_ ;
	wire _w25719_ ;
	wire _w25720_ ;
	wire _w25721_ ;
	wire _w25722_ ;
	wire _w25723_ ;
	wire _w25724_ ;
	wire _w25725_ ;
	wire _w25726_ ;
	wire _w25727_ ;
	wire _w25728_ ;
	wire _w25729_ ;
	wire _w25730_ ;
	wire _w25731_ ;
	wire _w25732_ ;
	wire _w25733_ ;
	wire _w25734_ ;
	wire _w25735_ ;
	wire _w25736_ ;
	wire _w25737_ ;
	wire _w25738_ ;
	wire _w25739_ ;
	wire _w25740_ ;
	wire _w25741_ ;
	wire _w25742_ ;
	wire _w25743_ ;
	wire _w25744_ ;
	wire _w25745_ ;
	wire _w25746_ ;
	wire _w25747_ ;
	wire _w25748_ ;
	wire _w25749_ ;
	wire _w25750_ ;
	wire _w25751_ ;
	wire _w25752_ ;
	wire _w25753_ ;
	wire _w25754_ ;
	wire _w25755_ ;
	wire _w25756_ ;
	wire _w25757_ ;
	wire _w25758_ ;
	wire _w25759_ ;
	wire _w25760_ ;
	wire _w25761_ ;
	wire _w25762_ ;
	wire _w25763_ ;
	wire _w25764_ ;
	wire _w25765_ ;
	wire _w25766_ ;
	wire _w25767_ ;
	wire _w25768_ ;
	wire _w25769_ ;
	wire _w25770_ ;
	wire _w25771_ ;
	wire _w25772_ ;
	wire _w25773_ ;
	wire _w25774_ ;
	wire _w25775_ ;
	wire _w25776_ ;
	wire _w25777_ ;
	wire _w25778_ ;
	wire _w25779_ ;
	wire _w25780_ ;
	wire _w25781_ ;
	wire _w25782_ ;
	wire _w25783_ ;
	wire _w25784_ ;
	wire _w25785_ ;
	wire _w25786_ ;
	wire _w25787_ ;
	wire _w25788_ ;
	wire _w25789_ ;
	wire _w25790_ ;
	wire _w25791_ ;
	wire _w25792_ ;
	wire _w25793_ ;
	wire _w25794_ ;
	wire _w25795_ ;
	wire _w25796_ ;
	wire _w25797_ ;
	wire _w25798_ ;
	wire _w25799_ ;
	wire _w25800_ ;
	wire _w25801_ ;
	wire _w25802_ ;
	wire _w25803_ ;
	wire _w25804_ ;
	wire _w25805_ ;
	wire _w25806_ ;
	wire _w25807_ ;
	wire _w25808_ ;
	wire _w25809_ ;
	wire _w25810_ ;
	wire _w25811_ ;
	wire _w25812_ ;
	wire _w25813_ ;
	wire _w25814_ ;
	wire _w25815_ ;
	wire _w25816_ ;
	wire _w25817_ ;
	wire _w25818_ ;
	wire _w25819_ ;
	wire _w25820_ ;
	wire _w25821_ ;
	wire _w25822_ ;
	wire _w25823_ ;
	wire _w25824_ ;
	wire _w25825_ ;
	wire _w25826_ ;
	wire _w25827_ ;
	wire _w25828_ ;
	wire _w25829_ ;
	wire _w25830_ ;
	wire _w25831_ ;
	wire _w25832_ ;
	wire _w25833_ ;
	wire _w25834_ ;
	wire _w25835_ ;
	wire _w25836_ ;
	wire _w25837_ ;
	wire _w25838_ ;
	wire _w25839_ ;
	wire _w25840_ ;
	wire _w25841_ ;
	wire _w25842_ ;
	wire _w25843_ ;
	wire _w25844_ ;
	wire _w25845_ ;
	wire _w25846_ ;
	wire _w25847_ ;
	wire _w25848_ ;
	wire _w25849_ ;
	wire _w25850_ ;
	wire _w25851_ ;
	wire _w25852_ ;
	wire _w25853_ ;
	wire _w25854_ ;
	wire _w25855_ ;
	wire _w25856_ ;
	wire _w25857_ ;
	wire _w25858_ ;
	wire _w25859_ ;
	wire _w25860_ ;
	wire _w25861_ ;
	wire _w25862_ ;
	wire _w25863_ ;
	wire _w25864_ ;
	wire _w25865_ ;
	wire _w25866_ ;
	wire _w25867_ ;
	wire _w25868_ ;
	wire _w25869_ ;
	wire _w25870_ ;
	wire _w25871_ ;
	wire _w25872_ ;
	wire _w25873_ ;
	wire _w25874_ ;
	wire _w25875_ ;
	wire _w25876_ ;
	wire _w25877_ ;
	wire _w25878_ ;
	wire _w25879_ ;
	wire _w25880_ ;
	wire _w25881_ ;
	wire _w25882_ ;
	wire _w25883_ ;
	wire _w25884_ ;
	wire _w25885_ ;
	wire _w25886_ ;
	wire _w25887_ ;
	wire _w25888_ ;
	wire _w25889_ ;
	wire _w25890_ ;
	wire _w25891_ ;
	wire _w25892_ ;
	wire _w25893_ ;
	wire _w25894_ ;
	wire _w25895_ ;
	wire _w25896_ ;
	wire _w25897_ ;
	wire _w25898_ ;
	wire _w25899_ ;
	wire _w25900_ ;
	wire _w25901_ ;
	wire _w25902_ ;
	wire _w25903_ ;
	wire _w25904_ ;
	wire _w25905_ ;
	wire _w25906_ ;
	wire _w25907_ ;
	wire _w25908_ ;
	wire _w25909_ ;
	wire _w25910_ ;
	wire _w25911_ ;
	wire _w25912_ ;
	wire _w25913_ ;
	wire _w25914_ ;
	wire _w25915_ ;
	wire _w25916_ ;
	wire _w25917_ ;
	wire _w25918_ ;
	wire _w25919_ ;
	wire _w25920_ ;
	wire _w25921_ ;
	wire _w25922_ ;
	wire _w25923_ ;
	wire _w25924_ ;
	wire _w25925_ ;
	wire _w25926_ ;
	wire _w25927_ ;
	wire _w25928_ ;
	wire _w25929_ ;
	wire _w25930_ ;
	wire _w25931_ ;
	wire _w25932_ ;
	wire _w25933_ ;
	wire _w25934_ ;
	wire _w25935_ ;
	wire _w25936_ ;
	wire _w25937_ ;
	wire _w25938_ ;
	wire _w25939_ ;
	wire _w25940_ ;
	wire _w25941_ ;
	wire _w25942_ ;
	wire _w25943_ ;
	wire _w25944_ ;
	wire _w25945_ ;
	wire _w25946_ ;
	wire _w25947_ ;
	wire _w25948_ ;
	wire _w25949_ ;
	wire _w25950_ ;
	wire _w25951_ ;
	wire _w25952_ ;
	wire _w25953_ ;
	wire _w25954_ ;
	wire _w25955_ ;
	wire _w25956_ ;
	wire _w25957_ ;
	wire _w25958_ ;
	wire _w25959_ ;
	wire _w25960_ ;
	wire _w25961_ ;
	wire _w25962_ ;
	wire _w25963_ ;
	wire _w25964_ ;
	wire _w25965_ ;
	wire _w25966_ ;
	wire _w25967_ ;
	wire _w25968_ ;
	wire _w25969_ ;
	wire _w25970_ ;
	wire _w25971_ ;
	wire _w25972_ ;
	wire _w25973_ ;
	wire _w25974_ ;
	wire _w25975_ ;
	wire _w25976_ ;
	wire _w25977_ ;
	wire _w25978_ ;
	wire _w25979_ ;
	wire _w25980_ ;
	wire _w25981_ ;
	wire _w25982_ ;
	wire _w25983_ ;
	wire _w25984_ ;
	wire _w25985_ ;
	wire _w25986_ ;
	wire _w25987_ ;
	wire _w25988_ ;
	wire _w25989_ ;
	wire _w25990_ ;
	wire _w25991_ ;
	wire _w25992_ ;
	wire _w25993_ ;
	wire _w25994_ ;
	wire _w25995_ ;
	wire _w25996_ ;
	wire _w25997_ ;
	wire _w25998_ ;
	wire _w25999_ ;
	wire _w26000_ ;
	wire _w26001_ ;
	wire _w26002_ ;
	wire _w26003_ ;
	wire _w26004_ ;
	wire _w26005_ ;
	wire _w26006_ ;
	wire _w26007_ ;
	wire _w26008_ ;
	wire _w26009_ ;
	wire _w26010_ ;
	wire _w26011_ ;
	wire _w26012_ ;
	wire _w26013_ ;
	wire _w26014_ ;
	wire _w26015_ ;
	wire _w26016_ ;
	wire _w26017_ ;
	wire _w26018_ ;
	wire _w26019_ ;
	wire _w26020_ ;
	wire _w26021_ ;
	wire _w26022_ ;
	wire _w26023_ ;
	wire _w26024_ ;
	wire _w26025_ ;
	wire _w26026_ ;
	wire _w26027_ ;
	wire _w26028_ ;
	wire _w26029_ ;
	wire _w26030_ ;
	wire _w26031_ ;
	wire _w26032_ ;
	wire _w26033_ ;
	wire _w26034_ ;
	wire _w26035_ ;
	wire _w26036_ ;
	wire _w26037_ ;
	wire _w26038_ ;
	wire _w26039_ ;
	wire _w26040_ ;
	wire _w26041_ ;
	wire _w26042_ ;
	wire _w26043_ ;
	wire _w26044_ ;
	wire _w26045_ ;
	wire _w26046_ ;
	wire _w26047_ ;
	wire _w26048_ ;
	wire _w26049_ ;
	wire _w26050_ ;
	wire _w26051_ ;
	wire _w26052_ ;
	wire _w26053_ ;
	wire _w26054_ ;
	wire _w26055_ ;
	wire _w26056_ ;
	wire _w26057_ ;
	wire _w26058_ ;
	wire _w26059_ ;
	wire _w26060_ ;
	wire _w26061_ ;
	wire _w26062_ ;
	wire _w26063_ ;
	wire _w26064_ ;
	wire _w26065_ ;
	wire _w26066_ ;
	wire _w26067_ ;
	wire _w26068_ ;
	wire _w26069_ ;
	wire _w26070_ ;
	wire _w26071_ ;
	wire _w26072_ ;
	wire _w26073_ ;
	wire _w26074_ ;
	wire _w26075_ ;
	wire _w26076_ ;
	wire _w26077_ ;
	wire _w26078_ ;
	wire _w26079_ ;
	wire _w26080_ ;
	wire _w26081_ ;
	wire _w26082_ ;
	wire _w26083_ ;
	wire _w26084_ ;
	wire _w26085_ ;
	wire _w26086_ ;
	wire _w26087_ ;
	wire _w26088_ ;
	wire _w26089_ ;
	wire _w26090_ ;
	wire _w26091_ ;
	wire _w26092_ ;
	wire _w26093_ ;
	wire _w26094_ ;
	wire _w26095_ ;
	wire _w26096_ ;
	wire _w26097_ ;
	wire _w26098_ ;
	wire _w26099_ ;
	wire _w26100_ ;
	wire _w26101_ ;
	wire _w26102_ ;
	wire _w26103_ ;
	wire _w26104_ ;
	wire _w26105_ ;
	wire _w26106_ ;
	wire _w26107_ ;
	wire _w26108_ ;
	wire _w26109_ ;
	wire _w26110_ ;
	wire _w26111_ ;
	wire _w26112_ ;
	wire _w26113_ ;
	wire _w26114_ ;
	wire _w26115_ ;
	wire _w26116_ ;
	wire _w26117_ ;
	wire _w26118_ ;
	wire _w26119_ ;
	wire _w26120_ ;
	wire _w26121_ ;
	wire _w26122_ ;
	wire _w26123_ ;
	wire _w26124_ ;
	wire _w26125_ ;
	wire _w26126_ ;
	wire _w26127_ ;
	wire _w26128_ ;
	wire _w26129_ ;
	wire _w26130_ ;
	wire _w26131_ ;
	wire _w26132_ ;
	wire _w26133_ ;
	wire _w26134_ ;
	wire _w26135_ ;
	wire _w26136_ ;
	wire _w26137_ ;
	wire _w26138_ ;
	wire _w26139_ ;
	wire _w26140_ ;
	wire _w26141_ ;
	wire _w26142_ ;
	wire _w26143_ ;
	wire _w26144_ ;
	wire _w26145_ ;
	wire _w26146_ ;
	wire _w26147_ ;
	wire _w26148_ ;
	wire _w26149_ ;
	wire _w26150_ ;
	wire _w26151_ ;
	wire _w26152_ ;
	wire _w26153_ ;
	wire _w26154_ ;
	wire _w26155_ ;
	wire _w26156_ ;
	wire _w26157_ ;
	wire _w26158_ ;
	wire _w26159_ ;
	wire _w26160_ ;
	wire _w26161_ ;
	wire _w26162_ ;
	wire _w26163_ ;
	wire _w26164_ ;
	wire _w26165_ ;
	wire _w26166_ ;
	wire _w26167_ ;
	wire _w26168_ ;
	wire _w26169_ ;
	wire _w26170_ ;
	wire _w26171_ ;
	wire _w26172_ ;
	wire _w26173_ ;
	wire _w26174_ ;
	wire _w26175_ ;
	wire _w26176_ ;
	wire _w26177_ ;
	wire _w26178_ ;
	wire _w26179_ ;
	wire _w26180_ ;
	wire _w26181_ ;
	wire _w26182_ ;
	wire _w26183_ ;
	wire _w26184_ ;
	wire _w26185_ ;
	wire _w26186_ ;
	wire _w26187_ ;
	wire _w26188_ ;
	wire _w26189_ ;
	wire _w26190_ ;
	wire _w26191_ ;
	wire _w26192_ ;
	wire _w26193_ ;
	wire _w26194_ ;
	wire _w26195_ ;
	wire _w26196_ ;
	wire _w26197_ ;
	wire _w26198_ ;
	wire _w26199_ ;
	wire _w26200_ ;
	wire _w26201_ ;
	wire _w26202_ ;
	wire _w26203_ ;
	wire _w26204_ ;
	wire _w26205_ ;
	wire _w26206_ ;
	wire _w26207_ ;
	wire _w26208_ ;
	wire _w26209_ ;
	wire _w26210_ ;
	wire _w26211_ ;
	wire _w26212_ ;
	wire _w26213_ ;
	wire _w26214_ ;
	wire _w26215_ ;
	wire _w26216_ ;
	wire _w26217_ ;
	wire _w26218_ ;
	wire _w26219_ ;
	wire _w26220_ ;
	wire _w26221_ ;
	wire _w26222_ ;
	wire _w26223_ ;
	wire _w26224_ ;
	wire _w26225_ ;
	wire _w26226_ ;
	wire _w26227_ ;
	wire _w26228_ ;
	wire _w26229_ ;
	wire _w26230_ ;
	wire _w26231_ ;
	wire _w26232_ ;
	wire _w26233_ ;
	wire _w26234_ ;
	wire _w26235_ ;
	wire _w26236_ ;
	wire _w26237_ ;
	wire _w26238_ ;
	wire _w26239_ ;
	wire _w26240_ ;
	wire _w26241_ ;
	wire _w26242_ ;
	wire _w26243_ ;
	wire _w26244_ ;
	wire _w26245_ ;
	wire _w26246_ ;
	wire _w26247_ ;
	wire _w26248_ ;
	wire _w26249_ ;
	wire _w26250_ ;
	wire _w26251_ ;
	wire _w26252_ ;
	wire _w26253_ ;
	wire _w26254_ ;
	wire _w26255_ ;
	wire _w26256_ ;
	wire _w26257_ ;
	wire _w26258_ ;
	wire _w26259_ ;
	wire _w26260_ ;
	wire _w26261_ ;
	wire _w26262_ ;
	wire _w26263_ ;
	wire _w26264_ ;
	wire _w26265_ ;
	wire _w26266_ ;
	wire _w26267_ ;
	wire _w26268_ ;
	wire _w26269_ ;
	wire _w26270_ ;
	wire _w26271_ ;
	wire _w26272_ ;
	wire _w26273_ ;
	wire _w26274_ ;
	wire _w26275_ ;
	wire _w26276_ ;
	wire _w26277_ ;
	wire _w26278_ ;
	wire _w26279_ ;
	wire _w26280_ ;
	wire _w26281_ ;
	wire _w26282_ ;
	wire _w26283_ ;
	wire _w26284_ ;
	wire _w26285_ ;
	wire _w26286_ ;
	wire _w26287_ ;
	wire _w26288_ ;
	wire _w26289_ ;
	wire _w26290_ ;
	wire _w26291_ ;
	wire _w26292_ ;
	wire _w26293_ ;
	wire _w26294_ ;
	wire _w26295_ ;
	wire _w26296_ ;
	wire _w26297_ ;
	wire _w26298_ ;
	wire _w26299_ ;
	wire _w26300_ ;
	wire _w26301_ ;
	wire _w26302_ ;
	wire _w26303_ ;
	wire _w26304_ ;
	wire _w26305_ ;
	wire _w26306_ ;
	wire _w26307_ ;
	wire _w26308_ ;
	wire _w26309_ ;
	wire _w26310_ ;
	wire _w26311_ ;
	wire _w26312_ ;
	wire _w26313_ ;
	wire _w26314_ ;
	wire _w26315_ ;
	wire _w26316_ ;
	wire _w26317_ ;
	wire _w26318_ ;
	wire _w26319_ ;
	wire _w26320_ ;
	wire _w26321_ ;
	wire _w26322_ ;
	wire _w26323_ ;
	wire _w26324_ ;
	wire _w26325_ ;
	wire _w26326_ ;
	wire _w26327_ ;
	wire _w26328_ ;
	wire _w26329_ ;
	wire _w26330_ ;
	wire _w26331_ ;
	wire _w26332_ ;
	wire _w26333_ ;
	wire _w26334_ ;
	wire _w26335_ ;
	wire _w26336_ ;
	wire _w26337_ ;
	wire _w26338_ ;
	wire _w26339_ ;
	wire _w26340_ ;
	wire _w26341_ ;
	wire _w26342_ ;
	wire _w26343_ ;
	wire _w26344_ ;
	wire _w26345_ ;
	wire _w26346_ ;
	wire _w26347_ ;
	wire _w26348_ ;
	wire _w26349_ ;
	wire _w26350_ ;
	wire _w26351_ ;
	wire _w26352_ ;
	wire _w26353_ ;
	wire _w26354_ ;
	wire _w26355_ ;
	wire _w26356_ ;
	wire _w26357_ ;
	wire _w26358_ ;
	wire _w26359_ ;
	wire _w26360_ ;
	wire _w26361_ ;
	wire _w26362_ ;
	wire _w26363_ ;
	wire _w26364_ ;
	wire _w26365_ ;
	wire _w26366_ ;
	wire _w26367_ ;
	wire _w26368_ ;
	wire _w26369_ ;
	wire _w26370_ ;
	wire _w26371_ ;
	wire _w26372_ ;
	wire _w26373_ ;
	wire _w26374_ ;
	wire _w26375_ ;
	wire _w26376_ ;
	wire _w26377_ ;
	wire _w26378_ ;
	wire _w26379_ ;
	wire _w26380_ ;
	wire _w26381_ ;
	wire _w26382_ ;
	wire _w26383_ ;
	wire _w26384_ ;
	wire _w26385_ ;
	wire _w26386_ ;
	wire _w26387_ ;
	wire _w26388_ ;
	wire _w26389_ ;
	wire _w26390_ ;
	wire _w26391_ ;
	wire _w26392_ ;
	wire _w26393_ ;
	wire _w26394_ ;
	wire _w26395_ ;
	wire _w26396_ ;
	wire _w26397_ ;
	wire _w26398_ ;
	wire _w26399_ ;
	wire _w26400_ ;
	wire _w26401_ ;
	wire _w26402_ ;
	wire _w26403_ ;
	wire _w26404_ ;
	wire _w26405_ ;
	wire _w26406_ ;
	wire _w26407_ ;
	wire _w26408_ ;
	wire _w26409_ ;
	wire _w26410_ ;
	wire _w26411_ ;
	wire _w26412_ ;
	wire _w26413_ ;
	wire _w26414_ ;
	wire _w26415_ ;
	wire _w26416_ ;
	wire _w26417_ ;
	wire _w26418_ ;
	wire _w26419_ ;
	wire _w26420_ ;
	wire _w26421_ ;
	wire _w26422_ ;
	wire _w26423_ ;
	wire _w26424_ ;
	wire _w26425_ ;
	wire _w26426_ ;
	wire _w26427_ ;
	wire _w26428_ ;
	wire _w26429_ ;
	wire _w26430_ ;
	wire _w26431_ ;
	wire _w26432_ ;
	wire _w26433_ ;
	wire _w26434_ ;
	wire _w26435_ ;
	wire _w26436_ ;
	wire _w26437_ ;
	wire _w26438_ ;
	wire _w26439_ ;
	wire _w26440_ ;
	wire _w26441_ ;
	wire _w26442_ ;
	wire _w26443_ ;
	wire _w26444_ ;
	wire _w26445_ ;
	wire _w26446_ ;
	wire _w26447_ ;
	wire _w26448_ ;
	wire _w26449_ ;
	wire _w26450_ ;
	wire _w26451_ ;
	wire _w26452_ ;
	wire _w26453_ ;
	wire _w26454_ ;
	wire _w26455_ ;
	wire _w26456_ ;
	wire _w26457_ ;
	wire _w26458_ ;
	wire _w26459_ ;
	wire _w26460_ ;
	wire _w26461_ ;
	wire _w26462_ ;
	wire _w26463_ ;
	wire _w26464_ ;
	wire _w26465_ ;
	wire _w26466_ ;
	wire _w26467_ ;
	wire _w26468_ ;
	wire _w26469_ ;
	wire _w26470_ ;
	wire _w26471_ ;
	wire _w26472_ ;
	wire _w26473_ ;
	wire _w26474_ ;
	wire _w26475_ ;
	wire _w26476_ ;
	wire _w26477_ ;
	wire _w26478_ ;
	wire _w26479_ ;
	wire _w26480_ ;
	wire _w26481_ ;
	wire _w26482_ ;
	wire _w26483_ ;
	wire _w26484_ ;
	wire _w26485_ ;
	wire _w26486_ ;
	wire _w26487_ ;
	wire _w26488_ ;
	wire _w26489_ ;
	wire _w26490_ ;
	wire _w26491_ ;
	wire _w26492_ ;
	wire _w26493_ ;
	wire _w26494_ ;
	wire _w26495_ ;
	wire _w26496_ ;
	wire _w26497_ ;
	wire _w26498_ ;
	wire _w26499_ ;
	wire _w26500_ ;
	wire _w26501_ ;
	wire _w26502_ ;
	wire _w26503_ ;
	wire _w26504_ ;
	wire _w26505_ ;
	wire _w26506_ ;
	wire _w26507_ ;
	wire _w26508_ ;
	wire _w26509_ ;
	wire _w26510_ ;
	wire _w26511_ ;
	wire _w26512_ ;
	wire _w26513_ ;
	wire _w26514_ ;
	wire _w26515_ ;
	wire _w26516_ ;
	wire _w26517_ ;
	wire _w26518_ ;
	wire _w26519_ ;
	wire _w26520_ ;
	wire _w26521_ ;
	wire _w26522_ ;
	wire _w26523_ ;
	wire _w26524_ ;
	wire _w26525_ ;
	wire _w26526_ ;
	wire _w26527_ ;
	wire _w26528_ ;
	wire _w26529_ ;
	wire _w26530_ ;
	wire _w26531_ ;
	wire _w26532_ ;
	wire _w26533_ ;
	wire _w26534_ ;
	wire _w26535_ ;
	wire _w26536_ ;
	wire _w26537_ ;
	wire _w26538_ ;
	wire _w26539_ ;
	wire _w26540_ ;
	wire _w26541_ ;
	wire _w26542_ ;
	wire _w26543_ ;
	wire _w26544_ ;
	wire _w26545_ ;
	wire _w26546_ ;
	wire _w26547_ ;
	wire _w26548_ ;
	wire _w26549_ ;
	wire _w26550_ ;
	wire _w26551_ ;
	wire _w26552_ ;
	wire _w26553_ ;
	wire _w26554_ ;
	wire _w26555_ ;
	wire _w26556_ ;
	wire _w26557_ ;
	wire _w26558_ ;
	wire _w26559_ ;
	wire _w26560_ ;
	wire _w26561_ ;
	wire _w26562_ ;
	wire _w26563_ ;
	wire _w26564_ ;
	wire _w26565_ ;
	wire _w26566_ ;
	wire _w26567_ ;
	wire _w26568_ ;
	wire _w26569_ ;
	wire _w26570_ ;
	wire _w26571_ ;
	wire _w26572_ ;
	wire _w26573_ ;
	wire _w26574_ ;
	wire _w26575_ ;
	wire _w26576_ ;
	wire _w26577_ ;
	wire _w26578_ ;
	wire _w26579_ ;
	wire _w26580_ ;
	wire _w26581_ ;
	wire _w26582_ ;
	wire _w26583_ ;
	wire _w26584_ ;
	wire _w26585_ ;
	wire _w26586_ ;
	wire _w26587_ ;
	wire _w26588_ ;
	wire _w26589_ ;
	wire _w26590_ ;
	wire _w26591_ ;
	wire _w26592_ ;
	wire _w26593_ ;
	wire _w26594_ ;
	wire _w26595_ ;
	wire _w26596_ ;
	wire _w26597_ ;
	wire _w26598_ ;
	wire _w26599_ ;
	wire _w26600_ ;
	wire _w26601_ ;
	wire _w26602_ ;
	wire _w26603_ ;
	wire _w26604_ ;
	wire _w26605_ ;
	wire _w26606_ ;
	wire _w26607_ ;
	wire _w26608_ ;
	wire _w26609_ ;
	wire _w26610_ ;
	wire _w26611_ ;
	wire _w26612_ ;
	wire _w26613_ ;
	wire _w26614_ ;
	wire _w26615_ ;
	wire _w26616_ ;
	wire _w26617_ ;
	wire _w26618_ ;
	wire _w26619_ ;
	wire _w26620_ ;
	wire _w26621_ ;
	wire _w26622_ ;
	wire _w26623_ ;
	wire _w26624_ ;
	wire _w26625_ ;
	wire _w26626_ ;
	wire _w26627_ ;
	wire _w26628_ ;
	wire _w26629_ ;
	wire _w26630_ ;
	wire _w26631_ ;
	wire _w26632_ ;
	wire _w26633_ ;
	wire _w26634_ ;
	wire _w26635_ ;
	wire _w26636_ ;
	wire _w26637_ ;
	wire _w26638_ ;
	wire _w26639_ ;
	wire _w26640_ ;
	wire _w26641_ ;
	wire _w26642_ ;
	wire _w26643_ ;
	wire _w26644_ ;
	wire _w26645_ ;
	wire _w26646_ ;
	wire _w26647_ ;
	wire _w26648_ ;
	wire _w26649_ ;
	wire _w26650_ ;
	wire _w26651_ ;
	wire _w26652_ ;
	wire _w26653_ ;
	wire _w26654_ ;
	wire _w26655_ ;
	wire _w26656_ ;
	wire _w26657_ ;
	wire _w26658_ ;
	wire _w26659_ ;
	wire _w26660_ ;
	wire _w26661_ ;
	wire _w26662_ ;
	wire _w26663_ ;
	wire _w26664_ ;
	wire _w26665_ ;
	wire _w26666_ ;
	wire _w26667_ ;
	wire _w26668_ ;
	wire _w26669_ ;
	wire _w26670_ ;
	wire _w26671_ ;
	wire _w26672_ ;
	wire _w26673_ ;
	wire _w26674_ ;
	wire _w26675_ ;
	wire _w26676_ ;
	wire _w26677_ ;
	wire _w26678_ ;
	wire _w26679_ ;
	wire _w26680_ ;
	wire _w26681_ ;
	wire _w26682_ ;
	wire _w26683_ ;
	wire _w26684_ ;
	wire _w26685_ ;
	wire _w26686_ ;
	wire _w26687_ ;
	wire _w26688_ ;
	wire _w26689_ ;
	wire _w26690_ ;
	wire _w26691_ ;
	wire _w26692_ ;
	wire _w26693_ ;
	wire _w26694_ ;
	wire _w26695_ ;
	wire _w26696_ ;
	wire _w26697_ ;
	wire _w26698_ ;
	wire _w26699_ ;
	wire _w26700_ ;
	wire _w26701_ ;
	wire _w26702_ ;
	wire _w26703_ ;
	wire _w26704_ ;
	wire _w26705_ ;
	wire _w26706_ ;
	wire _w26707_ ;
	wire _w26708_ ;
	wire _w26709_ ;
	wire _w26710_ ;
	wire _w26711_ ;
	wire _w26712_ ;
	wire _w26713_ ;
	wire _w26714_ ;
	wire _w26715_ ;
	wire _w26716_ ;
	wire _w26717_ ;
	wire _w26718_ ;
	wire _w26719_ ;
	wire _w26720_ ;
	wire _w26721_ ;
	wire _w26722_ ;
	wire _w26723_ ;
	wire _w26724_ ;
	wire _w26725_ ;
	wire _w26726_ ;
	wire _w26727_ ;
	wire _w26728_ ;
	wire _w26729_ ;
	wire _w26730_ ;
	wire _w26731_ ;
	wire _w26732_ ;
	wire _w26733_ ;
	wire _w26734_ ;
	wire _w26735_ ;
	wire _w26736_ ;
	wire _w26737_ ;
	wire _w26738_ ;
	wire _w26739_ ;
	wire _w26740_ ;
	wire _w26741_ ;
	wire _w26742_ ;
	wire _w26743_ ;
	wire _w26744_ ;
	wire _w26745_ ;
	wire _w26746_ ;
	wire _w26747_ ;
	wire _w26748_ ;
	wire _w26749_ ;
	wire _w26750_ ;
	wire _w26751_ ;
	wire _w26752_ ;
	wire _w26753_ ;
	wire _w26754_ ;
	wire _w26755_ ;
	wire _w26756_ ;
	wire _w26757_ ;
	wire _w26758_ ;
	wire _w26759_ ;
	wire _w26760_ ;
	wire _w26761_ ;
	wire _w26762_ ;
	wire _w26763_ ;
	wire _w26764_ ;
	wire _w26765_ ;
	wire _w26766_ ;
	wire _w26767_ ;
	wire _w26768_ ;
	wire _w26769_ ;
	wire _w26770_ ;
	wire _w26771_ ;
	wire _w26772_ ;
	wire _w26773_ ;
	wire _w26774_ ;
	wire _w26775_ ;
	wire _w26776_ ;
	wire _w26777_ ;
	wire _w26778_ ;
	wire _w26779_ ;
	wire _w26780_ ;
	wire _w26781_ ;
	wire _w26782_ ;
	wire _w26783_ ;
	wire _w26784_ ;
	wire _w26785_ ;
	wire _w26786_ ;
	wire _w26787_ ;
	wire _w26788_ ;
	wire _w26789_ ;
	wire _w26790_ ;
	wire _w26791_ ;
	wire _w26792_ ;
	wire _w26793_ ;
	wire _w26794_ ;
	wire _w26795_ ;
	wire _w26796_ ;
	wire _w26797_ ;
	wire _w26798_ ;
	wire _w26799_ ;
	wire _w26800_ ;
	wire _w26801_ ;
	wire _w26802_ ;
	wire _w26803_ ;
	wire _w26804_ ;
	wire _w26805_ ;
	wire _w26806_ ;
	wire _w26807_ ;
	wire _w26808_ ;
	wire _w26809_ ;
	wire _w26810_ ;
	wire _w26811_ ;
	wire _w26812_ ;
	wire _w26813_ ;
	wire _w26814_ ;
	wire _w26815_ ;
	wire _w26816_ ;
	wire _w26817_ ;
	wire _w26818_ ;
	wire _w26819_ ;
	wire _w26820_ ;
	wire _w26821_ ;
	wire _w26822_ ;
	wire _w26823_ ;
	wire _w26824_ ;
	wire _w26825_ ;
	wire _w26826_ ;
	wire _w26827_ ;
	wire _w26828_ ;
	wire _w26829_ ;
	wire _w26830_ ;
	wire _w26831_ ;
	wire _w26832_ ;
	wire _w26833_ ;
	wire _w26834_ ;
	wire _w26835_ ;
	wire _w26836_ ;
	wire _w26837_ ;
	wire _w26838_ ;
	wire _w26839_ ;
	wire _w26840_ ;
	wire _w26841_ ;
	wire _w26842_ ;
	wire _w26843_ ;
	wire _w26844_ ;
	wire _w26845_ ;
	wire _w26846_ ;
	wire _w26847_ ;
	wire _w26848_ ;
	wire _w26849_ ;
	wire _w26850_ ;
	wire _w26851_ ;
	wire _w26852_ ;
	wire _w26853_ ;
	wire _w26854_ ;
	wire _w26855_ ;
	wire _w26856_ ;
	wire _w26857_ ;
	wire _w26858_ ;
	wire _w26859_ ;
	wire _w26860_ ;
	wire _w26861_ ;
	wire _w26862_ ;
	wire _w26863_ ;
	wire _w26864_ ;
	wire _w26865_ ;
	wire _w26866_ ;
	wire _w26867_ ;
	wire _w26868_ ;
	wire _w26869_ ;
	wire _w26870_ ;
	wire _w26871_ ;
	wire _w26872_ ;
	wire _w26873_ ;
	wire _w26874_ ;
	wire _w26875_ ;
	wire _w26876_ ;
	wire _w26877_ ;
	wire _w26878_ ;
	wire _w26879_ ;
	wire _w26880_ ;
	wire _w26881_ ;
	wire _w26882_ ;
	wire _w26883_ ;
	wire _w26884_ ;
	wire _w26885_ ;
	wire _w26886_ ;
	wire _w26887_ ;
	wire _w26888_ ;
	wire _w26889_ ;
	wire _w26890_ ;
	wire _w26891_ ;
	wire _w26892_ ;
	wire _w26893_ ;
	wire _w26894_ ;
	wire _w26895_ ;
	wire _w26896_ ;
	wire _w26897_ ;
	wire _w26898_ ;
	wire _w26899_ ;
	wire _w26900_ ;
	wire _w26901_ ;
	wire _w26902_ ;
	wire _w26903_ ;
	wire _w26904_ ;
	wire _w26905_ ;
	wire _w26906_ ;
	wire _w26907_ ;
	wire _w26908_ ;
	wire _w26909_ ;
	wire _w26910_ ;
	wire _w26911_ ;
	wire _w26912_ ;
	wire _w26913_ ;
	wire _w26914_ ;
	wire _w26915_ ;
	wire _w26916_ ;
	wire _w26917_ ;
	wire _w26918_ ;
	wire _w26919_ ;
	wire _w26920_ ;
	wire _w26921_ ;
	wire _w26922_ ;
	wire _w26923_ ;
	wire _w26924_ ;
	wire _w26925_ ;
	wire _w26926_ ;
	wire _w26927_ ;
	wire _w26928_ ;
	wire _w26929_ ;
	wire _w26930_ ;
	wire _w26931_ ;
	wire _w26932_ ;
	wire _w26933_ ;
	wire _w26934_ ;
	wire _w26935_ ;
	wire _w26936_ ;
	wire _w26937_ ;
	wire _w26938_ ;
	wire _w26939_ ;
	wire _w26940_ ;
	wire _w26941_ ;
	wire _w26942_ ;
	wire _w26943_ ;
	wire _w26944_ ;
	wire _w26945_ ;
	wire _w26946_ ;
	wire _w26947_ ;
	wire _w26948_ ;
	wire _w26949_ ;
	wire _w26950_ ;
	wire _w26951_ ;
	wire _w26952_ ;
	wire _w26953_ ;
	wire _w26954_ ;
	wire _w26955_ ;
	wire _w26956_ ;
	wire _w26957_ ;
	wire _w26958_ ;
	wire _w26959_ ;
	wire _w26960_ ;
	wire _w26961_ ;
	wire _w26962_ ;
	wire _w26963_ ;
	wire _w26964_ ;
	wire _w26965_ ;
	wire _w26966_ ;
	wire _w26967_ ;
	wire _w26968_ ;
	wire _w26969_ ;
	wire _w26970_ ;
	wire _w26971_ ;
	wire _w26972_ ;
	wire _w26973_ ;
	wire _w26974_ ;
	wire _w26975_ ;
	wire _w26976_ ;
	wire _w26977_ ;
	wire _w26978_ ;
	wire _w26979_ ;
	wire _w26980_ ;
	wire _w26981_ ;
	wire _w26982_ ;
	wire _w26983_ ;
	wire _w26984_ ;
	wire _w26985_ ;
	wire _w26986_ ;
	wire _w26987_ ;
	wire _w26988_ ;
	wire _w26989_ ;
	wire _w26990_ ;
	wire _w26991_ ;
	wire _w26992_ ;
	wire _w26993_ ;
	wire _w26994_ ;
	wire _w26995_ ;
	wire _w26996_ ;
	wire _w26997_ ;
	wire _w26998_ ;
	wire _w26999_ ;
	wire _w27000_ ;
	wire _w27001_ ;
	wire _w27002_ ;
	wire _w27003_ ;
	wire _w27004_ ;
	wire _w27005_ ;
	wire _w27006_ ;
	wire _w27007_ ;
	wire _w27008_ ;
	wire _w27009_ ;
	wire _w27010_ ;
	wire _w27011_ ;
	wire _w27012_ ;
	wire _w27013_ ;
	wire _w27014_ ;
	wire _w27015_ ;
	wire _w27016_ ;
	wire _w27017_ ;
	wire _w27018_ ;
	wire _w27019_ ;
	wire _w27020_ ;
	wire _w27021_ ;
	wire _w27022_ ;
	wire _w27023_ ;
	wire _w27024_ ;
	wire _w27025_ ;
	wire _w27026_ ;
	wire _w27027_ ;
	wire _w27028_ ;
	wire _w27029_ ;
	wire _w27030_ ;
	wire _w27031_ ;
	wire _w27032_ ;
	wire _w27033_ ;
	wire _w27034_ ;
	wire _w27035_ ;
	wire _w27036_ ;
	wire _w27037_ ;
	wire _w27038_ ;
	wire _w27039_ ;
	wire _w27040_ ;
	wire _w27041_ ;
	wire _w27042_ ;
	wire _w27043_ ;
	wire _w27044_ ;
	wire _w27045_ ;
	wire _w27046_ ;
	wire _w27047_ ;
	wire _w27048_ ;
	wire _w27049_ ;
	wire _w27050_ ;
	wire _w27051_ ;
	wire _w27052_ ;
	wire _w27053_ ;
	wire _w27054_ ;
	wire _w27055_ ;
	wire _w27056_ ;
	wire _w27057_ ;
	wire _w27058_ ;
	wire _w27059_ ;
	wire _w27060_ ;
	wire _w27061_ ;
	wire _w27062_ ;
	wire _w27063_ ;
	wire _w27064_ ;
	wire _w27065_ ;
	wire _w27066_ ;
	wire _w27067_ ;
	wire _w27068_ ;
	wire _w27069_ ;
	wire _w27070_ ;
	wire _w27071_ ;
	wire _w27072_ ;
	wire _w27073_ ;
	wire _w27074_ ;
	wire _w27075_ ;
	wire _w27076_ ;
	wire _w27077_ ;
	wire _w27078_ ;
	wire _w27079_ ;
	wire _w27080_ ;
	wire _w27081_ ;
	wire _w27082_ ;
	wire _w27083_ ;
	wire _w27084_ ;
	wire _w27085_ ;
	wire _w27086_ ;
	wire _w27087_ ;
	wire _w27088_ ;
	wire _w27089_ ;
	wire _w27090_ ;
	wire _w27091_ ;
	wire _w27092_ ;
	wire _w27093_ ;
	wire _w27094_ ;
	wire _w27095_ ;
	wire _w27096_ ;
	wire _w27097_ ;
	wire _w27098_ ;
	wire _w27099_ ;
	wire _w27100_ ;
	wire _w27101_ ;
	wire _w27102_ ;
	wire _w27103_ ;
	wire _w27104_ ;
	wire _w27105_ ;
	wire _w27106_ ;
	wire _w27107_ ;
	wire _w27108_ ;
	wire _w27109_ ;
	wire _w27110_ ;
	wire _w27111_ ;
	wire _w27112_ ;
	wire _w27113_ ;
	wire _w27114_ ;
	wire _w27115_ ;
	wire _w27116_ ;
	wire _w27117_ ;
	wire _w27118_ ;
	wire _w27119_ ;
	wire _w27120_ ;
	wire _w27121_ ;
	wire _w27122_ ;
	wire _w27123_ ;
	wire _w27124_ ;
	wire _w27125_ ;
	wire _w27126_ ;
	wire _w27127_ ;
	wire _w27128_ ;
	wire _w27129_ ;
	wire _w27130_ ;
	wire _w27131_ ;
	wire _w27132_ ;
	wire _w27133_ ;
	wire _w27134_ ;
	wire _w27135_ ;
	wire _w27136_ ;
	wire _w27137_ ;
	wire _w27138_ ;
	wire _w27139_ ;
	wire _w27140_ ;
	wire _w27141_ ;
	wire _w27142_ ;
	wire _w27143_ ;
	wire _w27144_ ;
	wire _w27145_ ;
	wire _w27146_ ;
	wire _w27147_ ;
	wire _w27148_ ;
	wire _w27149_ ;
	wire _w27150_ ;
	wire _w27151_ ;
	wire _w27152_ ;
	wire _w27153_ ;
	wire _w27154_ ;
	wire _w27155_ ;
	wire _w27156_ ;
	wire _w27157_ ;
	wire _w27158_ ;
	wire _w27159_ ;
	wire _w27160_ ;
	wire _w27161_ ;
	wire _w27162_ ;
	wire _w27163_ ;
	wire _w27164_ ;
	wire _w27165_ ;
	wire _w27166_ ;
	wire _w27167_ ;
	wire _w27168_ ;
	wire _w27169_ ;
	wire _w27170_ ;
	wire _w27171_ ;
	wire _w27172_ ;
	wire _w27173_ ;
	wire _w27174_ ;
	wire _w27175_ ;
	wire _w27176_ ;
	wire _w27177_ ;
	wire _w27178_ ;
	wire _w27179_ ;
	wire _w27180_ ;
	wire _w27181_ ;
	wire _w27182_ ;
	wire _w27183_ ;
	wire _w27184_ ;
	wire _w27185_ ;
	wire _w27186_ ;
	wire _w27187_ ;
	wire _w27188_ ;
	wire _w27189_ ;
	wire _w27190_ ;
	wire _w27191_ ;
	wire _w27192_ ;
	wire _w27193_ ;
	wire _w27194_ ;
	wire _w27195_ ;
	wire _w27196_ ;
	wire _w27197_ ;
	wire _w27198_ ;
	wire _w27199_ ;
	wire _w27200_ ;
	wire _w27201_ ;
	wire _w27202_ ;
	wire _w27203_ ;
	wire _w27204_ ;
	wire _w27205_ ;
	wire _w27206_ ;
	wire _w27207_ ;
	wire _w27208_ ;
	wire _w27209_ ;
	wire _w27210_ ;
	wire _w27211_ ;
	wire _w27212_ ;
	wire _w27213_ ;
	wire _w27214_ ;
	wire _w27215_ ;
	wire _w27216_ ;
	wire _w27217_ ;
	wire _w27218_ ;
	wire _w27219_ ;
	wire _w27220_ ;
	wire _w27221_ ;
	wire _w27222_ ;
	wire _w27223_ ;
	wire _w27224_ ;
	wire _w27225_ ;
	wire _w27226_ ;
	wire _w27227_ ;
	wire _w27228_ ;
	wire _w27229_ ;
	wire _w27230_ ;
	wire _w27231_ ;
	wire _w27232_ ;
	wire _w27233_ ;
	wire _w27234_ ;
	wire _w27235_ ;
	wire _w27236_ ;
	wire _w27237_ ;
	wire _w27238_ ;
	wire _w27239_ ;
	wire _w27240_ ;
	wire _w27241_ ;
	wire _w27242_ ;
	wire _w27243_ ;
	wire _w27244_ ;
	wire _w27245_ ;
	wire _w27246_ ;
	wire _w27247_ ;
	wire _w27248_ ;
	wire _w27249_ ;
	wire _w27250_ ;
	wire _w27251_ ;
	wire _w27252_ ;
	wire _w27253_ ;
	wire _w27254_ ;
	wire _w27255_ ;
	wire _w27256_ ;
	wire _w27257_ ;
	wire _w27258_ ;
	wire _w27259_ ;
	wire _w27260_ ;
	wire _w27261_ ;
	wire _w27262_ ;
	wire _w27263_ ;
	wire _w27264_ ;
	wire _w27265_ ;
	wire _w27266_ ;
	wire _w27267_ ;
	wire _w27268_ ;
	wire _w27269_ ;
	wire _w27270_ ;
	wire _w27271_ ;
	wire _w27272_ ;
	wire _w27273_ ;
	wire _w27274_ ;
	wire _w27275_ ;
	wire _w27276_ ;
	wire _w27277_ ;
	wire _w27278_ ;
	wire _w27279_ ;
	wire _w27280_ ;
	wire _w27281_ ;
	wire _w27282_ ;
	wire _w27283_ ;
	wire _w27284_ ;
	wire _w27285_ ;
	wire _w27286_ ;
	wire _w27287_ ;
	wire _w27288_ ;
	wire _w27289_ ;
	wire _w27290_ ;
	wire _w27291_ ;
	wire _w27292_ ;
	wire _w27293_ ;
	wire _w27294_ ;
	wire _w27295_ ;
	wire _w27296_ ;
	wire _w27297_ ;
	wire _w27298_ ;
	wire _w27299_ ;
	wire _w27300_ ;
	wire _w27301_ ;
	wire _w27302_ ;
	wire _w27303_ ;
	wire _w27304_ ;
	wire _w27305_ ;
	wire _w27306_ ;
	wire _w27307_ ;
	wire _w27308_ ;
	wire _w27309_ ;
	wire _w27310_ ;
	wire _w27311_ ;
	wire _w27312_ ;
	wire _w27313_ ;
	wire _w27314_ ;
	wire _w27315_ ;
	wire _w27316_ ;
	wire _w27317_ ;
	wire _w27318_ ;
	wire _w27319_ ;
	wire _w27320_ ;
	wire _w27321_ ;
	wire _w27322_ ;
	wire _w27323_ ;
	wire _w27324_ ;
	wire _w27325_ ;
	wire _w27326_ ;
	wire _w27327_ ;
	wire _w27328_ ;
	wire _w27329_ ;
	wire _w27330_ ;
	wire _w27331_ ;
	wire _w27332_ ;
	wire _w27333_ ;
	wire _w27334_ ;
	wire _w27335_ ;
	wire _w27336_ ;
	wire _w27337_ ;
	wire _w27338_ ;
	wire _w27339_ ;
	wire _w27340_ ;
	wire _w27341_ ;
	wire _w27342_ ;
	wire _w27343_ ;
	wire _w27344_ ;
	wire _w27345_ ;
	wire _w27346_ ;
	wire _w27347_ ;
	wire _w27348_ ;
	wire _w27349_ ;
	wire _w27350_ ;
	wire _w27351_ ;
	wire _w27352_ ;
	wire _w27353_ ;
	wire _w27354_ ;
	wire _w27355_ ;
	wire _w27356_ ;
	wire _w27357_ ;
	wire _w27358_ ;
	wire _w27359_ ;
	wire _w27360_ ;
	wire _w27361_ ;
	wire _w27362_ ;
	wire _w27363_ ;
	wire _w27364_ ;
	wire _w27365_ ;
	wire _w27366_ ;
	wire _w27367_ ;
	wire _w27368_ ;
	wire _w27369_ ;
	wire _w27370_ ;
	wire _w27371_ ;
	wire _w27372_ ;
	wire _w27373_ ;
	wire _w27374_ ;
	wire _w27375_ ;
	wire _w27376_ ;
	wire _w27377_ ;
	wire _w27378_ ;
	wire _w27379_ ;
	wire _w27380_ ;
	wire _w27381_ ;
	wire _w27382_ ;
	wire _w27383_ ;
	wire _w27384_ ;
	wire _w27385_ ;
	wire _w27386_ ;
	wire _w27387_ ;
	wire _w27388_ ;
	wire _w27389_ ;
	wire _w27390_ ;
	wire _w27391_ ;
	wire _w27392_ ;
	wire _w27393_ ;
	wire _w27394_ ;
	wire _w27395_ ;
	wire _w27396_ ;
	wire _w27397_ ;
	wire _w27398_ ;
	wire _w27399_ ;
	wire _w27400_ ;
	wire _w27401_ ;
	wire _w27402_ ;
	wire _w27403_ ;
	wire _w27404_ ;
	wire _w27405_ ;
	wire _w27406_ ;
	wire _w27407_ ;
	wire _w27408_ ;
	wire _w27409_ ;
	wire _w27410_ ;
	wire _w27411_ ;
	wire _w27412_ ;
	wire _w27413_ ;
	wire _w27414_ ;
	wire _w27415_ ;
	wire _w27416_ ;
	wire _w27417_ ;
	wire _w27418_ ;
	wire _w27419_ ;
	wire _w27420_ ;
	wire _w27421_ ;
	wire _w27422_ ;
	wire _w27423_ ;
	wire _w27424_ ;
	wire _w27425_ ;
	wire _w27426_ ;
	wire _w27427_ ;
	wire _w27428_ ;
	wire _w27429_ ;
	wire _w27430_ ;
	wire _w27431_ ;
	wire _w27432_ ;
	wire _w27433_ ;
	wire _w27434_ ;
	wire _w27435_ ;
	wire _w27436_ ;
	wire _w27437_ ;
	wire _w27438_ ;
	wire _w27439_ ;
	wire _w27440_ ;
	wire _w27441_ ;
	wire _w27442_ ;
	wire _w27443_ ;
	wire _w27444_ ;
	wire _w27445_ ;
	wire _w27446_ ;
	wire _w27447_ ;
	wire _w27448_ ;
	wire _w27449_ ;
	wire _w27450_ ;
	wire _w27451_ ;
	wire _w27452_ ;
	wire _w27453_ ;
	wire _w27454_ ;
	wire _w27455_ ;
	wire _w27456_ ;
	wire _w27457_ ;
	wire _w27458_ ;
	wire _w27459_ ;
	wire _w27460_ ;
	wire _w27461_ ;
	wire _w27462_ ;
	wire _w27463_ ;
	wire _w27464_ ;
	wire _w27465_ ;
	wire _w27466_ ;
	wire _w27467_ ;
	wire _w27468_ ;
	wire _w27469_ ;
	wire _w27470_ ;
	wire _w27471_ ;
	wire _w27472_ ;
	wire _w27473_ ;
	wire _w27474_ ;
	wire _w27475_ ;
	wire _w27476_ ;
	wire _w27477_ ;
	wire _w27478_ ;
	wire _w27479_ ;
	wire _w27480_ ;
	wire _w27481_ ;
	wire _w27482_ ;
	wire _w27483_ ;
	wire _w27484_ ;
	wire _w27485_ ;
	wire _w27486_ ;
	wire _w27487_ ;
	wire _w27488_ ;
	wire _w27489_ ;
	wire _w27490_ ;
	wire _w27491_ ;
	wire _w27492_ ;
	wire _w27493_ ;
	wire _w27494_ ;
	wire _w27495_ ;
	wire _w27496_ ;
	wire _w27497_ ;
	wire _w27498_ ;
	wire _w27499_ ;
	wire _w27500_ ;
	wire _w27501_ ;
	wire _w27502_ ;
	wire _w27503_ ;
	wire _w27504_ ;
	wire _w27505_ ;
	wire _w27506_ ;
	wire _w27507_ ;
	wire _w27508_ ;
	wire _w27509_ ;
	wire _w27510_ ;
	wire _w27511_ ;
	wire _w27512_ ;
	wire _w27513_ ;
	wire _w27514_ ;
	wire _w27515_ ;
	wire _w27516_ ;
	wire _w27517_ ;
	wire _w27518_ ;
	wire _w27519_ ;
	wire _w27520_ ;
	wire _w27521_ ;
	wire _w27522_ ;
	wire _w27523_ ;
	wire _w27524_ ;
	wire _w27525_ ;
	wire _w27526_ ;
	wire _w27527_ ;
	wire _w27528_ ;
	wire _w27529_ ;
	wire _w27530_ ;
	wire _w27531_ ;
	wire _w27532_ ;
	wire _w27533_ ;
	wire _w27534_ ;
	wire _w27535_ ;
	wire _w27536_ ;
	wire _w27537_ ;
	wire _w27538_ ;
	wire _w27539_ ;
	wire _w27540_ ;
	wire _w27541_ ;
	wire _w27542_ ;
	wire _w27543_ ;
	wire _w27544_ ;
	wire _w27545_ ;
	wire _w27546_ ;
	wire _w27547_ ;
	wire _w27548_ ;
	wire _w27549_ ;
	wire _w27550_ ;
	wire _w27551_ ;
	wire _w27552_ ;
	wire _w27553_ ;
	wire _w27554_ ;
	wire _w27555_ ;
	wire _w27556_ ;
	wire _w27557_ ;
	wire _w27558_ ;
	wire _w27559_ ;
	wire _w27560_ ;
	wire _w27561_ ;
	wire _w27562_ ;
	wire _w27563_ ;
	wire _w27564_ ;
	wire _w27565_ ;
	wire _w27566_ ;
	wire _w27567_ ;
	wire _w27568_ ;
	wire _w27569_ ;
	wire _w27570_ ;
	wire _w27571_ ;
	wire _w27572_ ;
	wire _w27573_ ;
	wire _w27574_ ;
	wire _w27575_ ;
	wire _w27576_ ;
	wire _w27577_ ;
	wire _w27578_ ;
	wire _w27579_ ;
	wire _w27580_ ;
	wire _w27581_ ;
	wire _w27582_ ;
	wire _w27583_ ;
	wire _w27584_ ;
	wire _w27585_ ;
	wire _w27586_ ;
	wire _w27587_ ;
	wire _w27588_ ;
	wire _w27589_ ;
	wire _w27590_ ;
	wire _w27591_ ;
	wire _w27592_ ;
	wire _w27593_ ;
	wire _w27594_ ;
	wire _w27595_ ;
	wire _w27596_ ;
	wire _w27597_ ;
	wire _w27598_ ;
	wire _w27599_ ;
	wire _w27600_ ;
	wire _w27601_ ;
	wire _w27602_ ;
	wire _w27603_ ;
	wire _w27604_ ;
	wire _w27605_ ;
	wire _w27606_ ;
	wire _w27607_ ;
	wire _w27608_ ;
	wire _w27609_ ;
	wire _w27610_ ;
	wire _w27611_ ;
	wire _w27612_ ;
	wire _w27613_ ;
	wire _w27614_ ;
	wire _w27615_ ;
	wire _w27616_ ;
	wire _w27617_ ;
	wire _w27618_ ;
	wire _w27619_ ;
	wire _w27620_ ;
	wire _w27621_ ;
	wire _w27622_ ;
	wire _w27623_ ;
	wire _w27624_ ;
	wire _w27625_ ;
	wire _w27626_ ;
	wire _w27627_ ;
	wire _w27628_ ;
	wire _w27629_ ;
	wire _w27630_ ;
	wire _w27631_ ;
	wire _w27632_ ;
	wire _w27633_ ;
	wire _w27634_ ;
	wire _w27635_ ;
	wire _w27636_ ;
	wire _w27637_ ;
	wire _w27638_ ;
	wire _w27639_ ;
	wire _w27640_ ;
	wire _w27641_ ;
	wire _w27642_ ;
	wire _w27643_ ;
	wire _w27644_ ;
	wire _w27645_ ;
	wire _w27646_ ;
	wire _w27647_ ;
	wire _w27648_ ;
	wire _w27649_ ;
	wire _w27650_ ;
	wire _w27651_ ;
	wire _w27652_ ;
	wire _w27653_ ;
	wire _w27654_ ;
	wire _w27655_ ;
	wire _w27656_ ;
	wire _w27657_ ;
	wire _w27658_ ;
	wire _w27659_ ;
	wire _w27660_ ;
	wire _w27661_ ;
	wire _w27662_ ;
	wire _w27663_ ;
	wire _w27664_ ;
	wire _w27665_ ;
	wire _w27666_ ;
	wire _w27667_ ;
	wire _w27668_ ;
	wire _w27669_ ;
	wire _w27670_ ;
	wire _w27671_ ;
	wire _w27672_ ;
	wire _w27673_ ;
	wire _w27674_ ;
	wire _w27675_ ;
	wire _w27676_ ;
	wire _w27677_ ;
	wire _w27678_ ;
	wire _w27679_ ;
	wire _w27680_ ;
	wire _w27681_ ;
	wire _w27682_ ;
	wire _w27683_ ;
	wire _w27684_ ;
	wire _w27685_ ;
	wire _w27686_ ;
	wire _w27687_ ;
	wire _w27688_ ;
	wire _w27689_ ;
	wire _w27690_ ;
	wire _w27691_ ;
	wire _w27692_ ;
	wire _w27693_ ;
	wire _w27694_ ;
	wire _w27695_ ;
	wire _w27696_ ;
	wire _w27697_ ;
	wire _w27698_ ;
	wire _w27699_ ;
	wire _w27700_ ;
	wire _w27701_ ;
	wire _w27702_ ;
	wire _w27703_ ;
	wire _w27704_ ;
	wire _w27705_ ;
	wire _w27706_ ;
	wire _w27707_ ;
	wire _w27708_ ;
	wire _w27709_ ;
	wire _w27710_ ;
	wire _w27711_ ;
	wire _w27712_ ;
	wire _w27713_ ;
	wire _w27714_ ;
	wire _w27715_ ;
	wire _w27716_ ;
	wire _w27717_ ;
	wire _w27718_ ;
	wire _w27719_ ;
	wire _w27720_ ;
	wire _w27721_ ;
	wire _w27722_ ;
	wire _w27723_ ;
	wire _w27724_ ;
	wire _w27725_ ;
	wire _w27726_ ;
	wire _w27727_ ;
	wire _w27728_ ;
	wire _w27729_ ;
	wire _w27730_ ;
	wire _w27731_ ;
	wire _w27732_ ;
	wire _w27733_ ;
	wire _w27734_ ;
	wire _w27735_ ;
	wire _w27736_ ;
	wire _w27737_ ;
	wire _w27738_ ;
	wire _w27739_ ;
	wire _w27740_ ;
	wire _w27741_ ;
	wire _w27742_ ;
	wire _w27743_ ;
	wire _w27744_ ;
	wire _w27745_ ;
	wire _w27746_ ;
	wire _w27747_ ;
	wire _w27748_ ;
	wire _w27749_ ;
	wire _w27750_ ;
	wire _w27751_ ;
	wire _w27752_ ;
	wire _w27753_ ;
	wire _w27754_ ;
	wire _w27755_ ;
	wire _w27756_ ;
	wire _w27757_ ;
	wire _w27758_ ;
	wire _w27759_ ;
	wire _w27760_ ;
	wire _w27761_ ;
	wire _w27762_ ;
	wire _w27763_ ;
	wire _w27764_ ;
	wire _w27765_ ;
	wire _w27766_ ;
	wire _w27767_ ;
	wire _w27768_ ;
	wire _w27769_ ;
	wire _w27770_ ;
	wire _w27771_ ;
	wire _w27772_ ;
	wire _w27773_ ;
	wire _w27774_ ;
	wire _w27775_ ;
	wire _w27776_ ;
	wire _w27777_ ;
	wire _w27778_ ;
	wire _w27779_ ;
	wire _w27780_ ;
	wire _w27781_ ;
	wire _w27782_ ;
	wire _w27783_ ;
	wire _w27784_ ;
	wire _w27785_ ;
	wire _w27786_ ;
	wire _w27787_ ;
	wire _w27788_ ;
	wire _w27789_ ;
	wire _w27790_ ;
	wire _w27791_ ;
	wire _w27792_ ;
	wire _w27793_ ;
	wire _w27794_ ;
	wire _w27795_ ;
	wire _w27796_ ;
	wire _w27797_ ;
	wire _w27798_ ;
	wire _w27799_ ;
	wire _w27800_ ;
	wire _w27801_ ;
	wire _w27802_ ;
	wire _w27803_ ;
	wire _w27804_ ;
	wire _w27805_ ;
	wire _w27806_ ;
	wire _w27807_ ;
	wire _w27808_ ;
	wire _w27809_ ;
	wire _w27810_ ;
	wire _w27811_ ;
	wire _w27812_ ;
	wire _w27813_ ;
	wire _w27814_ ;
	wire _w27815_ ;
	wire _w27816_ ;
	wire _w27817_ ;
	wire _w27818_ ;
	wire _w27819_ ;
	wire _w27820_ ;
	wire _w27821_ ;
	wire _w27822_ ;
	wire _w27823_ ;
	wire _w27824_ ;
	wire _w27825_ ;
	wire _w27826_ ;
	wire _w27827_ ;
	wire _w27828_ ;
	wire _w27829_ ;
	wire _w27830_ ;
	wire _w27831_ ;
	wire _w27832_ ;
	wire _w27833_ ;
	wire _w27834_ ;
	wire _w27835_ ;
	wire _w27836_ ;
	wire _w27837_ ;
	wire _w27838_ ;
	wire _w27839_ ;
	wire _w27840_ ;
	wire _w27841_ ;
	wire _w27842_ ;
	wire _w27843_ ;
	wire _w27844_ ;
	wire _w27845_ ;
	wire _w27846_ ;
	wire _w27847_ ;
	wire _w27848_ ;
	wire _w27849_ ;
	wire _w27850_ ;
	wire _w27851_ ;
	wire _w27852_ ;
	wire _w27853_ ;
	wire _w27854_ ;
	wire _w27855_ ;
	wire _w27856_ ;
	wire _w27857_ ;
	wire _w27858_ ;
	wire _w27859_ ;
	wire _w27860_ ;
	wire _w27861_ ;
	wire _w27862_ ;
	wire _w27863_ ;
	wire _w27864_ ;
	wire _w27865_ ;
	wire _w27866_ ;
	wire _w27867_ ;
	wire _w27868_ ;
	wire _w27869_ ;
	wire _w27870_ ;
	wire _w27871_ ;
	wire _w27872_ ;
	wire _w27873_ ;
	wire _w27874_ ;
	wire _w27875_ ;
	wire _w27876_ ;
	wire _w27877_ ;
	wire _w27878_ ;
	wire _w27879_ ;
	wire _w27880_ ;
	wire _w27881_ ;
	wire _w27882_ ;
	wire _w27883_ ;
	wire _w27884_ ;
	wire _w27885_ ;
	wire _w27886_ ;
	wire _w27887_ ;
	wire _w27888_ ;
	wire _w27889_ ;
	wire _w27890_ ;
	wire _w27891_ ;
	wire _w27892_ ;
	wire _w27893_ ;
	wire _w27894_ ;
	wire _w27895_ ;
	wire _w27896_ ;
	wire _w27897_ ;
	wire _w27898_ ;
	wire _w27899_ ;
	wire _w27900_ ;
	wire _w27901_ ;
	wire _w27902_ ;
	wire _w27903_ ;
	wire _w27904_ ;
	wire _w27905_ ;
	wire _w27906_ ;
	wire _w27907_ ;
	wire _w27908_ ;
	wire _w27909_ ;
	wire _w27910_ ;
	wire _w27911_ ;
	wire _w27912_ ;
	wire _w27913_ ;
	wire _w27914_ ;
	wire _w27915_ ;
	wire _w27916_ ;
	wire _w27917_ ;
	wire _w27918_ ;
	wire _w27919_ ;
	wire _w27920_ ;
	wire _w27921_ ;
	wire _w27922_ ;
	wire _w27923_ ;
	wire _w27924_ ;
	wire _w27925_ ;
	wire _w27926_ ;
	wire _w27927_ ;
	wire _w27928_ ;
	wire _w27929_ ;
	wire _w27930_ ;
	wire _w27931_ ;
	wire _w27932_ ;
	wire _w27933_ ;
	wire _w27934_ ;
	wire _w27935_ ;
	wire _w27936_ ;
	wire _w27937_ ;
	wire _w27938_ ;
	wire _w27939_ ;
	wire _w27940_ ;
	wire _w27941_ ;
	wire _w27942_ ;
	wire _w27943_ ;
	wire _w27944_ ;
	wire _w27945_ ;
	wire _w27946_ ;
	wire _w27947_ ;
	wire _w27948_ ;
	wire _w27949_ ;
	wire _w27950_ ;
	wire _w27951_ ;
	wire _w27952_ ;
	wire _w27953_ ;
	wire _w27954_ ;
	wire _w27955_ ;
	wire _w27956_ ;
	wire _w27957_ ;
	wire _w27958_ ;
	wire _w27959_ ;
	wire _w27960_ ;
	wire _w27961_ ;
	wire _w27962_ ;
	wire _w27963_ ;
	wire _w27964_ ;
	wire _w27965_ ;
	wire _w27966_ ;
	wire _w27967_ ;
	wire _w27968_ ;
	wire _w27969_ ;
	wire _w27970_ ;
	wire _w27971_ ;
	wire _w27972_ ;
	wire _w27973_ ;
	wire _w27974_ ;
	wire _w27975_ ;
	wire _w27976_ ;
	wire _w27977_ ;
	wire _w27978_ ;
	wire _w27979_ ;
	wire _w27980_ ;
	wire _w27981_ ;
	wire _w27982_ ;
	wire _w27983_ ;
	wire _w27984_ ;
	wire _w27985_ ;
	wire _w27986_ ;
	wire _w27987_ ;
	wire _w27988_ ;
	wire _w27989_ ;
	wire _w27990_ ;
	wire _w27991_ ;
	wire _w27992_ ;
	wire _w27993_ ;
	wire _w27994_ ;
	wire _w27995_ ;
	wire _w27996_ ;
	wire _w27997_ ;
	wire _w27998_ ;
	wire _w27999_ ;
	wire _w28000_ ;
	wire _w28001_ ;
	wire _w28002_ ;
	wire _w28003_ ;
	wire _w28004_ ;
	wire _w28005_ ;
	wire _w28006_ ;
	wire _w28007_ ;
	wire _w28008_ ;
	wire _w28009_ ;
	wire _w28010_ ;
	wire _w28011_ ;
	wire _w28012_ ;
	wire _w28013_ ;
	wire _w28014_ ;
	wire _w28015_ ;
	wire _w28016_ ;
	wire _w28017_ ;
	wire _w28018_ ;
	wire _w28019_ ;
	wire _w28020_ ;
	wire _w28021_ ;
	wire _w28022_ ;
	wire _w28023_ ;
	wire _w28024_ ;
	wire _w28025_ ;
	wire _w28026_ ;
	wire _w28027_ ;
	wire _w28028_ ;
	wire _w28029_ ;
	wire _w28030_ ;
	wire _w28031_ ;
	wire _w28032_ ;
	wire _w28033_ ;
	wire _w28034_ ;
	wire _w28035_ ;
	wire _w28036_ ;
	wire _w28037_ ;
	wire _w28038_ ;
	wire _w28039_ ;
	wire _w28040_ ;
	wire _w28041_ ;
	wire _w28042_ ;
	wire _w28043_ ;
	wire _w28044_ ;
	wire _w28045_ ;
	wire _w28046_ ;
	wire _w28047_ ;
	wire _w28048_ ;
	wire _w28049_ ;
	wire _w28050_ ;
	wire _w28051_ ;
	wire _w28052_ ;
	wire _w28053_ ;
	wire _w28054_ ;
	wire _w28055_ ;
	wire _w28056_ ;
	wire _w28057_ ;
	wire _w28058_ ;
	wire _w28059_ ;
	wire _w28060_ ;
	wire _w28061_ ;
	wire _w28062_ ;
	wire _w28063_ ;
	wire _w28064_ ;
	wire _w28065_ ;
	wire _w28066_ ;
	wire _w28067_ ;
	wire _w28068_ ;
	wire _w28069_ ;
	wire _w28070_ ;
	wire _w28071_ ;
	wire _w28072_ ;
	wire _w28073_ ;
	wire _w28074_ ;
	wire _w28075_ ;
	wire _w28076_ ;
	wire _w28077_ ;
	wire _w28078_ ;
	wire _w28079_ ;
	wire _w28080_ ;
	wire _w28081_ ;
	wire _w28082_ ;
	wire _w28083_ ;
	wire _w28084_ ;
	wire _w28085_ ;
	wire _w28086_ ;
	wire _w28087_ ;
	wire _w28088_ ;
	wire _w28089_ ;
	wire _w28090_ ;
	wire _w28091_ ;
	wire _w28092_ ;
	wire _w28093_ ;
	wire _w28094_ ;
	wire _w28095_ ;
	wire _w28096_ ;
	wire _w28097_ ;
	wire _w28098_ ;
	wire _w28099_ ;
	wire _w28100_ ;
	wire _w28101_ ;
	wire _w28102_ ;
	wire _w28103_ ;
	wire _w28104_ ;
	wire _w28105_ ;
	wire _w28106_ ;
	wire _w28107_ ;
	wire _w28108_ ;
	wire _w28109_ ;
	wire _w28110_ ;
	wire _w28111_ ;
	wire _w28112_ ;
	wire _w28113_ ;
	wire _w28114_ ;
	wire _w28115_ ;
	wire _w28116_ ;
	wire _w28117_ ;
	wire _w28118_ ;
	wire _w28119_ ;
	wire _w28120_ ;
	wire _w28121_ ;
	wire _w28122_ ;
	wire _w28123_ ;
	wire _w28124_ ;
	wire _w28125_ ;
	wire _w28126_ ;
	wire _w28127_ ;
	wire _w28128_ ;
	wire _w28129_ ;
	wire _w28130_ ;
	wire _w28131_ ;
	wire _w28132_ ;
	wire _w28133_ ;
	wire _w28134_ ;
	wire _w28135_ ;
	wire _w28136_ ;
	wire _w28137_ ;
	wire _w28138_ ;
	wire _w28139_ ;
	wire _w28140_ ;
	wire _w28141_ ;
	wire _w28142_ ;
	wire _w28143_ ;
	wire _w28144_ ;
	wire _w28145_ ;
	wire _w28146_ ;
	wire _w28147_ ;
	wire _w28148_ ;
	wire _w28149_ ;
	wire _w28150_ ;
	wire _w28151_ ;
	wire _w28152_ ;
	wire _w28153_ ;
	wire _w28154_ ;
	wire _w28155_ ;
	wire _w28156_ ;
	wire _w28157_ ;
	wire _w28158_ ;
	wire _w28159_ ;
	wire _w28160_ ;
	wire _w28161_ ;
	wire _w28162_ ;
	wire _w28163_ ;
	wire _w28164_ ;
	wire _w28165_ ;
	wire _w28166_ ;
	wire _w28167_ ;
	wire _w28168_ ;
	wire _w28169_ ;
	wire _w28170_ ;
	wire _w28171_ ;
	wire _w28172_ ;
	wire _w28173_ ;
	wire _w28174_ ;
	wire _w28175_ ;
	wire _w28176_ ;
	wire _w28177_ ;
	wire _w28178_ ;
	wire _w28179_ ;
	wire _w28180_ ;
	wire _w28181_ ;
	wire _w28182_ ;
	wire _w28183_ ;
	wire _w28184_ ;
	wire _w28185_ ;
	wire _w28186_ ;
	wire _w28187_ ;
	wire _w28188_ ;
	wire _w28189_ ;
	wire _w28190_ ;
	wire _w28191_ ;
	wire _w28192_ ;
	wire _w28193_ ;
	wire _w28194_ ;
	wire _w28195_ ;
	wire _w28196_ ;
	wire _w28197_ ;
	wire _w28198_ ;
	wire _w28199_ ;
	wire _w28200_ ;
	wire _w28201_ ;
	wire _w28202_ ;
	wire _w28203_ ;
	wire _w28204_ ;
	wire _w28205_ ;
	wire _w28206_ ;
	wire _w28207_ ;
	wire _w28208_ ;
	wire _w28209_ ;
	wire _w28210_ ;
	wire _w28211_ ;
	wire _w28212_ ;
	wire _w28213_ ;
	wire _w28214_ ;
	wire _w28215_ ;
	wire _w28216_ ;
	wire _w28217_ ;
	wire _w28218_ ;
	wire _w28219_ ;
	wire _w28220_ ;
	wire _w28221_ ;
	wire _w28222_ ;
	wire _w28223_ ;
	wire _w28224_ ;
	wire _w28225_ ;
	wire _w28226_ ;
	wire _w28227_ ;
	wire _w28228_ ;
	wire _w28229_ ;
	wire _w28230_ ;
	wire _w28231_ ;
	wire _w28232_ ;
	wire _w28233_ ;
	wire _w28234_ ;
	wire _w28235_ ;
	wire _w28236_ ;
	wire _w28237_ ;
	wire _w28238_ ;
	wire _w28239_ ;
	wire _w28240_ ;
	wire _w28241_ ;
	wire _w28242_ ;
	wire _w28243_ ;
	wire _w28244_ ;
	wire _w28245_ ;
	wire _w28246_ ;
	wire _w28247_ ;
	wire _w28248_ ;
	wire _w28249_ ;
	wire _w28250_ ;
	wire _w28251_ ;
	wire _w28252_ ;
	wire _w28253_ ;
	wire _w28254_ ;
	wire _w28255_ ;
	wire _w28256_ ;
	wire _w28257_ ;
	wire _w28258_ ;
	wire _w28259_ ;
	wire _w28260_ ;
	wire _w28261_ ;
	wire _w28262_ ;
	wire _w28263_ ;
	wire _w28264_ ;
	wire _w28265_ ;
	wire _w28266_ ;
	wire _w28267_ ;
	wire _w28268_ ;
	wire _w28269_ ;
	wire _w28270_ ;
	wire _w28271_ ;
	wire _w28272_ ;
	wire _w28273_ ;
	wire _w28274_ ;
	wire _w28275_ ;
	wire _w28276_ ;
	wire _w28277_ ;
	wire _w28278_ ;
	wire _w28279_ ;
	wire _w28280_ ;
	wire _w28281_ ;
	wire _w28282_ ;
	wire _w28283_ ;
	wire _w28284_ ;
	wire _w28285_ ;
	wire _w28286_ ;
	wire _w28287_ ;
	wire _w28288_ ;
	wire _w28289_ ;
	wire _w28290_ ;
	wire _w28291_ ;
	wire _w28292_ ;
	wire _w28293_ ;
	wire _w28294_ ;
	wire _w28295_ ;
	wire _w28296_ ;
	wire _w28297_ ;
	wire _w28298_ ;
	wire _w28299_ ;
	wire _w28300_ ;
	wire _w28301_ ;
	wire _w28302_ ;
	wire _w28303_ ;
	wire _w28304_ ;
	wire _w28305_ ;
	wire _w28306_ ;
	wire _w28307_ ;
	wire _w28308_ ;
	wire _w28309_ ;
	wire _w28310_ ;
	wire _w28311_ ;
	wire _w28312_ ;
	wire _w28313_ ;
	wire _w28314_ ;
	wire _w28315_ ;
	wire _w28316_ ;
	wire _w28317_ ;
	wire _w28318_ ;
	wire _w28319_ ;
	wire _w28320_ ;
	wire _w28321_ ;
	wire _w28322_ ;
	wire _w28323_ ;
	wire _w28324_ ;
	wire _w28325_ ;
	wire _w28326_ ;
	wire _w28327_ ;
	wire _w28328_ ;
	wire _w28329_ ;
	wire _w28330_ ;
	wire _w28331_ ;
	wire _w28332_ ;
	wire _w28333_ ;
	wire _w28334_ ;
	wire _w28335_ ;
	wire _w28336_ ;
	wire _w28337_ ;
	wire _w28338_ ;
	wire _w28339_ ;
	wire _w28340_ ;
	wire _w28341_ ;
	wire _w28342_ ;
	wire _w28343_ ;
	wire _w28344_ ;
	wire _w28345_ ;
	wire _w28346_ ;
	wire _w28347_ ;
	wire _w28348_ ;
	wire _w28349_ ;
	wire _w28350_ ;
	wire _w28351_ ;
	wire _w28352_ ;
	wire _w28353_ ;
	wire _w28354_ ;
	wire _w28355_ ;
	wire _w28356_ ;
	wire _w28357_ ;
	wire _w28358_ ;
	wire _w28359_ ;
	wire _w28360_ ;
	wire _w28361_ ;
	wire _w28362_ ;
	wire _w28363_ ;
	wire _w28364_ ;
	wire _w28365_ ;
	wire _w28366_ ;
	wire _w28367_ ;
	wire _w28368_ ;
	wire _w28369_ ;
	wire _w28370_ ;
	wire _w28371_ ;
	wire _w28372_ ;
	wire _w28373_ ;
	wire _w28374_ ;
	wire _w28375_ ;
	wire _w28376_ ;
	wire _w28377_ ;
	wire _w28378_ ;
	wire _w28379_ ;
	wire _w28380_ ;
	wire _w28381_ ;
	wire _w28382_ ;
	wire _w28383_ ;
	wire _w28384_ ;
	wire _w28385_ ;
	wire _w28386_ ;
	wire _w28387_ ;
	wire _w28388_ ;
	wire _w28389_ ;
	wire _w28390_ ;
	wire _w28391_ ;
	wire _w28392_ ;
	wire _w28393_ ;
	wire _w28394_ ;
	wire _w28395_ ;
	wire _w28396_ ;
	wire _w28397_ ;
	wire _w28398_ ;
	wire _w28399_ ;
	wire _w28400_ ;
	wire _w28401_ ;
	wire _w28402_ ;
	wire _w28403_ ;
	wire _w28404_ ;
	wire _w28405_ ;
	wire _w28406_ ;
	wire _w28407_ ;
	wire _w28408_ ;
	wire _w28409_ ;
	wire _w28410_ ;
	wire _w28411_ ;
	wire _w28412_ ;
	wire _w28413_ ;
	wire _w28414_ ;
	wire _w28415_ ;
	wire _w28416_ ;
	wire _w28417_ ;
	wire _w28418_ ;
	wire _w28419_ ;
	wire _w28420_ ;
	wire _w28421_ ;
	wire _w28422_ ;
	wire _w28423_ ;
	wire _w28424_ ;
	wire _w28425_ ;
	wire _w28426_ ;
	wire _w28427_ ;
	wire _w28428_ ;
	wire _w28429_ ;
	wire _w28430_ ;
	wire _w28431_ ;
	wire _w28432_ ;
	wire _w28433_ ;
	wire _w28434_ ;
	wire _w28435_ ;
	wire _w28436_ ;
	wire _w28437_ ;
	wire _w28438_ ;
	wire _w28439_ ;
	wire _w28440_ ;
	wire _w28441_ ;
	wire _w28442_ ;
	wire _w28443_ ;
	wire _w28444_ ;
	wire _w28445_ ;
	wire _w28446_ ;
	wire _w28447_ ;
	wire _w28448_ ;
	wire _w28449_ ;
	wire _w28450_ ;
	wire _w28451_ ;
	wire _w28452_ ;
	wire _w28453_ ;
	wire _w28454_ ;
	wire _w28455_ ;
	wire _w28456_ ;
	wire _w28457_ ;
	wire _w28458_ ;
	wire _w28459_ ;
	wire _w28460_ ;
	wire _w28461_ ;
	wire _w28462_ ;
	wire _w28463_ ;
	wire _w28464_ ;
	wire _w28465_ ;
	wire _w28466_ ;
	wire _w28467_ ;
	wire _w28468_ ;
	wire _w28469_ ;
	wire _w28470_ ;
	wire _w28471_ ;
	wire _w28472_ ;
	wire _w28473_ ;
	wire _w28474_ ;
	wire _w28475_ ;
	wire _w28476_ ;
	wire _w28477_ ;
	wire _w28478_ ;
	wire _w28479_ ;
	wire _w28480_ ;
	wire _w28481_ ;
	wire _w28482_ ;
	wire _w28483_ ;
	wire _w28484_ ;
	wire _w28485_ ;
	wire _w28486_ ;
	wire _w28487_ ;
	wire _w28488_ ;
	wire _w28489_ ;
	wire _w28490_ ;
	wire _w28491_ ;
	wire _w28492_ ;
	wire _w28493_ ;
	wire _w28494_ ;
	wire _w28495_ ;
	wire _w28496_ ;
	wire _w28497_ ;
	wire _w28498_ ;
	wire _w28499_ ;
	wire _w28500_ ;
	wire _w28501_ ;
	wire _w28502_ ;
	wire _w28503_ ;
	wire _w28504_ ;
	wire _w28505_ ;
	wire _w28506_ ;
	wire _w28507_ ;
	wire _w28508_ ;
	wire _w28509_ ;
	wire _w28510_ ;
	wire _w28511_ ;
	wire _w28512_ ;
	wire _w28513_ ;
	wire _w28514_ ;
	wire _w28515_ ;
	wire _w28516_ ;
	wire _w28517_ ;
	wire _w28518_ ;
	wire _w28519_ ;
	wire _w28520_ ;
	wire _w28521_ ;
	wire _w28522_ ;
	wire _w28523_ ;
	wire _w28524_ ;
	wire _w28525_ ;
	wire _w28526_ ;
	wire _w28527_ ;
	wire _w28528_ ;
	wire _w28529_ ;
	wire _w28530_ ;
	wire _w28531_ ;
	wire _w28532_ ;
	wire _w28533_ ;
	wire _w28534_ ;
	wire _w28535_ ;
	wire _w28536_ ;
	wire _w28537_ ;
	wire _w28538_ ;
	wire _w28539_ ;
	wire _w28540_ ;
	wire _w28541_ ;
	wire _w28542_ ;
	wire _w28543_ ;
	wire _w28544_ ;
	wire _w28545_ ;
	wire _w28546_ ;
	wire _w28547_ ;
	wire _w28548_ ;
	wire _w28549_ ;
	wire _w28550_ ;
	wire _w28551_ ;
	wire _w28552_ ;
	wire _w28553_ ;
	wire _w28554_ ;
	wire _w28555_ ;
	wire _w28556_ ;
	wire _w28557_ ;
	wire _w28558_ ;
	wire _w28559_ ;
	wire _w28560_ ;
	wire _w28561_ ;
	wire _w28562_ ;
	wire _w28563_ ;
	wire _w28564_ ;
	wire _w28565_ ;
	wire _w28566_ ;
	wire _w28567_ ;
	wire _w28568_ ;
	wire _w28569_ ;
	wire _w28570_ ;
	wire _w28571_ ;
	wire _w28572_ ;
	wire _w28573_ ;
	wire _w28574_ ;
	wire _w28575_ ;
	wire _w28576_ ;
	wire _w28577_ ;
	wire _w28578_ ;
	wire _w28579_ ;
	wire _w28580_ ;
	wire _w28581_ ;
	wire _w28582_ ;
	wire _w28583_ ;
	wire _w28584_ ;
	wire _w28585_ ;
	wire _w28586_ ;
	wire _w28587_ ;
	wire _w28588_ ;
	wire _w28589_ ;
	wire _w28590_ ;
	wire _w28591_ ;
	wire _w28592_ ;
	wire _w28593_ ;
	wire _w28594_ ;
	wire _w28595_ ;
	wire _w28596_ ;
	wire _w28597_ ;
	wire _w28598_ ;
	wire _w28599_ ;
	wire _w28600_ ;
	wire _w28601_ ;
	wire _w28602_ ;
	wire _w28603_ ;
	wire _w28604_ ;
	wire _w28605_ ;
	wire _w28606_ ;
	wire _w28607_ ;
	wire _w28608_ ;
	wire _w28609_ ;
	wire _w28610_ ;
	wire _w28611_ ;
	wire _w28612_ ;
	wire _w28613_ ;
	wire _w28614_ ;
	wire _w28615_ ;
	wire _w28616_ ;
	wire _w28617_ ;
	wire _w28618_ ;
	wire _w28619_ ;
	wire _w28620_ ;
	wire _w28621_ ;
	wire _w28622_ ;
	wire _w28623_ ;
	wire _w28624_ ;
	wire _w28625_ ;
	wire _w28626_ ;
	wire _w28627_ ;
	wire _w28628_ ;
	wire _w28629_ ;
	wire _w28630_ ;
	wire _w28631_ ;
	wire _w28632_ ;
	wire _w28633_ ;
	wire _w28634_ ;
	wire _w28635_ ;
	wire _w28636_ ;
	wire _w28637_ ;
	wire _w28638_ ;
	wire _w28639_ ;
	wire _w28640_ ;
	wire _w28641_ ;
	wire _w28642_ ;
	wire _w28643_ ;
	wire _w28644_ ;
	wire _w28645_ ;
	wire _w28646_ ;
	wire _w28647_ ;
	wire _w28648_ ;
	wire _w28649_ ;
	wire _w28650_ ;
	wire _w28651_ ;
	wire _w28652_ ;
	wire _w28653_ ;
	wire _w28654_ ;
	wire _w28655_ ;
	wire _w28656_ ;
	wire _w28657_ ;
	wire _w28658_ ;
	wire _w28659_ ;
	wire _w28660_ ;
	wire _w28661_ ;
	wire _w28662_ ;
	wire _w28663_ ;
	wire _w28664_ ;
	wire _w28665_ ;
	wire _w28666_ ;
	wire _w28667_ ;
	wire _w28668_ ;
	wire _w28669_ ;
	wire _w28670_ ;
	wire _w28671_ ;
	wire _w28672_ ;
	wire _w28673_ ;
	wire _w28674_ ;
	wire _w28675_ ;
	wire _w28676_ ;
	wire _w28677_ ;
	wire _w28678_ ;
	wire _w28679_ ;
	wire _w28680_ ;
	wire _w28681_ ;
	wire _w28682_ ;
	wire _w28683_ ;
	wire _w28684_ ;
	wire _w28685_ ;
	wire _w28686_ ;
	wire _w28687_ ;
	wire _w28688_ ;
	wire _w28689_ ;
	wire _w28690_ ;
	wire _w28691_ ;
	wire _w28692_ ;
	wire _w28693_ ;
	wire _w28694_ ;
	wire _w28695_ ;
	wire _w28696_ ;
	wire _w28697_ ;
	wire _w28698_ ;
	wire _w28699_ ;
	wire _w28700_ ;
	wire _w28701_ ;
	wire _w28702_ ;
	wire _w28703_ ;
	wire _w28704_ ;
	wire _w28705_ ;
	wire _w28706_ ;
	wire _w28707_ ;
	wire _w28708_ ;
	wire _w28709_ ;
	wire _w28710_ ;
	wire _w28711_ ;
	wire _w28712_ ;
	wire _w28713_ ;
	wire _w28714_ ;
	wire _w28715_ ;
	wire _w28716_ ;
	wire _w28717_ ;
	wire _w28718_ ;
	wire _w28719_ ;
	wire _w28720_ ;
	wire _w28721_ ;
	wire _w28722_ ;
	wire _w28723_ ;
	wire _w28724_ ;
	wire _w28725_ ;
	wire _w28726_ ;
	wire _w28727_ ;
	wire _w28728_ ;
	wire _w28729_ ;
	wire _w28730_ ;
	wire _w28731_ ;
	wire _w28732_ ;
	wire _w28733_ ;
	wire _w28734_ ;
	wire _w28735_ ;
	wire _w28736_ ;
	wire _w28737_ ;
	wire _w28738_ ;
	wire _w28739_ ;
	wire _w28740_ ;
	wire _w28741_ ;
	wire _w28742_ ;
	wire _w28743_ ;
	wire _w28744_ ;
	wire _w28745_ ;
	wire _w28746_ ;
	wire _w28747_ ;
	wire _w28748_ ;
	wire _w28749_ ;
	wire _w28750_ ;
	wire _w28751_ ;
	wire _w28752_ ;
	wire _w28753_ ;
	wire _w28754_ ;
	wire _w28755_ ;
	wire _w28756_ ;
	wire _w28757_ ;
	wire _w28758_ ;
	wire _w28759_ ;
	wire _w28760_ ;
	wire _w28761_ ;
	wire _w28762_ ;
	wire _w28763_ ;
	wire _w28764_ ;
	wire _w28765_ ;
	wire _w28766_ ;
	wire _w28767_ ;
	wire _w28768_ ;
	wire _w28769_ ;
	wire _w28770_ ;
	wire _w28771_ ;
	wire _w28772_ ;
	wire _w28773_ ;
	wire _w28774_ ;
	wire _w28775_ ;
	wire _w28776_ ;
	wire _w28777_ ;
	wire _w28778_ ;
	wire _w28779_ ;
	wire _w28780_ ;
	wire _w28781_ ;
	wire _w28782_ ;
	wire _w28783_ ;
	wire _w28784_ ;
	wire _w28785_ ;
	wire _w28786_ ;
	wire _w28787_ ;
	wire _w28788_ ;
	wire _w28789_ ;
	wire _w28790_ ;
	wire _w28791_ ;
	wire _w28792_ ;
	wire _w28793_ ;
	wire _w28794_ ;
	wire _w28795_ ;
	wire _w28796_ ;
	wire _w28797_ ;
	wire _w28798_ ;
	wire _w28799_ ;
	wire _w28800_ ;
	wire _w28801_ ;
	wire _w28802_ ;
	wire _w28803_ ;
	wire _w28804_ ;
	wire _w28805_ ;
	wire _w28806_ ;
	wire _w28807_ ;
	wire _w28808_ ;
	wire _w28809_ ;
	wire _w28810_ ;
	wire _w28811_ ;
	wire _w28812_ ;
	wire _w28813_ ;
	wire _w28814_ ;
	wire _w28815_ ;
	wire _w28816_ ;
	wire _w28817_ ;
	wire _w28818_ ;
	wire _w28819_ ;
	wire _w28820_ ;
	wire _w28821_ ;
	wire _w28822_ ;
	wire _w28823_ ;
	wire _w28824_ ;
	wire _w28825_ ;
	wire _w28826_ ;
	wire _w28827_ ;
	wire _w28828_ ;
	wire _w28829_ ;
	wire _w28830_ ;
	wire _w28831_ ;
	wire _w28832_ ;
	wire _w28833_ ;
	wire _w28834_ ;
	wire _w28835_ ;
	wire _w28836_ ;
	wire _w28837_ ;
	wire _w28838_ ;
	wire _w28839_ ;
	wire _w28840_ ;
	wire _w28841_ ;
	wire _w28842_ ;
	wire _w28843_ ;
	wire _w28844_ ;
	wire _w28845_ ;
	wire _w28846_ ;
	wire _w28847_ ;
	wire _w28848_ ;
	wire _w28849_ ;
	wire _w28850_ ;
	wire _w28851_ ;
	wire _w28852_ ;
	wire _w28853_ ;
	wire _w28854_ ;
	wire _w28855_ ;
	wire _w28856_ ;
	wire _w28857_ ;
	wire _w28858_ ;
	wire _w28859_ ;
	wire _w28860_ ;
	wire _w28861_ ;
	wire _w28862_ ;
	wire _w28863_ ;
	wire _w28864_ ;
	wire _w28865_ ;
	wire _w28866_ ;
	wire _w28867_ ;
	wire _w28868_ ;
	wire _w28869_ ;
	wire _w28870_ ;
	wire _w28871_ ;
	wire _w28872_ ;
	wire _w28873_ ;
	wire _w28874_ ;
	wire _w28875_ ;
	wire _w28876_ ;
	wire _w28877_ ;
	wire _w28878_ ;
	wire _w28879_ ;
	wire _w28880_ ;
	wire _w28881_ ;
	wire _w28882_ ;
	wire _w28883_ ;
	wire _w28884_ ;
	wire _w28885_ ;
	wire _w28886_ ;
	wire _w28887_ ;
	wire _w28888_ ;
	wire _w28889_ ;
	wire _w28890_ ;
	wire _w28891_ ;
	wire _w28892_ ;
	wire _w28893_ ;
	wire _w28894_ ;
	wire _w28895_ ;
	wire _w28896_ ;
	wire _w28897_ ;
	wire _w28898_ ;
	wire _w28899_ ;
	wire _w28900_ ;
	wire _w28901_ ;
	wire _w28902_ ;
	wire _w28903_ ;
	wire _w28904_ ;
	wire _w28905_ ;
	wire _w28906_ ;
	wire _w28907_ ;
	wire _w28908_ ;
	wire _w28909_ ;
	wire _w28910_ ;
	wire _w28911_ ;
	wire _w28912_ ;
	wire _w28913_ ;
	wire _w28914_ ;
	wire _w28915_ ;
	wire _w28916_ ;
	wire _w28917_ ;
	wire _w28918_ ;
	wire _w28919_ ;
	wire _w28920_ ;
	wire _w28921_ ;
	wire _w28922_ ;
	wire _w28923_ ;
	wire _w28924_ ;
	wire _w28925_ ;
	wire _w28926_ ;
	wire _w28927_ ;
	wire _w28928_ ;
	wire _w28929_ ;
	wire _w28930_ ;
	wire _w28931_ ;
	wire _w28932_ ;
	wire _w28933_ ;
	wire _w28934_ ;
	wire _w28935_ ;
	wire _w28936_ ;
	wire _w28937_ ;
	wire _w28938_ ;
	wire _w28939_ ;
	wire _w28940_ ;
	wire _w28941_ ;
	wire _w28942_ ;
	wire _w28943_ ;
	wire _w28944_ ;
	wire _w28945_ ;
	wire _w28946_ ;
	wire _w28947_ ;
	wire _w28948_ ;
	wire _w28949_ ;
	wire _w28950_ ;
	wire _w28951_ ;
	wire _w28952_ ;
	wire _w28953_ ;
	wire _w28954_ ;
	wire _w28955_ ;
	wire _w28956_ ;
	wire _w28957_ ;
	wire _w28958_ ;
	wire _w28959_ ;
	wire _w28960_ ;
	wire _w28961_ ;
	wire _w28962_ ;
	wire _w28963_ ;
	wire _w28964_ ;
	wire _w28965_ ;
	wire _w28966_ ;
	wire _w28967_ ;
	wire _w28968_ ;
	wire _w28969_ ;
	wire _w28970_ ;
	wire _w28971_ ;
	wire _w28972_ ;
	wire _w28973_ ;
	wire _w28974_ ;
	wire _w28975_ ;
	wire _w28976_ ;
	wire _w28977_ ;
	wire _w28978_ ;
	wire _w28979_ ;
	wire _w28980_ ;
	wire _w28981_ ;
	wire _w28982_ ;
	wire _w28983_ ;
	wire _w28984_ ;
	wire _w28985_ ;
	wire _w28986_ ;
	wire _w28987_ ;
	wire _w28988_ ;
	wire _w28989_ ;
	wire _w28990_ ;
	wire _w28991_ ;
	wire _w28992_ ;
	wire _w28993_ ;
	wire _w28994_ ;
	wire _w28995_ ;
	wire _w28996_ ;
	wire _w28997_ ;
	wire _w28998_ ;
	wire _w28999_ ;
	wire _w29000_ ;
	wire _w29001_ ;
	wire _w29002_ ;
	wire _w29003_ ;
	wire _w29004_ ;
	wire _w29005_ ;
	wire _w29006_ ;
	wire _w29007_ ;
	wire _w29008_ ;
	wire _w29009_ ;
	wire _w29010_ ;
	wire _w29011_ ;
	wire _w29012_ ;
	wire _w29013_ ;
	wire _w29014_ ;
	wire _w29015_ ;
	wire _w29016_ ;
	wire _w29017_ ;
	wire _w29018_ ;
	wire _w29019_ ;
	wire _w29020_ ;
	wire _w29021_ ;
	wire _w29022_ ;
	wire _w29023_ ;
	wire _w29024_ ;
	wire _w29025_ ;
	wire _w29026_ ;
	wire _w29027_ ;
	wire _w29028_ ;
	wire _w29029_ ;
	wire _w29030_ ;
	wire _w29031_ ;
	wire _w29032_ ;
	wire _w29033_ ;
	wire _w29034_ ;
	wire _w29035_ ;
	wire _w29036_ ;
	wire _w29037_ ;
	wire _w29038_ ;
	wire _w29039_ ;
	wire _w29040_ ;
	wire _w29041_ ;
	wire _w29042_ ;
	wire _w29043_ ;
	wire _w29044_ ;
	wire _w29045_ ;
	wire _w29046_ ;
	wire _w29047_ ;
	wire _w29048_ ;
	wire _w29049_ ;
	wire _w29050_ ;
	wire _w29051_ ;
	wire _w29052_ ;
	wire _w29053_ ;
	wire _w29054_ ;
	wire _w29055_ ;
	wire _w29056_ ;
	wire _w29057_ ;
	wire _w29058_ ;
	wire _w29059_ ;
	wire _w29060_ ;
	wire _w29061_ ;
	wire _w29062_ ;
	wire _w29063_ ;
	wire _w29064_ ;
	wire _w29065_ ;
	wire _w29066_ ;
	wire _w29067_ ;
	wire _w29068_ ;
	wire _w29069_ ;
	wire _w29070_ ;
	wire _w29071_ ;
	wire _w29072_ ;
	wire _w29073_ ;
	wire _w29074_ ;
	wire _w29075_ ;
	wire _w29076_ ;
	wire _w29077_ ;
	wire _w29078_ ;
	wire _w29079_ ;
	wire _w29080_ ;
	wire _w29081_ ;
	wire _w29082_ ;
	wire _w29083_ ;
	wire _w29084_ ;
	wire _w29085_ ;
	wire _w29086_ ;
	wire _w29087_ ;
	wire _w29088_ ;
	wire _w29089_ ;
	wire _w29090_ ;
	wire _w29091_ ;
	wire _w29092_ ;
	wire _w29093_ ;
	wire _w29094_ ;
	wire _w29095_ ;
	wire _w29096_ ;
	wire _w29097_ ;
	wire _w29098_ ;
	wire _w29099_ ;
	wire _w29100_ ;
	wire _w29101_ ;
	wire _w29102_ ;
	wire _w29103_ ;
	wire _w29104_ ;
	wire _w29105_ ;
	wire _w29106_ ;
	wire _w29107_ ;
	wire _w29108_ ;
	wire _w29109_ ;
	wire _w29110_ ;
	wire _w29111_ ;
	wire _w29112_ ;
	wire _w29113_ ;
	wire _w29114_ ;
	wire _w29115_ ;
	wire _w29116_ ;
	wire _w29117_ ;
	wire _w29118_ ;
	wire _w29119_ ;
	wire _w29120_ ;
	wire _w29121_ ;
	wire _w29122_ ;
	wire _w29123_ ;
	wire _w29124_ ;
	wire _w29125_ ;
	wire _w29126_ ;
	wire _w29127_ ;
	wire _w29128_ ;
	wire _w29129_ ;
	wire _w29130_ ;
	wire _w29131_ ;
	wire _w29132_ ;
	wire _w29133_ ;
	wire _w29134_ ;
	wire _w29135_ ;
	wire _w29136_ ;
	wire _w29137_ ;
	wire _w29138_ ;
	wire _w29139_ ;
	wire _w29140_ ;
	wire _w29141_ ;
	wire _w29142_ ;
	wire _w29143_ ;
	wire _w29144_ ;
	wire _w29145_ ;
	wire _w29146_ ;
	wire _w29147_ ;
	wire _w29148_ ;
	wire _w29149_ ;
	wire _w29150_ ;
	wire _w29151_ ;
	wire _w29152_ ;
	wire _w29153_ ;
	wire _w29154_ ;
	wire _w29155_ ;
	wire _w29156_ ;
	wire _w29157_ ;
	wire _w29158_ ;
	wire _w29159_ ;
	wire _w29160_ ;
	wire _w29161_ ;
	wire _w29162_ ;
	wire _w29163_ ;
	wire _w29164_ ;
	wire _w29165_ ;
	wire _w29166_ ;
	wire _w29167_ ;
	wire _w29168_ ;
	wire _w29169_ ;
	wire _w29170_ ;
	wire _w29171_ ;
	wire _w29172_ ;
	wire _w29173_ ;
	wire _w29174_ ;
	wire _w29175_ ;
	wire _w29176_ ;
	wire _w29177_ ;
	wire _w29178_ ;
	wire _w29179_ ;
	wire _w29180_ ;
	wire _w29181_ ;
	wire _w29182_ ;
	wire _w29183_ ;
	wire _w29184_ ;
	wire _w29185_ ;
	wire _w29186_ ;
	wire _w29187_ ;
	wire _w29188_ ;
	wire _w29189_ ;
	wire _w29190_ ;
	wire _w29191_ ;
	wire _w29192_ ;
	wire _w29193_ ;
	wire _w29194_ ;
	wire _w29195_ ;
	wire _w29196_ ;
	wire _w29197_ ;
	wire _w29198_ ;
	wire _w29199_ ;
	wire _w29200_ ;
	wire _w29201_ ;
	wire _w29202_ ;
	wire _w29203_ ;
	wire _w29204_ ;
	wire _w29205_ ;
	wire _w29206_ ;
	wire _w29207_ ;
	wire _w29208_ ;
	wire _w29209_ ;
	wire _w29210_ ;
	wire _w29211_ ;
	wire _w29212_ ;
	wire _w29213_ ;
	wire _w29214_ ;
	wire _w29215_ ;
	wire _w29216_ ;
	wire _w29217_ ;
	wire _w29218_ ;
	wire _w29219_ ;
	wire _w29220_ ;
	wire _w29221_ ;
	wire _w29222_ ;
	wire _w29223_ ;
	wire _w29224_ ;
	wire _w29225_ ;
	wire _w29226_ ;
	wire _w29227_ ;
	wire _w29228_ ;
	wire _w29229_ ;
	wire _w29230_ ;
	wire _w29231_ ;
	wire _w29232_ ;
	wire _w29233_ ;
	wire _w29234_ ;
	wire _w29235_ ;
	wire _w29236_ ;
	wire _w29237_ ;
	wire _w29238_ ;
	wire _w29239_ ;
	wire _w29240_ ;
	wire _w29241_ ;
	wire _w29242_ ;
	wire _w29243_ ;
	wire _w29244_ ;
	wire _w29245_ ;
	wire _w29246_ ;
	wire _w29247_ ;
	wire _w29248_ ;
	wire _w29249_ ;
	wire _w29250_ ;
	wire _w29251_ ;
	wire _w29252_ ;
	wire _w29253_ ;
	wire _w29254_ ;
	wire _w29255_ ;
	wire _w29256_ ;
	wire _w29257_ ;
	wire _w29258_ ;
	wire _w29259_ ;
	wire _w29260_ ;
	wire _w29261_ ;
	wire _w29262_ ;
	wire _w29263_ ;
	wire _w29264_ ;
	wire _w29265_ ;
	wire _w29266_ ;
	wire _w29267_ ;
	wire _w29268_ ;
	wire _w29269_ ;
	wire _w29270_ ;
	wire _w29271_ ;
	wire _w29272_ ;
	wire _w29273_ ;
	wire _w29274_ ;
	wire _w29275_ ;
	wire _w29276_ ;
	wire _w29277_ ;
	wire _w29278_ ;
	wire _w29279_ ;
	wire _w29280_ ;
	wire _w29281_ ;
	wire _w29282_ ;
	wire _w29283_ ;
	wire _w29284_ ;
	wire _w29285_ ;
	wire _w29286_ ;
	wire _w29287_ ;
	wire _w29288_ ;
	wire _w29289_ ;
	wire _w29290_ ;
	wire _w29291_ ;
	wire _w29292_ ;
	wire _w29293_ ;
	wire _w29294_ ;
	wire _w29295_ ;
	wire _w29296_ ;
	wire _w29297_ ;
	wire _w29298_ ;
	wire _w29299_ ;
	wire _w29300_ ;
	wire _w29301_ ;
	wire _w29302_ ;
	wire _w29303_ ;
	wire _w29304_ ;
	wire _w29305_ ;
	wire _w29306_ ;
	wire _w29307_ ;
	wire _w29308_ ;
	wire _w29309_ ;
	wire _w29310_ ;
	wire _w29311_ ;
	wire _w29312_ ;
	wire _w29313_ ;
	wire _w29314_ ;
	wire _w29315_ ;
	wire _w29316_ ;
	wire _w29317_ ;
	wire _w29318_ ;
	wire _w29319_ ;
	wire _w29320_ ;
	wire _w29321_ ;
	wire _w29322_ ;
	wire _w29323_ ;
	wire _w29324_ ;
	wire _w29325_ ;
	wire _w29326_ ;
	wire _w29327_ ;
	wire _w29328_ ;
	wire _w29329_ ;
	wire _w29330_ ;
	wire _w29331_ ;
	wire _w29332_ ;
	wire _w29333_ ;
	wire _w29334_ ;
	wire _w29335_ ;
	wire _w29336_ ;
	wire _w29337_ ;
	wire _w29338_ ;
	wire _w29339_ ;
	wire _w29340_ ;
	wire _w29341_ ;
	wire _w29342_ ;
	wire _w29343_ ;
	wire _w29344_ ;
	wire _w29345_ ;
	wire _w29346_ ;
	wire _w29347_ ;
	wire _w29348_ ;
	wire _w29349_ ;
	wire _w29350_ ;
	wire _w29351_ ;
	wire _w29352_ ;
	wire _w29353_ ;
	wire _w29354_ ;
	wire _w29355_ ;
	wire _w29356_ ;
	wire _w29357_ ;
	wire _w29358_ ;
	wire _w29359_ ;
	wire _w29360_ ;
	wire _w29361_ ;
	wire _w29362_ ;
	wire _w29363_ ;
	wire _w29364_ ;
	wire _w29365_ ;
	wire _w29366_ ;
	wire _w29367_ ;
	wire _w29368_ ;
	wire _w29369_ ;
	wire _w29370_ ;
	wire _w29371_ ;
	wire _w29372_ ;
	wire _w29373_ ;
	wire _w29374_ ;
	wire _w29375_ ;
	wire _w29376_ ;
	wire _w29377_ ;
	wire _w29378_ ;
	wire _w29379_ ;
	wire _w29380_ ;
	wire _w29381_ ;
	wire _w29382_ ;
	wire _w29383_ ;
	wire _w29384_ ;
	wire _w29385_ ;
	wire _w29386_ ;
	wire _w29387_ ;
	wire _w29388_ ;
	wire _w29389_ ;
	wire _w29390_ ;
	wire _w29391_ ;
	wire _w29392_ ;
	wire _w29393_ ;
	wire _w29394_ ;
	wire _w29395_ ;
	wire _w29396_ ;
	wire _w29397_ ;
	wire _w29398_ ;
	wire _w29399_ ;
	wire _w29400_ ;
	wire _w29401_ ;
	wire _w29402_ ;
	wire _w29403_ ;
	wire _w29404_ ;
	wire _w29405_ ;
	wire _w29406_ ;
	wire _w29407_ ;
	wire _w29408_ ;
	wire _w29409_ ;
	wire _w29410_ ;
	wire _w29411_ ;
	wire _w29412_ ;
	wire _w29413_ ;
	wire _w29414_ ;
	wire _w29415_ ;
	wire _w29416_ ;
	wire _w29417_ ;
	wire _w29418_ ;
	wire _w29419_ ;
	wire _w29420_ ;
	wire _w29421_ ;
	wire _w29422_ ;
	wire _w29423_ ;
	wire _w29424_ ;
	wire _w29425_ ;
	wire _w29426_ ;
	wire _w29427_ ;
	wire _w29428_ ;
	wire _w29429_ ;
	wire _w29430_ ;
	wire _w29431_ ;
	wire _w29432_ ;
	wire _w29433_ ;
	wire _w29434_ ;
	wire _w29435_ ;
	wire _w29436_ ;
	wire _w29437_ ;
	wire _w29438_ ;
	wire _w29439_ ;
	wire _w29440_ ;
	wire _w29441_ ;
	wire _w29442_ ;
	wire _w29443_ ;
	wire _w29444_ ;
	wire _w29445_ ;
	wire _w29446_ ;
	wire _w29447_ ;
	wire _w29448_ ;
	wire _w29449_ ;
	wire _w29450_ ;
	wire _w29451_ ;
	wire _w29452_ ;
	wire _w29453_ ;
	wire _w29454_ ;
	wire _w29455_ ;
	wire _w29456_ ;
	wire _w29457_ ;
	wire _w29458_ ;
	wire _w29459_ ;
	wire _w29460_ ;
	wire _w29461_ ;
	wire _w29462_ ;
	wire _w29463_ ;
	wire _w29464_ ;
	wire _w29465_ ;
	wire _w29466_ ;
	wire _w29467_ ;
	wire _w29468_ ;
	wire _w29469_ ;
	wire _w29470_ ;
	wire _w29471_ ;
	wire _w29472_ ;
	wire _w29473_ ;
	wire _w29474_ ;
	wire _w29475_ ;
	wire _w29476_ ;
	wire _w29477_ ;
	wire _w29478_ ;
	wire _w29479_ ;
	wire _w29480_ ;
	wire _w29481_ ;
	wire _w29482_ ;
	wire _w29483_ ;
	wire _w29484_ ;
	wire _w29485_ ;
	wire _w29486_ ;
	wire _w29487_ ;
	wire _w29488_ ;
	wire _w29489_ ;
	wire _w29490_ ;
	wire _w29491_ ;
	wire _w29492_ ;
	wire _w29493_ ;
	wire _w29494_ ;
	wire _w29495_ ;
	wire _w29496_ ;
	wire _w29497_ ;
	wire _w29498_ ;
	wire _w29499_ ;
	wire _w29500_ ;
	wire _w29501_ ;
	wire _w29502_ ;
	wire _w29503_ ;
	wire _w29504_ ;
	wire _w29505_ ;
	wire _w29506_ ;
	wire _w29507_ ;
	wire _w29508_ ;
	wire _w29509_ ;
	wire _w29510_ ;
	wire _w29511_ ;
	wire _w29512_ ;
	wire _w29513_ ;
	wire _w29514_ ;
	wire _w29515_ ;
	wire _w29516_ ;
	wire _w29517_ ;
	wire _w29518_ ;
	wire _w29519_ ;
	wire _w29520_ ;
	wire _w29521_ ;
	wire _w29522_ ;
	wire _w29523_ ;
	wire _w29524_ ;
	wire _w29525_ ;
	wire _w29526_ ;
	wire _w29527_ ;
	wire _w29528_ ;
	wire _w29529_ ;
	wire _w29530_ ;
	wire _w29531_ ;
	wire _w29532_ ;
	wire _w29533_ ;
	wire _w29534_ ;
	wire _w29535_ ;
	wire _w29536_ ;
	wire _w29537_ ;
	wire _w29538_ ;
	wire _w29539_ ;
	wire _w29540_ ;
	wire _w29541_ ;
	wire _w29542_ ;
	wire _w29543_ ;
	wire _w29544_ ;
	wire _w29545_ ;
	wire _w29546_ ;
	wire _w29547_ ;
	wire _w29548_ ;
	wire _w29549_ ;
	wire _w29550_ ;
	wire _w29551_ ;
	wire _w29552_ ;
	wire _w29553_ ;
	wire _w29554_ ;
	wire _w29555_ ;
	wire _w29556_ ;
	wire _w29557_ ;
	wire _w29558_ ;
	wire _w29559_ ;
	wire _w29560_ ;
	wire _w29561_ ;
	wire _w29562_ ;
	wire _w29563_ ;
	wire _w29564_ ;
	wire _w29565_ ;
	wire _w29566_ ;
	wire _w29567_ ;
	wire _w29568_ ;
	wire _w29569_ ;
	wire _w29570_ ;
	wire _w29571_ ;
	wire _w29572_ ;
	wire _w29573_ ;
	wire _w29574_ ;
	wire _w29575_ ;
	wire _w29576_ ;
	wire _w29577_ ;
	wire _w29578_ ;
	wire _w29579_ ;
	wire _w29580_ ;
	wire _w29581_ ;
	wire _w29582_ ;
	wire _w29583_ ;
	wire _w29584_ ;
	wire _w29585_ ;
	wire _w29586_ ;
	wire _w29587_ ;
	wire _w29588_ ;
	wire _w29589_ ;
	wire _w29590_ ;
	wire _w29591_ ;
	wire _w29592_ ;
	wire _w29593_ ;
	wire _w29594_ ;
	wire _w29595_ ;
	wire _w29596_ ;
	wire _w29597_ ;
	wire _w29598_ ;
	wire _w29599_ ;
	wire _w29600_ ;
	wire _w29601_ ;
	wire _w29602_ ;
	wire _w29603_ ;
	wire _w29604_ ;
	wire _w29605_ ;
	wire _w29606_ ;
	wire _w29607_ ;
	wire _w29608_ ;
	wire _w29609_ ;
	wire _w29610_ ;
	wire _w29611_ ;
	wire _w29612_ ;
	wire _w29613_ ;
	wire _w29614_ ;
	wire _w29615_ ;
	wire _w29616_ ;
	wire _w29617_ ;
	wire _w29618_ ;
	wire _w29619_ ;
	wire _w29620_ ;
	wire _w29621_ ;
	wire _w29622_ ;
	wire _w29623_ ;
	wire _w29624_ ;
	wire _w29625_ ;
	wire _w29626_ ;
	wire _w29627_ ;
	wire _w29628_ ;
	wire _w29629_ ;
	wire _w29630_ ;
	wire _w29631_ ;
	wire _w29632_ ;
	wire _w29633_ ;
	wire _w29634_ ;
	wire _w29635_ ;
	wire _w29636_ ;
	wire _w29637_ ;
	wire _w29638_ ;
	wire _w29639_ ;
	wire _w29640_ ;
	wire _w29641_ ;
	wire _w29642_ ;
	wire _w29643_ ;
	wire _w29644_ ;
	wire _w29645_ ;
	wire _w29646_ ;
	wire _w29647_ ;
	wire _w29648_ ;
	wire _w29649_ ;
	wire _w29650_ ;
	wire _w29651_ ;
	wire _w29652_ ;
	wire _w29653_ ;
	wire _w29654_ ;
	wire _w29655_ ;
	wire _w29656_ ;
	wire _w29657_ ;
	wire _w29658_ ;
	wire _w29659_ ;
	wire _w29660_ ;
	wire _w29661_ ;
	wire _w29662_ ;
	wire _w29663_ ;
	wire _w29664_ ;
	wire _w29665_ ;
	wire _w29666_ ;
	wire _w29667_ ;
	wire _w29668_ ;
	wire _w29669_ ;
	wire _w29670_ ;
	wire _w29671_ ;
	wire _w29672_ ;
	wire _w29673_ ;
	wire _w29674_ ;
	wire _w29675_ ;
	wire _w29676_ ;
	wire _w29677_ ;
	wire _w29678_ ;
	wire _w29679_ ;
	wire _w29680_ ;
	wire _w29681_ ;
	wire _w29682_ ;
	wire _w29683_ ;
	wire _w29684_ ;
	wire _w29685_ ;
	wire _w29686_ ;
	wire _w29687_ ;
	wire _w29688_ ;
	wire _w29689_ ;
	wire _w29690_ ;
	wire _w29691_ ;
	wire _w29692_ ;
	wire _w29693_ ;
	wire _w29694_ ;
	wire _w29695_ ;
	wire _w29696_ ;
	wire _w29697_ ;
	wire _w29698_ ;
	wire _w29699_ ;
	wire _w29700_ ;
	wire _w29701_ ;
	wire _w29702_ ;
	wire _w29703_ ;
	wire _w29704_ ;
	wire _w29705_ ;
	wire _w29706_ ;
	wire _w29707_ ;
	wire _w29708_ ;
	wire _w29709_ ;
	wire _w29710_ ;
	wire _w29711_ ;
	wire _w29712_ ;
	wire _w29713_ ;
	wire _w29714_ ;
	wire _w29715_ ;
	wire _w29716_ ;
	wire _w29717_ ;
	wire _w29718_ ;
	wire _w29719_ ;
	wire _w29720_ ;
	wire _w29721_ ;
	wire _w29722_ ;
	wire _w29723_ ;
	wire _w29724_ ;
	wire _w29725_ ;
	wire _w29726_ ;
	wire _w29727_ ;
	wire _w29728_ ;
	wire _w29729_ ;
	wire _w29730_ ;
	wire _w29731_ ;
	wire _w29732_ ;
	wire _w29733_ ;
	wire _w29734_ ;
	wire _w29735_ ;
	wire _w29736_ ;
	wire _w29737_ ;
	wire _w29738_ ;
	wire _w29739_ ;
	wire _w29740_ ;
	wire _w29741_ ;
	wire _w29742_ ;
	wire _w29743_ ;
	wire _w29744_ ;
	wire _w29745_ ;
	wire _w29746_ ;
	wire _w29747_ ;
	wire _w29748_ ;
	wire _w29749_ ;
	wire _w29750_ ;
	wire _w29751_ ;
	wire _w29752_ ;
	wire _w29753_ ;
	wire _w29754_ ;
	wire _w29755_ ;
	wire _w29756_ ;
	wire _w29757_ ;
	wire _w29758_ ;
	wire _w29759_ ;
	wire _w29760_ ;
	wire _w29761_ ;
	wire _w29762_ ;
	wire _w29763_ ;
	wire _w29764_ ;
	wire _w29765_ ;
	wire _w29766_ ;
	wire _w29767_ ;
	wire _w29768_ ;
	wire _w29769_ ;
	wire _w29770_ ;
	wire _w29771_ ;
	wire _w29772_ ;
	wire _w29773_ ;
	wire _w29774_ ;
	wire _w29775_ ;
	wire _w29776_ ;
	wire _w29777_ ;
	wire _w29778_ ;
	wire _w29779_ ;
	wire _w29780_ ;
	wire _w29781_ ;
	wire _w29782_ ;
	wire _w29783_ ;
	wire _w29784_ ;
	wire _w29785_ ;
	wire _w29786_ ;
	wire _w29787_ ;
	wire _w29788_ ;
	wire _w29789_ ;
	wire _w29790_ ;
	wire _w29791_ ;
	wire _w29792_ ;
	wire _w29793_ ;
	wire _w29794_ ;
	wire _w29795_ ;
	wire _w29796_ ;
	wire _w29797_ ;
	wire _w29798_ ;
	wire _w29799_ ;
	wire _w29800_ ;
	wire _w29801_ ;
	wire _w29802_ ;
	wire _w29803_ ;
	wire _w29804_ ;
	wire _w29805_ ;
	wire _w29806_ ;
	wire _w29807_ ;
	wire _w29808_ ;
	wire _w29809_ ;
	wire _w29810_ ;
	wire _w29811_ ;
	wire _w29812_ ;
	wire _w29813_ ;
	wire _w29814_ ;
	wire _w29815_ ;
	wire _w29816_ ;
	wire _w29817_ ;
	wire _w29818_ ;
	wire _w29819_ ;
	wire _w29820_ ;
	wire _w29821_ ;
	wire _w29822_ ;
	wire _w29823_ ;
	wire _w29824_ ;
	wire _w29825_ ;
	wire _w29826_ ;
	wire _w29827_ ;
	wire _w29828_ ;
	wire _w29829_ ;
	wire _w29830_ ;
	wire _w29831_ ;
	wire _w29832_ ;
	wire _w29833_ ;
	wire _w29834_ ;
	wire _w29835_ ;
	wire _w29836_ ;
	wire _w29837_ ;
	wire _w29838_ ;
	wire _w29839_ ;
	wire _w29840_ ;
	wire _w29841_ ;
	wire _w29842_ ;
	wire _w29843_ ;
	wire _w29844_ ;
	wire _w29845_ ;
	wire _w29846_ ;
	wire _w29847_ ;
	wire _w29848_ ;
	wire _w29849_ ;
	wire _w29850_ ;
	wire _w29851_ ;
	wire _w29852_ ;
	wire _w29853_ ;
	wire _w29854_ ;
	wire _w29855_ ;
	wire _w29856_ ;
	wire _w29857_ ;
	wire _w29858_ ;
	wire _w29859_ ;
	wire _w29860_ ;
	wire _w29861_ ;
	wire _w29862_ ;
	wire _w29863_ ;
	wire _w29864_ ;
	wire _w29865_ ;
	wire _w29866_ ;
	wire _w29867_ ;
	wire _w29868_ ;
	wire _w29869_ ;
	wire _w29870_ ;
	wire _w29871_ ;
	wire _w29872_ ;
	wire _w29873_ ;
	wire _w29874_ ;
	wire _w29875_ ;
	wire _w29876_ ;
	wire _w29877_ ;
	wire _w29878_ ;
	wire _w29879_ ;
	wire _w29880_ ;
	wire _w29881_ ;
	wire _w29882_ ;
	wire _w29883_ ;
	wire _w29884_ ;
	wire _w29885_ ;
	wire _w29886_ ;
	wire _w29887_ ;
	wire _w29888_ ;
	wire _w29889_ ;
	wire _w29890_ ;
	wire _w29891_ ;
	wire _w29892_ ;
	wire _w29893_ ;
	wire _w29894_ ;
	wire _w29895_ ;
	wire _w29896_ ;
	wire _w29897_ ;
	wire _w29898_ ;
	wire _w29899_ ;
	wire _w29900_ ;
	wire _w29901_ ;
	wire _w29902_ ;
	wire _w29903_ ;
	wire _w29904_ ;
	wire _w29905_ ;
	wire _w29906_ ;
	wire _w29907_ ;
	wire _w29908_ ;
	wire _w29909_ ;
	wire _w29910_ ;
	wire _w29911_ ;
	wire _w29912_ ;
	wire _w29913_ ;
	wire _w29914_ ;
	wire _w29915_ ;
	wire _w29916_ ;
	wire _w29917_ ;
	wire _w29918_ ;
	wire _w29919_ ;
	wire _w29920_ ;
	wire _w29921_ ;
	wire _w29922_ ;
	wire _w29923_ ;
	wire _w29924_ ;
	wire _w29925_ ;
	wire _w29926_ ;
	wire _w29927_ ;
	wire _w29928_ ;
	wire _w29929_ ;
	wire _w29930_ ;
	wire _w29931_ ;
	wire _w29932_ ;
	wire _w29933_ ;
	wire _w29934_ ;
	wire _w29935_ ;
	wire _w29936_ ;
	wire _w29937_ ;
	wire _w29938_ ;
	wire _w29939_ ;
	wire _w29940_ ;
	wire _w29941_ ;
	wire _w29942_ ;
	wire _w29943_ ;
	wire _w29944_ ;
	wire _w29945_ ;
	wire _w29946_ ;
	wire _w29947_ ;
	wire _w29948_ ;
	wire _w29949_ ;
	wire _w29950_ ;
	wire _w29951_ ;
	wire _w29952_ ;
	wire _w29953_ ;
	wire _w29954_ ;
	wire _w29955_ ;
	wire _w29956_ ;
	wire _w29957_ ;
	wire _w29958_ ;
	wire _w29959_ ;
	wire _w29960_ ;
	wire _w29961_ ;
	wire _w29962_ ;
	wire _w29963_ ;
	wire _w29964_ ;
	wire _w29965_ ;
	wire _w29966_ ;
	wire _w29967_ ;
	wire _w29968_ ;
	wire _w29969_ ;
	wire _w29970_ ;
	wire _w29971_ ;
	wire _w29972_ ;
	wire _w29973_ ;
	wire _w29974_ ;
	wire _w29975_ ;
	wire _w29976_ ;
	wire _w29977_ ;
	wire _w29978_ ;
	wire _w29979_ ;
	wire _w29980_ ;
	wire _w29981_ ;
	wire _w29982_ ;
	wire _w29983_ ;
	wire _w29984_ ;
	wire _w29985_ ;
	wire _w29986_ ;
	wire _w29987_ ;
	wire _w29988_ ;
	wire _w29989_ ;
	wire _w29990_ ;
	wire _w29991_ ;
	wire _w29992_ ;
	wire _w29993_ ;
	wire _w29994_ ;
	wire _w29995_ ;
	wire _w29996_ ;
	wire _w29997_ ;
	wire _w29998_ ;
	wire _w29999_ ;
	wire _w30000_ ;
	wire _w30001_ ;
	wire _w30002_ ;
	wire _w30003_ ;
	wire _w30004_ ;
	wire _w30005_ ;
	wire _w30006_ ;
	wire _w30007_ ;
	wire _w30008_ ;
	wire _w30009_ ;
	wire _w30010_ ;
	wire _w30011_ ;
	wire _w30012_ ;
	wire _w30013_ ;
	wire _w30014_ ;
	wire _w30015_ ;
	wire _w30016_ ;
	wire _w30017_ ;
	wire _w30018_ ;
	wire _w30019_ ;
	wire _w30020_ ;
	wire _w30021_ ;
	wire _w30022_ ;
	wire _w30023_ ;
	wire _w30024_ ;
	wire _w30025_ ;
	wire _w30026_ ;
	wire _w30027_ ;
	wire _w30028_ ;
	wire _w30029_ ;
	wire _w30030_ ;
	wire _w30031_ ;
	wire _w30032_ ;
	wire _w30033_ ;
	wire _w30034_ ;
	wire _w30035_ ;
	wire _w30036_ ;
	wire _w30037_ ;
	wire _w30038_ ;
	wire _w30039_ ;
	wire _w30040_ ;
	wire _w30041_ ;
	wire _w30042_ ;
	wire _w30043_ ;
	wire _w30044_ ;
	wire _w30045_ ;
	wire _w30046_ ;
	wire _w30047_ ;
	wire _w30048_ ;
	wire _w30049_ ;
	wire _w30050_ ;
	wire _w30051_ ;
	wire _w30052_ ;
	wire _w30053_ ;
	wire _w30054_ ;
	wire _w30055_ ;
	wire _w30056_ ;
	wire _w30057_ ;
	wire _w30058_ ;
	wire _w30059_ ;
	wire _w30060_ ;
	wire _w30061_ ;
	wire _w30062_ ;
	wire _w30063_ ;
	wire _w30064_ ;
	wire _w30065_ ;
	wire _w30066_ ;
	wire _w30067_ ;
	wire _w30068_ ;
	wire _w30069_ ;
	wire _w30070_ ;
	wire _w30071_ ;
	wire _w30072_ ;
	wire _w30073_ ;
	wire _w30074_ ;
	wire _w30075_ ;
	wire _w30076_ ;
	wire _w30077_ ;
	wire _w30078_ ;
	wire _w30079_ ;
	wire _w30080_ ;
	wire _w30081_ ;
	wire _w30082_ ;
	wire _w30083_ ;
	wire _w30084_ ;
	wire _w30085_ ;
	wire _w30086_ ;
	wire _w30087_ ;
	wire _w30088_ ;
	wire _w30089_ ;
	wire _w30090_ ;
	wire _w30091_ ;
	wire _w30092_ ;
	wire _w30093_ ;
	wire _w30094_ ;
	wire _w30095_ ;
	wire _w30096_ ;
	wire _w30097_ ;
	wire _w30098_ ;
	wire _w30099_ ;
	wire _w30100_ ;
	wire _w30101_ ;
	wire _w30102_ ;
	wire _w30103_ ;
	wire _w30104_ ;
	wire _w30105_ ;
	wire _w30106_ ;
	wire _w30107_ ;
	wire _w30108_ ;
	wire _w30109_ ;
	wire _w30110_ ;
	wire _w30111_ ;
	wire _w30112_ ;
	wire _w30113_ ;
	wire _w30114_ ;
	wire _w30115_ ;
	wire _w30116_ ;
	wire _w30117_ ;
	wire _w30118_ ;
	wire _w30119_ ;
	wire _w30120_ ;
	wire _w30121_ ;
	wire _w30122_ ;
	wire _w30123_ ;
	wire _w30124_ ;
	wire _w30125_ ;
	wire _w30126_ ;
	wire _w30127_ ;
	wire _w30128_ ;
	wire _w30129_ ;
	wire _w30130_ ;
	wire _w30131_ ;
	wire _w30132_ ;
	wire _w30133_ ;
	wire _w30134_ ;
	wire _w30135_ ;
	wire _w30136_ ;
	wire _w30137_ ;
	wire _w30138_ ;
	wire _w30139_ ;
	wire _w30140_ ;
	wire _w30141_ ;
	wire _w30142_ ;
	wire _w30143_ ;
	wire _w30144_ ;
	wire _w30145_ ;
	wire _w30146_ ;
	wire _w30147_ ;
	wire _w30148_ ;
	wire _w30149_ ;
	wire _w30150_ ;
	wire _w30151_ ;
	wire _w30152_ ;
	wire _w30153_ ;
	wire _w30154_ ;
	wire _w30155_ ;
	wire _w30156_ ;
	wire _w30157_ ;
	wire _w30158_ ;
	wire _w30159_ ;
	wire _w30160_ ;
	wire _w30161_ ;
	wire _w30162_ ;
	wire _w30163_ ;
	wire _w30164_ ;
	wire _w30165_ ;
	wire _w30166_ ;
	wire _w30167_ ;
	wire _w30168_ ;
	wire _w30169_ ;
	wire _w30170_ ;
	wire _w30171_ ;
	wire _w30172_ ;
	wire _w30173_ ;
	wire _w30174_ ;
	wire _w30175_ ;
	wire _w30176_ ;
	wire _w30177_ ;
	wire _w30178_ ;
	wire _w30179_ ;
	wire _w30180_ ;
	wire _w30181_ ;
	wire _w30182_ ;
	wire _w30183_ ;
	wire _w30184_ ;
	wire _w30185_ ;
	wire _w30186_ ;
	wire _w30187_ ;
	wire _w30188_ ;
	wire _w30189_ ;
	wire _w30190_ ;
	wire _w30191_ ;
	wire _w30192_ ;
	wire _w30193_ ;
	wire _w30194_ ;
	wire _w30195_ ;
	wire _w30196_ ;
	wire _w30197_ ;
	wire _w30198_ ;
	wire _w30199_ ;
	wire _w30200_ ;
	wire _w30201_ ;
	wire _w30202_ ;
	wire _w30203_ ;
	wire _w30204_ ;
	wire _w30205_ ;
	wire _w30206_ ;
	wire _w30207_ ;
	wire _w30208_ ;
	wire _w30209_ ;
	wire _w30210_ ;
	wire _w30211_ ;
	wire _w30212_ ;
	wire _w30213_ ;
	wire _w30214_ ;
	wire _w30215_ ;
	wire _w30216_ ;
	wire _w30217_ ;
	wire _w30218_ ;
	wire _w30219_ ;
	wire _w30220_ ;
	wire _w30221_ ;
	wire _w30222_ ;
	wire _w30223_ ;
	wire _w30224_ ;
	wire _w30225_ ;
	wire _w30226_ ;
	wire _w30227_ ;
	wire _w30228_ ;
	wire _w30229_ ;
	wire _w30230_ ;
	wire _w30231_ ;
	wire _w30232_ ;
	wire _w30233_ ;
	wire _w30234_ ;
	wire _w30235_ ;
	wire _w30236_ ;
	wire _w30237_ ;
	wire _w30238_ ;
	wire _w30239_ ;
	wire _w30240_ ;
	wire _w30241_ ;
	wire _w30242_ ;
	wire _w30243_ ;
	wire _w30244_ ;
	wire _w30245_ ;
	wire _w30246_ ;
	wire _w30247_ ;
	wire _w30248_ ;
	wire _w30249_ ;
	wire _w30250_ ;
	wire _w30251_ ;
	wire _w30252_ ;
	wire _w30253_ ;
	wire _w30254_ ;
	wire _w30255_ ;
	wire _w30256_ ;
	wire _w30257_ ;
	wire _w30258_ ;
	wire _w30259_ ;
	wire _w30260_ ;
	wire _w30261_ ;
	wire _w30262_ ;
	wire _w30263_ ;
	wire _w30264_ ;
	wire _w30265_ ;
	wire _w30266_ ;
	wire _w30267_ ;
	wire _w30268_ ;
	wire _w30269_ ;
	wire _w30270_ ;
	wire _w30271_ ;
	wire _w30272_ ;
	wire _w30273_ ;
	wire _w30274_ ;
	wire _w30275_ ;
	wire _w30276_ ;
	wire _w30277_ ;
	wire _w30278_ ;
	wire _w30279_ ;
	wire _w30280_ ;
	wire _w30281_ ;
	wire _w30282_ ;
	wire _w30283_ ;
	wire _w30284_ ;
	wire _w30285_ ;
	wire _w30286_ ;
	wire _w30287_ ;
	wire _w30288_ ;
	wire _w30289_ ;
	wire _w30290_ ;
	wire _w30291_ ;
	wire _w30292_ ;
	wire _w30293_ ;
	wire _w30294_ ;
	wire _w30295_ ;
	wire _w30296_ ;
	wire _w30297_ ;
	wire _w30298_ ;
	wire _w30299_ ;
	wire _w30300_ ;
	wire _w30301_ ;
	wire _w30302_ ;
	wire _w30303_ ;
	wire _w30304_ ;
	wire _w30305_ ;
	wire _w30306_ ;
	wire _w30307_ ;
	wire _w30308_ ;
	wire _w30309_ ;
	wire _w30310_ ;
	wire _w30311_ ;
	wire _w30312_ ;
	wire _w30313_ ;
	wire _w30314_ ;
	wire _w30315_ ;
	wire _w30316_ ;
	wire _w30317_ ;
	wire _w30318_ ;
	wire _w30319_ ;
	wire _w30320_ ;
	wire _w30321_ ;
	wire _w30322_ ;
	wire _w30323_ ;
	wire _w30324_ ;
	wire _w30325_ ;
	wire _w30326_ ;
	wire _w30327_ ;
	wire _w30328_ ;
	wire _w30329_ ;
	wire _w30330_ ;
	wire _w30331_ ;
	wire _w30332_ ;
	wire _w30333_ ;
	wire _w30334_ ;
	wire _w30335_ ;
	wire _w30336_ ;
	wire _w30337_ ;
	wire _w30338_ ;
	wire _w30339_ ;
	wire _w30340_ ;
	wire _w30341_ ;
	wire _w30342_ ;
	wire _w30343_ ;
	wire _w30344_ ;
	wire _w30345_ ;
	wire _w30346_ ;
	wire _w30347_ ;
	wire _w30348_ ;
	wire _w30349_ ;
	wire _w30350_ ;
	wire _w30351_ ;
	wire _w30352_ ;
	wire _w30353_ ;
	wire _w30354_ ;
	wire _w30355_ ;
	wire _w30356_ ;
	wire _w30357_ ;
	wire _w30358_ ;
	wire _w30359_ ;
	wire _w30360_ ;
	wire _w30361_ ;
	wire _w30362_ ;
	wire _w30363_ ;
	wire _w30364_ ;
	wire _w30365_ ;
	wire _w30366_ ;
	wire _w30367_ ;
	wire _w30368_ ;
	wire _w30369_ ;
	wire _w30370_ ;
	wire _w30371_ ;
	wire _w30372_ ;
	wire _w30373_ ;
	wire _w30374_ ;
	wire _w30375_ ;
	wire _w30376_ ;
	wire _w30377_ ;
	wire _w30378_ ;
	wire _w30379_ ;
	wire _w30380_ ;
	wire _w30381_ ;
	wire _w30382_ ;
	wire _w30383_ ;
	wire _w30384_ ;
	wire _w30385_ ;
	wire _w30386_ ;
	wire _w30387_ ;
	wire _w30388_ ;
	wire _w30389_ ;
	wire _w30390_ ;
	wire _w30391_ ;
	wire _w30392_ ;
	wire _w30393_ ;
	wire _w30394_ ;
	wire _w30395_ ;
	wire _w30396_ ;
	wire _w30397_ ;
	wire _w30398_ ;
	wire _w30399_ ;
	wire _w30400_ ;
	wire _w30401_ ;
	wire _w30402_ ;
	wire _w30403_ ;
	wire _w30404_ ;
	wire _w30405_ ;
	wire _w30406_ ;
	wire _w30407_ ;
	wire _w30408_ ;
	wire _w30409_ ;
	wire _w30410_ ;
	wire _w30411_ ;
	wire _w30412_ ;
	wire _w30413_ ;
	wire _w30414_ ;
	wire _w30415_ ;
	wire _w30416_ ;
	wire _w30417_ ;
	wire _w30418_ ;
	wire _w30419_ ;
	wire _w30420_ ;
	wire _w30421_ ;
	wire _w30422_ ;
	wire _w30423_ ;
	wire _w30424_ ;
	wire _w30425_ ;
	wire _w30426_ ;
	wire _w30427_ ;
	wire _w30428_ ;
	wire _w30429_ ;
	wire _w30430_ ;
	wire _w30431_ ;
	wire _w30432_ ;
	wire _w30433_ ;
	wire _w30434_ ;
	wire _w30435_ ;
	wire _w30436_ ;
	wire _w30437_ ;
	wire _w30438_ ;
	wire _w30439_ ;
	wire _w30440_ ;
	wire _w30441_ ;
	wire _w30442_ ;
	wire _w30443_ ;
	wire _w30444_ ;
	wire _w30445_ ;
	wire _w30446_ ;
	wire _w30447_ ;
	wire _w30448_ ;
	wire _w30449_ ;
	wire _w30450_ ;
	wire _w30451_ ;
	wire _w30452_ ;
	wire _w30453_ ;
	wire _w30454_ ;
	wire _w30455_ ;
	wire _w30456_ ;
	wire _w30457_ ;
	wire _w30458_ ;
	wire _w30459_ ;
	wire _w30460_ ;
	wire _w30461_ ;
	wire _w30462_ ;
	wire _w30463_ ;
	wire _w30464_ ;
	wire _w30465_ ;
	wire _w30466_ ;
	wire _w30467_ ;
	wire _w30468_ ;
	wire _w30469_ ;
	wire _w30470_ ;
	wire _w30471_ ;
	wire _w30472_ ;
	wire _w30473_ ;
	wire _w30474_ ;
	wire _w30475_ ;
	wire _w30476_ ;
	wire _w30477_ ;
	wire _w30478_ ;
	wire _w30479_ ;
	wire _w30480_ ;
	wire _w30481_ ;
	wire _w30482_ ;
	wire _w30483_ ;
	wire _w30484_ ;
	wire _w30485_ ;
	wire _w30486_ ;
	wire _w30487_ ;
	wire _w30488_ ;
	wire _w30489_ ;
	wire _w30490_ ;
	wire _w30491_ ;
	wire _w30492_ ;
	wire _w30493_ ;
	wire _w30494_ ;
	wire _w30495_ ;
	wire _w30496_ ;
	wire _w30497_ ;
	wire _w30498_ ;
	wire _w30499_ ;
	wire _w30500_ ;
	wire _w30501_ ;
	wire _w30502_ ;
	wire _w30503_ ;
	wire _w30504_ ;
	wire _w30505_ ;
	wire _w30506_ ;
	wire _w30507_ ;
	wire _w30508_ ;
	wire _w30509_ ;
	wire _w30510_ ;
	wire _w30511_ ;
	wire _w30512_ ;
	wire _w30513_ ;
	wire _w30514_ ;
	wire _w30515_ ;
	wire _w30516_ ;
	wire _w30517_ ;
	wire _w30518_ ;
	wire _w30519_ ;
	wire _w30520_ ;
	wire _w30521_ ;
	wire _w30522_ ;
	wire _w30523_ ;
	wire _w30524_ ;
	wire _w30525_ ;
	wire _w30526_ ;
	wire _w30527_ ;
	wire _w30528_ ;
	wire _w30529_ ;
	wire _w30530_ ;
	wire _w30531_ ;
	wire _w30532_ ;
	wire _w30533_ ;
	wire _w30534_ ;
	wire _w30535_ ;
	wire _w30536_ ;
	wire _w30537_ ;
	wire _w30538_ ;
	wire _w30539_ ;
	wire _w30540_ ;
	wire _w30541_ ;
	wire _w30542_ ;
	wire _w30543_ ;
	wire _w30544_ ;
	wire _w30545_ ;
	wire _w30546_ ;
	wire _w30547_ ;
	wire _w30548_ ;
	wire _w30549_ ;
	wire _w30550_ ;
	wire _w30551_ ;
	wire _w30552_ ;
	wire _w30553_ ;
	wire _w30554_ ;
	wire _w30555_ ;
	wire _w30556_ ;
	wire _w30557_ ;
	wire _w30558_ ;
	wire _w30559_ ;
	wire _w30560_ ;
	wire _w30561_ ;
	wire _w30562_ ;
	wire _w30563_ ;
	wire _w30564_ ;
	wire _w30565_ ;
	wire _w30566_ ;
	wire _w30567_ ;
	wire _w30568_ ;
	wire _w30569_ ;
	wire _w30570_ ;
	wire _w30571_ ;
	wire _w30572_ ;
	wire _w30573_ ;
	wire _w30574_ ;
	wire _w30575_ ;
	wire _w30576_ ;
	wire _w30577_ ;
	wire _w30578_ ;
	wire _w30579_ ;
	wire _w30580_ ;
	wire _w30581_ ;
	wire _w30582_ ;
	wire _w30583_ ;
	wire _w30584_ ;
	wire _w30585_ ;
	wire _w30586_ ;
	wire _w30587_ ;
	wire _w30588_ ;
	wire _w30589_ ;
	wire _w30590_ ;
	wire _w30591_ ;
	wire _w30592_ ;
	wire _w30593_ ;
	wire _w30594_ ;
	wire _w30595_ ;
	wire _w30596_ ;
	wire _w30597_ ;
	wire _w30598_ ;
	wire _w30599_ ;
	wire _w30600_ ;
	wire _w30601_ ;
	wire _w30602_ ;
	wire _w30603_ ;
	wire _w30604_ ;
	wire _w30605_ ;
	wire _w30606_ ;
	wire _w30607_ ;
	wire _w30608_ ;
	wire _w30609_ ;
	wire _w30610_ ;
	wire _w30611_ ;
	wire _w30612_ ;
	wire _w30613_ ;
	wire _w30614_ ;
	wire _w30615_ ;
	wire _w30616_ ;
	wire _w30617_ ;
	wire _w30618_ ;
	wire _w30619_ ;
	wire _w30620_ ;
	wire _w30621_ ;
	wire _w30622_ ;
	wire _w30623_ ;
	wire _w30624_ ;
	wire _w30625_ ;
	wire _w30626_ ;
	wire _w30627_ ;
	wire _w30628_ ;
	wire _w30629_ ;
	wire _w30630_ ;
	wire _w30631_ ;
	wire _w30632_ ;
	wire _w30633_ ;
	wire _w30634_ ;
	wire _w30635_ ;
	wire _w30636_ ;
	wire _w30637_ ;
	wire _w30638_ ;
	wire _w30639_ ;
	wire _w30640_ ;
	wire _w30641_ ;
	wire _w30642_ ;
	wire _w30643_ ;
	wire _w30644_ ;
	wire _w30645_ ;
	wire _w30646_ ;
	wire _w30647_ ;
	wire _w30648_ ;
	wire _w30649_ ;
	wire _w30650_ ;
	wire _w30651_ ;
	wire _w30652_ ;
	wire _w30653_ ;
	wire _w30654_ ;
	wire _w30655_ ;
	wire _w30656_ ;
	wire _w30657_ ;
	wire _w30658_ ;
	wire _w30659_ ;
	wire _w30660_ ;
	wire _w30661_ ;
	wire _w30662_ ;
	wire _w30663_ ;
	wire _w30664_ ;
	wire _w30665_ ;
	wire _w30666_ ;
	wire _w30667_ ;
	wire _w30668_ ;
	wire _w30669_ ;
	wire _w30670_ ;
	wire _w30671_ ;
	wire _w30672_ ;
	wire _w30673_ ;
	wire _w30674_ ;
	wire _w30675_ ;
	wire _w30676_ ;
	wire _w30677_ ;
	wire _w30678_ ;
	wire _w30679_ ;
	wire _w30680_ ;
	wire _w30681_ ;
	wire _w30682_ ;
	wire _w30683_ ;
	wire _w30684_ ;
	wire _w30685_ ;
	wire _w30686_ ;
	wire _w30687_ ;
	wire _w30688_ ;
	wire _w30689_ ;
	wire _w30690_ ;
	wire _w30691_ ;
	wire _w30692_ ;
	wire _w30693_ ;
	wire _w30694_ ;
	wire _w30695_ ;
	wire _w30696_ ;
	wire _w30697_ ;
	wire _w30698_ ;
	wire _w30699_ ;
	wire _w30700_ ;
	wire _w30701_ ;
	wire _w30702_ ;
	wire _w30703_ ;
	wire _w30704_ ;
	wire _w30705_ ;
	wire _w30706_ ;
	wire _w30707_ ;
	wire _w30708_ ;
	wire _w30709_ ;
	wire _w30710_ ;
	wire _w30711_ ;
	wire _w30712_ ;
	wire _w30713_ ;
	wire _w30714_ ;
	wire _w30715_ ;
	wire _w30716_ ;
	wire _w30717_ ;
	wire _w30718_ ;
	wire _w30719_ ;
	wire _w30720_ ;
	wire _w30721_ ;
	wire _w30722_ ;
	wire _w30723_ ;
	wire _w30724_ ;
	wire _w30725_ ;
	wire _w30726_ ;
	wire _w30727_ ;
	wire _w30728_ ;
	wire _w30729_ ;
	wire _w30730_ ;
	wire _w30731_ ;
	wire _w30732_ ;
	wire _w30733_ ;
	wire _w30734_ ;
	wire _w30735_ ;
	wire _w30736_ ;
	wire _w30737_ ;
	wire _w30738_ ;
	wire _w30739_ ;
	wire _w30740_ ;
	wire _w30741_ ;
	wire _w30742_ ;
	wire _w30743_ ;
	wire _w30744_ ;
	wire _w30745_ ;
	wire _w30746_ ;
	wire _w30747_ ;
	wire _w30748_ ;
	wire _w30749_ ;
	wire _w30750_ ;
	wire _w30751_ ;
	wire _w30752_ ;
	wire _w30753_ ;
	wire _w30754_ ;
	wire _w30755_ ;
	wire _w30756_ ;
	wire _w30757_ ;
	wire _w30758_ ;
	wire _w30759_ ;
	wire _w30760_ ;
	wire _w30761_ ;
	wire _w30762_ ;
	wire _w30763_ ;
	wire _w30764_ ;
	wire _w30765_ ;
	wire _w30766_ ;
	wire _w30767_ ;
	wire _w30768_ ;
	wire _w30769_ ;
	wire _w30770_ ;
	wire _w30771_ ;
	wire _w30772_ ;
	wire _w30773_ ;
	wire _w30774_ ;
	wire _w30775_ ;
	wire _w30776_ ;
	wire _w30777_ ;
	wire _w30778_ ;
	wire _w30779_ ;
	wire _w30780_ ;
	wire _w30781_ ;
	wire _w30782_ ;
	wire _w30783_ ;
	wire _w30784_ ;
	wire _w30785_ ;
	wire _w30786_ ;
	wire _w30787_ ;
	wire _w30788_ ;
	wire _w30789_ ;
	wire _w30790_ ;
	wire _w30791_ ;
	wire _w30792_ ;
	wire _w30793_ ;
	wire _w30794_ ;
	wire _w30795_ ;
	wire _w30796_ ;
	wire _w30797_ ;
	wire _w30798_ ;
	wire _w30799_ ;
	wire _w30800_ ;
	wire _w30801_ ;
	wire _w30802_ ;
	wire _w30803_ ;
	wire _w30804_ ;
	wire _w30805_ ;
	wire _w30806_ ;
	wire _w30807_ ;
	wire _w30808_ ;
	wire _w30809_ ;
	wire _w30810_ ;
	wire _w30811_ ;
	wire _w30812_ ;
	wire _w30813_ ;
	wire _w30814_ ;
	wire _w30815_ ;
	wire _w30816_ ;
	wire _w30817_ ;
	wire _w30818_ ;
	wire _w30819_ ;
	wire _w30820_ ;
	wire _w30821_ ;
	wire _w30822_ ;
	wire _w30823_ ;
	wire _w30824_ ;
	wire _w30825_ ;
	wire _w30826_ ;
	wire _w30827_ ;
	wire _w30828_ ;
	wire _w30829_ ;
	wire _w30830_ ;
	wire _w30831_ ;
	wire _w30832_ ;
	wire _w30833_ ;
	wire _w30834_ ;
	wire _w30835_ ;
	wire _w30836_ ;
	wire _w30837_ ;
	wire _w30838_ ;
	wire _w30839_ ;
	wire _w30840_ ;
	wire _w30841_ ;
	wire _w30842_ ;
	wire _w30843_ ;
	wire _w30844_ ;
	wire _w30845_ ;
	wire _w30846_ ;
	wire _w30847_ ;
	wire _w30848_ ;
	wire _w30849_ ;
	wire _w30850_ ;
	wire _w30851_ ;
	wire _w30852_ ;
	wire _w30853_ ;
	wire _w30854_ ;
	wire _w30855_ ;
	wire _w30856_ ;
	wire _w30857_ ;
	wire _w30858_ ;
	wire _w30859_ ;
	wire _w30860_ ;
	wire _w30861_ ;
	wire _w30862_ ;
	wire _w30863_ ;
	wire _w30864_ ;
	wire _w30865_ ;
	wire _w30866_ ;
	wire _w30867_ ;
	wire _w30868_ ;
	wire _w30869_ ;
	wire _w30870_ ;
	wire _w30871_ ;
	wire _w30872_ ;
	wire _w30873_ ;
	wire _w30874_ ;
	wire _w30875_ ;
	wire _w30876_ ;
	wire _w30877_ ;
	wire _w30878_ ;
	wire _w30879_ ;
	wire _w30880_ ;
	wire _w30881_ ;
	wire _w30882_ ;
	wire _w30883_ ;
	wire _w30884_ ;
	wire _w30885_ ;
	wire _w30886_ ;
	wire _w30887_ ;
	wire _w30888_ ;
	wire _w30889_ ;
	wire _w30890_ ;
	wire _w30891_ ;
	wire _w30892_ ;
	wire _w30893_ ;
	wire _w30894_ ;
	wire _w30895_ ;
	wire _w30896_ ;
	wire _w30897_ ;
	wire _w30898_ ;
	wire _w30899_ ;
	wire _w30900_ ;
	wire _w30901_ ;
	wire _w30902_ ;
	wire _w30903_ ;
	wire _w30904_ ;
	wire _w30905_ ;
	wire _w30906_ ;
	wire _w30907_ ;
	wire _w30908_ ;
	wire _w30909_ ;
	wire _w30910_ ;
	wire _w30911_ ;
	wire _w30912_ ;
	wire _w30913_ ;
	wire _w30914_ ;
	wire _w30915_ ;
	wire _w30916_ ;
	wire _w30917_ ;
	wire _w30918_ ;
	wire _w30919_ ;
	wire _w30920_ ;
	wire _w30921_ ;
	wire _w30922_ ;
	wire _w30923_ ;
	wire _w30924_ ;
	wire _w30925_ ;
	wire _w30926_ ;
	wire _w30927_ ;
	wire _w30928_ ;
	wire _w30929_ ;
	wire _w30930_ ;
	wire _w30931_ ;
	wire _w30932_ ;
	wire _w30933_ ;
	wire _w30934_ ;
	wire _w30935_ ;
	wire _w30936_ ;
	wire _w30937_ ;
	wire _w30938_ ;
	wire _w30939_ ;
	wire _w30940_ ;
	wire _w30941_ ;
	wire _w30942_ ;
	wire _w30943_ ;
	wire _w30944_ ;
	wire _w30945_ ;
	wire _w30946_ ;
	wire _w30947_ ;
	wire _w30948_ ;
	wire _w30949_ ;
	wire _w30950_ ;
	wire _w30951_ ;
	wire _w30952_ ;
	wire _w30953_ ;
	wire _w30954_ ;
	wire _w30955_ ;
	wire _w30956_ ;
	wire _w30957_ ;
	wire _w30958_ ;
	wire _w30959_ ;
	wire _w30960_ ;
	wire _w30961_ ;
	wire _w30962_ ;
	wire _w30963_ ;
	wire _w30964_ ;
	wire _w30965_ ;
	wire _w30966_ ;
	wire _w30967_ ;
	wire _w30968_ ;
	wire _w30969_ ;
	wire _w30970_ ;
	wire _w30971_ ;
	wire _w30972_ ;
	wire _w30973_ ;
	wire _w30974_ ;
	wire _w30975_ ;
	wire _w30976_ ;
	wire _w30977_ ;
	wire _w30978_ ;
	wire _w30979_ ;
	wire _w30980_ ;
	wire _w30981_ ;
	wire _w30982_ ;
	wire _w30983_ ;
	wire _w30984_ ;
	wire _w30985_ ;
	wire _w30986_ ;
	wire _w30987_ ;
	wire _w30988_ ;
	wire _w30989_ ;
	wire _w30990_ ;
	wire _w30991_ ;
	wire _w30992_ ;
	wire _w30993_ ;
	wire _w30994_ ;
	wire _w30995_ ;
	wire _w30996_ ;
	wire _w30997_ ;
	wire _w30998_ ;
	wire _w30999_ ;
	wire _w31000_ ;
	wire _w31001_ ;
	wire _w31002_ ;
	wire _w31003_ ;
	wire _w31004_ ;
	wire _w31005_ ;
	wire _w31006_ ;
	wire _w31007_ ;
	wire _w31008_ ;
	wire _w31009_ ;
	wire _w31010_ ;
	wire _w31011_ ;
	wire _w31012_ ;
	wire _w31013_ ;
	wire _w31014_ ;
	wire _w31015_ ;
	wire _w31016_ ;
	wire _w31017_ ;
	wire _w31018_ ;
	wire _w31019_ ;
	wire _w31020_ ;
	wire _w31021_ ;
	wire _w31022_ ;
	wire _w31023_ ;
	wire _w31024_ ;
	wire _w31025_ ;
	wire _w31026_ ;
	wire _w31027_ ;
	wire _w31028_ ;
	wire _w31029_ ;
	wire _w31030_ ;
	wire _w31031_ ;
	wire _w31032_ ;
	wire _w31033_ ;
	wire _w31034_ ;
	wire _w31035_ ;
	wire _w31036_ ;
	wire _w31037_ ;
	wire _w31038_ ;
	wire _w31039_ ;
	wire _w31040_ ;
	wire _w31041_ ;
	wire _w31042_ ;
	wire _w31043_ ;
	wire _w31044_ ;
	wire _w31045_ ;
	wire _w31046_ ;
	wire _w31047_ ;
	wire _w31048_ ;
	wire _w31049_ ;
	wire _w31050_ ;
	wire _w31051_ ;
	wire _w31052_ ;
	wire _w31053_ ;
	wire _w31054_ ;
	wire _w31055_ ;
	wire _w31056_ ;
	wire _w31057_ ;
	wire _w31058_ ;
	wire _w31059_ ;
	wire _w31060_ ;
	wire _w31061_ ;
	wire _w31062_ ;
	wire _w31063_ ;
	wire _w31064_ ;
	wire _w31065_ ;
	wire _w31066_ ;
	wire _w31067_ ;
	wire _w31068_ ;
	wire _w31069_ ;
	wire _w31070_ ;
	wire _w31071_ ;
	wire _w31072_ ;
	wire _w31073_ ;
	wire _w31074_ ;
	wire _w31075_ ;
	wire _w31076_ ;
	wire _w31077_ ;
	wire _w31078_ ;
	wire _w31079_ ;
	wire _w31080_ ;
	wire _w31081_ ;
	wire _w31082_ ;
	wire _w31083_ ;
	wire _w31084_ ;
	wire _w31085_ ;
	wire _w31086_ ;
	wire _w31087_ ;
	wire _w31088_ ;
	wire _w31089_ ;
	wire _w31090_ ;
	wire _w31091_ ;
	wire _w31092_ ;
	wire _w31093_ ;
	wire _w31094_ ;
	wire _w31095_ ;
	wire _w31096_ ;
	wire _w31097_ ;
	wire _w31098_ ;
	wire _w31099_ ;
	wire _w31100_ ;
	wire _w31101_ ;
	wire _w31102_ ;
	wire _w31103_ ;
	wire _w31104_ ;
	wire _w31105_ ;
	wire _w31106_ ;
	wire _w31107_ ;
	wire _w31108_ ;
	wire _w31109_ ;
	wire _w31110_ ;
	wire _w31111_ ;
	wire _w31112_ ;
	wire _w31113_ ;
	wire _w31114_ ;
	wire _w31115_ ;
	wire _w31116_ ;
	wire _w31117_ ;
	wire _w31118_ ;
	wire _w31119_ ;
	wire _w31120_ ;
	wire _w31121_ ;
	wire _w31122_ ;
	wire _w31123_ ;
	wire _w31124_ ;
	wire _w31125_ ;
	wire _w31126_ ;
	wire _w31127_ ;
	wire _w31128_ ;
	wire _w31129_ ;
	wire _w31130_ ;
	wire _w31131_ ;
	wire _w31132_ ;
	wire _w31133_ ;
	wire _w31134_ ;
	wire _w31135_ ;
	wire _w31136_ ;
	wire _w31137_ ;
	wire _w31138_ ;
	wire _w31139_ ;
	wire _w31140_ ;
	wire _w31141_ ;
	wire _w31142_ ;
	wire _w31143_ ;
	wire _w31144_ ;
	wire _w31145_ ;
	wire _w31146_ ;
	wire _w31147_ ;
	wire _w31148_ ;
	wire _w31149_ ;
	wire _w31150_ ;
	wire _w31151_ ;
	wire _w31152_ ;
	wire _w31153_ ;
	wire _w31154_ ;
	wire _w31155_ ;
	wire _w31156_ ;
	wire _w31157_ ;
	wire _w31158_ ;
	wire _w31159_ ;
	wire _w31160_ ;
	wire _w31161_ ;
	wire _w31162_ ;
	wire _w31163_ ;
	wire _w31164_ ;
	wire _w31165_ ;
	wire _w31166_ ;
	wire _w31167_ ;
	wire _w31168_ ;
	wire _w31169_ ;
	wire _w31170_ ;
	wire _w31171_ ;
	wire _w31172_ ;
	wire _w31173_ ;
	wire _w31174_ ;
	wire _w31175_ ;
	wire _w31176_ ;
	wire _w31177_ ;
	wire _w31178_ ;
	wire _w31179_ ;
	wire _w31180_ ;
	wire _w31181_ ;
	wire _w31182_ ;
	wire _w31183_ ;
	wire _w31184_ ;
	wire _w31185_ ;
	wire _w31186_ ;
	wire _w31187_ ;
	wire _w31188_ ;
	wire _w31189_ ;
	wire _w31190_ ;
	wire _w31191_ ;
	wire _w31192_ ;
	wire _w31193_ ;
	wire _w31194_ ;
	wire _w31195_ ;
	wire _w31196_ ;
	wire _w31197_ ;
	wire _w31198_ ;
	wire _w31199_ ;
	wire _w31200_ ;
	wire _w31201_ ;
	wire _w31202_ ;
	wire _w31203_ ;
	wire _w31204_ ;
	wire _w31205_ ;
	wire _w31206_ ;
	wire _w31207_ ;
	wire _w31208_ ;
	wire _w31209_ ;
	wire _w31210_ ;
	wire _w31211_ ;
	wire _w31212_ ;
	wire _w31213_ ;
	wire _w31214_ ;
	wire _w31215_ ;
	wire _w31216_ ;
	wire _w31217_ ;
	wire _w31218_ ;
	wire _w31219_ ;
	wire _w31220_ ;
	wire _w31221_ ;
	wire _w31222_ ;
	wire _w31223_ ;
	wire _w31224_ ;
	wire _w31225_ ;
	wire _w31226_ ;
	wire _w31227_ ;
	wire _w31228_ ;
	wire _w31229_ ;
	wire _w31230_ ;
	wire _w31231_ ;
	wire _w31232_ ;
	wire _w31233_ ;
	wire _w31234_ ;
	wire _w31235_ ;
	wire _w31236_ ;
	wire _w31237_ ;
	wire _w31238_ ;
	wire _w31239_ ;
	wire _w31240_ ;
	wire _w31241_ ;
	wire _w31242_ ;
	wire _w31243_ ;
	wire _w31244_ ;
	wire _w31245_ ;
	wire _w31246_ ;
	wire _w31247_ ;
	wire _w31248_ ;
	wire _w31249_ ;
	wire _w31250_ ;
	wire _w31251_ ;
	wire _w31252_ ;
	wire _w31253_ ;
	wire _w31254_ ;
	wire _w31255_ ;
	wire _w31256_ ;
	wire _w31257_ ;
	wire _w31258_ ;
	wire _w31259_ ;
	wire _w31260_ ;
	wire _w31261_ ;
	wire _w31262_ ;
	wire _w31263_ ;
	wire _w31264_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10512_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10513_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10514_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10515_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10516_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10517_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10518_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10519_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w10518_,
		_w10519_,
		_w10520_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w10516_,
		_w10517_,
		_w10521_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w10514_,
		_w10515_,
		_w10522_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w10521_,
		_w10522_,
		_w10523_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w10520_,
		_w10523_,
		_w10524_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10524_,
		_w10525_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10525_,
		_w10526_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w10513_,
		_w10526_,
		_w10527_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w10528_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\rxethmac1_crcrx_Crc_reg[0]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		_w10529_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		_w10530_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10531_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[16]/NET0131 ,
		_w10532_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\rxethmac1_crcrx_Crc_reg[17]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w10533_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[1]/NET0131 ,
		_w10534_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w10535_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\rxethmac1_crcrx_Crc_reg[22]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		_w10536_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w10537_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		_w10538_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w10539_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[3]/NET0131 ,
		_w10540_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\rxethmac1_crcrx_Crc_reg[4]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w10541_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\rxethmac1_crcrx_Crc_reg[6]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[7]/NET0131 ,
		_w10542_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\rxethmac1_crcrx_Crc_reg[8]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[9]/NET0131 ,
		_w10543_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w10542_,
		_w10543_,
		_w10544_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w10540_,
		_w10541_,
		_w10545_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w10538_,
		_w10539_,
		_w10546_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w10536_,
		_w10537_,
		_w10547_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w10534_,
		_w10535_,
		_w10548_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w10532_,
		_w10533_,
		_w10549_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w10530_,
		_w10531_,
		_w10550_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w10528_,
		_w10529_,
		_w10551_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w10550_,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w10548_,
		_w10549_,
		_w10553_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w10546_,
		_w10547_,
		_w10554_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w10544_,
		_w10545_,
		_w10555_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w10554_,
		_w10555_,
		_w10556_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w10552_,
		_w10553_,
		_w10557_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w10556_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w10527_,
		_w10558_,
		_w10559_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10559_,
		_w10560_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10512_,
		_w10561_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w10560_,
		_w10561_,
		_w10562_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		wb_rst_i_pad,
		_w10563_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10564_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10565_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10524_,
		_w10566_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w10564_,
		_w10565_,
		_w10567_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		_w10568_,
		_w10569_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		_w10568_,
		_w10570_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w10563_,
		_w10569_,
		_w10571_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w10570_,
		_w10571_,
		_w10572_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w10573_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w10573_,
		_w10574_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w10574_,
		_w10575_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w10576_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w10573_,
		_w10576_,
		_w10577_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w10577_,
		_w10578_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w10575_,
		_w10578_,
		_w10579_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w10579_,
		_w10580_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\rxethmac1_crcrx_Crc_reg[27]/NET0131 ,
		_w10580_,
		_w10581_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10582_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mtxen_pad_o_pad,
		_w10583_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\RxEnSync_reg/NET0131 ,
		mrxdv_pad_i_pad,
		_w10584_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		_w10584_,
		_w10585_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w10583_,
		_w10585_,
		_w10586_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10587_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10588_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10589_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10590_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10591_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10592_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10593_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10594_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10595_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10596_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10597_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10598_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10599_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w10600_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10601_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10602_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10603_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w10604_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w10603_,
		_w10604_,
		_w10605_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10606_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10607_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10608_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10609_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w10610_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10611_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10612_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w10613_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w10614_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10615_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w10616_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10617_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10618_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10619_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w10587_,
		_w10620_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w10588_,
		_w10589_,
		_w10621_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w10590_,
		_w10591_,
		_w10622_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w10592_,
		_w10593_,
		_w10623_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w10594_,
		_w10595_,
		_w10624_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w10596_,
		_w10597_,
		_w10625_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w10598_,
		_w10599_,
		_w10626_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w10600_,
		_w10601_,
		_w10627_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w10602_,
		_w10606_,
		_w10628_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w10607_,
		_w10608_,
		_w10629_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w10609_,
		_w10610_,
		_w10630_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w10611_,
		_w10612_,
		_w10631_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w10613_,
		_w10614_,
		_w10632_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w10615_,
		_w10616_,
		_w10633_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w10617_,
		_w10618_,
		_w10634_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w10619_,
		_w10634_,
		_w10635_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w10632_,
		_w10633_,
		_w10636_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w10630_,
		_w10631_,
		_w10637_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w10628_,
		_w10629_,
		_w10638_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w10626_,
		_w10627_,
		_w10639_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w10624_,
		_w10625_,
		_w10640_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		_w10622_,
		_w10623_,
		_w10641_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w10620_,
		_w10621_,
		_w10642_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w10605_,
		_w10642_,
		_w10643_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w10640_,
		_w10641_,
		_w10644_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w10638_,
		_w10639_,
		_w10645_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w10636_,
		_w10637_,
		_w10646_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w10635_,
		_w10646_,
		_w10647_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w10644_,
		_w10645_,
		_w10648_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w10643_,
		_w10648_,
		_w10649_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w10647_,
		_w10649_,
		_w10650_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w10586_,
		_w10650_,
		_w10651_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w10582_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mtxd_pad_o[2]_pad ,
		_w10653_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[2]_pad ,
		_w10654_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w10653_,
		_w10654_,
		_w10655_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		_w10655_,
		_w10656_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		_w10655_,
		_w10657_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w10656_,
		_w10657_,
		_w10658_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w10652_,
		_w10658_,
		_w10659_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		_w10659_,
		_w10660_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		\rxethmac1_crcrx_Crc_reg[23]/NET0131 ,
		_w10659_,
		_w10661_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w10580_,
		_w10660_,
		_w10662_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mtxd_pad_o[1]_pad ,
		_w10664_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[1]_pad ,
		_w10665_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w10664_,
		_w10665_,
		_w10666_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		_w10666_,
		_w10667_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		_w10666_,
		_w10668_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w10667_,
		_w10668_,
		_w10669_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w10652_,
		_w10669_,
		_w10670_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		_w10670_,
		_w10671_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\rxethmac1_crcrx_Crc_reg[24]/NET0131 ,
		_w10670_,
		_w10672_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		_w10580_,
		_w10671_,
		_w10673_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		_w10672_,
		_w10673_,
		_w10674_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w10568_,
		_w10675_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		_w10568_,
		_w10676_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		_w10563_,
		_w10675_,
		_w10677_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w10676_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\ethreg1_MODER_1_DataOut_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		_w10679_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		\wishbone_TxStatus_reg[11]/NET0131 ,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w10681_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		_w10682_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w10681_,
		_w10682_,
		_w10683_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\Collision_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w10684_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w10684_,
		_w10685_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w10683_,
		_w10685_,
		_w10686_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10687_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10688_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w10687_,
		_w10688_,
		_w10689_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w10689_,
		_w10690_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w10689_,
		_w10691_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w10690_,
		_w10691_,
		_w10692_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w10693_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10694_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w10687_,
		_w10694_,
		_w10695_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w10693_,
		_w10695_,
		_w10696_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w10692_,
		_w10696_,
		_w10697_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10697_,
		_w10698_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10699_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w10689_,
		_w10699_,
		_w10700_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10700_,
		_w10701_
	);
	LUT2 #(
		.INIT('h2)
	) name190 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10700_,
		_w10702_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w10701_,
		_w10702_,
		_w10703_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10703_,
		_w10704_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w10698_,
		_w10704_,
		_w10705_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10706_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w10700_,
		_w10706_,
		_w10707_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w10707_,
		_w10708_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w10707_,
		_w10709_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w10708_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w10705_,
		_w10710_,
		_w10711_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w10705_,
		_w10710_,
		_w10712_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w10711_,
		_w10712_,
		_w10713_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10713_,
		_w10714_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w10696_,
		_w10715_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w10690_,
		_w10716_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w10700_,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w10715_,
		_w10717_,
		_w10718_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w10718_,
		_w10719_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w10701_,
		_w10720_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w10707_,
		_w10720_,
		_w10721_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w10719_,
		_w10721_,
		_w10722_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w10705_,
		_w10722_,
		_w10723_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10723_,
		_w10724_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w10714_,
		_w10724_,
		_w10725_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w10698_,
		_w10703_,
		_w10726_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w10719_,
		_w10726_,
		_w10727_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10727_,
		_w10728_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w10727_,
		_w10729_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w10715_,
		_w10717_,
		_w10730_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w10718_,
		_w10730_,
		_w10731_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w10731_,
		_w10732_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w10729_,
		_w10732_,
		_w10733_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w10728_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		_w10725_,
		_w10734_,
		_w10735_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w10713_,
		_w10736_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w10723_,
		_w10737_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w10714_,
		_w10737_,
		_w10738_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w10736_,
		_w10738_,
		_w10739_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w10735_,
		_w10739_,
		_w10740_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10741_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w10707_,
		_w10741_,
		_w10742_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10742_,
		_w10743_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10743_,
		_w10744_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w10744_,
		_w10745_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w10744_,
		_w10746_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w10745_,
		_w10746_,
		_w10747_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10710_,
		_w10748_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w10705_,
		_w10748_,
		_w10749_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10742_,
		_w10750_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w10743_,
		_w10750_,
		_w10751_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10751_,
		_w10752_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w10749_,
		_w10752_,
		_w10753_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w10747_,
		_w10753_,
		_w10754_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w10747_,
		_w10753_,
		_w10755_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w10754_,
		_w10755_,
		_w10756_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10756_,
		_w10757_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w10743_,
		_w10758_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w10744_,
		_w10758_,
		_w10759_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w10721_,
		_w10760_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w10719_,
		_w10760_,
		_w10761_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w10708_,
		_w10762_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w10742_,
		_w10762_,
		_w10763_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w10761_,
		_w10764_,
		_w10765_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w10759_,
		_w10765_,
		_w10766_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w10759_,
		_w10765_,
		_w10767_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w10766_,
		_w10767_,
		_w10768_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10768_,
		_w10769_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w10757_,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w10749_,
		_w10751_,
		_w10771_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w10749_,
		_w10751_,
		_w10772_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w10771_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w10773_,
		_w10774_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w10761_,
		_w10763_,
		_w10775_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w10761_,
		_w10763_,
		_w10776_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w10775_,
		_w10776_,
		_w10777_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w10774_,
		_w10778_,
		_w10779_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w10770_,
		_w10779_,
		_w10780_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		_w10740_,
		_w10780_,
		_w10781_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w10692_,
		_w10696_,
		_w10782_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w10697_,
		_w10782_,
		_w10783_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w10783_,
		_w10784_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w10693_,
		_w10785_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w10786_,
		_w10787_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10787_,
		_w10788_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w10787_,
		_w10789_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w10788_,
		_w10789_,
		_w10790_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10790_,
		_w10791_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w10786_,
		_w10792_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w10787_,
		_w10792_,
		_w10793_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10793_,
		_w10795_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w10785_,
		_w10796_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w10786_,
		_w10796_,
		_w10797_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10797_,
		_w10799_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w10693_,
		_w10800_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w10785_,
		_w10800_,
		_w10801_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10801_,
		_w10802_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w10803_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w10693_,
		_w10803_,
		_w10804_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10806_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10807_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		_w10807_,
		_w10808_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w10806_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w10805_,
		_w10809_,
		_w10810_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10801_,
		_w10811_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10804_,
		_w10812_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w10810_,
		_w10812_,
		_w10813_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w10811_,
		_w10813_,
		_w10814_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w10799_,
		_w10802_,
		_w10815_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w10814_,
		_w10815_,
		_w10816_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w10795_,
		_w10798_,
		_w10817_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w10816_,
		_w10817_,
		_w10818_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w10791_,
		_w10794_,
		_w10819_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w10818_,
		_w10819_,
		_w10820_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w10783_,
		_w10821_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10790_,
		_w10822_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w10821_,
		_w10822_,
		_w10823_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		_w10820_,
		_w10823_,
		_w10824_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w10784_,
		_w10824_,
		_w10825_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w10731_,
		_w10826_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w10729_,
		_w10826_,
		_w10827_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w10725_,
		_w10827_,
		_w10828_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w10825_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w10780_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w10777_,
		_w10831_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w10774_,
		_w10831_,
		_w10832_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w10770_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w10756_,
		_w10834_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w10768_,
		_w10835_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w10757_,
		_w10835_,
		_w10836_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w10773_,
		_w10837_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w10770_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w10834_,
		_w10836_,
		_w10839_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w10833_,
		_w10839_,
		_w10840_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w10838_,
		_w10840_,
		_w10841_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w10781_,
		_w10830_,
		_w10842_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w10841_,
		_w10842_,
		_w10843_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w10746_,
		_w10766_,
		_w10844_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w10745_,
		_w10844_,
		_w10845_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w10845_,
		_w10846_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w10754_,
		_w10847_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w10845_,
		_w10847_,
		_w10848_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w10846_,
		_w10848_,
		_w10849_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w10843_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		\ethreg1_MODER_1_DataOut_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		_w10851_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		\wishbone_TxStatus_reg[12]/NET0131 ,
		_w10851_,
		_w10852_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w10850_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w10680_,
		_w10686_,
		_w10854_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w10853_,
		_w10854_,
		_w10855_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10806_,
		_w10856_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w10684_,
		_w10857_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w10856_,
		_w10857_,
		_w10858_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w10855_,
		_w10858_,
		_w10859_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w10684_,
		_w10860_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10860_,
		_w10861_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w10857_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w10863_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10864_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10865_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w10866_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10867_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10868_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10869_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10870_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10871_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w10872_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w10873_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10874_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10875_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w10876_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10877_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		_w10878_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w10879_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10880_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w10881_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w10882_
	);
	LUT2 #(
		.INIT('h2)
	) name371 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10883_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w10884_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10885_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w10886_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w10887_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w10888_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w10889_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w10890_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10891_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w10892_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w10893_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w10894_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w10863_,
		_w10895_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w10864_,
		_w10865_,
		_w10896_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w10866_,
		_w10867_,
		_w10897_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w10868_,
		_w10869_,
		_w10898_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w10870_,
		_w10871_,
		_w10899_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w10872_,
		_w10873_,
		_w10900_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w10874_,
		_w10875_,
		_w10901_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w10876_,
		_w10877_,
		_w10902_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w10878_,
		_w10879_,
		_w10903_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w10880_,
		_w10881_,
		_w10904_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w10882_,
		_w10883_,
		_w10905_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w10884_,
		_w10885_,
		_w10906_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w10886_,
		_w10887_,
		_w10907_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w10888_,
		_w10889_,
		_w10908_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w10890_,
		_w10891_,
		_w10909_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w10892_,
		_w10893_,
		_w10910_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w10894_,
		_w10910_,
		_w10911_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w10908_,
		_w10909_,
		_w10912_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w10906_,
		_w10907_,
		_w10913_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		_w10904_,
		_w10905_,
		_w10914_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w10902_,
		_w10903_,
		_w10915_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w10900_,
		_w10901_,
		_w10916_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w10898_,
		_w10899_,
		_w10917_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w10896_,
		_w10897_,
		_w10918_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w10895_,
		_w10918_,
		_w10919_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w10916_,
		_w10917_,
		_w10920_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w10914_,
		_w10915_,
		_w10921_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w10912_,
		_w10913_,
		_w10922_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w10911_,
		_w10922_,
		_w10923_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w10920_,
		_w10921_,
		_w10924_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w10919_,
		_w10924_,
		_w10925_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w10923_,
		_w10925_,
		_w10926_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w10862_,
		_w10926_,
		_w10927_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		_w10859_,
		_w10927_,
		_w10928_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10929_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10930_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10931_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10932_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10933_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10934_
	);
	LUT2 #(
		.INIT('h4)
	) name423 (
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10935_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10936_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w10937_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10937_,
		_w10938_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10939_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10937_,
		_w10940_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		\ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 ,
		_w10940_,
		_w10941_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w10938_,
		_w10939_,
		_w10942_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		_w10941_,
		_w10942_,
		_w10943_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w10935_,
		_w10936_,
		_w10944_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w10943_,
		_w10944_,
		_w10945_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w10933_,
		_w10934_,
		_w10946_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w10945_,
		_w10946_,
		_w10947_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w10931_,
		_w10932_,
		_w10948_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w10947_,
		_w10948_,
		_w10949_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w10929_,
		_w10930_,
		_w10950_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w10949_,
		_w10950_,
		_w10951_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10952_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w10953_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10954_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10955_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w10954_,
		_w10955_,
		_w10956_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w10957_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10958_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w10957_,
		_w10958_,
		_w10959_
	);
	LUT2 #(
		.INIT('h2)
	) name448 (
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w10960_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10961_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w10960_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w10963_
	);
	LUT2 #(
		.INIT('h2)
	) name452 (
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10964_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10965_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w10964_,
		_w10965_,
		_w10966_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w10967_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w10968_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w10967_,
		_w10968_,
		_w10969_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w10970_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w10971_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10972_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w10963_,
		_w10970_,
		_w10973_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w10971_,
		_w10972_,
		_w10974_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w10973_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w10956_,
		_w10959_,
		_w10976_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w10962_,
		_w10966_,
		_w10977_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w10969_,
		_w10977_,
		_w10978_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w10975_,
		_w10976_,
		_w10979_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w10978_,
		_w10979_,
		_w10980_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w10981_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w10952_,
		_w10981_,
		_w10982_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w10953_,
		_w10982_,
		_w10983_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w10980_,
		_w10983_,
		_w10984_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		_w10951_,
		_w10984_,
		_w10985_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w10856_,
		_w10986_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w10987_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w10988_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w10987_,
		_w10988_,
		_w10989_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w10990_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w10991_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w10992_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w10993_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		_w10994_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		_w10995_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w10994_,
		_w10995_,
		_w10996_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w10990_,
		_w10991_,
		_w10997_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w10992_,
		_w10993_,
		_w10998_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w10997_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w10989_,
		_w10996_,
		_w11000_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		_w10999_,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w11001_,
		_w11002_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		_w11003_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		_w11004_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		_w11005_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		_w11006_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		_w11007_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		_w11006_,
		_w11007_,
		_w11008_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w11004_,
		_w11005_,
		_w11009_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w11003_,
		_w11009_,
		_w11010_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w11008_,
		_w11010_,
		_w11011_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		\ethreg1_MODER_1_DataOut_reg[0]/NET0131 ,
		_w11011_,
		_w11012_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w11002_,
		_w11012_,
		_w11013_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w10986_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w11015_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11016_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w10856_,
		_w11017_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w11018_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		_w11019_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w11018_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w11017_,
		_w11020_,
		_w11021_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11022_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\txethmac1_random1_RandomLatched_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w11023_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11024_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11025_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11026_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11027_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11028_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		\txethmac1_random1_RandomLatched_reg[7]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11029_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11030_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11031_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11032_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11033_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w11032_,
		_w11033_,
		_w11034_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11035_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11036_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11037_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11038_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11039_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11040_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w11015_,
		_w11016_,
		_w11041_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w11022_,
		_w11023_,
		_w11042_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w11024_,
		_w11025_,
		_w11043_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w11026_,
		_w11027_,
		_w11044_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w11028_,
		_w11029_,
		_w11045_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w11030_,
		_w11031_,
		_w11046_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w11035_,
		_w11036_,
		_w11047_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w11037_,
		_w11038_,
		_w11048_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w11039_,
		_w11040_,
		_w11049_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		_w11048_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w11046_,
		_w11047_,
		_w11051_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		_w11044_,
		_w11045_,
		_w11052_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		_w11042_,
		_w11043_,
		_w11053_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w11034_,
		_w11041_,
		_w11054_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		_w11053_,
		_w11054_,
		_w11055_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		_w11051_,
		_w11052_,
		_w11056_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w11050_,
		_w11056_,
		_w11057_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		_w11021_,
		_w11055_,
		_w11058_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w11057_,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w10953_,
		_w11060_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w11061_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w11060_,
		_w11061_,
		_w11062_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		_w11059_,
		_w11062_,
		_w11063_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w11014_,
		_w11063_,
		_w11064_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		_w10985_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		_w10928_,
		_w11065_,
		_w11066_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w10860_,
		_w11067_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w10684_,
		_w11067_,
		_w11068_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w11069_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w11070_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11017_,
		_w11071_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		_w11069_,
		_w11070_,
		_w11072_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w11071_,
		_w11072_,
		_w11073_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w11068_,
		_w11073_,
		_w11074_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w10680_,
		_w10686_,
		_w11075_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		_w10853_,
		_w11075_,
		_w11076_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w10684_,
		_w11077_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w10680_,
		_w11077_,
		_w11078_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w10850_,
		_w11078_,
		_w11079_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w11076_,
		_w11079_,
		_w11080_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		_w11074_,
		_w11080_,
		_w11081_
	);
	LUT2 #(
		.INIT('h4)
	) name570 (
		\ethreg1_MODER_1_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w11082_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w11083_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w11084_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w11085_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w11086_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		_w11085_,
		_w11086_,
		_w11087_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		_w11083_,
		_w11084_,
		_w11088_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w11018_,
		_w11082_,
		_w11089_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w11088_,
		_w11089_,
		_w11090_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		_w10856_,
		_w11087_,
		_w11091_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		_w11090_,
		_w11091_,
		_w11092_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w11092_,
		_w11093_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w10953_,
		_w11093_,
		_w11094_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w11092_,
		_w11095_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w11096_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11097_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w11096_,
		_w11098_,
		_w11099_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		_w11095_,
		_w11099_,
		_w11100_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w10986_,
		_w11101_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w11071_,
		_w11101_,
		_w11102_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w11094_,
		_w11102_,
		_w11103_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w11100_,
		_w11103_,
		_w11104_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w11081_,
		_w11104_,
		_w11105_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		_w11066_,
		_w11105_,
		_w11106_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		_w11093_,
		_w11099_,
		_w11107_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11070_,
		_w11108_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		_w11069_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w11109_,
		_w11110_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w11111_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		_w11110_,
		_w11111_,
		_w11112_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w11107_,
		_w11112_,
		_w11113_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w11113_,
		_w11114_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w11113_,
		_w11115_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w11114_,
		_w11115_,
		_w11116_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		_w11106_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		_w11017_,
		_w11113_,
		_w11118_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		_w11018_,
		_w11118_,
		_w11119_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w11119_,
		_w11120_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w11120_,
		_w11121_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w11121_,
		_w11122_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w11122_,
		_w11123_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w11123_,
		_w11124_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w11124_,
		_w11125_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\txethmac1_txcounters1_NibCnt_reg[11]/NET0131 ,
		_w11124_,
		_w11126_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w11125_,
		_w11126_,
		_w11127_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		_w11106_,
		_w11127_,
		_w11128_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w11126_,
		_w11129_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\txethmac1_txcounters1_NibCnt_reg[12]/NET0131 ,
		_w11126_,
		_w11130_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w11129_,
		_w11130_,
		_w11131_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w11106_,
		_w11131_,
		_w11132_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		\txethmac1_txcounters1_NibCnt_reg[10]/NET0131 ,
		_w11123_,
		_w11133_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		_w11124_,
		_w11133_,
		_w11134_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		_w11106_,
		_w11134_,
		_w11135_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w11130_,
		_w11136_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\txethmac1_txcounters1_NibCnt_reg[13]/NET0131 ,
		_w11130_,
		_w11137_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		_w11136_,
		_w11137_,
		_w11138_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		_w11106_,
		_w11138_,
		_w11139_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w11137_,
		_w11140_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\txethmac1_txcounters1_NibCnt_reg[14]/NET0131 ,
		_w11137_,
		_w11141_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w11140_,
		_w11141_,
		_w11142_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		_w11106_,
		_w11142_,
		_w11143_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w11141_,
		_w11144_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		\txethmac1_txcounters1_NibCnt_reg[15]/NET0131 ,
		_w11141_,
		_w11145_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w11144_,
		_w11145_,
		_w11146_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		_w11106_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w11114_,
		_w11148_
	);
	LUT2 #(
		.INIT('h2)
	) name637 (
		_w10806_,
		_w11113_,
		_w11149_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w11148_,
		_w11149_,
		_w11150_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		_w11106_,
		_w11150_,
		_w11151_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w11149_,
		_w11152_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w10856_,
		_w11113_,
		_w11153_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w11152_,
		_w11153_,
		_w11154_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		_w11106_,
		_w11154_,
		_w11155_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w11153_,
		_w11156_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w11118_,
		_w11156_,
		_w11157_
	);
	LUT2 #(
		.INIT('h8)
	) name646 (
		_w11106_,
		_w11157_,
		_w11158_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w11118_,
		_w11159_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w11118_,
		_w11160_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		_w11159_,
		_w11160_,
		_w11161_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w11106_,
		_w11161_,
		_w11162_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w11159_,
		_w11163_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w11119_,
		_w11163_,
		_w11164_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		_w11106_,
		_w11164_,
		_w11165_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w11119_,
		_w11166_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w11120_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w11106_,
		_w11167_,
		_w11168_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		\txethmac1_txcounters1_NibCnt_reg[7]/NET0131 ,
		_w11120_,
		_w11169_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w11121_,
		_w11169_,
		_w11170_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		_w11106_,
		_w11170_,
		_w11171_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\txethmac1_txcounters1_NibCnt_reg[8]/NET0131 ,
		_w11121_,
		_w11172_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w11122_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h8)
	) name662 (
		_w11106_,
		_w11173_,
		_w11174_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		\txethmac1_txcounters1_NibCnt_reg[9]/NET0131 ,
		_w11122_,
		_w11175_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w11123_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		_w11106_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w11178_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w11178_,
		_w11179_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11180_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w11179_,
		_w11180_,
		_w11181_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		\txethmac1_txcrc_Crc_reg[26]/NET0131 ,
		_w11181_,
		_w11182_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		\txethmac1_txcrc_Crc_reg[27]/NET0131 ,
		_w11181_,
		_w11183_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		_w10959_,
		_w10969_,
		_w11184_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		_w10966_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w10972_,
		_w11185_,
		_w11186_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w10971_,
		_w11186_,
		_w11187_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		_w10956_,
		_w11187_,
		_w11188_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		_w10962_,
		_w11188_,
		_w11189_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		_w10970_,
		_w11190_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		_w11189_,
		_w11190_,
		_w11191_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w11192_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w11193_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[5]/NET0131 ,
		_w11194_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w11195_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w11196_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[4]/NET0131 ,
		_w11197_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[3]/NET0131 ,
		_w11198_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w11199_
	);
	LUT2 #(
		.INIT('h2)
	) name688 (
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[2]/NET0131 ,
		_w11200_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w11201_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[1]/NET0131 ,
		_w11202_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		\ethreg1_IPGT_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w11203_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w11202_,
		_w11203_,
		_w11204_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w11200_,
		_w11201_,
		_w11205_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w11204_,
		_w11205_,
		_w11206_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w11198_,
		_w11199_,
		_w11207_
	);
	LUT2 #(
		.INIT('h4)
	) name696 (
		_w11206_,
		_w11207_,
		_w11208_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w11196_,
		_w11197_,
		_w11209_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		_w11208_,
		_w11209_,
		_w11210_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w11194_,
		_w11195_,
		_w11211_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w11210_,
		_w11211_,
		_w11212_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w11192_,
		_w11193_,
		_w11213_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w11212_,
		_w11213_,
		_w11214_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		\txethmac1_txcounters1_NibCnt_reg[6]/NET0131 ,
		_w11215_
	);
	LUT2 #(
		.INIT('h2)
	) name704 (
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		_w11215_,
		_w11216_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w11214_,
		_w11216_,
		_w11217_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w11217_,
		_w11218_
	);
	LUT2 #(
		.INIT('h4)
	) name707 (
		_w11191_,
		_w11218_,
		_w11219_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w11219_,
		_w11220_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w11099_,
		_w11221_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w10953_,
		_w11221_,
		_w11222_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w11220_,
		_w11222_,
		_w11223_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w11066_,
		_w11223_,
		_w11224_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		\txethmac1_txstatem1_StateDefer_reg/NET0131 ,
		_w11066_,
		_w11225_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w11094_,
		_w11225_,
		_w11226_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mtxd_pad_o[3]_pad ,
		_w11227_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[3]_pad ,
		_w11228_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w11227_,
		_w11228_,
		_w11229_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		_w11229_,
		_w11230_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		_w11229_,
		_w11231_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w11230_,
		_w11231_,
		_w11232_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w10658_,
		_w11232_,
		_w11233_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		_w10658_,
		_w11232_,
		_w11234_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w11233_,
		_w11234_,
		_w11235_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		_w10652_,
		_w11235_,
		_w11236_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		_w11236_,
		_w11237_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		\rxethmac1_crcrx_Crc_reg[19]/NET0131 ,
		_w11236_,
		_w11238_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w10580_,
		_w11237_,
		_w11239_
	);
	LUT2 #(
		.INIT('h4)
	) name728 (
		_w11238_,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		_w10658_,
		_w10669_,
		_w11241_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w10658_,
		_w10669_,
		_w11242_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w11241_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h2)
	) name732 (
		_w10652_,
		_w11243_,
		_w11244_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		_w11244_,
		_w11245_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		\rxethmac1_crcrx_Crc_reg[20]/NET0131 ,
		_w11244_,
		_w11246_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		_w10580_,
		_w11245_,
		_w11247_
	);
	LUT2 #(
		.INIT('h4)
	) name736 (
		_w11246_,
		_w11247_,
		_w11248_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		\rxethmac1_crcrx_Crc_reg[26]/NET0131 ,
		_w10580_,
		_w11249_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11080_,
		_w11250_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w11074_,
		_w11250_,
		_w11251_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		_w11066_,
		_w11251_,
		_w11252_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w11074_,
		_w11253_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w10986_,
		_w11013_,
		_w11254_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w11253_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		_w11066_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		_w10686_,
		_w10853_,
		_w11257_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		\txethmac1_txstatem1_StatePAD_reg/NET0131 ,
		_w11257_,
		_w11258_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		_w11081_,
		_w11258_,
		_w11259_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w10986_,
		_w11260_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w11012_,
		_w11260_,
		_w11261_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w11059_,
		_w11261_,
		_w11262_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		_w11262_,
		_w11263_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		_w11262_,
		_w11264_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		_w10986_,
		_w11002_,
		_w11265_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		\txethmac1_StopExcessiveDeferOccured_reg/NET0131 ,
		_w11095_,
		_w11266_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		_w11099_,
		_w11266_,
		_w11267_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w11265_,
		_w11268_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w11267_,
		_w11268_,
		_w11269_
	);
	LUT2 #(
		.INIT('h8)
	) name758 (
		_w10928_,
		_w11269_,
		_w11270_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w11263_,
		_w11264_,
		_w11271_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w11270_,
		_w11271_,
		_w11272_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w11273_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		_w11262_,
		_w11273_,
		_w11274_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w11274_,
		_w11275_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w11274_,
		_w11276_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w11275_,
		_w11276_,
		_w11277_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w11270_,
		_w11277_,
		_w11278_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w11276_,
		_w11279_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w11276_,
		_w11280_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w11279_,
		_w11280_,
		_w11281_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w11270_,
		_w11281_,
		_w11282_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w11263_,
		_w11283_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w11274_,
		_w11283_,
		_w11284_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w11270_,
		_w11284_,
		_w11285_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w11286_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[7]/NET0131 ,
		_w11287_
	);
	LUT2 #(
		.INIT('h4)
	) name776 (
		\maccontrol1_transmitcontrol1_ControlData_reg[7]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11288_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		_w11286_,
		_w11287_,
		_w11289_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w11288_,
		_w11289_,
		_w11290_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[3]/NET0131 ,
		_w11291_
	);
	LUT2 #(
		.INIT('h4)
	) name780 (
		\maccontrol1_transmitcontrol1_ControlData_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11292_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11291_,
		_w11293_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w11292_,
		_w11293_,
		_w11294_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w11290_,
		_w11294_,
		_w11295_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		_w11295_,
		_w11296_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		_w11295_,
		_w11297_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		_w11296_,
		_w11297_,
		_w11298_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[4]/NET0131 ,
		_w11299_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		\maccontrol1_transmitcontrol1_ControlData_reg[4]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11300_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		_w11286_,
		_w11299_,
		_w11301_
	);
	LUT2 #(
		.INIT('h4)
	) name790 (
		_w11300_,
		_w11301_,
		_w11302_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[0]/NET0131 ,
		_w11303_
	);
	LUT2 #(
		.INIT('h4)
	) name792 (
		\maccontrol1_transmitcontrol1_ControlData_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11304_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11303_,
		_w11305_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w11304_,
		_w11305_,
		_w11306_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w11302_,
		_w11306_,
		_w11307_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w11307_,
		_w11309_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w11308_,
		_w11309_,
		_w11310_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		_w11298_,
		_w11310_,
		_w11311_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		_w11298_,
		_w11310_,
		_w11312_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11311_,
		_w11313_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		_w11312_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\txethmac1_txcrc_Crc_reg[22]/NET0131 ,
		_w11314_,
		_w11315_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		\txethmac1_txcrc_Crc_reg[22]/NET0131 ,
		_w11314_,
		_w11316_
	);
	LUT2 #(
		.INIT('h2)
	) name805 (
		_w11181_,
		_w11315_,
		_w11317_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w11316_,
		_w11317_,
		_w11318_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[2]/NET0131 ,
		_w11319_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		\maccontrol1_transmitcontrol1_ControlData_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11320_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11319_,
		_w11321_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		_w11320_,
		_w11321_,
		_w11322_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[6]/NET0131 ,
		_w11323_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		\maccontrol1_transmitcontrol1_ControlData_reg[6]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11324_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		_w11286_,
		_w11323_,
		_w11325_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w11324_,
		_w11325_,
		_w11326_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w11322_,
		_w11326_,
		_w11327_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11327_,
		_w11328_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11327_,
		_w11329_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w11328_,
		_w11329_,
		_w11330_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11330_,
		_w11331_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		\txethmac1_txcrc_Crc_reg[23]/NET0131 ,
		_w11331_,
		_w11332_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		\txethmac1_txcrc_Crc_reg[23]/NET0131 ,
		_w11331_,
		_w11333_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		_w11181_,
		_w11332_,
		_w11334_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		_w11333_,
		_w11334_,
		_w11335_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[5]/NET0131 ,
		_w11336_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		\maccontrol1_transmitcontrol1_ControlData_reg[5]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11337_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w11336_,
		_w11338_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w11337_,
		_w11338_,
		_w11339_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11339_,
		_w11340_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\wishbone_TxData_reg[1]/NET0131 ,
		_w11341_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		\maccontrol1_transmitcontrol1_ControlData_reg[1]/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w11342_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w11341_,
		_w11343_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		_w11342_,
		_w11343_,
		_w11344_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w11340_,
		_w11344_,
		_w11345_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		_w11345_,
		_w11346_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		_w11345_,
		_w11347_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w11346_,
		_w11347_,
		_w11348_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11348_,
		_w11349_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\txethmac1_txcrc_Crc_reg[24]/NET0131 ,
		_w11349_,
		_w11350_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		\txethmac1_txcrc_Crc_reg[24]/NET0131 ,
		_w11349_,
		_w11351_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		_w11181_,
		_w11350_,
		_w11352_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		_w11351_,
		_w11352_,
		_w11353_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w11094_,
		_w11354_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w11219_,
		_w11354_,
		_w11355_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		_w11066_,
		_w11355_,
		_w11356_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		_w11254_,
		_w11357_
	);
	LUT2 #(
		.INIT('h2)
	) name846 (
		_w11066_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mtxd_pad_o[0]_pad ,
		_w11359_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		\mrxd_pad_i[0]_pad ,
		_w11360_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w11359_,
		_w11360_,
		_w11361_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w11361_,
		_w11362_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w11361_,
		_w11363_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w11362_,
		_w11363_,
		_w11364_
	);
	LUT2 #(
		.INIT('h4)
	) name853 (
		_w11232_,
		_w11364_,
		_w11365_
	);
	LUT2 #(
		.INIT('h2)
	) name854 (
		_w11232_,
		_w11364_,
		_w11366_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		_w11365_,
		_w11366_,
		_w11367_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		_w10652_,
		_w11367_,
		_w11368_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		\rxethmac1_crcrx_Crc_reg[22]/NET0131 ,
		_w11368_,
		_w11369_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		\rxethmac1_crcrx_Crc_reg[22]/NET0131 ,
		_w11368_,
		_w11370_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w11369_,
		_w11370_,
		_w11371_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		_w10580_,
		_w11371_,
		_w11372_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11310_,
		_w11373_
	);
	LUT2 #(
		.INIT('h2)
	) name862 (
		\txethmac1_txcrc_Crc_reg[25]/NET0131 ,
		_w11373_,
		_w11374_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		\txethmac1_txcrc_Crc_reg[25]/NET0131 ,
		_w11373_,
		_w11375_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		_w11181_,
		_w11374_,
		_w11376_
	);
	LUT2 #(
		.INIT('h4)
	) name865 (
		_w11375_,
		_w11376_,
		_w11377_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w11067_,
		_w11378_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		_w11074_,
		_w11378_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w10927_,
		_w11067_,
		_w11380_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		\txethmac1_ColWindow_reg/NET0131 ,
		_w11001_,
		_w11381_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		_w11074_,
		_w11381_,
		_w11382_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w11267_,
		_w11379_,
		_w11383_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w11382_,
		_w11383_,
		_w11384_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		_w11380_,
		_w11384_,
		_w11385_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		_w10859_,
		_w11385_,
		_w11386_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		\txethmac1_TxDone_reg/NET0131 ,
		_w10859_,
		_w11387_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		\txethmac1_StatusLatch_reg/NET0131 ,
		_w11099_,
		_w11388_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w11387_,
		_w11388_,
		_w11389_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		\ethreg1_ResetTxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetTxCIrq_txclk_reg/NET0131 ,
		_w11390_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		\maccontrol1_transmitcontrol1_TxCtrlEndFrm_reg/NET0131 ,
		_w11391_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w10859_,
		_w11391_,
		_w11392_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w11390_,
		_w11392_,
		_w11393_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w10652_,
		_w11364_,
		_w11394_
	);
	LUT2 #(
		.INIT('h2)
	) name883 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		_w11394_,
		_w11395_
	);
	LUT2 #(
		.INIT('h4)
	) name884 (
		\rxethmac1_crcrx_Crc_reg[15]/NET0131 ,
		_w11394_,
		_w11396_
	);
	LUT2 #(
		.INIT('h2)
	) name885 (
		_w10580_,
		_w11395_,
		_w11397_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w11396_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		\rxethmac1_crcrx_Crc_reg[16]/NET0131 ,
		_w10580_,
		_w11399_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11298_,
		_w11400_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		\txethmac1_txcrc_Crc_reg[18]/NET0131 ,
		_w11400_,
		_w11401_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		\txethmac1_txcrc_Crc_reg[18]/NET0131 ,
		_w11400_,
		_w11402_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w11181_,
		_w11401_,
		_w11403_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		_w11402_,
		_w11403_,
		_w11404_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11405_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w11406_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w11405_,
		_w11406_,
		_w11407_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w11295_,
		_w11327_,
		_w11408_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		_w11295_,
		_w11327_,
		_w11409_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w11408_,
		_w11409_,
		_w11410_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w11407_,
		_w11410_,
		_w11411_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		_w11407_,
		_w11410_,
		_w11412_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11411_,
		_w11413_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		_w11412_,
		_w11413_,
		_w11414_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		\txethmac1_txcrc_Crc_reg[19]/NET0131 ,
		_w11414_,
		_w11415_
	);
	LUT2 #(
		.INIT('h4)
	) name904 (
		\txethmac1_txcrc_Crc_reg[19]/NET0131 ,
		_w11414_,
		_w11416_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		_w11181_,
		_w11415_,
		_w11417_
	);
	LUT2 #(
		.INIT('h4)
	) name906 (
		_w11416_,
		_w11417_,
		_w11418_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		_w11330_,
		_w11348_,
		_w11419_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w11330_,
		_w11348_,
		_w11420_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		_w11419_,
		_w11420_,
		_w11421_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11421_,
		_w11422_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\txethmac1_txcrc_Crc_reg[20]/NET0131 ,
		_w11422_,
		_w11423_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		\txethmac1_txcrc_Crc_reg[20]/NET0131 ,
		_w11422_,
		_w11424_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		_w11181_,
		_w11423_,
		_w11425_
	);
	LUT2 #(
		.INIT('h4)
	) name914 (
		_w11424_,
		_w11425_,
		_w11426_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		_w10652_,
		_w11232_,
		_w11427_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		_w11427_,
		_w11428_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		\rxethmac1_crcrx_Crc_reg[12]/NET0131 ,
		_w11427_,
		_w11429_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		_w10580_,
		_w11428_,
		_w11430_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		_w11429_,
		_w11430_,
		_w11431_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w11427_,
		_w11432_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		\rxethmac1_crcrx_Crc_reg[18]/NET0131 ,
		_w11427_,
		_w11433_
	);
	LUT2 #(
		.INIT('h2)
	) name922 (
		_w10580_,
		_w11432_,
		_w11434_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w11433_,
		_w11434_,
		_w11435_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		_w11310_,
		_w11348_,
		_w11436_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w11310_,
		_w11348_,
		_w11437_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w11436_,
		_w11438_
	);
	LUT2 #(
		.INIT('h4)
	) name927 (
		_w11437_,
		_w11438_,
		_w11439_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		\txethmac1_txcrc_Crc_reg[21]/NET0131 ,
		_w11439_,
		_w11440_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		\txethmac1_txcrc_Crc_reg[21]/NET0131 ,
		_w11439_,
		_w11441_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		_w11181_,
		_w11440_,
		_w11442_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w11441_,
		_w11442_,
		_w11443_
	);
	LUT2 #(
		.INIT('h2)
	) name932 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		_w11394_,
		_w11444_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		\rxethmac1_crcrx_Crc_reg[11]/NET0131 ,
		_w11394_,
		_w11445_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		_w10580_,
		_w11444_,
		_w11446_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w11445_,
		_w11446_,
		_w11447_
	);
	LUT2 #(
		.INIT('h2)
	) name936 (
		\ethreg1_ResetRxCIrq_sync2_reg/NET0131 ,
		\ethreg1_ResetRxCIrq_sync3_reg/NET0131 ,
		_w11448_
	);
	LUT2 #(
		.INIT('h2)
	) name937 (
		\ethreg1_SetRxCIrq_rxclk_reg/NET0131 ,
		_w11448_,
		_w11449_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11450_
	);
	LUT2 #(
		.INIT('h8)
	) name939 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w11450_,
		_w11451_
	);
	LUT2 #(
		.INIT('h8)
	) name940 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11451_,
		_w11452_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11453_,
		_w11454_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11454_,
		_w11455_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11455_,
		_w11456_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11456_,
		_w11457_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11457_,
		_w11458_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11458_,
		_w11459_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11459_,
		_w11460_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11460_,
		_w11461_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11461_,
		_w11462_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11462_,
		_w11463_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w11462_,
		_w11464_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		_w11463_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		_w11465_,
		_w11466_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		_w11465_,
		_w11467_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w11461_,
		_w11468_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w11462_,
		_w11468_,
		_w11469_
	);
	LUT2 #(
		.INIT('h2)
	) name958 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		_w11469_,
		_w11470_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w11460_,
		_w11471_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w11461_,
		_w11471_,
		_w11472_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		_w11472_,
		_w11473_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		_w11469_,
		_w11474_
	);
	LUT2 #(
		.INIT('h2)
	) name963 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		_w11472_,
		_w11475_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w11459_,
		_w11476_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w11460_,
		_w11476_,
		_w11477_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		_w11477_,
		_w11479_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w11458_,
		_w11480_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w11459_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		_w11481_,
		_w11482_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w11457_,
		_w11483_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w11458_,
		_w11483_,
		_w11484_
	);
	LUT2 #(
		.INIT('h2)
	) name973 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		_w11484_,
		_w11485_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		_w11481_,
		_w11486_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11451_,
		_w11487_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w11452_,
		_w11487_,
		_w11488_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w11489_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11490_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w11490_,
		_w11491_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		_w11451_,
		_w11491_,
		_w11492_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w11493_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w11490_,
		_w11494_,
		_w11495_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w10589_,
		_w10605_,
		_w11496_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		_w11496_,
		_w11497_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w11495_,
		_w11497_,
		_w11498_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w11499_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		_w11496_,
		_w11500_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w11499_,
		_w11500_,
		_w11501_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		_w11498_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w11489_,
		_w11493_,
		_w11503_
	);
	LUT2 #(
		.INIT('h4)
	) name992 (
		_w11502_,
		_w11503_,
		_w11504_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w11452_,
		_w11505_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w11453_,
		_w11505_,
		_w11506_
	);
	LUT2 #(
		.INIT('h2)
	) name995 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w11507_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w11508_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w11507_,
		_w11508_,
		_w11509_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w11504_,
		_w11509_,
		_w11510_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w11453_,
		_w11511_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w11454_,
		_w11511_,
		_w11512_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		_w11512_,
		_w11513_
	);
	LUT2 #(
		.INIT('h4)
	) name1002 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w11514_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w11513_,
		_w11514_,
		_w11515_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w11510_,
		_w11515_,
		_w11516_
	);
	LUT2 #(
		.INIT('h1)
	) name1005 (
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w11454_,
		_w11517_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w11455_,
		_w11517_,
		_w11518_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		_w11518_,
		_w11519_
	);
	LUT2 #(
		.INIT('h2)
	) name1008 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		_w11512_,
		_w11520_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w11519_,
		_w11520_,
		_w11521_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w11516_,
		_w11521_,
		_w11522_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		_w11518_,
		_w11523_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w11455_,
		_w11524_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w11456_,
		_w11524_,
		_w11525_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		_w11525_,
		_w11526_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w11523_,
		_w11526_,
		_w11527_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w11522_,
		_w11527_,
		_w11528_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		_w11525_,
		_w11529_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w11456_,
		_w11530_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w11457_,
		_w11530_,
		_w11531_
	);
	LUT2 #(
		.INIT('h2)
	) name1020 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		_w11531_,
		_w11532_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w11529_,
		_w11532_,
		_w11533_
	);
	LUT2 #(
		.INIT('h4)
	) name1022 (
		_w11528_,
		_w11533_,
		_w11534_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		_w11484_,
		_w11535_
	);
	LUT2 #(
		.INIT('h4)
	) name1024 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		_w11531_,
		_w11536_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w11535_,
		_w11536_,
		_w11537_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w11534_,
		_w11537_,
		_w11538_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w11485_,
		_w11486_,
		_w11539_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w11538_,
		_w11539_,
		_w11540_
	);
	LUT2 #(
		.INIT('h1)
	) name1029 (
		_w11479_,
		_w11482_,
		_w11541_
	);
	LUT2 #(
		.INIT('h4)
	) name1030 (
		_w11540_,
		_w11541_,
		_w11542_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w11475_,
		_w11478_,
		_w11543_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w11542_,
		_w11543_,
		_w11544_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w11473_,
		_w11474_,
		_w11545_
	);
	LUT2 #(
		.INIT('h4)
	) name1034 (
		_w11544_,
		_w11545_,
		_w11546_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w11470_,
		_w11546_,
		_w11547_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w11467_,
		_w11547_,
		_w11548_
	);
	LUT2 #(
		.INIT('h1)
	) name1037 (
		_w11466_,
		_w11548_,
		_w11549_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w11472_,
		_w11550_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w11477_,
		_w11551_
	);
	LUT2 #(
		.INIT('h2)
	) name1040 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w11481_,
		_w11552_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w11477_,
		_w11553_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w11481_,
		_w11554_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w11484_,
		_w11555_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w11484_,
		_w11556_
	);
	LUT2 #(
		.INIT('h2)
	) name1045 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w11531_,
		_w11557_
	);
	LUT2 #(
		.INIT('h2)
	) name1046 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w11525_,
		_w11558_
	);
	LUT2 #(
		.INIT('h2)
	) name1047 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w11559_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w11495_,
		_w11560_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11561_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w11562_
	);
	LUT2 #(
		.INIT('h2)
	) name1051 (
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w11563_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w11562_,
		_w11563_,
		_w11564_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w11495_,
		_w11565_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w11561_,
		_w11564_,
		_w11566_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		_w11565_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w11559_,
		_w11560_,
		_w11568_
	);
	LUT2 #(
		.INIT('h4)
	) name1057 (
		_w11567_,
		_w11568_,
		_w11569_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w11570_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w11571_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w11570_,
		_w11571_,
		_w11572_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w11569_,
		_w11572_,
		_w11573_
	);
	LUT2 #(
		.INIT('h2)
	) name1062 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w11574_
	);
	LUT2 #(
		.INIT('h2)
	) name1063 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w11575_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w11574_,
		_w11575_,
		_w11576_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w11573_,
		_w11576_,
		_w11577_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w11512_,
		_w11579_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		_w11578_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('h4)
	) name1069 (
		_w11577_,
		_w11580_,
		_w11581_
	);
	LUT2 #(
		.INIT('h2)
	) name1070 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w11518_,
		_w11582_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w11512_,
		_w11583_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w11582_,
		_w11583_,
		_w11584_
	);
	LUT2 #(
		.INIT('h4)
	) name1073 (
		_w11581_,
		_w11584_,
		_w11585_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w11518_,
		_w11586_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w11585_,
		_w11586_,
		_w11587_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w11558_,
		_w11587_,
		_w11588_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w11525_,
		_w11589_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w11531_,
		_w11590_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w11589_,
		_w11590_,
		_w11591_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		_w11588_,
		_w11591_,
		_w11592_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w11556_,
		_w11557_,
		_w11593_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w11592_,
		_w11593_,
		_w11594_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w11554_,
		_w11555_,
		_w11595_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w11594_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w11552_,
		_w11553_,
		_w11597_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w11596_,
		_w11597_,
		_w11598_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w11550_,
		_w11551_,
		_w11599_
	);
	LUT2 #(
		.INIT('h4)
	) name1088 (
		_w11598_,
		_w11599_,
		_w11600_
	);
	LUT2 #(
		.INIT('h2)
	) name1089 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w11469_,
		_w11601_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w11465_,
		_w11602_
	);
	LUT2 #(
		.INIT('h2)
	) name1091 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w11472_,
		_w11603_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w11601_,
		_w11603_,
		_w11604_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w11602_,
		_w11604_,
		_w11605_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w11600_,
		_w11605_,
		_w11606_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w11465_,
		_w11607_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w11469_,
		_w11608_
	);
	LUT2 #(
		.INIT('h4)
	) name1097 (
		_w11602_,
		_w11608_,
		_w11609_
	);
	LUT2 #(
		.INIT('h1)
	) name1098 (
		_w11607_,
		_w11609_,
		_w11610_
	);
	LUT2 #(
		.INIT('h4)
	) name1099 (
		_w11606_,
		_w11610_,
		_w11611_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w11612_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w11613_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w11612_,
		_w11613_,
		_w11614_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w11611_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h4)
	) name1104 (
		_w11549_,
		_w11615_,
		_w11616_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w11449_,
		_w11616_,
		_w11617_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_Divider2_reg/NET0131 ,
		_w11618_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		\maccontrol1_receivecontrol1_Pause_reg/NET0131 ,
		_w11618_,
		_w11619_
	);
	LUT2 #(
		.INIT('h8)
	) name1108 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 ,
		_w11619_,
		_w11620_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		_w11620_,
		_w11621_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 ,
		_w11621_,
		_w11622_
	);
	LUT2 #(
		.INIT('h8)
	) name1111 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 ,
		_w11622_,
		_w11623_
	);
	LUT2 #(
		.INIT('h8)
	) name1112 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 ,
		_w11623_,
		_w11624_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 ,
		_w11624_,
		_w11625_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 ,
		_w11626_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		_w11627_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		_w11628_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11629_
	);
	LUT2 #(
		.INIT('h8)
	) name1118 (
		_w11628_,
		_w11629_,
		_w11630_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		_w11627_,
		_w11630_,
		_w11631_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 ,
		_w11632_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		_w11633_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		_w11634_
	);
	LUT2 #(
		.INIT('h1)
	) name1123 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11635_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		_w11634_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w11632_,
		_w11633_,
		_w11637_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		_w11626_,
		_w11637_,
		_w11638_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w11636_,
		_w11638_,
		_w11639_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		_w11631_,
		_w11639_,
		_w11640_
	);
	LUT2 #(
		.INIT('h2)
	) name1129 (
		_w11625_,
		_w11640_,
		_w11641_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		_w11641_,
		_w11642_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		_w11642_,
		_w11643_
	);
	LUT2 #(
		.INIT('h4)
	) name1132 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		_w11643_,
		_w11644_
	);
	LUT2 #(
		.INIT('h2)
	) name1133 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		_w11644_,
		_w11645_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[3]/NET0131 ,
		_w11644_,
		_w11646_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w11645_,
		_w11646_,
		_w11647_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w11616_,
		_w11647_,
		_w11648_
	);
	LUT2 #(
		.INIT('h4)
	) name1137 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 ,
		_w11616_,
		_w11649_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w11648_,
		_w11649_,
		_w11650_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[0]/NET0131 ,
		_w11641_,
		_w11651_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w11642_,
		_w11651_,
		_w11652_
	);
	LUT2 #(
		.INIT('h4)
	) name1141 (
		_w11616_,
		_w11652_,
		_w11653_
	);
	LUT2 #(
		.INIT('h4)
	) name1142 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 ,
		_w11616_,
		_w11654_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w11653_,
		_w11654_,
		_w11655_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		_w11626_,
		_w11646_,
		_w11656_
	);
	LUT2 #(
		.INIT('h4)
	) name1145 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		_w11656_,
		_w11657_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		_w11657_,
		_w11658_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11658_,
		_w11659_
	);
	LUT2 #(
		.INIT('h4)
	) name1148 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11659_,
		_w11660_
	);
	LUT2 #(
		.INIT('h2)
	) name1149 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		_w11660_,
		_w11661_
	);
	LUT2 #(
		.INIT('h4)
	) name1150 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[10]/NET0131 ,
		_w11660_,
		_w11662_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w11661_,
		_w11662_,
		_w11663_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w11616_,
		_w11663_,
		_w11664_
	);
	LUT2 #(
		.INIT('h4)
	) name1153 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 ,
		_w11616_,
		_w11665_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w11664_,
		_w11665_,
		_w11666_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w11627_,
		_w11660_,
		_w11667_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		_w11667_,
		_w11668_
	);
	LUT2 #(
		.INIT('h2)
	) name1157 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		_w11668_,
		_w11669_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[13]/NET0131 ,
		_w11668_,
		_w11670_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w11616_,
		_w11669_,
		_w11671_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w11670_,
		_w11671_,
		_w11672_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 ,
		_w11616_,
		_w11673_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w11672_,
		_w11673_,
		_w11674_
	);
	LUT2 #(
		.INIT('h2)
	) name1163 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[11]/NET0131 ,
		_w11662_,
		_w11675_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		_w11667_,
		_w11675_,
		_w11676_
	);
	LUT2 #(
		.INIT('h4)
	) name1165 (
		_w11616_,
		_w11676_,
		_w11677_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 ,
		_w11616_,
		_w11678_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w11677_,
		_w11678_,
		_w11679_
	);
	LUT2 #(
		.INIT('h2)
	) name1168 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[1]/NET0131 ,
		_w11642_,
		_w11680_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w11643_,
		_w11680_,
		_w11681_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w11616_,
		_w11681_,
		_w11682_
	);
	LUT2 #(
		.INIT('h4)
	) name1171 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 ,
		_w11616_,
		_w11683_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w11682_,
		_w11683_,
		_w11684_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		_w11631_,
		_w11659_,
		_w11685_
	);
	LUT2 #(
		.INIT('h2)
	) name1174 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[15]/NET0131 ,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		_w11616_,
		_w11686_,
		_w11687_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 ,
		_w11616_,
		_w11688_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w11687_,
		_w11688_,
		_w11689_
	);
	LUT2 #(
		.INIT('h2)
	) name1178 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[2]/NET0131 ,
		_w11643_,
		_w11690_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w11644_,
		_w11690_,
		_w11691_
	);
	LUT2 #(
		.INIT('h4)
	) name1180 (
		_w11616_,
		_w11691_,
		_w11692_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 ,
		_w11616_,
		_w11693_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w11692_,
		_w11693_,
		_w11694_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[7]/NET0131 ,
		_w11657_,
		_w11695_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w11658_,
		_w11695_,
		_w11696_
	);
	LUT2 #(
		.INIT('h4)
	) name1185 (
		_w11616_,
		_w11696_,
		_w11697_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 ,
		_w11616_,
		_w11698_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w11697_,
		_w11698_,
		_w11699_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[9]/NET0131 ,
		_w11659_,
		_w11700_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w11660_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w11616_,
		_w11701_,
		_w11702_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 ,
		_w11616_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		_w11646_,
		_w11705_
	);
	LUT2 #(
		.INIT('h2)
	) name1194 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[4]/NET0131 ,
		_w11646_,
		_w11706_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		_w11705_,
		_w11706_,
		_w11707_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		_w11616_,
		_w11707_,
		_w11708_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 ,
		_w11616_,
		_w11709_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w11708_,
		_w11709_,
		_w11710_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[5]/NET0131 ,
		_w11705_,
		_w11711_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w11656_,
		_w11711_,
		_w11712_
	);
	LUT2 #(
		.INIT('h4)
	) name1201 (
		_w11616_,
		_w11712_,
		_w11713_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 ,
		_w11616_,
		_w11714_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		_w11713_,
		_w11714_,
		_w11715_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 ,
		_w11670_,
		_w11716_
	);
	LUT2 #(
		.INIT('h8)
	) name1205 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[14]/NET0131 ,
		_w11670_,
		_w11717_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w11716_,
		_w11717_,
		_w11718_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w11616_,
		_w11718_,
		_w11719_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 ,
		_w11616_,
		_w11720_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w11719_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[8]/NET0131 ,
		_w11658_,
		_w11722_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w11659_,
		_w11722_,
		_w11723_
	);
	LUT2 #(
		.INIT('h4)
	) name1212 (
		_w11616_,
		_w11723_,
		_w11724_
	);
	LUT2 #(
		.INIT('h4)
	) name1213 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 ,
		_w11616_,
		_w11725_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w11724_,
		_w11725_,
		_w11726_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[12]/NET0131 ,
		_w11667_,
		_w11727_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w11668_,
		_w11727_,
		_w11728_
	);
	LUT2 #(
		.INIT('h4)
	) name1217 (
		_w11616_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 ,
		_w11616_,
		_w11730_
	);
	LUT2 #(
		.INIT('h1)
	) name1219 (
		_w11729_,
		_w11730_,
		_w11731_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		\maccontrol1_receivecontrol1_PauseTimer_reg[6]/NET0131 ,
		_w11656_,
		_w11732_
	);
	LUT2 #(
		.INIT('h1)
	) name1221 (
		_w11657_,
		_w11732_,
		_w11733_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		_w11616_,
		_w11733_,
		_w11734_
	);
	LUT2 #(
		.INIT('h4)
	) name1223 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 ,
		_w11616_,
		_w11735_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w11734_,
		_w11735_,
		_w11736_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		_w10669_,
		_w11364_,
		_w11737_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w10669_,
		_w11364_,
		_w11738_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w11737_,
		_w11738_,
		_w11739_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		_w10658_,
		_w11739_,
		_w11740_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w10658_,
		_w11739_,
		_w11741_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w11740_,
		_w11741_,
		_w11742_
	);
	LUT2 #(
		.INIT('h8)
	) name1231 (
		_w10652_,
		_w11742_,
		_w11743_
	);
	LUT2 #(
		.INIT('h2)
	) name1232 (
		\rxethmac1_crcrx_Crc_reg[9]/NET0131 ,
		_w11743_,
		_w11744_
	);
	LUT2 #(
		.INIT('h4)
	) name1233 (
		\rxethmac1_crcrx_Crc_reg[9]/NET0131 ,
		_w11743_,
		_w11745_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		_w10580_,
		_w11744_,
		_w11746_
	);
	LUT2 #(
		.INIT('h4)
	) name1235 (
		_w11745_,
		_w11746_,
		_w11747_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\txethmac1_txcrc_Crc_reg[14]/NET0131 ,
		_w11349_,
		_w11748_
	);
	LUT2 #(
		.INIT('h4)
	) name1237 (
		\txethmac1_txcrc_Crc_reg[14]/NET0131 ,
		_w11349_,
		_w11749_
	);
	LUT2 #(
		.INIT('h2)
	) name1238 (
		_w11181_,
		_w11748_,
		_w11750_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w11749_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		\txethmac1_txcrc_Crc_reg[15]/NET0131 ,
		_w11373_,
		_w11752_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\txethmac1_txcrc_Crc_reg[15]/NET0131 ,
		_w11373_,
		_w11753_
	);
	LUT2 #(
		.INIT('h2)
	) name1242 (
		_w11181_,
		_w11752_,
		_w11754_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		_w11753_,
		_w11754_,
		_w11755_
	);
	LUT2 #(
		.INIT('h4)
	) name1244 (
		\txethmac1_txcrc_Crc_reg[16]/NET0131 ,
		_w11181_,
		_w11756_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10586_,
		_w11757_
	);
	LUT2 #(
		.INIT('h2)
	) name1246 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10651_,
		_w11758_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w11757_,
		_w11758_,
		_w11759_
	);
	LUT2 #(
		.INIT('h4)
	) name1248 (
		\macstatus1_ShortFrame_reg/NET0131 ,
		_w11759_,
		_w11760_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w11611_,
		_w11759_,
		_w11761_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11760_,
		_w11762_
	);
	LUT2 #(
		.INIT('h4)
	) name1251 (
		_w11761_,
		_w11762_,
		_w11763_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w11232_,
		_w11243_,
		_w11764_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		_w11232_,
		_w11243_,
		_w11765_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w11764_,
		_w11765_,
		_w11766_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		_w10652_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		\rxethmac1_crcrx_Crc_reg[8]/NET0131 ,
		_w11767_,
		_w11768_
	);
	LUT2 #(
		.INIT('h4)
	) name1257 (
		\rxethmac1_crcrx_Crc_reg[8]/NET0131 ,
		_w11767_,
		_w11769_
	);
	LUT2 #(
		.INIT('h2)
	) name1258 (
		_w10580_,
		_w11768_,
		_w11770_
	);
	LUT2 #(
		.INIT('h4)
	) name1259 (
		_w11769_,
		_w11770_,
		_w11771_
	);
	LUT2 #(
		.INIT('h2)
	) name1260 (
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10670_,
		_w11772_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		\rxethmac1_crcrx_Crc_reg[14]/NET0131 ,
		_w10670_,
		_w11773_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		_w10580_,
		_w11772_,
		_w11774_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w11773_,
		_w11774_,
		_w11775_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		\txethmac1_txcrc_Crc_reg[17]/NET0131 ,
		_w11181_,
		_w11776_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		\macstatus1_ReceivedPacketTooBig_reg/NET0131 ,
		_w11759_,
		_w11777_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w11759_,
		_w11778_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w11549_,
		_w11778_,
		_w11779_
	);
	LUT2 #(
		.INIT('h1)
	) name1268 (
		_w11777_,
		_w11779_,
		_w11780_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11780_,
		_w11781_
	);
	LUT2 #(
		.INIT('h2)
	) name1270 (
		\txethmac1_txcrc_Crc_reg[12]/NET0131 ,
		_w11400_,
		_w11782_
	);
	LUT2 #(
		.INIT('h4)
	) name1271 (
		\txethmac1_txcrc_Crc_reg[12]/NET0131 ,
		_w11400_,
		_w11783_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		_w11181_,
		_w11782_,
		_w11784_
	);
	LUT2 #(
		.INIT('h4)
	) name1273 (
		_w11783_,
		_w11784_,
		_w11785_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w10655_,
		_w11361_,
		_w11786_
	);
	LUT2 #(
		.INIT('h2)
	) name1275 (
		_w10655_,
		_w11361_,
		_w11787_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w11786_,
		_w11787_,
		_w11788_
	);
	LUT2 #(
		.INIT('h2)
	) name1277 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w11789_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w10528_,
		_w11789_,
		_w11790_
	);
	LUT2 #(
		.INIT('h2)
	) name1279 (
		_w11232_,
		_w11790_,
		_w11791_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w11232_,
		_w11790_,
		_w11792_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w11791_,
		_w11792_,
		_w11793_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w11788_,
		_w11793_,
		_w11794_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w11788_,
		_w11793_,
		_w11795_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w11794_,
		_w11795_,
		_w11796_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w10652_,
		_w11796_,
		_w11797_
	);
	LUT2 #(
		.INIT('h2)
	) name1286 (
		\rxethmac1_crcrx_Crc_reg[7]/NET0131 ,
		_w11797_,
		_w11798_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		\rxethmac1_crcrx_Crc_reg[7]/NET0131 ,
		_w11797_,
		_w11799_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w10580_,
		_w11798_,
		_w11800_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w11799_,
		_w11800_,
		_w11801_
	);
	LUT2 #(
		.INIT('h2)
	) name1290 (
		\txethmac1_txcrc_Crc_reg[13]/NET0131 ,
		_w11331_,
		_w11802_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		\txethmac1_txcrc_Crc_reg[13]/NET0131 ,
		_w11331_,
		_w11803_
	);
	LUT2 #(
		.INIT('h2)
	) name1292 (
		_w11181_,
		_w11802_,
		_w11804_
	);
	LUT2 #(
		.INIT('h4)
	) name1293 (
		_w11803_,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h2)
	) name1294 (
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w11244_,
		_w11806_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		\rxethmac1_crcrx_Crc_reg[5]/NET0131 ,
		_w11244_,
		_w11807_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		_w10580_,
		_w11806_,
		_w11808_
	);
	LUT2 #(
		.INIT('h4)
	) name1297 (
		_w11807_,
		_w11808_,
		_w11809_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		\txethmac1_txcrc_Crc_reg[10]/NET0131 ,
		_w11439_,
		_w11810_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		\txethmac1_txcrc_Crc_reg[10]/NET0131 ,
		_w11439_,
		_w11811_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		_w11181_,
		_w11810_,
		_w11812_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		_w11811_,
		_w11812_,
		_w11813_
	);
	LUT2 #(
		.INIT('h2)
	) name1302 (
		\txethmac1_txcrc_Crc_reg[11]/NET0131 ,
		_w11373_,
		_w11814_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		\txethmac1_txcrc_Crc_reg[11]/NET0131 ,
		_w11373_,
		_w11815_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w11181_,
		_w11814_,
		_w11816_
	);
	LUT2 #(
		.INIT('h4)
	) name1305 (
		_w11815_,
		_w11816_,
		_w11817_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		_w10652_,
		_w11739_,
		_w11818_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		_w11818_,
		_w11819_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		\rxethmac1_crcrx_Crc_reg[10]/NET0131 ,
		_w11818_,
		_w11820_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		_w10580_,
		_w11819_,
		_w11821_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		_w11820_,
		_w11821_,
		_w11822_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		\rxethmac1_crcrx_Crc_reg[4]/NET0131 ,
		_w11797_,
		_w11823_
	);
	LUT2 #(
		.INIT('h4)
	) name1312 (
		\rxethmac1_crcrx_Crc_reg[4]/NET0131 ,
		_w11797_,
		_w11824_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		_w10580_,
		_w11823_,
		_w11825_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		_w11824_,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11827_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w11828_
	);
	LUT2 #(
		.INIT('h4)
	) name1317 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w11828_,
		_w11829_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w11827_,
		_w11829_,
		_w11830_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11831_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11832_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11833_
	);
	LUT2 #(
		.INIT('h4)
	) name1322 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11833_,
		_w11834_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11832_,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name1324 (
		_w11834_,
		_w11835_,
		_w11836_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11837_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		_w11836_,
		_w11837_,
		_w11838_
	);
	LUT2 #(
		.INIT('h4)
	) name1327 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11839_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11840_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11841_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w11840_,
		_w11841_,
		_w11842_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name1332 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11844_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11845_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11846_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w11845_,
		_w11846_,
		_w11847_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11848_
	);
	LUT2 #(
		.INIT('h2)
	) name1337 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11849_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11850_
	);
	LUT2 #(
		.INIT('h4)
	) name1339 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11851_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11852_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11853_
	);
	LUT2 #(
		.INIT('h2)
	) name1342 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11854_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11855_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11856_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w11839_,
		_w11843_,
		_w11857_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w11844_,
		_w11848_,
		_w11858_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w11849_,
		_w11850_,
		_w11859_
	);
	LUT2 #(
		.INIT('h1)
	) name1348 (
		_w11851_,
		_w11852_,
		_w11860_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w11853_,
		_w11854_,
		_w11861_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w11855_,
		_w11856_,
		_w11862_
	);
	LUT2 #(
		.INIT('h8)
	) name1351 (
		_w11861_,
		_w11862_,
		_w11863_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		_w11859_,
		_w11860_,
		_w11864_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		_w11857_,
		_w11858_,
		_w11865_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w11842_,
		_w11847_,
		_w11866_
	);
	LUT2 #(
		.INIT('h8)
	) name1355 (
		_w11865_,
		_w11866_,
		_w11867_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w11863_,
		_w11864_,
		_w11868_
	);
	LUT2 #(
		.INIT('h8)
	) name1357 (
		_w11867_,
		_w11868_,
		_w11869_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w11838_,
		_w11869_,
		_w11870_
	);
	LUT2 #(
		.INIT('h2)
	) name1359 (
		_w11831_,
		_w11870_,
		_w11871_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11834_,
		_w11872_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11873_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w11832_,
		_w11873_,
		_w11874_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w11872_,
		_w11874_,
		_w11875_
	);
	LUT2 #(
		.INIT('h4)
	) name1364 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11876_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11877_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11878_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w11877_,
		_w11878_,
		_w11879_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11880_
	);
	LUT2 #(
		.INIT('h4)
	) name1369 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11881_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11882_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11883_
	);
	LUT2 #(
		.INIT('h1)
	) name1372 (
		_w11882_,
		_w11883_,
		_w11884_
	);
	LUT2 #(
		.INIT('h4)
	) name1373 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11885_
	);
	LUT2 #(
		.INIT('h2)
	) name1374 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11886_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11887_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11888_
	);
	LUT2 #(
		.INIT('h4)
	) name1377 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11889_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11890_
	);
	LUT2 #(
		.INIT('h2)
	) name1379 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11891_
	);
	LUT2 #(
		.INIT('h4)
	) name1380 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11892_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11893_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w11876_,
		_w11880_,
		_w11894_
	);
	LUT2 #(
		.INIT('h1)
	) name1383 (
		_w11881_,
		_w11885_,
		_w11895_
	);
	LUT2 #(
		.INIT('h1)
	) name1384 (
		_w11886_,
		_w11887_,
		_w11896_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		_w11888_,
		_w11889_,
		_w11897_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		_w11890_,
		_w11891_,
		_w11898_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w11892_,
		_w11893_,
		_w11899_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w11898_,
		_w11899_,
		_w11900_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w11896_,
		_w11897_,
		_w11901_
	);
	LUT2 #(
		.INIT('h8)
	) name1390 (
		_w11894_,
		_w11895_,
		_w11902_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w11879_,
		_w11884_,
		_w11903_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		_w11902_,
		_w11903_,
		_w11904_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		_w11900_,
		_w11901_,
		_w11905_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		_w11904_,
		_w11905_,
		_w11906_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w11875_,
		_w11906_,
		_w11907_
	);
	LUT2 #(
		.INIT('h2)
	) name1396 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11908_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w11908_,
		_w11909_
	);
	LUT2 #(
		.INIT('h4)
	) name1398 (
		_w11907_,
		_w11909_,
		_w11910_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w11871_,
		_w11910_,
		_w11911_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		_w11830_,
		_w11911_,
		_w11912_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		_w11829_,
		_w11913_
	);
	LUT2 #(
		.INIT('h4)
	) name1402 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11913_,
		_w11914_
	);
	LUT2 #(
		.INIT('h4)
	) name1403 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11914_,
		_w11915_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w11915_,
		_w11916_
	);
	LUT2 #(
		.INIT('h4)
	) name1405 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11917_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11918_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11919_
	);
	LUT2 #(
		.INIT('h1)
	) name1408 (
		_w11918_,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h2)
	) name1409 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11921_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11922_
	);
	LUT2 #(
		.INIT('h1)
	) name1411 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11923_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11924_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w11923_,
		_w11924_,
		_w11925_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11926_
	);
	LUT2 #(
		.INIT('h2)
	) name1415 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11927_
	);
	LUT2 #(
		.INIT('h2)
	) name1416 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11928_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11929_
	);
	LUT2 #(
		.INIT('h4)
	) name1418 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11930_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11931_
	);
	LUT2 #(
		.INIT('h2)
	) name1420 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11932_
	);
	LUT2 #(
		.INIT('h4)
	) name1421 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11933_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11934_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w11917_,
		_w11921_,
		_w11935_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w11922_,
		_w11926_,
		_w11936_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w11927_,
		_w11928_,
		_w11937_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w11929_,
		_w11930_,
		_w11938_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w11931_,
		_w11932_,
		_w11939_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w11933_,
		_w11934_,
		_w11940_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		_w11939_,
		_w11940_,
		_w11941_
	);
	LUT2 #(
		.INIT('h8)
	) name1430 (
		_w11937_,
		_w11938_,
		_w11942_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w11935_,
		_w11936_,
		_w11943_
	);
	LUT2 #(
		.INIT('h1)
	) name1432 (
		_w11920_,
		_w11925_,
		_w11944_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		_w11943_,
		_w11944_,
		_w11945_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		_w11941_,
		_w11942_,
		_w11946_
	);
	LUT2 #(
		.INIT('h8)
	) name1435 (
		_w11945_,
		_w11946_,
		_w11947_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w11838_,
		_w11947_,
		_w11948_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		_w11908_,
		_w11948_,
		_w11949_
	);
	LUT2 #(
		.INIT('h8)
	) name1438 (
		_w11836_,
		_w11873_,
		_w11950_
	);
	LUT2 #(
		.INIT('h4)
	) name1439 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11951_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11952_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11953_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w11952_,
		_w11953_,
		_w11954_
	);
	LUT2 #(
		.INIT('h2)
	) name1443 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11955_
	);
	LUT2 #(
		.INIT('h4)
	) name1444 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w11956_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11957_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11958_
	);
	LUT2 #(
		.INIT('h1)
	) name1447 (
		_w11957_,
		_w11958_,
		_w11959_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11960_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11961_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11962_
	);
	LUT2 #(
		.INIT('h4)
	) name1451 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11963_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11964_
	);
	LUT2 #(
		.INIT('h2)
	) name1453 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11965_
	);
	LUT2 #(
		.INIT('h2)
	) name1454 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11966_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w11967_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11968_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w11951_,
		_w11955_,
		_w11969_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		_w11956_,
		_w11960_,
		_w11970_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w11961_,
		_w11962_,
		_w11971_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w11963_,
		_w11964_,
		_w11972_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w11965_,
		_w11966_,
		_w11973_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w11967_,
		_w11968_,
		_w11974_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		_w11973_,
		_w11974_,
		_w11975_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		_w11971_,
		_w11972_,
		_w11976_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		_w11969_,
		_w11970_,
		_w11977_
	);
	LUT2 #(
		.INIT('h1)
	) name1466 (
		_w11954_,
		_w11959_,
		_w11978_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		_w11977_,
		_w11978_,
		_w11979_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w11975_,
		_w11976_,
		_w11980_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		_w11979_,
		_w11980_,
		_w11981_
	);
	LUT2 #(
		.INIT('h1)
	) name1470 (
		_w11950_,
		_w11981_,
		_w11982_
	);
	LUT2 #(
		.INIT('h2)
	) name1471 (
		_w11831_,
		_w11982_,
		_w11983_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w11949_,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		_w11914_,
		_w11984_,
		_w11985_
	);
	LUT2 #(
		.INIT('h1)
	) name1474 (
		_w11916_,
		_w11985_,
		_w11986_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w11830_,
		_w11986_,
		_w11987_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w11988_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11989_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w11990_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w11989_,
		_w11990_,
		_w11991_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11992_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w11993_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11994_
	);
	LUT2 #(
		.INIT('h8)
	) name1483 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w11995_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w11994_,
		_w11995_,
		_w11996_
	);
	LUT2 #(
		.INIT('h4)
	) name1485 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11997_
	);
	LUT2 #(
		.INIT('h2)
	) name1486 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w11998_
	);
	LUT2 #(
		.INIT('h2)
	) name1487 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w11999_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w12000_
	);
	LUT2 #(
		.INIT('h4)
	) name1489 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w12001_
	);
	LUT2 #(
		.INIT('h2)
	) name1490 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w12002_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w12003_
	);
	LUT2 #(
		.INIT('h4)
	) name1492 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w12004_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w12005_
	);
	LUT2 #(
		.INIT('h1)
	) name1494 (
		_w11988_,
		_w11992_,
		_w12006_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		_w11993_,
		_w11997_,
		_w12007_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w11998_,
		_w11999_,
		_w12008_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		_w12000_,
		_w12001_,
		_w12009_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w12002_,
		_w12003_,
		_w12010_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		_w12004_,
		_w12005_,
		_w12011_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		_w12008_,
		_w12009_,
		_w12013_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		_w12006_,
		_w12007_,
		_w12014_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w11991_,
		_w11996_,
		_w12015_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		_w12014_,
		_w12015_,
		_w12016_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w12012_,
		_w12013_,
		_w12017_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w12016_,
		_w12017_,
		_w12018_
	);
	LUT2 #(
		.INIT('h2)
	) name1507 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w11950_,
		_w12019_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		_w12018_,
		_w12019_,
		_w12020_
	);
	LUT2 #(
		.INIT('h4)
	) name1509 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w12021_
	);
	LUT2 #(
		.INIT('h1)
	) name1510 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w12022_
	);
	LUT2 #(
		.INIT('h8)
	) name1511 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w12023_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		_w12022_,
		_w12023_,
		_w12024_
	);
	LUT2 #(
		.INIT('h2)
	) name1513 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w12025_
	);
	LUT2 #(
		.INIT('h4)
	) name1514 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w12026_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w12027_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w12028_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w12027_,
		_w12028_,
		_w12029_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w12030_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w12031_
	);
	LUT2 #(
		.INIT('h2)
	) name1520 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w12032_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w12033_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w12034_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w12035_
	);
	LUT2 #(
		.INIT('h2)
	) name1524 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w12036_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w12037_
	);
	LUT2 #(
		.INIT('h2)
	) name1526 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w12038_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		_w12021_,
		_w12025_,
		_w12039_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w12026_,
		_w12030_,
		_w12040_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w12031_,
		_w12032_,
		_w12041_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w12033_,
		_w12034_,
		_w12042_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		_w12035_,
		_w12036_,
		_w12043_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w12037_,
		_w12038_,
		_w12044_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		_w12043_,
		_w12044_,
		_w12045_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		_w12041_,
		_w12042_,
		_w12046_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		_w12039_,
		_w12040_,
		_w12047_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		_w12024_,
		_w12029_,
		_w12048_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		_w12047_,
		_w12048_,
		_w12049_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		_w12045_,
		_w12046_,
		_w12050_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		_w12049_,
		_w12050_,
		_w12051_
	);
	LUT2 #(
		.INIT('h2)
	) name1540 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w12052_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w12053_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w12052_,
		_w12053_,
		_w12054_
	);
	LUT2 #(
		.INIT('h8)
	) name1543 (
		_w11833_,
		_w11873_,
		_w12055_
	);
	LUT2 #(
		.INIT('h8)
	) name1544 (
		_w12054_,
		_w12055_,
		_w12056_
	);
	LUT2 #(
		.INIT('h1)
	) name1545 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w12056_,
		_w12057_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		_w12051_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11830_,
		_w12059_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		_w12020_,
		_w12059_,
		_w12060_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		_w12058_,
		_w12060_,
		_w12061_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w11987_,
		_w12061_,
		_w12062_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w12062_,
		_w12063_
	);
	LUT2 #(
		.INIT('h1)
	) name1552 (
		_w11912_,
		_w12063_,
		_w12064_
	);
	LUT2 #(
		.INIT('h2)
	) name1553 (
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w11394_,
		_w12065_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		\rxethmac1_crcrx_Crc_reg[25]/NET0131 ,
		_w11394_,
		_w12066_
	);
	LUT2 #(
		.INIT('h2)
	) name1555 (
		_w10580_,
		_w12065_,
		_w12067_
	);
	LUT2 #(
		.INIT('h4)
	) name1556 (
		_w12066_,
		_w12067_,
		_w12068_
	);
	LUT2 #(
		.INIT('h4)
	) name1557 (
		_w10655_,
		_w10666_,
		_w12069_
	);
	LUT2 #(
		.INIT('h4)
	) name1558 (
		_w11361_,
		_w12069_,
		_w12070_
	);
	LUT2 #(
		.INIT('h8)
	) name1559 (
		_w11229_,
		_w12070_,
		_w12071_
	);
	LUT2 #(
		.INIT('h2)
	) name1560 (
		\WillTransmit_q2_reg/P0001 ,
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w12072_
	);
	LUT2 #(
		.INIT('h2)
	) name1561 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w12072_,
		_w12073_
	);
	LUT2 #(
		.INIT('h4)
	) name1562 (
		_w10586_,
		_w12073_,
		_w12074_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		_w12071_,
		_w12074_,
		_w12075_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w11229_,
		_w12076_
	);
	LUT2 #(
		.INIT('h8)
	) name1565 (
		_w12070_,
		_w12076_,
		_w12077_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		_w12078_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		_w12079_
	);
	LUT2 #(
		.INIT('h8)
	) name1568 (
		\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 ,
		_w12079_,
		_w12080_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w12078_,
		_w12080_,
		_w12081_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w12081_,
		_w12082_
	);
	LUT2 #(
		.INIT('h2)
	) name1571 (
		_w12077_,
		_w12082_,
		_w12083_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w12083_,
		_w12084_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w10586_,
		_w12084_,
		_w12085_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		_w12086_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w12086_,
		_w12087_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		_w10582_,
		_w12087_,
		_w12088_
	);
	LUT2 #(
		.INIT('h2)
	) name1577 (
		_w10586_,
		_w12088_,
		_w12089_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10650_,
		_w12090_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w12072_,
		_w12091_
	);
	LUT2 #(
		.INIT('h8)
	) name1580 (
		_w12077_,
		_w12082_,
		_w12092_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w12091_,
		_w12092_,
		_w12093_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		_w12090_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('h1)
	) name1583 (
		_w10586_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w12089_,
		_w12095_,
		_w12096_
	);
	LUT2 #(
		.INIT('h4)
	) name1585 (
		_w12085_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		_w12073_,
		_w12098_
	);
	LUT2 #(
		.INIT('h4)
	) name1587 (
		_w10586_,
		_w12071_,
		_w12099_
	);
	LUT2 #(
		.INIT('h4)
	) name1588 (
		_w12098_,
		_w12099_,
		_w12100_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w12100_,
		_w12101_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w12075_,
		_w12101_,
		_w12102_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w12097_,
		_w12102_,
		_w12103_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		_w11298_,
		_w11421_,
		_w12104_
	);
	LUT2 #(
		.INIT('h4)
	) name1593 (
		_w11298_,
		_w11421_,
		_w12105_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w12104_,
		_w12106_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		_w12105_,
		_w12106_,
		_w12107_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		\txethmac1_txcrc_Crc_reg[8]/NET0131 ,
		_w12107_,
		_w12108_
	);
	LUT2 #(
		.INIT('h4)
	) name1597 (
		\txethmac1_txcrc_Crc_reg[8]/NET0131 ,
		_w12107_,
		_w12109_
	);
	LUT2 #(
		.INIT('h2)
	) name1598 (
		_w11181_,
		_w12108_,
		_w12110_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w12109_,
		_w12110_,
		_w12111_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		_w11232_,
		_w11739_,
		_w12112_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		_w11232_,
		_w11739_,
		_w12113_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w12112_,
		_w12113_,
		_w12114_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w10652_,
		_w12114_,
		_w12115_
	);
	LUT2 #(
		.INIT('h2)
	) name1604 (
		\rxethmac1_crcrx_Crc_reg[3]/NET0131 ,
		_w12115_,
		_w12116_
	);
	LUT2 #(
		.INIT('h4)
	) name1605 (
		\rxethmac1_crcrx_Crc_reg[3]/NET0131 ,
		_w12115_,
		_w12117_
	);
	LUT2 #(
		.INIT('h2)
	) name1606 (
		_w10580_,
		_w12116_,
		_w12118_
	);
	LUT2 #(
		.INIT('h4)
	) name1607 (
		_w12117_,
		_w12118_,
		_w12119_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w12077_,
		_w12090_,
		_w12120_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		_w10586_,
		_w12120_,
		_w12121_
	);
	LUT2 #(
		.INIT('h4)
	) name1610 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w12098_,
		_w12122_
	);
	LUT2 #(
		.INIT('h8)
	) name1611 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w11450_,
		_w12123_
	);
	LUT2 #(
		.INIT('h8)
	) name1612 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w12124_
	);
	LUT2 #(
		.INIT('h8)
	) name1613 (
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w12124_,
		_w12125_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		_w12123_,
		_w12125_,
		_w12126_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w12127_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w12127_,
		_w12128_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w12129_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w12129_,
		_w12130_
	);
	LUT2 #(
		.INIT('h8)
	) name1619 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w12128_,
		_w12131_
	);
	LUT2 #(
		.INIT('h8)
	) name1620 (
		_w12130_,
		_w12131_,
		_w12132_
	);
	LUT2 #(
		.INIT('h8)
	) name1621 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w12133_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		_w12126_,
		_w12134_,
		_w12135_
	);
	LUT2 #(
		.INIT('h8)
	) name1624 (
		_w12132_,
		_w12135_,
		_w12136_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w10578_,
		_w12137_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w12136_,
		_w12137_,
		_w12138_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		_w12122_,
		_w12138_,
		_w12139_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w10586_,
		_w12139_,
		_w12140_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		_w12120_,
		_w12140_,
		_w12141_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w12141_,
		_w12143_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w12121_,
		_w12142_,
		_w12144_
	);
	LUT2 #(
		.INIT('h4)
	) name1633 (
		_w12143_,
		_w12144_,
		_w12145_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		_w12133_,
		_w12141_,
		_w12146_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w12126_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w12147_,
		_w12148_
	);
	LUT2 #(
		.INIT('h8)
	) name1637 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		\rxethmac1_rxcounters1_ByteCnt_reg[10]/NET0131 ,
		_w12149_,
		_w12150_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		_w12128_,
		_w12147_,
		_w12151_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w12121_,
		_w12151_,
		_w12152_
	);
	LUT2 #(
		.INIT('h4)
	) name1641 (
		_w12150_,
		_w12152_,
		_w12153_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w12151_,
		_w12154_
	);
	LUT2 #(
		.INIT('h8)
	) name1643 (
		\rxethmac1_rxcounters1_ByteCnt_reg[11]/NET0131 ,
		_w12151_,
		_w12155_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w12121_,
		_w12154_,
		_w12156_
	);
	LUT2 #(
		.INIT('h4)
	) name1645 (
		_w12155_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h8)
	) name1646 (
		_w12130_,
		_w12151_,
		_w12158_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		_w12129_,
		_w12151_,
		_w12159_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		\rxethmac1_rxcounters1_ByteCnt_reg[13]/NET0131 ,
		_w12159_,
		_w12160_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w12121_,
		_w12158_,
		_w12161_
	);
	LUT2 #(
		.INIT('h4)
	) name1650 (
		_w12160_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		\rxethmac1_rxcounters1_ByteCnt_reg[12]/NET0131 ,
		_w12155_,
		_w12163_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		_w12121_,
		_w12159_,
		_w12164_
	);
	LUT2 #(
		.INIT('h4)
	) name1653 (
		_w12163_,
		_w12164_,
		_w12165_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		\rxethmac1_rxcounters1_ByteCnt_reg[14]/NET0131 ,
		_w12158_,
		_w12166_
	);
	LUT2 #(
		.INIT('h8)
	) name1655 (
		_w12132_,
		_w12147_,
		_w12167_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		_w12121_,
		_w12167_,
		_w12168_
	);
	LUT2 #(
		.INIT('h4)
	) name1657 (
		_w12166_,
		_w12168_,
		_w12169_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w12167_,
		_w12170_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		\rxethmac1_rxcounters1_ByteCnt_reg[15]/NET0131 ,
		_w12167_,
		_w12171_
	);
	LUT2 #(
		.INIT('h1)
	) name1660 (
		_w12121_,
		_w12170_,
		_w12172_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w12171_,
		_w12172_,
		_w12173_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w12143_,
		_w12174_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w12121_,
		_w12146_,
		_w12175_
	);
	LUT2 #(
		.INIT('h4)
	) name1664 (
		_w12174_,
		_w12175_,
		_w12176_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w12146_,
		_w12177_
	);
	LUT2 #(
		.INIT('h8)
	) name1666 (
		\rxethmac1_rxcounters1_ByteCnt_reg[2]/NET0131 ,
		_w12133_,
		_w12178_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w12141_,
		_w12178_,
		_w12179_
	);
	LUT2 #(
		.INIT('h1)
	) name1668 (
		_w12121_,
		_w12179_,
		_w12180_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		_w12177_,
		_w12180_,
		_w12181_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w12179_,
		_w12182_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w12179_,
		_w12183_
	);
	LUT2 #(
		.INIT('h1)
	) name1672 (
		_w12121_,
		_w12182_,
		_w12184_
	);
	LUT2 #(
		.INIT('h4)
	) name1673 (
		_w12183_,
		_w12184_,
		_w12185_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w12123_,
		_w12146_,
		_w12186_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		\rxethmac1_rxcounters1_ByteCnt_reg[4]/NET0131 ,
		_w12183_,
		_w12187_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w12121_,
		_w12186_,
		_w12188_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w12187_,
		_w12188_,
		_w12189_
	);
	LUT2 #(
		.INIT('h8)
	) name1678 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w12186_,
		_w12190_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		\rxethmac1_rxcounters1_ByteCnt_reg[5]/NET0131 ,
		_w12186_,
		_w12191_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		_w12121_,
		_w12190_,
		_w12192_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		_w12191_,
		_w12192_,
		_w12193_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w12190_,
		_w12194_
	);
	LUT2 #(
		.INIT('h8)
	) name1683 (
		\rxethmac1_rxcounters1_ByteCnt_reg[6]/NET0131 ,
		_w12190_,
		_w12195_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w12121_,
		_w12194_,
		_w12196_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		_w12195_,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h1)
	) name1686 (
		\rxethmac1_rxcounters1_ByteCnt_reg[7]/NET0131 ,
		_w12195_,
		_w12198_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		_w12121_,
		_w12147_,
		_w12199_
	);
	LUT2 #(
		.INIT('h4)
	) name1688 (
		_w12198_,
		_w12199_,
		_w12200_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		\rxethmac1_rxcounters1_ByteCnt_reg[8]/NET0131 ,
		_w12147_,
		_w12201_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		_w12121_,
		_w12148_,
		_w12202_
	);
	LUT2 #(
		.INIT('h4)
	) name1691 (
		_w12201_,
		_w12202_,
		_w12203_
	);
	LUT2 #(
		.INIT('h1)
	) name1692 (
		\rxethmac1_rxcounters1_ByteCnt_reg[9]/NET0131 ,
		_w12148_,
		_w12204_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w12121_,
		_w12149_,
		_w12205_
	);
	LUT2 #(
		.INIT('h4)
	) name1694 (
		_w12204_,
		_w12205_,
		_w12206_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w11310_,
		_w11421_,
		_w12207_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w11310_,
		_w11421_,
		_w12208_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w12207_,
		_w12209_
	);
	LUT2 #(
		.INIT('h4)
	) name1698 (
		_w12208_,
		_w12209_,
		_w12210_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		\txethmac1_txcrc_Crc_reg[9]/NET0131 ,
		_w12210_,
		_w12211_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		\txethmac1_txcrc_Crc_reg[9]/NET0131 ,
		_w12210_,
		_w12212_
	);
	LUT2 #(
		.INIT('h2)
	) name1701 (
		_w11181_,
		_w12211_,
		_w12213_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w12212_,
		_w12213_,
		_w12214_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10651_,
		_w12215_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w12097_,
		_w12216_,
		_w12217_
	);
	LUT2 #(
		.INIT('h4)
	) name1706 (
		_w10586_,
		_w12077_,
		_w12218_
	);
	LUT2 #(
		.INIT('h1)
	) name1707 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w12218_,
		_w12219_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w12087_,
		_w12220_
	);
	LUT2 #(
		.INIT('h2)
	) name1709 (
		_w12082_,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		_w12219_,
		_w12221_,
		_w12222_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		_w12222_,
		_w12223_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		_w12223_,
		_w12224_
	);
	LUT2 #(
		.INIT('h8)
	) name1713 (
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		_w12224_,
		_w12225_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 ,
		_w12226_,
		_w12227_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\rxethmac1_rxcounters1_IFGCounter_reg[4]/NET0131 ,
		_w12226_,
		_w12228_
	);
	LUT2 #(
		.INIT('h2)
	) name1717 (
		_w12219_,
		_w12227_,
		_w12229_
	);
	LUT2 #(
		.INIT('h4)
	) name1718 (
		_w12228_,
		_w12229_,
		_w12230_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		\rxethmac1_rxcounters1_IFGCounter_reg[2]/NET0131 ,
		_w12224_,
		_w12231_
	);
	LUT2 #(
		.INIT('h2)
	) name1720 (
		_w12219_,
		_w12225_,
		_w12232_
	);
	LUT2 #(
		.INIT('h4)
	) name1721 (
		_w12231_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		\rxethmac1_rxcounters1_IFGCounter_reg[3]/NET0131 ,
		_w12225_,
		_w12234_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		_w12219_,
		_w12226_,
		_w12235_
	);
	LUT2 #(
		.INIT('h4)
	) name1724 (
		_w12234_,
		_w12235_,
		_w12236_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		\rxethmac1_rxcounters1_IFGCounter_reg[0]/NET0131 ,
		_w12222_,
		_w12237_
	);
	LUT2 #(
		.INIT('h2)
	) name1726 (
		_w12219_,
		_w12223_,
		_w12238_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w12237_,
		_w12238_,
		_w12239_
	);
	LUT2 #(
		.INIT('h4)
	) name1728 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w12240_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w12241_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w12240_,
		_w12242_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		_w12241_,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		\wishbone_tx_fifo_data_out_reg[25]/P0001 ,
		_w12243_,
		_w12244_
	);
	LUT2 #(
		.INIT('h4)
	) name1733 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		\wishbone_TxStartFrm_sync2_reg/NET0131 ,
		_w12245_
	);
	LUT2 #(
		.INIT('h8)
	) name1734 (
		\wishbone_Flop_reg/NET0131 ,
		_w12240_,
		_w12246_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w12247_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		\wishbone_TxDataLatched_reg[1]/NET0131 ,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w12249_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		\wishbone_TxDataLatched_reg[17]/NET0131 ,
		_w12249_,
		_w12250_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w12251_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		\wishbone_TxDataLatched_reg[9]/NET0131 ,
		_w12251_,
		_w12252_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w12253_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		\wishbone_TxDataLatched_reg[25]/NET0131 ,
		_w12253_,
		_w12254_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w12248_,
		_w12250_,
		_w12255_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w12252_,
		_w12254_,
		_w12256_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		_w12255_,
		_w12256_,
		_w12257_
	);
	LUT2 #(
		.INIT('h2)
	) name1746 (
		_w12246_,
		_w12257_,
		_w12258_
	);
	LUT2 #(
		.INIT('h2)
	) name1747 (
		\wishbone_TxData_reg[1]/NET0131 ,
		_w12246_,
		_w12259_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w12258_,
		_w12259_,
		_w12260_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w12243_,
		_w12260_,
		_w12261_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w12244_,
		_w12245_,
		_w12262_
	);
	LUT2 #(
		.INIT('h4)
	) name1751 (
		_w12261_,
		_w12262_,
		_w12263_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w12264_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		\wishbone_tx_fifo_data_out_reg[25]/P0001 ,
		_w12264_,
		_w12265_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		\wishbone_tx_fifo_data_out_reg[1]/P0001 ,
		_w12241_,
		_w12266_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w12267_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\wishbone_tx_fifo_data_out_reg[17]/P0001 ,
		_w12267_,
		_w12268_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w12269_
	);
	LUT2 #(
		.INIT('h8)
	) name1758 (
		\wishbone_tx_fifo_data_out_reg[9]/P0001 ,
		_w12269_,
		_w12270_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		_w12245_,
		_w12265_,
		_w12271_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w12266_,
		_w12268_,
		_w12272_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		_w12270_,
		_w12272_,
		_w12273_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w12271_,
		_w12273_,
		_w12274_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w12263_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		\wishbone_tx_fifo_data_out_reg[26]/P0001 ,
		_w12243_,
		_w12276_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\wishbone_TxDataLatched_reg[10]/NET0131 ,
		_w12251_,
		_w12277_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\wishbone_TxDataLatched_reg[26]/NET0131 ,
		_w12253_,
		_w12278_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		\wishbone_TxDataLatched_reg[2]/NET0131 ,
		_w12247_,
		_w12279_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\wishbone_TxDataLatched_reg[18]/NET0131 ,
		_w12249_,
		_w12280_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w12277_,
		_w12278_,
		_w12281_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w12279_,
		_w12280_,
		_w12282_
	);
	LUT2 #(
		.INIT('h8)
	) name1771 (
		_w12281_,
		_w12282_,
		_w12283_
	);
	LUT2 #(
		.INIT('h2)
	) name1772 (
		_w12246_,
		_w12283_,
		_w12284_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		\wishbone_TxData_reg[2]/NET0131 ,
		_w12246_,
		_w12285_
	);
	LUT2 #(
		.INIT('h1)
	) name1774 (
		_w12284_,
		_w12285_,
		_w12286_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w12243_,
		_w12286_,
		_w12287_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w12245_,
		_w12276_,
		_w12288_
	);
	LUT2 #(
		.INIT('h4)
	) name1777 (
		_w12287_,
		_w12288_,
		_w12289_
	);
	LUT2 #(
		.INIT('h8)
	) name1778 (
		\wishbone_tx_fifo_data_out_reg[26]/P0001 ,
		_w12264_,
		_w12290_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		\wishbone_tx_fifo_data_out_reg[2]/P0001 ,
		_w12241_,
		_w12291_
	);
	LUT2 #(
		.INIT('h8)
	) name1780 (
		\wishbone_tx_fifo_data_out_reg[18]/P0001 ,
		_w12267_,
		_w12292_
	);
	LUT2 #(
		.INIT('h8)
	) name1781 (
		\wishbone_tx_fifo_data_out_reg[10]/P0001 ,
		_w12269_,
		_w12293_
	);
	LUT2 #(
		.INIT('h2)
	) name1782 (
		_w12245_,
		_w12290_,
		_w12294_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w12291_,
		_w12292_,
		_w12295_
	);
	LUT2 #(
		.INIT('h4)
	) name1784 (
		_w12293_,
		_w12295_,
		_w12296_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		_w12294_,
		_w12296_,
		_w12297_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w12289_,
		_w12297_,
		_w12298_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		\wishbone_tx_fifo_data_out_reg[27]/P0001 ,
		_w12243_,
		_w12299_
	);
	LUT2 #(
		.INIT('h8)
	) name1788 (
		\wishbone_TxDataLatched_reg[3]/NET0131 ,
		_w12247_,
		_w12300_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\wishbone_TxDataLatched_reg[19]/NET0131 ,
		_w12249_,
		_w12301_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		\wishbone_TxDataLatched_reg[11]/NET0131 ,
		_w12251_,
		_w12302_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		\wishbone_TxDataLatched_reg[27]/NET0131 ,
		_w12253_,
		_w12303_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w12300_,
		_w12301_,
		_w12304_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w12302_,
		_w12303_,
		_w12305_
	);
	LUT2 #(
		.INIT('h8)
	) name1794 (
		_w12304_,
		_w12305_,
		_w12306_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		_w12246_,
		_w12306_,
		_w12307_
	);
	LUT2 #(
		.INIT('h2)
	) name1796 (
		\wishbone_TxData_reg[3]/NET0131 ,
		_w12246_,
		_w12308_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w12307_,
		_w12308_,
		_w12309_
	);
	LUT2 #(
		.INIT('h1)
	) name1798 (
		_w12243_,
		_w12309_,
		_w12310_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w12245_,
		_w12299_,
		_w12311_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		_w12310_,
		_w12311_,
		_w12312_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		\wishbone_tx_fifo_data_out_reg[27]/P0001 ,
		_w12264_,
		_w12313_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		\wishbone_tx_fifo_data_out_reg[3]/P0001 ,
		_w12241_,
		_w12314_
	);
	LUT2 #(
		.INIT('h8)
	) name1803 (
		\wishbone_tx_fifo_data_out_reg[19]/P0001 ,
		_w12267_,
		_w12315_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		\wishbone_tx_fifo_data_out_reg[11]/P0001 ,
		_w12269_,
		_w12316_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		_w12245_,
		_w12313_,
		_w12317_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w12314_,
		_w12315_,
		_w12318_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		_w12316_,
		_w12318_,
		_w12319_
	);
	LUT2 #(
		.INIT('h8)
	) name1808 (
		_w12317_,
		_w12319_,
		_w12320_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w12312_,
		_w12320_,
		_w12321_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\wishbone_tx_fifo_data_out_reg[28]/P0001 ,
		_w12243_,
		_w12322_
	);
	LUT2 #(
		.INIT('h8)
	) name1811 (
		\wishbone_TxDataLatched_reg[4]/NET0131 ,
		_w12247_,
		_w12323_
	);
	LUT2 #(
		.INIT('h8)
	) name1812 (
		\wishbone_TxDataLatched_reg[20]/NET0131 ,
		_w12249_,
		_w12324_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		\wishbone_TxDataLatched_reg[12]/NET0131 ,
		_w12251_,
		_w12325_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		\wishbone_TxDataLatched_reg[28]/NET0131 ,
		_w12253_,
		_w12326_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w12323_,
		_w12324_,
		_w12327_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w12325_,
		_w12326_,
		_w12328_
	);
	LUT2 #(
		.INIT('h8)
	) name1817 (
		_w12327_,
		_w12328_,
		_w12329_
	);
	LUT2 #(
		.INIT('h2)
	) name1818 (
		_w12246_,
		_w12329_,
		_w12330_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		\wishbone_TxData_reg[4]/NET0131 ,
		_w12246_,
		_w12331_
	);
	LUT2 #(
		.INIT('h1)
	) name1820 (
		_w12330_,
		_w12331_,
		_w12332_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w12243_,
		_w12332_,
		_w12333_
	);
	LUT2 #(
		.INIT('h1)
	) name1822 (
		_w12245_,
		_w12322_,
		_w12334_
	);
	LUT2 #(
		.INIT('h4)
	) name1823 (
		_w12333_,
		_w12334_,
		_w12335_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		\wishbone_tx_fifo_data_out_reg[28]/P0001 ,
		_w12264_,
		_w12336_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		\wishbone_tx_fifo_data_out_reg[4]/P0001 ,
		_w12241_,
		_w12337_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		\wishbone_tx_fifo_data_out_reg[20]/P0001 ,
		_w12267_,
		_w12338_
	);
	LUT2 #(
		.INIT('h8)
	) name1827 (
		\wishbone_tx_fifo_data_out_reg[12]/P0001 ,
		_w12269_,
		_w12339_
	);
	LUT2 #(
		.INIT('h2)
	) name1828 (
		_w12245_,
		_w12336_,
		_w12340_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w12337_,
		_w12338_,
		_w12341_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		_w12339_,
		_w12341_,
		_w12342_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		_w12340_,
		_w12342_,
		_w12343_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w12335_,
		_w12343_,
		_w12344_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		\wishbone_tx_fifo_data_out_reg[24]/P0001 ,
		_w12243_,
		_w12345_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		\wishbone_TxDataLatched_reg[8]/NET0131 ,
		_w12251_,
		_w12346_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		\wishbone_TxDataLatched_reg[24]/NET0131 ,
		_w12253_,
		_w12347_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		\wishbone_TxDataLatched_reg[0]/NET0131 ,
		_w12247_,
		_w12348_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		\wishbone_TxDataLatched_reg[16]/NET0131 ,
		_w12249_,
		_w12349_
	);
	LUT2 #(
		.INIT('h1)
	) name1838 (
		_w12346_,
		_w12347_,
		_w12350_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w12348_,
		_w12349_,
		_w12351_
	);
	LUT2 #(
		.INIT('h8)
	) name1840 (
		_w12350_,
		_w12351_,
		_w12352_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w12246_,
		_w12352_,
		_w12353_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		\wishbone_TxData_reg[0]/NET0131 ,
		_w12246_,
		_w12354_
	);
	LUT2 #(
		.INIT('h1)
	) name1843 (
		_w12353_,
		_w12354_,
		_w12355_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w12243_,
		_w12355_,
		_w12356_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w12245_,
		_w12345_,
		_w12357_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		_w12356_,
		_w12357_,
		_w12358_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		\wishbone_tx_fifo_data_out_reg[24]/P0001 ,
		_w12264_,
		_w12359_
	);
	LUT2 #(
		.INIT('h8)
	) name1848 (
		\wishbone_tx_fifo_data_out_reg[0]/P0001 ,
		_w12241_,
		_w12360_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		\wishbone_tx_fifo_data_out_reg[16]/P0001 ,
		_w12267_,
		_w12361_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		\wishbone_tx_fifo_data_out_reg[8]/P0001 ,
		_w12269_,
		_w12362_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		_w12245_,
		_w12359_,
		_w12363_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w12360_,
		_w12361_,
		_w12364_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		_w12362_,
		_w12364_,
		_w12365_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w12363_,
		_w12365_,
		_w12366_
	);
	LUT2 #(
		.INIT('h1)
	) name1855 (
		_w12358_,
		_w12366_,
		_w12367_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		\wishbone_tx_fifo_data_out_reg[30]/P0001 ,
		_w12243_,
		_w12368_
	);
	LUT2 #(
		.INIT('h8)
	) name1857 (
		\wishbone_TxDataLatched_reg[6]/NET0131 ,
		_w12247_,
		_w12369_
	);
	LUT2 #(
		.INIT('h8)
	) name1858 (
		\wishbone_TxDataLatched_reg[22]/NET0131 ,
		_w12249_,
		_w12370_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		\wishbone_TxDataLatched_reg[14]/NET0131 ,
		_w12251_,
		_w12371_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		\wishbone_TxDataLatched_reg[30]/NET0131 ,
		_w12253_,
		_w12372_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		_w12369_,
		_w12370_,
		_w12373_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w12371_,
		_w12372_,
		_w12374_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		_w12373_,
		_w12374_,
		_w12375_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		_w12246_,
		_w12375_,
		_w12376_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		\wishbone_TxData_reg[6]/NET0131 ,
		_w12246_,
		_w12377_
	);
	LUT2 #(
		.INIT('h1)
	) name1866 (
		_w12376_,
		_w12377_,
		_w12378_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w12243_,
		_w12378_,
		_w12379_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w12245_,
		_w12368_,
		_w12380_
	);
	LUT2 #(
		.INIT('h4)
	) name1869 (
		_w12379_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		\wishbone_tx_fifo_data_out_reg[30]/P0001 ,
		_w12264_,
		_w12382_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		\wishbone_tx_fifo_data_out_reg[6]/P0001 ,
		_w12241_,
		_w12383_
	);
	LUT2 #(
		.INIT('h8)
	) name1872 (
		\wishbone_tx_fifo_data_out_reg[22]/P0001 ,
		_w12267_,
		_w12384_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		\wishbone_tx_fifo_data_out_reg[14]/P0001 ,
		_w12269_,
		_w12385_
	);
	LUT2 #(
		.INIT('h2)
	) name1874 (
		_w12245_,
		_w12382_,
		_w12386_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w12383_,
		_w12384_,
		_w12387_
	);
	LUT2 #(
		.INIT('h4)
	) name1876 (
		_w12385_,
		_w12387_,
		_w12388_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		_w12386_,
		_w12388_,
		_w12389_
	);
	LUT2 #(
		.INIT('h1)
	) name1878 (
		_w12381_,
		_w12389_,
		_w12390_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		\wishbone_tx_fifo_data_out_reg[29]/P0001 ,
		_w12243_,
		_w12391_
	);
	LUT2 #(
		.INIT('h8)
	) name1880 (
		\wishbone_TxDataLatched_reg[5]/NET0131 ,
		_w12247_,
		_w12392_
	);
	LUT2 #(
		.INIT('h8)
	) name1881 (
		\wishbone_TxDataLatched_reg[21]/NET0131 ,
		_w12249_,
		_w12393_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		\wishbone_TxDataLatched_reg[13]/NET0131 ,
		_w12251_,
		_w12394_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		\wishbone_TxDataLatched_reg[29]/NET0131 ,
		_w12253_,
		_w12395_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w12392_,
		_w12393_,
		_w12396_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w12394_,
		_w12395_,
		_w12397_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		_w12396_,
		_w12397_,
		_w12398_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		_w12246_,
		_w12398_,
		_w12399_
	);
	LUT2 #(
		.INIT('h2)
	) name1888 (
		\wishbone_TxData_reg[5]/NET0131 ,
		_w12246_,
		_w12400_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w12399_,
		_w12400_,
		_w12401_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w12243_,
		_w12401_,
		_w12402_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w12245_,
		_w12391_,
		_w12403_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		_w12402_,
		_w12403_,
		_w12404_
	);
	LUT2 #(
		.INIT('h8)
	) name1893 (
		\wishbone_tx_fifo_data_out_reg[29]/P0001 ,
		_w12264_,
		_w12405_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		\wishbone_tx_fifo_data_out_reg[5]/P0001 ,
		_w12241_,
		_w12406_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		\wishbone_tx_fifo_data_out_reg[21]/P0001 ,
		_w12267_,
		_w12407_
	);
	LUT2 #(
		.INIT('h8)
	) name1896 (
		\wishbone_tx_fifo_data_out_reg[13]/P0001 ,
		_w12269_,
		_w12408_
	);
	LUT2 #(
		.INIT('h2)
	) name1897 (
		_w12245_,
		_w12405_,
		_w12409_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w12406_,
		_w12407_,
		_w12410_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w12408_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		_w12409_,
		_w12411_,
		_w12412_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w12404_,
		_w12412_,
		_w12413_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		\wishbone_tx_fifo_data_out_reg[31]/P0001 ,
		_w12243_,
		_w12414_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		\wishbone_TxDataLatched_reg[7]/NET0131 ,
		_w12247_,
		_w12415_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		\wishbone_TxDataLatched_reg[23]/NET0131 ,
		_w12249_,
		_w12416_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		\wishbone_TxDataLatched_reg[15]/NET0131 ,
		_w12251_,
		_w12417_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		\wishbone_TxDataLatched_reg[31]/NET0131 ,
		_w12253_,
		_w12418_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w12415_,
		_w12416_,
		_w12419_
	);
	LUT2 #(
		.INIT('h1)
	) name1908 (
		_w12417_,
		_w12418_,
		_w12420_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		_w12419_,
		_w12420_,
		_w12421_
	);
	LUT2 #(
		.INIT('h2)
	) name1910 (
		_w12246_,
		_w12421_,
		_w12422_
	);
	LUT2 #(
		.INIT('h2)
	) name1911 (
		\wishbone_TxData_reg[7]/NET0131 ,
		_w12246_,
		_w12423_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		_w12422_,
		_w12423_,
		_w12424_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w12243_,
		_w12424_,
		_w12425_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		_w12245_,
		_w12414_,
		_w12426_
	);
	LUT2 #(
		.INIT('h4)
	) name1915 (
		_w12425_,
		_w12426_,
		_w12427_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		\wishbone_tx_fifo_data_out_reg[31]/P0001 ,
		_w12264_,
		_w12428_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		\wishbone_tx_fifo_data_out_reg[7]/P0001 ,
		_w12241_,
		_w12429_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		\wishbone_tx_fifo_data_out_reg[23]/P0001 ,
		_w12267_,
		_w12430_
	);
	LUT2 #(
		.INIT('h8)
	) name1919 (
		\wishbone_tx_fifo_data_out_reg[15]/P0001 ,
		_w12269_,
		_w12431_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		_w12245_,
		_w12428_,
		_w12432_
	);
	LUT2 #(
		.INIT('h1)
	) name1921 (
		_w12429_,
		_w12430_,
		_w12433_
	);
	LUT2 #(
		.INIT('h4)
	) name1922 (
		_w12431_,
		_w12433_,
		_w12434_
	);
	LUT2 #(
		.INIT('h8)
	) name1923 (
		_w12432_,
		_w12434_,
		_w12435_
	);
	LUT2 #(
		.INIT('h1)
	) name1924 (
		_w12427_,
		_w12435_,
		_w12436_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		\rxethmac1_crcrx_Crc_reg[1]/NET0131 ,
		_w11797_,
		_w12437_
	);
	LUT2 #(
		.INIT('h4)
	) name1926 (
		\rxethmac1_crcrx_Crc_reg[1]/NET0131 ,
		_w11797_,
		_w12438_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w10580_,
		_w12437_,
		_w12439_
	);
	LUT2 #(
		.INIT('h4)
	) name1928 (
		_w12438_,
		_w12439_,
		_w12440_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		\rxethmac1_rxcounters1_IFGCounter_reg[1]/NET0131 ,
		_w12223_,
		_w12441_
	);
	LUT2 #(
		.INIT('h2)
	) name1930 (
		_w12219_,
		_w12224_,
		_w12442_
	);
	LUT2 #(
		.INIT('h4)
	) name1931 (
		_w12441_,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w12088_,
		_w12444_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w10586_,
		_w12444_,
		_w12445_
	);
	LUT2 #(
		.INIT('h2)
	) name1934 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w12446_
	);
	LUT2 #(
		.INIT('h4)
	) name1935 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w12447_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w12446_,
		_w12447_,
		_w12448_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w11298_,
		_w11307_,
		_w12449_
	);
	LUT2 #(
		.INIT('h8)
	) name1938 (
		_w11298_,
		_w11307_,
		_w12450_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w12449_,
		_w12450_,
		_w12451_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w11345_,
		_w12451_,
		_w12452_
	);
	LUT2 #(
		.INIT('h8)
	) name1941 (
		_w11345_,
		_w12451_,
		_w12453_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w12452_,
		_w12453_,
		_w12454_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w12448_,
		_w12454_,
		_w12455_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		_w12448_,
		_w12454_,
		_w12456_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w12455_,
		_w12457_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		_w12456_,
		_w12457_,
		_w12458_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		\txethmac1_txcrc_Crc_reg[6]/NET0131 ,
		_w12458_,
		_w12459_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		\txethmac1_txcrc_Crc_reg[6]/NET0131 ,
		_w12458_,
		_w12460_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		_w11181_,
		_w12459_,
		_w12461_
	);
	LUT2 #(
		.INIT('h4)
	) name1950 (
		_w12460_,
		_w12461_,
		_w12462_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w12463_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w12464_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w12463_,
		_w12464_,
		_w12465_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w11327_,
		_w12451_,
		_w12466_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		_w11327_,
		_w12451_,
		_w12467_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w12466_,
		_w12467_,
		_w12468_
	);
	LUT2 #(
		.INIT('h1)
	) name1957 (
		_w12465_,
		_w12468_,
		_w12469_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		_w12465_,
		_w12468_,
		_w12470_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w12469_,
		_w12471_
	);
	LUT2 #(
		.INIT('h4)
	) name1960 (
		_w12470_,
		_w12471_,
		_w12472_
	);
	LUT2 #(
		.INIT('h2)
	) name1961 (
		\txethmac1_txcrc_Crc_reg[7]/NET0131 ,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('h4)
	) name1962 (
		\txethmac1_txcrc_Crc_reg[7]/NET0131 ,
		_w12472_,
		_w12474_
	);
	LUT2 #(
		.INIT('h2)
	) name1963 (
		_w11181_,
		_w12473_,
		_w12475_
	);
	LUT2 #(
		.INIT('h4)
	) name1964 (
		_w12474_,
		_w12475_,
		_w12476_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w12477_
	);
	LUT2 #(
		.INIT('h8)
	) name1966 (
		\rxethmac1_Broadcast_reg/NET0131 ,
		_w12477_,
		_w12478_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		\rxethmac1_LatchedByte_reg[4]/NET0131 ,
		\rxethmac1_LatchedByte_reg[5]/NET0131 ,
		_w12479_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		\rxethmac1_LatchedByte_reg[6]/NET0131 ,
		\rxethmac1_LatchedByte_reg[7]/NET0131 ,
		_w12480_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		_w12479_,
		_w12480_,
		_w12481_
	);
	LUT2 #(
		.INIT('h2)
	) name1970 (
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w12482_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		_w10564_,
		_w12482_,
		_w12483_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		_w10525_,
		_w12483_,
		_w12484_
	);
	LUT2 #(
		.INIT('h8)
	) name1973 (
		_w12481_,
		_w12484_,
		_w12485_
	);
	LUT2 #(
		.INIT('h1)
	) name1974 (
		_w12478_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h8)
	) name1975 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		\rxethmac1_LatchedByte_reg[1]/NET0131 ,
		_w12487_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		\rxethmac1_LatchedByte_reg[2]/NET0131 ,
		\rxethmac1_LatchedByte_reg[3]/NET0131 ,
		_w12488_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w12487_,
		_w12488_,
		_w12489_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		_w12481_,
		_w12489_,
		_w12490_
	);
	LUT2 #(
		.INIT('h2)
	) name1979 (
		_w10564_,
		_w12178_,
		_w12491_
	);
	LUT2 #(
		.INIT('h4)
	) name1980 (
		_w12490_,
		_w12491_,
		_w12492_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w10524_,
		_w12492_,
		_w12493_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w12486_,
		_w12493_,
		_w12494_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w12085_,
		_w12495_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		_w12215_,
		_w12495_,
		_w12496_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		_w12096_,
		_w12496_,
		_w12497_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		\rxethmac1_rxstatem1_StatePreamble_reg/NET0131 ,
		_w12075_,
		_w12498_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		_w12099_,
		_w12498_,
		_w12499_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		_w12096_,
		_w12499_,
		_w12500_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w10565_,
		_w10582_,
		_w12501_
	);
	LUT2 #(
		.INIT('h8)
	) name1990 (
		_w10526_,
		_w12501_,
		_w12502_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		_w10582_,
		_w12133_,
		_w12503_
	);
	LUT2 #(
		.INIT('h8)
	) name1992 (
		_w10526_,
		_w12503_,
		_w12504_
	);
	LUT2 #(
		.INIT('h4)
	) name1993 (
		_w11906_,
		_w12504_,
		_w12505_
	);
	LUT2 #(
		.INIT('h1)
	) name1994 (
		\rxethmac1_rxcounters1_ByteCnt_reg[3]/NET0131 ,
		_w10582_,
		_w12506_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		_w10566_,
		_w12506_,
		_w12507_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		_w10513_,
		_w12507_,
		_w12508_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		_w12051_,
		_w12508_,
		_w12509_
	);
	LUT2 #(
		.INIT('h8)
	) name1998 (
		_w12482_,
		_w12507_,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		_w10565_,
		_w12507_,
		_w12511_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w12133_,
		_w12507_,
		_w12512_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w12477_,
		_w12512_,
		_w12513_
	);
	LUT2 #(
		.INIT('h4)
	) name2002 (
		_w11947_,
		_w12512_,
		_w12514_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w12511_,
		_w12513_,
		_w12515_
	);
	LUT2 #(
		.INIT('h4)
	) name2004 (
		_w12514_,
		_w12515_,
		_w12516_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		_w11981_,
		_w12511_,
		_w12517_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		_w12516_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w12510_,
		_w12518_,
		_w12519_
	);
	LUT2 #(
		.INIT('h8)
	) name2008 (
		_w12018_,
		_w12510_,
		_w12520_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		_w12519_,
		_w12520_,
		_w12521_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		_w12508_,
		_w12521_,
		_w12522_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w12504_,
		_w12509_,
		_w12523_
	);
	LUT2 #(
		.INIT('h4)
	) name2012 (
		_w12522_,
		_w12523_,
		_w12524_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		\rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 ,
		_w12505_,
		_w12525_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w12524_,
		_w12525_,
		_w12526_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		_w12502_,
		_w12526_,
		_w12527_
	);
	LUT2 #(
		.INIT('h4)
	) name2016 (
		_w11869_,
		_w12502_,
		_w12528_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w12527_,
		_w12528_,
		_w12529_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		\rxethmac1_rxstatem1_StateDrop_reg/NET0131 ,
		_w12094_,
		_w12530_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		_w10586_,
		_w12530_,
		_w12531_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		_w12532_
	);
	LUT2 #(
		.INIT('h4)
	) name2021 (
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		\macstatus1_ShortFrame_reg/NET0131 ,
		_w12533_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		\RxAbortRst_reg/NET0131 ,
		\RxAbort_latch_reg/NET0131 ,
		_w12534_
	);
	LUT2 #(
		.INIT('h4)
	) name2023 (
		\macstatus1_InvalidSymbol_reg/NET0131 ,
		\macstatus1_LatchedMRxErr_reg/NET0131 ,
		_w12535_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		\rxethmac1_rxaddrcheck1_RxAbort_reg/NET0131 ,
		_w12532_,
		_w12536_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		_w12533_,
		_w12534_,
		_w12537_
	);
	LUT2 #(
		.INIT('h4)
	) name2026 (
		_w12535_,
		_w12537_,
		_w12538_
	);
	LUT2 #(
		.INIT('h8)
	) name2027 (
		_w12536_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		m_wb_ack_i_pad,
		m_wb_err_i_pad,
		_w12540_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w12540_,
		_w12541_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w12540_,
		_w12542_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		_w12541_,
		_w12542_,
		_w12543_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12543_,
		_w12544_
	);
	LUT2 #(
		.INIT('h2)
	) name2033 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12544_,
		_w12545_
	);
	LUT2 #(
		.INIT('h4)
	) name2034 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w12546_
	);
	LUT2 #(
		.INIT('h2)
	) name2035 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w12547_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		_w12540_,
		_w12546_,
		_w12548_
	);
	LUT2 #(
		.INIT('h4)
	) name2037 (
		_w12547_,
		_w12548_,
		_w12549_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12549_,
		_w12550_
	);
	LUT2 #(
		.INIT('h1)
	) name2039 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w12551_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w12553_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w12552_,
		_w12553_,
		_w12554_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12554_,
		_w12555_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		_w12540_,
		_w12555_,
		_w12556_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		_w12557_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w12557_,
		_w12558_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w12550_,
		_w12558_,
		_w12559_
	);
	LUT2 #(
		.INIT('h4)
	) name2048 (
		_w12545_,
		_w12559_,
		_w12560_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w12556_,
		_w12560_,
		_w12561_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w12557_,
		_w12562_
	);
	LUT2 #(
		.INIT('h1)
	) name2051 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12563_
	);
	LUT2 #(
		.INIT('h4)
	) name2052 (
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w12540_,
		_w12564_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		_w12563_,
		_w12564_,
		_w12565_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w12554_,
		_w12565_,
		_w12566_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12567_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w12563_,
		_w12567_,
		_w12568_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		_w12541_,
		_w12568_,
		_w12569_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w12555_,
		_w12569_,
		_w12570_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w12566_,
		_w12570_,
		_w12571_
	);
	LUT2 #(
		.INIT('h2)
	) name2060 (
		_w12562_,
		_w12571_,
		_w12572_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w12561_,
		_w12572_,
		_w12573_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		_w12574_
	);
	LUT2 #(
		.INIT('h4)
	) name2063 (
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w12574_,
		_w12575_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w12572_,
		_w12575_,
		_w12576_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w12573_,
		_w12576_,
		_w12577_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w12577_,
		_w12578_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		_w12579_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		\m_wb_adr_o[4]_pad ,
		_w12579_,
		_w12580_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		\m_wb_adr_o[5]_pad ,
		_w12580_,
		_w12581_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		\m_wb_adr_o[6]_pad ,
		_w12581_,
		_w12582_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		\m_wb_adr_o[7]_pad ,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\m_wb_adr_o[8]_pad ,
		_w12583_,
		_w12584_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		\m_wb_adr_o[9]_pad ,
		_w12584_,
		_w12585_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		\m_wb_adr_o[10]_pad ,
		_w12585_,
		_w12586_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		\m_wb_adr_o[11]_pad ,
		_w12586_,
		_w12587_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		\m_wb_adr_o[12]_pad ,
		_w12587_,
		_w12588_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		\m_wb_adr_o[13]_pad ,
		\m_wb_adr_o[14]_pad ,
		_w12589_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		_w12588_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		\m_wb_adr_o[15]_pad ,
		_w12590_,
		_w12591_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		\m_wb_adr_o[16]_pad ,
		_w12591_,
		_w12592_
	);
	LUT2 #(
		.INIT('h8)
	) name2081 (
		\m_wb_adr_o[17]_pad ,
		\m_wb_adr_o[18]_pad ,
		_w12593_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w12592_,
		_w12593_,
		_w12594_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		\m_wb_adr_o[19]_pad ,
		_w12594_,
		_w12595_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		\m_wb_adr_o[20]_pad ,
		_w12595_,
		_w12596_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\m_wb_adr_o[21]_pad ,
		_w12596_,
		_w12597_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		\m_wb_adr_o[22]_pad ,
		\m_wb_adr_o[23]_pad ,
		_w12598_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		\m_wb_adr_o[24]_pad ,
		_w12598_,
		_w12599_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		\m_wb_adr_o[25]_pad ,
		\m_wb_adr_o[26]_pad ,
		_w12600_
	);
	LUT2 #(
		.INIT('h8)
	) name2089 (
		_w12599_,
		_w12600_,
		_w12601_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		_w12597_,
		_w12601_,
		_w12602_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		\m_wb_adr_o[27]_pad ,
		\m_wb_adr_o[28]_pad ,
		_w12603_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		_w12602_,
		_w12603_,
		_w12604_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		\m_wb_adr_o[29]_pad ,
		_w12604_,
		_w12605_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		\m_wb_adr_o[30]_pad ,
		_w12605_,
		_w12606_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		_w12607_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w12607_,
		_w12608_
	);
	LUT2 #(
		.INIT('h4)
	) name2097 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w12608_,
		_w12609_
	);
	LUT2 #(
		.INIT('h4)
	) name2098 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12546_,
		_w12610_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w12554_,
		_w12611_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12543_,
		_w12612_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12557_,
		_w12613_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w12540_,
		_w12613_,
		_w12614_
	);
	LUT2 #(
		.INIT('h1)
	) name2103 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12540_,
		_w12615_
	);
	LUT2 #(
		.INIT('h2)
	) name2104 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12546_,
		_w12616_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w12610_,
		_w12615_,
		_w12617_
	);
	LUT2 #(
		.INIT('h4)
	) name2106 (
		_w12616_,
		_w12617_,
		_w12618_
	);
	LUT2 #(
		.INIT('h4)
	) name2107 (
		_w12614_,
		_w12618_,
		_w12619_
	);
	LUT2 #(
		.INIT('h2)
	) name2108 (
		_w12611_,
		_w12612_,
		_w12620_
	);
	LUT2 #(
		.INIT('h8)
	) name2109 (
		_w12619_,
		_w12620_,
		_w12621_
	);
	LUT2 #(
		.INIT('h4)
	) name2110 (
		_w12609_,
		_w12621_,
		_w12622_
	);
	LUT2 #(
		.INIT('h2)
	) name2111 (
		_w12561_,
		_w12575_,
		_w12623_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w12622_,
		_w12623_,
		_w12624_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		\m_wb_adr_o[30]_pad ,
		_w12605_,
		_w12625_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w12606_,
		_w12624_,
		_w12626_
	);
	LUT2 #(
		.INIT('h4)
	) name2115 (
		_w12625_,
		_w12626_,
		_w12627_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w12554_,
		_w12628_
	);
	LUT2 #(
		.INIT('h2)
	) name2117 (
		_w12569_,
		_w12613_,
		_w12629_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		_w12565_,
		_w12629_,
		_w12630_
	);
	LUT2 #(
		.INIT('h2)
	) name2119 (
		_w12628_,
		_w12630_,
		_w12631_
	);
	LUT2 #(
		.INIT('h1)
	) name2120 (
		_w12621_,
		_w12631_,
		_w12632_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		_w12608_,
		_w12631_,
		_w12633_
	);
	LUT2 #(
		.INIT('h1)
	) name2122 (
		_w12632_,
		_w12633_,
		_w12634_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w12634_,
		_w12635_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		_w12573_,
		_w12632_,
		_w12636_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		\m_wb_adr_o[30]_pad ,
		_w12636_,
		_w12637_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		_w12578_,
		_w12635_,
		_w12638_
	);
	LUT2 #(
		.INIT('h4)
	) name2127 (
		_w12637_,
		_w12638_,
		_w12639_
	);
	LUT2 #(
		.INIT('h4)
	) name2128 (
		_w12627_,
		_w12639_,
		_w12640_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w11913_,
		_w12641_
	);
	LUT2 #(
		.INIT('h2)
	) name2130 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h2)
	) name2131 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w11838_,
		_w12643_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w12643_,
		_w12644_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w11827_,
		_w12645_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		\rxethmac1_RxValid_reg/NET0131 ,
		_w12645_,
		_w12646_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w12646_,
		_w12647_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w12642_,
		_w12647_,
		_w12648_
	);
	LUT2 #(
		.INIT('h4)
	) name2137 (
		_w12644_,
		_w12648_,
		_w12649_
	);
	LUT2 #(
		.INIT('h2)
	) name2138 (
		\maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 ,
		_w12649_,
		_w12650_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w12651_
	);
	LUT2 #(
		.INIT('h8)
	) name2140 (
		_w11950_,
		_w12651_,
		_w12652_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		_w12641_,
		_w12652_,
		_w12653_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w12650_,
		_w12653_,
		_w12654_
	);
	LUT2 #(
		.INIT('h8)
	) name2143 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxEn_reg/NET0131 ,
		_w12655_
	);
	LUT2 #(
		.INIT('h8)
	) name2144 (
		\wishbone_TxBDRead_reg/NET0131 ,
		_w12655_,
		_w12656_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w12657_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w12656_,
		_w12657_,
		_w12658_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w12658_,
		_w12659_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w12660_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		_w12661_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		_w12660_,
		_w12661_,
		_w12662_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		_w12663_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w12664_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		_w12663_,
		_w12664_,
		_w12665_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		_w12662_,
		_w12665_,
		_w12666_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		\wishbone_bd_ram_mem3_reg[4][28]/P0001 ,
		_w12666_,
		_w12667_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		_w12668_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w12660_,
		_w12668_,
		_w12669_
	);
	LUT2 #(
		.INIT('h8)
	) name2158 (
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w12670_
	);
	LUT2 #(
		.INIT('h4)
	) name2159 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		_w12671_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w12670_,
		_w12671_,
		_w12672_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		_w12669_,
		_w12672_,
		_w12673_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		\wishbone_bd_ram_mem3_reg[62][28]/P0001 ,
		_w12673_,
		_w12674_
	);
	LUT2 #(
		.INIT('h2)
	) name2163 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		_w12675_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		_w12660_,
		_w12675_,
		_w12676_
	);
	LUT2 #(
		.INIT('h1)
	) name2165 (
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w12677_
	);
	LUT2 #(
		.INIT('h8)
	) name2166 (
		_w12671_,
		_w12677_,
		_w12678_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		_w12676_,
		_w12678_,
		_w12679_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		\wishbone_bd_ram_mem3_reg[18][28]/P0001 ,
		_w12679_,
		_w12680_
	);
	LUT2 #(
		.INIT('h2)
	) name2169 (
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w12681_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		\wishbone_bd_ram_raddr_reg[4]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[5]/NET0131 ,
		_w12682_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		_w12681_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h8)
	) name2172 (
		_w12664_,
		_w12671_,
		_w12684_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		_w12683_,
		_w12684_,
		_w12685_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		\wishbone_bd_ram_mem3_reg[102][28]/P0001 ,
		_w12685_,
		_w12686_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		_w12675_,
		_w12681_,
		_w12687_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		_w12663_,
		_w12677_,
		_w12688_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		_w12687_,
		_w12688_,
		_w12689_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		\wishbone_bd_ram_mem3_reg[80][28]/P0001 ,
		_w12689_,
		_w12690_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		_w12691_
	);
	LUT2 #(
		.INIT('h4)
	) name2180 (
		\wishbone_bd_ram_raddr_reg[2]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[3]/P0001 ,
		_w12692_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w12691_,
		_w12692_,
		_w12693_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w12694_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		_w12682_,
		_w12694_,
		_w12695_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		_w12693_,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		\wishbone_bd_ram_mem3_reg[235][28]/P0001 ,
		_w12696_,
		_w12697_
	);
	LUT2 #(
		.INIT('h8)
	) name2186 (
		_w12671_,
		_w12692_,
		_w12698_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		_w12676_,
		_w12698_,
		_w12699_
	);
	LUT2 #(
		.INIT('h8)
	) name2188 (
		\wishbone_bd_ram_mem3_reg[26][28]/P0001 ,
		_w12699_,
		_w12700_
	);
	LUT2 #(
		.INIT('h8)
	) name2189 (
		_w12677_,
		_w12691_,
		_w12701_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		_w12660_,
		_w12682_,
		_w12702_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		_w12701_,
		_w12702_,
		_w12703_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		\wishbone_bd_ram_mem3_reg[35][28]/P0001 ,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		_w12668_,
		_w12681_,
		_w12705_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		_w12663_,
		_w12692_,
		_w12706_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		_w12705_,
		_w12706_,
		_w12707_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		\wishbone_bd_ram_mem3_reg[120][28]/P0001 ,
		_w12707_,
		_w12708_
	);
	LUT2 #(
		.INIT('h2)
	) name2197 (
		\wishbone_bd_ram_raddr_reg[0]/P0001 ,
		\wishbone_bd_ram_raddr_reg[1]/NET0131 ,
		_w12709_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		_w12664_,
		_w12709_,
		_w12710_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		_w12695_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		\wishbone_bd_ram_mem3_reg[229][28]/P0001 ,
		_w12711_,
		_w12712_
	);
	LUT2 #(
		.INIT('h8)
	) name2201 (
		_w12683_,
		_w12698_,
		_w12713_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		\wishbone_bd_ram_mem3_reg[106][28]/P0001 ,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h8)
	) name2203 (
		_w12705_,
		_w12710_,
		_w12715_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		\wishbone_bd_ram_mem3_reg[117][28]/P0001 ,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		_w12662_,
		_w12688_,
		_w12717_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		\wishbone_bd_ram_mem3_reg[0][28]/P0001 ,
		_w12717_,
		_w12718_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		_w12692_,
		_w12709_,
		_w12719_
	);
	LUT2 #(
		.INIT('h4)
	) name2208 (
		\wishbone_bd_ram_raddr_reg[6]/NET0131 ,
		\wishbone_bd_ram_raddr_reg[7]/NET0131 ,
		_w12720_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		_w12682_,
		_w12720_,
		_w12721_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		_w12719_,
		_w12721_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name2211 (
		\wishbone_bd_ram_mem3_reg[169][28]/P0001 ,
		_w12722_,
		_w12723_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		_w12670_,
		_w12709_,
		_w12724_
	);
	LUT2 #(
		.INIT('h8)
	) name2213 (
		_w12669_,
		_w12724_,
		_w12725_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		\wishbone_bd_ram_mem3_reg[61][28]/P0001 ,
		_w12725_,
		_w12726_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		_w12664_,
		_w12691_,
		_w12727_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		_w12662_,
		_w12727_,
		_w12728_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		\wishbone_bd_ram_mem3_reg[7][28]/P0001 ,
		_w12728_,
		_w12729_
	);
	LUT2 #(
		.INIT('h8)
	) name2218 (
		_w12663_,
		_w12670_,
		_w12730_
	);
	LUT2 #(
		.INIT('h8)
	) name2219 (
		_w12695_,
		_w12730_,
		_w12731_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		\wishbone_bd_ram_mem3_reg[236][28]/P0001 ,
		_w12731_,
		_w12732_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		_w12688_,
		_w12705_,
		_w12733_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		\wishbone_bd_ram_mem3_reg[112][28]/P0001 ,
		_w12733_,
		_w12734_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		_w12684_,
		_w12687_,
		_w12735_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		\wishbone_bd_ram_mem3_reg[86][28]/P0001 ,
		_w12735_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w12661_,
		_w12681_,
		_w12737_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		_w12710_,
		_w12737_,
		_w12738_
	);
	LUT2 #(
		.INIT('h8)
	) name2227 (
		\wishbone_bd_ram_mem3_reg[69][28]/P0001 ,
		_w12738_,
		_w12739_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		_w12675_,
		_w12720_,
		_w12740_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		_w12710_,
		_w12740_,
		_w12741_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		\wishbone_bd_ram_mem3_reg[149][28]/P0001 ,
		_w12741_,
		_w12742_
	);
	LUT2 #(
		.INIT('h8)
	) name2231 (
		_w12670_,
		_w12691_,
		_w12743_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		_w12683_,
		_w12743_,
		_w12744_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		\wishbone_bd_ram_mem3_reg[111][28]/P0001 ,
		_w12744_,
		_w12745_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		_w12668_,
		_w12694_,
		_w12746_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		_w12665_,
		_w12746_,
		_w12747_
	);
	LUT2 #(
		.INIT('h8)
	) name2236 (
		\wishbone_bd_ram_mem3_reg[244][28]/P0001 ,
		_w12747_,
		_w12748_
	);
	LUT2 #(
		.INIT('h8)
	) name2237 (
		_w12683_,
		_w12693_,
		_w12749_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		\wishbone_bd_ram_mem3_reg[107][28]/P0001 ,
		_w12749_,
		_w12750_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		_w12683_,
		_w12719_,
		_w12751_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		\wishbone_bd_ram_mem3_reg[105][28]/P0001 ,
		_w12751_,
		_w12752_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		_w12677_,
		_w12709_,
		_w12753_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		_w12721_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h8)
	) name2243 (
		\wishbone_bd_ram_mem3_reg[161][28]/P0001 ,
		_w12754_,
		_w12755_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		_w12688_,
		_w12740_,
		_w12756_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		\wishbone_bd_ram_mem3_reg[144][28]/P0001 ,
		_w12756_,
		_w12757_
	);
	LUT2 #(
		.INIT('h8)
	) name2246 (
		_w12695_,
		_w12706_,
		_w12758_
	);
	LUT2 #(
		.INIT('h8)
	) name2247 (
		\wishbone_bd_ram_mem3_reg[232][28]/P0001 ,
		_w12758_,
		_w12759_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		_w12661_,
		_w12720_,
		_w12760_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		_w12710_,
		_w12760_,
		_w12761_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		\wishbone_bd_ram_mem3_reg[133][28]/P0001 ,
		_w12761_,
		_w12762_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		_w12684_,
		_w12760_,
		_w12763_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		\wishbone_bd_ram_mem3_reg[134][28]/P0001 ,
		_w12763_,
		_w12764_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		_w12665_,
		_w12695_,
		_w12765_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		\wishbone_bd_ram_mem3_reg[228][28]/P0001 ,
		_w12765_,
		_w12766_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		_w12661_,
		_w12694_,
		_w12767_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		_w12727_,
		_w12767_,
		_w12768_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		\wishbone_bd_ram_mem3_reg[199][28]/P0001 ,
		_w12768_,
		_w12769_
	);
	LUT2 #(
		.INIT('h8)
	) name2258 (
		_w12669_,
		_w12684_,
		_w12770_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		\wishbone_bd_ram_mem3_reg[54][28]/P0001 ,
		_w12770_,
		_w12771_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		_w12678_,
		_w12767_,
		_w12772_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		\wishbone_bd_ram_mem3_reg[194][28]/P0001 ,
		_w12772_,
		_w12773_
	);
	LUT2 #(
		.INIT('h8)
	) name2262 (
		_w12740_,
		_w12743_,
		_w12774_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		\wishbone_bd_ram_mem3_reg[159][28]/P0001 ,
		_w12774_,
		_w12775_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		_w12753_,
		_w12760_,
		_w12776_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		\wishbone_bd_ram_mem3_reg[129][28]/P0001 ,
		_w12776_,
		_w12777_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w12669_,
		_w12706_,
		_w12778_
	);
	LUT2 #(
		.INIT('h8)
	) name2267 (
		\wishbone_bd_ram_mem3_reg[56][28]/P0001 ,
		_w12778_,
		_w12779_
	);
	LUT2 #(
		.INIT('h8)
	) name2268 (
		_w12669_,
		_w12693_,
		_w12780_
	);
	LUT2 #(
		.INIT('h8)
	) name2269 (
		\wishbone_bd_ram_mem3_reg[59][28]/P0001 ,
		_w12780_,
		_w12781_
	);
	LUT2 #(
		.INIT('h8)
	) name2270 (
		_w12668_,
		_w12720_,
		_w12782_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		_w12698_,
		_w12782_,
		_w12783_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		\wishbone_bd_ram_mem3_reg[186][28]/P0001 ,
		_w12783_,
		_w12784_
	);
	LUT2 #(
		.INIT('h8)
	) name2273 (
		_w12669_,
		_w12727_,
		_w12785_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		\wishbone_bd_ram_mem3_reg[55][28]/P0001 ,
		_w12785_,
		_w12786_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		_w12727_,
		_w12782_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name2276 (
		\wishbone_bd_ram_mem3_reg[183][28]/P0001 ,
		_w12787_,
		_w12788_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		_w12706_,
		_w12746_,
		_w12789_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		\wishbone_bd_ram_mem3_reg[248][28]/P0001 ,
		_w12789_,
		_w12790_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w12665_,
		_w12782_,
		_w12791_
	);
	LUT2 #(
		.INIT('h8)
	) name2280 (
		\wishbone_bd_ram_mem3_reg[180][28]/P0001 ,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		_w12688_,
		_w12760_,
		_w12793_
	);
	LUT2 #(
		.INIT('h8)
	) name2282 (
		\wishbone_bd_ram_mem3_reg[128][28]/P0001 ,
		_w12793_,
		_w12794_
	);
	LUT2 #(
		.INIT('h8)
	) name2283 (
		_w12675_,
		_w12694_,
		_w12795_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		_w12665_,
		_w12795_,
		_w12796_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		\wishbone_bd_ram_mem3_reg[212][28]/P0001 ,
		_w12796_,
		_w12797_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		_w12727_,
		_w12737_,
		_w12798_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		\wishbone_bd_ram_mem3_reg[71][28]/P0001 ,
		_w12798_,
		_w12799_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		_w12665_,
		_w12702_,
		_w12800_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		\wishbone_bd_ram_mem3_reg[36][28]/P0001 ,
		_w12800_,
		_w12801_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		_w12724_,
		_w12795_,
		_w12802_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		\wishbone_bd_ram_mem3_reg[221][28]/P0001 ,
		_w12802_,
		_w12803_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w12701_,
		_w12746_,
		_w12804_
	);
	LUT2 #(
		.INIT('h8)
	) name2293 (
		\wishbone_bd_ram_mem3_reg[243][28]/P0001 ,
		_w12804_,
		_w12805_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w12693_,
		_w12795_,
		_w12806_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		\wishbone_bd_ram_mem3_reg[219][28]/P0001 ,
		_w12806_,
		_w12807_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		_w12662_,
		_w12719_,
		_w12808_
	);
	LUT2 #(
		.INIT('h8)
	) name2297 (
		\wishbone_bd_ram_mem3_reg[9][28]/P0001 ,
		_w12808_,
		_w12809_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		_w12706_,
		_w12737_,
		_w12810_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		\wishbone_bd_ram_mem3_reg[72][28]/P0001 ,
		_w12810_,
		_w12811_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		_w12698_,
		_w12737_,
		_w12812_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		\wishbone_bd_ram_mem3_reg[74][28]/P0001 ,
		_w12812_,
		_w12813_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w12693_,
		_w12760_,
		_w12814_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		\wishbone_bd_ram_mem3_reg[139][28]/P0001 ,
		_w12814_,
		_w12815_
	);
	LUT2 #(
		.INIT('h8)
	) name2304 (
		_w12678_,
		_w12683_,
		_w12816_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		\wishbone_bd_ram_mem3_reg[98][28]/P0001 ,
		_w12816_,
		_w12817_
	);
	LUT2 #(
		.INIT('h8)
	) name2306 (
		_w12727_,
		_w12746_,
		_w12818_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		\wishbone_bd_ram_mem3_reg[247][28]/P0001 ,
		_w12818_,
		_w12819_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		_w12684_,
		_w12782_,
		_w12820_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		\wishbone_bd_ram_mem3_reg[182][28]/P0001 ,
		_w12820_,
		_w12821_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		_w12719_,
		_w12767_,
		_w12822_
	);
	LUT2 #(
		.INIT('h8)
	) name2311 (
		\wishbone_bd_ram_mem3_reg[201][28]/P0001 ,
		_w12822_,
		_w12823_
	);
	LUT2 #(
		.INIT('h8)
	) name2312 (
		_w12678_,
		_w12737_,
		_w12824_
	);
	LUT2 #(
		.INIT('h8)
	) name2313 (
		\wishbone_bd_ram_mem3_reg[66][28]/P0001 ,
		_w12824_,
		_w12825_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		_w12693_,
		_w12737_,
		_w12826_
	);
	LUT2 #(
		.INIT('h8)
	) name2315 (
		\wishbone_bd_ram_mem3_reg[75][28]/P0001 ,
		_w12826_,
		_w12827_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		_w12710_,
		_w12782_,
		_w12828_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		\wishbone_bd_ram_mem3_reg[181][28]/P0001 ,
		_w12828_,
		_w12829_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		_w12684_,
		_w12705_,
		_w12830_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		\wishbone_bd_ram_mem3_reg[118][28]/P0001 ,
		_w12830_,
		_w12831_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		_w12684_,
		_w12767_,
		_w12832_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		\wishbone_bd_ram_mem3_reg[198][28]/P0001 ,
		_w12832_,
		_w12833_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		_w12710_,
		_w12767_,
		_w12834_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		\wishbone_bd_ram_mem3_reg[197][28]/P0001 ,
		_w12834_,
		_w12835_
	);
	LUT2 #(
		.INIT('h8)
	) name2324 (
		_w12695_,
		_w12719_,
		_w12836_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		\wishbone_bd_ram_mem3_reg[233][28]/P0001 ,
		_w12836_,
		_w12837_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w12743_,
		_w12795_,
		_w12838_
	);
	LUT2 #(
		.INIT('h8)
	) name2327 (
		\wishbone_bd_ram_mem3_reg[223][28]/P0001 ,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		_w12684_,
		_w12737_,
		_w12840_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		\wishbone_bd_ram_mem3_reg[70][28]/P0001 ,
		_w12840_,
		_w12841_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		_w12698_,
		_w12702_,
		_w12842_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		\wishbone_bd_ram_mem3_reg[42][28]/P0001 ,
		_w12842_,
		_w12843_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		_w12687_,
		_w12743_,
		_w12844_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		\wishbone_bd_ram_mem3_reg[95][28]/P0001 ,
		_w12844_,
		_w12845_
	);
	LUT2 #(
		.INIT('h8)
	) name2334 (
		_w12683_,
		_w12727_,
		_w12846_
	);
	LUT2 #(
		.INIT('h8)
	) name2335 (
		\wishbone_bd_ram_mem3_reg[103][28]/P0001 ,
		_w12846_,
		_w12847_
	);
	LUT2 #(
		.INIT('h8)
	) name2336 (
		_w12676_,
		_w12753_,
		_w12848_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		\wishbone_bd_ram_mem3_reg[17][28]/P0001 ,
		_w12848_,
		_w12849_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		_w12669_,
		_w12743_,
		_w12850_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		\wishbone_bd_ram_mem3_reg[63][28]/P0001 ,
		_w12850_,
		_w12851_
	);
	LUT2 #(
		.INIT('h8)
	) name2340 (
		_w12701_,
		_w12760_,
		_w12852_
	);
	LUT2 #(
		.INIT('h8)
	) name2341 (
		\wishbone_bd_ram_mem3_reg[131][28]/P0001 ,
		_w12852_,
		_w12853_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		_w12721_,
		_w12724_,
		_w12854_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		\wishbone_bd_ram_mem3_reg[173][28]/P0001 ,
		_w12854_,
		_w12855_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		_w12695_,
		_w12727_,
		_w12856_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		\wishbone_bd_ram_mem3_reg[231][28]/P0001 ,
		_w12856_,
		_w12857_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		_w12672_,
		_w12782_,
		_w12858_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		\wishbone_bd_ram_mem3_reg[190][28]/P0001 ,
		_w12858_,
		_w12859_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		_w12687_,
		_w12706_,
		_w12860_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		\wishbone_bd_ram_mem3_reg[88][28]/P0001 ,
		_w12860_,
		_w12861_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		_w12695_,
		_w12743_,
		_w12862_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		\wishbone_bd_ram_mem3_reg[239][28]/P0001 ,
		_w12862_,
		_w12863_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w12688_,
		_w12746_,
		_w12864_
	);
	LUT2 #(
		.INIT('h8)
	) name2353 (
		\wishbone_bd_ram_mem3_reg[240][28]/P0001 ,
		_w12864_,
		_w12865_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		_w12662_,
		_w12701_,
		_w12866_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		\wishbone_bd_ram_mem3_reg[3][28]/P0001 ,
		_w12866_,
		_w12867_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		_w12688_,
		_w12782_,
		_w12868_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		\wishbone_bd_ram_mem3_reg[176][28]/P0001 ,
		_w12868_,
		_w12869_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		_w12698_,
		_w12767_,
		_w12870_
	);
	LUT2 #(
		.INIT('h8)
	) name2359 (
		\wishbone_bd_ram_mem3_reg[202][28]/P0001 ,
		_w12870_,
		_w12871_
	);
	LUT2 #(
		.INIT('h8)
	) name2360 (
		_w12688_,
		_w12721_,
		_w12872_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		\wishbone_bd_ram_mem3_reg[160][28]/P0001 ,
		_w12872_,
		_w12873_
	);
	LUT2 #(
		.INIT('h8)
	) name2362 (
		_w12672_,
		_w12737_,
		_w12874_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		\wishbone_bd_ram_mem3_reg[78][28]/P0001 ,
		_w12874_,
		_w12875_
	);
	LUT2 #(
		.INIT('h8)
	) name2364 (
		_w12665_,
		_w12721_,
		_w12876_
	);
	LUT2 #(
		.INIT('h8)
	) name2365 (
		\wishbone_bd_ram_mem3_reg[164][28]/P0001 ,
		_w12876_,
		_w12877_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		_w12662_,
		_w12710_,
		_w12878_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		\wishbone_bd_ram_mem3_reg[5][28]/P0001 ,
		_w12878_,
		_w12879_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		_w12676_,
		_w12693_,
		_w12880_
	);
	LUT2 #(
		.INIT('h8)
	) name2369 (
		\wishbone_bd_ram_mem3_reg[27][28]/P0001 ,
		_w12880_,
		_w12881_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		_w12701_,
		_w12721_,
		_w12882_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		\wishbone_bd_ram_mem3_reg[163][28]/P0001 ,
		_w12882_,
		_w12883_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		_w12672_,
		_w12702_,
		_w12884_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		\wishbone_bd_ram_mem3_reg[46][28]/P0001 ,
		_w12884_,
		_w12885_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		_w12678_,
		_w12782_,
		_w12886_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		\wishbone_bd_ram_mem3_reg[178][28]/P0001 ,
		_w12886_,
		_w12887_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		_w12683_,
		_w12724_,
		_w12888_
	);
	LUT2 #(
		.INIT('h8)
	) name2377 (
		\wishbone_bd_ram_mem3_reg[109][28]/P0001 ,
		_w12888_,
		_w12889_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		_w12719_,
		_w12740_,
		_w12890_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		\wishbone_bd_ram_mem3_reg[153][28]/P0001 ,
		_w12890_,
		_w12891_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		_w12672_,
		_w12746_,
		_w12892_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		\wishbone_bd_ram_mem3_reg[254][28]/P0001 ,
		_w12892_,
		_w12893_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		_w12730_,
		_w12760_,
		_w12894_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		\wishbone_bd_ram_mem3_reg[140][28]/P0001 ,
		_w12894_,
		_w12895_
	);
	LUT2 #(
		.INIT('h8)
	) name2384 (
		_w12702_,
		_w12730_,
		_w12896_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\wishbone_bd_ram_mem3_reg[44][28]/P0001 ,
		_w12896_,
		_w12897_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		_w12672_,
		_w12740_,
		_w12898_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		\wishbone_bd_ram_mem3_reg[158][28]/P0001 ,
		_w12898_,
		_w12899_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		_w12719_,
		_w12746_,
		_w12900_
	);
	LUT2 #(
		.INIT('h8)
	) name2389 (
		\wishbone_bd_ram_mem3_reg[249][28]/P0001 ,
		_w12900_,
		_w12901_
	);
	LUT2 #(
		.INIT('h8)
	) name2390 (
		_w12688_,
		_w12695_,
		_w12902_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		\wishbone_bd_ram_mem3_reg[224][28]/P0001 ,
		_w12902_,
		_w12903_
	);
	LUT2 #(
		.INIT('h8)
	) name2392 (
		_w12702_,
		_w12743_,
		_w12904_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		\wishbone_bd_ram_mem3_reg[47][28]/P0001 ,
		_w12904_,
		_w12905_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		_w12676_,
		_w12710_,
		_w12906_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		\wishbone_bd_ram_mem3_reg[21][28]/P0001 ,
		_w12906_,
		_w12907_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		_w12702_,
		_w12724_,
		_w12908_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		\wishbone_bd_ram_mem3_reg[45][28]/P0001 ,
		_w12908_,
		_w12909_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		_w12693_,
		_w12721_,
		_w12910_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		\wishbone_bd_ram_mem3_reg[171][28]/P0001 ,
		_w12910_,
		_w12911_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		_w12683_,
		_w12688_,
		_w12912_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		\wishbone_bd_ram_mem3_reg[96][28]/P0001 ,
		_w12912_,
		_w12913_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		_w12678_,
		_w12760_,
		_w12914_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		\wishbone_bd_ram_mem3_reg[130][28]/P0001 ,
		_w12914_,
		_w12915_
	);
	LUT2 #(
		.INIT('h8)
	) name2404 (
		_w12687_,
		_w12701_,
		_w12916_
	);
	LUT2 #(
		.INIT('h8)
	) name2405 (
		\wishbone_bd_ram_mem3_reg[83][28]/P0001 ,
		_w12916_,
		_w12917_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		_w12719_,
		_w12737_,
		_w12918_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		\wishbone_bd_ram_mem3_reg[73][28]/P0001 ,
		_w12918_,
		_w12919_
	);
	LUT2 #(
		.INIT('h8)
	) name2408 (
		_w12662_,
		_w12706_,
		_w12920_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		\wishbone_bd_ram_mem3_reg[8][28]/P0001 ,
		_w12920_,
		_w12921_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		_w12743_,
		_w12760_,
		_w12922_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		\wishbone_bd_ram_mem3_reg[143][28]/P0001 ,
		_w12922_,
		_w12923_
	);
	LUT2 #(
		.INIT('h8)
	) name2412 (
		_w12678_,
		_w12795_,
		_w12924_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		\wishbone_bd_ram_mem3_reg[210][28]/P0001 ,
		_w12924_,
		_w12925_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		_w12724_,
		_w12740_,
		_w12926_
	);
	LUT2 #(
		.INIT('h8)
	) name2415 (
		\wishbone_bd_ram_mem3_reg[157][28]/P0001 ,
		_w12926_,
		_w12927_
	);
	LUT2 #(
		.INIT('h8)
	) name2416 (
		_w12672_,
		_w12760_,
		_w12928_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		\wishbone_bd_ram_mem3_reg[142][28]/P0001 ,
		_w12928_,
		_w12929_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		_w12678_,
		_w12702_,
		_w12930_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		\wishbone_bd_ram_mem3_reg[34][28]/P0001 ,
		_w12930_,
		_w12931_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		_w12678_,
		_w12746_,
		_w12932_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		\wishbone_bd_ram_mem3_reg[242][28]/P0001 ,
		_w12932_,
		_w12933_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		_w12665_,
		_w12687_,
		_w12934_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		\wishbone_bd_ram_mem3_reg[84][28]/P0001 ,
		_w12934_,
		_w12935_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		_w12695_,
		_w12701_,
		_w12936_
	);
	LUT2 #(
		.INIT('h8)
	) name2425 (
		\wishbone_bd_ram_mem3_reg[227][28]/P0001 ,
		_w12936_,
		_w12937_
	);
	LUT2 #(
		.INIT('h8)
	) name2426 (
		_w12688_,
		_w12767_,
		_w12938_
	);
	LUT2 #(
		.INIT('h8)
	) name2427 (
		\wishbone_bd_ram_mem3_reg[192][28]/P0001 ,
		_w12938_,
		_w12939_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		_w12719_,
		_w12782_,
		_w12940_
	);
	LUT2 #(
		.INIT('h8)
	) name2429 (
		\wishbone_bd_ram_mem3_reg[185][28]/P0001 ,
		_w12940_,
		_w12941_
	);
	LUT2 #(
		.INIT('h8)
	) name2430 (
		_w12678_,
		_w12687_,
		_w12942_
	);
	LUT2 #(
		.INIT('h8)
	) name2431 (
		\wishbone_bd_ram_mem3_reg[82][28]/P0001 ,
		_w12942_,
		_w12943_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		_w12721_,
		_w12730_,
		_w12944_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		\wishbone_bd_ram_mem3_reg[172][28]/P0001 ,
		_w12944_,
		_w12945_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		_w12665_,
		_w12737_,
		_w12946_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		\wishbone_bd_ram_mem3_reg[68][28]/P0001 ,
		_w12946_,
		_w12947_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		_w12730_,
		_w12782_,
		_w12948_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		\wishbone_bd_ram_mem3_reg[188][28]/P0001 ,
		_w12948_,
		_w12949_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		_w12687_,
		_w12753_,
		_w12950_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		\wishbone_bd_ram_mem3_reg[81][28]/P0001 ,
		_w12950_,
		_w12951_
	);
	LUT2 #(
		.INIT('h8)
	) name2440 (
		_w12676_,
		_w12724_,
		_w12952_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		\wishbone_bd_ram_mem3_reg[29][28]/P0001 ,
		_w12952_,
		_w12953_
	);
	LUT2 #(
		.INIT('h8)
	) name2442 (
		_w12672_,
		_w12767_,
		_w12954_
	);
	LUT2 #(
		.INIT('h8)
	) name2443 (
		\wishbone_bd_ram_mem3_reg[206][28]/P0001 ,
		_w12954_,
		_w12955_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		_w12705_,
		_w12724_,
		_w12956_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		\wishbone_bd_ram_mem3_reg[125][28]/P0001 ,
		_w12956_,
		_w12957_
	);
	LUT2 #(
		.INIT('h8)
	) name2446 (
		_w12698_,
		_w12760_,
		_w12958_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		\wishbone_bd_ram_mem3_reg[138][28]/P0001 ,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		_w12665_,
		_w12683_,
		_w12960_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		\wishbone_bd_ram_mem3_reg[100][28]/P0001 ,
		_w12960_,
		_w12961_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		_w12698_,
		_w12740_,
		_w12962_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		\wishbone_bd_ram_mem3_reg[154][28]/P0001 ,
		_w12962_,
		_w12963_
	);
	LUT2 #(
		.INIT('h8)
	) name2452 (
		_w12687_,
		_w12719_,
		_w12964_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		\wishbone_bd_ram_mem3_reg[89][28]/P0001 ,
		_w12964_,
		_w12965_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w12706_,
		_w12740_,
		_w12966_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		\wishbone_bd_ram_mem3_reg[152][28]/P0001 ,
		_w12966_,
		_w12967_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		_w12662_,
		_w12684_,
		_w12968_
	);
	LUT2 #(
		.INIT('h8)
	) name2457 (
		\wishbone_bd_ram_mem3_reg[6][28]/P0001 ,
		_w12968_,
		_w12969_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		_w12669_,
		_w12688_,
		_w12970_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\wishbone_bd_ram_mem3_reg[48][28]/P0001 ,
		_w12970_,
		_w12971_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		_w12672_,
		_w12721_,
		_w12972_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		\wishbone_bd_ram_mem3_reg[174][28]/P0001 ,
		_w12972_,
		_w12973_
	);
	LUT2 #(
		.INIT('h8)
	) name2462 (
		_w12727_,
		_w12795_,
		_w12974_
	);
	LUT2 #(
		.INIT('h8)
	) name2463 (
		\wishbone_bd_ram_mem3_reg[215][28]/P0001 ,
		_w12974_,
		_w12975_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		_w12688_,
		_w12737_,
		_w12976_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		\wishbone_bd_ram_mem3_reg[64][28]/P0001 ,
		_w12976_,
		_w12977_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		_w12687_,
		_w12698_,
		_w12978_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		\wishbone_bd_ram_mem3_reg[90][28]/P0001 ,
		_w12978_,
		_w12979_
	);
	LUT2 #(
		.INIT('h8)
	) name2468 (
		_w12702_,
		_w12753_,
		_w12980_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		\wishbone_bd_ram_mem3_reg[33][28]/P0001 ,
		_w12980_,
		_w12981_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w12724_,
		_w12737_,
		_w12982_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		\wishbone_bd_ram_mem3_reg[77][28]/P0001 ,
		_w12982_,
		_w12983_
	);
	LUT2 #(
		.INIT('h8)
	) name2472 (
		_w12684_,
		_w12795_,
		_w12984_
	);
	LUT2 #(
		.INIT('h8)
	) name2473 (
		\wishbone_bd_ram_mem3_reg[214][28]/P0001 ,
		_w12984_,
		_w12985_
	);
	LUT2 #(
		.INIT('h8)
	) name2474 (
		_w12721_,
		_w12727_,
		_w12986_
	);
	LUT2 #(
		.INIT('h8)
	) name2475 (
		\wishbone_bd_ram_mem3_reg[167][28]/P0001 ,
		_w12986_,
		_w12987_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		_w12706_,
		_w12767_,
		_w12988_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		\wishbone_bd_ram_mem3_reg[200][28]/P0001 ,
		_w12988_,
		_w12989_
	);
	LUT2 #(
		.INIT('h8)
	) name2478 (
		_w12695_,
		_w12724_,
		_w12990_
	);
	LUT2 #(
		.INIT('h8)
	) name2479 (
		\wishbone_bd_ram_mem3_reg[237][28]/P0001 ,
		_w12990_,
		_w12991_
	);
	LUT2 #(
		.INIT('h8)
	) name2480 (
		_w12665_,
		_w12760_,
		_w12992_
	);
	LUT2 #(
		.INIT('h8)
	) name2481 (
		\wishbone_bd_ram_mem3_reg[132][28]/P0001 ,
		_w12992_,
		_w12993_
	);
	LUT2 #(
		.INIT('h8)
	) name2482 (
		_w12669_,
		_w12753_,
		_w12994_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		\wishbone_bd_ram_mem3_reg[49][28]/P0001 ,
		_w12994_,
		_w12995_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		_w12753_,
		_w12782_,
		_w12996_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		\wishbone_bd_ram_mem3_reg[177][28]/P0001 ,
		_w12996_,
		_w12997_
	);
	LUT2 #(
		.INIT('h8)
	) name2486 (
		_w12665_,
		_w12705_,
		_w12998_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		\wishbone_bd_ram_mem3_reg[116][28]/P0001 ,
		_w12998_,
		_w12999_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		_w12665_,
		_w12740_,
		_w13000_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		\wishbone_bd_ram_mem3_reg[148][28]/P0001 ,
		_w13000_,
		_w13001_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		_w12710_,
		_w12795_,
		_w13002_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		\wishbone_bd_ram_mem3_reg[213][28]/P0001 ,
		_w13002_,
		_w13003_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		_w12724_,
		_w12760_,
		_w13004_
	);
	LUT2 #(
		.INIT('h8)
	) name2493 (
		\wishbone_bd_ram_mem3_reg[141][28]/P0001 ,
		_w13004_,
		_w13005_
	);
	LUT2 #(
		.INIT('h8)
	) name2494 (
		_w12746_,
		_w12753_,
		_w13006_
	);
	LUT2 #(
		.INIT('h8)
	) name2495 (
		\wishbone_bd_ram_mem3_reg[241][28]/P0001 ,
		_w13006_,
		_w13007_
	);
	LUT2 #(
		.INIT('h8)
	) name2496 (
		_w12676_,
		_w12727_,
		_w13008_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		\wishbone_bd_ram_mem3_reg[23][28]/P0001 ,
		_w13008_,
		_w13009_
	);
	LUT2 #(
		.INIT('h8)
	) name2498 (
		_w12687_,
		_w12730_,
		_w13010_
	);
	LUT2 #(
		.INIT('h8)
	) name2499 (
		\wishbone_bd_ram_mem3_reg[92][28]/P0001 ,
		_w13010_,
		_w13011_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		_w12676_,
		_w12701_,
		_w13012_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\wishbone_bd_ram_mem3_reg[19][28]/P0001 ,
		_w13012_,
		_w13013_
	);
	LUT2 #(
		.INIT('h8)
	) name2502 (
		_w12662_,
		_w12753_,
		_w13014_
	);
	LUT2 #(
		.INIT('h8)
	) name2503 (
		\wishbone_bd_ram_mem3_reg[1][28]/P0001 ,
		_w13014_,
		_w13015_
	);
	LUT2 #(
		.INIT('h8)
	) name2504 (
		_w12687_,
		_w12724_,
		_w13016_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		\wishbone_bd_ram_mem3_reg[93][28]/P0001 ,
		_w13016_,
		_w13017_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w12702_,
		_w12727_,
		_w13018_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		\wishbone_bd_ram_mem3_reg[39][28]/P0001 ,
		_w13018_,
		_w13019_
	);
	LUT2 #(
		.INIT('h8)
	) name2508 (
		_w12669_,
		_w12710_,
		_w13020_
	);
	LUT2 #(
		.INIT('h8)
	) name2509 (
		\wishbone_bd_ram_mem3_reg[53][28]/P0001 ,
		_w13020_,
		_w13021_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		_w12710_,
		_w12746_,
		_w13022_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		\wishbone_bd_ram_mem3_reg[245][28]/P0001 ,
		_w13022_,
		_w13023_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		_w12669_,
		_w12701_,
		_w13024_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		\wishbone_bd_ram_mem3_reg[51][28]/P0001 ,
		_w13024_,
		_w13025_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		_w12705_,
		_w12753_,
		_w13026_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		\wishbone_bd_ram_mem3_reg[113][28]/P0001 ,
		_w13026_,
		_w13027_
	);
	LUT2 #(
		.INIT('h8)
	) name2516 (
		_w12706_,
		_w12795_,
		_w13028_
	);
	LUT2 #(
		.INIT('h8)
	) name2517 (
		\wishbone_bd_ram_mem3_reg[216][28]/P0001 ,
		_w13028_,
		_w13029_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		_w12698_,
		_w12721_,
		_w13030_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		\wishbone_bd_ram_mem3_reg[170][28]/P0001 ,
		_w13030_,
		_w13031_
	);
	LUT2 #(
		.INIT('h8)
	) name2520 (
		_w12688_,
		_w12795_,
		_w13032_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\wishbone_bd_ram_mem3_reg[208][28]/P0001 ,
		_w13032_,
		_w13033_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		_w12743_,
		_w12782_,
		_w13034_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		\wishbone_bd_ram_mem3_reg[191][28]/P0001 ,
		_w13034_,
		_w13035_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		_w12684_,
		_w12695_,
		_w13036_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		\wishbone_bd_ram_mem3_reg[230][28]/P0001 ,
		_w13036_,
		_w13037_
	);
	LUT2 #(
		.INIT('h8)
	) name2526 (
		_w12683_,
		_w12701_,
		_w13038_
	);
	LUT2 #(
		.INIT('h8)
	) name2527 (
		\wishbone_bd_ram_mem3_reg[99][28]/P0001 ,
		_w13038_,
		_w13039_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		_w12684_,
		_w12721_,
		_w13040_
	);
	LUT2 #(
		.INIT('h8)
	) name2529 (
		\wishbone_bd_ram_mem3_reg[166][28]/P0001 ,
		_w13040_,
		_w13041_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		_w12724_,
		_w12782_,
		_w13042_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		\wishbone_bd_ram_mem3_reg[189][28]/P0001 ,
		_w13042_,
		_w13043_
	);
	LUT2 #(
		.INIT('h8)
	) name2532 (
		_w12710_,
		_w12721_,
		_w13044_
	);
	LUT2 #(
		.INIT('h8)
	) name2533 (
		\wishbone_bd_ram_mem3_reg[165][28]/P0001 ,
		_w13044_,
		_w13045_
	);
	LUT2 #(
		.INIT('h8)
	) name2534 (
		_w12672_,
		_w12683_,
		_w13046_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		\wishbone_bd_ram_mem3_reg[110][28]/P0001 ,
		_w13046_,
		_w13047_
	);
	LUT2 #(
		.INIT('h8)
	) name2536 (
		_w12705_,
		_w12727_,
		_w13048_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		\wishbone_bd_ram_mem3_reg[119][28]/P0001 ,
		_w13048_,
		_w13049_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		_w12701_,
		_w12782_,
		_w13050_
	);
	LUT2 #(
		.INIT('h8)
	) name2539 (
		\wishbone_bd_ram_mem3_reg[179][28]/P0001 ,
		_w13050_,
		_w13051_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		_w12702_,
		_w12719_,
		_w13052_
	);
	LUT2 #(
		.INIT('h8)
	) name2541 (
		\wishbone_bd_ram_mem3_reg[41][28]/P0001 ,
		_w13052_,
		_w13053_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		_w12693_,
		_w12746_,
		_w13054_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		\wishbone_bd_ram_mem3_reg[251][28]/P0001 ,
		_w13054_,
		_w13055_
	);
	LUT2 #(
		.INIT('h8)
	) name2544 (
		_w12753_,
		_w12767_,
		_w13056_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		\wishbone_bd_ram_mem3_reg[193][28]/P0001 ,
		_w13056_,
		_w13057_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		_w12705_,
		_w12730_,
		_w13058_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		\wishbone_bd_ram_mem3_reg[124][28]/P0001 ,
		_w13058_,
		_w13059_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		_w12678_,
		_w12740_,
		_w13060_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		\wishbone_bd_ram_mem3_reg[146][28]/P0001 ,
		_w13060_,
		_w13061_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		_w12706_,
		_w12782_,
		_w13062_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		\wishbone_bd_ram_mem3_reg[184][28]/P0001 ,
		_w13062_,
		_w13063_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		_w12706_,
		_w12760_,
		_w13064_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		\wishbone_bd_ram_mem3_reg[136][28]/P0001 ,
		_w13064_,
		_w13065_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		_w12730_,
		_w12795_,
		_w13066_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		\wishbone_bd_ram_mem3_reg[220][28]/P0001 ,
		_w13066_,
		_w13067_
	);
	LUT2 #(
		.INIT('h8)
	) name2556 (
		_w12724_,
		_w12767_,
		_w13068_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		\wishbone_bd_ram_mem3_reg[205][28]/P0001 ,
		_w13068_,
		_w13069_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		_w12669_,
		_w12698_,
		_w13070_
	);
	LUT2 #(
		.INIT('h8)
	) name2559 (
		\wishbone_bd_ram_mem3_reg[58][28]/P0001 ,
		_w13070_,
		_w13071_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		_w12743_,
		_w12746_,
		_w13072_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		\wishbone_bd_ram_mem3_reg[255][28]/P0001 ,
		_w13072_,
		_w13073_
	);
	LUT2 #(
		.INIT('h8)
	) name2562 (
		_w12687_,
		_w12693_,
		_w13074_
	);
	LUT2 #(
		.INIT('h8)
	) name2563 (
		\wishbone_bd_ram_mem3_reg[91][28]/P0001 ,
		_w13074_,
		_w13075_
	);
	LUT2 #(
		.INIT('h8)
	) name2564 (
		_w12684_,
		_w12746_,
		_w13076_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		\wishbone_bd_ram_mem3_reg[246][28]/P0001 ,
		_w13076_,
		_w13077_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		_w12705_,
		_w12719_,
		_w13078_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\wishbone_bd_ram_mem3_reg[121][28]/P0001 ,
		_w13078_,
		_w13079_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		_w12730_,
		_w12746_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		\wishbone_bd_ram_mem3_reg[252][28]/P0001 ,
		_w13080_,
		_w13081_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		_w12665_,
		_w12669_,
		_w13082_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		\wishbone_bd_ram_mem3_reg[52][28]/P0001 ,
		_w13082_,
		_w13083_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		_w12676_,
		_w12706_,
		_w13084_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		\wishbone_bd_ram_mem3_reg[24][28]/P0001 ,
		_w13084_,
		_w13085_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		_w12662_,
		_w12672_,
		_w13086_
	);
	LUT2 #(
		.INIT('h8)
	) name2575 (
		\wishbone_bd_ram_mem3_reg[14][28]/P0001 ,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h8)
	) name2576 (
		_w12662_,
		_w12678_,
		_w13088_
	);
	LUT2 #(
		.INIT('h8)
	) name2577 (
		\wishbone_bd_ram_mem3_reg[2][28]/P0001 ,
		_w13088_,
		_w13089_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		_w12665_,
		_w12767_,
		_w13090_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		\wishbone_bd_ram_mem3_reg[196][28]/P0001 ,
		_w13090_,
		_w13091_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		_w12695_,
		_w12753_,
		_w13092_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		\wishbone_bd_ram_mem3_reg[225][28]/P0001 ,
		_w13092_,
		_w13093_
	);
	LUT2 #(
		.INIT('h8)
	) name2582 (
		_w12672_,
		_w12795_,
		_w13094_
	);
	LUT2 #(
		.INIT('h8)
	) name2583 (
		\wishbone_bd_ram_mem3_reg[222][28]/P0001 ,
		_w13094_,
		_w13095_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		_w12683_,
		_w12753_,
		_w13096_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		\wishbone_bd_ram_mem3_reg[97][28]/P0001 ,
		_w13096_,
		_w13097_
	);
	LUT2 #(
		.INIT('h8)
	) name2586 (
		_w12678_,
		_w12721_,
		_w13098_
	);
	LUT2 #(
		.INIT('h8)
	) name2587 (
		\wishbone_bd_ram_mem3_reg[162][28]/P0001 ,
		_w13098_,
		_w13099_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		_w12724_,
		_w12746_,
		_w13100_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\wishbone_bd_ram_mem3_reg[253][28]/P0001 ,
		_w13100_,
		_w13101_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		_w12702_,
		_w12710_,
		_w13102_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		\wishbone_bd_ram_mem3_reg[37][28]/P0001 ,
		_w13102_,
		_w13103_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		_w12672_,
		_w12676_,
		_w13104_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		\wishbone_bd_ram_mem3_reg[30][28]/P0001 ,
		_w13104_,
		_w13105_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		_w12740_,
		_w12753_,
		_w13106_
	);
	LUT2 #(
		.INIT('h8)
	) name2595 (
		\wishbone_bd_ram_mem3_reg[145][28]/P0001 ,
		_w13106_,
		_w13107_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		_w12676_,
		_w12719_,
		_w13108_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		\wishbone_bd_ram_mem3_reg[25][28]/P0001 ,
		_w13108_,
		_w13109_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w12676_,
		_w12684_,
		_w13110_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		\wishbone_bd_ram_mem3_reg[22][28]/P0001 ,
		_w13110_,
		_w13111_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		_w12701_,
		_w12705_,
		_w13112_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		\wishbone_bd_ram_mem3_reg[115][28]/P0001 ,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		_w12693_,
		_w12705_,
		_w13114_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		\wishbone_bd_ram_mem3_reg[123][28]/P0001 ,
		_w13114_,
		_w13115_
	);
	LUT2 #(
		.INIT('h8)
	) name2604 (
		_w12669_,
		_w12719_,
		_w13116_
	);
	LUT2 #(
		.INIT('h8)
	) name2605 (
		\wishbone_bd_ram_mem3_reg[57][28]/P0001 ,
		_w13116_,
		_w13117_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		_w12662_,
		_w12730_,
		_w13118_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		\wishbone_bd_ram_mem3_reg[12][28]/P0001 ,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		_w12688_,
		_w12702_,
		_w13120_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		\wishbone_bd_ram_mem3_reg[32][28]/P0001 ,
		_w13120_,
		_w13121_
	);
	LUT2 #(
		.INIT('h8)
	) name2610 (
		_w12693_,
		_w12740_,
		_w13122_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		\wishbone_bd_ram_mem3_reg[155][28]/P0001 ,
		_w13122_,
		_w13123_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		_w12727_,
		_w12760_,
		_w13124_
	);
	LUT2 #(
		.INIT('h8)
	) name2613 (
		\wishbone_bd_ram_mem3_reg[135][28]/P0001 ,
		_w13124_,
		_w13125_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		_w12721_,
		_w12743_,
		_w13126_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		\wishbone_bd_ram_mem3_reg[175][28]/P0001 ,
		_w13126_,
		_w13127_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		_w12698_,
		_w12746_,
		_w13128_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		\wishbone_bd_ram_mem3_reg[250][28]/P0001 ,
		_w13128_,
		_w13129_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		_w12698_,
		_w12705_,
		_w13130_
	);
	LUT2 #(
		.INIT('h8)
	) name2619 (
		\wishbone_bd_ram_mem3_reg[122][28]/P0001 ,
		_w13130_,
		_w13131_
	);
	LUT2 #(
		.INIT('h8)
	) name2620 (
		_w12702_,
		_w12706_,
		_w13132_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		\wishbone_bd_ram_mem3_reg[40][28]/P0001 ,
		_w13132_,
		_w13133_
	);
	LUT2 #(
		.INIT('h8)
	) name2622 (
		_w12701_,
		_w12737_,
		_w13134_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		\wishbone_bd_ram_mem3_reg[67][28]/P0001 ,
		_w13134_,
		_w13135_
	);
	LUT2 #(
		.INIT('h8)
	) name2624 (
		_w12684_,
		_w12740_,
		_w13136_
	);
	LUT2 #(
		.INIT('h8)
	) name2625 (
		\wishbone_bd_ram_mem3_reg[150][28]/P0001 ,
		_w13136_,
		_w13137_
	);
	LUT2 #(
		.INIT('h8)
	) name2626 (
		_w12678_,
		_w12695_,
		_w13138_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		\wishbone_bd_ram_mem3_reg[226][28]/P0001 ,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		_w12676_,
		_w12688_,
		_w13140_
	);
	LUT2 #(
		.INIT('h8)
	) name2629 (
		\wishbone_bd_ram_mem3_reg[16][28]/P0001 ,
		_w13140_,
		_w13141_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		_w12727_,
		_w12740_,
		_w13142_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		\wishbone_bd_ram_mem3_reg[151][28]/P0001 ,
		_w13142_,
		_w13143_
	);
	LUT2 #(
		.INIT('h8)
	) name2632 (
		_w12701_,
		_w12767_,
		_w13144_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		\wishbone_bd_ram_mem3_reg[195][28]/P0001 ,
		_w13144_,
		_w13145_
	);
	LUT2 #(
		.INIT('h8)
	) name2634 (
		_w12701_,
		_w12740_,
		_w13146_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		\wishbone_bd_ram_mem3_reg[147][28]/P0001 ,
		_w13146_,
		_w13147_
	);
	LUT2 #(
		.INIT('h8)
	) name2636 (
		_w12683_,
		_w12706_,
		_w13148_
	);
	LUT2 #(
		.INIT('h8)
	) name2637 (
		\wishbone_bd_ram_mem3_reg[104][28]/P0001 ,
		_w13148_,
		_w13149_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		_w12669_,
		_w12678_,
		_w13150_
	);
	LUT2 #(
		.INIT('h8)
	) name2639 (
		\wishbone_bd_ram_mem3_reg[50][28]/P0001 ,
		_w13150_,
		_w13151_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		_w12753_,
		_w12795_,
		_w13152_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		\wishbone_bd_ram_mem3_reg[209][28]/P0001 ,
		_w13152_,
		_w13153_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		_w12687_,
		_w12727_,
		_w13154_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		\wishbone_bd_ram_mem3_reg[87][28]/P0001 ,
		_w13154_,
		_w13155_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		_w12683_,
		_w12730_,
		_w13156_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		\wishbone_bd_ram_mem3_reg[108][28]/P0001 ,
		_w13156_,
		_w13157_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		_w12693_,
		_w12767_,
		_w13158_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\wishbone_bd_ram_mem3_reg[203][28]/P0001 ,
		_w13158_,
		_w13159_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		_w12672_,
		_w12695_,
		_w13160_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		\wishbone_bd_ram_mem3_reg[238][28]/P0001 ,
		_w13160_,
		_w13161_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		_w12730_,
		_w12767_,
		_w13162_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		\wishbone_bd_ram_mem3_reg[204][28]/P0001 ,
		_w13162_,
		_w13163_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		_w12705_,
		_w12743_,
		_w13164_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		\wishbone_bd_ram_mem3_reg[127][28]/P0001 ,
		_w13164_,
		_w13165_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		_w12701_,
		_w12795_,
		_w13166_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		\wishbone_bd_ram_mem3_reg[211][28]/P0001 ,
		_w13166_,
		_w13167_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		_w12719_,
		_w12760_,
		_w13168_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		\wishbone_bd_ram_mem3_reg[137][28]/P0001 ,
		_w13168_,
		_w13169_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		_w12676_,
		_w12730_,
		_w13170_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		\wishbone_bd_ram_mem3_reg[28][28]/P0001 ,
		_w13170_,
		_w13171_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		_w12662_,
		_w12698_,
		_w13172_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		\wishbone_bd_ram_mem3_reg[10][28]/P0001 ,
		_w13172_,
		_w13173_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		_w12665_,
		_w12676_,
		_w13174_
	);
	LUT2 #(
		.INIT('h8)
	) name2663 (
		\wishbone_bd_ram_mem3_reg[20][28]/P0001 ,
		_w13174_,
		_w13175_
	);
	LUT2 #(
		.INIT('h8)
	) name2664 (
		_w12737_,
		_w12753_,
		_w13176_
	);
	LUT2 #(
		.INIT('h8)
	) name2665 (
		\wishbone_bd_ram_mem3_reg[65][28]/P0001 ,
		_w13176_,
		_w13177_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		_w12662_,
		_w12724_,
		_w13178_
	);
	LUT2 #(
		.INIT('h8)
	) name2667 (
		\wishbone_bd_ram_mem3_reg[13][28]/P0001 ,
		_w13178_,
		_w13179_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		_w12743_,
		_w12767_,
		_w13180_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		\wishbone_bd_ram_mem3_reg[207][28]/P0001 ,
		_w13180_,
		_w13181_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		_w12684_,
		_w12702_,
		_w13182_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		\wishbone_bd_ram_mem3_reg[38][28]/P0001 ,
		_w13182_,
		_w13183_
	);
	LUT2 #(
		.INIT('h8)
	) name2672 (
		_w12730_,
		_w12737_,
		_w13184_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		\wishbone_bd_ram_mem3_reg[76][28]/P0001 ,
		_w13184_,
		_w13185_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		_w12672_,
		_w12687_,
		_w13186_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		\wishbone_bd_ram_mem3_reg[94][28]/P0001 ,
		_w13186_,
		_w13187_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		_w12719_,
		_w12795_,
		_w13188_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		\wishbone_bd_ram_mem3_reg[217][28]/P0001 ,
		_w13188_,
		_w13189_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		_w12730_,
		_w12740_,
		_w13190_
	);
	LUT2 #(
		.INIT('h8)
	) name2679 (
		\wishbone_bd_ram_mem3_reg[156][28]/P0001 ,
		_w13190_,
		_w13191_
	);
	LUT2 #(
		.INIT('h8)
	) name2680 (
		_w12683_,
		_w12710_,
		_w13192_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		\wishbone_bd_ram_mem3_reg[101][28]/P0001 ,
		_w13192_,
		_w13193_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		_w12662_,
		_w12693_,
		_w13194_
	);
	LUT2 #(
		.INIT('h8)
	) name2683 (
		\wishbone_bd_ram_mem3_reg[11][28]/P0001 ,
		_w13194_,
		_w13195_
	);
	LUT2 #(
		.INIT('h8)
	) name2684 (
		_w12693_,
		_w12782_,
		_w13196_
	);
	LUT2 #(
		.INIT('h8)
	) name2685 (
		\wishbone_bd_ram_mem3_reg[187][28]/P0001 ,
		_w13196_,
		_w13197_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		_w12676_,
		_w12743_,
		_w13198_
	);
	LUT2 #(
		.INIT('h8)
	) name2687 (
		\wishbone_bd_ram_mem3_reg[31][28]/P0001 ,
		_w13198_,
		_w13199_
	);
	LUT2 #(
		.INIT('h8)
	) name2688 (
		_w12693_,
		_w12702_,
		_w13200_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		\wishbone_bd_ram_mem3_reg[43][28]/P0001 ,
		_w13200_,
		_w13201_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		_w12678_,
		_w12705_,
		_w13202_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		\wishbone_bd_ram_mem3_reg[114][28]/P0001 ,
		_w13202_,
		_w13203_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		_w12669_,
		_w12730_,
		_w13204_
	);
	LUT2 #(
		.INIT('h8)
	) name2693 (
		\wishbone_bd_ram_mem3_reg[60][28]/P0001 ,
		_w13204_,
		_w13205_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		_w12698_,
		_w12795_,
		_w13206_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		\wishbone_bd_ram_mem3_reg[218][28]/P0001 ,
		_w13206_,
		_w13207_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		_w12706_,
		_w12721_,
		_w13208_
	);
	LUT2 #(
		.INIT('h8)
	) name2697 (
		\wishbone_bd_ram_mem3_reg[168][28]/P0001 ,
		_w13208_,
		_w13209_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		_w12662_,
		_w12743_,
		_w13210_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		\wishbone_bd_ram_mem3_reg[15][28]/P0001 ,
		_w13210_,
		_w13211_
	);
	LUT2 #(
		.INIT('h8)
	) name2700 (
		_w12737_,
		_w12743_,
		_w13212_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		\wishbone_bd_ram_mem3_reg[79][28]/P0001 ,
		_w13212_,
		_w13213_
	);
	LUT2 #(
		.INIT('h8)
	) name2702 (
		_w12695_,
		_w12698_,
		_w13214_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		\wishbone_bd_ram_mem3_reg[234][28]/P0001 ,
		_w13214_,
		_w13215_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w12687_,
		_w12710_,
		_w13216_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		\wishbone_bd_ram_mem3_reg[85][28]/P0001 ,
		_w13216_,
		_w13217_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		_w12672_,
		_w12705_,
		_w13218_
	);
	LUT2 #(
		.INIT('h8)
	) name2707 (
		\wishbone_bd_ram_mem3_reg[126][28]/P0001 ,
		_w13218_,
		_w13219_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w12667_,
		_w12674_,
		_w13220_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w12680_,
		_w12686_,
		_w13221_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w12690_,
		_w12697_,
		_w13222_
	);
	LUT2 #(
		.INIT('h1)
	) name2711 (
		_w12700_,
		_w12704_,
		_w13223_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w12708_,
		_w12712_,
		_w13224_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w12714_,
		_w12716_,
		_w13225_
	);
	LUT2 #(
		.INIT('h1)
	) name2714 (
		_w12718_,
		_w12723_,
		_w13226_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w12726_,
		_w12729_,
		_w13227_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w12732_,
		_w12734_,
		_w13228_
	);
	LUT2 #(
		.INIT('h1)
	) name2717 (
		_w12736_,
		_w12739_,
		_w13229_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w12742_,
		_w12745_,
		_w13230_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w12748_,
		_w12750_,
		_w13231_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w12752_,
		_w12755_,
		_w13232_
	);
	LUT2 #(
		.INIT('h1)
	) name2721 (
		_w12757_,
		_w12759_,
		_w13233_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w12762_,
		_w12764_,
		_w13234_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w12766_,
		_w12769_,
		_w13235_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w12771_,
		_w12773_,
		_w13236_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		_w12775_,
		_w12777_,
		_w13237_
	);
	LUT2 #(
		.INIT('h1)
	) name2726 (
		_w12779_,
		_w12781_,
		_w13238_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w12784_,
		_w12786_,
		_w13239_
	);
	LUT2 #(
		.INIT('h1)
	) name2728 (
		_w12788_,
		_w12790_,
		_w13240_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w12792_,
		_w12794_,
		_w13241_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w12797_,
		_w12799_,
		_w13242_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		_w12801_,
		_w12803_,
		_w13243_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		_w12805_,
		_w12807_,
		_w13244_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w12809_,
		_w12811_,
		_w13245_
	);
	LUT2 #(
		.INIT('h1)
	) name2734 (
		_w12813_,
		_w12815_,
		_w13246_
	);
	LUT2 #(
		.INIT('h1)
	) name2735 (
		_w12817_,
		_w12819_,
		_w13247_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w12821_,
		_w12823_,
		_w13248_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		_w12825_,
		_w12827_,
		_w13249_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w12829_,
		_w12831_,
		_w13250_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w12833_,
		_w12835_,
		_w13251_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w12837_,
		_w12839_,
		_w13252_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w12841_,
		_w12843_,
		_w13253_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w12845_,
		_w12847_,
		_w13254_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		_w12849_,
		_w12851_,
		_w13255_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w12853_,
		_w12855_,
		_w13256_
	);
	LUT2 #(
		.INIT('h1)
	) name2745 (
		_w12857_,
		_w12859_,
		_w13257_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w12861_,
		_w12863_,
		_w13258_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		_w12865_,
		_w12867_,
		_w13259_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w12869_,
		_w12871_,
		_w13260_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w12873_,
		_w12875_,
		_w13261_
	);
	LUT2 #(
		.INIT('h1)
	) name2750 (
		_w12877_,
		_w12879_,
		_w13262_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w12881_,
		_w12883_,
		_w13263_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w12885_,
		_w12887_,
		_w13264_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w12889_,
		_w12891_,
		_w13265_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w12893_,
		_w12895_,
		_w13266_
	);
	LUT2 #(
		.INIT('h1)
	) name2755 (
		_w12897_,
		_w12899_,
		_w13267_
	);
	LUT2 #(
		.INIT('h1)
	) name2756 (
		_w12901_,
		_w12903_,
		_w13268_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w12905_,
		_w12907_,
		_w13269_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w12909_,
		_w12911_,
		_w13270_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		_w12913_,
		_w12915_,
		_w13271_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w12917_,
		_w12919_,
		_w13272_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w12921_,
		_w12923_,
		_w13273_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		_w12925_,
		_w12927_,
		_w13274_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w12929_,
		_w12931_,
		_w13275_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w12933_,
		_w12935_,
		_w13276_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w12937_,
		_w12939_,
		_w13277_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w12941_,
		_w12943_,
		_w13278_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w12945_,
		_w12947_,
		_w13279_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w12949_,
		_w12951_,
		_w13280_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w12953_,
		_w12955_,
		_w13281_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w12957_,
		_w12959_,
		_w13282_
	);
	LUT2 #(
		.INIT('h1)
	) name2771 (
		_w12961_,
		_w12963_,
		_w13283_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w12965_,
		_w12967_,
		_w13284_
	);
	LUT2 #(
		.INIT('h1)
	) name2773 (
		_w12969_,
		_w12971_,
		_w13285_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		_w12973_,
		_w12975_,
		_w13286_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w12977_,
		_w12979_,
		_w13287_
	);
	LUT2 #(
		.INIT('h1)
	) name2776 (
		_w12981_,
		_w12983_,
		_w13288_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		_w12985_,
		_w12987_,
		_w13289_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w12989_,
		_w12991_,
		_w13290_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w12993_,
		_w12995_,
		_w13291_
	);
	LUT2 #(
		.INIT('h1)
	) name2780 (
		_w12997_,
		_w12999_,
		_w13292_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w13001_,
		_w13003_,
		_w13293_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w13005_,
		_w13007_,
		_w13294_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		_w13009_,
		_w13011_,
		_w13295_
	);
	LUT2 #(
		.INIT('h1)
	) name2784 (
		_w13013_,
		_w13015_,
		_w13296_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w13017_,
		_w13019_,
		_w13297_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w13021_,
		_w13023_,
		_w13298_
	);
	LUT2 #(
		.INIT('h1)
	) name2787 (
		_w13025_,
		_w13027_,
		_w13299_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w13029_,
		_w13031_,
		_w13300_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w13033_,
		_w13035_,
		_w13301_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w13037_,
		_w13039_,
		_w13302_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w13041_,
		_w13043_,
		_w13303_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		_w13045_,
		_w13047_,
		_w13304_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		_w13049_,
		_w13051_,
		_w13305_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w13053_,
		_w13055_,
		_w13306_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w13057_,
		_w13059_,
		_w13307_
	);
	LUT2 #(
		.INIT('h1)
	) name2796 (
		_w13061_,
		_w13063_,
		_w13308_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w13065_,
		_w13067_,
		_w13309_
	);
	LUT2 #(
		.INIT('h1)
	) name2798 (
		_w13069_,
		_w13071_,
		_w13310_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		_w13073_,
		_w13075_,
		_w13311_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w13077_,
		_w13079_,
		_w13312_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w13081_,
		_w13083_,
		_w13313_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w13085_,
		_w13087_,
		_w13314_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w13089_,
		_w13091_,
		_w13315_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		_w13093_,
		_w13095_,
		_w13316_
	);
	LUT2 #(
		.INIT('h1)
	) name2805 (
		_w13097_,
		_w13099_,
		_w13317_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w13101_,
		_w13103_,
		_w13318_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w13105_,
		_w13107_,
		_w13319_
	);
	LUT2 #(
		.INIT('h1)
	) name2808 (
		_w13109_,
		_w13111_,
		_w13320_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w13113_,
		_w13115_,
		_w13321_
	);
	LUT2 #(
		.INIT('h1)
	) name2810 (
		_w13117_,
		_w13119_,
		_w13322_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w13121_,
		_w13123_,
		_w13323_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w13125_,
		_w13127_,
		_w13324_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w13129_,
		_w13131_,
		_w13325_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w13133_,
		_w13135_,
		_w13326_
	);
	LUT2 #(
		.INIT('h1)
	) name2815 (
		_w13137_,
		_w13139_,
		_w13327_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w13141_,
		_w13143_,
		_w13328_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w13145_,
		_w13147_,
		_w13329_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w13149_,
		_w13151_,
		_w13330_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w13153_,
		_w13155_,
		_w13331_
	);
	LUT2 #(
		.INIT('h1)
	) name2820 (
		_w13157_,
		_w13159_,
		_w13332_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w13161_,
		_w13163_,
		_w13333_
	);
	LUT2 #(
		.INIT('h1)
	) name2822 (
		_w13165_,
		_w13167_,
		_w13334_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		_w13169_,
		_w13171_,
		_w13335_
	);
	LUT2 #(
		.INIT('h1)
	) name2824 (
		_w13173_,
		_w13175_,
		_w13336_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w13177_,
		_w13179_,
		_w13337_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w13181_,
		_w13183_,
		_w13338_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w13185_,
		_w13187_,
		_w13339_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w13189_,
		_w13191_,
		_w13340_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w13193_,
		_w13195_,
		_w13341_
	);
	LUT2 #(
		.INIT('h1)
	) name2830 (
		_w13197_,
		_w13199_,
		_w13342_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w13201_,
		_w13203_,
		_w13343_
	);
	LUT2 #(
		.INIT('h1)
	) name2832 (
		_w13205_,
		_w13207_,
		_w13344_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w13209_,
		_w13211_,
		_w13345_
	);
	LUT2 #(
		.INIT('h1)
	) name2834 (
		_w13213_,
		_w13215_,
		_w13346_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w13217_,
		_w13219_,
		_w13347_
	);
	LUT2 #(
		.INIT('h8)
	) name2836 (
		_w13346_,
		_w13347_,
		_w13348_
	);
	LUT2 #(
		.INIT('h8)
	) name2837 (
		_w13344_,
		_w13345_,
		_w13349_
	);
	LUT2 #(
		.INIT('h8)
	) name2838 (
		_w13342_,
		_w13343_,
		_w13350_
	);
	LUT2 #(
		.INIT('h8)
	) name2839 (
		_w13340_,
		_w13341_,
		_w13351_
	);
	LUT2 #(
		.INIT('h8)
	) name2840 (
		_w13338_,
		_w13339_,
		_w13352_
	);
	LUT2 #(
		.INIT('h8)
	) name2841 (
		_w13336_,
		_w13337_,
		_w13353_
	);
	LUT2 #(
		.INIT('h8)
	) name2842 (
		_w13334_,
		_w13335_,
		_w13354_
	);
	LUT2 #(
		.INIT('h8)
	) name2843 (
		_w13332_,
		_w13333_,
		_w13355_
	);
	LUT2 #(
		.INIT('h8)
	) name2844 (
		_w13330_,
		_w13331_,
		_w13356_
	);
	LUT2 #(
		.INIT('h8)
	) name2845 (
		_w13328_,
		_w13329_,
		_w13357_
	);
	LUT2 #(
		.INIT('h8)
	) name2846 (
		_w13326_,
		_w13327_,
		_w13358_
	);
	LUT2 #(
		.INIT('h8)
	) name2847 (
		_w13324_,
		_w13325_,
		_w13359_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		_w13322_,
		_w13323_,
		_w13360_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		_w13320_,
		_w13321_,
		_w13361_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		_w13318_,
		_w13319_,
		_w13362_
	);
	LUT2 #(
		.INIT('h8)
	) name2851 (
		_w13316_,
		_w13317_,
		_w13363_
	);
	LUT2 #(
		.INIT('h8)
	) name2852 (
		_w13314_,
		_w13315_,
		_w13364_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		_w13312_,
		_w13313_,
		_w13365_
	);
	LUT2 #(
		.INIT('h8)
	) name2854 (
		_w13310_,
		_w13311_,
		_w13366_
	);
	LUT2 #(
		.INIT('h8)
	) name2855 (
		_w13308_,
		_w13309_,
		_w13367_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		_w13306_,
		_w13307_,
		_w13368_
	);
	LUT2 #(
		.INIT('h8)
	) name2857 (
		_w13304_,
		_w13305_,
		_w13369_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		_w13302_,
		_w13303_,
		_w13370_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		_w13300_,
		_w13301_,
		_w13371_
	);
	LUT2 #(
		.INIT('h8)
	) name2860 (
		_w13298_,
		_w13299_,
		_w13372_
	);
	LUT2 #(
		.INIT('h8)
	) name2861 (
		_w13296_,
		_w13297_,
		_w13373_
	);
	LUT2 #(
		.INIT('h8)
	) name2862 (
		_w13294_,
		_w13295_,
		_w13374_
	);
	LUT2 #(
		.INIT('h8)
	) name2863 (
		_w13292_,
		_w13293_,
		_w13375_
	);
	LUT2 #(
		.INIT('h8)
	) name2864 (
		_w13290_,
		_w13291_,
		_w13376_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w13288_,
		_w13289_,
		_w13377_
	);
	LUT2 #(
		.INIT('h8)
	) name2866 (
		_w13286_,
		_w13287_,
		_w13378_
	);
	LUT2 #(
		.INIT('h8)
	) name2867 (
		_w13284_,
		_w13285_,
		_w13379_
	);
	LUT2 #(
		.INIT('h8)
	) name2868 (
		_w13282_,
		_w13283_,
		_w13380_
	);
	LUT2 #(
		.INIT('h8)
	) name2869 (
		_w13280_,
		_w13281_,
		_w13381_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w13278_,
		_w13279_,
		_w13382_
	);
	LUT2 #(
		.INIT('h8)
	) name2871 (
		_w13276_,
		_w13277_,
		_w13383_
	);
	LUT2 #(
		.INIT('h8)
	) name2872 (
		_w13274_,
		_w13275_,
		_w13384_
	);
	LUT2 #(
		.INIT('h8)
	) name2873 (
		_w13272_,
		_w13273_,
		_w13385_
	);
	LUT2 #(
		.INIT('h8)
	) name2874 (
		_w13270_,
		_w13271_,
		_w13386_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		_w13268_,
		_w13269_,
		_w13387_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		_w13266_,
		_w13267_,
		_w13388_
	);
	LUT2 #(
		.INIT('h8)
	) name2877 (
		_w13264_,
		_w13265_,
		_w13389_
	);
	LUT2 #(
		.INIT('h8)
	) name2878 (
		_w13262_,
		_w13263_,
		_w13390_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w13260_,
		_w13261_,
		_w13391_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		_w13258_,
		_w13259_,
		_w13392_
	);
	LUT2 #(
		.INIT('h8)
	) name2881 (
		_w13256_,
		_w13257_,
		_w13393_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w13254_,
		_w13255_,
		_w13394_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		_w13252_,
		_w13253_,
		_w13395_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w13250_,
		_w13251_,
		_w13396_
	);
	LUT2 #(
		.INIT('h8)
	) name2885 (
		_w13248_,
		_w13249_,
		_w13397_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		_w13246_,
		_w13247_,
		_w13398_
	);
	LUT2 #(
		.INIT('h8)
	) name2887 (
		_w13244_,
		_w13245_,
		_w13399_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		_w13242_,
		_w13243_,
		_w13400_
	);
	LUT2 #(
		.INIT('h8)
	) name2889 (
		_w13240_,
		_w13241_,
		_w13401_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		_w13238_,
		_w13239_,
		_w13402_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		_w13236_,
		_w13237_,
		_w13403_
	);
	LUT2 #(
		.INIT('h8)
	) name2892 (
		_w13234_,
		_w13235_,
		_w13404_
	);
	LUT2 #(
		.INIT('h8)
	) name2893 (
		_w13232_,
		_w13233_,
		_w13405_
	);
	LUT2 #(
		.INIT('h8)
	) name2894 (
		_w13230_,
		_w13231_,
		_w13406_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w13228_,
		_w13229_,
		_w13407_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w13226_,
		_w13227_,
		_w13408_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		_w13224_,
		_w13225_,
		_w13409_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		_w13222_,
		_w13223_,
		_w13410_
	);
	LUT2 #(
		.INIT('h8)
	) name2899 (
		_w13220_,
		_w13221_,
		_w13411_
	);
	LUT2 #(
		.INIT('h8)
	) name2900 (
		_w13410_,
		_w13411_,
		_w13412_
	);
	LUT2 #(
		.INIT('h8)
	) name2901 (
		_w13408_,
		_w13409_,
		_w13413_
	);
	LUT2 #(
		.INIT('h8)
	) name2902 (
		_w13406_,
		_w13407_,
		_w13414_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w13404_,
		_w13405_,
		_w13415_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w13402_,
		_w13403_,
		_w13416_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		_w13400_,
		_w13401_,
		_w13417_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		_w13398_,
		_w13399_,
		_w13418_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		_w13396_,
		_w13397_,
		_w13419_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		_w13394_,
		_w13395_,
		_w13420_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		_w13392_,
		_w13393_,
		_w13421_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w13390_,
		_w13391_,
		_w13422_
	);
	LUT2 #(
		.INIT('h8)
	) name2911 (
		_w13388_,
		_w13389_,
		_w13423_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		_w13386_,
		_w13387_,
		_w13424_
	);
	LUT2 #(
		.INIT('h8)
	) name2913 (
		_w13384_,
		_w13385_,
		_w13425_
	);
	LUT2 #(
		.INIT('h8)
	) name2914 (
		_w13382_,
		_w13383_,
		_w13426_
	);
	LUT2 #(
		.INIT('h8)
	) name2915 (
		_w13380_,
		_w13381_,
		_w13427_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		_w13378_,
		_w13379_,
		_w13428_
	);
	LUT2 #(
		.INIT('h8)
	) name2917 (
		_w13376_,
		_w13377_,
		_w13429_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		_w13374_,
		_w13375_,
		_w13430_
	);
	LUT2 #(
		.INIT('h8)
	) name2919 (
		_w13372_,
		_w13373_,
		_w13431_
	);
	LUT2 #(
		.INIT('h8)
	) name2920 (
		_w13370_,
		_w13371_,
		_w13432_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		_w13368_,
		_w13369_,
		_w13433_
	);
	LUT2 #(
		.INIT('h8)
	) name2922 (
		_w13366_,
		_w13367_,
		_w13434_
	);
	LUT2 #(
		.INIT('h8)
	) name2923 (
		_w13364_,
		_w13365_,
		_w13435_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		_w13362_,
		_w13363_,
		_w13436_
	);
	LUT2 #(
		.INIT('h8)
	) name2925 (
		_w13360_,
		_w13361_,
		_w13437_
	);
	LUT2 #(
		.INIT('h8)
	) name2926 (
		_w13358_,
		_w13359_,
		_w13438_
	);
	LUT2 #(
		.INIT('h8)
	) name2927 (
		_w13356_,
		_w13357_,
		_w13439_
	);
	LUT2 #(
		.INIT('h8)
	) name2928 (
		_w13354_,
		_w13355_,
		_w13440_
	);
	LUT2 #(
		.INIT('h8)
	) name2929 (
		_w13352_,
		_w13353_,
		_w13441_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		_w13350_,
		_w13351_,
		_w13442_
	);
	LUT2 #(
		.INIT('h8)
	) name2931 (
		_w13348_,
		_w13349_,
		_w13443_
	);
	LUT2 #(
		.INIT('h8)
	) name2932 (
		_w13442_,
		_w13443_,
		_w13444_
	);
	LUT2 #(
		.INIT('h8)
	) name2933 (
		_w13440_,
		_w13441_,
		_w13445_
	);
	LUT2 #(
		.INIT('h8)
	) name2934 (
		_w13438_,
		_w13439_,
		_w13446_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		_w13436_,
		_w13437_,
		_w13447_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		_w13434_,
		_w13435_,
		_w13448_
	);
	LUT2 #(
		.INIT('h8)
	) name2937 (
		_w13432_,
		_w13433_,
		_w13449_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w13430_,
		_w13431_,
		_w13450_
	);
	LUT2 #(
		.INIT('h8)
	) name2939 (
		_w13428_,
		_w13429_,
		_w13451_
	);
	LUT2 #(
		.INIT('h8)
	) name2940 (
		_w13426_,
		_w13427_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		_w13424_,
		_w13425_,
		_w13453_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		_w13422_,
		_w13423_,
		_w13454_
	);
	LUT2 #(
		.INIT('h8)
	) name2943 (
		_w13420_,
		_w13421_,
		_w13455_
	);
	LUT2 #(
		.INIT('h8)
	) name2944 (
		_w13418_,
		_w13419_,
		_w13456_
	);
	LUT2 #(
		.INIT('h8)
	) name2945 (
		_w13416_,
		_w13417_,
		_w13457_
	);
	LUT2 #(
		.INIT('h8)
	) name2946 (
		_w13414_,
		_w13415_,
		_w13458_
	);
	LUT2 #(
		.INIT('h8)
	) name2947 (
		_w13412_,
		_w13413_,
		_w13459_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		_w13458_,
		_w13459_,
		_w13460_
	);
	LUT2 #(
		.INIT('h8)
	) name2949 (
		_w13456_,
		_w13457_,
		_w13461_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		_w13454_,
		_w13455_,
		_w13462_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		_w13452_,
		_w13453_,
		_w13463_
	);
	LUT2 #(
		.INIT('h8)
	) name2952 (
		_w13450_,
		_w13451_,
		_w13464_
	);
	LUT2 #(
		.INIT('h8)
	) name2953 (
		_w13448_,
		_w13449_,
		_w13465_
	);
	LUT2 #(
		.INIT('h8)
	) name2954 (
		_w13446_,
		_w13447_,
		_w13466_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		_w13444_,
		_w13445_,
		_w13467_
	);
	LUT2 #(
		.INIT('h8)
	) name2956 (
		_w13466_,
		_w13467_,
		_w13468_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		_w13464_,
		_w13465_,
		_w13469_
	);
	LUT2 #(
		.INIT('h8)
	) name2958 (
		_w13462_,
		_w13463_,
		_w13470_
	);
	LUT2 #(
		.INIT('h8)
	) name2959 (
		_w13460_,
		_w13461_,
		_w13471_
	);
	LUT2 #(
		.INIT('h8)
	) name2960 (
		_w13470_,
		_w13471_,
		_w13472_
	);
	LUT2 #(
		.INIT('h8)
	) name2961 (
		_w13468_,
		_w13469_,
		_w13473_
	);
	LUT2 #(
		.INIT('h8)
	) name2962 (
		_w13472_,
		_w13473_,
		_w13474_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		wb_rst_i_pad,
		_w13474_,
		_w13475_
	);
	LUT2 #(
		.INIT('h8)
	) name2964 (
		_w12656_,
		_w13475_,
		_w13476_
	);
	LUT2 #(
		.INIT('h1)
	) name2965 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		\wishbone_TxLength_reg[11]/NET0131 ,
		_w13477_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		\wishbone_TxLength_reg[8]/NET0131 ,
		_w13478_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w13478_,
		_w13479_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w13480_
	);
	LUT2 #(
		.INIT('h4)
	) name2969 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w13480_,
		_w13481_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w13482_
	);
	LUT2 #(
		.INIT('h8)
	) name2971 (
		_w13481_,
		_w13482_,
		_w13483_
	);
	LUT2 #(
		.INIT('h8)
	) name2972 (
		_w13479_,
		_w13483_,
		_w13484_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w13485_
	);
	LUT2 #(
		.INIT('h1)
	) name2974 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w13485_,
		_w13486_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w13485_,
		_w13487_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w13487_,
		_w13488_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w13486_,
		_w13488_,
		_w13489_
	);
	LUT2 #(
		.INIT('h8)
	) name2978 (
		_w13477_,
		_w13484_,
		_w13490_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		_w13489_,
		_w13490_,
		_w13491_
	);
	LUT2 #(
		.INIT('h4)
	) name2980 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w13491_,
		_w13492_
	);
	LUT2 #(
		.INIT('h2)
	) name2981 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		_w13491_,
		_w13493_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		_w13492_,
		_w13493_,
		_w13494_
	);
	LUT2 #(
		.INIT('h1)
	) name2983 (
		\wishbone_TxLength_reg[12]/NET0131 ,
		\wishbone_TxLength_reg[13]/NET0131 ,
		_w13495_
	);
	LUT2 #(
		.INIT('h4)
	) name2984 (
		\wishbone_TxLength_reg[14]/NET0131 ,
		_w13477_,
		_w13496_
	);
	LUT2 #(
		.INIT('h8)
	) name2985 (
		_w13495_,
		_w13496_,
		_w13497_
	);
	LUT2 #(
		.INIT('h4)
	) name2986 (
		\wishbone_TxLength_reg[15]/NET0131 ,
		_w13497_,
		_w13498_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		_w13484_,
		_w13498_,
		_w13499_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		_w12657_,
		_w13499_,
		_w13500_
	);
	LUT2 #(
		.INIT('h4)
	) name2989 (
		_w12656_,
		_w13500_,
		_w13501_
	);
	LUT2 #(
		.INIT('h4)
	) name2990 (
		_w13494_,
		_w13501_,
		_w13502_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		_w12659_,
		_w13502_,
		_w13503_
	);
	LUT2 #(
		.INIT('h4)
	) name2992 (
		_w13476_,
		_w13503_,
		_w13504_
	);
	LUT2 #(
		.INIT('h4)
	) name2993 (
		_w13492_,
		_w13501_,
		_w13505_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		_w12658_,
		_w13505_,
		_w13506_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		\wishbone_TxLength_reg[13]/NET0131 ,
		_w13506_,
		_w13507_
	);
	LUT2 #(
		.INIT('h8)
	) name2996 (
		\wishbone_bd_ram_mem3_reg[175][29]/P0001 ,
		_w13126_,
		_w13508_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		\wishbone_bd_ram_mem3_reg[141][29]/P0001 ,
		_w13004_,
		_w13509_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		\wishbone_bd_ram_mem3_reg[189][29]/P0001 ,
		_w13042_,
		_w13510_
	);
	LUT2 #(
		.INIT('h8)
	) name2999 (
		\wishbone_bd_ram_mem3_reg[185][29]/P0001 ,
		_w12940_,
		_w13511_
	);
	LUT2 #(
		.INIT('h8)
	) name3000 (
		\wishbone_bd_ram_mem3_reg[144][29]/P0001 ,
		_w12756_,
		_w13512_
	);
	LUT2 #(
		.INIT('h8)
	) name3001 (
		\wishbone_bd_ram_mem3_reg[61][29]/P0001 ,
		_w12725_,
		_w13513_
	);
	LUT2 #(
		.INIT('h8)
	) name3002 (
		\wishbone_bd_ram_mem3_reg[135][29]/P0001 ,
		_w13124_,
		_w13514_
	);
	LUT2 #(
		.INIT('h8)
	) name3003 (
		\wishbone_bd_ram_mem3_reg[66][29]/P0001 ,
		_w12824_,
		_w13515_
	);
	LUT2 #(
		.INIT('h8)
	) name3004 (
		\wishbone_bd_ram_mem3_reg[103][29]/P0001 ,
		_w12846_,
		_w13516_
	);
	LUT2 #(
		.INIT('h8)
	) name3005 (
		\wishbone_bd_ram_mem3_reg[240][29]/P0001 ,
		_w12864_,
		_w13517_
	);
	LUT2 #(
		.INIT('h8)
	) name3006 (
		\wishbone_bd_ram_mem3_reg[170][29]/P0001 ,
		_w13030_,
		_w13518_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		\wishbone_bd_ram_mem3_reg[136][29]/P0001 ,
		_w13064_,
		_w13519_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\wishbone_bd_ram_mem3_reg[13][29]/P0001 ,
		_w13178_,
		_w13520_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\wishbone_bd_ram_mem3_reg[162][29]/P0001 ,
		_w13098_,
		_w13521_
	);
	LUT2 #(
		.INIT('h8)
	) name3010 (
		\wishbone_bd_ram_mem3_reg[131][29]/P0001 ,
		_w12852_,
		_w13522_
	);
	LUT2 #(
		.INIT('h8)
	) name3011 (
		\wishbone_bd_ram_mem3_reg[22][29]/P0001 ,
		_w13110_,
		_w13523_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		\wishbone_bd_ram_mem3_reg[247][29]/P0001 ,
		_w12818_,
		_w13524_
	);
	LUT2 #(
		.INIT('h8)
	) name3013 (
		\wishbone_bd_ram_mem3_reg[222][29]/P0001 ,
		_w13094_,
		_w13525_
	);
	LUT2 #(
		.INIT('h8)
	) name3014 (
		\wishbone_bd_ram_mem3_reg[34][29]/P0001 ,
		_w12930_,
		_w13526_
	);
	LUT2 #(
		.INIT('h8)
	) name3015 (
		\wishbone_bd_ram_mem3_reg[17][29]/P0001 ,
		_w12848_,
		_w13527_
	);
	LUT2 #(
		.INIT('h8)
	) name3016 (
		\wishbone_bd_ram_mem3_reg[80][29]/P0001 ,
		_w12689_,
		_w13528_
	);
	LUT2 #(
		.INIT('h8)
	) name3017 (
		\wishbone_bd_ram_mem3_reg[91][29]/P0001 ,
		_w13074_,
		_w13529_
	);
	LUT2 #(
		.INIT('h8)
	) name3018 (
		\wishbone_bd_ram_mem3_reg[212][29]/P0001 ,
		_w12796_,
		_w13530_
	);
	LUT2 #(
		.INIT('h8)
	) name3019 (
		\wishbone_bd_ram_mem3_reg[107][29]/P0001 ,
		_w12749_,
		_w13531_
	);
	LUT2 #(
		.INIT('h8)
	) name3020 (
		\wishbone_bd_ram_mem3_reg[169][29]/P0001 ,
		_w12722_,
		_w13532_
	);
	LUT2 #(
		.INIT('h8)
	) name3021 (
		\wishbone_bd_ram_mem3_reg[149][29]/P0001 ,
		_w12741_,
		_w13533_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		\wishbone_bd_ram_mem3_reg[182][29]/P0001 ,
		_w12820_,
		_w13534_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		\wishbone_bd_ram_mem3_reg[154][29]/P0001 ,
		_w12962_,
		_w13535_
	);
	LUT2 #(
		.INIT('h8)
	) name3024 (
		\wishbone_bd_ram_mem3_reg[139][29]/P0001 ,
		_w12814_,
		_w13536_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		\wishbone_bd_ram_mem3_reg[142][29]/P0001 ,
		_w12928_,
		_w13537_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		\wishbone_bd_ram_mem3_reg[198][29]/P0001 ,
		_w12832_,
		_w13538_
	);
	LUT2 #(
		.INIT('h8)
	) name3027 (
		\wishbone_bd_ram_mem3_reg[244][29]/P0001 ,
		_w12747_,
		_w13539_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		\wishbone_bd_ram_mem3_reg[101][29]/P0001 ,
		_w13192_,
		_w13540_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		\wishbone_bd_ram_mem3_reg[226][29]/P0001 ,
		_w13138_,
		_w13541_
	);
	LUT2 #(
		.INIT('h8)
	) name3030 (
		\wishbone_bd_ram_mem3_reg[159][29]/P0001 ,
		_w12774_,
		_w13542_
	);
	LUT2 #(
		.INIT('h8)
	) name3031 (
		\wishbone_bd_ram_mem3_reg[116][29]/P0001 ,
		_w12998_,
		_w13543_
	);
	LUT2 #(
		.INIT('h8)
	) name3032 (
		\wishbone_bd_ram_mem3_reg[38][29]/P0001 ,
		_w13182_,
		_w13544_
	);
	LUT2 #(
		.INIT('h8)
	) name3033 (
		\wishbone_bd_ram_mem3_reg[45][29]/P0001 ,
		_w12908_,
		_w13545_
	);
	LUT2 #(
		.INIT('h8)
	) name3034 (
		\wishbone_bd_ram_mem3_reg[195][29]/P0001 ,
		_w13144_,
		_w13546_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		\wishbone_bd_ram_mem3_reg[196][29]/P0001 ,
		_w13090_,
		_w13547_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		\wishbone_bd_ram_mem3_reg[183][29]/P0001 ,
		_w12787_,
		_w13548_
	);
	LUT2 #(
		.INIT('h8)
	) name3037 (
		\wishbone_bd_ram_mem3_reg[252][29]/P0001 ,
		_w13080_,
		_w13549_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		\wishbone_bd_ram_mem3_reg[180][29]/P0001 ,
		_w12791_,
		_w13550_
	);
	LUT2 #(
		.INIT('h8)
	) name3039 (
		\wishbone_bd_ram_mem3_reg[29][29]/P0001 ,
		_w12952_,
		_w13551_
	);
	LUT2 #(
		.INIT('h8)
	) name3040 (
		\wishbone_bd_ram_mem3_reg[203][29]/P0001 ,
		_w13158_,
		_w13552_
	);
	LUT2 #(
		.INIT('h8)
	) name3041 (
		\wishbone_bd_ram_mem3_reg[117][29]/P0001 ,
		_w12715_,
		_w13553_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		\wishbone_bd_ram_mem3_reg[73][29]/P0001 ,
		_w12918_,
		_w13554_
	);
	LUT2 #(
		.INIT('h8)
	) name3043 (
		\wishbone_bd_ram_mem3_reg[251][29]/P0001 ,
		_w13054_,
		_w13555_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		\wishbone_bd_ram_mem3_reg[220][29]/P0001 ,
		_w13066_,
		_w13556_
	);
	LUT2 #(
		.INIT('h8)
	) name3045 (
		\wishbone_bd_ram_mem3_reg[216][29]/P0001 ,
		_w13028_,
		_w13557_
	);
	LUT2 #(
		.INIT('h8)
	) name3046 (
		\wishbone_bd_ram_mem3_reg[12][29]/P0001 ,
		_w13118_,
		_w13558_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		\wishbone_bd_ram_mem3_reg[56][29]/P0001 ,
		_w12778_,
		_w13559_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		\wishbone_bd_ram_mem3_reg[6][29]/P0001 ,
		_w12968_,
		_w13560_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		\wishbone_bd_ram_mem3_reg[110][29]/P0001 ,
		_w13046_,
		_w13561_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		\wishbone_bd_ram_mem3_reg[89][29]/P0001 ,
		_w12964_,
		_w13562_
	);
	LUT2 #(
		.INIT('h8)
	) name3051 (
		\wishbone_bd_ram_mem3_reg[64][29]/P0001 ,
		_w12976_,
		_w13563_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		\wishbone_bd_ram_mem3_reg[171][29]/P0001 ,
		_w12910_,
		_w13564_
	);
	LUT2 #(
		.INIT('h8)
	) name3053 (
		\wishbone_bd_ram_mem3_reg[239][29]/P0001 ,
		_w12862_,
		_w13565_
	);
	LUT2 #(
		.INIT('h8)
	) name3054 (
		\wishbone_bd_ram_mem3_reg[93][29]/P0001 ,
		_w13016_,
		_w13566_
	);
	LUT2 #(
		.INIT('h8)
	) name3055 (
		\wishbone_bd_ram_mem3_reg[59][29]/P0001 ,
		_w12780_,
		_w13567_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		\wishbone_bd_ram_mem3_reg[194][29]/P0001 ,
		_w12772_,
		_w13568_
	);
	LUT2 #(
		.INIT('h8)
	) name3057 (
		\wishbone_bd_ram_mem3_reg[39][29]/P0001 ,
		_w13018_,
		_w13569_
	);
	LUT2 #(
		.INIT('h8)
	) name3058 (
		\wishbone_bd_ram_mem3_reg[237][29]/P0001 ,
		_w12990_,
		_w13570_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		\wishbone_bd_ram_mem3_reg[204][29]/P0001 ,
		_w13162_,
		_w13571_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		\wishbone_bd_ram_mem3_reg[233][29]/P0001 ,
		_w12836_,
		_w13572_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		\wishbone_bd_ram_mem3_reg[191][29]/P0001 ,
		_w13034_,
		_w13573_
	);
	LUT2 #(
		.INIT('h8)
	) name3062 (
		\wishbone_bd_ram_mem3_reg[83][29]/P0001 ,
		_w12916_,
		_w13574_
	);
	LUT2 #(
		.INIT('h8)
	) name3063 (
		\wishbone_bd_ram_mem3_reg[27][29]/P0001 ,
		_w12880_,
		_w13575_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		\wishbone_bd_ram_mem3_reg[125][29]/P0001 ,
		_w12956_,
		_w13576_
	);
	LUT2 #(
		.INIT('h8)
	) name3065 (
		\wishbone_bd_ram_mem3_reg[121][29]/P0001 ,
		_w13078_,
		_w13577_
	);
	LUT2 #(
		.INIT('h8)
	) name3066 (
		\wishbone_bd_ram_mem3_reg[4][29]/P0001 ,
		_w12666_,
		_w13578_
	);
	LUT2 #(
		.INIT('h8)
	) name3067 (
		\wishbone_bd_ram_mem3_reg[81][29]/P0001 ,
		_w12950_,
		_w13579_
	);
	LUT2 #(
		.INIT('h8)
	) name3068 (
		\wishbone_bd_ram_mem3_reg[67][29]/P0001 ,
		_w13134_,
		_w13580_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		\wishbone_bd_ram_mem3_reg[106][29]/P0001 ,
		_w12713_,
		_w13581_
	);
	LUT2 #(
		.INIT('h8)
	) name3070 (
		\wishbone_bd_ram_mem3_reg[174][29]/P0001 ,
		_w12972_,
		_w13582_
	);
	LUT2 #(
		.INIT('h8)
	) name3071 (
		\wishbone_bd_ram_mem3_reg[181][29]/P0001 ,
		_w12828_,
		_w13583_
	);
	LUT2 #(
		.INIT('h8)
	) name3072 (
		\wishbone_bd_ram_mem3_reg[104][29]/P0001 ,
		_w13148_,
		_w13584_
	);
	LUT2 #(
		.INIT('h8)
	) name3073 (
		\wishbone_bd_ram_mem3_reg[201][29]/P0001 ,
		_w12822_,
		_w13585_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		\wishbone_bd_ram_mem3_reg[75][29]/P0001 ,
		_w12826_,
		_w13586_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		\wishbone_bd_ram_mem3_reg[2][29]/P0001 ,
		_w13088_,
		_w13587_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		\wishbone_bd_ram_mem3_reg[202][29]/P0001 ,
		_w12870_,
		_w13588_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		\wishbone_bd_ram_mem3_reg[111][29]/P0001 ,
		_w12744_,
		_w13589_
	);
	LUT2 #(
		.INIT('h8)
	) name3078 (
		\wishbone_bd_ram_mem3_reg[160][29]/P0001 ,
		_w12872_,
		_w13590_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		\wishbone_bd_ram_mem3_reg[127][29]/P0001 ,
		_w13164_,
		_w13591_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		\wishbone_bd_ram_mem3_reg[77][29]/P0001 ,
		_w12982_,
		_w13592_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		\wishbone_bd_ram_mem3_reg[42][29]/P0001 ,
		_w12842_,
		_w13593_
	);
	LUT2 #(
		.INIT('h8)
	) name3082 (
		\wishbone_bd_ram_mem3_reg[65][29]/P0001 ,
		_w13176_,
		_w13594_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		\wishbone_bd_ram_mem3_reg[70][29]/P0001 ,
		_w12840_,
		_w13595_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		\wishbone_bd_ram_mem3_reg[46][29]/P0001 ,
		_w12884_,
		_w13596_
	);
	LUT2 #(
		.INIT('h8)
	) name3085 (
		\wishbone_bd_ram_mem3_reg[112][29]/P0001 ,
		_w12733_,
		_w13597_
	);
	LUT2 #(
		.INIT('h8)
	) name3086 (
		\wishbone_bd_ram_mem3_reg[36][29]/P0001 ,
		_w12800_,
		_w13598_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		\wishbone_bd_ram_mem3_reg[90][29]/P0001 ,
		_w12978_,
		_w13599_
	);
	LUT2 #(
		.INIT('h8)
	) name3088 (
		\wishbone_bd_ram_mem3_reg[71][29]/P0001 ,
		_w12798_,
		_w13600_
	);
	LUT2 #(
		.INIT('h8)
	) name3089 (
		\wishbone_bd_ram_mem3_reg[113][29]/P0001 ,
		_w13026_,
		_w13601_
	);
	LUT2 #(
		.INIT('h8)
	) name3090 (
		\wishbone_bd_ram_mem3_reg[86][29]/P0001 ,
		_w12735_,
		_w13602_
	);
	LUT2 #(
		.INIT('h8)
	) name3091 (
		\wishbone_bd_ram_mem3_reg[158][29]/P0001 ,
		_w12898_,
		_w13603_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		\wishbone_bd_ram_mem3_reg[253][29]/P0001 ,
		_w13100_,
		_w13604_
	);
	LUT2 #(
		.INIT('h8)
	) name3093 (
		\wishbone_bd_ram_mem3_reg[243][29]/P0001 ,
		_w12804_,
		_w13605_
	);
	LUT2 #(
		.INIT('h8)
	) name3094 (
		\wishbone_bd_ram_mem3_reg[57][29]/P0001 ,
		_w13116_,
		_w13606_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		\wishbone_bd_ram_mem3_reg[44][29]/P0001 ,
		_w12896_,
		_w13607_
	);
	LUT2 #(
		.INIT('h8)
	) name3096 (
		\wishbone_bd_ram_mem3_reg[123][29]/P0001 ,
		_w13114_,
		_w13608_
	);
	LUT2 #(
		.INIT('h8)
	) name3097 (
		\wishbone_bd_ram_mem3_reg[192][29]/P0001 ,
		_w12938_,
		_w13609_
	);
	LUT2 #(
		.INIT('h8)
	) name3098 (
		\wishbone_bd_ram_mem3_reg[173][29]/P0001 ,
		_w12854_,
		_w13610_
	);
	LUT2 #(
		.INIT('h8)
	) name3099 (
		\wishbone_bd_ram_mem3_reg[120][29]/P0001 ,
		_w12707_,
		_w13611_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		\wishbone_bd_ram_mem3_reg[48][29]/P0001 ,
		_w12970_,
		_w13612_
	);
	LUT2 #(
		.INIT('h8)
	) name3101 (
		\wishbone_bd_ram_mem3_reg[35][29]/P0001 ,
		_w12703_,
		_w13613_
	);
	LUT2 #(
		.INIT('h8)
	) name3102 (
		\wishbone_bd_ram_mem3_reg[24][29]/P0001 ,
		_w13084_,
		_w13614_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		\wishbone_bd_ram_mem3_reg[231][29]/P0001 ,
		_w12856_,
		_w13615_
	);
	LUT2 #(
		.INIT('h8)
	) name3104 (
		\wishbone_bd_ram_mem3_reg[210][29]/P0001 ,
		_w12924_,
		_w13616_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		\wishbone_bd_ram_mem3_reg[85][29]/P0001 ,
		_w13216_,
		_w13617_
	);
	LUT2 #(
		.INIT('h8)
	) name3106 (
		\wishbone_bd_ram_mem3_reg[134][29]/P0001 ,
		_w12763_,
		_w13618_
	);
	LUT2 #(
		.INIT('h8)
	) name3107 (
		\wishbone_bd_ram_mem3_reg[95][29]/P0001 ,
		_w12844_,
		_w13619_
	);
	LUT2 #(
		.INIT('h8)
	) name3108 (
		\wishbone_bd_ram_mem3_reg[199][29]/P0001 ,
		_w12768_,
		_w13620_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		\wishbone_bd_ram_mem3_reg[49][29]/P0001 ,
		_w12994_,
		_w13621_
	);
	LUT2 #(
		.INIT('h8)
	) name3110 (
		\wishbone_bd_ram_mem3_reg[250][29]/P0001 ,
		_w13128_,
		_w13622_
	);
	LUT2 #(
		.INIT('h8)
	) name3111 (
		\wishbone_bd_ram_mem3_reg[126][29]/P0001 ,
		_w13218_,
		_w13623_
	);
	LUT2 #(
		.INIT('h8)
	) name3112 (
		\wishbone_bd_ram_mem3_reg[224][29]/P0001 ,
		_w12902_,
		_w13624_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		\wishbone_bd_ram_mem3_reg[188][29]/P0001 ,
		_w12948_,
		_w13625_
	);
	LUT2 #(
		.INIT('h8)
	) name3114 (
		\wishbone_bd_ram_mem3_reg[105][29]/P0001 ,
		_w12751_,
		_w13626_
	);
	LUT2 #(
		.INIT('h8)
	) name3115 (
		\wishbone_bd_ram_mem3_reg[58][29]/P0001 ,
		_w13070_,
		_w13627_
	);
	LUT2 #(
		.INIT('h8)
	) name3116 (
		\wishbone_bd_ram_mem3_reg[193][29]/P0001 ,
		_w13056_,
		_w13628_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		\wishbone_bd_ram_mem3_reg[178][29]/P0001 ,
		_w12886_,
		_w13629_
	);
	LUT2 #(
		.INIT('h8)
	) name3118 (
		\wishbone_bd_ram_mem3_reg[47][29]/P0001 ,
		_w12904_,
		_w13630_
	);
	LUT2 #(
		.INIT('h8)
	) name3119 (
		\wishbone_bd_ram_mem3_reg[225][29]/P0001 ,
		_w13092_,
		_w13631_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		\wishbone_bd_ram_mem3_reg[143][29]/P0001 ,
		_w12922_,
		_w13632_
	);
	LUT2 #(
		.INIT('h8)
	) name3121 (
		\wishbone_bd_ram_mem3_reg[147][29]/P0001 ,
		_w13146_,
		_w13633_
	);
	LUT2 #(
		.INIT('h8)
	) name3122 (
		\wishbone_bd_ram_mem3_reg[100][29]/P0001 ,
		_w12960_,
		_w13634_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		\wishbone_bd_ram_mem3_reg[94][29]/P0001 ,
		_w13186_,
		_w13635_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		\wishbone_bd_ram_mem3_reg[102][29]/P0001 ,
		_w12685_,
		_w13636_
	);
	LUT2 #(
		.INIT('h8)
	) name3125 (
		\wishbone_bd_ram_mem3_reg[129][29]/P0001 ,
		_w12776_,
		_w13637_
	);
	LUT2 #(
		.INIT('h8)
	) name3126 (
		\wishbone_bd_ram_mem3_reg[10][29]/P0001 ,
		_w13172_,
		_w13638_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		\wishbone_bd_ram_mem3_reg[163][29]/P0001 ,
		_w12882_,
		_w13639_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		\wishbone_bd_ram_mem3_reg[151][29]/P0001 ,
		_w13142_,
		_w13640_
	);
	LUT2 #(
		.INIT('h8)
	) name3129 (
		\wishbone_bd_ram_mem3_reg[14][29]/P0001 ,
		_w13086_,
		_w13641_
	);
	LUT2 #(
		.INIT('h8)
	) name3130 (
		\wishbone_bd_ram_mem3_reg[26][29]/P0001 ,
		_w12699_,
		_w13642_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		\wishbone_bd_ram_mem3_reg[200][29]/P0001 ,
		_w12988_,
		_w13643_
	);
	LUT2 #(
		.INIT('h8)
	) name3132 (
		\wishbone_bd_ram_mem3_reg[18][29]/P0001 ,
		_w12679_,
		_w13644_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		\wishbone_bd_ram_mem3_reg[88][29]/P0001 ,
		_w12860_,
		_w13645_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		\wishbone_bd_ram_mem3_reg[219][29]/P0001 ,
		_w12806_,
		_w13646_
	);
	LUT2 #(
		.INIT('h8)
	) name3135 (
		\wishbone_bd_ram_mem3_reg[167][29]/P0001 ,
		_w12986_,
		_w13647_
	);
	LUT2 #(
		.INIT('h8)
	) name3136 (
		\wishbone_bd_ram_mem3_reg[205][29]/P0001 ,
		_w13068_,
		_w13648_
	);
	LUT2 #(
		.INIT('h8)
	) name3137 (
		\wishbone_bd_ram_mem3_reg[176][29]/P0001 ,
		_w12868_,
		_w13649_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		\wishbone_bd_ram_mem3_reg[23][29]/P0001 ,
		_w13008_,
		_w13650_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		\wishbone_bd_ram_mem3_reg[164][29]/P0001 ,
		_w12876_,
		_w13651_
	);
	LUT2 #(
		.INIT('h8)
	) name3140 (
		\wishbone_bd_ram_mem3_reg[146][29]/P0001 ,
		_w13060_,
		_w13652_
	);
	LUT2 #(
		.INIT('h8)
	) name3141 (
		\wishbone_bd_ram_mem3_reg[54][29]/P0001 ,
		_w12770_,
		_w13653_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		\wishbone_bd_ram_mem3_reg[128][29]/P0001 ,
		_w12793_,
		_w13654_
	);
	LUT2 #(
		.INIT('h8)
	) name3143 (
		\wishbone_bd_ram_mem3_reg[229][29]/P0001 ,
		_w12711_,
		_w13655_
	);
	LUT2 #(
		.INIT('h8)
	) name3144 (
		\wishbone_bd_ram_mem3_reg[62][29]/P0001 ,
		_w12673_,
		_w13656_
	);
	LUT2 #(
		.INIT('h8)
	) name3145 (
		\wishbone_bd_ram_mem3_reg[248][29]/P0001 ,
		_w12789_,
		_w13657_
	);
	LUT2 #(
		.INIT('h8)
	) name3146 (
		\wishbone_bd_ram_mem3_reg[152][29]/P0001 ,
		_w12966_,
		_w13658_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		\wishbone_bd_ram_mem3_reg[172][29]/P0001 ,
		_w12944_,
		_w13659_
	);
	LUT2 #(
		.INIT('h8)
	) name3148 (
		\wishbone_bd_ram_mem3_reg[28][29]/P0001 ,
		_w13170_,
		_w13660_
	);
	LUT2 #(
		.INIT('h8)
	) name3149 (
		\wishbone_bd_ram_mem3_reg[3][29]/P0001 ,
		_w12866_,
		_w13661_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		\wishbone_bd_ram_mem3_reg[137][29]/P0001 ,
		_w13168_,
		_w13662_
	);
	LUT2 #(
		.INIT('h8)
	) name3151 (
		\wishbone_bd_ram_mem3_reg[78][29]/P0001 ,
		_w12874_,
		_w13663_
	);
	LUT2 #(
		.INIT('h8)
	) name3152 (
		\wishbone_bd_ram_mem3_reg[165][29]/P0001 ,
		_w13044_,
		_w13664_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		\wishbone_bd_ram_mem3_reg[254][29]/P0001 ,
		_w12892_,
		_w13665_
	);
	LUT2 #(
		.INIT('h8)
	) name3154 (
		\wishbone_bd_ram_mem3_reg[76][29]/P0001 ,
		_w13184_,
		_w13666_
	);
	LUT2 #(
		.INIT('h8)
	) name3155 (
		\wishbone_bd_ram_mem3_reg[179][29]/P0001 ,
		_w13050_,
		_w13667_
	);
	LUT2 #(
		.INIT('h8)
	) name3156 (
		\wishbone_bd_ram_mem3_reg[217][29]/P0001 ,
		_w13188_,
		_w13668_
	);
	LUT2 #(
		.INIT('h8)
	) name3157 (
		\wishbone_bd_ram_mem3_reg[209][29]/P0001 ,
		_w13152_,
		_w13669_
	);
	LUT2 #(
		.INIT('h8)
	) name3158 (
		\wishbone_bd_ram_mem3_reg[150][29]/P0001 ,
		_w13136_,
		_w13670_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		\wishbone_bd_ram_mem3_reg[223][29]/P0001 ,
		_w12838_,
		_w13671_
	);
	LUT2 #(
		.INIT('h8)
	) name3160 (
		\wishbone_bd_ram_mem3_reg[153][29]/P0001 ,
		_w12890_,
		_w13672_
	);
	LUT2 #(
		.INIT('h8)
	) name3161 (
		\wishbone_bd_ram_mem3_reg[155][29]/P0001 ,
		_w13122_,
		_w13673_
	);
	LUT2 #(
		.INIT('h8)
	) name3162 (
		\wishbone_bd_ram_mem3_reg[96][29]/P0001 ,
		_w12912_,
		_w13674_
	);
	LUT2 #(
		.INIT('h8)
	) name3163 (
		\wishbone_bd_ram_mem3_reg[156][29]/P0001 ,
		_w13190_,
		_w13675_
	);
	LUT2 #(
		.INIT('h8)
	) name3164 (
		\wishbone_bd_ram_mem3_reg[92][29]/P0001 ,
		_w13010_,
		_w13676_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		\wishbone_bd_ram_mem3_reg[132][29]/P0001 ,
		_w12992_,
		_w13677_
	);
	LUT2 #(
		.INIT('h8)
	) name3166 (
		\wishbone_bd_ram_mem3_reg[37][29]/P0001 ,
		_w13102_,
		_w13678_
	);
	LUT2 #(
		.INIT('h8)
	) name3167 (
		\wishbone_bd_ram_mem3_reg[197][29]/P0001 ,
		_w12834_,
		_w13679_
	);
	LUT2 #(
		.INIT('h8)
	) name3168 (
		\wishbone_bd_ram_mem3_reg[55][29]/P0001 ,
		_w12785_,
		_w13680_
	);
	LUT2 #(
		.INIT('h8)
	) name3169 (
		\wishbone_bd_ram_mem3_reg[99][29]/P0001 ,
		_w13038_,
		_w13681_
	);
	LUT2 #(
		.INIT('h8)
	) name3170 (
		\wishbone_bd_ram_mem3_reg[234][29]/P0001 ,
		_w13214_,
		_w13682_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		\wishbone_bd_ram_mem3_reg[187][29]/P0001 ,
		_w13196_,
		_w13683_
	);
	LUT2 #(
		.INIT('h8)
	) name3172 (
		\wishbone_bd_ram_mem3_reg[177][29]/P0001 ,
		_w12996_,
		_w13684_
	);
	LUT2 #(
		.INIT('h8)
	) name3173 (
		\wishbone_bd_ram_mem3_reg[133][29]/P0001 ,
		_w12761_,
		_w13685_
	);
	LUT2 #(
		.INIT('h8)
	) name3174 (
		\wishbone_bd_ram_mem3_reg[218][29]/P0001 ,
		_w13206_,
		_w13686_
	);
	LUT2 #(
		.INIT('h8)
	) name3175 (
		\wishbone_bd_ram_mem3_reg[235][29]/P0001 ,
		_w12696_,
		_w13687_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		\wishbone_bd_ram_mem3_reg[236][29]/P0001 ,
		_w12731_,
		_w13688_
	);
	LUT2 #(
		.INIT('h8)
	) name3177 (
		\wishbone_bd_ram_mem3_reg[79][29]/P0001 ,
		_w13212_,
		_w13689_
	);
	LUT2 #(
		.INIT('h8)
	) name3178 (
		\wishbone_bd_ram_mem3_reg[140][29]/P0001 ,
		_w12894_,
		_w13690_
	);
	LUT2 #(
		.INIT('h8)
	) name3179 (
		\wishbone_bd_ram_mem3_reg[124][29]/P0001 ,
		_w13058_,
		_w13691_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		\wishbone_bd_ram_mem3_reg[245][29]/P0001 ,
		_w13022_,
		_w13692_
	);
	LUT2 #(
		.INIT('h8)
	) name3181 (
		\wishbone_bd_ram_mem3_reg[16][29]/P0001 ,
		_w13140_,
		_w13693_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		\wishbone_bd_ram_mem3_reg[227][29]/P0001 ,
		_w12936_,
		_w13694_
	);
	LUT2 #(
		.INIT('h8)
	) name3183 (
		\wishbone_bd_ram_mem3_reg[52][29]/P0001 ,
		_w13082_,
		_w13695_
	);
	LUT2 #(
		.INIT('h8)
	) name3184 (
		\wishbone_bd_ram_mem3_reg[5][29]/P0001 ,
		_w12878_,
		_w13696_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		\wishbone_bd_ram_mem3_reg[31][29]/P0001 ,
		_w13198_,
		_w13697_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		\wishbone_bd_ram_mem3_reg[30][29]/P0001 ,
		_w13104_,
		_w13698_
	);
	LUT2 #(
		.INIT('h8)
	) name3187 (
		\wishbone_bd_ram_mem3_reg[184][29]/P0001 ,
		_w13062_,
		_w13699_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		\wishbone_bd_ram_mem3_reg[190][29]/P0001 ,
		_w12858_,
		_w13700_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		\wishbone_bd_ram_mem3_reg[232][29]/P0001 ,
		_w12758_,
		_w13701_
	);
	LUT2 #(
		.INIT('h8)
	) name3190 (
		\wishbone_bd_ram_mem3_reg[228][29]/P0001 ,
		_w12765_,
		_w13702_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		\wishbone_bd_ram_mem3_reg[214][29]/P0001 ,
		_w12984_,
		_w13703_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		\wishbone_bd_ram_mem3_reg[221][29]/P0001 ,
		_w12802_,
		_w13704_
	);
	LUT2 #(
		.INIT('h8)
	) name3193 (
		\wishbone_bd_ram_mem3_reg[0][29]/P0001 ,
		_w12717_,
		_w13705_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		\wishbone_bd_ram_mem3_reg[50][29]/P0001 ,
		_w13150_,
		_w13706_
	);
	LUT2 #(
		.INIT('h8)
	) name3195 (
		\wishbone_bd_ram_mem3_reg[230][29]/P0001 ,
		_w13036_,
		_w13707_
	);
	LUT2 #(
		.INIT('h8)
	) name3196 (
		\wishbone_bd_ram_mem3_reg[32][29]/P0001 ,
		_w13120_,
		_w13708_
	);
	LUT2 #(
		.INIT('h8)
	) name3197 (
		\wishbone_bd_ram_mem3_reg[41][29]/P0001 ,
		_w13052_,
		_w13709_
	);
	LUT2 #(
		.INIT('h8)
	) name3198 (
		\wishbone_bd_ram_mem3_reg[51][29]/P0001 ,
		_w13024_,
		_w13710_
	);
	LUT2 #(
		.INIT('h8)
	) name3199 (
		\wishbone_bd_ram_mem3_reg[208][29]/P0001 ,
		_w13032_,
		_w13711_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		\wishbone_bd_ram_mem3_reg[119][29]/P0001 ,
		_w13048_,
		_w13712_
	);
	LUT2 #(
		.INIT('h8)
	) name3201 (
		\wishbone_bd_ram_mem3_reg[9][29]/P0001 ,
		_w12808_,
		_w13713_
	);
	LUT2 #(
		.INIT('h8)
	) name3202 (
		\wishbone_bd_ram_mem3_reg[215][29]/P0001 ,
		_w12974_,
		_w13714_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		\wishbone_bd_ram_mem3_reg[74][29]/P0001 ,
		_w12812_,
		_w13715_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		\wishbone_bd_ram_mem3_reg[157][29]/P0001 ,
		_w12926_,
		_w13716_
	);
	LUT2 #(
		.INIT('h8)
	) name3205 (
		\wishbone_bd_ram_mem3_reg[8][29]/P0001 ,
		_w12920_,
		_w13717_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		\wishbone_bd_ram_mem3_reg[213][29]/P0001 ,
		_w13002_,
		_w13718_
	);
	LUT2 #(
		.INIT('h8)
	) name3207 (
		\wishbone_bd_ram_mem3_reg[63][29]/P0001 ,
		_w12850_,
		_w13719_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		\wishbone_bd_ram_mem3_reg[40][29]/P0001 ,
		_w13132_,
		_w13720_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		\wishbone_bd_ram_mem3_reg[1][29]/P0001 ,
		_w13014_,
		_w13721_
	);
	LUT2 #(
		.INIT('h8)
	) name3210 (
		\wishbone_bd_ram_mem3_reg[82][29]/P0001 ,
		_w12942_,
		_w13722_
	);
	LUT2 #(
		.INIT('h8)
	) name3211 (
		\wishbone_bd_ram_mem3_reg[206][29]/P0001 ,
		_w12954_,
		_w13723_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		\wishbone_bd_ram_mem3_reg[148][29]/P0001 ,
		_w13000_,
		_w13724_
	);
	LUT2 #(
		.INIT('h8)
	) name3213 (
		\wishbone_bd_ram_mem3_reg[98][29]/P0001 ,
		_w12816_,
		_w13725_
	);
	LUT2 #(
		.INIT('h8)
	) name3214 (
		\wishbone_bd_ram_mem3_reg[186][29]/P0001 ,
		_w12783_,
		_w13726_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		\wishbone_bd_ram_mem3_reg[7][29]/P0001 ,
		_w12728_,
		_w13727_
	);
	LUT2 #(
		.INIT('h8)
	) name3216 (
		\wishbone_bd_ram_mem3_reg[166][29]/P0001 ,
		_w13040_,
		_w13728_
	);
	LUT2 #(
		.INIT('h8)
	) name3217 (
		\wishbone_bd_ram_mem3_reg[69][29]/P0001 ,
		_w12738_,
		_w13729_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		\wishbone_bd_ram_mem3_reg[84][29]/P0001 ,
		_w12934_,
		_w13730_
	);
	LUT2 #(
		.INIT('h8)
	) name3219 (
		\wishbone_bd_ram_mem3_reg[53][29]/P0001 ,
		_w13020_,
		_w13731_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		\wishbone_bd_ram_mem3_reg[145][29]/P0001 ,
		_w13106_,
		_w13732_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		\wishbone_bd_ram_mem3_reg[114][29]/P0001 ,
		_w13202_,
		_w13733_
	);
	LUT2 #(
		.INIT('h8)
	) name3222 (
		\wishbone_bd_ram_mem3_reg[246][29]/P0001 ,
		_w13076_,
		_w13734_
	);
	LUT2 #(
		.INIT('h8)
	) name3223 (
		\wishbone_bd_ram_mem3_reg[255][29]/P0001 ,
		_w13072_,
		_w13735_
	);
	LUT2 #(
		.INIT('h8)
	) name3224 (
		\wishbone_bd_ram_mem3_reg[108][29]/P0001 ,
		_w13156_,
		_w13736_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		\wishbone_bd_ram_mem3_reg[211][29]/P0001 ,
		_w13166_,
		_w13737_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		\wishbone_bd_ram_mem3_reg[97][29]/P0001 ,
		_w13096_,
		_w13738_
	);
	LUT2 #(
		.INIT('h8)
	) name3227 (
		\wishbone_bd_ram_mem3_reg[19][29]/P0001 ,
		_w13012_,
		_w13739_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		\wishbone_bd_ram_mem3_reg[11][29]/P0001 ,
		_w13194_,
		_w13740_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		\wishbone_bd_ram_mem3_reg[161][29]/P0001 ,
		_w12754_,
		_w13741_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\wishbone_bd_ram_mem3_reg[21][29]/P0001 ,
		_w12906_,
		_w13742_
	);
	LUT2 #(
		.INIT('h8)
	) name3231 (
		\wishbone_bd_ram_mem3_reg[33][29]/P0001 ,
		_w12980_,
		_w13743_
	);
	LUT2 #(
		.INIT('h8)
	) name3232 (
		\wishbone_bd_ram_mem3_reg[207][29]/P0001 ,
		_w13180_,
		_w13744_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		\wishbone_bd_ram_mem3_reg[20][29]/P0001 ,
		_w13174_,
		_w13745_
	);
	LUT2 #(
		.INIT('h8)
	) name3234 (
		\wishbone_bd_ram_mem3_reg[25][29]/P0001 ,
		_w13108_,
		_w13746_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		\wishbone_bd_ram_mem3_reg[238][29]/P0001 ,
		_w13160_,
		_w13747_
	);
	LUT2 #(
		.INIT('h8)
	) name3236 (
		\wishbone_bd_ram_mem3_reg[87][29]/P0001 ,
		_w13154_,
		_w13748_
	);
	LUT2 #(
		.INIT('h8)
	) name3237 (
		\wishbone_bd_ram_mem3_reg[130][29]/P0001 ,
		_w12914_,
		_w13749_
	);
	LUT2 #(
		.INIT('h8)
	) name3238 (
		\wishbone_bd_ram_mem3_reg[138][29]/P0001 ,
		_w12958_,
		_w13750_
	);
	LUT2 #(
		.INIT('h8)
	) name3239 (
		\wishbone_bd_ram_mem3_reg[115][29]/P0001 ,
		_w13112_,
		_w13751_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		\wishbone_bd_ram_mem3_reg[249][29]/P0001 ,
		_w12900_,
		_w13752_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		\wishbone_bd_ram_mem3_reg[15][29]/P0001 ,
		_w13210_,
		_w13753_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		\wishbone_bd_ram_mem3_reg[68][29]/P0001 ,
		_w12946_,
		_w13754_
	);
	LUT2 #(
		.INIT('h8)
	) name3243 (
		\wishbone_bd_ram_mem3_reg[72][29]/P0001 ,
		_w12810_,
		_w13755_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		\wishbone_bd_ram_mem3_reg[60][29]/P0001 ,
		_w13204_,
		_w13756_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		\wishbone_bd_ram_mem3_reg[168][29]/P0001 ,
		_w13208_,
		_w13757_
	);
	LUT2 #(
		.INIT('h8)
	) name3246 (
		\wishbone_bd_ram_mem3_reg[122][29]/P0001 ,
		_w13130_,
		_w13758_
	);
	LUT2 #(
		.INIT('h8)
	) name3247 (
		\wishbone_bd_ram_mem3_reg[109][29]/P0001 ,
		_w12888_,
		_w13759_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		\wishbone_bd_ram_mem3_reg[43][29]/P0001 ,
		_w13200_,
		_w13760_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		\wishbone_bd_ram_mem3_reg[241][29]/P0001 ,
		_w13006_,
		_w13761_
	);
	LUT2 #(
		.INIT('h8)
	) name3250 (
		\wishbone_bd_ram_mem3_reg[118][29]/P0001 ,
		_w12830_,
		_w13762_
	);
	LUT2 #(
		.INIT('h8)
	) name3251 (
		\wishbone_bd_ram_mem3_reg[242][29]/P0001 ,
		_w12932_,
		_w13763_
	);
	LUT2 #(
		.INIT('h1)
	) name3252 (
		_w13508_,
		_w13509_,
		_w13764_
	);
	LUT2 #(
		.INIT('h1)
	) name3253 (
		_w13510_,
		_w13511_,
		_w13765_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w13512_,
		_w13513_,
		_w13766_
	);
	LUT2 #(
		.INIT('h1)
	) name3255 (
		_w13514_,
		_w13515_,
		_w13767_
	);
	LUT2 #(
		.INIT('h1)
	) name3256 (
		_w13516_,
		_w13517_,
		_w13768_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w13518_,
		_w13519_,
		_w13769_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w13520_,
		_w13521_,
		_w13770_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w13522_,
		_w13523_,
		_w13771_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		_w13524_,
		_w13525_,
		_w13772_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w13526_,
		_w13527_,
		_w13773_
	);
	LUT2 #(
		.INIT('h1)
	) name3262 (
		_w13528_,
		_w13529_,
		_w13774_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		_w13530_,
		_w13531_,
		_w13775_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		_w13532_,
		_w13533_,
		_w13776_
	);
	LUT2 #(
		.INIT('h1)
	) name3265 (
		_w13534_,
		_w13535_,
		_w13777_
	);
	LUT2 #(
		.INIT('h1)
	) name3266 (
		_w13536_,
		_w13537_,
		_w13778_
	);
	LUT2 #(
		.INIT('h1)
	) name3267 (
		_w13538_,
		_w13539_,
		_w13779_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w13540_,
		_w13541_,
		_w13780_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w13542_,
		_w13543_,
		_w13781_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w13544_,
		_w13545_,
		_w13782_
	);
	LUT2 #(
		.INIT('h1)
	) name3271 (
		_w13546_,
		_w13547_,
		_w13783_
	);
	LUT2 #(
		.INIT('h1)
	) name3272 (
		_w13548_,
		_w13549_,
		_w13784_
	);
	LUT2 #(
		.INIT('h1)
	) name3273 (
		_w13550_,
		_w13551_,
		_w13785_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		_w13552_,
		_w13553_,
		_w13786_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w13554_,
		_w13555_,
		_w13787_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w13556_,
		_w13557_,
		_w13788_
	);
	LUT2 #(
		.INIT('h1)
	) name3277 (
		_w13558_,
		_w13559_,
		_w13789_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w13560_,
		_w13561_,
		_w13790_
	);
	LUT2 #(
		.INIT('h1)
	) name3279 (
		_w13562_,
		_w13563_,
		_w13791_
	);
	LUT2 #(
		.INIT('h1)
	) name3280 (
		_w13564_,
		_w13565_,
		_w13792_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w13566_,
		_w13567_,
		_w13793_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w13568_,
		_w13569_,
		_w13794_
	);
	LUT2 #(
		.INIT('h1)
	) name3283 (
		_w13570_,
		_w13571_,
		_w13795_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w13572_,
		_w13573_,
		_w13796_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w13574_,
		_w13575_,
		_w13797_
	);
	LUT2 #(
		.INIT('h1)
	) name3286 (
		_w13576_,
		_w13577_,
		_w13798_
	);
	LUT2 #(
		.INIT('h1)
	) name3287 (
		_w13578_,
		_w13579_,
		_w13799_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w13580_,
		_w13581_,
		_w13800_
	);
	LUT2 #(
		.INIT('h1)
	) name3289 (
		_w13582_,
		_w13583_,
		_w13801_
	);
	LUT2 #(
		.INIT('h1)
	) name3290 (
		_w13584_,
		_w13585_,
		_w13802_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w13586_,
		_w13587_,
		_w13803_
	);
	LUT2 #(
		.INIT('h1)
	) name3292 (
		_w13588_,
		_w13589_,
		_w13804_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		_w13590_,
		_w13591_,
		_w13805_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w13592_,
		_w13593_,
		_w13806_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w13594_,
		_w13595_,
		_w13807_
	);
	LUT2 #(
		.INIT('h1)
	) name3296 (
		_w13596_,
		_w13597_,
		_w13808_
	);
	LUT2 #(
		.INIT('h1)
	) name3297 (
		_w13598_,
		_w13599_,
		_w13809_
	);
	LUT2 #(
		.INIT('h1)
	) name3298 (
		_w13600_,
		_w13601_,
		_w13810_
	);
	LUT2 #(
		.INIT('h1)
	) name3299 (
		_w13602_,
		_w13603_,
		_w13811_
	);
	LUT2 #(
		.INIT('h1)
	) name3300 (
		_w13604_,
		_w13605_,
		_w13812_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w13606_,
		_w13607_,
		_w13813_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		_w13608_,
		_w13609_,
		_w13814_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w13610_,
		_w13611_,
		_w13815_
	);
	LUT2 #(
		.INIT('h1)
	) name3304 (
		_w13612_,
		_w13613_,
		_w13816_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		_w13614_,
		_w13615_,
		_w13817_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w13616_,
		_w13617_,
		_w13818_
	);
	LUT2 #(
		.INIT('h1)
	) name3307 (
		_w13618_,
		_w13619_,
		_w13819_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w13620_,
		_w13621_,
		_w13820_
	);
	LUT2 #(
		.INIT('h1)
	) name3309 (
		_w13622_,
		_w13623_,
		_w13821_
	);
	LUT2 #(
		.INIT('h1)
	) name3310 (
		_w13624_,
		_w13625_,
		_w13822_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		_w13626_,
		_w13627_,
		_w13823_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w13628_,
		_w13629_,
		_w13824_
	);
	LUT2 #(
		.INIT('h1)
	) name3313 (
		_w13630_,
		_w13631_,
		_w13825_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		_w13632_,
		_w13633_,
		_w13826_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w13634_,
		_w13635_,
		_w13827_
	);
	LUT2 #(
		.INIT('h1)
	) name3316 (
		_w13636_,
		_w13637_,
		_w13828_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		_w13638_,
		_w13639_,
		_w13829_
	);
	LUT2 #(
		.INIT('h1)
	) name3318 (
		_w13640_,
		_w13641_,
		_w13830_
	);
	LUT2 #(
		.INIT('h1)
	) name3319 (
		_w13642_,
		_w13643_,
		_w13831_
	);
	LUT2 #(
		.INIT('h1)
	) name3320 (
		_w13644_,
		_w13645_,
		_w13832_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		_w13646_,
		_w13647_,
		_w13833_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		_w13648_,
		_w13649_,
		_w13834_
	);
	LUT2 #(
		.INIT('h1)
	) name3323 (
		_w13650_,
		_w13651_,
		_w13835_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		_w13652_,
		_w13653_,
		_w13836_
	);
	LUT2 #(
		.INIT('h1)
	) name3325 (
		_w13654_,
		_w13655_,
		_w13837_
	);
	LUT2 #(
		.INIT('h1)
	) name3326 (
		_w13656_,
		_w13657_,
		_w13838_
	);
	LUT2 #(
		.INIT('h1)
	) name3327 (
		_w13658_,
		_w13659_,
		_w13839_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w13660_,
		_w13661_,
		_w13840_
	);
	LUT2 #(
		.INIT('h1)
	) name3329 (
		_w13662_,
		_w13663_,
		_w13841_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		_w13664_,
		_w13665_,
		_w13842_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w13666_,
		_w13667_,
		_w13843_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w13668_,
		_w13669_,
		_w13844_
	);
	LUT2 #(
		.INIT('h1)
	) name3333 (
		_w13670_,
		_w13671_,
		_w13845_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		_w13672_,
		_w13673_,
		_w13846_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w13674_,
		_w13675_,
		_w13847_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w13676_,
		_w13677_,
		_w13848_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w13678_,
		_w13679_,
		_w13849_
	);
	LUT2 #(
		.INIT('h1)
	) name3338 (
		_w13680_,
		_w13681_,
		_w13850_
	);
	LUT2 #(
		.INIT('h1)
	) name3339 (
		_w13682_,
		_w13683_,
		_w13851_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w13684_,
		_w13685_,
		_w13852_
	);
	LUT2 #(
		.INIT('h1)
	) name3341 (
		_w13686_,
		_w13687_,
		_w13853_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w13688_,
		_w13689_,
		_w13854_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w13690_,
		_w13691_,
		_w13855_
	);
	LUT2 #(
		.INIT('h1)
	) name3344 (
		_w13692_,
		_w13693_,
		_w13856_
	);
	LUT2 #(
		.INIT('h1)
	) name3345 (
		_w13694_,
		_w13695_,
		_w13857_
	);
	LUT2 #(
		.INIT('h1)
	) name3346 (
		_w13696_,
		_w13697_,
		_w13858_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w13698_,
		_w13699_,
		_w13859_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w13700_,
		_w13701_,
		_w13860_
	);
	LUT2 #(
		.INIT('h1)
	) name3349 (
		_w13702_,
		_w13703_,
		_w13861_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w13704_,
		_w13705_,
		_w13862_
	);
	LUT2 #(
		.INIT('h1)
	) name3351 (
		_w13706_,
		_w13707_,
		_w13863_
	);
	LUT2 #(
		.INIT('h1)
	) name3352 (
		_w13708_,
		_w13709_,
		_w13864_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w13710_,
		_w13711_,
		_w13865_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w13712_,
		_w13713_,
		_w13866_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w13714_,
		_w13715_,
		_w13867_
	);
	LUT2 #(
		.INIT('h1)
	) name3356 (
		_w13716_,
		_w13717_,
		_w13868_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w13718_,
		_w13719_,
		_w13869_
	);
	LUT2 #(
		.INIT('h1)
	) name3358 (
		_w13720_,
		_w13721_,
		_w13870_
	);
	LUT2 #(
		.INIT('h1)
	) name3359 (
		_w13722_,
		_w13723_,
		_w13871_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		_w13724_,
		_w13725_,
		_w13872_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w13726_,
		_w13727_,
		_w13873_
	);
	LUT2 #(
		.INIT('h1)
	) name3362 (
		_w13728_,
		_w13729_,
		_w13874_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		_w13730_,
		_w13731_,
		_w13875_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w13732_,
		_w13733_,
		_w13876_
	);
	LUT2 #(
		.INIT('h1)
	) name3365 (
		_w13734_,
		_w13735_,
		_w13877_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		_w13736_,
		_w13737_,
		_w13878_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w13738_,
		_w13739_,
		_w13879_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w13740_,
		_w13741_,
		_w13880_
	);
	LUT2 #(
		.INIT('h1)
	) name3369 (
		_w13742_,
		_w13743_,
		_w13881_
	);
	LUT2 #(
		.INIT('h1)
	) name3370 (
		_w13744_,
		_w13745_,
		_w13882_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w13746_,
		_w13747_,
		_w13883_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		_w13748_,
		_w13749_,
		_w13884_
	);
	LUT2 #(
		.INIT('h1)
	) name3373 (
		_w13750_,
		_w13751_,
		_w13885_
	);
	LUT2 #(
		.INIT('h1)
	) name3374 (
		_w13752_,
		_w13753_,
		_w13886_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w13754_,
		_w13755_,
		_w13887_
	);
	LUT2 #(
		.INIT('h1)
	) name3376 (
		_w13756_,
		_w13757_,
		_w13888_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		_w13758_,
		_w13759_,
		_w13889_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w13760_,
		_w13761_,
		_w13890_
	);
	LUT2 #(
		.INIT('h1)
	) name3379 (
		_w13762_,
		_w13763_,
		_w13891_
	);
	LUT2 #(
		.INIT('h8)
	) name3380 (
		_w13890_,
		_w13891_,
		_w13892_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		_w13888_,
		_w13889_,
		_w13893_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		_w13886_,
		_w13887_,
		_w13894_
	);
	LUT2 #(
		.INIT('h8)
	) name3383 (
		_w13884_,
		_w13885_,
		_w13895_
	);
	LUT2 #(
		.INIT('h8)
	) name3384 (
		_w13882_,
		_w13883_,
		_w13896_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		_w13880_,
		_w13881_,
		_w13897_
	);
	LUT2 #(
		.INIT('h8)
	) name3386 (
		_w13878_,
		_w13879_,
		_w13898_
	);
	LUT2 #(
		.INIT('h8)
	) name3387 (
		_w13876_,
		_w13877_,
		_w13899_
	);
	LUT2 #(
		.INIT('h8)
	) name3388 (
		_w13874_,
		_w13875_,
		_w13900_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w13872_,
		_w13873_,
		_w13901_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		_w13870_,
		_w13871_,
		_w13902_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w13868_,
		_w13869_,
		_w13903_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		_w13866_,
		_w13867_,
		_w13904_
	);
	LUT2 #(
		.INIT('h8)
	) name3393 (
		_w13864_,
		_w13865_,
		_w13905_
	);
	LUT2 #(
		.INIT('h8)
	) name3394 (
		_w13862_,
		_w13863_,
		_w13906_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		_w13860_,
		_w13861_,
		_w13907_
	);
	LUT2 #(
		.INIT('h8)
	) name3396 (
		_w13858_,
		_w13859_,
		_w13908_
	);
	LUT2 #(
		.INIT('h8)
	) name3397 (
		_w13856_,
		_w13857_,
		_w13909_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		_w13854_,
		_w13855_,
		_w13910_
	);
	LUT2 #(
		.INIT('h8)
	) name3399 (
		_w13852_,
		_w13853_,
		_w13911_
	);
	LUT2 #(
		.INIT('h8)
	) name3400 (
		_w13850_,
		_w13851_,
		_w13912_
	);
	LUT2 #(
		.INIT('h8)
	) name3401 (
		_w13848_,
		_w13849_,
		_w13913_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		_w13846_,
		_w13847_,
		_w13914_
	);
	LUT2 #(
		.INIT('h8)
	) name3403 (
		_w13844_,
		_w13845_,
		_w13915_
	);
	LUT2 #(
		.INIT('h8)
	) name3404 (
		_w13842_,
		_w13843_,
		_w13916_
	);
	LUT2 #(
		.INIT('h8)
	) name3405 (
		_w13840_,
		_w13841_,
		_w13917_
	);
	LUT2 #(
		.INIT('h8)
	) name3406 (
		_w13838_,
		_w13839_,
		_w13918_
	);
	LUT2 #(
		.INIT('h8)
	) name3407 (
		_w13836_,
		_w13837_,
		_w13919_
	);
	LUT2 #(
		.INIT('h8)
	) name3408 (
		_w13834_,
		_w13835_,
		_w13920_
	);
	LUT2 #(
		.INIT('h8)
	) name3409 (
		_w13832_,
		_w13833_,
		_w13921_
	);
	LUT2 #(
		.INIT('h8)
	) name3410 (
		_w13830_,
		_w13831_,
		_w13922_
	);
	LUT2 #(
		.INIT('h8)
	) name3411 (
		_w13828_,
		_w13829_,
		_w13923_
	);
	LUT2 #(
		.INIT('h8)
	) name3412 (
		_w13826_,
		_w13827_,
		_w13924_
	);
	LUT2 #(
		.INIT('h8)
	) name3413 (
		_w13824_,
		_w13825_,
		_w13925_
	);
	LUT2 #(
		.INIT('h8)
	) name3414 (
		_w13822_,
		_w13823_,
		_w13926_
	);
	LUT2 #(
		.INIT('h8)
	) name3415 (
		_w13820_,
		_w13821_,
		_w13927_
	);
	LUT2 #(
		.INIT('h8)
	) name3416 (
		_w13818_,
		_w13819_,
		_w13928_
	);
	LUT2 #(
		.INIT('h8)
	) name3417 (
		_w13816_,
		_w13817_,
		_w13929_
	);
	LUT2 #(
		.INIT('h8)
	) name3418 (
		_w13814_,
		_w13815_,
		_w13930_
	);
	LUT2 #(
		.INIT('h8)
	) name3419 (
		_w13812_,
		_w13813_,
		_w13931_
	);
	LUT2 #(
		.INIT('h8)
	) name3420 (
		_w13810_,
		_w13811_,
		_w13932_
	);
	LUT2 #(
		.INIT('h8)
	) name3421 (
		_w13808_,
		_w13809_,
		_w13933_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		_w13806_,
		_w13807_,
		_w13934_
	);
	LUT2 #(
		.INIT('h8)
	) name3423 (
		_w13804_,
		_w13805_,
		_w13935_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		_w13802_,
		_w13803_,
		_w13936_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		_w13800_,
		_w13801_,
		_w13937_
	);
	LUT2 #(
		.INIT('h8)
	) name3426 (
		_w13798_,
		_w13799_,
		_w13938_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		_w13796_,
		_w13797_,
		_w13939_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		_w13794_,
		_w13795_,
		_w13940_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		_w13792_,
		_w13793_,
		_w13941_
	);
	LUT2 #(
		.INIT('h8)
	) name3430 (
		_w13790_,
		_w13791_,
		_w13942_
	);
	LUT2 #(
		.INIT('h8)
	) name3431 (
		_w13788_,
		_w13789_,
		_w13943_
	);
	LUT2 #(
		.INIT('h8)
	) name3432 (
		_w13786_,
		_w13787_,
		_w13944_
	);
	LUT2 #(
		.INIT('h8)
	) name3433 (
		_w13784_,
		_w13785_,
		_w13945_
	);
	LUT2 #(
		.INIT('h8)
	) name3434 (
		_w13782_,
		_w13783_,
		_w13946_
	);
	LUT2 #(
		.INIT('h8)
	) name3435 (
		_w13780_,
		_w13781_,
		_w13947_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		_w13778_,
		_w13779_,
		_w13948_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w13776_,
		_w13777_,
		_w13949_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w13774_,
		_w13775_,
		_w13950_
	);
	LUT2 #(
		.INIT('h8)
	) name3439 (
		_w13772_,
		_w13773_,
		_w13951_
	);
	LUT2 #(
		.INIT('h8)
	) name3440 (
		_w13770_,
		_w13771_,
		_w13952_
	);
	LUT2 #(
		.INIT('h8)
	) name3441 (
		_w13768_,
		_w13769_,
		_w13953_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		_w13766_,
		_w13767_,
		_w13954_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		_w13764_,
		_w13765_,
		_w13955_
	);
	LUT2 #(
		.INIT('h8)
	) name3444 (
		_w13954_,
		_w13955_,
		_w13956_
	);
	LUT2 #(
		.INIT('h8)
	) name3445 (
		_w13952_,
		_w13953_,
		_w13957_
	);
	LUT2 #(
		.INIT('h8)
	) name3446 (
		_w13950_,
		_w13951_,
		_w13958_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		_w13948_,
		_w13949_,
		_w13959_
	);
	LUT2 #(
		.INIT('h8)
	) name3448 (
		_w13946_,
		_w13947_,
		_w13960_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		_w13944_,
		_w13945_,
		_w13961_
	);
	LUT2 #(
		.INIT('h8)
	) name3450 (
		_w13942_,
		_w13943_,
		_w13962_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		_w13940_,
		_w13941_,
		_w13963_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		_w13938_,
		_w13939_,
		_w13964_
	);
	LUT2 #(
		.INIT('h8)
	) name3453 (
		_w13936_,
		_w13937_,
		_w13965_
	);
	LUT2 #(
		.INIT('h8)
	) name3454 (
		_w13934_,
		_w13935_,
		_w13966_
	);
	LUT2 #(
		.INIT('h8)
	) name3455 (
		_w13932_,
		_w13933_,
		_w13967_
	);
	LUT2 #(
		.INIT('h8)
	) name3456 (
		_w13930_,
		_w13931_,
		_w13968_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		_w13928_,
		_w13929_,
		_w13969_
	);
	LUT2 #(
		.INIT('h8)
	) name3458 (
		_w13926_,
		_w13927_,
		_w13970_
	);
	LUT2 #(
		.INIT('h8)
	) name3459 (
		_w13924_,
		_w13925_,
		_w13971_
	);
	LUT2 #(
		.INIT('h8)
	) name3460 (
		_w13922_,
		_w13923_,
		_w13972_
	);
	LUT2 #(
		.INIT('h8)
	) name3461 (
		_w13920_,
		_w13921_,
		_w13973_
	);
	LUT2 #(
		.INIT('h8)
	) name3462 (
		_w13918_,
		_w13919_,
		_w13974_
	);
	LUT2 #(
		.INIT('h8)
	) name3463 (
		_w13916_,
		_w13917_,
		_w13975_
	);
	LUT2 #(
		.INIT('h8)
	) name3464 (
		_w13914_,
		_w13915_,
		_w13976_
	);
	LUT2 #(
		.INIT('h8)
	) name3465 (
		_w13912_,
		_w13913_,
		_w13977_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		_w13910_,
		_w13911_,
		_w13978_
	);
	LUT2 #(
		.INIT('h8)
	) name3467 (
		_w13908_,
		_w13909_,
		_w13979_
	);
	LUT2 #(
		.INIT('h8)
	) name3468 (
		_w13906_,
		_w13907_,
		_w13980_
	);
	LUT2 #(
		.INIT('h8)
	) name3469 (
		_w13904_,
		_w13905_,
		_w13981_
	);
	LUT2 #(
		.INIT('h8)
	) name3470 (
		_w13902_,
		_w13903_,
		_w13982_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		_w13900_,
		_w13901_,
		_w13983_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		_w13898_,
		_w13899_,
		_w13984_
	);
	LUT2 #(
		.INIT('h8)
	) name3473 (
		_w13896_,
		_w13897_,
		_w13985_
	);
	LUT2 #(
		.INIT('h8)
	) name3474 (
		_w13894_,
		_w13895_,
		_w13986_
	);
	LUT2 #(
		.INIT('h8)
	) name3475 (
		_w13892_,
		_w13893_,
		_w13987_
	);
	LUT2 #(
		.INIT('h8)
	) name3476 (
		_w13986_,
		_w13987_,
		_w13988_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		_w13984_,
		_w13985_,
		_w13989_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		_w13982_,
		_w13983_,
		_w13990_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		_w13980_,
		_w13981_,
		_w13991_
	);
	LUT2 #(
		.INIT('h8)
	) name3480 (
		_w13978_,
		_w13979_,
		_w13992_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		_w13976_,
		_w13977_,
		_w13993_
	);
	LUT2 #(
		.INIT('h8)
	) name3482 (
		_w13974_,
		_w13975_,
		_w13994_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w13972_,
		_w13973_,
		_w13995_
	);
	LUT2 #(
		.INIT('h8)
	) name3484 (
		_w13970_,
		_w13971_,
		_w13996_
	);
	LUT2 #(
		.INIT('h8)
	) name3485 (
		_w13968_,
		_w13969_,
		_w13997_
	);
	LUT2 #(
		.INIT('h8)
	) name3486 (
		_w13966_,
		_w13967_,
		_w13998_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		_w13964_,
		_w13965_,
		_w13999_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		_w13962_,
		_w13963_,
		_w14000_
	);
	LUT2 #(
		.INIT('h8)
	) name3489 (
		_w13960_,
		_w13961_,
		_w14001_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		_w13958_,
		_w13959_,
		_w14002_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		_w13956_,
		_w13957_,
		_w14003_
	);
	LUT2 #(
		.INIT('h8)
	) name3492 (
		_w14002_,
		_w14003_,
		_w14004_
	);
	LUT2 #(
		.INIT('h8)
	) name3493 (
		_w14000_,
		_w14001_,
		_w14005_
	);
	LUT2 #(
		.INIT('h8)
	) name3494 (
		_w13998_,
		_w13999_,
		_w14006_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		_w13996_,
		_w13997_,
		_w14007_
	);
	LUT2 #(
		.INIT('h8)
	) name3496 (
		_w13994_,
		_w13995_,
		_w14008_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		_w13992_,
		_w13993_,
		_w14009_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		_w13990_,
		_w13991_,
		_w14010_
	);
	LUT2 #(
		.INIT('h8)
	) name3499 (
		_w13988_,
		_w13989_,
		_w14011_
	);
	LUT2 #(
		.INIT('h8)
	) name3500 (
		_w14010_,
		_w14011_,
		_w14012_
	);
	LUT2 #(
		.INIT('h8)
	) name3501 (
		_w14008_,
		_w14009_,
		_w14013_
	);
	LUT2 #(
		.INIT('h8)
	) name3502 (
		_w14006_,
		_w14007_,
		_w14014_
	);
	LUT2 #(
		.INIT('h8)
	) name3503 (
		_w14004_,
		_w14005_,
		_w14015_
	);
	LUT2 #(
		.INIT('h8)
	) name3504 (
		_w14014_,
		_w14015_,
		_w14016_
	);
	LUT2 #(
		.INIT('h8)
	) name3505 (
		_w14012_,
		_w14013_,
		_w14017_
	);
	LUT2 #(
		.INIT('h8)
	) name3506 (
		_w14016_,
		_w14017_,
		_w14018_
	);
	LUT2 #(
		.INIT('h1)
	) name3507 (
		wb_rst_i_pad,
		_w14018_,
		_w14019_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		_w12656_,
		_w14019_,
		_w14020_
	);
	LUT2 #(
		.INIT('h8)
	) name3509 (
		_w13491_,
		_w13495_,
		_w14021_
	);
	LUT2 #(
		.INIT('h8)
	) name3510 (
		_w13501_,
		_w14021_,
		_w14022_
	);
	LUT2 #(
		.INIT('h1)
	) name3511 (
		_w13507_,
		_w14022_,
		_w14023_
	);
	LUT2 #(
		.INIT('h4)
	) name3512 (
		_w14020_,
		_w14023_,
		_w14024_
	);
	LUT2 #(
		.INIT('h8)
	) name3513 (
		\wishbone_bd_ram_mem3_reg[164][30]/P0001 ,
		_w12876_,
		_w14025_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		\wishbone_bd_ram_mem3_reg[135][30]/P0001 ,
		_w13124_,
		_w14026_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		\wishbone_bd_ram_mem3_reg[19][30]/P0001 ,
		_w13012_,
		_w14027_
	);
	LUT2 #(
		.INIT('h8)
	) name3516 (
		\wishbone_bd_ram_mem3_reg[103][30]/P0001 ,
		_w12846_,
		_w14028_
	);
	LUT2 #(
		.INIT('h8)
	) name3517 (
		\wishbone_bd_ram_mem3_reg[20][30]/P0001 ,
		_w13174_,
		_w14029_
	);
	LUT2 #(
		.INIT('h8)
	) name3518 (
		\wishbone_bd_ram_mem3_reg[224][30]/P0001 ,
		_w12902_,
		_w14030_
	);
	LUT2 #(
		.INIT('h8)
	) name3519 (
		\wishbone_bd_ram_mem3_reg[60][30]/P0001 ,
		_w13204_,
		_w14031_
	);
	LUT2 #(
		.INIT('h8)
	) name3520 (
		\wishbone_bd_ram_mem3_reg[36][30]/P0001 ,
		_w12800_,
		_w14032_
	);
	LUT2 #(
		.INIT('h8)
	) name3521 (
		\wishbone_bd_ram_mem3_reg[89][30]/P0001 ,
		_w12964_,
		_w14033_
	);
	LUT2 #(
		.INIT('h8)
	) name3522 (
		\wishbone_bd_ram_mem3_reg[250][30]/P0001 ,
		_w13128_,
		_w14034_
	);
	LUT2 #(
		.INIT('h8)
	) name3523 (
		\wishbone_bd_ram_mem3_reg[185][30]/P0001 ,
		_w12940_,
		_w14035_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		\wishbone_bd_ram_mem3_reg[100][30]/P0001 ,
		_w12960_,
		_w14036_
	);
	LUT2 #(
		.INIT('h8)
	) name3525 (
		\wishbone_bd_ram_mem3_reg[9][30]/P0001 ,
		_w12808_,
		_w14037_
	);
	LUT2 #(
		.INIT('h8)
	) name3526 (
		\wishbone_bd_ram_mem3_reg[97][30]/P0001 ,
		_w13096_,
		_w14038_
	);
	LUT2 #(
		.INIT('h8)
	) name3527 (
		\wishbone_bd_ram_mem3_reg[149][30]/P0001 ,
		_w12741_,
		_w14039_
	);
	LUT2 #(
		.INIT('h8)
	) name3528 (
		\wishbone_bd_ram_mem3_reg[28][30]/P0001 ,
		_w13170_,
		_w14040_
	);
	LUT2 #(
		.INIT('h8)
	) name3529 (
		\wishbone_bd_ram_mem3_reg[255][30]/P0001 ,
		_w13072_,
		_w14041_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		\wishbone_bd_ram_mem3_reg[87][30]/P0001 ,
		_w13154_,
		_w14042_
	);
	LUT2 #(
		.INIT('h8)
	) name3531 (
		\wishbone_bd_ram_mem3_reg[0][30]/P0001 ,
		_w12717_,
		_w14043_
	);
	LUT2 #(
		.INIT('h8)
	) name3532 (
		\wishbone_bd_ram_mem3_reg[18][30]/P0001 ,
		_w12679_,
		_w14044_
	);
	LUT2 #(
		.INIT('h8)
	) name3533 (
		\wishbone_bd_ram_mem3_reg[34][30]/P0001 ,
		_w12930_,
		_w14045_
	);
	LUT2 #(
		.INIT('h8)
	) name3534 (
		\wishbone_bd_ram_mem3_reg[169][30]/P0001 ,
		_w12722_,
		_w14046_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		\wishbone_bd_ram_mem3_reg[200][30]/P0001 ,
		_w12988_,
		_w14047_
	);
	LUT2 #(
		.INIT('h8)
	) name3536 (
		\wishbone_bd_ram_mem3_reg[230][30]/P0001 ,
		_w13036_,
		_w14048_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		\wishbone_bd_ram_mem3_reg[112][30]/P0001 ,
		_w12733_,
		_w14049_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		\wishbone_bd_ram_mem3_reg[86][30]/P0001 ,
		_w12735_,
		_w14050_
	);
	LUT2 #(
		.INIT('h8)
	) name3539 (
		\wishbone_bd_ram_mem3_reg[153][30]/P0001 ,
		_w12890_,
		_w14051_
	);
	LUT2 #(
		.INIT('h8)
	) name3540 (
		\wishbone_bd_ram_mem3_reg[234][30]/P0001 ,
		_w13214_,
		_w14052_
	);
	LUT2 #(
		.INIT('h8)
	) name3541 (
		\wishbone_bd_ram_mem3_reg[186][30]/P0001 ,
		_w12783_,
		_w14053_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		\wishbone_bd_ram_mem3_reg[136][30]/P0001 ,
		_w13064_,
		_w14054_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		\wishbone_bd_ram_mem3_reg[158][30]/P0001 ,
		_w12898_,
		_w14055_
	);
	LUT2 #(
		.INIT('h8)
	) name3544 (
		\wishbone_bd_ram_mem3_reg[212][30]/P0001 ,
		_w12796_,
		_w14056_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		\wishbone_bd_ram_mem3_reg[59][30]/P0001 ,
		_w12780_,
		_w14057_
	);
	LUT2 #(
		.INIT('h8)
	) name3546 (
		\wishbone_bd_ram_mem3_reg[134][30]/P0001 ,
		_w12763_,
		_w14058_
	);
	LUT2 #(
		.INIT('h8)
	) name3547 (
		\wishbone_bd_ram_mem3_reg[23][30]/P0001 ,
		_w13008_,
		_w14059_
	);
	LUT2 #(
		.INIT('h8)
	) name3548 (
		\wishbone_bd_ram_mem3_reg[142][30]/P0001 ,
		_w12928_,
		_w14060_
	);
	LUT2 #(
		.INIT('h8)
	) name3549 (
		\wishbone_bd_ram_mem3_reg[47][30]/P0001 ,
		_w12904_,
		_w14061_
	);
	LUT2 #(
		.INIT('h8)
	) name3550 (
		\wishbone_bd_ram_mem3_reg[54][30]/P0001 ,
		_w12770_,
		_w14062_
	);
	LUT2 #(
		.INIT('h8)
	) name3551 (
		\wishbone_bd_ram_mem3_reg[139][30]/P0001 ,
		_w12814_,
		_w14063_
	);
	LUT2 #(
		.INIT('h8)
	) name3552 (
		\wishbone_bd_ram_mem3_reg[239][30]/P0001 ,
		_w12862_,
		_w14064_
	);
	LUT2 #(
		.INIT('h8)
	) name3553 (
		\wishbone_bd_ram_mem3_reg[243][30]/P0001 ,
		_w12804_,
		_w14065_
	);
	LUT2 #(
		.INIT('h8)
	) name3554 (
		\wishbone_bd_ram_mem3_reg[219][30]/P0001 ,
		_w12806_,
		_w14066_
	);
	LUT2 #(
		.INIT('h8)
	) name3555 (
		\wishbone_bd_ram_mem3_reg[189][30]/P0001 ,
		_w13042_,
		_w14067_
	);
	LUT2 #(
		.INIT('h8)
	) name3556 (
		\wishbone_bd_ram_mem3_reg[141][30]/P0001 ,
		_w13004_,
		_w14068_
	);
	LUT2 #(
		.INIT('h8)
	) name3557 (
		\wishbone_bd_ram_mem3_reg[179][30]/P0001 ,
		_w13050_,
		_w14069_
	);
	LUT2 #(
		.INIT('h8)
	) name3558 (
		\wishbone_bd_ram_mem3_reg[53][30]/P0001 ,
		_w13020_,
		_w14070_
	);
	LUT2 #(
		.INIT('h8)
	) name3559 (
		\wishbone_bd_ram_mem3_reg[6][30]/P0001 ,
		_w12968_,
		_w14071_
	);
	LUT2 #(
		.INIT('h8)
	) name3560 (
		\wishbone_bd_ram_mem3_reg[254][30]/P0001 ,
		_w12892_,
		_w14072_
	);
	LUT2 #(
		.INIT('h8)
	) name3561 (
		\wishbone_bd_ram_mem3_reg[236][30]/P0001 ,
		_w12731_,
		_w14073_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\wishbone_bd_ram_mem3_reg[187][30]/P0001 ,
		_w13196_,
		_w14074_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		\wishbone_bd_ram_mem3_reg[13][30]/P0001 ,
		_w13178_,
		_w14075_
	);
	LUT2 #(
		.INIT('h8)
	) name3564 (
		\wishbone_bd_ram_mem3_reg[26][30]/P0001 ,
		_w12699_,
		_w14076_
	);
	LUT2 #(
		.INIT('h8)
	) name3565 (
		\wishbone_bd_ram_mem3_reg[129][30]/P0001 ,
		_w12776_,
		_w14077_
	);
	LUT2 #(
		.INIT('h8)
	) name3566 (
		\wishbone_bd_ram_mem3_reg[91][30]/P0001 ,
		_w13074_,
		_w14078_
	);
	LUT2 #(
		.INIT('h8)
	) name3567 (
		\wishbone_bd_ram_mem3_reg[166][30]/P0001 ,
		_w13040_,
		_w14079_
	);
	LUT2 #(
		.INIT('h8)
	) name3568 (
		\wishbone_bd_ram_mem3_reg[204][30]/P0001 ,
		_w13162_,
		_w14080_
	);
	LUT2 #(
		.INIT('h8)
	) name3569 (
		\wishbone_bd_ram_mem3_reg[96][30]/P0001 ,
		_w12912_,
		_w14081_
	);
	LUT2 #(
		.INIT('h8)
	) name3570 (
		\wishbone_bd_ram_mem3_reg[190][30]/P0001 ,
		_w12858_,
		_w14082_
	);
	LUT2 #(
		.INIT('h8)
	) name3571 (
		\wishbone_bd_ram_mem3_reg[92][30]/P0001 ,
		_w13010_,
		_w14083_
	);
	LUT2 #(
		.INIT('h8)
	) name3572 (
		\wishbone_bd_ram_mem3_reg[117][30]/P0001 ,
		_w12715_,
		_w14084_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		\wishbone_bd_ram_mem3_reg[178][30]/P0001 ,
		_w12886_,
		_w14085_
	);
	LUT2 #(
		.INIT('h8)
	) name3574 (
		\wishbone_bd_ram_mem3_reg[157][30]/P0001 ,
		_w12926_,
		_w14086_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		\wishbone_bd_ram_mem3_reg[176][30]/P0001 ,
		_w12868_,
		_w14087_
	);
	LUT2 #(
		.INIT('h8)
	) name3576 (
		\wishbone_bd_ram_mem3_reg[235][30]/P0001 ,
		_w12696_,
		_w14088_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		\wishbone_bd_ram_mem3_reg[226][30]/P0001 ,
		_w13138_,
		_w14089_
	);
	LUT2 #(
		.INIT('h8)
	) name3578 (
		\wishbone_bd_ram_mem3_reg[199][30]/P0001 ,
		_w12768_,
		_w14090_
	);
	LUT2 #(
		.INIT('h8)
	) name3579 (
		\wishbone_bd_ram_mem3_reg[32][30]/P0001 ,
		_w13120_,
		_w14091_
	);
	LUT2 #(
		.INIT('h8)
	) name3580 (
		\wishbone_bd_ram_mem3_reg[67][30]/P0001 ,
		_w13134_,
		_w14092_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		\wishbone_bd_ram_mem3_reg[104][30]/P0001 ,
		_w13148_,
		_w14093_
	);
	LUT2 #(
		.INIT('h8)
	) name3582 (
		\wishbone_bd_ram_mem3_reg[102][30]/P0001 ,
		_w12685_,
		_w14094_
	);
	LUT2 #(
		.INIT('h8)
	) name3583 (
		\wishbone_bd_ram_mem3_reg[50][30]/P0001 ,
		_w13150_,
		_w14095_
	);
	LUT2 #(
		.INIT('h8)
	) name3584 (
		\wishbone_bd_ram_mem3_reg[163][30]/P0001 ,
		_w12882_,
		_w14096_
	);
	LUT2 #(
		.INIT('h8)
	) name3585 (
		\wishbone_bd_ram_mem3_reg[58][30]/P0001 ,
		_w13070_,
		_w14097_
	);
	LUT2 #(
		.INIT('h8)
	) name3586 (
		\wishbone_bd_ram_mem3_reg[205][30]/P0001 ,
		_w13068_,
		_w14098_
	);
	LUT2 #(
		.INIT('h8)
	) name3587 (
		\wishbone_bd_ram_mem3_reg[144][30]/P0001 ,
		_w12756_,
		_w14099_
	);
	LUT2 #(
		.INIT('h8)
	) name3588 (
		\wishbone_bd_ram_mem3_reg[215][30]/P0001 ,
		_w12974_,
		_w14100_
	);
	LUT2 #(
		.INIT('h8)
	) name3589 (
		\wishbone_bd_ram_mem3_reg[182][30]/P0001 ,
		_w12820_,
		_w14101_
	);
	LUT2 #(
		.INIT('h8)
	) name3590 (
		\wishbone_bd_ram_mem3_reg[227][30]/P0001 ,
		_w12936_,
		_w14102_
	);
	LUT2 #(
		.INIT('h8)
	) name3591 (
		\wishbone_bd_ram_mem3_reg[216][30]/P0001 ,
		_w13028_,
		_w14103_
	);
	LUT2 #(
		.INIT('h8)
	) name3592 (
		\wishbone_bd_ram_mem3_reg[43][30]/P0001 ,
		_w13200_,
		_w14104_
	);
	LUT2 #(
		.INIT('h8)
	) name3593 (
		\wishbone_bd_ram_mem3_reg[132][30]/P0001 ,
		_w12992_,
		_w14105_
	);
	LUT2 #(
		.INIT('h8)
	) name3594 (
		\wishbone_bd_ram_mem3_reg[237][30]/P0001 ,
		_w12990_,
		_w14106_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		\wishbone_bd_ram_mem3_reg[119][30]/P0001 ,
		_w13048_,
		_w14107_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		\wishbone_bd_ram_mem3_reg[242][30]/P0001 ,
		_w12932_,
		_w14108_
	);
	LUT2 #(
		.INIT('h8)
	) name3597 (
		\wishbone_bd_ram_mem3_reg[64][30]/P0001 ,
		_w12976_,
		_w14109_
	);
	LUT2 #(
		.INIT('h8)
	) name3598 (
		\wishbone_bd_ram_mem3_reg[211][30]/P0001 ,
		_w13166_,
		_w14110_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		\wishbone_bd_ram_mem3_reg[1][30]/P0001 ,
		_w13014_,
		_w14111_
	);
	LUT2 #(
		.INIT('h8)
	) name3600 (
		\wishbone_bd_ram_mem3_reg[10][30]/P0001 ,
		_w13172_,
		_w14112_
	);
	LUT2 #(
		.INIT('h8)
	) name3601 (
		\wishbone_bd_ram_mem3_reg[109][30]/P0001 ,
		_w12888_,
		_w14113_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		\wishbone_bd_ram_mem3_reg[181][30]/P0001 ,
		_w12828_,
		_w14114_
	);
	LUT2 #(
		.INIT('h8)
	) name3603 (
		\wishbone_bd_ram_mem3_reg[74][30]/P0001 ,
		_w12812_,
		_w14115_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		\wishbone_bd_ram_mem3_reg[192][30]/P0001 ,
		_w12938_,
		_w14116_
	);
	LUT2 #(
		.INIT('h8)
	) name3605 (
		\wishbone_bd_ram_mem3_reg[206][30]/P0001 ,
		_w12954_,
		_w14117_
	);
	LUT2 #(
		.INIT('h8)
	) name3606 (
		\wishbone_bd_ram_mem3_reg[175][30]/P0001 ,
		_w13126_,
		_w14118_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\wishbone_bd_ram_mem3_reg[77][30]/P0001 ,
		_w12982_,
		_w14119_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		\wishbone_bd_ram_mem3_reg[232][30]/P0001 ,
		_w12758_,
		_w14120_
	);
	LUT2 #(
		.INIT('h8)
	) name3609 (
		\wishbone_bd_ram_mem3_reg[210][30]/P0001 ,
		_w12924_,
		_w14121_
	);
	LUT2 #(
		.INIT('h8)
	) name3610 (
		\wishbone_bd_ram_mem3_reg[180][30]/P0001 ,
		_w12791_,
		_w14122_
	);
	LUT2 #(
		.INIT('h8)
	) name3611 (
		\wishbone_bd_ram_mem3_reg[56][30]/P0001 ,
		_w12778_,
		_w14123_
	);
	LUT2 #(
		.INIT('h8)
	) name3612 (
		\wishbone_bd_ram_mem3_reg[27][30]/P0001 ,
		_w12880_,
		_w14124_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		\wishbone_bd_ram_mem3_reg[83][30]/P0001 ,
		_w12916_,
		_w14125_
	);
	LUT2 #(
		.INIT('h8)
	) name3614 (
		\wishbone_bd_ram_mem3_reg[130][30]/P0001 ,
		_w12914_,
		_w14126_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		\wishbone_bd_ram_mem3_reg[98][30]/P0001 ,
		_w12816_,
		_w14127_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		\wishbone_bd_ram_mem3_reg[146][30]/P0001 ,
		_w13060_,
		_w14128_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		\wishbone_bd_ram_mem3_reg[66][30]/P0001 ,
		_w12824_,
		_w14129_
	);
	LUT2 #(
		.INIT('h8)
	) name3618 (
		\wishbone_bd_ram_mem3_reg[15][30]/P0001 ,
		_w13210_,
		_w14130_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		\wishbone_bd_ram_mem3_reg[33][30]/P0001 ,
		_w12980_,
		_w14131_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		\wishbone_bd_ram_mem3_reg[174][30]/P0001 ,
		_w12972_,
		_w14132_
	);
	LUT2 #(
		.INIT('h8)
	) name3621 (
		\wishbone_bd_ram_mem3_reg[196][30]/P0001 ,
		_w13090_,
		_w14133_
	);
	LUT2 #(
		.INIT('h8)
	) name3622 (
		\wishbone_bd_ram_mem3_reg[61][30]/P0001 ,
		_w12725_,
		_w14134_
	);
	LUT2 #(
		.INIT('h8)
	) name3623 (
		\wishbone_bd_ram_mem3_reg[116][30]/P0001 ,
		_w12998_,
		_w14135_
	);
	LUT2 #(
		.INIT('h8)
	) name3624 (
		\wishbone_bd_ram_mem3_reg[148][30]/P0001 ,
		_w13000_,
		_w14136_
	);
	LUT2 #(
		.INIT('h8)
	) name3625 (
		\wishbone_bd_ram_mem3_reg[183][30]/P0001 ,
		_w12787_,
		_w14137_
	);
	LUT2 #(
		.INIT('h8)
	) name3626 (
		\wishbone_bd_ram_mem3_reg[131][30]/P0001 ,
		_w12852_,
		_w14138_
	);
	LUT2 #(
		.INIT('h8)
	) name3627 (
		\wishbone_bd_ram_mem3_reg[213][30]/P0001 ,
		_w13002_,
		_w14139_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		\wishbone_bd_ram_mem3_reg[156][30]/P0001 ,
		_w13190_,
		_w14140_
	);
	LUT2 #(
		.INIT('h8)
	) name3629 (
		\wishbone_bd_ram_mem3_reg[173][30]/P0001 ,
		_w12854_,
		_w14141_
	);
	LUT2 #(
		.INIT('h8)
	) name3630 (
		\wishbone_bd_ram_mem3_reg[123][30]/P0001 ,
		_w13114_,
		_w14142_
	);
	LUT2 #(
		.INIT('h8)
	) name3631 (
		\wishbone_bd_ram_mem3_reg[193][30]/P0001 ,
		_w13056_,
		_w14143_
	);
	LUT2 #(
		.INIT('h8)
	) name3632 (
		\wishbone_bd_ram_mem3_reg[3][30]/P0001 ,
		_w12866_,
		_w14144_
	);
	LUT2 #(
		.INIT('h8)
	) name3633 (
		\wishbone_bd_ram_mem3_reg[154][30]/P0001 ,
		_w12962_,
		_w14145_
	);
	LUT2 #(
		.INIT('h8)
	) name3634 (
		\wishbone_bd_ram_mem3_reg[252][30]/P0001 ,
		_w13080_,
		_w14146_
	);
	LUT2 #(
		.INIT('h8)
	) name3635 (
		\wishbone_bd_ram_mem3_reg[72][30]/P0001 ,
		_w12810_,
		_w14147_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		\wishbone_bd_ram_mem3_reg[229][30]/P0001 ,
		_w12711_,
		_w14148_
	);
	LUT2 #(
		.INIT('h8)
	) name3637 (
		\wishbone_bd_ram_mem3_reg[107][30]/P0001 ,
		_w12749_,
		_w14149_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		\wishbone_bd_ram_mem3_reg[73][30]/P0001 ,
		_w12918_,
		_w14150_
	);
	LUT2 #(
		.INIT('h8)
	) name3639 (
		\wishbone_bd_ram_mem3_reg[208][30]/P0001 ,
		_w13032_,
		_w14151_
	);
	LUT2 #(
		.INIT('h8)
	) name3640 (
		\wishbone_bd_ram_mem3_reg[241][30]/P0001 ,
		_w13006_,
		_w14152_
	);
	LUT2 #(
		.INIT('h8)
	) name3641 (
		\wishbone_bd_ram_mem3_reg[125][30]/P0001 ,
		_w12956_,
		_w14153_
	);
	LUT2 #(
		.INIT('h8)
	) name3642 (
		\wishbone_bd_ram_mem3_reg[122][30]/P0001 ,
		_w13130_,
		_w14154_
	);
	LUT2 #(
		.INIT('h8)
	) name3643 (
		\wishbone_bd_ram_mem3_reg[147][30]/P0001 ,
		_w13146_,
		_w14155_
	);
	LUT2 #(
		.INIT('h8)
	) name3644 (
		\wishbone_bd_ram_mem3_reg[31][30]/P0001 ,
		_w13198_,
		_w14156_
	);
	LUT2 #(
		.INIT('h8)
	) name3645 (
		\wishbone_bd_ram_mem3_reg[121][30]/P0001 ,
		_w13078_,
		_w14157_
	);
	LUT2 #(
		.INIT('h8)
	) name3646 (
		\wishbone_bd_ram_mem3_reg[11][30]/P0001 ,
		_w13194_,
		_w14158_
	);
	LUT2 #(
		.INIT('h8)
	) name3647 (
		\wishbone_bd_ram_mem3_reg[49][30]/P0001 ,
		_w12994_,
		_w14159_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		\wishbone_bd_ram_mem3_reg[145][30]/P0001 ,
		_w13106_,
		_w14160_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		\wishbone_bd_ram_mem3_reg[8][30]/P0001 ,
		_w12920_,
		_w14161_
	);
	LUT2 #(
		.INIT('h8)
	) name3650 (
		\wishbone_bd_ram_mem3_reg[39][30]/P0001 ,
		_w13018_,
		_w14162_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		\wishbone_bd_ram_mem3_reg[246][30]/P0001 ,
		_w13076_,
		_w14163_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		\wishbone_bd_ram_mem3_reg[138][30]/P0001 ,
		_w12958_,
		_w14164_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		\wishbone_bd_ram_mem3_reg[220][30]/P0001 ,
		_w13066_,
		_w14165_
	);
	LUT2 #(
		.INIT('h8)
	) name3654 (
		\wishbone_bd_ram_mem3_reg[188][30]/P0001 ,
		_w12948_,
		_w14166_
	);
	LUT2 #(
		.INIT('h8)
	) name3655 (
		\wishbone_bd_ram_mem3_reg[12][30]/P0001 ,
		_w13118_,
		_w14167_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		\wishbone_bd_ram_mem3_reg[38][30]/P0001 ,
		_w13182_,
		_w14168_
	);
	LUT2 #(
		.INIT('h8)
	) name3657 (
		\wishbone_bd_ram_mem3_reg[143][30]/P0001 ,
		_w12922_,
		_w14169_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		\wishbone_bd_ram_mem3_reg[75][30]/P0001 ,
		_w12826_,
		_w14170_
	);
	LUT2 #(
		.INIT('h8)
	) name3659 (
		\wishbone_bd_ram_mem3_reg[118][30]/P0001 ,
		_w12830_,
		_w14171_
	);
	LUT2 #(
		.INIT('h8)
	) name3660 (
		\wishbone_bd_ram_mem3_reg[194][30]/P0001 ,
		_w12772_,
		_w14172_
	);
	LUT2 #(
		.INIT('h8)
	) name3661 (
		\wishbone_bd_ram_mem3_reg[29][30]/P0001 ,
		_w12952_,
		_w14173_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		\wishbone_bd_ram_mem3_reg[184][30]/P0001 ,
		_w13062_,
		_w14174_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		\wishbone_bd_ram_mem3_reg[82][30]/P0001 ,
		_w12942_,
		_w14175_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		\wishbone_bd_ram_mem3_reg[63][30]/P0001 ,
		_w12850_,
		_w14176_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		\wishbone_bd_ram_mem3_reg[115][30]/P0001 ,
		_w13112_,
		_w14177_
	);
	LUT2 #(
		.INIT('h8)
	) name3666 (
		\wishbone_bd_ram_mem3_reg[37][30]/P0001 ,
		_w13102_,
		_w14178_
	);
	LUT2 #(
		.INIT('h8)
	) name3667 (
		\wishbone_bd_ram_mem3_reg[7][30]/P0001 ,
		_w12728_,
		_w14179_
	);
	LUT2 #(
		.INIT('h8)
	) name3668 (
		\wishbone_bd_ram_mem3_reg[68][30]/P0001 ,
		_w12946_,
		_w14180_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		\wishbone_bd_ram_mem3_reg[45][30]/P0001 ,
		_w12908_,
		_w14181_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		\wishbone_bd_ram_mem3_reg[225][30]/P0001 ,
		_w13092_,
		_w14182_
	);
	LUT2 #(
		.INIT('h8)
	) name3671 (
		\wishbone_bd_ram_mem3_reg[35][30]/P0001 ,
		_w12703_,
		_w14183_
	);
	LUT2 #(
		.INIT('h8)
	) name3672 (
		\wishbone_bd_ram_mem3_reg[127][30]/P0001 ,
		_w13164_,
		_w14184_
	);
	LUT2 #(
		.INIT('h8)
	) name3673 (
		\wishbone_bd_ram_mem3_reg[248][30]/P0001 ,
		_w12789_,
		_w14185_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		\wishbone_bd_ram_mem3_reg[126][30]/P0001 ,
		_w13218_,
		_w14186_
	);
	LUT2 #(
		.INIT('h8)
	) name3675 (
		\wishbone_bd_ram_mem3_reg[93][30]/P0001 ,
		_w13016_,
		_w14187_
	);
	LUT2 #(
		.INIT('h8)
	) name3676 (
		\wishbone_bd_ram_mem3_reg[140][30]/P0001 ,
		_w12894_,
		_w14188_
	);
	LUT2 #(
		.INIT('h8)
	) name3677 (
		\wishbone_bd_ram_mem3_reg[171][30]/P0001 ,
		_w12910_,
		_w14189_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		\wishbone_bd_ram_mem3_reg[150][30]/P0001 ,
		_w13136_,
		_w14190_
	);
	LUT2 #(
		.INIT('h8)
	) name3679 (
		\wishbone_bd_ram_mem3_reg[95][30]/P0001 ,
		_w12844_,
		_w14191_
	);
	LUT2 #(
		.INIT('h8)
	) name3680 (
		\wishbone_bd_ram_mem3_reg[90][30]/P0001 ,
		_w12978_,
		_w14192_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		\wishbone_bd_ram_mem3_reg[71][30]/P0001 ,
		_w12798_,
		_w14193_
	);
	LUT2 #(
		.INIT('h8)
	) name3682 (
		\wishbone_bd_ram_mem3_reg[124][30]/P0001 ,
		_w13058_,
		_w14194_
	);
	LUT2 #(
		.INIT('h8)
	) name3683 (
		\wishbone_bd_ram_mem3_reg[65][30]/P0001 ,
		_w13176_,
		_w14195_
	);
	LUT2 #(
		.INIT('h8)
	) name3684 (
		\wishbone_bd_ram_mem3_reg[177][30]/P0001 ,
		_w12996_,
		_w14196_
	);
	LUT2 #(
		.INIT('h8)
	) name3685 (
		\wishbone_bd_ram_mem3_reg[14][30]/P0001 ,
		_w13086_,
		_w14197_
	);
	LUT2 #(
		.INIT('h8)
	) name3686 (
		\wishbone_bd_ram_mem3_reg[249][30]/P0001 ,
		_w12900_,
		_w14198_
	);
	LUT2 #(
		.INIT('h8)
	) name3687 (
		\wishbone_bd_ram_mem3_reg[162][30]/P0001 ,
		_w13098_,
		_w14199_
	);
	LUT2 #(
		.INIT('h8)
	) name3688 (
		\wishbone_bd_ram_mem3_reg[110][30]/P0001 ,
		_w13046_,
		_w14200_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		\wishbone_bd_ram_mem3_reg[120][30]/P0001 ,
		_w12707_,
		_w14201_
	);
	LUT2 #(
		.INIT('h8)
	) name3690 (
		\wishbone_bd_ram_mem3_reg[202][30]/P0001 ,
		_w12870_,
		_w14202_
	);
	LUT2 #(
		.INIT('h8)
	) name3691 (
		\wishbone_bd_ram_mem3_reg[168][30]/P0001 ,
		_w13208_,
		_w14203_
	);
	LUT2 #(
		.INIT('h8)
	) name3692 (
		\wishbone_bd_ram_mem3_reg[247][30]/P0001 ,
		_w12818_,
		_w14204_
	);
	LUT2 #(
		.INIT('h8)
	) name3693 (
		\wishbone_bd_ram_mem3_reg[209][30]/P0001 ,
		_w13152_,
		_w14205_
	);
	LUT2 #(
		.INIT('h8)
	) name3694 (
		\wishbone_bd_ram_mem3_reg[4][30]/P0001 ,
		_w12666_,
		_w14206_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		\wishbone_bd_ram_mem3_reg[191][30]/P0001 ,
		_w13034_,
		_w14207_
	);
	LUT2 #(
		.INIT('h8)
	) name3696 (
		\wishbone_bd_ram_mem3_reg[228][30]/P0001 ,
		_w12765_,
		_w14208_
	);
	LUT2 #(
		.INIT('h8)
	) name3697 (
		\wishbone_bd_ram_mem3_reg[217][30]/P0001 ,
		_w13188_,
		_w14209_
	);
	LUT2 #(
		.INIT('h8)
	) name3698 (
		\wishbone_bd_ram_mem3_reg[62][30]/P0001 ,
		_w12673_,
		_w14210_
	);
	LUT2 #(
		.INIT('h8)
	) name3699 (
		\wishbone_bd_ram_mem3_reg[207][30]/P0001 ,
		_w13180_,
		_w14211_
	);
	LUT2 #(
		.INIT('h8)
	) name3700 (
		\wishbone_bd_ram_mem3_reg[16][30]/P0001 ,
		_w13140_,
		_w14212_
	);
	LUT2 #(
		.INIT('h8)
	) name3701 (
		\wishbone_bd_ram_mem3_reg[88][30]/P0001 ,
		_w12860_,
		_w14213_
	);
	LUT2 #(
		.INIT('h8)
	) name3702 (
		\wishbone_bd_ram_mem3_reg[41][30]/P0001 ,
		_w13052_,
		_w14214_
	);
	LUT2 #(
		.INIT('h8)
	) name3703 (
		\wishbone_bd_ram_mem3_reg[40][30]/P0001 ,
		_w13132_,
		_w14215_
	);
	LUT2 #(
		.INIT('h8)
	) name3704 (
		\wishbone_bd_ram_mem3_reg[94][30]/P0001 ,
		_w13186_,
		_w14216_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		\wishbone_bd_ram_mem3_reg[201][30]/P0001 ,
		_w12822_,
		_w14217_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		\wishbone_bd_ram_mem3_reg[167][30]/P0001 ,
		_w12986_,
		_w14218_
	);
	LUT2 #(
		.INIT('h8)
	) name3707 (
		\wishbone_bd_ram_mem3_reg[105][30]/P0001 ,
		_w12751_,
		_w14219_
	);
	LUT2 #(
		.INIT('h8)
	) name3708 (
		\wishbone_bd_ram_mem3_reg[111][30]/P0001 ,
		_w12744_,
		_w14220_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		\wishbone_bd_ram_mem3_reg[245][30]/P0001 ,
		_w13022_,
		_w14221_
	);
	LUT2 #(
		.INIT('h8)
	) name3710 (
		\wishbone_bd_ram_mem3_reg[17][30]/P0001 ,
		_w12848_,
		_w14222_
	);
	LUT2 #(
		.INIT('h8)
	) name3711 (
		\wishbone_bd_ram_mem3_reg[69][30]/P0001 ,
		_w12738_,
		_w14223_
	);
	LUT2 #(
		.INIT('h8)
	) name3712 (
		\wishbone_bd_ram_mem3_reg[160][30]/P0001 ,
		_w12872_,
		_w14224_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		\wishbone_bd_ram_mem3_reg[51][30]/P0001 ,
		_w13024_,
		_w14225_
	);
	LUT2 #(
		.INIT('h8)
	) name3714 (
		\wishbone_bd_ram_mem3_reg[81][30]/P0001 ,
		_w12950_,
		_w14226_
	);
	LUT2 #(
		.INIT('h8)
	) name3715 (
		\wishbone_bd_ram_mem3_reg[76][30]/P0001 ,
		_w13184_,
		_w14227_
	);
	LUT2 #(
		.INIT('h8)
	) name3716 (
		\wishbone_bd_ram_mem3_reg[159][30]/P0001 ,
		_w12774_,
		_w14228_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		\wishbone_bd_ram_mem3_reg[223][30]/P0001 ,
		_w12838_,
		_w14229_
	);
	LUT2 #(
		.INIT('h8)
	) name3718 (
		\wishbone_bd_ram_mem3_reg[30][30]/P0001 ,
		_w13104_,
		_w14230_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		\wishbone_bd_ram_mem3_reg[165][30]/P0001 ,
		_w13044_,
		_w14231_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		\wishbone_bd_ram_mem3_reg[70][30]/P0001 ,
		_w12840_,
		_w14232_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		\wishbone_bd_ram_mem3_reg[85][30]/P0001 ,
		_w13216_,
		_w14233_
	);
	LUT2 #(
		.INIT('h8)
	) name3722 (
		\wishbone_bd_ram_mem3_reg[2][30]/P0001 ,
		_w13088_,
		_w14234_
	);
	LUT2 #(
		.INIT('h8)
	) name3723 (
		\wishbone_bd_ram_mem3_reg[238][30]/P0001 ,
		_w13160_,
		_w14235_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		\wishbone_bd_ram_mem3_reg[218][30]/P0001 ,
		_w13206_,
		_w14236_
	);
	LUT2 #(
		.INIT('h8)
	) name3725 (
		\wishbone_bd_ram_mem3_reg[42][30]/P0001 ,
		_w12842_,
		_w14237_
	);
	LUT2 #(
		.INIT('h8)
	) name3726 (
		\wishbone_bd_ram_mem3_reg[128][30]/P0001 ,
		_w12793_,
		_w14238_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		\wishbone_bd_ram_mem3_reg[137][30]/P0001 ,
		_w13168_,
		_w14239_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		\wishbone_bd_ram_mem3_reg[251][30]/P0001 ,
		_w13054_,
		_w14240_
	);
	LUT2 #(
		.INIT('h8)
	) name3729 (
		\wishbone_bd_ram_mem3_reg[80][30]/P0001 ,
		_w12689_,
		_w14241_
	);
	LUT2 #(
		.INIT('h8)
	) name3730 (
		\wishbone_bd_ram_mem3_reg[231][30]/P0001 ,
		_w12856_,
		_w14242_
	);
	LUT2 #(
		.INIT('h8)
	) name3731 (
		\wishbone_bd_ram_mem3_reg[198][30]/P0001 ,
		_w12832_,
		_w14243_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		\wishbone_bd_ram_mem3_reg[25][30]/P0001 ,
		_w13108_,
		_w14244_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		\wishbone_bd_ram_mem3_reg[108][30]/P0001 ,
		_w13156_,
		_w14245_
	);
	LUT2 #(
		.INIT('h8)
	) name3734 (
		\wishbone_bd_ram_mem3_reg[21][30]/P0001 ,
		_w12906_,
		_w14246_
	);
	LUT2 #(
		.INIT('h8)
	) name3735 (
		\wishbone_bd_ram_mem3_reg[114][30]/P0001 ,
		_w13202_,
		_w14247_
	);
	LUT2 #(
		.INIT('h8)
	) name3736 (
		\wishbone_bd_ram_mem3_reg[155][30]/P0001 ,
		_w13122_,
		_w14248_
	);
	LUT2 #(
		.INIT('h8)
	) name3737 (
		\wishbone_bd_ram_mem3_reg[84][30]/P0001 ,
		_w12934_,
		_w14249_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		\wishbone_bd_ram_mem3_reg[244][30]/P0001 ,
		_w12747_,
		_w14250_
	);
	LUT2 #(
		.INIT('h8)
	) name3739 (
		\wishbone_bd_ram_mem3_reg[221][30]/P0001 ,
		_w12802_,
		_w14251_
	);
	LUT2 #(
		.INIT('h8)
	) name3740 (
		\wishbone_bd_ram_mem3_reg[203][30]/P0001 ,
		_w13158_,
		_w14252_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		\wishbone_bd_ram_mem3_reg[113][30]/P0001 ,
		_w13026_,
		_w14253_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		\wishbone_bd_ram_mem3_reg[197][30]/P0001 ,
		_w12834_,
		_w14254_
	);
	LUT2 #(
		.INIT('h8)
	) name3743 (
		\wishbone_bd_ram_mem3_reg[152][30]/P0001 ,
		_w12966_,
		_w14255_
	);
	LUT2 #(
		.INIT('h8)
	) name3744 (
		\wishbone_bd_ram_mem3_reg[22][30]/P0001 ,
		_w13110_,
		_w14256_
	);
	LUT2 #(
		.INIT('h8)
	) name3745 (
		\wishbone_bd_ram_mem3_reg[48][30]/P0001 ,
		_w12970_,
		_w14257_
	);
	LUT2 #(
		.INIT('h8)
	) name3746 (
		\wishbone_bd_ram_mem3_reg[52][30]/P0001 ,
		_w13082_,
		_w14258_
	);
	LUT2 #(
		.INIT('h8)
	) name3747 (
		\wishbone_bd_ram_mem3_reg[5][30]/P0001 ,
		_w12878_,
		_w14259_
	);
	LUT2 #(
		.INIT('h8)
	) name3748 (
		\wishbone_bd_ram_mem3_reg[78][30]/P0001 ,
		_w12874_,
		_w14260_
	);
	LUT2 #(
		.INIT('h8)
	) name3749 (
		\wishbone_bd_ram_mem3_reg[253][30]/P0001 ,
		_w13100_,
		_w14261_
	);
	LUT2 #(
		.INIT('h8)
	) name3750 (
		\wishbone_bd_ram_mem3_reg[79][30]/P0001 ,
		_w13212_,
		_w14262_
	);
	LUT2 #(
		.INIT('h8)
	) name3751 (
		\wishbone_bd_ram_mem3_reg[55][30]/P0001 ,
		_w12785_,
		_w14263_
	);
	LUT2 #(
		.INIT('h8)
	) name3752 (
		\wishbone_bd_ram_mem3_reg[222][30]/P0001 ,
		_w13094_,
		_w14264_
	);
	LUT2 #(
		.INIT('h8)
	) name3753 (
		\wishbone_bd_ram_mem3_reg[240][30]/P0001 ,
		_w12864_,
		_w14265_
	);
	LUT2 #(
		.INIT('h8)
	) name3754 (
		\wishbone_bd_ram_mem3_reg[151][30]/P0001 ,
		_w13142_,
		_w14266_
	);
	LUT2 #(
		.INIT('h8)
	) name3755 (
		\wishbone_bd_ram_mem3_reg[195][30]/P0001 ,
		_w13144_,
		_w14267_
	);
	LUT2 #(
		.INIT('h8)
	) name3756 (
		\wishbone_bd_ram_mem3_reg[46][30]/P0001 ,
		_w12884_,
		_w14268_
	);
	LUT2 #(
		.INIT('h8)
	) name3757 (
		\wishbone_bd_ram_mem3_reg[214][30]/P0001 ,
		_w12984_,
		_w14269_
	);
	LUT2 #(
		.INIT('h8)
	) name3758 (
		\wishbone_bd_ram_mem3_reg[172][30]/P0001 ,
		_w12944_,
		_w14270_
	);
	LUT2 #(
		.INIT('h8)
	) name3759 (
		\wishbone_bd_ram_mem3_reg[24][30]/P0001 ,
		_w13084_,
		_w14271_
	);
	LUT2 #(
		.INIT('h8)
	) name3760 (
		\wishbone_bd_ram_mem3_reg[170][30]/P0001 ,
		_w13030_,
		_w14272_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		\wishbone_bd_ram_mem3_reg[161][30]/P0001 ,
		_w12754_,
		_w14273_
	);
	LUT2 #(
		.INIT('h8)
	) name3762 (
		\wishbone_bd_ram_mem3_reg[99][30]/P0001 ,
		_w13038_,
		_w14274_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		\wishbone_bd_ram_mem3_reg[101][30]/P0001 ,
		_w13192_,
		_w14275_
	);
	LUT2 #(
		.INIT('h8)
	) name3764 (
		\wishbone_bd_ram_mem3_reg[233][30]/P0001 ,
		_w12836_,
		_w14276_
	);
	LUT2 #(
		.INIT('h8)
	) name3765 (
		\wishbone_bd_ram_mem3_reg[44][30]/P0001 ,
		_w12896_,
		_w14277_
	);
	LUT2 #(
		.INIT('h8)
	) name3766 (
		\wishbone_bd_ram_mem3_reg[133][30]/P0001 ,
		_w12761_,
		_w14278_
	);
	LUT2 #(
		.INIT('h8)
	) name3767 (
		\wishbone_bd_ram_mem3_reg[57][30]/P0001 ,
		_w13116_,
		_w14279_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		\wishbone_bd_ram_mem3_reg[106][30]/P0001 ,
		_w12713_,
		_w14280_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w14025_,
		_w14026_,
		_w14281_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		_w14027_,
		_w14028_,
		_w14282_
	);
	LUT2 #(
		.INIT('h1)
	) name3771 (
		_w14029_,
		_w14030_,
		_w14283_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w14031_,
		_w14032_,
		_w14284_
	);
	LUT2 #(
		.INIT('h1)
	) name3773 (
		_w14033_,
		_w14034_,
		_w14285_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w14035_,
		_w14036_,
		_w14286_
	);
	LUT2 #(
		.INIT('h1)
	) name3775 (
		_w14037_,
		_w14038_,
		_w14287_
	);
	LUT2 #(
		.INIT('h1)
	) name3776 (
		_w14039_,
		_w14040_,
		_w14288_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w14041_,
		_w14042_,
		_w14289_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w14043_,
		_w14044_,
		_w14290_
	);
	LUT2 #(
		.INIT('h1)
	) name3779 (
		_w14045_,
		_w14046_,
		_w14291_
	);
	LUT2 #(
		.INIT('h1)
	) name3780 (
		_w14047_,
		_w14048_,
		_w14292_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w14049_,
		_w14050_,
		_w14293_
	);
	LUT2 #(
		.INIT('h1)
	) name3782 (
		_w14051_,
		_w14052_,
		_w14294_
	);
	LUT2 #(
		.INIT('h1)
	) name3783 (
		_w14053_,
		_w14054_,
		_w14295_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		_w14055_,
		_w14056_,
		_w14296_
	);
	LUT2 #(
		.INIT('h1)
	) name3785 (
		_w14057_,
		_w14058_,
		_w14297_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w14059_,
		_w14060_,
		_w14298_
	);
	LUT2 #(
		.INIT('h1)
	) name3787 (
		_w14061_,
		_w14062_,
		_w14299_
	);
	LUT2 #(
		.INIT('h1)
	) name3788 (
		_w14063_,
		_w14064_,
		_w14300_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		_w14065_,
		_w14066_,
		_w14301_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w14067_,
		_w14068_,
		_w14302_
	);
	LUT2 #(
		.INIT('h1)
	) name3791 (
		_w14069_,
		_w14070_,
		_w14303_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		_w14071_,
		_w14072_,
		_w14304_
	);
	LUT2 #(
		.INIT('h1)
	) name3793 (
		_w14073_,
		_w14074_,
		_w14305_
	);
	LUT2 #(
		.INIT('h1)
	) name3794 (
		_w14075_,
		_w14076_,
		_w14306_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w14077_,
		_w14078_,
		_w14307_
	);
	LUT2 #(
		.INIT('h1)
	) name3796 (
		_w14079_,
		_w14080_,
		_w14308_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w14081_,
		_w14082_,
		_w14309_
	);
	LUT2 #(
		.INIT('h1)
	) name3798 (
		_w14083_,
		_w14084_,
		_w14310_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		_w14085_,
		_w14086_,
		_w14311_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		_w14087_,
		_w14088_,
		_w14312_
	);
	LUT2 #(
		.INIT('h1)
	) name3801 (
		_w14089_,
		_w14090_,
		_w14313_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w14091_,
		_w14092_,
		_w14314_
	);
	LUT2 #(
		.INIT('h1)
	) name3803 (
		_w14093_,
		_w14094_,
		_w14315_
	);
	LUT2 #(
		.INIT('h1)
	) name3804 (
		_w14095_,
		_w14096_,
		_w14316_
	);
	LUT2 #(
		.INIT('h1)
	) name3805 (
		_w14097_,
		_w14098_,
		_w14317_
	);
	LUT2 #(
		.INIT('h1)
	) name3806 (
		_w14099_,
		_w14100_,
		_w14318_
	);
	LUT2 #(
		.INIT('h1)
	) name3807 (
		_w14101_,
		_w14102_,
		_w14319_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		_w14103_,
		_w14104_,
		_w14320_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w14105_,
		_w14106_,
		_w14321_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		_w14107_,
		_w14108_,
		_w14322_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w14109_,
		_w14110_,
		_w14323_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w14111_,
		_w14112_,
		_w14324_
	);
	LUT2 #(
		.INIT('h1)
	) name3813 (
		_w14113_,
		_w14114_,
		_w14325_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		_w14115_,
		_w14116_,
		_w14326_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w14117_,
		_w14118_,
		_w14327_
	);
	LUT2 #(
		.INIT('h1)
	) name3816 (
		_w14119_,
		_w14120_,
		_w14328_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w14121_,
		_w14122_,
		_w14329_
	);
	LUT2 #(
		.INIT('h1)
	) name3818 (
		_w14123_,
		_w14124_,
		_w14330_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w14125_,
		_w14126_,
		_w14331_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w14127_,
		_w14128_,
		_w14332_
	);
	LUT2 #(
		.INIT('h1)
	) name3821 (
		_w14129_,
		_w14130_,
		_w14333_
	);
	LUT2 #(
		.INIT('h1)
	) name3822 (
		_w14131_,
		_w14132_,
		_w14334_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		_w14133_,
		_w14134_,
		_w14335_
	);
	LUT2 #(
		.INIT('h1)
	) name3824 (
		_w14135_,
		_w14136_,
		_w14336_
	);
	LUT2 #(
		.INIT('h1)
	) name3825 (
		_w14137_,
		_w14138_,
		_w14337_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w14139_,
		_w14140_,
		_w14338_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w14141_,
		_w14142_,
		_w14339_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		_w14143_,
		_w14144_,
		_w14340_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w14145_,
		_w14146_,
		_w14341_
	);
	LUT2 #(
		.INIT('h1)
	) name3830 (
		_w14147_,
		_w14148_,
		_w14342_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w14149_,
		_w14150_,
		_w14343_
	);
	LUT2 #(
		.INIT('h1)
	) name3832 (
		_w14151_,
		_w14152_,
		_w14344_
	);
	LUT2 #(
		.INIT('h1)
	) name3833 (
		_w14153_,
		_w14154_,
		_w14345_
	);
	LUT2 #(
		.INIT('h1)
	) name3834 (
		_w14155_,
		_w14156_,
		_w14346_
	);
	LUT2 #(
		.INIT('h1)
	) name3835 (
		_w14157_,
		_w14158_,
		_w14347_
	);
	LUT2 #(
		.INIT('h1)
	) name3836 (
		_w14159_,
		_w14160_,
		_w14348_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w14161_,
		_w14162_,
		_w14349_
	);
	LUT2 #(
		.INIT('h1)
	) name3838 (
		_w14163_,
		_w14164_,
		_w14350_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w14165_,
		_w14166_,
		_w14351_
	);
	LUT2 #(
		.INIT('h1)
	) name3840 (
		_w14167_,
		_w14168_,
		_w14352_
	);
	LUT2 #(
		.INIT('h1)
	) name3841 (
		_w14169_,
		_w14170_,
		_w14353_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w14171_,
		_w14172_,
		_w14354_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w14173_,
		_w14174_,
		_w14355_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		_w14175_,
		_w14176_,
		_w14356_
	);
	LUT2 #(
		.INIT('h1)
	) name3845 (
		_w14177_,
		_w14178_,
		_w14357_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w14179_,
		_w14180_,
		_w14358_
	);
	LUT2 #(
		.INIT('h1)
	) name3847 (
		_w14181_,
		_w14182_,
		_w14359_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w14183_,
		_w14184_,
		_w14360_
	);
	LUT2 #(
		.INIT('h1)
	) name3849 (
		_w14185_,
		_w14186_,
		_w14361_
	);
	LUT2 #(
		.INIT('h1)
	) name3850 (
		_w14187_,
		_w14188_,
		_w14362_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w14189_,
		_w14190_,
		_w14363_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w14191_,
		_w14192_,
		_w14364_
	);
	LUT2 #(
		.INIT('h1)
	) name3853 (
		_w14193_,
		_w14194_,
		_w14365_
	);
	LUT2 #(
		.INIT('h1)
	) name3854 (
		_w14195_,
		_w14196_,
		_w14366_
	);
	LUT2 #(
		.INIT('h1)
	) name3855 (
		_w14197_,
		_w14198_,
		_w14367_
	);
	LUT2 #(
		.INIT('h1)
	) name3856 (
		_w14199_,
		_w14200_,
		_w14368_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w14201_,
		_w14202_,
		_w14369_
	);
	LUT2 #(
		.INIT('h1)
	) name3858 (
		_w14203_,
		_w14204_,
		_w14370_
	);
	LUT2 #(
		.INIT('h1)
	) name3859 (
		_w14205_,
		_w14206_,
		_w14371_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		_w14207_,
		_w14208_,
		_w14372_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w14209_,
		_w14210_,
		_w14373_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w14211_,
		_w14212_,
		_w14374_
	);
	LUT2 #(
		.INIT('h1)
	) name3863 (
		_w14213_,
		_w14214_,
		_w14375_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w14215_,
		_w14216_,
		_w14376_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w14217_,
		_w14218_,
		_w14377_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		_w14219_,
		_w14220_,
		_w14378_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w14221_,
		_w14222_,
		_w14379_
	);
	LUT2 #(
		.INIT('h1)
	) name3868 (
		_w14223_,
		_w14224_,
		_w14380_
	);
	LUT2 #(
		.INIT('h1)
	) name3869 (
		_w14225_,
		_w14226_,
		_w14381_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w14227_,
		_w14228_,
		_w14382_
	);
	LUT2 #(
		.INIT('h1)
	) name3871 (
		_w14229_,
		_w14230_,
		_w14383_
	);
	LUT2 #(
		.INIT('h1)
	) name3872 (
		_w14231_,
		_w14232_,
		_w14384_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w14233_,
		_w14234_,
		_w14385_
	);
	LUT2 #(
		.INIT('h1)
	) name3874 (
		_w14235_,
		_w14236_,
		_w14386_
	);
	LUT2 #(
		.INIT('h1)
	) name3875 (
		_w14237_,
		_w14238_,
		_w14387_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		_w14239_,
		_w14240_,
		_w14388_
	);
	LUT2 #(
		.INIT('h1)
	) name3877 (
		_w14241_,
		_w14242_,
		_w14389_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w14243_,
		_w14244_,
		_w14390_
	);
	LUT2 #(
		.INIT('h1)
	) name3879 (
		_w14245_,
		_w14246_,
		_w14391_
	);
	LUT2 #(
		.INIT('h1)
	) name3880 (
		_w14247_,
		_w14248_,
		_w14392_
	);
	LUT2 #(
		.INIT('h1)
	) name3881 (
		_w14249_,
		_w14250_,
		_w14393_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		_w14251_,
		_w14252_,
		_w14394_
	);
	LUT2 #(
		.INIT('h1)
	) name3883 (
		_w14253_,
		_w14254_,
		_w14395_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w14255_,
		_w14256_,
		_w14396_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w14257_,
		_w14258_,
		_w14397_
	);
	LUT2 #(
		.INIT('h1)
	) name3886 (
		_w14259_,
		_w14260_,
		_w14398_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w14261_,
		_w14262_,
		_w14399_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		_w14263_,
		_w14264_,
		_w14400_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w14265_,
		_w14266_,
		_w14401_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		_w14267_,
		_w14268_,
		_w14402_
	);
	LUT2 #(
		.INIT('h1)
	) name3891 (
		_w14269_,
		_w14270_,
		_w14403_
	);
	LUT2 #(
		.INIT('h1)
	) name3892 (
		_w14271_,
		_w14272_,
		_w14404_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w14273_,
		_w14274_,
		_w14405_
	);
	LUT2 #(
		.INIT('h1)
	) name3894 (
		_w14275_,
		_w14276_,
		_w14406_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w14277_,
		_w14278_,
		_w14407_
	);
	LUT2 #(
		.INIT('h1)
	) name3896 (
		_w14279_,
		_w14280_,
		_w14408_
	);
	LUT2 #(
		.INIT('h8)
	) name3897 (
		_w14407_,
		_w14408_,
		_w14409_
	);
	LUT2 #(
		.INIT('h8)
	) name3898 (
		_w14405_,
		_w14406_,
		_w14410_
	);
	LUT2 #(
		.INIT('h8)
	) name3899 (
		_w14403_,
		_w14404_,
		_w14411_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		_w14401_,
		_w14402_,
		_w14412_
	);
	LUT2 #(
		.INIT('h8)
	) name3901 (
		_w14399_,
		_w14400_,
		_w14413_
	);
	LUT2 #(
		.INIT('h8)
	) name3902 (
		_w14397_,
		_w14398_,
		_w14414_
	);
	LUT2 #(
		.INIT('h8)
	) name3903 (
		_w14395_,
		_w14396_,
		_w14415_
	);
	LUT2 #(
		.INIT('h8)
	) name3904 (
		_w14393_,
		_w14394_,
		_w14416_
	);
	LUT2 #(
		.INIT('h8)
	) name3905 (
		_w14391_,
		_w14392_,
		_w14417_
	);
	LUT2 #(
		.INIT('h8)
	) name3906 (
		_w14389_,
		_w14390_,
		_w14418_
	);
	LUT2 #(
		.INIT('h8)
	) name3907 (
		_w14387_,
		_w14388_,
		_w14419_
	);
	LUT2 #(
		.INIT('h8)
	) name3908 (
		_w14385_,
		_w14386_,
		_w14420_
	);
	LUT2 #(
		.INIT('h8)
	) name3909 (
		_w14383_,
		_w14384_,
		_w14421_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		_w14381_,
		_w14382_,
		_w14422_
	);
	LUT2 #(
		.INIT('h8)
	) name3911 (
		_w14379_,
		_w14380_,
		_w14423_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		_w14377_,
		_w14378_,
		_w14424_
	);
	LUT2 #(
		.INIT('h8)
	) name3913 (
		_w14375_,
		_w14376_,
		_w14425_
	);
	LUT2 #(
		.INIT('h8)
	) name3914 (
		_w14373_,
		_w14374_,
		_w14426_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		_w14371_,
		_w14372_,
		_w14427_
	);
	LUT2 #(
		.INIT('h8)
	) name3916 (
		_w14369_,
		_w14370_,
		_w14428_
	);
	LUT2 #(
		.INIT('h8)
	) name3917 (
		_w14367_,
		_w14368_,
		_w14429_
	);
	LUT2 #(
		.INIT('h8)
	) name3918 (
		_w14365_,
		_w14366_,
		_w14430_
	);
	LUT2 #(
		.INIT('h8)
	) name3919 (
		_w14363_,
		_w14364_,
		_w14431_
	);
	LUT2 #(
		.INIT('h8)
	) name3920 (
		_w14361_,
		_w14362_,
		_w14432_
	);
	LUT2 #(
		.INIT('h8)
	) name3921 (
		_w14359_,
		_w14360_,
		_w14433_
	);
	LUT2 #(
		.INIT('h8)
	) name3922 (
		_w14357_,
		_w14358_,
		_w14434_
	);
	LUT2 #(
		.INIT('h8)
	) name3923 (
		_w14355_,
		_w14356_,
		_w14435_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		_w14353_,
		_w14354_,
		_w14436_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		_w14351_,
		_w14352_,
		_w14437_
	);
	LUT2 #(
		.INIT('h8)
	) name3926 (
		_w14349_,
		_w14350_,
		_w14438_
	);
	LUT2 #(
		.INIT('h8)
	) name3927 (
		_w14347_,
		_w14348_,
		_w14439_
	);
	LUT2 #(
		.INIT('h8)
	) name3928 (
		_w14345_,
		_w14346_,
		_w14440_
	);
	LUT2 #(
		.INIT('h8)
	) name3929 (
		_w14343_,
		_w14344_,
		_w14441_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w14341_,
		_w14342_,
		_w14442_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		_w14339_,
		_w14340_,
		_w14443_
	);
	LUT2 #(
		.INIT('h8)
	) name3932 (
		_w14337_,
		_w14338_,
		_w14444_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		_w14335_,
		_w14336_,
		_w14445_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w14333_,
		_w14334_,
		_w14446_
	);
	LUT2 #(
		.INIT('h8)
	) name3935 (
		_w14331_,
		_w14332_,
		_w14447_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w14329_,
		_w14330_,
		_w14448_
	);
	LUT2 #(
		.INIT('h8)
	) name3937 (
		_w14327_,
		_w14328_,
		_w14449_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w14325_,
		_w14326_,
		_w14450_
	);
	LUT2 #(
		.INIT('h8)
	) name3939 (
		_w14323_,
		_w14324_,
		_w14451_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w14321_,
		_w14322_,
		_w14452_
	);
	LUT2 #(
		.INIT('h8)
	) name3941 (
		_w14319_,
		_w14320_,
		_w14453_
	);
	LUT2 #(
		.INIT('h8)
	) name3942 (
		_w14317_,
		_w14318_,
		_w14454_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		_w14315_,
		_w14316_,
		_w14455_
	);
	LUT2 #(
		.INIT('h8)
	) name3944 (
		_w14313_,
		_w14314_,
		_w14456_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w14311_,
		_w14312_,
		_w14457_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		_w14309_,
		_w14310_,
		_w14458_
	);
	LUT2 #(
		.INIT('h8)
	) name3947 (
		_w14307_,
		_w14308_,
		_w14459_
	);
	LUT2 #(
		.INIT('h8)
	) name3948 (
		_w14305_,
		_w14306_,
		_w14460_
	);
	LUT2 #(
		.INIT('h8)
	) name3949 (
		_w14303_,
		_w14304_,
		_w14461_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w14301_,
		_w14302_,
		_w14462_
	);
	LUT2 #(
		.INIT('h8)
	) name3951 (
		_w14299_,
		_w14300_,
		_w14463_
	);
	LUT2 #(
		.INIT('h8)
	) name3952 (
		_w14297_,
		_w14298_,
		_w14464_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		_w14295_,
		_w14296_,
		_w14465_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		_w14293_,
		_w14294_,
		_w14466_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w14291_,
		_w14292_,
		_w14467_
	);
	LUT2 #(
		.INIT('h8)
	) name3956 (
		_w14289_,
		_w14290_,
		_w14468_
	);
	LUT2 #(
		.INIT('h8)
	) name3957 (
		_w14287_,
		_w14288_,
		_w14469_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		_w14285_,
		_w14286_,
		_w14470_
	);
	LUT2 #(
		.INIT('h8)
	) name3959 (
		_w14283_,
		_w14284_,
		_w14471_
	);
	LUT2 #(
		.INIT('h8)
	) name3960 (
		_w14281_,
		_w14282_,
		_w14472_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		_w14471_,
		_w14472_,
		_w14473_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		_w14469_,
		_w14470_,
		_w14474_
	);
	LUT2 #(
		.INIT('h8)
	) name3963 (
		_w14467_,
		_w14468_,
		_w14475_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		_w14465_,
		_w14466_,
		_w14476_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		_w14463_,
		_w14464_,
		_w14477_
	);
	LUT2 #(
		.INIT('h8)
	) name3966 (
		_w14461_,
		_w14462_,
		_w14478_
	);
	LUT2 #(
		.INIT('h8)
	) name3967 (
		_w14459_,
		_w14460_,
		_w14479_
	);
	LUT2 #(
		.INIT('h8)
	) name3968 (
		_w14457_,
		_w14458_,
		_w14480_
	);
	LUT2 #(
		.INIT('h8)
	) name3969 (
		_w14455_,
		_w14456_,
		_w14481_
	);
	LUT2 #(
		.INIT('h8)
	) name3970 (
		_w14453_,
		_w14454_,
		_w14482_
	);
	LUT2 #(
		.INIT('h8)
	) name3971 (
		_w14451_,
		_w14452_,
		_w14483_
	);
	LUT2 #(
		.INIT('h8)
	) name3972 (
		_w14449_,
		_w14450_,
		_w14484_
	);
	LUT2 #(
		.INIT('h8)
	) name3973 (
		_w14447_,
		_w14448_,
		_w14485_
	);
	LUT2 #(
		.INIT('h8)
	) name3974 (
		_w14445_,
		_w14446_,
		_w14486_
	);
	LUT2 #(
		.INIT('h8)
	) name3975 (
		_w14443_,
		_w14444_,
		_w14487_
	);
	LUT2 #(
		.INIT('h8)
	) name3976 (
		_w14441_,
		_w14442_,
		_w14488_
	);
	LUT2 #(
		.INIT('h8)
	) name3977 (
		_w14439_,
		_w14440_,
		_w14489_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		_w14437_,
		_w14438_,
		_w14490_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		_w14435_,
		_w14436_,
		_w14491_
	);
	LUT2 #(
		.INIT('h8)
	) name3980 (
		_w14433_,
		_w14434_,
		_w14492_
	);
	LUT2 #(
		.INIT('h8)
	) name3981 (
		_w14431_,
		_w14432_,
		_w14493_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		_w14429_,
		_w14430_,
		_w14494_
	);
	LUT2 #(
		.INIT('h8)
	) name3983 (
		_w14427_,
		_w14428_,
		_w14495_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		_w14425_,
		_w14426_,
		_w14496_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		_w14423_,
		_w14424_,
		_w14497_
	);
	LUT2 #(
		.INIT('h8)
	) name3986 (
		_w14421_,
		_w14422_,
		_w14498_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		_w14419_,
		_w14420_,
		_w14499_
	);
	LUT2 #(
		.INIT('h8)
	) name3988 (
		_w14417_,
		_w14418_,
		_w14500_
	);
	LUT2 #(
		.INIT('h8)
	) name3989 (
		_w14415_,
		_w14416_,
		_w14501_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		_w14413_,
		_w14414_,
		_w14502_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		_w14411_,
		_w14412_,
		_w14503_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		_w14409_,
		_w14410_,
		_w14504_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		_w14503_,
		_w14504_,
		_w14505_
	);
	LUT2 #(
		.INIT('h8)
	) name3994 (
		_w14501_,
		_w14502_,
		_w14506_
	);
	LUT2 #(
		.INIT('h8)
	) name3995 (
		_w14499_,
		_w14500_,
		_w14507_
	);
	LUT2 #(
		.INIT('h8)
	) name3996 (
		_w14497_,
		_w14498_,
		_w14508_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		_w14495_,
		_w14496_,
		_w14509_
	);
	LUT2 #(
		.INIT('h8)
	) name3998 (
		_w14493_,
		_w14494_,
		_w14510_
	);
	LUT2 #(
		.INIT('h8)
	) name3999 (
		_w14491_,
		_w14492_,
		_w14511_
	);
	LUT2 #(
		.INIT('h8)
	) name4000 (
		_w14489_,
		_w14490_,
		_w14512_
	);
	LUT2 #(
		.INIT('h8)
	) name4001 (
		_w14487_,
		_w14488_,
		_w14513_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		_w14485_,
		_w14486_,
		_w14514_
	);
	LUT2 #(
		.INIT('h8)
	) name4003 (
		_w14483_,
		_w14484_,
		_w14515_
	);
	LUT2 #(
		.INIT('h8)
	) name4004 (
		_w14481_,
		_w14482_,
		_w14516_
	);
	LUT2 #(
		.INIT('h8)
	) name4005 (
		_w14479_,
		_w14480_,
		_w14517_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w14477_,
		_w14478_,
		_w14518_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		_w14475_,
		_w14476_,
		_w14519_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		_w14473_,
		_w14474_,
		_w14520_
	);
	LUT2 #(
		.INIT('h8)
	) name4009 (
		_w14519_,
		_w14520_,
		_w14521_
	);
	LUT2 #(
		.INIT('h8)
	) name4010 (
		_w14517_,
		_w14518_,
		_w14522_
	);
	LUT2 #(
		.INIT('h8)
	) name4011 (
		_w14515_,
		_w14516_,
		_w14523_
	);
	LUT2 #(
		.INIT('h8)
	) name4012 (
		_w14513_,
		_w14514_,
		_w14524_
	);
	LUT2 #(
		.INIT('h8)
	) name4013 (
		_w14511_,
		_w14512_,
		_w14525_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		_w14509_,
		_w14510_,
		_w14526_
	);
	LUT2 #(
		.INIT('h8)
	) name4015 (
		_w14507_,
		_w14508_,
		_w14527_
	);
	LUT2 #(
		.INIT('h8)
	) name4016 (
		_w14505_,
		_w14506_,
		_w14528_
	);
	LUT2 #(
		.INIT('h8)
	) name4017 (
		_w14527_,
		_w14528_,
		_w14529_
	);
	LUT2 #(
		.INIT('h8)
	) name4018 (
		_w14525_,
		_w14526_,
		_w14530_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w14523_,
		_w14524_,
		_w14531_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		_w14521_,
		_w14522_,
		_w14532_
	);
	LUT2 #(
		.INIT('h8)
	) name4021 (
		_w14531_,
		_w14532_,
		_w14533_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		_w14529_,
		_w14530_,
		_w14534_
	);
	LUT2 #(
		.INIT('h8)
	) name4023 (
		_w14533_,
		_w14534_,
		_w14535_
	);
	LUT2 #(
		.INIT('h1)
	) name4024 (
		wb_rst_i_pad,
		_w14535_,
		_w14536_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		_w12656_,
		_w14536_,
		_w14537_
	);
	LUT2 #(
		.INIT('h2)
	) name4026 (
		_w13501_,
		_w14021_,
		_w14538_
	);
	LUT2 #(
		.INIT('h1)
	) name4027 (
		_w12658_,
		_w14538_,
		_w14539_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		\wishbone_TxLength_reg[14]/NET0131 ,
		_w14539_,
		_w14540_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		\wishbone_TxLength_reg[14]/NET0131 ,
		_w14022_,
		_w14541_
	);
	LUT2 #(
		.INIT('h1)
	) name4030 (
		_w14540_,
		_w14541_,
		_w14542_
	);
	LUT2 #(
		.INIT('h4)
	) name4031 (
		_w14537_,
		_w14542_,
		_w14543_
	);
	LUT2 #(
		.INIT('h2)
	) name4032 (
		\rxethmac1_crcrx_Crc_reg[6]/NET0131 ,
		_w12115_,
		_w14544_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		\rxethmac1_crcrx_Crc_reg[6]/NET0131 ,
		_w12115_,
		_w14545_
	);
	LUT2 #(
		.INIT('h2)
	) name4034 (
		_w10580_,
		_w14544_,
		_w14546_
	);
	LUT2 #(
		.INIT('h4)
	) name4035 (
		_w14545_,
		_w14546_,
		_w14547_
	);
	LUT2 #(
		.INIT('h2)
	) name4036 (
		\rxethmac1_crcrx_Crc_reg[0]/NET0131 ,
		_w12115_,
		_w14548_
	);
	LUT2 #(
		.INIT('h4)
	) name4037 (
		\rxethmac1_crcrx_Crc_reg[0]/NET0131 ,
		_w12115_,
		_w14549_
	);
	LUT2 #(
		.INIT('h2)
	) name4038 (
		_w10580_,
		_w14548_,
		_w14550_
	);
	LUT2 #(
		.INIT('h4)
	) name4039 (
		_w14549_,
		_w14550_,
		_w14551_
	);
	LUT2 #(
		.INIT('h8)
	) name4040 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w14552_
	);
	LUT2 #(
		.INIT('h8)
	) name4041 (
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w14552_,
		_w14553_
	);
	LUT2 #(
		.INIT('h8)
	) name4042 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w14554_
	);
	LUT2 #(
		.INIT('h8)
	) name4043 (
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w14555_
	);
	LUT2 #(
		.INIT('h8)
	) name4044 (
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w14555_,
		_w14556_
	);
	LUT2 #(
		.INIT('h8)
	) name4045 (
		_w14554_,
		_w14556_,
		_w14557_
	);
	LUT2 #(
		.INIT('h2)
	) name4046 (
		\txethmac1_txcounters1_NibCnt_reg[0]/NET0131 ,
		_w11069_,
		_w14558_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w14558_,
		_w14559_
	);
	LUT2 #(
		.INIT('h8)
	) name4048 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w14560_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w14561_
	);
	LUT2 #(
		.INIT('h8)
	) name4050 (
		_w14560_,
		_w14561_,
		_w14562_
	);
	LUT2 #(
		.INIT('h8)
	) name4051 (
		_w14557_,
		_w14562_,
		_w14563_
	);
	LUT2 #(
		.INIT('h8)
	) name4052 (
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w14563_,
		_w14564_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w14565_
	);
	LUT2 #(
		.INIT('h8)
	) name4054 (
		_w14564_,
		_w14565_,
		_w14566_
	);
	LUT2 #(
		.INIT('h8)
	) name4055 (
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w14553_,
		_w14567_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		_w14566_,
		_w14567_,
		_w14568_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w14559_,
		_w14568_,
		_w14569_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w11021_,
		_w14569_,
		_w14570_
	);
	LUT2 #(
		.INIT('h2)
	) name4059 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w14570_,
		_w14571_
	);
	LUT2 #(
		.INIT('h8)
	) name4060 (
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w14571_,
		_w14572_
	);
	LUT2 #(
		.INIT('h8)
	) name4061 (
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w14573_,
		_w14574_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		_w14557_,
		_w14574_,
		_w14575_
	);
	LUT2 #(
		.INIT('h8)
	) name4064 (
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w14575_,
		_w14576_
	);
	LUT2 #(
		.INIT('h8)
	) name4065 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		_w14576_,
		_w14577_
	);
	LUT2 #(
		.INIT('h8)
	) name4066 (
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w14577_,
		_w14578_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		_w14553_,
		_w14578_,
		_w14579_
	);
	LUT2 #(
		.INIT('h1)
	) name4068 (
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w14579_,
		_w14580_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		_w11221_,
		_w14581_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		_w11254_,
		_w14581_,
		_w14582_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		\txethmac1_txcounters1_ByteCnt_reg[15]/NET0131 ,
		_w14579_,
		_w14583_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		_w14580_,
		_w14582_,
		_w14584_
	);
	LUT2 #(
		.INIT('h4)
	) name4073 (
		_w14583_,
		_w14584_,
		_w14585_
	);
	LUT2 #(
		.INIT('h8)
	) name4074 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w12577_,
		_w14586_
	);
	LUT2 #(
		.INIT('h4)
	) name4075 (
		\m_wb_adr_o[2]_pad ,
		_w12621_,
		_w14587_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		_w12634_,
		_w14587_,
		_w14588_
	);
	LUT2 #(
		.INIT('h2)
	) name4077 (
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		_w14588_,
		_w14589_
	);
	LUT2 #(
		.INIT('h4)
	) name4078 (
		_w12608_,
		_w12621_,
		_w14590_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		_w12623_,
		_w14590_,
		_w14591_
	);
	LUT2 #(
		.INIT('h8)
	) name4080 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w12561_,
		_w14592_
	);
	LUT2 #(
		.INIT('h2)
	) name4081 (
		_w14591_,
		_w14592_,
		_w14593_
	);
	LUT2 #(
		.INIT('h1)
	) name4082 (
		\m_wb_adr_o[2]_pad ,
		_w14593_,
		_w14594_
	);
	LUT2 #(
		.INIT('h8)
	) name4083 (
		\m_wb_adr_o[2]_pad ,
		_w12636_,
		_w14595_
	);
	LUT2 #(
		.INIT('h1)
	) name4084 (
		_w14586_,
		_w14589_,
		_w14596_
	);
	LUT2 #(
		.INIT('h4)
	) name4085 (
		_w14595_,
		_w14596_,
		_w14597_
	);
	LUT2 #(
		.INIT('h4)
	) name4086 (
		_w14594_,
		_w14597_,
		_w14598_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		\wishbone_bd_ram_mem3_reg[78][24]/P0001 ,
		_w12874_,
		_w14599_
	);
	LUT2 #(
		.INIT('h8)
	) name4088 (
		\wishbone_bd_ram_mem3_reg[157][24]/P0001 ,
		_w12926_,
		_w14600_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		\wishbone_bd_ram_mem3_reg[17][24]/P0001 ,
		_w12848_,
		_w14601_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		\wishbone_bd_ram_mem3_reg[0][24]/P0001 ,
		_w12717_,
		_w14602_
	);
	LUT2 #(
		.INIT('h8)
	) name4091 (
		\wishbone_bd_ram_mem3_reg[3][24]/P0001 ,
		_w12866_,
		_w14603_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		\wishbone_bd_ram_mem3_reg[126][24]/P0001 ,
		_w13218_,
		_w14604_
	);
	LUT2 #(
		.INIT('h8)
	) name4093 (
		\wishbone_bd_ram_mem3_reg[34][24]/P0001 ,
		_w12930_,
		_w14605_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		\wishbone_bd_ram_mem3_reg[55][24]/P0001 ,
		_w12785_,
		_w14606_
	);
	LUT2 #(
		.INIT('h8)
	) name4095 (
		\wishbone_bd_ram_mem3_reg[104][24]/P0001 ,
		_w13148_,
		_w14607_
	);
	LUT2 #(
		.INIT('h8)
	) name4096 (
		\wishbone_bd_ram_mem3_reg[252][24]/P0001 ,
		_w13080_,
		_w14608_
	);
	LUT2 #(
		.INIT('h8)
	) name4097 (
		\wishbone_bd_ram_mem3_reg[197][24]/P0001 ,
		_w12834_,
		_w14609_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		\wishbone_bd_ram_mem3_reg[137][24]/P0001 ,
		_w13168_,
		_w14610_
	);
	LUT2 #(
		.INIT('h8)
	) name4099 (
		\wishbone_bd_ram_mem3_reg[144][24]/P0001 ,
		_w12756_,
		_w14611_
	);
	LUT2 #(
		.INIT('h8)
	) name4100 (
		\wishbone_bd_ram_mem3_reg[227][24]/P0001 ,
		_w12936_,
		_w14612_
	);
	LUT2 #(
		.INIT('h8)
	) name4101 (
		\wishbone_bd_ram_mem3_reg[57][24]/P0001 ,
		_w13116_,
		_w14613_
	);
	LUT2 #(
		.INIT('h8)
	) name4102 (
		\wishbone_bd_ram_mem3_reg[188][24]/P0001 ,
		_w12948_,
		_w14614_
	);
	LUT2 #(
		.INIT('h8)
	) name4103 (
		\wishbone_bd_ram_mem3_reg[205][24]/P0001 ,
		_w13068_,
		_w14615_
	);
	LUT2 #(
		.INIT('h8)
	) name4104 (
		\wishbone_bd_ram_mem3_reg[176][24]/P0001 ,
		_w12868_,
		_w14616_
	);
	LUT2 #(
		.INIT('h8)
	) name4105 (
		\wishbone_bd_ram_mem3_reg[131][24]/P0001 ,
		_w12852_,
		_w14617_
	);
	LUT2 #(
		.INIT('h8)
	) name4106 (
		\wishbone_bd_ram_mem3_reg[39][24]/P0001 ,
		_w13018_,
		_w14618_
	);
	LUT2 #(
		.INIT('h8)
	) name4107 (
		\wishbone_bd_ram_mem3_reg[201][24]/P0001 ,
		_w12822_,
		_w14619_
	);
	LUT2 #(
		.INIT('h8)
	) name4108 (
		\wishbone_bd_ram_mem3_reg[91][24]/P0001 ,
		_w13074_,
		_w14620_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		\wishbone_bd_ram_mem3_reg[211][24]/P0001 ,
		_w13166_,
		_w14621_
	);
	LUT2 #(
		.INIT('h8)
	) name4110 (
		\wishbone_bd_ram_mem3_reg[149][24]/P0001 ,
		_w12741_,
		_w14622_
	);
	LUT2 #(
		.INIT('h8)
	) name4111 (
		\wishbone_bd_ram_mem3_reg[196][24]/P0001 ,
		_w13090_,
		_w14623_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		\wishbone_bd_ram_mem3_reg[84][24]/P0001 ,
		_w12934_,
		_w14624_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		\wishbone_bd_ram_mem3_reg[121][24]/P0001 ,
		_w13078_,
		_w14625_
	);
	LUT2 #(
		.INIT('h8)
	) name4114 (
		\wishbone_bd_ram_mem3_reg[83][24]/P0001 ,
		_w12916_,
		_w14626_
	);
	LUT2 #(
		.INIT('h8)
	) name4115 (
		\wishbone_bd_ram_mem3_reg[35][24]/P0001 ,
		_w12703_,
		_w14627_
	);
	LUT2 #(
		.INIT('h8)
	) name4116 (
		\wishbone_bd_ram_mem3_reg[218][24]/P0001 ,
		_w13206_,
		_w14628_
	);
	LUT2 #(
		.INIT('h8)
	) name4117 (
		\wishbone_bd_ram_mem3_reg[241][24]/P0001 ,
		_w13006_,
		_w14629_
	);
	LUT2 #(
		.INIT('h8)
	) name4118 (
		\wishbone_bd_ram_mem3_reg[170][24]/P0001 ,
		_w13030_,
		_w14630_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\wishbone_bd_ram_mem3_reg[100][24]/P0001 ,
		_w12960_,
		_w14631_
	);
	LUT2 #(
		.INIT('h8)
	) name4120 (
		\wishbone_bd_ram_mem3_reg[229][24]/P0001 ,
		_w12711_,
		_w14632_
	);
	LUT2 #(
		.INIT('h8)
	) name4121 (
		\wishbone_bd_ram_mem3_reg[110][24]/P0001 ,
		_w13046_,
		_w14633_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		\wishbone_bd_ram_mem3_reg[99][24]/P0001 ,
		_w13038_,
		_w14634_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		\wishbone_bd_ram_mem3_reg[130][24]/P0001 ,
		_w12914_,
		_w14635_
	);
	LUT2 #(
		.INIT('h8)
	) name4124 (
		\wishbone_bd_ram_mem3_reg[133][24]/P0001 ,
		_w12761_,
		_w14636_
	);
	LUT2 #(
		.INIT('h8)
	) name4125 (
		\wishbone_bd_ram_mem3_reg[152][24]/P0001 ,
		_w12966_,
		_w14637_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		\wishbone_bd_ram_mem3_reg[25][24]/P0001 ,
		_w13108_,
		_w14638_
	);
	LUT2 #(
		.INIT('h8)
	) name4127 (
		\wishbone_bd_ram_mem3_reg[220][24]/P0001 ,
		_w13066_,
		_w14639_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		\wishbone_bd_ram_mem3_reg[245][24]/P0001 ,
		_w13022_,
		_w14640_
	);
	LUT2 #(
		.INIT('h8)
	) name4129 (
		\wishbone_bd_ram_mem3_reg[33][24]/P0001 ,
		_w12980_,
		_w14641_
	);
	LUT2 #(
		.INIT('h8)
	) name4130 (
		\wishbone_bd_ram_mem3_reg[61][24]/P0001 ,
		_w12725_,
		_w14642_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		\wishbone_bd_ram_mem3_reg[114][24]/P0001 ,
		_w13202_,
		_w14643_
	);
	LUT2 #(
		.INIT('h8)
	) name4132 (
		\wishbone_bd_ram_mem3_reg[93][24]/P0001 ,
		_w13016_,
		_w14644_
	);
	LUT2 #(
		.INIT('h8)
	) name4133 (
		\wishbone_bd_ram_mem3_reg[141][24]/P0001 ,
		_w13004_,
		_w14645_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\wishbone_bd_ram_mem3_reg[146][24]/P0001 ,
		_w13060_,
		_w14646_
	);
	LUT2 #(
		.INIT('h8)
	) name4135 (
		\wishbone_bd_ram_mem3_reg[173][24]/P0001 ,
		_w12854_,
		_w14647_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		\wishbone_bd_ram_mem3_reg[226][24]/P0001 ,
		_w13138_,
		_w14648_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		\wishbone_bd_ram_mem3_reg[204][24]/P0001 ,
		_w13162_,
		_w14649_
	);
	LUT2 #(
		.INIT('h8)
	) name4138 (
		\wishbone_bd_ram_mem3_reg[24][24]/P0001 ,
		_w13084_,
		_w14650_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		\wishbone_bd_ram_mem3_reg[66][24]/P0001 ,
		_w12824_,
		_w14651_
	);
	LUT2 #(
		.INIT('h8)
	) name4140 (
		\wishbone_bd_ram_mem3_reg[105][24]/P0001 ,
		_w12751_,
		_w14652_
	);
	LUT2 #(
		.INIT('h8)
	) name4141 (
		\wishbone_bd_ram_mem3_reg[89][24]/P0001 ,
		_w12964_,
		_w14653_
	);
	LUT2 #(
		.INIT('h8)
	) name4142 (
		\wishbone_bd_ram_mem3_reg[224][24]/P0001 ,
		_w12902_,
		_w14654_
	);
	LUT2 #(
		.INIT('h8)
	) name4143 (
		\wishbone_bd_ram_mem3_reg[90][24]/P0001 ,
		_w12978_,
		_w14655_
	);
	LUT2 #(
		.INIT('h8)
	) name4144 (
		\wishbone_bd_ram_mem3_reg[184][24]/P0001 ,
		_w13062_,
		_w14656_
	);
	LUT2 #(
		.INIT('h8)
	) name4145 (
		\wishbone_bd_ram_mem3_reg[73][24]/P0001 ,
		_w12918_,
		_w14657_
	);
	LUT2 #(
		.INIT('h8)
	) name4146 (
		\wishbone_bd_ram_mem3_reg[31][24]/P0001 ,
		_w13198_,
		_w14658_
	);
	LUT2 #(
		.INIT('h8)
	) name4147 (
		\wishbone_bd_ram_mem3_reg[158][24]/P0001 ,
		_w12898_,
		_w14659_
	);
	LUT2 #(
		.INIT('h8)
	) name4148 (
		\wishbone_bd_ram_mem3_reg[26][24]/P0001 ,
		_w12699_,
		_w14660_
	);
	LUT2 #(
		.INIT('h8)
	) name4149 (
		\wishbone_bd_ram_mem3_reg[165][24]/P0001 ,
		_w13044_,
		_w14661_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		\wishbone_bd_ram_mem3_reg[209][24]/P0001 ,
		_w13152_,
		_w14662_
	);
	LUT2 #(
		.INIT('h8)
	) name4151 (
		\wishbone_bd_ram_mem3_reg[181][24]/P0001 ,
		_w12828_,
		_w14663_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		\wishbone_bd_ram_mem3_reg[244][24]/P0001 ,
		_w12747_,
		_w14664_
	);
	LUT2 #(
		.INIT('h8)
	) name4153 (
		\wishbone_bd_ram_mem3_reg[109][24]/P0001 ,
		_w12888_,
		_w14665_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		\wishbone_bd_ram_mem3_reg[88][24]/P0001 ,
		_w12860_,
		_w14666_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		\wishbone_bd_ram_mem3_reg[171][24]/P0001 ,
		_w12910_,
		_w14667_
	);
	LUT2 #(
		.INIT('h8)
	) name4156 (
		\wishbone_bd_ram_mem3_reg[40][24]/P0001 ,
		_w13132_,
		_w14668_
	);
	LUT2 #(
		.INIT('h8)
	) name4157 (
		\wishbone_bd_ram_mem3_reg[2][24]/P0001 ,
		_w13088_,
		_w14669_
	);
	LUT2 #(
		.INIT('h8)
	) name4158 (
		\wishbone_bd_ram_mem3_reg[75][24]/P0001 ,
		_w12826_,
		_w14670_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		\wishbone_bd_ram_mem3_reg[80][24]/P0001 ,
		_w12689_,
		_w14671_
	);
	LUT2 #(
		.INIT('h8)
	) name4160 (
		\wishbone_bd_ram_mem3_reg[140][24]/P0001 ,
		_w12894_,
		_w14672_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		\wishbone_bd_ram_mem3_reg[160][24]/P0001 ,
		_w12872_,
		_w14673_
	);
	LUT2 #(
		.INIT('h8)
	) name4162 (
		\wishbone_bd_ram_mem3_reg[219][24]/P0001 ,
		_w12806_,
		_w14674_
	);
	LUT2 #(
		.INIT('h8)
	) name4163 (
		\wishbone_bd_ram_mem3_reg[120][24]/P0001 ,
		_w12707_,
		_w14675_
	);
	LUT2 #(
		.INIT('h8)
	) name4164 (
		\wishbone_bd_ram_mem3_reg[250][24]/P0001 ,
		_w13128_,
		_w14676_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		\wishbone_bd_ram_mem3_reg[215][24]/P0001 ,
		_w12974_,
		_w14677_
	);
	LUT2 #(
		.INIT('h8)
	) name4166 (
		\wishbone_bd_ram_mem3_reg[67][24]/P0001 ,
		_w13134_,
		_w14678_
	);
	LUT2 #(
		.INIT('h8)
	) name4167 (
		\wishbone_bd_ram_mem3_reg[111][24]/P0001 ,
		_w12744_,
		_w14679_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		\wishbone_bd_ram_mem3_reg[228][24]/P0001 ,
		_w12765_,
		_w14680_
	);
	LUT2 #(
		.INIT('h8)
	) name4169 (
		\wishbone_bd_ram_mem3_reg[47][24]/P0001 ,
		_w12904_,
		_w14681_
	);
	LUT2 #(
		.INIT('h8)
	) name4170 (
		\wishbone_bd_ram_mem3_reg[185][24]/P0001 ,
		_w12940_,
		_w14682_
	);
	LUT2 #(
		.INIT('h8)
	) name4171 (
		\wishbone_bd_ram_mem3_reg[143][24]/P0001 ,
		_w12922_,
		_w14683_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\wishbone_bd_ram_mem3_reg[8][24]/P0001 ,
		_w12920_,
		_w14684_
	);
	LUT2 #(
		.INIT('h8)
	) name4173 (
		\wishbone_bd_ram_mem3_reg[142][24]/P0001 ,
		_w12928_,
		_w14685_
	);
	LUT2 #(
		.INIT('h8)
	) name4174 (
		\wishbone_bd_ram_mem3_reg[115][24]/P0001 ,
		_w13112_,
		_w14686_
	);
	LUT2 #(
		.INIT('h8)
	) name4175 (
		\wishbone_bd_ram_mem3_reg[154][24]/P0001 ,
		_w12962_,
		_w14687_
	);
	LUT2 #(
		.INIT('h8)
	) name4176 (
		\wishbone_bd_ram_mem3_reg[129][24]/P0001 ,
		_w12776_,
		_w14688_
	);
	LUT2 #(
		.INIT('h8)
	) name4177 (
		\wishbone_bd_ram_mem3_reg[172][24]/P0001 ,
		_w12944_,
		_w14689_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		\wishbone_bd_ram_mem3_reg[28][24]/P0001 ,
		_w13170_,
		_w14690_
	);
	LUT2 #(
		.INIT('h8)
	) name4179 (
		\wishbone_bd_ram_mem3_reg[249][24]/P0001 ,
		_w12900_,
		_w14691_
	);
	LUT2 #(
		.INIT('h8)
	) name4180 (
		\wishbone_bd_ram_mem3_reg[106][24]/P0001 ,
		_w12713_,
		_w14692_
	);
	LUT2 #(
		.INIT('h8)
	) name4181 (
		\wishbone_bd_ram_mem3_reg[65][24]/P0001 ,
		_w13176_,
		_w14693_
	);
	LUT2 #(
		.INIT('h8)
	) name4182 (
		\wishbone_bd_ram_mem3_reg[150][24]/P0001 ,
		_w13136_,
		_w14694_
	);
	LUT2 #(
		.INIT('h8)
	) name4183 (
		\wishbone_bd_ram_mem3_reg[178][24]/P0001 ,
		_w12886_,
		_w14695_
	);
	LUT2 #(
		.INIT('h8)
	) name4184 (
		\wishbone_bd_ram_mem3_reg[127][24]/P0001 ,
		_w13164_,
		_w14696_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		\wishbone_bd_ram_mem3_reg[60][24]/P0001 ,
		_w13204_,
		_w14697_
	);
	LUT2 #(
		.INIT('h8)
	) name4186 (
		\wishbone_bd_ram_mem3_reg[18][24]/P0001 ,
		_w12679_,
		_w14698_
	);
	LUT2 #(
		.INIT('h8)
	) name4187 (
		\wishbone_bd_ram_mem3_reg[168][24]/P0001 ,
		_w13208_,
		_w14699_
	);
	LUT2 #(
		.INIT('h8)
	) name4188 (
		\wishbone_bd_ram_mem3_reg[182][24]/P0001 ,
		_w12820_,
		_w14700_
	);
	LUT2 #(
		.INIT('h8)
	) name4189 (
		\wishbone_bd_ram_mem3_reg[230][24]/P0001 ,
		_w13036_,
		_w14701_
	);
	LUT2 #(
		.INIT('h8)
	) name4190 (
		\wishbone_bd_ram_mem3_reg[21][24]/P0001 ,
		_w12906_,
		_w14702_
	);
	LUT2 #(
		.INIT('h8)
	) name4191 (
		\wishbone_bd_ram_mem3_reg[22][24]/P0001 ,
		_w13110_,
		_w14703_
	);
	LUT2 #(
		.INIT('h8)
	) name4192 (
		\wishbone_bd_ram_mem3_reg[97][24]/P0001 ,
		_w13096_,
		_w14704_
	);
	LUT2 #(
		.INIT('h8)
	) name4193 (
		\wishbone_bd_ram_mem3_reg[255][24]/P0001 ,
		_w13072_,
		_w14705_
	);
	LUT2 #(
		.INIT('h8)
	) name4194 (
		\wishbone_bd_ram_mem3_reg[164][24]/P0001 ,
		_w12876_,
		_w14706_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		\wishbone_bd_ram_mem3_reg[41][24]/P0001 ,
		_w13052_,
		_w14707_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		\wishbone_bd_ram_mem3_reg[52][24]/P0001 ,
		_w13082_,
		_w14708_
	);
	LUT2 #(
		.INIT('h8)
	) name4197 (
		\wishbone_bd_ram_mem3_reg[147][24]/P0001 ,
		_w13146_,
		_w14709_
	);
	LUT2 #(
		.INIT('h8)
	) name4198 (
		\wishbone_bd_ram_mem3_reg[20][24]/P0001 ,
		_w13174_,
		_w14710_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		\wishbone_bd_ram_mem3_reg[247][24]/P0001 ,
		_w12818_,
		_w14711_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		\wishbone_bd_ram_mem3_reg[29][24]/P0001 ,
		_w12952_,
		_w14712_
	);
	LUT2 #(
		.INIT('h8)
	) name4201 (
		\wishbone_bd_ram_mem3_reg[216][24]/P0001 ,
		_w13028_,
		_w14713_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		\wishbone_bd_ram_mem3_reg[145][24]/P0001 ,
		_w13106_,
		_w14714_
	);
	LUT2 #(
		.INIT('h8)
	) name4203 (
		\wishbone_bd_ram_mem3_reg[212][24]/P0001 ,
		_w12796_,
		_w14715_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		\wishbone_bd_ram_mem3_reg[10][24]/P0001 ,
		_w13172_,
		_w14716_
	);
	LUT2 #(
		.INIT('h8)
	) name4205 (
		\wishbone_bd_ram_mem3_reg[139][24]/P0001 ,
		_w12814_,
		_w14717_
	);
	LUT2 #(
		.INIT('h8)
	) name4206 (
		\wishbone_bd_ram_mem3_reg[30][24]/P0001 ,
		_w13104_,
		_w14718_
	);
	LUT2 #(
		.INIT('h8)
	) name4207 (
		\wishbone_bd_ram_mem3_reg[132][24]/P0001 ,
		_w12992_,
		_w14719_
	);
	LUT2 #(
		.INIT('h8)
	) name4208 (
		\wishbone_bd_ram_mem3_reg[187][24]/P0001 ,
		_w13196_,
		_w14720_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		\wishbone_bd_ram_mem3_reg[43][24]/P0001 ,
		_w13200_,
		_w14721_
	);
	LUT2 #(
		.INIT('h8)
	) name4210 (
		\wishbone_bd_ram_mem3_reg[239][24]/P0001 ,
		_w12862_,
		_w14722_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		\wishbone_bd_ram_mem3_reg[192][24]/P0001 ,
		_w12938_,
		_w14723_
	);
	LUT2 #(
		.INIT('h8)
	) name4212 (
		\wishbone_bd_ram_mem3_reg[162][24]/P0001 ,
		_w13098_,
		_w14724_
	);
	LUT2 #(
		.INIT('h8)
	) name4213 (
		\wishbone_bd_ram_mem3_reg[36][24]/P0001 ,
		_w12800_,
		_w14725_
	);
	LUT2 #(
		.INIT('h8)
	) name4214 (
		\wishbone_bd_ram_mem3_reg[9][24]/P0001 ,
		_w12808_,
		_w14726_
	);
	LUT2 #(
		.INIT('h8)
	) name4215 (
		\wishbone_bd_ram_mem3_reg[108][24]/P0001 ,
		_w13156_,
		_w14727_
	);
	LUT2 #(
		.INIT('h8)
	) name4216 (
		\wishbone_bd_ram_mem3_reg[19][24]/P0001 ,
		_w13012_,
		_w14728_
	);
	LUT2 #(
		.INIT('h8)
	) name4217 (
		\wishbone_bd_ram_mem3_reg[15][24]/P0001 ,
		_w13210_,
		_w14729_
	);
	LUT2 #(
		.INIT('h8)
	) name4218 (
		\wishbone_bd_ram_mem3_reg[23][24]/P0001 ,
		_w13008_,
		_w14730_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		\wishbone_bd_ram_mem3_reg[98][24]/P0001 ,
		_w12816_,
		_w14731_
	);
	LUT2 #(
		.INIT('h8)
	) name4220 (
		\wishbone_bd_ram_mem3_reg[45][24]/P0001 ,
		_w12908_,
		_w14732_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		\wishbone_bd_ram_mem3_reg[86][24]/P0001 ,
		_w12735_,
		_w14733_
	);
	LUT2 #(
		.INIT('h8)
	) name4222 (
		\wishbone_bd_ram_mem3_reg[64][24]/P0001 ,
		_w12976_,
		_w14734_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		\wishbone_bd_ram_mem3_reg[183][24]/P0001 ,
		_w12787_,
		_w14735_
	);
	LUT2 #(
		.INIT('h8)
	) name4224 (
		\wishbone_bd_ram_mem3_reg[161][24]/P0001 ,
		_w12754_,
		_w14736_
	);
	LUT2 #(
		.INIT('h8)
	) name4225 (
		\wishbone_bd_ram_mem3_reg[190][24]/P0001 ,
		_w12858_,
		_w14737_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		\wishbone_bd_ram_mem3_reg[54][24]/P0001 ,
		_w12770_,
		_w14738_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		\wishbone_bd_ram_mem3_reg[179][24]/P0001 ,
		_w13050_,
		_w14739_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		\wishbone_bd_ram_mem3_reg[167][24]/P0001 ,
		_w12986_,
		_w14740_
	);
	LUT2 #(
		.INIT('h8)
	) name4229 (
		\wishbone_bd_ram_mem3_reg[202][24]/P0001 ,
		_w12870_,
		_w14741_
	);
	LUT2 #(
		.INIT('h8)
	) name4230 (
		\wishbone_bd_ram_mem3_reg[119][24]/P0001 ,
		_w13048_,
		_w14742_
	);
	LUT2 #(
		.INIT('h8)
	) name4231 (
		\wishbone_bd_ram_mem3_reg[231][24]/P0001 ,
		_w12856_,
		_w14743_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		\wishbone_bd_ram_mem3_reg[48][24]/P0001 ,
		_w12970_,
		_w14744_
	);
	LUT2 #(
		.INIT('h8)
	) name4233 (
		\wishbone_bd_ram_mem3_reg[12][24]/P0001 ,
		_w13118_,
		_w14745_
	);
	LUT2 #(
		.INIT('h8)
	) name4234 (
		\wishbone_bd_ram_mem3_reg[240][24]/P0001 ,
		_w12864_,
		_w14746_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		\wishbone_bd_ram_mem3_reg[37][24]/P0001 ,
		_w13102_,
		_w14747_
	);
	LUT2 #(
		.INIT('h8)
	) name4236 (
		\wishbone_bd_ram_mem3_reg[222][24]/P0001 ,
		_w13094_,
		_w14748_
	);
	LUT2 #(
		.INIT('h8)
	) name4237 (
		\wishbone_bd_ram_mem3_reg[92][24]/P0001 ,
		_w13010_,
		_w14749_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		\wishbone_bd_ram_mem3_reg[208][24]/P0001 ,
		_w13032_,
		_w14750_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		\wishbone_bd_ram_mem3_reg[51][24]/P0001 ,
		_w13024_,
		_w14751_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		\wishbone_bd_ram_mem3_reg[5][24]/P0001 ,
		_w12878_,
		_w14752_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		\wishbone_bd_ram_mem3_reg[155][24]/P0001 ,
		_w13122_,
		_w14753_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		\wishbone_bd_ram_mem3_reg[72][24]/P0001 ,
		_w12810_,
		_w14754_
	);
	LUT2 #(
		.INIT('h8)
	) name4243 (
		\wishbone_bd_ram_mem3_reg[138][24]/P0001 ,
		_w12958_,
		_w14755_
	);
	LUT2 #(
		.INIT('h8)
	) name4244 (
		\wishbone_bd_ram_mem3_reg[246][24]/P0001 ,
		_w13076_,
		_w14756_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		\wishbone_bd_ram_mem3_reg[210][24]/P0001 ,
		_w12924_,
		_w14757_
	);
	LUT2 #(
		.INIT('h8)
	) name4246 (
		\wishbone_bd_ram_mem3_reg[107][24]/P0001 ,
		_w12749_,
		_w14758_
	);
	LUT2 #(
		.INIT('h8)
	) name4247 (
		\wishbone_bd_ram_mem3_reg[136][24]/P0001 ,
		_w13064_,
		_w14759_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		\wishbone_bd_ram_mem3_reg[135][24]/P0001 ,
		_w13124_,
		_w14760_
	);
	LUT2 #(
		.INIT('h8)
	) name4249 (
		\wishbone_bd_ram_mem3_reg[87][24]/P0001 ,
		_w13154_,
		_w14761_
	);
	LUT2 #(
		.INIT('h8)
	) name4250 (
		\wishbone_bd_ram_mem3_reg[156][24]/P0001 ,
		_w13190_,
		_w14762_
	);
	LUT2 #(
		.INIT('h8)
	) name4251 (
		\wishbone_bd_ram_mem3_reg[79][24]/P0001 ,
		_w13212_,
		_w14763_
	);
	LUT2 #(
		.INIT('h8)
	) name4252 (
		\wishbone_bd_ram_mem3_reg[101][24]/P0001 ,
		_w13192_,
		_w14764_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		\wishbone_bd_ram_mem3_reg[199][24]/P0001 ,
		_w12768_,
		_w14765_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		\wishbone_bd_ram_mem3_reg[58][24]/P0001 ,
		_w13070_,
		_w14766_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		\wishbone_bd_ram_mem3_reg[198][24]/P0001 ,
		_w12832_,
		_w14767_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		\wishbone_bd_ram_mem3_reg[46][24]/P0001 ,
		_w12884_,
		_w14768_
	);
	LUT2 #(
		.INIT('h8)
	) name4257 (
		\wishbone_bd_ram_mem3_reg[96][24]/P0001 ,
		_w12912_,
		_w14769_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		\wishbone_bd_ram_mem3_reg[203][24]/P0001 ,
		_w13158_,
		_w14770_
	);
	LUT2 #(
		.INIT('h8)
	) name4259 (
		\wishbone_bd_ram_mem3_reg[207][24]/P0001 ,
		_w13180_,
		_w14771_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		\wishbone_bd_ram_mem3_reg[248][24]/P0001 ,
		_w12789_,
		_w14772_
	);
	LUT2 #(
		.INIT('h8)
	) name4261 (
		\wishbone_bd_ram_mem3_reg[94][24]/P0001 ,
		_w13186_,
		_w14773_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		\wishbone_bd_ram_mem3_reg[7][24]/P0001 ,
		_w12728_,
		_w14774_
	);
	LUT2 #(
		.INIT('h8)
	) name4263 (
		\wishbone_bd_ram_mem3_reg[148][24]/P0001 ,
		_w13000_,
		_w14775_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		\wishbone_bd_ram_mem3_reg[134][24]/P0001 ,
		_w12763_,
		_w14776_
	);
	LUT2 #(
		.INIT('h8)
	) name4265 (
		\wishbone_bd_ram_mem3_reg[163][24]/P0001 ,
		_w12882_,
		_w14777_
	);
	LUT2 #(
		.INIT('h8)
	) name4266 (
		\wishbone_bd_ram_mem3_reg[186][24]/P0001 ,
		_w12783_,
		_w14778_
	);
	LUT2 #(
		.INIT('h8)
	) name4267 (
		\wishbone_bd_ram_mem3_reg[235][24]/P0001 ,
		_w12696_,
		_w14779_
	);
	LUT2 #(
		.INIT('h8)
	) name4268 (
		\wishbone_bd_ram_mem3_reg[42][24]/P0001 ,
		_w12842_,
		_w14780_
	);
	LUT2 #(
		.INIT('h8)
	) name4269 (
		\wishbone_bd_ram_mem3_reg[200][24]/P0001 ,
		_w12988_,
		_w14781_
	);
	LUT2 #(
		.INIT('h8)
	) name4270 (
		\wishbone_bd_ram_mem3_reg[112][24]/P0001 ,
		_w12733_,
		_w14782_
	);
	LUT2 #(
		.INIT('h8)
	) name4271 (
		\wishbone_bd_ram_mem3_reg[251][24]/P0001 ,
		_w13054_,
		_w14783_
	);
	LUT2 #(
		.INIT('h8)
	) name4272 (
		\wishbone_bd_ram_mem3_reg[151][24]/P0001 ,
		_w13142_,
		_w14784_
	);
	LUT2 #(
		.INIT('h8)
	) name4273 (
		\wishbone_bd_ram_mem3_reg[254][24]/P0001 ,
		_w12892_,
		_w14785_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		\wishbone_bd_ram_mem3_reg[103][24]/P0001 ,
		_w12846_,
		_w14786_
	);
	LUT2 #(
		.INIT('h8)
	) name4275 (
		\wishbone_bd_ram_mem3_reg[69][24]/P0001 ,
		_w12738_,
		_w14787_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		\wishbone_bd_ram_mem3_reg[225][24]/P0001 ,
		_w13092_,
		_w14788_
	);
	LUT2 #(
		.INIT('h8)
	) name4277 (
		\wishbone_bd_ram_mem3_reg[1][24]/P0001 ,
		_w13014_,
		_w14789_
	);
	LUT2 #(
		.INIT('h8)
	) name4278 (
		\wishbone_bd_ram_mem3_reg[70][24]/P0001 ,
		_w12840_,
		_w14790_
	);
	LUT2 #(
		.INIT('h8)
	) name4279 (
		\wishbone_bd_ram_mem3_reg[238][24]/P0001 ,
		_w13160_,
		_w14791_
	);
	LUT2 #(
		.INIT('h8)
	) name4280 (
		\wishbone_bd_ram_mem3_reg[124][24]/P0001 ,
		_w13058_,
		_w14792_
	);
	LUT2 #(
		.INIT('h8)
	) name4281 (
		\wishbone_bd_ram_mem3_reg[234][24]/P0001 ,
		_w13214_,
		_w14793_
	);
	LUT2 #(
		.INIT('h8)
	) name4282 (
		\wishbone_bd_ram_mem3_reg[232][24]/P0001 ,
		_w12758_,
		_w14794_
	);
	LUT2 #(
		.INIT('h8)
	) name4283 (
		\wishbone_bd_ram_mem3_reg[214][24]/P0001 ,
		_w12984_,
		_w14795_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		\wishbone_bd_ram_mem3_reg[177][24]/P0001 ,
		_w12996_,
		_w14796_
	);
	LUT2 #(
		.INIT('h8)
	) name4285 (
		\wishbone_bd_ram_mem3_reg[166][24]/P0001 ,
		_w13040_,
		_w14797_
	);
	LUT2 #(
		.INIT('h8)
	) name4286 (
		\wishbone_bd_ram_mem3_reg[102][24]/P0001 ,
		_w12685_,
		_w14798_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		\wishbone_bd_ram_mem3_reg[11][24]/P0001 ,
		_w13194_,
		_w14799_
	);
	LUT2 #(
		.INIT('h8)
	) name4288 (
		\wishbone_bd_ram_mem3_reg[53][24]/P0001 ,
		_w13020_,
		_w14800_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		\wishbone_bd_ram_mem3_reg[169][24]/P0001 ,
		_w12722_,
		_w14801_
	);
	LUT2 #(
		.INIT('h8)
	) name4290 (
		\wishbone_bd_ram_mem3_reg[59][24]/P0001 ,
		_w12780_,
		_w14802_
	);
	LUT2 #(
		.INIT('h8)
	) name4291 (
		\wishbone_bd_ram_mem3_reg[118][24]/P0001 ,
		_w12830_,
		_w14803_
	);
	LUT2 #(
		.INIT('h8)
	) name4292 (
		\wishbone_bd_ram_mem3_reg[50][24]/P0001 ,
		_w13150_,
		_w14804_
	);
	LUT2 #(
		.INIT('h8)
	) name4293 (
		\wishbone_bd_ram_mem3_reg[81][24]/P0001 ,
		_w12950_,
		_w14805_
	);
	LUT2 #(
		.INIT('h8)
	) name4294 (
		\wishbone_bd_ram_mem3_reg[82][24]/P0001 ,
		_w12942_,
		_w14806_
	);
	LUT2 #(
		.INIT('h8)
	) name4295 (
		\wishbone_bd_ram_mem3_reg[68][24]/P0001 ,
		_w12946_,
		_w14807_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		\wishbone_bd_ram_mem3_reg[38][24]/P0001 ,
		_w13182_,
		_w14808_
	);
	LUT2 #(
		.INIT('h8)
	) name4297 (
		\wishbone_bd_ram_mem3_reg[233][24]/P0001 ,
		_w12836_,
		_w14809_
	);
	LUT2 #(
		.INIT('h8)
	) name4298 (
		\wishbone_bd_ram_mem3_reg[117][24]/P0001 ,
		_w12715_,
		_w14810_
	);
	LUT2 #(
		.INIT('h8)
	) name4299 (
		\wishbone_bd_ram_mem3_reg[153][24]/P0001 ,
		_w12890_,
		_w14811_
	);
	LUT2 #(
		.INIT('h8)
	) name4300 (
		\wishbone_bd_ram_mem3_reg[44][24]/P0001 ,
		_w12896_,
		_w14812_
	);
	LUT2 #(
		.INIT('h8)
	) name4301 (
		\wishbone_bd_ram_mem3_reg[191][24]/P0001 ,
		_w13034_,
		_w14813_
	);
	LUT2 #(
		.INIT('h8)
	) name4302 (
		\wishbone_bd_ram_mem3_reg[217][24]/P0001 ,
		_w13188_,
		_w14814_
	);
	LUT2 #(
		.INIT('h8)
	) name4303 (
		\wishbone_bd_ram_mem3_reg[77][24]/P0001 ,
		_w12982_,
		_w14815_
	);
	LUT2 #(
		.INIT('h8)
	) name4304 (
		\wishbone_bd_ram_mem3_reg[125][24]/P0001 ,
		_w12956_,
		_w14816_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		\wishbone_bd_ram_mem3_reg[237][24]/P0001 ,
		_w12990_,
		_w14817_
	);
	LUT2 #(
		.INIT('h8)
	) name4306 (
		\wishbone_bd_ram_mem3_reg[195][24]/P0001 ,
		_w13144_,
		_w14818_
	);
	LUT2 #(
		.INIT('h8)
	) name4307 (
		\wishbone_bd_ram_mem3_reg[189][24]/P0001 ,
		_w13042_,
		_w14819_
	);
	LUT2 #(
		.INIT('h8)
	) name4308 (
		\wishbone_bd_ram_mem3_reg[180][24]/P0001 ,
		_w12791_,
		_w14820_
	);
	LUT2 #(
		.INIT('h8)
	) name4309 (
		\wishbone_bd_ram_mem3_reg[243][24]/P0001 ,
		_w12804_,
		_w14821_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		\wishbone_bd_ram_mem3_reg[116][24]/P0001 ,
		_w12998_,
		_w14822_
	);
	LUT2 #(
		.INIT('h8)
	) name4311 (
		\wishbone_bd_ram_mem3_reg[174][24]/P0001 ,
		_w12972_,
		_w14823_
	);
	LUT2 #(
		.INIT('h8)
	) name4312 (
		\wishbone_bd_ram_mem3_reg[242][24]/P0001 ,
		_w12932_,
		_w14824_
	);
	LUT2 #(
		.INIT('h8)
	) name4313 (
		\wishbone_bd_ram_mem3_reg[194][24]/P0001 ,
		_w12772_,
		_w14825_
	);
	LUT2 #(
		.INIT('h8)
	) name4314 (
		\wishbone_bd_ram_mem3_reg[223][24]/P0001 ,
		_w12838_,
		_w14826_
	);
	LUT2 #(
		.INIT('h8)
	) name4315 (
		\wishbone_bd_ram_mem3_reg[128][24]/P0001 ,
		_w12793_,
		_w14827_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\wishbone_bd_ram_mem3_reg[113][24]/P0001 ,
		_w13026_,
		_w14828_
	);
	LUT2 #(
		.INIT('h8)
	) name4317 (
		\wishbone_bd_ram_mem3_reg[123][24]/P0001 ,
		_w13114_,
		_w14829_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		\wishbone_bd_ram_mem3_reg[206][24]/P0001 ,
		_w12954_,
		_w14830_
	);
	LUT2 #(
		.INIT('h8)
	) name4319 (
		\wishbone_bd_ram_mem3_reg[74][24]/P0001 ,
		_w12812_,
		_w14831_
	);
	LUT2 #(
		.INIT('h8)
	) name4320 (
		\wishbone_bd_ram_mem3_reg[56][24]/P0001 ,
		_w12778_,
		_w14832_
	);
	LUT2 #(
		.INIT('h8)
	) name4321 (
		\wishbone_bd_ram_mem3_reg[95][24]/P0001 ,
		_w12844_,
		_w14833_
	);
	LUT2 #(
		.INIT('h8)
	) name4322 (
		\wishbone_bd_ram_mem3_reg[49][24]/P0001 ,
		_w12994_,
		_w14834_
	);
	LUT2 #(
		.INIT('h8)
	) name4323 (
		\wishbone_bd_ram_mem3_reg[221][24]/P0001 ,
		_w12802_,
		_w14835_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		\wishbone_bd_ram_mem3_reg[85][24]/P0001 ,
		_w13216_,
		_w14836_
	);
	LUT2 #(
		.INIT('h8)
	) name4325 (
		\wishbone_bd_ram_mem3_reg[63][24]/P0001 ,
		_w12850_,
		_w14837_
	);
	LUT2 #(
		.INIT('h8)
	) name4326 (
		\wishbone_bd_ram_mem3_reg[71][24]/P0001 ,
		_w12798_,
		_w14838_
	);
	LUT2 #(
		.INIT('h8)
	) name4327 (
		\wishbone_bd_ram_mem3_reg[253][24]/P0001 ,
		_w13100_,
		_w14839_
	);
	LUT2 #(
		.INIT('h8)
	) name4328 (
		\wishbone_bd_ram_mem3_reg[62][24]/P0001 ,
		_w12673_,
		_w14840_
	);
	LUT2 #(
		.INIT('h8)
	) name4329 (
		\wishbone_bd_ram_mem3_reg[122][24]/P0001 ,
		_w13130_,
		_w14841_
	);
	LUT2 #(
		.INIT('h8)
	) name4330 (
		\wishbone_bd_ram_mem3_reg[6][24]/P0001 ,
		_w12968_,
		_w14842_
	);
	LUT2 #(
		.INIT('h8)
	) name4331 (
		\wishbone_bd_ram_mem3_reg[213][24]/P0001 ,
		_w13002_,
		_w14843_
	);
	LUT2 #(
		.INIT('h8)
	) name4332 (
		\wishbone_bd_ram_mem3_reg[76][24]/P0001 ,
		_w13184_,
		_w14844_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		\wishbone_bd_ram_mem3_reg[16][24]/P0001 ,
		_w13140_,
		_w14845_
	);
	LUT2 #(
		.INIT('h8)
	) name4334 (
		\wishbone_bd_ram_mem3_reg[175][24]/P0001 ,
		_w13126_,
		_w14846_
	);
	LUT2 #(
		.INIT('h8)
	) name4335 (
		\wishbone_bd_ram_mem3_reg[27][24]/P0001 ,
		_w12880_,
		_w14847_
	);
	LUT2 #(
		.INIT('h8)
	) name4336 (
		\wishbone_bd_ram_mem3_reg[159][24]/P0001 ,
		_w12774_,
		_w14848_
	);
	LUT2 #(
		.INIT('h8)
	) name4337 (
		\wishbone_bd_ram_mem3_reg[32][24]/P0001 ,
		_w13120_,
		_w14849_
	);
	LUT2 #(
		.INIT('h8)
	) name4338 (
		\wishbone_bd_ram_mem3_reg[14][24]/P0001 ,
		_w13086_,
		_w14850_
	);
	LUT2 #(
		.INIT('h8)
	) name4339 (
		\wishbone_bd_ram_mem3_reg[13][24]/P0001 ,
		_w13178_,
		_w14851_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		\wishbone_bd_ram_mem3_reg[193][24]/P0001 ,
		_w13056_,
		_w14852_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		\wishbone_bd_ram_mem3_reg[4][24]/P0001 ,
		_w12666_,
		_w14853_
	);
	LUT2 #(
		.INIT('h8)
	) name4342 (
		\wishbone_bd_ram_mem3_reg[236][24]/P0001 ,
		_w12731_,
		_w14854_
	);
	LUT2 #(
		.INIT('h1)
	) name4343 (
		_w14599_,
		_w14600_,
		_w14855_
	);
	LUT2 #(
		.INIT('h1)
	) name4344 (
		_w14601_,
		_w14602_,
		_w14856_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		_w14603_,
		_w14604_,
		_w14857_
	);
	LUT2 #(
		.INIT('h1)
	) name4346 (
		_w14605_,
		_w14606_,
		_w14858_
	);
	LUT2 #(
		.INIT('h1)
	) name4347 (
		_w14607_,
		_w14608_,
		_w14859_
	);
	LUT2 #(
		.INIT('h1)
	) name4348 (
		_w14609_,
		_w14610_,
		_w14860_
	);
	LUT2 #(
		.INIT('h1)
	) name4349 (
		_w14611_,
		_w14612_,
		_w14861_
	);
	LUT2 #(
		.INIT('h1)
	) name4350 (
		_w14613_,
		_w14614_,
		_w14862_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w14615_,
		_w14616_,
		_w14863_
	);
	LUT2 #(
		.INIT('h1)
	) name4352 (
		_w14617_,
		_w14618_,
		_w14864_
	);
	LUT2 #(
		.INIT('h1)
	) name4353 (
		_w14619_,
		_w14620_,
		_w14865_
	);
	LUT2 #(
		.INIT('h1)
	) name4354 (
		_w14621_,
		_w14622_,
		_w14866_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w14623_,
		_w14624_,
		_w14867_
	);
	LUT2 #(
		.INIT('h1)
	) name4356 (
		_w14625_,
		_w14626_,
		_w14868_
	);
	LUT2 #(
		.INIT('h1)
	) name4357 (
		_w14627_,
		_w14628_,
		_w14869_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w14629_,
		_w14630_,
		_w14870_
	);
	LUT2 #(
		.INIT('h1)
	) name4359 (
		_w14631_,
		_w14632_,
		_w14871_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w14633_,
		_w14634_,
		_w14872_
	);
	LUT2 #(
		.INIT('h1)
	) name4361 (
		_w14635_,
		_w14636_,
		_w14873_
	);
	LUT2 #(
		.INIT('h1)
	) name4362 (
		_w14637_,
		_w14638_,
		_w14874_
	);
	LUT2 #(
		.INIT('h1)
	) name4363 (
		_w14639_,
		_w14640_,
		_w14875_
	);
	LUT2 #(
		.INIT('h1)
	) name4364 (
		_w14641_,
		_w14642_,
		_w14876_
	);
	LUT2 #(
		.INIT('h1)
	) name4365 (
		_w14643_,
		_w14644_,
		_w14877_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w14645_,
		_w14646_,
		_w14878_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w14647_,
		_w14648_,
		_w14879_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w14649_,
		_w14650_,
		_w14880_
	);
	LUT2 #(
		.INIT('h1)
	) name4369 (
		_w14651_,
		_w14652_,
		_w14881_
	);
	LUT2 #(
		.INIT('h1)
	) name4370 (
		_w14653_,
		_w14654_,
		_w14882_
	);
	LUT2 #(
		.INIT('h1)
	) name4371 (
		_w14655_,
		_w14656_,
		_w14883_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w14657_,
		_w14658_,
		_w14884_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w14659_,
		_w14660_,
		_w14885_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w14661_,
		_w14662_,
		_w14886_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w14663_,
		_w14664_,
		_w14887_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w14665_,
		_w14666_,
		_w14888_
	);
	LUT2 #(
		.INIT('h1)
	) name4377 (
		_w14667_,
		_w14668_,
		_w14889_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		_w14669_,
		_w14670_,
		_w14890_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w14671_,
		_w14672_,
		_w14891_
	);
	LUT2 #(
		.INIT('h1)
	) name4380 (
		_w14673_,
		_w14674_,
		_w14892_
	);
	LUT2 #(
		.INIT('h1)
	) name4381 (
		_w14675_,
		_w14676_,
		_w14893_
	);
	LUT2 #(
		.INIT('h1)
	) name4382 (
		_w14677_,
		_w14678_,
		_w14894_
	);
	LUT2 #(
		.INIT('h1)
	) name4383 (
		_w14679_,
		_w14680_,
		_w14895_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		_w14681_,
		_w14682_,
		_w14896_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		_w14683_,
		_w14684_,
		_w14897_
	);
	LUT2 #(
		.INIT('h1)
	) name4386 (
		_w14685_,
		_w14686_,
		_w14898_
	);
	LUT2 #(
		.INIT('h1)
	) name4387 (
		_w14687_,
		_w14688_,
		_w14899_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w14689_,
		_w14690_,
		_w14900_
	);
	LUT2 #(
		.INIT('h1)
	) name4389 (
		_w14691_,
		_w14692_,
		_w14901_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w14693_,
		_w14694_,
		_w14902_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w14695_,
		_w14696_,
		_w14903_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		_w14697_,
		_w14698_,
		_w14904_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w14699_,
		_w14700_,
		_w14905_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w14701_,
		_w14702_,
		_w14906_
	);
	LUT2 #(
		.INIT('h1)
	) name4395 (
		_w14703_,
		_w14704_,
		_w14907_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w14705_,
		_w14706_,
		_w14908_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w14707_,
		_w14708_,
		_w14909_
	);
	LUT2 #(
		.INIT('h1)
	) name4398 (
		_w14709_,
		_w14710_,
		_w14910_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w14711_,
		_w14712_,
		_w14911_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w14713_,
		_w14714_,
		_w14912_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w14715_,
		_w14716_,
		_w14913_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		_w14717_,
		_w14718_,
		_w14914_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w14719_,
		_w14720_,
		_w14915_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w14721_,
		_w14722_,
		_w14916_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w14723_,
		_w14724_,
		_w14917_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w14725_,
		_w14726_,
		_w14918_
	);
	LUT2 #(
		.INIT('h1)
	) name4407 (
		_w14727_,
		_w14728_,
		_w14919_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w14729_,
		_w14730_,
		_w14920_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w14731_,
		_w14732_,
		_w14921_
	);
	LUT2 #(
		.INIT('h1)
	) name4410 (
		_w14733_,
		_w14734_,
		_w14922_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w14735_,
		_w14736_,
		_w14923_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w14737_,
		_w14738_,
		_w14924_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w14739_,
		_w14740_,
		_w14925_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		_w14741_,
		_w14742_,
		_w14926_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w14743_,
		_w14744_,
		_w14927_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		_w14745_,
		_w14746_,
		_w14928_
	);
	LUT2 #(
		.INIT('h1)
	) name4417 (
		_w14747_,
		_w14748_,
		_w14929_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		_w14749_,
		_w14750_,
		_w14930_
	);
	LUT2 #(
		.INIT('h1)
	) name4419 (
		_w14751_,
		_w14752_,
		_w14931_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		_w14753_,
		_w14754_,
		_w14932_
	);
	LUT2 #(
		.INIT('h1)
	) name4421 (
		_w14755_,
		_w14756_,
		_w14933_
	);
	LUT2 #(
		.INIT('h1)
	) name4422 (
		_w14757_,
		_w14758_,
		_w14934_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w14759_,
		_w14760_,
		_w14935_
	);
	LUT2 #(
		.INIT('h1)
	) name4424 (
		_w14761_,
		_w14762_,
		_w14936_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		_w14763_,
		_w14764_,
		_w14937_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w14765_,
		_w14766_,
		_w14938_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w14767_,
		_w14768_,
		_w14939_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w14769_,
		_w14770_,
		_w14940_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w14771_,
		_w14772_,
		_w14941_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w14773_,
		_w14774_,
		_w14942_
	);
	LUT2 #(
		.INIT('h1)
	) name4431 (
		_w14775_,
		_w14776_,
		_w14943_
	);
	LUT2 #(
		.INIT('h1)
	) name4432 (
		_w14777_,
		_w14778_,
		_w14944_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w14779_,
		_w14780_,
		_w14945_
	);
	LUT2 #(
		.INIT('h1)
	) name4434 (
		_w14781_,
		_w14782_,
		_w14946_
	);
	LUT2 #(
		.INIT('h1)
	) name4435 (
		_w14783_,
		_w14784_,
		_w14947_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w14785_,
		_w14786_,
		_w14948_
	);
	LUT2 #(
		.INIT('h1)
	) name4437 (
		_w14787_,
		_w14788_,
		_w14949_
	);
	LUT2 #(
		.INIT('h1)
	) name4438 (
		_w14789_,
		_w14790_,
		_w14950_
	);
	LUT2 #(
		.INIT('h1)
	) name4439 (
		_w14791_,
		_w14792_,
		_w14951_
	);
	LUT2 #(
		.INIT('h1)
	) name4440 (
		_w14793_,
		_w14794_,
		_w14952_
	);
	LUT2 #(
		.INIT('h1)
	) name4441 (
		_w14795_,
		_w14796_,
		_w14953_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		_w14797_,
		_w14798_,
		_w14954_
	);
	LUT2 #(
		.INIT('h1)
	) name4443 (
		_w14799_,
		_w14800_,
		_w14955_
	);
	LUT2 #(
		.INIT('h1)
	) name4444 (
		_w14801_,
		_w14802_,
		_w14956_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		_w14803_,
		_w14804_,
		_w14957_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w14805_,
		_w14806_,
		_w14958_
	);
	LUT2 #(
		.INIT('h1)
	) name4447 (
		_w14807_,
		_w14808_,
		_w14959_
	);
	LUT2 #(
		.INIT('h1)
	) name4448 (
		_w14809_,
		_w14810_,
		_w14960_
	);
	LUT2 #(
		.INIT('h1)
	) name4449 (
		_w14811_,
		_w14812_,
		_w14961_
	);
	LUT2 #(
		.INIT('h1)
	) name4450 (
		_w14813_,
		_w14814_,
		_w14962_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w14815_,
		_w14816_,
		_w14963_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w14817_,
		_w14818_,
		_w14964_
	);
	LUT2 #(
		.INIT('h1)
	) name4453 (
		_w14819_,
		_w14820_,
		_w14965_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w14821_,
		_w14822_,
		_w14966_
	);
	LUT2 #(
		.INIT('h1)
	) name4455 (
		_w14823_,
		_w14824_,
		_w14967_
	);
	LUT2 #(
		.INIT('h1)
	) name4456 (
		_w14825_,
		_w14826_,
		_w14968_
	);
	LUT2 #(
		.INIT('h1)
	) name4457 (
		_w14827_,
		_w14828_,
		_w14969_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w14829_,
		_w14830_,
		_w14970_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w14831_,
		_w14832_,
		_w14971_
	);
	LUT2 #(
		.INIT('h1)
	) name4460 (
		_w14833_,
		_w14834_,
		_w14972_
	);
	LUT2 #(
		.INIT('h1)
	) name4461 (
		_w14835_,
		_w14836_,
		_w14973_
	);
	LUT2 #(
		.INIT('h1)
	) name4462 (
		_w14837_,
		_w14838_,
		_w14974_
	);
	LUT2 #(
		.INIT('h1)
	) name4463 (
		_w14839_,
		_w14840_,
		_w14975_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		_w14841_,
		_w14842_,
		_w14976_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		_w14843_,
		_w14844_,
		_w14977_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		_w14845_,
		_w14846_,
		_w14978_
	);
	LUT2 #(
		.INIT('h1)
	) name4467 (
		_w14847_,
		_w14848_,
		_w14979_
	);
	LUT2 #(
		.INIT('h1)
	) name4468 (
		_w14849_,
		_w14850_,
		_w14980_
	);
	LUT2 #(
		.INIT('h1)
	) name4469 (
		_w14851_,
		_w14852_,
		_w14981_
	);
	LUT2 #(
		.INIT('h1)
	) name4470 (
		_w14853_,
		_w14854_,
		_w14982_
	);
	LUT2 #(
		.INIT('h8)
	) name4471 (
		_w14981_,
		_w14982_,
		_w14983_
	);
	LUT2 #(
		.INIT('h8)
	) name4472 (
		_w14979_,
		_w14980_,
		_w14984_
	);
	LUT2 #(
		.INIT('h8)
	) name4473 (
		_w14977_,
		_w14978_,
		_w14985_
	);
	LUT2 #(
		.INIT('h8)
	) name4474 (
		_w14975_,
		_w14976_,
		_w14986_
	);
	LUT2 #(
		.INIT('h8)
	) name4475 (
		_w14973_,
		_w14974_,
		_w14987_
	);
	LUT2 #(
		.INIT('h8)
	) name4476 (
		_w14971_,
		_w14972_,
		_w14988_
	);
	LUT2 #(
		.INIT('h8)
	) name4477 (
		_w14969_,
		_w14970_,
		_w14989_
	);
	LUT2 #(
		.INIT('h8)
	) name4478 (
		_w14967_,
		_w14968_,
		_w14990_
	);
	LUT2 #(
		.INIT('h8)
	) name4479 (
		_w14965_,
		_w14966_,
		_w14991_
	);
	LUT2 #(
		.INIT('h8)
	) name4480 (
		_w14963_,
		_w14964_,
		_w14992_
	);
	LUT2 #(
		.INIT('h8)
	) name4481 (
		_w14961_,
		_w14962_,
		_w14993_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w14959_,
		_w14960_,
		_w14994_
	);
	LUT2 #(
		.INIT('h8)
	) name4483 (
		_w14957_,
		_w14958_,
		_w14995_
	);
	LUT2 #(
		.INIT('h8)
	) name4484 (
		_w14955_,
		_w14956_,
		_w14996_
	);
	LUT2 #(
		.INIT('h8)
	) name4485 (
		_w14953_,
		_w14954_,
		_w14997_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		_w14951_,
		_w14952_,
		_w14998_
	);
	LUT2 #(
		.INIT('h8)
	) name4487 (
		_w14949_,
		_w14950_,
		_w14999_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		_w14947_,
		_w14948_,
		_w15000_
	);
	LUT2 #(
		.INIT('h8)
	) name4489 (
		_w14945_,
		_w14946_,
		_w15001_
	);
	LUT2 #(
		.INIT('h8)
	) name4490 (
		_w14943_,
		_w14944_,
		_w15002_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		_w14941_,
		_w14942_,
		_w15003_
	);
	LUT2 #(
		.INIT('h8)
	) name4492 (
		_w14939_,
		_w14940_,
		_w15004_
	);
	LUT2 #(
		.INIT('h8)
	) name4493 (
		_w14937_,
		_w14938_,
		_w15005_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		_w14935_,
		_w14936_,
		_w15006_
	);
	LUT2 #(
		.INIT('h8)
	) name4495 (
		_w14933_,
		_w14934_,
		_w15007_
	);
	LUT2 #(
		.INIT('h8)
	) name4496 (
		_w14931_,
		_w14932_,
		_w15008_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		_w14929_,
		_w14930_,
		_w15009_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		_w14927_,
		_w14928_,
		_w15010_
	);
	LUT2 #(
		.INIT('h8)
	) name4499 (
		_w14925_,
		_w14926_,
		_w15011_
	);
	LUT2 #(
		.INIT('h8)
	) name4500 (
		_w14923_,
		_w14924_,
		_w15012_
	);
	LUT2 #(
		.INIT('h8)
	) name4501 (
		_w14921_,
		_w14922_,
		_w15013_
	);
	LUT2 #(
		.INIT('h8)
	) name4502 (
		_w14919_,
		_w14920_,
		_w15014_
	);
	LUT2 #(
		.INIT('h8)
	) name4503 (
		_w14917_,
		_w14918_,
		_w15015_
	);
	LUT2 #(
		.INIT('h8)
	) name4504 (
		_w14915_,
		_w14916_,
		_w15016_
	);
	LUT2 #(
		.INIT('h8)
	) name4505 (
		_w14913_,
		_w14914_,
		_w15017_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		_w14911_,
		_w14912_,
		_w15018_
	);
	LUT2 #(
		.INIT('h8)
	) name4507 (
		_w14909_,
		_w14910_,
		_w15019_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		_w14907_,
		_w14908_,
		_w15020_
	);
	LUT2 #(
		.INIT('h8)
	) name4509 (
		_w14905_,
		_w14906_,
		_w15021_
	);
	LUT2 #(
		.INIT('h8)
	) name4510 (
		_w14903_,
		_w14904_,
		_w15022_
	);
	LUT2 #(
		.INIT('h8)
	) name4511 (
		_w14901_,
		_w14902_,
		_w15023_
	);
	LUT2 #(
		.INIT('h8)
	) name4512 (
		_w14899_,
		_w14900_,
		_w15024_
	);
	LUT2 #(
		.INIT('h8)
	) name4513 (
		_w14897_,
		_w14898_,
		_w15025_
	);
	LUT2 #(
		.INIT('h8)
	) name4514 (
		_w14895_,
		_w14896_,
		_w15026_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		_w14893_,
		_w14894_,
		_w15027_
	);
	LUT2 #(
		.INIT('h8)
	) name4516 (
		_w14891_,
		_w14892_,
		_w15028_
	);
	LUT2 #(
		.INIT('h8)
	) name4517 (
		_w14889_,
		_w14890_,
		_w15029_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		_w14887_,
		_w14888_,
		_w15030_
	);
	LUT2 #(
		.INIT('h8)
	) name4519 (
		_w14885_,
		_w14886_,
		_w15031_
	);
	LUT2 #(
		.INIT('h8)
	) name4520 (
		_w14883_,
		_w14884_,
		_w15032_
	);
	LUT2 #(
		.INIT('h8)
	) name4521 (
		_w14881_,
		_w14882_,
		_w15033_
	);
	LUT2 #(
		.INIT('h8)
	) name4522 (
		_w14879_,
		_w14880_,
		_w15034_
	);
	LUT2 #(
		.INIT('h8)
	) name4523 (
		_w14877_,
		_w14878_,
		_w15035_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		_w14875_,
		_w14876_,
		_w15036_
	);
	LUT2 #(
		.INIT('h8)
	) name4525 (
		_w14873_,
		_w14874_,
		_w15037_
	);
	LUT2 #(
		.INIT('h8)
	) name4526 (
		_w14871_,
		_w14872_,
		_w15038_
	);
	LUT2 #(
		.INIT('h8)
	) name4527 (
		_w14869_,
		_w14870_,
		_w15039_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		_w14867_,
		_w14868_,
		_w15040_
	);
	LUT2 #(
		.INIT('h8)
	) name4529 (
		_w14865_,
		_w14866_,
		_w15041_
	);
	LUT2 #(
		.INIT('h8)
	) name4530 (
		_w14863_,
		_w14864_,
		_w15042_
	);
	LUT2 #(
		.INIT('h8)
	) name4531 (
		_w14861_,
		_w14862_,
		_w15043_
	);
	LUT2 #(
		.INIT('h8)
	) name4532 (
		_w14859_,
		_w14860_,
		_w15044_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		_w14857_,
		_w14858_,
		_w15045_
	);
	LUT2 #(
		.INIT('h8)
	) name4534 (
		_w14855_,
		_w14856_,
		_w15046_
	);
	LUT2 #(
		.INIT('h8)
	) name4535 (
		_w15045_,
		_w15046_,
		_w15047_
	);
	LUT2 #(
		.INIT('h8)
	) name4536 (
		_w15043_,
		_w15044_,
		_w15048_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		_w15041_,
		_w15042_,
		_w15049_
	);
	LUT2 #(
		.INIT('h8)
	) name4538 (
		_w15039_,
		_w15040_,
		_w15050_
	);
	LUT2 #(
		.INIT('h8)
	) name4539 (
		_w15037_,
		_w15038_,
		_w15051_
	);
	LUT2 #(
		.INIT('h8)
	) name4540 (
		_w15035_,
		_w15036_,
		_w15052_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		_w15033_,
		_w15034_,
		_w15053_
	);
	LUT2 #(
		.INIT('h8)
	) name4542 (
		_w15031_,
		_w15032_,
		_w15054_
	);
	LUT2 #(
		.INIT('h8)
	) name4543 (
		_w15029_,
		_w15030_,
		_w15055_
	);
	LUT2 #(
		.INIT('h8)
	) name4544 (
		_w15027_,
		_w15028_,
		_w15056_
	);
	LUT2 #(
		.INIT('h8)
	) name4545 (
		_w15025_,
		_w15026_,
		_w15057_
	);
	LUT2 #(
		.INIT('h8)
	) name4546 (
		_w15023_,
		_w15024_,
		_w15058_
	);
	LUT2 #(
		.INIT('h8)
	) name4547 (
		_w15021_,
		_w15022_,
		_w15059_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		_w15019_,
		_w15020_,
		_w15060_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		_w15017_,
		_w15018_,
		_w15061_
	);
	LUT2 #(
		.INIT('h8)
	) name4550 (
		_w15015_,
		_w15016_,
		_w15062_
	);
	LUT2 #(
		.INIT('h8)
	) name4551 (
		_w15013_,
		_w15014_,
		_w15063_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		_w15011_,
		_w15012_,
		_w15064_
	);
	LUT2 #(
		.INIT('h8)
	) name4553 (
		_w15009_,
		_w15010_,
		_w15065_
	);
	LUT2 #(
		.INIT('h8)
	) name4554 (
		_w15007_,
		_w15008_,
		_w15066_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		_w15005_,
		_w15006_,
		_w15067_
	);
	LUT2 #(
		.INIT('h8)
	) name4556 (
		_w15003_,
		_w15004_,
		_w15068_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		_w15001_,
		_w15002_,
		_w15069_
	);
	LUT2 #(
		.INIT('h8)
	) name4558 (
		_w14999_,
		_w15000_,
		_w15070_
	);
	LUT2 #(
		.INIT('h8)
	) name4559 (
		_w14997_,
		_w14998_,
		_w15071_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		_w14995_,
		_w14996_,
		_w15072_
	);
	LUT2 #(
		.INIT('h8)
	) name4561 (
		_w14993_,
		_w14994_,
		_w15073_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		_w14991_,
		_w14992_,
		_w15074_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		_w14989_,
		_w14990_,
		_w15075_
	);
	LUT2 #(
		.INIT('h8)
	) name4564 (
		_w14987_,
		_w14988_,
		_w15076_
	);
	LUT2 #(
		.INIT('h8)
	) name4565 (
		_w14985_,
		_w14986_,
		_w15077_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		_w14983_,
		_w14984_,
		_w15078_
	);
	LUT2 #(
		.INIT('h8)
	) name4567 (
		_w15077_,
		_w15078_,
		_w15079_
	);
	LUT2 #(
		.INIT('h8)
	) name4568 (
		_w15075_,
		_w15076_,
		_w15080_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		_w15073_,
		_w15074_,
		_w15081_
	);
	LUT2 #(
		.INIT('h8)
	) name4570 (
		_w15071_,
		_w15072_,
		_w15082_
	);
	LUT2 #(
		.INIT('h8)
	) name4571 (
		_w15069_,
		_w15070_,
		_w15083_
	);
	LUT2 #(
		.INIT('h8)
	) name4572 (
		_w15067_,
		_w15068_,
		_w15084_
	);
	LUT2 #(
		.INIT('h8)
	) name4573 (
		_w15065_,
		_w15066_,
		_w15085_
	);
	LUT2 #(
		.INIT('h8)
	) name4574 (
		_w15063_,
		_w15064_,
		_w15086_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		_w15061_,
		_w15062_,
		_w15087_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		_w15059_,
		_w15060_,
		_w15088_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		_w15057_,
		_w15058_,
		_w15089_
	);
	LUT2 #(
		.INIT('h8)
	) name4578 (
		_w15055_,
		_w15056_,
		_w15090_
	);
	LUT2 #(
		.INIT('h8)
	) name4579 (
		_w15053_,
		_w15054_,
		_w15091_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		_w15051_,
		_w15052_,
		_w15092_
	);
	LUT2 #(
		.INIT('h8)
	) name4581 (
		_w15049_,
		_w15050_,
		_w15093_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		_w15047_,
		_w15048_,
		_w15094_
	);
	LUT2 #(
		.INIT('h8)
	) name4583 (
		_w15093_,
		_w15094_,
		_w15095_
	);
	LUT2 #(
		.INIT('h8)
	) name4584 (
		_w15091_,
		_w15092_,
		_w15096_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		_w15089_,
		_w15090_,
		_w15097_
	);
	LUT2 #(
		.INIT('h8)
	) name4586 (
		_w15087_,
		_w15088_,
		_w15098_
	);
	LUT2 #(
		.INIT('h8)
	) name4587 (
		_w15085_,
		_w15086_,
		_w15099_
	);
	LUT2 #(
		.INIT('h8)
	) name4588 (
		_w15083_,
		_w15084_,
		_w15100_
	);
	LUT2 #(
		.INIT('h8)
	) name4589 (
		_w15081_,
		_w15082_,
		_w15101_
	);
	LUT2 #(
		.INIT('h8)
	) name4590 (
		_w15079_,
		_w15080_,
		_w15102_
	);
	LUT2 #(
		.INIT('h8)
	) name4591 (
		_w15101_,
		_w15102_,
		_w15103_
	);
	LUT2 #(
		.INIT('h8)
	) name4592 (
		_w15099_,
		_w15100_,
		_w15104_
	);
	LUT2 #(
		.INIT('h8)
	) name4593 (
		_w15097_,
		_w15098_,
		_w15105_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		_w15095_,
		_w15096_,
		_w15106_
	);
	LUT2 #(
		.INIT('h8)
	) name4595 (
		_w15105_,
		_w15106_,
		_w15107_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		_w15103_,
		_w15104_,
		_w15108_
	);
	LUT2 #(
		.INIT('h8)
	) name4597 (
		_w15107_,
		_w15108_,
		_w15109_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		wb_rst_i_pad,
		_w15109_,
		_w15110_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		_w12656_,
		_w15110_,
		_w15111_
	);
	LUT2 #(
		.INIT('h4)
	) name4600 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		_w13483_,
		_w15112_
	);
	LUT2 #(
		.INIT('h4)
	) name4601 (
		_w13489_,
		_w15112_,
		_w15113_
	);
	LUT2 #(
		.INIT('h8)
	) name4602 (
		_w13500_,
		_w15113_,
		_w15114_
	);
	LUT2 #(
		.INIT('h1)
	) name4603 (
		\wishbone_TxLength_reg[8]/NET0131 ,
		_w15114_,
		_w15115_
	);
	LUT2 #(
		.INIT('h1)
	) name4604 (
		_w13499_,
		_w15113_,
		_w15116_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		\wishbone_TxLength_reg[8]/NET0131 ,
		_w12657_,
		_w15117_
	);
	LUT2 #(
		.INIT('h4)
	) name4606 (
		_w15116_,
		_w15117_,
		_w15118_
	);
	LUT2 #(
		.INIT('h1)
	) name4607 (
		_w12656_,
		_w15118_,
		_w15119_
	);
	LUT2 #(
		.INIT('h4)
	) name4608 (
		_w15115_,
		_w15119_,
		_w15120_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		_w15111_,
		_w15120_,
		_w15121_
	);
	LUT2 #(
		.INIT('h8)
	) name4610 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w12577_,
		_w15122_
	);
	LUT2 #(
		.INIT('h8)
	) name4611 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w12561_,
		_w15123_
	);
	LUT2 #(
		.INIT('h2)
	) name4612 (
		_w14591_,
		_w15123_,
		_w15124_
	);
	LUT2 #(
		.INIT('h8)
	) name4613 (
		_w12597_,
		_w12599_,
		_w15125_
	);
	LUT2 #(
		.INIT('h8)
	) name4614 (
		\m_wb_adr_o[25]_pad ,
		_w15125_,
		_w15126_
	);
	LUT2 #(
		.INIT('h1)
	) name4615 (
		\m_wb_adr_o[26]_pad ,
		_w15126_,
		_w15127_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w12602_,
		_w15124_,
		_w15128_
	);
	LUT2 #(
		.INIT('h4)
	) name4617 (
		_w15127_,
		_w15128_,
		_w15129_
	);
	LUT2 #(
		.INIT('h8)
	) name4618 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		_w12634_,
		_w15130_
	);
	LUT2 #(
		.INIT('h8)
	) name4619 (
		\m_wb_adr_o[26]_pad ,
		_w12636_,
		_w15131_
	);
	LUT2 #(
		.INIT('h1)
	) name4620 (
		_w15122_,
		_w15130_,
		_w15132_
	);
	LUT2 #(
		.INIT('h4)
	) name4621 (
		_w15131_,
		_w15132_,
		_w15133_
	);
	LUT2 #(
		.INIT('h4)
	) name4622 (
		_w15129_,
		_w15133_,
		_w15134_
	);
	LUT2 #(
		.INIT('h8)
	) name4623 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		_w15135_
	);
	LUT2 #(
		.INIT('h8)
	) name4624 (
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15135_,
		_w15136_
	);
	LUT2 #(
		.INIT('h8)
	) name4625 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w15136_,
		_w15137_
	);
	LUT2 #(
		.INIT('h8)
	) name4626 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w15138_
	);
	LUT2 #(
		.INIT('h8)
	) name4627 (
		\wishbone_RxReady_reg/NET0131 ,
		_w15138_,
		_w15139_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		_w15139_,
		_w15140_
	);
	LUT2 #(
		.INIT('h8)
	) name4629 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w15140_,
		_w15141_
	);
	LUT2 #(
		.INIT('h4)
	) name4630 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w15142_
	);
	LUT2 #(
		.INIT('h8)
	) name4631 (
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w15142_,
		_w15143_
	);
	LUT2 #(
		.INIT('h8)
	) name4632 (
		\wishbone_RxReady_reg/NET0131 ,
		_w15135_,
		_w15144_
	);
	LUT2 #(
		.INIT('h8)
	) name4633 (
		_w15143_,
		_w15144_,
		_w15145_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		_w15141_,
		_w15145_,
		_w15146_
	);
	LUT2 #(
		.INIT('h4)
	) name4635 (
		_w15137_,
		_w15146_,
		_w15147_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w15147_,
		_w15148_
	);
	LUT2 #(
		.INIT('h1)
	) name4637 (
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w15146_,
		_w15149_
	);
	LUT2 #(
		.INIT('h1)
	) name4638 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15150_
	);
	LUT2 #(
		.INIT('h8)
	) name4639 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w15151_
	);
	LUT2 #(
		.INIT('h1)
	) name4640 (
		_w15150_,
		_w15151_,
		_w15152_
	);
	LUT2 #(
		.INIT('h4)
	) name4641 (
		_w15149_,
		_w15152_,
		_w15153_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w15147_,
		_w15153_,
		_w15154_
	);
	LUT2 #(
		.INIT('h8)
	) name4643 (
		\wishbone_RxDataLatched1_reg[10]/NET0131 ,
		_w15154_,
		_w15155_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w15148_,
		_w15155_,
		_w15156_
	);
	LUT2 #(
		.INIT('h8)
	) name4645 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		_w15147_,
		_w15157_
	);
	LUT2 #(
		.INIT('h8)
	) name4646 (
		\wishbone_RxDataLatched1_reg[11]/NET0131 ,
		_w15154_,
		_w15158_
	);
	LUT2 #(
		.INIT('h1)
	) name4647 (
		_w15157_,
		_w15158_,
		_w15159_
	);
	LUT2 #(
		.INIT('h8)
	) name4648 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		_w15147_,
		_w15160_
	);
	LUT2 #(
		.INIT('h8)
	) name4649 (
		\wishbone_RxDataLatched1_reg[12]/NET0131 ,
		_w15154_,
		_w15161_
	);
	LUT2 #(
		.INIT('h1)
	) name4650 (
		_w15160_,
		_w15161_,
		_w15162_
	);
	LUT2 #(
		.INIT('h8)
	) name4651 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		_w15147_,
		_w15163_
	);
	LUT2 #(
		.INIT('h8)
	) name4652 (
		\wishbone_RxDataLatched1_reg[13]/NET0131 ,
		_w15154_,
		_w15164_
	);
	LUT2 #(
		.INIT('h1)
	) name4653 (
		_w15163_,
		_w15164_,
		_w15165_
	);
	LUT2 #(
		.INIT('h8)
	) name4654 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w15147_,
		_w15166_
	);
	LUT2 #(
		.INIT('h8)
	) name4655 (
		\wishbone_RxDataLatched1_reg[14]/NET0131 ,
		_w15154_,
		_w15167_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w15166_,
		_w15167_,
		_w15168_
	);
	LUT2 #(
		.INIT('h8)
	) name4657 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		_w15147_,
		_w15169_
	);
	LUT2 #(
		.INIT('h8)
	) name4658 (
		\wishbone_RxDataLatched1_reg[15]/NET0131 ,
		_w15154_,
		_w15170_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w15169_,
		_w15170_,
		_w15171_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		_w15147_,
		_w15172_
	);
	LUT2 #(
		.INIT('h8)
	) name4661 (
		\wishbone_RxDataLatched1_reg[8]/NET0131 ,
		_w15154_,
		_w15173_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w15172_,
		_w15173_,
		_w15174_
	);
	LUT2 #(
		.INIT('h8)
	) name4663 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_RxEn_reg/NET0131 ,
		_w15175_
	);
	LUT2 #(
		.INIT('h8)
	) name4664 (
		\wishbone_RxBDRead_reg/NET0131 ,
		_w15175_,
		_w15176_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		\wishbone_RxBDReady_reg/NET0131 ,
		_w15176_,
		_w15177_
	);
	LUT2 #(
		.INIT('h8)
	) name4666 (
		\wishbone_bd_ram_mem1_reg[156][15]/P0001 ,
		_w13190_,
		_w15178_
	);
	LUT2 #(
		.INIT('h8)
	) name4667 (
		\wishbone_bd_ram_mem1_reg[242][15]/P0001 ,
		_w12932_,
		_w15179_
	);
	LUT2 #(
		.INIT('h8)
	) name4668 (
		\wishbone_bd_ram_mem1_reg[199][15]/P0001 ,
		_w12768_,
		_w15180_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		\wishbone_bd_ram_mem1_reg[173][15]/P0001 ,
		_w12854_,
		_w15181_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		\wishbone_bd_ram_mem1_reg[212][15]/P0001 ,
		_w12796_,
		_w15182_
	);
	LUT2 #(
		.INIT('h8)
	) name4671 (
		\wishbone_bd_ram_mem1_reg[85][15]/P0001 ,
		_w13216_,
		_w15183_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		\wishbone_bd_ram_mem1_reg[120][15]/P0001 ,
		_w12707_,
		_w15184_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		\wishbone_bd_ram_mem1_reg[169][15]/P0001 ,
		_w12722_,
		_w15185_
	);
	LUT2 #(
		.INIT('h8)
	) name4674 (
		\wishbone_bd_ram_mem1_reg[191][15]/P0001 ,
		_w13034_,
		_w15186_
	);
	LUT2 #(
		.INIT('h8)
	) name4675 (
		\wishbone_bd_ram_mem1_reg[217][15]/P0001 ,
		_w13188_,
		_w15187_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		\wishbone_bd_ram_mem1_reg[108][15]/P0001 ,
		_w13156_,
		_w15188_
	);
	LUT2 #(
		.INIT('h8)
	) name4677 (
		\wishbone_bd_ram_mem1_reg[139][15]/P0001 ,
		_w12814_,
		_w15189_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		\wishbone_bd_ram_mem1_reg[197][15]/P0001 ,
		_w12834_,
		_w15190_
	);
	LUT2 #(
		.INIT('h8)
	) name4679 (
		\wishbone_bd_ram_mem1_reg[155][15]/P0001 ,
		_w13122_,
		_w15191_
	);
	LUT2 #(
		.INIT('h8)
	) name4680 (
		\wishbone_bd_ram_mem1_reg[164][15]/P0001 ,
		_w12876_,
		_w15192_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		\wishbone_bd_ram_mem1_reg[226][15]/P0001 ,
		_w13138_,
		_w15193_
	);
	LUT2 #(
		.INIT('h8)
	) name4682 (
		\wishbone_bd_ram_mem1_reg[80][15]/P0001 ,
		_w12689_,
		_w15194_
	);
	LUT2 #(
		.INIT('h8)
	) name4683 (
		\wishbone_bd_ram_mem1_reg[237][15]/P0001 ,
		_w12990_,
		_w15195_
	);
	LUT2 #(
		.INIT('h8)
	) name4684 (
		\wishbone_bd_ram_mem1_reg[235][15]/P0001 ,
		_w12696_,
		_w15196_
	);
	LUT2 #(
		.INIT('h8)
	) name4685 (
		\wishbone_bd_ram_mem1_reg[86][15]/P0001 ,
		_w12735_,
		_w15197_
	);
	LUT2 #(
		.INIT('h8)
	) name4686 (
		\wishbone_bd_ram_mem1_reg[203][15]/P0001 ,
		_w13158_,
		_w15198_
	);
	LUT2 #(
		.INIT('h8)
	) name4687 (
		\wishbone_bd_ram_mem1_reg[147][15]/P0001 ,
		_w13146_,
		_w15199_
	);
	LUT2 #(
		.INIT('h8)
	) name4688 (
		\wishbone_bd_ram_mem1_reg[1][15]/P0001 ,
		_w13014_,
		_w15200_
	);
	LUT2 #(
		.INIT('h8)
	) name4689 (
		\wishbone_bd_ram_mem1_reg[179][15]/P0001 ,
		_w13050_,
		_w15201_
	);
	LUT2 #(
		.INIT('h8)
	) name4690 (
		\wishbone_bd_ram_mem1_reg[45][15]/P0001 ,
		_w12908_,
		_w15202_
	);
	LUT2 #(
		.INIT('h8)
	) name4691 (
		\wishbone_bd_ram_mem1_reg[180][15]/P0001 ,
		_w12791_,
		_w15203_
	);
	LUT2 #(
		.INIT('h8)
	) name4692 (
		\wishbone_bd_ram_mem1_reg[68][15]/P0001 ,
		_w12946_,
		_w15204_
	);
	LUT2 #(
		.INIT('h8)
	) name4693 (
		\wishbone_bd_ram_mem1_reg[233][15]/P0001 ,
		_w12836_,
		_w15205_
	);
	LUT2 #(
		.INIT('h8)
	) name4694 (
		\wishbone_bd_ram_mem1_reg[138][15]/P0001 ,
		_w12958_,
		_w15206_
	);
	LUT2 #(
		.INIT('h8)
	) name4695 (
		\wishbone_bd_ram_mem1_reg[252][15]/P0001 ,
		_w13080_,
		_w15207_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		\wishbone_bd_ram_mem1_reg[22][15]/P0001 ,
		_w13110_,
		_w15208_
	);
	LUT2 #(
		.INIT('h8)
	) name4697 (
		\wishbone_bd_ram_mem1_reg[62][15]/P0001 ,
		_w12673_,
		_w15209_
	);
	LUT2 #(
		.INIT('h8)
	) name4698 (
		\wishbone_bd_ram_mem1_reg[188][15]/P0001 ,
		_w12948_,
		_w15210_
	);
	LUT2 #(
		.INIT('h8)
	) name4699 (
		\wishbone_bd_ram_mem1_reg[198][15]/P0001 ,
		_w12832_,
		_w15211_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		\wishbone_bd_ram_mem1_reg[249][15]/P0001 ,
		_w12900_,
		_w15212_
	);
	LUT2 #(
		.INIT('h8)
	) name4701 (
		\wishbone_bd_ram_mem1_reg[196][15]/P0001 ,
		_w13090_,
		_w15213_
	);
	LUT2 #(
		.INIT('h8)
	) name4702 (
		\wishbone_bd_ram_mem1_reg[88][15]/P0001 ,
		_w12860_,
		_w15214_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		\wishbone_bd_ram_mem1_reg[172][15]/P0001 ,
		_w12944_,
		_w15215_
	);
	LUT2 #(
		.INIT('h8)
	) name4704 (
		\wishbone_bd_ram_mem1_reg[129][15]/P0001 ,
		_w12776_,
		_w15216_
	);
	LUT2 #(
		.INIT('h8)
	) name4705 (
		\wishbone_bd_ram_mem1_reg[227][15]/P0001 ,
		_w12936_,
		_w15217_
	);
	LUT2 #(
		.INIT('h8)
	) name4706 (
		\wishbone_bd_ram_mem1_reg[18][15]/P0001 ,
		_w12679_,
		_w15218_
	);
	LUT2 #(
		.INIT('h8)
	) name4707 (
		\wishbone_bd_ram_mem1_reg[181][15]/P0001 ,
		_w12828_,
		_w15219_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		\wishbone_bd_ram_mem1_reg[20][15]/P0001 ,
		_w13174_,
		_w15220_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		\wishbone_bd_ram_mem1_reg[189][15]/P0001 ,
		_w13042_,
		_w15221_
	);
	LUT2 #(
		.INIT('h8)
	) name4710 (
		\wishbone_bd_ram_mem1_reg[67][15]/P0001 ,
		_w13134_,
		_w15222_
	);
	LUT2 #(
		.INIT('h8)
	) name4711 (
		\wishbone_bd_ram_mem1_reg[41][15]/P0001 ,
		_w13052_,
		_w15223_
	);
	LUT2 #(
		.INIT('h8)
	) name4712 (
		\wishbone_bd_ram_mem1_reg[122][15]/P0001 ,
		_w13130_,
		_w15224_
	);
	LUT2 #(
		.INIT('h8)
	) name4713 (
		\wishbone_bd_ram_mem1_reg[25][15]/P0001 ,
		_w13108_,
		_w15225_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		\wishbone_bd_ram_mem1_reg[52][15]/P0001 ,
		_w13082_,
		_w15226_
	);
	LUT2 #(
		.INIT('h8)
	) name4715 (
		\wishbone_bd_ram_mem1_reg[112][15]/P0001 ,
		_w12733_,
		_w15227_
	);
	LUT2 #(
		.INIT('h8)
	) name4716 (
		\wishbone_bd_ram_mem1_reg[255][15]/P0001 ,
		_w13072_,
		_w15228_
	);
	LUT2 #(
		.INIT('h8)
	) name4717 (
		\wishbone_bd_ram_mem1_reg[175][15]/P0001 ,
		_w13126_,
		_w15229_
	);
	LUT2 #(
		.INIT('h8)
	) name4718 (
		\wishbone_bd_ram_mem1_reg[73][15]/P0001 ,
		_w12918_,
		_w15230_
	);
	LUT2 #(
		.INIT('h8)
	) name4719 (
		\wishbone_bd_ram_mem1_reg[201][15]/P0001 ,
		_w12822_,
		_w15231_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		\wishbone_bd_ram_mem1_reg[37][15]/P0001 ,
		_w13102_,
		_w15232_
	);
	LUT2 #(
		.INIT('h8)
	) name4721 (
		\wishbone_bd_ram_mem1_reg[104][15]/P0001 ,
		_w13148_,
		_w15233_
	);
	LUT2 #(
		.INIT('h8)
	) name4722 (
		\wishbone_bd_ram_mem1_reg[27][15]/P0001 ,
		_w12880_,
		_w15234_
	);
	LUT2 #(
		.INIT('h8)
	) name4723 (
		\wishbone_bd_ram_mem1_reg[7][15]/P0001 ,
		_w12728_,
		_w15235_
	);
	LUT2 #(
		.INIT('h8)
	) name4724 (
		\wishbone_bd_ram_mem1_reg[150][15]/P0001 ,
		_w13136_,
		_w15236_
	);
	LUT2 #(
		.INIT('h8)
	) name4725 (
		\wishbone_bd_ram_mem1_reg[215][15]/P0001 ,
		_w12974_,
		_w15237_
	);
	LUT2 #(
		.INIT('h8)
	) name4726 (
		\wishbone_bd_ram_mem1_reg[238][15]/P0001 ,
		_w13160_,
		_w15238_
	);
	LUT2 #(
		.INIT('h8)
	) name4727 (
		\wishbone_bd_ram_mem1_reg[58][15]/P0001 ,
		_w13070_,
		_w15239_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		\wishbone_bd_ram_mem1_reg[195][15]/P0001 ,
		_w13144_,
		_w15240_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		\wishbone_bd_ram_mem1_reg[60][15]/P0001 ,
		_w13204_,
		_w15241_
	);
	LUT2 #(
		.INIT('h8)
	) name4730 (
		\wishbone_bd_ram_mem1_reg[15][15]/P0001 ,
		_w13210_,
		_w15242_
	);
	LUT2 #(
		.INIT('h8)
	) name4731 (
		\wishbone_bd_ram_mem1_reg[26][15]/P0001 ,
		_w12699_,
		_w15243_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		\wishbone_bd_ram_mem1_reg[97][15]/P0001 ,
		_w13096_,
		_w15244_
	);
	LUT2 #(
		.INIT('h8)
	) name4733 (
		\wishbone_bd_ram_mem1_reg[160][15]/P0001 ,
		_w12872_,
		_w15245_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		\wishbone_bd_ram_mem1_reg[47][15]/P0001 ,
		_w12904_,
		_w15246_
	);
	LUT2 #(
		.INIT('h8)
	) name4735 (
		\wishbone_bd_ram_mem1_reg[21][15]/P0001 ,
		_w12906_,
		_w15247_
	);
	LUT2 #(
		.INIT('h8)
	) name4736 (
		\wishbone_bd_ram_mem1_reg[77][15]/P0001 ,
		_w12982_,
		_w15248_
	);
	LUT2 #(
		.INIT('h8)
	) name4737 (
		\wishbone_bd_ram_mem1_reg[206][15]/P0001 ,
		_w12954_,
		_w15249_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		\wishbone_bd_ram_mem1_reg[153][15]/P0001 ,
		_w12890_,
		_w15250_
	);
	LUT2 #(
		.INIT('h8)
	) name4739 (
		\wishbone_bd_ram_mem1_reg[98][15]/P0001 ,
		_w12816_,
		_w15251_
	);
	LUT2 #(
		.INIT('h8)
	) name4740 (
		\wishbone_bd_ram_mem1_reg[192][15]/P0001 ,
		_w12938_,
		_w15252_
	);
	LUT2 #(
		.INIT('h8)
	) name4741 (
		\wishbone_bd_ram_mem1_reg[142][15]/P0001 ,
		_w12928_,
		_w15253_
	);
	LUT2 #(
		.INIT('h8)
	) name4742 (
		\wishbone_bd_ram_mem1_reg[4][15]/P0001 ,
		_w12666_,
		_w15254_
	);
	LUT2 #(
		.INIT('h8)
	) name4743 (
		\wishbone_bd_ram_mem1_reg[117][15]/P0001 ,
		_w12715_,
		_w15255_
	);
	LUT2 #(
		.INIT('h8)
	) name4744 (
		\wishbone_bd_ram_mem1_reg[152][15]/P0001 ,
		_w12966_,
		_w15256_
	);
	LUT2 #(
		.INIT('h8)
	) name4745 (
		\wishbone_bd_ram_mem1_reg[103][15]/P0001 ,
		_w12846_,
		_w15257_
	);
	LUT2 #(
		.INIT('h8)
	) name4746 (
		\wishbone_bd_ram_mem1_reg[234][15]/P0001 ,
		_w13214_,
		_w15258_
	);
	LUT2 #(
		.INIT('h8)
	) name4747 (
		\wishbone_bd_ram_mem1_reg[162][15]/P0001 ,
		_w13098_,
		_w15259_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		\wishbone_bd_ram_mem1_reg[145][15]/P0001 ,
		_w13106_,
		_w15260_
	);
	LUT2 #(
		.INIT('h8)
	) name4749 (
		\wishbone_bd_ram_mem1_reg[72][15]/P0001 ,
		_w12810_,
		_w15261_
	);
	LUT2 #(
		.INIT('h8)
	) name4750 (
		\wishbone_bd_ram_mem1_reg[44][15]/P0001 ,
		_w12896_,
		_w15262_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		\wishbone_bd_ram_mem1_reg[243][15]/P0001 ,
		_w12804_,
		_w15263_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		\wishbone_bd_ram_mem1_reg[118][15]/P0001 ,
		_w12830_,
		_w15264_
	);
	LUT2 #(
		.INIT('h8)
	) name4753 (
		\wishbone_bd_ram_mem1_reg[193][15]/P0001 ,
		_w13056_,
		_w15265_
	);
	LUT2 #(
		.INIT('h8)
	) name4754 (
		\wishbone_bd_ram_mem1_reg[132][15]/P0001 ,
		_w12992_,
		_w15266_
	);
	LUT2 #(
		.INIT('h8)
	) name4755 (
		\wishbone_bd_ram_mem1_reg[83][15]/P0001 ,
		_w12916_,
		_w15267_
	);
	LUT2 #(
		.INIT('h8)
	) name4756 (
		\wishbone_bd_ram_mem1_reg[167][15]/P0001 ,
		_w12986_,
		_w15268_
	);
	LUT2 #(
		.INIT('h8)
	) name4757 (
		\wishbone_bd_ram_mem1_reg[151][15]/P0001 ,
		_w13142_,
		_w15269_
	);
	LUT2 #(
		.INIT('h8)
	) name4758 (
		\wishbone_bd_ram_mem1_reg[105][15]/P0001 ,
		_w12751_,
		_w15270_
	);
	LUT2 #(
		.INIT('h8)
	) name4759 (
		\wishbone_bd_ram_mem1_reg[141][15]/P0001 ,
		_w13004_,
		_w15271_
	);
	LUT2 #(
		.INIT('h8)
	) name4760 (
		\wishbone_bd_ram_mem1_reg[149][15]/P0001 ,
		_w12741_,
		_w15272_
	);
	LUT2 #(
		.INIT('h8)
	) name4761 (
		\wishbone_bd_ram_mem1_reg[194][15]/P0001 ,
		_w12772_,
		_w15273_
	);
	LUT2 #(
		.INIT('h8)
	) name4762 (
		\wishbone_bd_ram_mem1_reg[109][15]/P0001 ,
		_w12888_,
		_w15274_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		\wishbone_bd_ram_mem1_reg[42][15]/P0001 ,
		_w12842_,
		_w15275_
	);
	LUT2 #(
		.INIT('h8)
	) name4764 (
		\wishbone_bd_ram_mem1_reg[144][15]/P0001 ,
		_w12756_,
		_w15276_
	);
	LUT2 #(
		.INIT('h8)
	) name4765 (
		\wishbone_bd_ram_mem1_reg[166][15]/P0001 ,
		_w13040_,
		_w15277_
	);
	LUT2 #(
		.INIT('h8)
	) name4766 (
		\wishbone_bd_ram_mem1_reg[218][15]/P0001 ,
		_w13206_,
		_w15278_
	);
	LUT2 #(
		.INIT('h8)
	) name4767 (
		\wishbone_bd_ram_mem1_reg[90][15]/P0001 ,
		_w12978_,
		_w15279_
	);
	LUT2 #(
		.INIT('h8)
	) name4768 (
		\wishbone_bd_ram_mem1_reg[126][15]/P0001 ,
		_w13218_,
		_w15280_
	);
	LUT2 #(
		.INIT('h8)
	) name4769 (
		\wishbone_bd_ram_mem1_reg[119][15]/P0001 ,
		_w13048_,
		_w15281_
	);
	LUT2 #(
		.INIT('h8)
	) name4770 (
		\wishbone_bd_ram_mem1_reg[240][15]/P0001 ,
		_w12864_,
		_w15282_
	);
	LUT2 #(
		.INIT('h8)
	) name4771 (
		\wishbone_bd_ram_mem1_reg[76][15]/P0001 ,
		_w13184_,
		_w15283_
	);
	LUT2 #(
		.INIT('h8)
	) name4772 (
		\wishbone_bd_ram_mem1_reg[84][15]/P0001 ,
		_w12934_,
		_w15284_
	);
	LUT2 #(
		.INIT('h8)
	) name4773 (
		\wishbone_bd_ram_mem1_reg[177][15]/P0001 ,
		_w12996_,
		_w15285_
	);
	LUT2 #(
		.INIT('h8)
	) name4774 (
		\wishbone_bd_ram_mem1_reg[123][15]/P0001 ,
		_w13114_,
		_w15286_
	);
	LUT2 #(
		.INIT('h8)
	) name4775 (
		\wishbone_bd_ram_mem1_reg[247][15]/P0001 ,
		_w12818_,
		_w15287_
	);
	LUT2 #(
		.INIT('h8)
	) name4776 (
		\wishbone_bd_ram_mem1_reg[133][15]/P0001 ,
		_w12761_,
		_w15288_
	);
	LUT2 #(
		.INIT('h8)
	) name4777 (
		\wishbone_bd_ram_mem1_reg[49][15]/P0001 ,
		_w12994_,
		_w15289_
	);
	LUT2 #(
		.INIT('h8)
	) name4778 (
		\wishbone_bd_ram_mem1_reg[29][15]/P0001 ,
		_w12952_,
		_w15290_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		\wishbone_bd_ram_mem1_reg[39][15]/P0001 ,
		_w13018_,
		_w15291_
	);
	LUT2 #(
		.INIT('h8)
	) name4780 (
		\wishbone_bd_ram_mem1_reg[134][15]/P0001 ,
		_w12763_,
		_w15292_
	);
	LUT2 #(
		.INIT('h8)
	) name4781 (
		\wishbone_bd_ram_mem1_reg[43][15]/P0001 ,
		_w13200_,
		_w15293_
	);
	LUT2 #(
		.INIT('h8)
	) name4782 (
		\wishbone_bd_ram_mem1_reg[50][15]/P0001 ,
		_w13150_,
		_w15294_
	);
	LUT2 #(
		.INIT('h8)
	) name4783 (
		\wishbone_bd_ram_mem1_reg[213][15]/P0001 ,
		_w13002_,
		_w15295_
	);
	LUT2 #(
		.INIT('h8)
	) name4784 (
		\wishbone_bd_ram_mem1_reg[32][15]/P0001 ,
		_w13120_,
		_w15296_
	);
	LUT2 #(
		.INIT('h8)
	) name4785 (
		\wishbone_bd_ram_mem1_reg[182][15]/P0001 ,
		_w12820_,
		_w15297_
	);
	LUT2 #(
		.INIT('h8)
	) name4786 (
		\wishbone_bd_ram_mem1_reg[163][15]/P0001 ,
		_w12882_,
		_w15298_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		\wishbone_bd_ram_mem1_reg[75][15]/P0001 ,
		_w12826_,
		_w15299_
	);
	LUT2 #(
		.INIT('h8)
	) name4788 (
		\wishbone_bd_ram_mem1_reg[9][15]/P0001 ,
		_w12808_,
		_w15300_
	);
	LUT2 #(
		.INIT('h8)
	) name4789 (
		\wishbone_bd_ram_mem1_reg[14][15]/P0001 ,
		_w13086_,
		_w15301_
	);
	LUT2 #(
		.INIT('h8)
	) name4790 (
		\wishbone_bd_ram_mem1_reg[13][15]/P0001 ,
		_w13178_,
		_w15302_
	);
	LUT2 #(
		.INIT('h8)
	) name4791 (
		\wishbone_bd_ram_mem1_reg[46][15]/P0001 ,
		_w12884_,
		_w15303_
	);
	LUT2 #(
		.INIT('h8)
	) name4792 (
		\wishbone_bd_ram_mem1_reg[101][15]/P0001 ,
		_w13192_,
		_w15304_
	);
	LUT2 #(
		.INIT('h8)
	) name4793 (
		\wishbone_bd_ram_mem1_reg[202][15]/P0001 ,
		_w12870_,
		_w15305_
	);
	LUT2 #(
		.INIT('h8)
	) name4794 (
		\wishbone_bd_ram_mem1_reg[78][15]/P0001 ,
		_w12874_,
		_w15306_
	);
	LUT2 #(
		.INIT('h8)
	) name4795 (
		\wishbone_bd_ram_mem1_reg[178][15]/P0001 ,
		_w12886_,
		_w15307_
	);
	LUT2 #(
		.INIT('h8)
	) name4796 (
		\wishbone_bd_ram_mem1_reg[219][15]/P0001 ,
		_w12806_,
		_w15308_
	);
	LUT2 #(
		.INIT('h8)
	) name4797 (
		\wishbone_bd_ram_mem1_reg[187][15]/P0001 ,
		_w13196_,
		_w15309_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		\wishbone_bd_ram_mem1_reg[171][15]/P0001 ,
		_w12910_,
		_w15310_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		\wishbone_bd_ram_mem1_reg[91][15]/P0001 ,
		_w13074_,
		_w15311_
	);
	LUT2 #(
		.INIT('h8)
	) name4800 (
		\wishbone_bd_ram_mem1_reg[33][15]/P0001 ,
		_w12980_,
		_w15312_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		\wishbone_bd_ram_mem1_reg[174][15]/P0001 ,
		_w12972_,
		_w15313_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		\wishbone_bd_ram_mem1_reg[61][15]/P0001 ,
		_w12725_,
		_w15314_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		\wishbone_bd_ram_mem1_reg[64][15]/P0001 ,
		_w12976_,
		_w15315_
	);
	LUT2 #(
		.INIT('h8)
	) name4804 (
		\wishbone_bd_ram_mem1_reg[111][15]/P0001 ,
		_w12744_,
		_w15316_
	);
	LUT2 #(
		.INIT('h8)
	) name4805 (
		\wishbone_bd_ram_mem1_reg[222][15]/P0001 ,
		_w13094_,
		_w15317_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		\wishbone_bd_ram_mem1_reg[170][15]/P0001 ,
		_w13030_,
		_w15318_
	);
	LUT2 #(
		.INIT('h8)
	) name4807 (
		\wishbone_bd_ram_mem1_reg[241][15]/P0001 ,
		_w13006_,
		_w15319_
	);
	LUT2 #(
		.INIT('h8)
	) name4808 (
		\wishbone_bd_ram_mem1_reg[115][15]/P0001 ,
		_w13112_,
		_w15320_
	);
	LUT2 #(
		.INIT('h8)
	) name4809 (
		\wishbone_bd_ram_mem1_reg[24][15]/P0001 ,
		_w13084_,
		_w15321_
	);
	LUT2 #(
		.INIT('h8)
	) name4810 (
		\wishbone_bd_ram_mem1_reg[125][15]/P0001 ,
		_w12956_,
		_w15322_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		\wishbone_bd_ram_mem1_reg[28][15]/P0001 ,
		_w13170_,
		_w15323_
	);
	LUT2 #(
		.INIT('h8)
	) name4812 (
		\wishbone_bd_ram_mem1_reg[127][15]/P0001 ,
		_w13164_,
		_w15324_
	);
	LUT2 #(
		.INIT('h8)
	) name4813 (
		\wishbone_bd_ram_mem1_reg[74][15]/P0001 ,
		_w12812_,
		_w15325_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		\wishbone_bd_ram_mem1_reg[130][15]/P0001 ,
		_w12914_,
		_w15326_
	);
	LUT2 #(
		.INIT('h8)
	) name4815 (
		\wishbone_bd_ram_mem1_reg[48][15]/P0001 ,
		_w12970_,
		_w15327_
	);
	LUT2 #(
		.INIT('h8)
	) name4816 (
		\wishbone_bd_ram_mem1_reg[207][15]/P0001 ,
		_w13180_,
		_w15328_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		\wishbone_bd_ram_mem1_reg[71][15]/P0001 ,
		_w12798_,
		_w15329_
	);
	LUT2 #(
		.INIT('h8)
	) name4818 (
		\wishbone_bd_ram_mem1_reg[11][15]/P0001 ,
		_w13194_,
		_w15330_
	);
	LUT2 #(
		.INIT('h8)
	) name4819 (
		\wishbone_bd_ram_mem1_reg[106][15]/P0001 ,
		_w12713_,
		_w15331_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		\wishbone_bd_ram_mem1_reg[251][15]/P0001 ,
		_w13054_,
		_w15332_
	);
	LUT2 #(
		.INIT('h8)
	) name4821 (
		\wishbone_bd_ram_mem1_reg[204][15]/P0001 ,
		_w13162_,
		_w15333_
	);
	LUT2 #(
		.INIT('h8)
	) name4822 (
		\wishbone_bd_ram_mem1_reg[31][15]/P0001 ,
		_w13198_,
		_w15334_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		\wishbone_bd_ram_mem1_reg[82][15]/P0001 ,
		_w12942_,
		_w15335_
	);
	LUT2 #(
		.INIT('h8)
	) name4824 (
		\wishbone_bd_ram_mem1_reg[137][15]/P0001 ,
		_w13168_,
		_w15336_
	);
	LUT2 #(
		.INIT('h8)
	) name4825 (
		\wishbone_bd_ram_mem1_reg[200][15]/P0001 ,
		_w12988_,
		_w15337_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\wishbone_bd_ram_mem1_reg[246][15]/P0001 ,
		_w13076_,
		_w15338_
	);
	LUT2 #(
		.INIT('h8)
	) name4827 (
		\wishbone_bd_ram_mem1_reg[205][15]/P0001 ,
		_w13068_,
		_w15339_
	);
	LUT2 #(
		.INIT('h8)
	) name4828 (
		\wishbone_bd_ram_mem1_reg[210][15]/P0001 ,
		_w12924_,
		_w15340_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		\wishbone_bd_ram_mem1_reg[0][15]/P0001 ,
		_w12717_,
		_w15341_
	);
	LUT2 #(
		.INIT('h8)
	) name4830 (
		\wishbone_bd_ram_mem1_reg[211][15]/P0001 ,
		_w13166_,
		_w15342_
	);
	LUT2 #(
		.INIT('h8)
	) name4831 (
		\wishbone_bd_ram_mem1_reg[165][15]/P0001 ,
		_w13044_,
		_w15343_
	);
	LUT2 #(
		.INIT('h8)
	) name4832 (
		\wishbone_bd_ram_mem1_reg[131][15]/P0001 ,
		_w12852_,
		_w15344_
	);
	LUT2 #(
		.INIT('h8)
	) name4833 (
		\wishbone_bd_ram_mem1_reg[107][15]/P0001 ,
		_w12749_,
		_w15345_
	);
	LUT2 #(
		.INIT('h8)
	) name4834 (
		\wishbone_bd_ram_mem1_reg[66][15]/P0001 ,
		_w12824_,
		_w15346_
	);
	LUT2 #(
		.INIT('h8)
	) name4835 (
		\wishbone_bd_ram_mem1_reg[35][15]/P0001 ,
		_w12703_,
		_w15347_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		\wishbone_bd_ram_mem1_reg[40][15]/P0001 ,
		_w13132_,
		_w15348_
	);
	LUT2 #(
		.INIT('h8)
	) name4837 (
		\wishbone_bd_ram_mem1_reg[143][15]/P0001 ,
		_w12922_,
		_w15349_
	);
	LUT2 #(
		.INIT('h8)
	) name4838 (
		\wishbone_bd_ram_mem1_reg[99][15]/P0001 ,
		_w13038_,
		_w15350_
	);
	LUT2 #(
		.INIT('h8)
	) name4839 (
		\wishbone_bd_ram_mem1_reg[168][15]/P0001 ,
		_w13208_,
		_w15351_
	);
	LUT2 #(
		.INIT('h8)
	) name4840 (
		\wishbone_bd_ram_mem1_reg[36][15]/P0001 ,
		_w12800_,
		_w15352_
	);
	LUT2 #(
		.INIT('h8)
	) name4841 (
		\wishbone_bd_ram_mem1_reg[214][15]/P0001 ,
		_w12984_,
		_w15353_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		\wishbone_bd_ram_mem1_reg[128][15]/P0001 ,
		_w12793_,
		_w15354_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		\wishbone_bd_ram_mem1_reg[124][15]/P0001 ,
		_w13058_,
		_w15355_
	);
	LUT2 #(
		.INIT('h8)
	) name4844 (
		\wishbone_bd_ram_mem1_reg[239][15]/P0001 ,
		_w12862_,
		_w15356_
	);
	LUT2 #(
		.INIT('h8)
	) name4845 (
		\wishbone_bd_ram_mem1_reg[17][15]/P0001 ,
		_w12848_,
		_w15357_
	);
	LUT2 #(
		.INIT('h8)
	) name4846 (
		\wishbone_bd_ram_mem1_reg[220][15]/P0001 ,
		_w13066_,
		_w15358_
	);
	LUT2 #(
		.INIT('h8)
	) name4847 (
		\wishbone_bd_ram_mem1_reg[95][15]/P0001 ,
		_w12844_,
		_w15359_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		\wishbone_bd_ram_mem1_reg[16][15]/P0001 ,
		_w13140_,
		_w15360_
	);
	LUT2 #(
		.INIT('h8)
	) name4849 (
		\wishbone_bd_ram_mem1_reg[81][15]/P0001 ,
		_w12950_,
		_w15361_
	);
	LUT2 #(
		.INIT('h8)
	) name4850 (
		\wishbone_bd_ram_mem1_reg[221][15]/P0001 ,
		_w12802_,
		_w15362_
	);
	LUT2 #(
		.INIT('h8)
	) name4851 (
		\wishbone_bd_ram_mem1_reg[30][15]/P0001 ,
		_w13104_,
		_w15363_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		\wishbone_bd_ram_mem1_reg[116][15]/P0001 ,
		_w12998_,
		_w15364_
	);
	LUT2 #(
		.INIT('h8)
	) name4853 (
		\wishbone_bd_ram_mem1_reg[224][15]/P0001 ,
		_w12902_,
		_w15365_
	);
	LUT2 #(
		.INIT('h8)
	) name4854 (
		\wishbone_bd_ram_mem1_reg[244][15]/P0001 ,
		_w12747_,
		_w15366_
	);
	LUT2 #(
		.INIT('h8)
	) name4855 (
		\wishbone_bd_ram_mem1_reg[87][15]/P0001 ,
		_w13154_,
		_w15367_
	);
	LUT2 #(
		.INIT('h8)
	) name4856 (
		\wishbone_bd_ram_mem1_reg[140][15]/P0001 ,
		_w12894_,
		_w15368_
	);
	LUT2 #(
		.INIT('h8)
	) name4857 (
		\wishbone_bd_ram_mem1_reg[158][15]/P0001 ,
		_w12898_,
		_w15369_
	);
	LUT2 #(
		.INIT('h8)
	) name4858 (
		\wishbone_bd_ram_mem1_reg[23][15]/P0001 ,
		_w13008_,
		_w15370_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		\wishbone_bd_ram_mem1_reg[208][15]/P0001 ,
		_w13032_,
		_w15371_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		\wishbone_bd_ram_mem1_reg[54][15]/P0001 ,
		_w12770_,
		_w15372_
	);
	LUT2 #(
		.INIT('h8)
	) name4861 (
		\wishbone_bd_ram_mem1_reg[248][15]/P0001 ,
		_w12789_,
		_w15373_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		\wishbone_bd_ram_mem1_reg[159][15]/P0001 ,
		_w12774_,
		_w15374_
	);
	LUT2 #(
		.INIT('h8)
	) name4863 (
		\wishbone_bd_ram_mem1_reg[56][15]/P0001 ,
		_w12778_,
		_w15375_
	);
	LUT2 #(
		.INIT('h8)
	) name4864 (
		\wishbone_bd_ram_mem1_reg[12][15]/P0001 ,
		_w13118_,
		_w15376_
	);
	LUT2 #(
		.INIT('h8)
	) name4865 (
		\wishbone_bd_ram_mem1_reg[161][15]/P0001 ,
		_w12754_,
		_w15377_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		\wishbone_bd_ram_mem1_reg[92][15]/P0001 ,
		_w13010_,
		_w15378_
	);
	LUT2 #(
		.INIT('h8)
	) name4867 (
		\wishbone_bd_ram_mem1_reg[186][15]/P0001 ,
		_w12783_,
		_w15379_
	);
	LUT2 #(
		.INIT('h8)
	) name4868 (
		\wishbone_bd_ram_mem1_reg[19][15]/P0001 ,
		_w13012_,
		_w15380_
	);
	LUT2 #(
		.INIT('h8)
	) name4869 (
		\wishbone_bd_ram_mem1_reg[232][15]/P0001 ,
		_w12758_,
		_w15381_
	);
	LUT2 #(
		.INIT('h8)
	) name4870 (
		\wishbone_bd_ram_mem1_reg[135][15]/P0001 ,
		_w13124_,
		_w15382_
	);
	LUT2 #(
		.INIT('h8)
	) name4871 (
		\wishbone_bd_ram_mem1_reg[2][15]/P0001 ,
		_w13088_,
		_w15383_
	);
	LUT2 #(
		.INIT('h8)
	) name4872 (
		\wishbone_bd_ram_mem1_reg[184][15]/P0001 ,
		_w13062_,
		_w15384_
	);
	LUT2 #(
		.INIT('h8)
	) name4873 (
		\wishbone_bd_ram_mem1_reg[154][15]/P0001 ,
		_w12962_,
		_w15385_
	);
	LUT2 #(
		.INIT('h8)
	) name4874 (
		\wishbone_bd_ram_mem1_reg[223][15]/P0001 ,
		_w12838_,
		_w15386_
	);
	LUT2 #(
		.INIT('h8)
	) name4875 (
		\wishbone_bd_ram_mem1_reg[89][15]/P0001 ,
		_w12964_,
		_w15387_
	);
	LUT2 #(
		.INIT('h8)
	) name4876 (
		\wishbone_bd_ram_mem1_reg[6][15]/P0001 ,
		_w12968_,
		_w15388_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		\wishbone_bd_ram_mem1_reg[70][15]/P0001 ,
		_w12840_,
		_w15389_
	);
	LUT2 #(
		.INIT('h8)
	) name4878 (
		\wishbone_bd_ram_mem1_reg[121][15]/P0001 ,
		_w13078_,
		_w15390_
	);
	LUT2 #(
		.INIT('h8)
	) name4879 (
		\wishbone_bd_ram_mem1_reg[65][15]/P0001 ,
		_w13176_,
		_w15391_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		\wishbone_bd_ram_mem1_reg[229][15]/P0001 ,
		_w12711_,
		_w15392_
	);
	LUT2 #(
		.INIT('h8)
	) name4881 (
		\wishbone_bd_ram_mem1_reg[100][15]/P0001 ,
		_w12960_,
		_w15393_
	);
	LUT2 #(
		.INIT('h8)
	) name4882 (
		\wishbone_bd_ram_mem1_reg[183][15]/P0001 ,
		_w12787_,
		_w15394_
	);
	LUT2 #(
		.INIT('h8)
	) name4883 (
		\wishbone_bd_ram_mem1_reg[96][15]/P0001 ,
		_w12912_,
		_w15395_
	);
	LUT2 #(
		.INIT('h8)
	) name4884 (
		\wishbone_bd_ram_mem1_reg[228][15]/P0001 ,
		_w12765_,
		_w15396_
	);
	LUT2 #(
		.INIT('h8)
	) name4885 (
		\wishbone_bd_ram_mem1_reg[59][15]/P0001 ,
		_w12780_,
		_w15397_
	);
	LUT2 #(
		.INIT('h8)
	) name4886 (
		\wishbone_bd_ram_mem1_reg[38][15]/P0001 ,
		_w13182_,
		_w15398_
	);
	LUT2 #(
		.INIT('h8)
	) name4887 (
		\wishbone_bd_ram_mem1_reg[34][15]/P0001 ,
		_w12930_,
		_w15399_
	);
	LUT2 #(
		.INIT('h8)
	) name4888 (
		\wishbone_bd_ram_mem1_reg[3][15]/P0001 ,
		_w12866_,
		_w15400_
	);
	LUT2 #(
		.INIT('h8)
	) name4889 (
		\wishbone_bd_ram_mem1_reg[63][15]/P0001 ,
		_w12850_,
		_w15401_
	);
	LUT2 #(
		.INIT('h8)
	) name4890 (
		\wishbone_bd_ram_mem1_reg[231][15]/P0001 ,
		_w12856_,
		_w15402_
	);
	LUT2 #(
		.INIT('h8)
	) name4891 (
		\wishbone_bd_ram_mem1_reg[209][15]/P0001 ,
		_w13152_,
		_w15403_
	);
	LUT2 #(
		.INIT('h8)
	) name4892 (
		\wishbone_bd_ram_mem1_reg[216][15]/P0001 ,
		_w13028_,
		_w15404_
	);
	LUT2 #(
		.INIT('h8)
	) name4893 (
		\wishbone_bd_ram_mem1_reg[8][15]/P0001 ,
		_w12920_,
		_w15405_
	);
	LUT2 #(
		.INIT('h8)
	) name4894 (
		\wishbone_bd_ram_mem1_reg[79][15]/P0001 ,
		_w13212_,
		_w15406_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		\wishbone_bd_ram_mem1_reg[5][15]/P0001 ,
		_w12878_,
		_w15407_
	);
	LUT2 #(
		.INIT('h8)
	) name4896 (
		\wishbone_bd_ram_mem1_reg[53][15]/P0001 ,
		_w13020_,
		_w15408_
	);
	LUT2 #(
		.INIT('h8)
	) name4897 (
		\wishbone_bd_ram_mem1_reg[225][15]/P0001 ,
		_w13092_,
		_w15409_
	);
	LUT2 #(
		.INIT('h8)
	) name4898 (
		\wishbone_bd_ram_mem1_reg[110][15]/P0001 ,
		_w13046_,
		_w15410_
	);
	LUT2 #(
		.INIT('h8)
	) name4899 (
		\wishbone_bd_ram_mem1_reg[230][15]/P0001 ,
		_w13036_,
		_w15411_
	);
	LUT2 #(
		.INIT('h8)
	) name4900 (
		\wishbone_bd_ram_mem1_reg[69][15]/P0001 ,
		_w12738_,
		_w15412_
	);
	LUT2 #(
		.INIT('h8)
	) name4901 (
		\wishbone_bd_ram_mem1_reg[146][15]/P0001 ,
		_w13060_,
		_w15413_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		\wishbone_bd_ram_mem1_reg[55][15]/P0001 ,
		_w12785_,
		_w15414_
	);
	LUT2 #(
		.INIT('h8)
	) name4903 (
		\wishbone_bd_ram_mem1_reg[157][15]/P0001 ,
		_w12926_,
		_w15415_
	);
	LUT2 #(
		.INIT('h8)
	) name4904 (
		\wishbone_bd_ram_mem1_reg[93][15]/P0001 ,
		_w13016_,
		_w15416_
	);
	LUT2 #(
		.INIT('h8)
	) name4905 (
		\wishbone_bd_ram_mem1_reg[176][15]/P0001 ,
		_w12868_,
		_w15417_
	);
	LUT2 #(
		.INIT('h8)
	) name4906 (
		\wishbone_bd_ram_mem1_reg[10][15]/P0001 ,
		_w13172_,
		_w15418_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		\wishbone_bd_ram_mem1_reg[102][15]/P0001 ,
		_w12685_,
		_w15419_
	);
	LUT2 #(
		.INIT('h8)
	) name4908 (
		\wishbone_bd_ram_mem1_reg[136][15]/P0001 ,
		_w13064_,
		_w15420_
	);
	LUT2 #(
		.INIT('h8)
	) name4909 (
		\wishbone_bd_ram_mem1_reg[190][15]/P0001 ,
		_w12858_,
		_w15421_
	);
	LUT2 #(
		.INIT('h8)
	) name4910 (
		\wishbone_bd_ram_mem1_reg[51][15]/P0001 ,
		_w13024_,
		_w15422_
	);
	LUT2 #(
		.INIT('h8)
	) name4911 (
		\wishbone_bd_ram_mem1_reg[250][15]/P0001 ,
		_w13128_,
		_w15423_
	);
	LUT2 #(
		.INIT('h8)
	) name4912 (
		\wishbone_bd_ram_mem1_reg[185][15]/P0001 ,
		_w12940_,
		_w15424_
	);
	LUT2 #(
		.INIT('h8)
	) name4913 (
		\wishbone_bd_ram_mem1_reg[148][15]/P0001 ,
		_w13000_,
		_w15425_
	);
	LUT2 #(
		.INIT('h8)
	) name4914 (
		\wishbone_bd_ram_mem1_reg[57][15]/P0001 ,
		_w13116_,
		_w15426_
	);
	LUT2 #(
		.INIT('h8)
	) name4915 (
		\wishbone_bd_ram_mem1_reg[254][15]/P0001 ,
		_w12892_,
		_w15427_
	);
	LUT2 #(
		.INIT('h8)
	) name4916 (
		\wishbone_bd_ram_mem1_reg[245][15]/P0001 ,
		_w13022_,
		_w15428_
	);
	LUT2 #(
		.INIT('h8)
	) name4917 (
		\wishbone_bd_ram_mem1_reg[253][15]/P0001 ,
		_w13100_,
		_w15429_
	);
	LUT2 #(
		.INIT('h8)
	) name4918 (
		\wishbone_bd_ram_mem1_reg[114][15]/P0001 ,
		_w13202_,
		_w15430_
	);
	LUT2 #(
		.INIT('h8)
	) name4919 (
		\wishbone_bd_ram_mem1_reg[94][15]/P0001 ,
		_w13186_,
		_w15431_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		\wishbone_bd_ram_mem1_reg[236][15]/P0001 ,
		_w12731_,
		_w15432_
	);
	LUT2 #(
		.INIT('h8)
	) name4921 (
		\wishbone_bd_ram_mem1_reg[113][15]/P0001 ,
		_w13026_,
		_w15433_
	);
	LUT2 #(
		.INIT('h1)
	) name4922 (
		_w15178_,
		_w15179_,
		_w15434_
	);
	LUT2 #(
		.INIT('h1)
	) name4923 (
		_w15180_,
		_w15181_,
		_w15435_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w15182_,
		_w15183_,
		_w15436_
	);
	LUT2 #(
		.INIT('h1)
	) name4925 (
		_w15184_,
		_w15185_,
		_w15437_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w15186_,
		_w15187_,
		_w15438_
	);
	LUT2 #(
		.INIT('h1)
	) name4927 (
		_w15188_,
		_w15189_,
		_w15439_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		_w15190_,
		_w15191_,
		_w15440_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w15192_,
		_w15193_,
		_w15441_
	);
	LUT2 #(
		.INIT('h1)
	) name4930 (
		_w15194_,
		_w15195_,
		_w15442_
	);
	LUT2 #(
		.INIT('h1)
	) name4931 (
		_w15196_,
		_w15197_,
		_w15443_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w15198_,
		_w15199_,
		_w15444_
	);
	LUT2 #(
		.INIT('h1)
	) name4933 (
		_w15200_,
		_w15201_,
		_w15445_
	);
	LUT2 #(
		.INIT('h1)
	) name4934 (
		_w15202_,
		_w15203_,
		_w15446_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w15204_,
		_w15205_,
		_w15447_
	);
	LUT2 #(
		.INIT('h1)
	) name4936 (
		_w15206_,
		_w15207_,
		_w15448_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w15208_,
		_w15209_,
		_w15449_
	);
	LUT2 #(
		.INIT('h1)
	) name4938 (
		_w15210_,
		_w15211_,
		_w15450_
	);
	LUT2 #(
		.INIT('h1)
	) name4939 (
		_w15212_,
		_w15213_,
		_w15451_
	);
	LUT2 #(
		.INIT('h1)
	) name4940 (
		_w15214_,
		_w15215_,
		_w15452_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w15216_,
		_w15217_,
		_w15453_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w15218_,
		_w15219_,
		_w15454_
	);
	LUT2 #(
		.INIT('h1)
	) name4943 (
		_w15220_,
		_w15221_,
		_w15455_
	);
	LUT2 #(
		.INIT('h1)
	) name4944 (
		_w15222_,
		_w15223_,
		_w15456_
	);
	LUT2 #(
		.INIT('h1)
	) name4945 (
		_w15224_,
		_w15225_,
		_w15457_
	);
	LUT2 #(
		.INIT('h1)
	) name4946 (
		_w15226_,
		_w15227_,
		_w15458_
	);
	LUT2 #(
		.INIT('h1)
	) name4947 (
		_w15228_,
		_w15229_,
		_w15459_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		_w15230_,
		_w15231_,
		_w15460_
	);
	LUT2 #(
		.INIT('h1)
	) name4949 (
		_w15232_,
		_w15233_,
		_w15461_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		_w15234_,
		_w15235_,
		_w15462_
	);
	LUT2 #(
		.INIT('h1)
	) name4951 (
		_w15236_,
		_w15237_,
		_w15463_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w15238_,
		_w15239_,
		_w15464_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		_w15240_,
		_w15241_,
		_w15465_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		_w15242_,
		_w15243_,
		_w15466_
	);
	LUT2 #(
		.INIT('h1)
	) name4955 (
		_w15244_,
		_w15245_,
		_w15467_
	);
	LUT2 #(
		.INIT('h1)
	) name4956 (
		_w15246_,
		_w15247_,
		_w15468_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		_w15248_,
		_w15249_,
		_w15469_
	);
	LUT2 #(
		.INIT('h1)
	) name4958 (
		_w15250_,
		_w15251_,
		_w15470_
	);
	LUT2 #(
		.INIT('h1)
	) name4959 (
		_w15252_,
		_w15253_,
		_w15471_
	);
	LUT2 #(
		.INIT('h1)
	) name4960 (
		_w15254_,
		_w15255_,
		_w15472_
	);
	LUT2 #(
		.INIT('h1)
	) name4961 (
		_w15256_,
		_w15257_,
		_w15473_
	);
	LUT2 #(
		.INIT('h1)
	) name4962 (
		_w15258_,
		_w15259_,
		_w15474_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		_w15260_,
		_w15261_,
		_w15475_
	);
	LUT2 #(
		.INIT('h1)
	) name4964 (
		_w15262_,
		_w15263_,
		_w15476_
	);
	LUT2 #(
		.INIT('h1)
	) name4965 (
		_w15264_,
		_w15265_,
		_w15477_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w15266_,
		_w15267_,
		_w15478_
	);
	LUT2 #(
		.INIT('h1)
	) name4967 (
		_w15268_,
		_w15269_,
		_w15479_
	);
	LUT2 #(
		.INIT('h1)
	) name4968 (
		_w15270_,
		_w15271_,
		_w15480_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		_w15272_,
		_w15273_,
		_w15481_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		_w15274_,
		_w15275_,
		_w15482_
	);
	LUT2 #(
		.INIT('h1)
	) name4971 (
		_w15276_,
		_w15277_,
		_w15483_
	);
	LUT2 #(
		.INIT('h1)
	) name4972 (
		_w15278_,
		_w15279_,
		_w15484_
	);
	LUT2 #(
		.INIT('h1)
	) name4973 (
		_w15280_,
		_w15281_,
		_w15485_
	);
	LUT2 #(
		.INIT('h1)
	) name4974 (
		_w15282_,
		_w15283_,
		_w15486_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w15284_,
		_w15285_,
		_w15487_
	);
	LUT2 #(
		.INIT('h1)
	) name4976 (
		_w15286_,
		_w15287_,
		_w15488_
	);
	LUT2 #(
		.INIT('h1)
	) name4977 (
		_w15288_,
		_w15289_,
		_w15489_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w15290_,
		_w15291_,
		_w15490_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		_w15292_,
		_w15293_,
		_w15491_
	);
	LUT2 #(
		.INIT('h1)
	) name4980 (
		_w15294_,
		_w15295_,
		_w15492_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		_w15296_,
		_w15297_,
		_w15493_
	);
	LUT2 #(
		.INIT('h1)
	) name4982 (
		_w15298_,
		_w15299_,
		_w15494_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w15300_,
		_w15301_,
		_w15495_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w15302_,
		_w15303_,
		_w15496_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w15304_,
		_w15305_,
		_w15497_
	);
	LUT2 #(
		.INIT('h1)
	) name4986 (
		_w15306_,
		_w15307_,
		_w15498_
	);
	LUT2 #(
		.INIT('h1)
	) name4987 (
		_w15308_,
		_w15309_,
		_w15499_
	);
	LUT2 #(
		.INIT('h1)
	) name4988 (
		_w15310_,
		_w15311_,
		_w15500_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		_w15312_,
		_w15313_,
		_w15501_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w15314_,
		_w15315_,
		_w15502_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		_w15316_,
		_w15317_,
		_w15503_
	);
	LUT2 #(
		.INIT('h1)
	) name4992 (
		_w15318_,
		_w15319_,
		_w15504_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w15320_,
		_w15321_,
		_w15505_
	);
	LUT2 #(
		.INIT('h1)
	) name4994 (
		_w15322_,
		_w15323_,
		_w15506_
	);
	LUT2 #(
		.INIT('h1)
	) name4995 (
		_w15324_,
		_w15325_,
		_w15507_
	);
	LUT2 #(
		.INIT('h1)
	) name4996 (
		_w15326_,
		_w15327_,
		_w15508_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w15328_,
		_w15329_,
		_w15509_
	);
	LUT2 #(
		.INIT('h1)
	) name4998 (
		_w15330_,
		_w15331_,
		_w15510_
	);
	LUT2 #(
		.INIT('h1)
	) name4999 (
		_w15332_,
		_w15333_,
		_w15511_
	);
	LUT2 #(
		.INIT('h1)
	) name5000 (
		_w15334_,
		_w15335_,
		_w15512_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		_w15336_,
		_w15337_,
		_w15513_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w15338_,
		_w15339_,
		_w15514_
	);
	LUT2 #(
		.INIT('h1)
	) name5003 (
		_w15340_,
		_w15341_,
		_w15515_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w15342_,
		_w15343_,
		_w15516_
	);
	LUT2 #(
		.INIT('h1)
	) name5005 (
		_w15344_,
		_w15345_,
		_w15517_
	);
	LUT2 #(
		.INIT('h1)
	) name5006 (
		_w15346_,
		_w15347_,
		_w15518_
	);
	LUT2 #(
		.INIT('h1)
	) name5007 (
		_w15348_,
		_w15349_,
		_w15519_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		_w15350_,
		_w15351_,
		_w15520_
	);
	LUT2 #(
		.INIT('h1)
	) name5009 (
		_w15352_,
		_w15353_,
		_w15521_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w15354_,
		_w15355_,
		_w15522_
	);
	LUT2 #(
		.INIT('h1)
	) name5011 (
		_w15356_,
		_w15357_,
		_w15523_
	);
	LUT2 #(
		.INIT('h1)
	) name5012 (
		_w15358_,
		_w15359_,
		_w15524_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		_w15360_,
		_w15361_,
		_w15525_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w15362_,
		_w15363_,
		_w15526_
	);
	LUT2 #(
		.INIT('h1)
	) name5015 (
		_w15364_,
		_w15365_,
		_w15527_
	);
	LUT2 #(
		.INIT('h1)
	) name5016 (
		_w15366_,
		_w15367_,
		_w15528_
	);
	LUT2 #(
		.INIT('h1)
	) name5017 (
		_w15368_,
		_w15369_,
		_w15529_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		_w15370_,
		_w15371_,
		_w15530_
	);
	LUT2 #(
		.INIT('h1)
	) name5019 (
		_w15372_,
		_w15373_,
		_w15531_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w15374_,
		_w15375_,
		_w15532_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		_w15376_,
		_w15377_,
		_w15533_
	);
	LUT2 #(
		.INIT('h1)
	) name5022 (
		_w15378_,
		_w15379_,
		_w15534_
	);
	LUT2 #(
		.INIT('h1)
	) name5023 (
		_w15380_,
		_w15381_,
		_w15535_
	);
	LUT2 #(
		.INIT('h1)
	) name5024 (
		_w15382_,
		_w15383_,
		_w15536_
	);
	LUT2 #(
		.INIT('h1)
	) name5025 (
		_w15384_,
		_w15385_,
		_w15537_
	);
	LUT2 #(
		.INIT('h1)
	) name5026 (
		_w15386_,
		_w15387_,
		_w15538_
	);
	LUT2 #(
		.INIT('h1)
	) name5027 (
		_w15388_,
		_w15389_,
		_w15539_
	);
	LUT2 #(
		.INIT('h1)
	) name5028 (
		_w15390_,
		_w15391_,
		_w15540_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		_w15392_,
		_w15393_,
		_w15541_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w15394_,
		_w15395_,
		_w15542_
	);
	LUT2 #(
		.INIT('h1)
	) name5031 (
		_w15396_,
		_w15397_,
		_w15543_
	);
	LUT2 #(
		.INIT('h1)
	) name5032 (
		_w15398_,
		_w15399_,
		_w15544_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		_w15400_,
		_w15401_,
		_w15545_
	);
	LUT2 #(
		.INIT('h1)
	) name5034 (
		_w15402_,
		_w15403_,
		_w15546_
	);
	LUT2 #(
		.INIT('h1)
	) name5035 (
		_w15404_,
		_w15405_,
		_w15547_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w15406_,
		_w15407_,
		_w15548_
	);
	LUT2 #(
		.INIT('h1)
	) name5037 (
		_w15408_,
		_w15409_,
		_w15549_
	);
	LUT2 #(
		.INIT('h1)
	) name5038 (
		_w15410_,
		_w15411_,
		_w15550_
	);
	LUT2 #(
		.INIT('h1)
	) name5039 (
		_w15412_,
		_w15413_,
		_w15551_
	);
	LUT2 #(
		.INIT('h1)
	) name5040 (
		_w15414_,
		_w15415_,
		_w15552_
	);
	LUT2 #(
		.INIT('h1)
	) name5041 (
		_w15416_,
		_w15417_,
		_w15553_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w15418_,
		_w15419_,
		_w15554_
	);
	LUT2 #(
		.INIT('h1)
	) name5043 (
		_w15420_,
		_w15421_,
		_w15555_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w15422_,
		_w15423_,
		_w15556_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w15424_,
		_w15425_,
		_w15557_
	);
	LUT2 #(
		.INIT('h1)
	) name5046 (
		_w15426_,
		_w15427_,
		_w15558_
	);
	LUT2 #(
		.INIT('h1)
	) name5047 (
		_w15428_,
		_w15429_,
		_w15559_
	);
	LUT2 #(
		.INIT('h1)
	) name5048 (
		_w15430_,
		_w15431_,
		_w15560_
	);
	LUT2 #(
		.INIT('h1)
	) name5049 (
		_w15432_,
		_w15433_,
		_w15561_
	);
	LUT2 #(
		.INIT('h8)
	) name5050 (
		_w15560_,
		_w15561_,
		_w15562_
	);
	LUT2 #(
		.INIT('h8)
	) name5051 (
		_w15558_,
		_w15559_,
		_w15563_
	);
	LUT2 #(
		.INIT('h8)
	) name5052 (
		_w15556_,
		_w15557_,
		_w15564_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		_w15554_,
		_w15555_,
		_w15565_
	);
	LUT2 #(
		.INIT('h8)
	) name5054 (
		_w15552_,
		_w15553_,
		_w15566_
	);
	LUT2 #(
		.INIT('h8)
	) name5055 (
		_w15550_,
		_w15551_,
		_w15567_
	);
	LUT2 #(
		.INIT('h8)
	) name5056 (
		_w15548_,
		_w15549_,
		_w15568_
	);
	LUT2 #(
		.INIT('h8)
	) name5057 (
		_w15546_,
		_w15547_,
		_w15569_
	);
	LUT2 #(
		.INIT('h8)
	) name5058 (
		_w15544_,
		_w15545_,
		_w15570_
	);
	LUT2 #(
		.INIT('h8)
	) name5059 (
		_w15542_,
		_w15543_,
		_w15571_
	);
	LUT2 #(
		.INIT('h8)
	) name5060 (
		_w15540_,
		_w15541_,
		_w15572_
	);
	LUT2 #(
		.INIT('h8)
	) name5061 (
		_w15538_,
		_w15539_,
		_w15573_
	);
	LUT2 #(
		.INIT('h8)
	) name5062 (
		_w15536_,
		_w15537_,
		_w15574_
	);
	LUT2 #(
		.INIT('h8)
	) name5063 (
		_w15534_,
		_w15535_,
		_w15575_
	);
	LUT2 #(
		.INIT('h8)
	) name5064 (
		_w15532_,
		_w15533_,
		_w15576_
	);
	LUT2 #(
		.INIT('h8)
	) name5065 (
		_w15530_,
		_w15531_,
		_w15577_
	);
	LUT2 #(
		.INIT('h8)
	) name5066 (
		_w15528_,
		_w15529_,
		_w15578_
	);
	LUT2 #(
		.INIT('h8)
	) name5067 (
		_w15526_,
		_w15527_,
		_w15579_
	);
	LUT2 #(
		.INIT('h8)
	) name5068 (
		_w15524_,
		_w15525_,
		_w15580_
	);
	LUT2 #(
		.INIT('h8)
	) name5069 (
		_w15522_,
		_w15523_,
		_w15581_
	);
	LUT2 #(
		.INIT('h8)
	) name5070 (
		_w15520_,
		_w15521_,
		_w15582_
	);
	LUT2 #(
		.INIT('h8)
	) name5071 (
		_w15518_,
		_w15519_,
		_w15583_
	);
	LUT2 #(
		.INIT('h8)
	) name5072 (
		_w15516_,
		_w15517_,
		_w15584_
	);
	LUT2 #(
		.INIT('h8)
	) name5073 (
		_w15514_,
		_w15515_,
		_w15585_
	);
	LUT2 #(
		.INIT('h8)
	) name5074 (
		_w15512_,
		_w15513_,
		_w15586_
	);
	LUT2 #(
		.INIT('h8)
	) name5075 (
		_w15510_,
		_w15511_,
		_w15587_
	);
	LUT2 #(
		.INIT('h8)
	) name5076 (
		_w15508_,
		_w15509_,
		_w15588_
	);
	LUT2 #(
		.INIT('h8)
	) name5077 (
		_w15506_,
		_w15507_,
		_w15589_
	);
	LUT2 #(
		.INIT('h8)
	) name5078 (
		_w15504_,
		_w15505_,
		_w15590_
	);
	LUT2 #(
		.INIT('h8)
	) name5079 (
		_w15502_,
		_w15503_,
		_w15591_
	);
	LUT2 #(
		.INIT('h8)
	) name5080 (
		_w15500_,
		_w15501_,
		_w15592_
	);
	LUT2 #(
		.INIT('h8)
	) name5081 (
		_w15498_,
		_w15499_,
		_w15593_
	);
	LUT2 #(
		.INIT('h8)
	) name5082 (
		_w15496_,
		_w15497_,
		_w15594_
	);
	LUT2 #(
		.INIT('h8)
	) name5083 (
		_w15494_,
		_w15495_,
		_w15595_
	);
	LUT2 #(
		.INIT('h8)
	) name5084 (
		_w15492_,
		_w15493_,
		_w15596_
	);
	LUT2 #(
		.INIT('h8)
	) name5085 (
		_w15490_,
		_w15491_,
		_w15597_
	);
	LUT2 #(
		.INIT('h8)
	) name5086 (
		_w15488_,
		_w15489_,
		_w15598_
	);
	LUT2 #(
		.INIT('h8)
	) name5087 (
		_w15486_,
		_w15487_,
		_w15599_
	);
	LUT2 #(
		.INIT('h8)
	) name5088 (
		_w15484_,
		_w15485_,
		_w15600_
	);
	LUT2 #(
		.INIT('h8)
	) name5089 (
		_w15482_,
		_w15483_,
		_w15601_
	);
	LUT2 #(
		.INIT('h8)
	) name5090 (
		_w15480_,
		_w15481_,
		_w15602_
	);
	LUT2 #(
		.INIT('h8)
	) name5091 (
		_w15478_,
		_w15479_,
		_w15603_
	);
	LUT2 #(
		.INIT('h8)
	) name5092 (
		_w15476_,
		_w15477_,
		_w15604_
	);
	LUT2 #(
		.INIT('h8)
	) name5093 (
		_w15474_,
		_w15475_,
		_w15605_
	);
	LUT2 #(
		.INIT('h8)
	) name5094 (
		_w15472_,
		_w15473_,
		_w15606_
	);
	LUT2 #(
		.INIT('h8)
	) name5095 (
		_w15470_,
		_w15471_,
		_w15607_
	);
	LUT2 #(
		.INIT('h8)
	) name5096 (
		_w15468_,
		_w15469_,
		_w15608_
	);
	LUT2 #(
		.INIT('h8)
	) name5097 (
		_w15466_,
		_w15467_,
		_w15609_
	);
	LUT2 #(
		.INIT('h8)
	) name5098 (
		_w15464_,
		_w15465_,
		_w15610_
	);
	LUT2 #(
		.INIT('h8)
	) name5099 (
		_w15462_,
		_w15463_,
		_w15611_
	);
	LUT2 #(
		.INIT('h8)
	) name5100 (
		_w15460_,
		_w15461_,
		_w15612_
	);
	LUT2 #(
		.INIT('h8)
	) name5101 (
		_w15458_,
		_w15459_,
		_w15613_
	);
	LUT2 #(
		.INIT('h8)
	) name5102 (
		_w15456_,
		_w15457_,
		_w15614_
	);
	LUT2 #(
		.INIT('h8)
	) name5103 (
		_w15454_,
		_w15455_,
		_w15615_
	);
	LUT2 #(
		.INIT('h8)
	) name5104 (
		_w15452_,
		_w15453_,
		_w15616_
	);
	LUT2 #(
		.INIT('h8)
	) name5105 (
		_w15450_,
		_w15451_,
		_w15617_
	);
	LUT2 #(
		.INIT('h8)
	) name5106 (
		_w15448_,
		_w15449_,
		_w15618_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		_w15446_,
		_w15447_,
		_w15619_
	);
	LUT2 #(
		.INIT('h8)
	) name5108 (
		_w15444_,
		_w15445_,
		_w15620_
	);
	LUT2 #(
		.INIT('h8)
	) name5109 (
		_w15442_,
		_w15443_,
		_w15621_
	);
	LUT2 #(
		.INIT('h8)
	) name5110 (
		_w15440_,
		_w15441_,
		_w15622_
	);
	LUT2 #(
		.INIT('h8)
	) name5111 (
		_w15438_,
		_w15439_,
		_w15623_
	);
	LUT2 #(
		.INIT('h8)
	) name5112 (
		_w15436_,
		_w15437_,
		_w15624_
	);
	LUT2 #(
		.INIT('h8)
	) name5113 (
		_w15434_,
		_w15435_,
		_w15625_
	);
	LUT2 #(
		.INIT('h8)
	) name5114 (
		_w15624_,
		_w15625_,
		_w15626_
	);
	LUT2 #(
		.INIT('h8)
	) name5115 (
		_w15622_,
		_w15623_,
		_w15627_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		_w15620_,
		_w15621_,
		_w15628_
	);
	LUT2 #(
		.INIT('h8)
	) name5117 (
		_w15618_,
		_w15619_,
		_w15629_
	);
	LUT2 #(
		.INIT('h8)
	) name5118 (
		_w15616_,
		_w15617_,
		_w15630_
	);
	LUT2 #(
		.INIT('h8)
	) name5119 (
		_w15614_,
		_w15615_,
		_w15631_
	);
	LUT2 #(
		.INIT('h8)
	) name5120 (
		_w15612_,
		_w15613_,
		_w15632_
	);
	LUT2 #(
		.INIT('h8)
	) name5121 (
		_w15610_,
		_w15611_,
		_w15633_
	);
	LUT2 #(
		.INIT('h8)
	) name5122 (
		_w15608_,
		_w15609_,
		_w15634_
	);
	LUT2 #(
		.INIT('h8)
	) name5123 (
		_w15606_,
		_w15607_,
		_w15635_
	);
	LUT2 #(
		.INIT('h8)
	) name5124 (
		_w15604_,
		_w15605_,
		_w15636_
	);
	LUT2 #(
		.INIT('h8)
	) name5125 (
		_w15602_,
		_w15603_,
		_w15637_
	);
	LUT2 #(
		.INIT('h8)
	) name5126 (
		_w15600_,
		_w15601_,
		_w15638_
	);
	LUT2 #(
		.INIT('h8)
	) name5127 (
		_w15598_,
		_w15599_,
		_w15639_
	);
	LUT2 #(
		.INIT('h8)
	) name5128 (
		_w15596_,
		_w15597_,
		_w15640_
	);
	LUT2 #(
		.INIT('h8)
	) name5129 (
		_w15594_,
		_w15595_,
		_w15641_
	);
	LUT2 #(
		.INIT('h8)
	) name5130 (
		_w15592_,
		_w15593_,
		_w15642_
	);
	LUT2 #(
		.INIT('h8)
	) name5131 (
		_w15590_,
		_w15591_,
		_w15643_
	);
	LUT2 #(
		.INIT('h8)
	) name5132 (
		_w15588_,
		_w15589_,
		_w15644_
	);
	LUT2 #(
		.INIT('h8)
	) name5133 (
		_w15586_,
		_w15587_,
		_w15645_
	);
	LUT2 #(
		.INIT('h8)
	) name5134 (
		_w15584_,
		_w15585_,
		_w15646_
	);
	LUT2 #(
		.INIT('h8)
	) name5135 (
		_w15582_,
		_w15583_,
		_w15647_
	);
	LUT2 #(
		.INIT('h8)
	) name5136 (
		_w15580_,
		_w15581_,
		_w15648_
	);
	LUT2 #(
		.INIT('h8)
	) name5137 (
		_w15578_,
		_w15579_,
		_w15649_
	);
	LUT2 #(
		.INIT('h8)
	) name5138 (
		_w15576_,
		_w15577_,
		_w15650_
	);
	LUT2 #(
		.INIT('h8)
	) name5139 (
		_w15574_,
		_w15575_,
		_w15651_
	);
	LUT2 #(
		.INIT('h8)
	) name5140 (
		_w15572_,
		_w15573_,
		_w15652_
	);
	LUT2 #(
		.INIT('h8)
	) name5141 (
		_w15570_,
		_w15571_,
		_w15653_
	);
	LUT2 #(
		.INIT('h8)
	) name5142 (
		_w15568_,
		_w15569_,
		_w15654_
	);
	LUT2 #(
		.INIT('h8)
	) name5143 (
		_w15566_,
		_w15567_,
		_w15655_
	);
	LUT2 #(
		.INIT('h8)
	) name5144 (
		_w15564_,
		_w15565_,
		_w15656_
	);
	LUT2 #(
		.INIT('h8)
	) name5145 (
		_w15562_,
		_w15563_,
		_w15657_
	);
	LUT2 #(
		.INIT('h8)
	) name5146 (
		_w15656_,
		_w15657_,
		_w15658_
	);
	LUT2 #(
		.INIT('h8)
	) name5147 (
		_w15654_,
		_w15655_,
		_w15659_
	);
	LUT2 #(
		.INIT('h8)
	) name5148 (
		_w15652_,
		_w15653_,
		_w15660_
	);
	LUT2 #(
		.INIT('h8)
	) name5149 (
		_w15650_,
		_w15651_,
		_w15661_
	);
	LUT2 #(
		.INIT('h8)
	) name5150 (
		_w15648_,
		_w15649_,
		_w15662_
	);
	LUT2 #(
		.INIT('h8)
	) name5151 (
		_w15646_,
		_w15647_,
		_w15663_
	);
	LUT2 #(
		.INIT('h8)
	) name5152 (
		_w15644_,
		_w15645_,
		_w15664_
	);
	LUT2 #(
		.INIT('h8)
	) name5153 (
		_w15642_,
		_w15643_,
		_w15665_
	);
	LUT2 #(
		.INIT('h8)
	) name5154 (
		_w15640_,
		_w15641_,
		_w15666_
	);
	LUT2 #(
		.INIT('h8)
	) name5155 (
		_w15638_,
		_w15639_,
		_w15667_
	);
	LUT2 #(
		.INIT('h8)
	) name5156 (
		_w15636_,
		_w15637_,
		_w15668_
	);
	LUT2 #(
		.INIT('h8)
	) name5157 (
		_w15634_,
		_w15635_,
		_w15669_
	);
	LUT2 #(
		.INIT('h8)
	) name5158 (
		_w15632_,
		_w15633_,
		_w15670_
	);
	LUT2 #(
		.INIT('h8)
	) name5159 (
		_w15630_,
		_w15631_,
		_w15671_
	);
	LUT2 #(
		.INIT('h8)
	) name5160 (
		_w15628_,
		_w15629_,
		_w15672_
	);
	LUT2 #(
		.INIT('h8)
	) name5161 (
		_w15626_,
		_w15627_,
		_w15673_
	);
	LUT2 #(
		.INIT('h8)
	) name5162 (
		_w15672_,
		_w15673_,
		_w15674_
	);
	LUT2 #(
		.INIT('h8)
	) name5163 (
		_w15670_,
		_w15671_,
		_w15675_
	);
	LUT2 #(
		.INIT('h8)
	) name5164 (
		_w15668_,
		_w15669_,
		_w15676_
	);
	LUT2 #(
		.INIT('h8)
	) name5165 (
		_w15666_,
		_w15667_,
		_w15677_
	);
	LUT2 #(
		.INIT('h8)
	) name5166 (
		_w15664_,
		_w15665_,
		_w15678_
	);
	LUT2 #(
		.INIT('h8)
	) name5167 (
		_w15662_,
		_w15663_,
		_w15679_
	);
	LUT2 #(
		.INIT('h8)
	) name5168 (
		_w15660_,
		_w15661_,
		_w15680_
	);
	LUT2 #(
		.INIT('h8)
	) name5169 (
		_w15658_,
		_w15659_,
		_w15681_
	);
	LUT2 #(
		.INIT('h8)
	) name5170 (
		_w15680_,
		_w15681_,
		_w15682_
	);
	LUT2 #(
		.INIT('h8)
	) name5171 (
		_w15678_,
		_w15679_,
		_w15683_
	);
	LUT2 #(
		.INIT('h8)
	) name5172 (
		_w15676_,
		_w15677_,
		_w15684_
	);
	LUT2 #(
		.INIT('h8)
	) name5173 (
		_w15674_,
		_w15675_,
		_w15685_
	);
	LUT2 #(
		.INIT('h8)
	) name5174 (
		_w15684_,
		_w15685_,
		_w15686_
	);
	LUT2 #(
		.INIT('h8)
	) name5175 (
		_w15682_,
		_w15683_,
		_w15687_
	);
	LUT2 #(
		.INIT('h8)
	) name5176 (
		_w15686_,
		_w15687_,
		_w15688_
	);
	LUT2 #(
		.INIT('h1)
	) name5177 (
		wb_rst_i_pad,
		_w15688_,
		_w15689_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		_w15176_,
		_w15689_,
		_w15690_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w15177_,
		_w15691_
	);
	LUT2 #(
		.INIT('h4)
	) name5180 (
		_w15690_,
		_w15691_,
		_w15692_
	);
	LUT2 #(
		.INIT('h8)
	) name5181 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w15147_,
		_w15693_
	);
	LUT2 #(
		.INIT('h8)
	) name5182 (
		\wishbone_RxDataLatched1_reg[9]/NET0131 ,
		_w15154_,
		_w15694_
	);
	LUT2 #(
		.INIT('h1)
	) name5183 (
		_w15693_,
		_w15694_,
		_w15695_
	);
	LUT2 #(
		.INIT('h8)
	) name5184 (
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w15175_,
		_w15696_
	);
	LUT2 #(
		.INIT('h1)
	) name5185 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w15696_,
		_w15697_
	);
	LUT2 #(
		.INIT('h8)
	) name5186 (
		m_wb_ack_i_pad,
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w15698_
	);
	LUT2 #(
		.INIT('h8)
	) name5187 (
		\wishbone_bd_ram_mem0_reg[108][1]/P0001 ,
		_w13156_,
		_w15699_
	);
	LUT2 #(
		.INIT('h8)
	) name5188 (
		\wishbone_bd_ram_mem0_reg[200][1]/P0001 ,
		_w12988_,
		_w15700_
	);
	LUT2 #(
		.INIT('h8)
	) name5189 (
		\wishbone_bd_ram_mem0_reg[90][1]/P0001 ,
		_w12978_,
		_w15701_
	);
	LUT2 #(
		.INIT('h8)
	) name5190 (
		\wishbone_bd_ram_mem0_reg[247][1]/P0001 ,
		_w12818_,
		_w15702_
	);
	LUT2 #(
		.INIT('h8)
	) name5191 (
		\wishbone_bd_ram_mem0_reg[197][1]/P0001 ,
		_w12834_,
		_w15703_
	);
	LUT2 #(
		.INIT('h8)
	) name5192 (
		\wishbone_bd_ram_mem0_reg[16][1]/P0001 ,
		_w13140_,
		_w15704_
	);
	LUT2 #(
		.INIT('h8)
	) name5193 (
		\wishbone_bd_ram_mem0_reg[2][1]/P0001 ,
		_w13088_,
		_w15705_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		\wishbone_bd_ram_mem0_reg[198][1]/P0001 ,
		_w12832_,
		_w15706_
	);
	LUT2 #(
		.INIT('h8)
	) name5195 (
		\wishbone_bd_ram_mem0_reg[60][1]/P0001 ,
		_w13204_,
		_w15707_
	);
	LUT2 #(
		.INIT('h8)
	) name5196 (
		\wishbone_bd_ram_mem0_reg[229][1]/P0001 ,
		_w12711_,
		_w15708_
	);
	LUT2 #(
		.INIT('h8)
	) name5197 (
		\wishbone_bd_ram_mem0_reg[104][1]/P0001 ,
		_w13148_,
		_w15709_
	);
	LUT2 #(
		.INIT('h8)
	) name5198 (
		\wishbone_bd_ram_mem0_reg[11][1]/P0001 ,
		_w13194_,
		_w15710_
	);
	LUT2 #(
		.INIT('h8)
	) name5199 (
		\wishbone_bd_ram_mem0_reg[72][1]/P0001 ,
		_w12810_,
		_w15711_
	);
	LUT2 #(
		.INIT('h8)
	) name5200 (
		\wishbone_bd_ram_mem0_reg[163][1]/P0001 ,
		_w12882_,
		_w15712_
	);
	LUT2 #(
		.INIT('h8)
	) name5201 (
		\wishbone_bd_ram_mem0_reg[161][1]/P0001 ,
		_w12754_,
		_w15713_
	);
	LUT2 #(
		.INIT('h8)
	) name5202 (
		\wishbone_bd_ram_mem0_reg[75][1]/P0001 ,
		_w12826_,
		_w15714_
	);
	LUT2 #(
		.INIT('h8)
	) name5203 (
		\wishbone_bd_ram_mem0_reg[230][1]/P0001 ,
		_w13036_,
		_w15715_
	);
	LUT2 #(
		.INIT('h8)
	) name5204 (
		\wishbone_bd_ram_mem0_reg[111][1]/P0001 ,
		_w12744_,
		_w15716_
	);
	LUT2 #(
		.INIT('h8)
	) name5205 (
		\wishbone_bd_ram_mem0_reg[199][1]/P0001 ,
		_w12768_,
		_w15717_
	);
	LUT2 #(
		.INIT('h8)
	) name5206 (
		\wishbone_bd_ram_mem0_reg[146][1]/P0001 ,
		_w13060_,
		_w15718_
	);
	LUT2 #(
		.INIT('h8)
	) name5207 (
		\wishbone_bd_ram_mem0_reg[231][1]/P0001 ,
		_w12856_,
		_w15719_
	);
	LUT2 #(
		.INIT('h8)
	) name5208 (
		\wishbone_bd_ram_mem0_reg[45][1]/P0001 ,
		_w12908_,
		_w15720_
	);
	LUT2 #(
		.INIT('h8)
	) name5209 (
		\wishbone_bd_ram_mem0_reg[220][1]/P0001 ,
		_w13066_,
		_w15721_
	);
	LUT2 #(
		.INIT('h8)
	) name5210 (
		\wishbone_bd_ram_mem0_reg[145][1]/P0001 ,
		_w13106_,
		_w15722_
	);
	LUT2 #(
		.INIT('h8)
	) name5211 (
		\wishbone_bd_ram_mem0_reg[53][1]/P0001 ,
		_w13020_,
		_w15723_
	);
	LUT2 #(
		.INIT('h8)
	) name5212 (
		\wishbone_bd_ram_mem0_reg[69][1]/P0001 ,
		_w12738_,
		_w15724_
	);
	LUT2 #(
		.INIT('h8)
	) name5213 (
		\wishbone_bd_ram_mem0_reg[42][1]/P0001 ,
		_w12842_,
		_w15725_
	);
	LUT2 #(
		.INIT('h8)
	) name5214 (
		\wishbone_bd_ram_mem0_reg[213][1]/P0001 ,
		_w13002_,
		_w15726_
	);
	LUT2 #(
		.INIT('h8)
	) name5215 (
		\wishbone_bd_ram_mem0_reg[215][1]/P0001 ,
		_w12974_,
		_w15727_
	);
	LUT2 #(
		.INIT('h8)
	) name5216 (
		\wishbone_bd_ram_mem0_reg[238][1]/P0001 ,
		_w13160_,
		_w15728_
	);
	LUT2 #(
		.INIT('h8)
	) name5217 (
		\wishbone_bd_ram_mem0_reg[252][1]/P0001 ,
		_w13080_,
		_w15729_
	);
	LUT2 #(
		.INIT('h8)
	) name5218 (
		\wishbone_bd_ram_mem0_reg[52][1]/P0001 ,
		_w13082_,
		_w15730_
	);
	LUT2 #(
		.INIT('h8)
	) name5219 (
		\wishbone_bd_ram_mem0_reg[54][1]/P0001 ,
		_w12770_,
		_w15731_
	);
	LUT2 #(
		.INIT('h8)
	) name5220 (
		\wishbone_bd_ram_mem0_reg[73][1]/P0001 ,
		_w12918_,
		_w15732_
	);
	LUT2 #(
		.INIT('h8)
	) name5221 (
		\wishbone_bd_ram_mem0_reg[129][1]/P0001 ,
		_w12776_,
		_w15733_
	);
	LUT2 #(
		.INIT('h8)
	) name5222 (
		\wishbone_bd_ram_mem0_reg[91][1]/P0001 ,
		_w13074_,
		_w15734_
	);
	LUT2 #(
		.INIT('h8)
	) name5223 (
		\wishbone_bd_ram_mem0_reg[34][1]/P0001 ,
		_w12930_,
		_w15735_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		\wishbone_bd_ram_mem0_reg[137][1]/P0001 ,
		_w13168_,
		_w15736_
	);
	LUT2 #(
		.INIT('h8)
	) name5225 (
		\wishbone_bd_ram_mem0_reg[59][1]/P0001 ,
		_w12780_,
		_w15737_
	);
	LUT2 #(
		.INIT('h8)
	) name5226 (
		\wishbone_bd_ram_mem0_reg[94][1]/P0001 ,
		_w13186_,
		_w15738_
	);
	LUT2 #(
		.INIT('h8)
	) name5227 (
		\wishbone_bd_ram_mem0_reg[5][1]/P0001 ,
		_w12878_,
		_w15739_
	);
	LUT2 #(
		.INIT('h8)
	) name5228 (
		\wishbone_bd_ram_mem0_reg[155][1]/P0001 ,
		_w13122_,
		_w15740_
	);
	LUT2 #(
		.INIT('h8)
	) name5229 (
		\wishbone_bd_ram_mem0_reg[255][1]/P0001 ,
		_w13072_,
		_w15741_
	);
	LUT2 #(
		.INIT('h8)
	) name5230 (
		\wishbone_bd_ram_mem0_reg[89][1]/P0001 ,
		_w12964_,
		_w15742_
	);
	LUT2 #(
		.INIT('h8)
	) name5231 (
		\wishbone_bd_ram_mem0_reg[141][1]/P0001 ,
		_w13004_,
		_w15743_
	);
	LUT2 #(
		.INIT('h8)
	) name5232 (
		\wishbone_bd_ram_mem0_reg[193][1]/P0001 ,
		_w13056_,
		_w15744_
	);
	LUT2 #(
		.INIT('h8)
	) name5233 (
		\wishbone_bd_ram_mem0_reg[51][1]/P0001 ,
		_w13024_,
		_w15745_
	);
	LUT2 #(
		.INIT('h8)
	) name5234 (
		\wishbone_bd_ram_mem0_reg[218][1]/P0001 ,
		_w13206_,
		_w15746_
	);
	LUT2 #(
		.INIT('h8)
	) name5235 (
		\wishbone_bd_ram_mem0_reg[174][1]/P0001 ,
		_w12972_,
		_w15747_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		\wishbone_bd_ram_mem0_reg[105][1]/P0001 ,
		_w12751_,
		_w15748_
	);
	LUT2 #(
		.INIT('h8)
	) name5237 (
		\wishbone_bd_ram_mem0_reg[127][1]/P0001 ,
		_w13164_,
		_w15749_
	);
	LUT2 #(
		.INIT('h8)
	) name5238 (
		\wishbone_bd_ram_mem0_reg[140][1]/P0001 ,
		_w12894_,
		_w15750_
	);
	LUT2 #(
		.INIT('h8)
	) name5239 (
		\wishbone_bd_ram_mem0_reg[115][1]/P0001 ,
		_w13112_,
		_w15751_
	);
	LUT2 #(
		.INIT('h8)
	) name5240 (
		\wishbone_bd_ram_mem0_reg[100][1]/P0001 ,
		_w12960_,
		_w15752_
	);
	LUT2 #(
		.INIT('h8)
	) name5241 (
		\wishbone_bd_ram_mem0_reg[38][1]/P0001 ,
		_w13182_,
		_w15753_
	);
	LUT2 #(
		.INIT('h8)
	) name5242 (
		\wishbone_bd_ram_mem0_reg[12][1]/P0001 ,
		_w13118_,
		_w15754_
	);
	LUT2 #(
		.INIT('h8)
	) name5243 (
		\wishbone_bd_ram_mem0_reg[95][1]/P0001 ,
		_w12844_,
		_w15755_
	);
	LUT2 #(
		.INIT('h8)
	) name5244 (
		\wishbone_bd_ram_mem0_reg[14][1]/P0001 ,
		_w13086_,
		_w15756_
	);
	LUT2 #(
		.INIT('h8)
	) name5245 (
		\wishbone_bd_ram_mem0_reg[248][1]/P0001 ,
		_w12789_,
		_w15757_
	);
	LUT2 #(
		.INIT('h8)
	) name5246 (
		\wishbone_bd_ram_mem0_reg[190][1]/P0001 ,
		_w12858_,
		_w15758_
	);
	LUT2 #(
		.INIT('h8)
	) name5247 (
		\wishbone_bd_ram_mem0_reg[181][1]/P0001 ,
		_w12828_,
		_w15759_
	);
	LUT2 #(
		.INIT('h8)
	) name5248 (
		\wishbone_bd_ram_mem0_reg[151][1]/P0001 ,
		_w13142_,
		_w15760_
	);
	LUT2 #(
		.INIT('h8)
	) name5249 (
		\wishbone_bd_ram_mem0_reg[167][1]/P0001 ,
		_w12986_,
		_w15761_
	);
	LUT2 #(
		.INIT('h8)
	) name5250 (
		\wishbone_bd_ram_mem0_reg[171][1]/P0001 ,
		_w12910_,
		_w15762_
	);
	LUT2 #(
		.INIT('h8)
	) name5251 (
		\wishbone_bd_ram_mem0_reg[7][1]/P0001 ,
		_w12728_,
		_w15763_
	);
	LUT2 #(
		.INIT('h8)
	) name5252 (
		\wishbone_bd_ram_mem0_reg[21][1]/P0001 ,
		_w12906_,
		_w15764_
	);
	LUT2 #(
		.INIT('h8)
	) name5253 (
		\wishbone_bd_ram_mem0_reg[217][1]/P0001 ,
		_w13188_,
		_w15765_
	);
	LUT2 #(
		.INIT('h8)
	) name5254 (
		\wishbone_bd_ram_mem0_reg[85][1]/P0001 ,
		_w13216_,
		_w15766_
	);
	LUT2 #(
		.INIT('h8)
	) name5255 (
		\wishbone_bd_ram_mem0_reg[44][1]/P0001 ,
		_w12896_,
		_w15767_
	);
	LUT2 #(
		.INIT('h8)
	) name5256 (
		\wishbone_bd_ram_mem0_reg[33][1]/P0001 ,
		_w12980_,
		_w15768_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		\wishbone_bd_ram_mem0_reg[17][1]/P0001 ,
		_w12848_,
		_w15769_
	);
	LUT2 #(
		.INIT('h8)
	) name5258 (
		\wishbone_bd_ram_mem0_reg[31][1]/P0001 ,
		_w13198_,
		_w15770_
	);
	LUT2 #(
		.INIT('h8)
	) name5259 (
		\wishbone_bd_ram_mem0_reg[3][1]/P0001 ,
		_w12866_,
		_w15771_
	);
	LUT2 #(
		.INIT('h8)
	) name5260 (
		\wishbone_bd_ram_mem0_reg[79][1]/P0001 ,
		_w13212_,
		_w15772_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		\wishbone_bd_ram_mem0_reg[149][1]/P0001 ,
		_w12741_,
		_w15773_
	);
	LUT2 #(
		.INIT('h8)
	) name5262 (
		\wishbone_bd_ram_mem0_reg[46][1]/P0001 ,
		_w12884_,
		_w15774_
	);
	LUT2 #(
		.INIT('h8)
	) name5263 (
		\wishbone_bd_ram_mem0_reg[84][1]/P0001 ,
		_w12934_,
		_w15775_
	);
	LUT2 #(
		.INIT('h8)
	) name5264 (
		\wishbone_bd_ram_mem0_reg[35][1]/P0001 ,
		_w12703_,
		_w15776_
	);
	LUT2 #(
		.INIT('h8)
	) name5265 (
		\wishbone_bd_ram_mem0_reg[187][1]/P0001 ,
		_w13196_,
		_w15777_
	);
	LUT2 #(
		.INIT('h8)
	) name5266 (
		\wishbone_bd_ram_mem0_reg[205][1]/P0001 ,
		_w13068_,
		_w15778_
	);
	LUT2 #(
		.INIT('h8)
	) name5267 (
		\wishbone_bd_ram_mem0_reg[201][1]/P0001 ,
		_w12822_,
		_w15779_
	);
	LUT2 #(
		.INIT('h8)
	) name5268 (
		\wishbone_bd_ram_mem0_reg[122][1]/P0001 ,
		_w13130_,
		_w15780_
	);
	LUT2 #(
		.INIT('h8)
	) name5269 (
		\wishbone_bd_ram_mem0_reg[130][1]/P0001 ,
		_w12914_,
		_w15781_
	);
	LUT2 #(
		.INIT('h8)
	) name5270 (
		\wishbone_bd_ram_mem0_reg[13][1]/P0001 ,
		_w13178_,
		_w15782_
	);
	LUT2 #(
		.INIT('h8)
	) name5271 (
		\wishbone_bd_ram_mem0_reg[166][1]/P0001 ,
		_w13040_,
		_w15783_
	);
	LUT2 #(
		.INIT('h8)
	) name5272 (
		\wishbone_bd_ram_mem0_reg[57][1]/P0001 ,
		_w13116_,
		_w15784_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		\wishbone_bd_ram_mem0_reg[50][1]/P0001 ,
		_w13150_,
		_w15785_
	);
	LUT2 #(
		.INIT('h8)
	) name5274 (
		\wishbone_bd_ram_mem0_reg[216][1]/P0001 ,
		_w13028_,
		_w15786_
	);
	LUT2 #(
		.INIT('h8)
	) name5275 (
		\wishbone_bd_ram_mem0_reg[249][1]/P0001 ,
		_w12900_,
		_w15787_
	);
	LUT2 #(
		.INIT('h8)
	) name5276 (
		\wishbone_bd_ram_mem0_reg[241][1]/P0001 ,
		_w13006_,
		_w15788_
	);
	LUT2 #(
		.INIT('h8)
	) name5277 (
		\wishbone_bd_ram_mem0_reg[168][1]/P0001 ,
		_w13208_,
		_w15789_
	);
	LUT2 #(
		.INIT('h8)
	) name5278 (
		\wishbone_bd_ram_mem0_reg[244][1]/P0001 ,
		_w12747_,
		_w15790_
	);
	LUT2 #(
		.INIT('h8)
	) name5279 (
		\wishbone_bd_ram_mem0_reg[19][1]/P0001 ,
		_w13012_,
		_w15791_
	);
	LUT2 #(
		.INIT('h8)
	) name5280 (
		\wishbone_bd_ram_mem0_reg[40][1]/P0001 ,
		_w13132_,
		_w15792_
	);
	LUT2 #(
		.INIT('h8)
	) name5281 (
		\wishbone_bd_ram_mem0_reg[126][1]/P0001 ,
		_w13218_,
		_w15793_
	);
	LUT2 #(
		.INIT('h8)
	) name5282 (
		\wishbone_bd_ram_mem0_reg[222][1]/P0001 ,
		_w13094_,
		_w15794_
	);
	LUT2 #(
		.INIT('h8)
	) name5283 (
		\wishbone_bd_ram_mem0_reg[55][1]/P0001 ,
		_w12785_,
		_w15795_
	);
	LUT2 #(
		.INIT('h8)
	) name5284 (
		\wishbone_bd_ram_mem0_reg[18][1]/P0001 ,
		_w12679_,
		_w15796_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		\wishbone_bd_ram_mem0_reg[47][1]/P0001 ,
		_w12904_,
		_w15797_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		\wishbone_bd_ram_mem0_reg[143][1]/P0001 ,
		_w12922_,
		_w15798_
	);
	LUT2 #(
		.INIT('h8)
	) name5287 (
		\wishbone_bd_ram_mem0_reg[63][1]/P0001 ,
		_w12850_,
		_w15799_
	);
	LUT2 #(
		.INIT('h8)
	) name5288 (
		\wishbone_bd_ram_mem0_reg[135][1]/P0001 ,
		_w13124_,
		_w15800_
	);
	LUT2 #(
		.INIT('h8)
	) name5289 (
		\wishbone_bd_ram_mem0_reg[58][1]/P0001 ,
		_w13070_,
		_w15801_
	);
	LUT2 #(
		.INIT('h8)
	) name5290 (
		\wishbone_bd_ram_mem0_reg[175][1]/P0001 ,
		_w13126_,
		_w15802_
	);
	LUT2 #(
		.INIT('h8)
	) name5291 (
		\wishbone_bd_ram_mem0_reg[214][1]/P0001 ,
		_w12984_,
		_w15803_
	);
	LUT2 #(
		.INIT('h8)
	) name5292 (
		\wishbone_bd_ram_mem0_reg[196][1]/P0001 ,
		_w13090_,
		_w15804_
	);
	LUT2 #(
		.INIT('h8)
	) name5293 (
		\wishbone_bd_ram_mem0_reg[1][1]/P0001 ,
		_w13014_,
		_w15805_
	);
	LUT2 #(
		.INIT('h8)
	) name5294 (
		\wishbone_bd_ram_mem0_reg[160][1]/P0001 ,
		_w12872_,
		_w15806_
	);
	LUT2 #(
		.INIT('h8)
	) name5295 (
		\wishbone_bd_ram_mem0_reg[225][1]/P0001 ,
		_w13092_,
		_w15807_
	);
	LUT2 #(
		.INIT('h8)
	) name5296 (
		\wishbone_bd_ram_mem0_reg[27][1]/P0001 ,
		_w12880_,
		_w15808_
	);
	LUT2 #(
		.INIT('h8)
	) name5297 (
		\wishbone_bd_ram_mem0_reg[124][1]/P0001 ,
		_w13058_,
		_w15809_
	);
	LUT2 #(
		.INIT('h8)
	) name5298 (
		\wishbone_bd_ram_mem0_reg[177][1]/P0001 ,
		_w12996_,
		_w15810_
	);
	LUT2 #(
		.INIT('h8)
	) name5299 (
		\wishbone_bd_ram_mem0_reg[125][1]/P0001 ,
		_w12956_,
		_w15811_
	);
	LUT2 #(
		.INIT('h8)
	) name5300 (
		\wishbone_bd_ram_mem0_reg[88][1]/P0001 ,
		_w12860_,
		_w15812_
	);
	LUT2 #(
		.INIT('h8)
	) name5301 (
		\wishbone_bd_ram_mem0_reg[159][1]/P0001 ,
		_w12774_,
		_w15813_
	);
	LUT2 #(
		.INIT('h8)
	) name5302 (
		\wishbone_bd_ram_mem0_reg[62][1]/P0001 ,
		_w12673_,
		_w15814_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		\wishbone_bd_ram_mem0_reg[114][1]/P0001 ,
		_w13202_,
		_w15815_
	);
	LUT2 #(
		.INIT('h8)
	) name5304 (
		\wishbone_bd_ram_mem0_reg[226][1]/P0001 ,
		_w13138_,
		_w15816_
	);
	LUT2 #(
		.INIT('h8)
	) name5305 (
		\wishbone_bd_ram_mem0_reg[87][1]/P0001 ,
		_w13154_,
		_w15817_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		\wishbone_bd_ram_mem0_reg[170][1]/P0001 ,
		_w13030_,
		_w15818_
	);
	LUT2 #(
		.INIT('h8)
	) name5307 (
		\wishbone_bd_ram_mem0_reg[109][1]/P0001 ,
		_w12888_,
		_w15819_
	);
	LUT2 #(
		.INIT('h8)
	) name5308 (
		\wishbone_bd_ram_mem0_reg[22][1]/P0001 ,
		_w13110_,
		_w15820_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		\wishbone_bd_ram_mem0_reg[107][1]/P0001 ,
		_w12749_,
		_w15821_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		\wishbone_bd_ram_mem0_reg[184][1]/P0001 ,
		_w13062_,
		_w15822_
	);
	LUT2 #(
		.INIT('h8)
	) name5311 (
		\wishbone_bd_ram_mem0_reg[242][1]/P0001 ,
		_w12932_,
		_w15823_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		\wishbone_bd_ram_mem0_reg[245][1]/P0001 ,
		_w13022_,
		_w15824_
	);
	LUT2 #(
		.INIT('h8)
	) name5313 (
		\wishbone_bd_ram_mem0_reg[123][1]/P0001 ,
		_w13114_,
		_w15825_
	);
	LUT2 #(
		.INIT('h8)
	) name5314 (
		\wishbone_bd_ram_mem0_reg[250][1]/P0001 ,
		_w13128_,
		_w15826_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\wishbone_bd_ram_mem0_reg[29][1]/P0001 ,
		_w12952_,
		_w15827_
	);
	LUT2 #(
		.INIT('h8)
	) name5316 (
		\wishbone_bd_ram_mem0_reg[152][1]/P0001 ,
		_w12966_,
		_w15828_
	);
	LUT2 #(
		.INIT('h8)
	) name5317 (
		\wishbone_bd_ram_mem0_reg[239][1]/P0001 ,
		_w12862_,
		_w15829_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		\wishbone_bd_ram_mem0_reg[219][1]/P0001 ,
		_w12806_,
		_w15830_
	);
	LUT2 #(
		.INIT('h8)
	) name5319 (
		\wishbone_bd_ram_mem0_reg[191][1]/P0001 ,
		_w13034_,
		_w15831_
	);
	LUT2 #(
		.INIT('h8)
	) name5320 (
		\wishbone_bd_ram_mem0_reg[139][1]/P0001 ,
		_w12814_,
		_w15832_
	);
	LUT2 #(
		.INIT('h8)
	) name5321 (
		\wishbone_bd_ram_mem0_reg[182][1]/P0001 ,
		_w12820_,
		_w15833_
	);
	LUT2 #(
		.INIT('h8)
	) name5322 (
		\wishbone_bd_ram_mem0_reg[119][1]/P0001 ,
		_w13048_,
		_w15834_
	);
	LUT2 #(
		.INIT('h8)
	) name5323 (
		\wishbone_bd_ram_mem0_reg[103][1]/P0001 ,
		_w12846_,
		_w15835_
	);
	LUT2 #(
		.INIT('h8)
	) name5324 (
		\wishbone_bd_ram_mem0_reg[96][1]/P0001 ,
		_w12912_,
		_w15836_
	);
	LUT2 #(
		.INIT('h8)
	) name5325 (
		\wishbone_bd_ram_mem0_reg[83][1]/P0001 ,
		_w12916_,
		_w15837_
	);
	LUT2 #(
		.INIT('h8)
	) name5326 (
		\wishbone_bd_ram_mem0_reg[133][1]/P0001 ,
		_w12761_,
		_w15838_
	);
	LUT2 #(
		.INIT('h8)
	) name5327 (
		\wishbone_bd_ram_mem0_reg[243][1]/P0001 ,
		_w12804_,
		_w15839_
	);
	LUT2 #(
		.INIT('h8)
	) name5328 (
		\wishbone_bd_ram_mem0_reg[150][1]/P0001 ,
		_w13136_,
		_w15840_
	);
	LUT2 #(
		.INIT('h8)
	) name5329 (
		\wishbone_bd_ram_mem0_reg[251][1]/P0001 ,
		_w13054_,
		_w15841_
	);
	LUT2 #(
		.INIT('h8)
	) name5330 (
		\wishbone_bd_ram_mem0_reg[43][1]/P0001 ,
		_w13200_,
		_w15842_
	);
	LUT2 #(
		.INIT('h8)
	) name5331 (
		\wishbone_bd_ram_mem0_reg[61][1]/P0001 ,
		_w12725_,
		_w15843_
	);
	LUT2 #(
		.INIT('h8)
	) name5332 (
		\wishbone_bd_ram_mem0_reg[158][1]/P0001 ,
		_w12898_,
		_w15844_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		\wishbone_bd_ram_mem0_reg[148][1]/P0001 ,
		_w13000_,
		_w15845_
	);
	LUT2 #(
		.INIT('h8)
	) name5334 (
		\wishbone_bd_ram_mem0_reg[142][1]/P0001 ,
		_w12928_,
		_w15846_
	);
	LUT2 #(
		.INIT('h8)
	) name5335 (
		\wishbone_bd_ram_mem0_reg[102][1]/P0001 ,
		_w12685_,
		_w15847_
	);
	LUT2 #(
		.INIT('h8)
	) name5336 (
		\wishbone_bd_ram_mem0_reg[134][1]/P0001 ,
		_w12763_,
		_w15848_
	);
	LUT2 #(
		.INIT('h8)
	) name5337 (
		\wishbone_bd_ram_mem0_reg[93][1]/P0001 ,
		_w13016_,
		_w15849_
	);
	LUT2 #(
		.INIT('h8)
	) name5338 (
		\wishbone_bd_ram_mem0_reg[162][1]/P0001 ,
		_w13098_,
		_w15850_
	);
	LUT2 #(
		.INIT('h8)
	) name5339 (
		\wishbone_bd_ram_mem0_reg[188][1]/P0001 ,
		_w12948_,
		_w15851_
	);
	LUT2 #(
		.INIT('h8)
	) name5340 (
		\wishbone_bd_ram_mem0_reg[223][1]/P0001 ,
		_w12838_,
		_w15852_
	);
	LUT2 #(
		.INIT('h8)
	) name5341 (
		\wishbone_bd_ram_mem0_reg[227][1]/P0001 ,
		_w12936_,
		_w15853_
	);
	LUT2 #(
		.INIT('h8)
	) name5342 (
		\wishbone_bd_ram_mem0_reg[24][1]/P0001 ,
		_w13084_,
		_w15854_
	);
	LUT2 #(
		.INIT('h8)
	) name5343 (
		\wishbone_bd_ram_mem0_reg[48][1]/P0001 ,
		_w12970_,
		_w15855_
	);
	LUT2 #(
		.INIT('h8)
	) name5344 (
		\wishbone_bd_ram_mem0_reg[232][1]/P0001 ,
		_w12758_,
		_w15856_
	);
	LUT2 #(
		.INIT('h8)
	) name5345 (
		\wishbone_bd_ram_mem0_reg[154][1]/P0001 ,
		_w12962_,
		_w15857_
	);
	LUT2 #(
		.INIT('h8)
	) name5346 (
		\wishbone_bd_ram_mem0_reg[113][1]/P0001 ,
		_w13026_,
		_w15858_
	);
	LUT2 #(
		.INIT('h8)
	) name5347 (
		\wishbone_bd_ram_mem0_reg[165][1]/P0001 ,
		_w13044_,
		_w15859_
	);
	LUT2 #(
		.INIT('h8)
	) name5348 (
		\wishbone_bd_ram_mem0_reg[164][1]/P0001 ,
		_w12876_,
		_w15860_
	);
	LUT2 #(
		.INIT('h8)
	) name5349 (
		\wishbone_bd_ram_mem0_reg[76][1]/P0001 ,
		_w13184_,
		_w15861_
	);
	LUT2 #(
		.INIT('h8)
	) name5350 (
		\wishbone_bd_ram_mem0_reg[8][1]/P0001 ,
		_w12920_,
		_w15862_
	);
	LUT2 #(
		.INIT('h8)
	) name5351 (
		\wishbone_bd_ram_mem0_reg[212][1]/P0001 ,
		_w12796_,
		_w15863_
	);
	LUT2 #(
		.INIT('h8)
	) name5352 (
		\wishbone_bd_ram_mem0_reg[208][1]/P0001 ,
		_w13032_,
		_w15864_
	);
	LUT2 #(
		.INIT('h8)
	) name5353 (
		\wishbone_bd_ram_mem0_reg[68][1]/P0001 ,
		_w12946_,
		_w15865_
	);
	LUT2 #(
		.INIT('h8)
	) name5354 (
		\wishbone_bd_ram_mem0_reg[67][1]/P0001 ,
		_w13134_,
		_w15866_
	);
	LUT2 #(
		.INIT('h8)
	) name5355 (
		\wishbone_bd_ram_mem0_reg[169][1]/P0001 ,
		_w12722_,
		_w15867_
	);
	LUT2 #(
		.INIT('h8)
	) name5356 (
		\wishbone_bd_ram_mem0_reg[41][1]/P0001 ,
		_w13052_,
		_w15868_
	);
	LUT2 #(
		.INIT('h8)
	) name5357 (
		\wishbone_bd_ram_mem0_reg[236][1]/P0001 ,
		_w12731_,
		_w15869_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		\wishbone_bd_ram_mem0_reg[65][1]/P0001 ,
		_w13176_,
		_w15870_
	);
	LUT2 #(
		.INIT('h8)
	) name5359 (
		\wishbone_bd_ram_mem0_reg[110][1]/P0001 ,
		_w13046_,
		_w15871_
	);
	LUT2 #(
		.INIT('h8)
	) name5360 (
		\wishbone_bd_ram_mem0_reg[23][1]/P0001 ,
		_w13008_,
		_w15872_
	);
	LUT2 #(
		.INIT('h8)
	) name5361 (
		\wishbone_bd_ram_mem0_reg[97][1]/P0001 ,
		_w13096_,
		_w15873_
	);
	LUT2 #(
		.INIT('h8)
	) name5362 (
		\wishbone_bd_ram_mem0_reg[254][1]/P0001 ,
		_w12892_,
		_w15874_
	);
	LUT2 #(
		.INIT('h8)
	) name5363 (
		\wishbone_bd_ram_mem0_reg[56][1]/P0001 ,
		_w12778_,
		_w15875_
	);
	LUT2 #(
		.INIT('h8)
	) name5364 (
		\wishbone_bd_ram_mem0_reg[147][1]/P0001 ,
		_w13146_,
		_w15876_
	);
	LUT2 #(
		.INIT('h8)
	) name5365 (
		\wishbone_bd_ram_mem0_reg[210][1]/P0001 ,
		_w12924_,
		_w15877_
	);
	LUT2 #(
		.INIT('h8)
	) name5366 (
		\wishbone_bd_ram_mem0_reg[157][1]/P0001 ,
		_w12926_,
		_w15878_
	);
	LUT2 #(
		.INIT('h8)
	) name5367 (
		\wishbone_bd_ram_mem0_reg[64][1]/P0001 ,
		_w12976_,
		_w15879_
	);
	LUT2 #(
		.INIT('h8)
	) name5368 (
		\wishbone_bd_ram_mem0_reg[209][1]/P0001 ,
		_w13152_,
		_w15880_
	);
	LUT2 #(
		.INIT('h8)
	) name5369 (
		\wishbone_bd_ram_mem0_reg[78][1]/P0001 ,
		_w12874_,
		_w15881_
	);
	LUT2 #(
		.INIT('h8)
	) name5370 (
		\wishbone_bd_ram_mem0_reg[116][1]/P0001 ,
		_w12998_,
		_w15882_
	);
	LUT2 #(
		.INIT('h8)
	) name5371 (
		\wishbone_bd_ram_mem0_reg[71][1]/P0001 ,
		_w12798_,
		_w15883_
	);
	LUT2 #(
		.INIT('h8)
	) name5372 (
		\wishbone_bd_ram_mem0_reg[235][1]/P0001 ,
		_w12696_,
		_w15884_
	);
	LUT2 #(
		.INIT('h8)
	) name5373 (
		\wishbone_bd_ram_mem0_reg[228][1]/P0001 ,
		_w12765_,
		_w15885_
	);
	LUT2 #(
		.INIT('h8)
	) name5374 (
		\wishbone_bd_ram_mem0_reg[128][1]/P0001 ,
		_w12793_,
		_w15886_
	);
	LUT2 #(
		.INIT('h8)
	) name5375 (
		\wishbone_bd_ram_mem0_reg[4][1]/P0001 ,
		_w12666_,
		_w15887_
	);
	LUT2 #(
		.INIT('h8)
	) name5376 (
		\wishbone_bd_ram_mem0_reg[6][1]/P0001 ,
		_w12968_,
		_w15888_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		\wishbone_bd_ram_mem0_reg[26][1]/P0001 ,
		_w12699_,
		_w15889_
	);
	LUT2 #(
		.INIT('h8)
	) name5378 (
		\wishbone_bd_ram_mem0_reg[74][1]/P0001 ,
		_w12812_,
		_w15890_
	);
	LUT2 #(
		.INIT('h8)
	) name5379 (
		\wishbone_bd_ram_mem0_reg[81][1]/P0001 ,
		_w12950_,
		_w15891_
	);
	LUT2 #(
		.INIT('h8)
	) name5380 (
		\wishbone_bd_ram_mem0_reg[132][1]/P0001 ,
		_w12992_,
		_w15892_
	);
	LUT2 #(
		.INIT('h8)
	) name5381 (
		\wishbone_bd_ram_mem0_reg[66][1]/P0001 ,
		_w12824_,
		_w15893_
	);
	LUT2 #(
		.INIT('h8)
	) name5382 (
		\wishbone_bd_ram_mem0_reg[70][1]/P0001 ,
		_w12840_,
		_w15894_
	);
	LUT2 #(
		.INIT('h8)
	) name5383 (
		\wishbone_bd_ram_mem0_reg[176][1]/P0001 ,
		_w12868_,
		_w15895_
	);
	LUT2 #(
		.INIT('h8)
	) name5384 (
		\wishbone_bd_ram_mem0_reg[204][1]/P0001 ,
		_w13162_,
		_w15896_
	);
	LUT2 #(
		.INIT('h8)
	) name5385 (
		\wishbone_bd_ram_mem0_reg[211][1]/P0001 ,
		_w13166_,
		_w15897_
	);
	LUT2 #(
		.INIT('h8)
	) name5386 (
		\wishbone_bd_ram_mem0_reg[121][1]/P0001 ,
		_w13078_,
		_w15898_
	);
	LUT2 #(
		.INIT('h8)
	) name5387 (
		\wishbone_bd_ram_mem0_reg[25][1]/P0001 ,
		_w13108_,
		_w15899_
	);
	LUT2 #(
		.INIT('h8)
	) name5388 (
		\wishbone_bd_ram_mem0_reg[207][1]/P0001 ,
		_w13180_,
		_w15900_
	);
	LUT2 #(
		.INIT('h8)
	) name5389 (
		\wishbone_bd_ram_mem0_reg[233][1]/P0001 ,
		_w12836_,
		_w15901_
	);
	LUT2 #(
		.INIT('h8)
	) name5390 (
		\wishbone_bd_ram_mem0_reg[194][1]/P0001 ,
		_w12772_,
		_w15902_
	);
	LUT2 #(
		.INIT('h8)
	) name5391 (
		\wishbone_bd_ram_mem0_reg[80][1]/P0001 ,
		_w12689_,
		_w15903_
	);
	LUT2 #(
		.INIT('h8)
	) name5392 (
		\wishbone_bd_ram_mem0_reg[144][1]/P0001 ,
		_w12756_,
		_w15904_
	);
	LUT2 #(
		.INIT('h8)
	) name5393 (
		\wishbone_bd_ram_mem0_reg[112][1]/P0001 ,
		_w12733_,
		_w15905_
	);
	LUT2 #(
		.INIT('h8)
	) name5394 (
		\wishbone_bd_ram_mem0_reg[10][1]/P0001 ,
		_w13172_,
		_w15906_
	);
	LUT2 #(
		.INIT('h8)
	) name5395 (
		\wishbone_bd_ram_mem0_reg[180][1]/P0001 ,
		_w12791_,
		_w15907_
	);
	LUT2 #(
		.INIT('h8)
	) name5396 (
		\wishbone_bd_ram_mem0_reg[120][1]/P0001 ,
		_w12707_,
		_w15908_
	);
	LUT2 #(
		.INIT('h8)
	) name5397 (
		\wishbone_bd_ram_mem0_reg[221][1]/P0001 ,
		_w12802_,
		_w15909_
	);
	LUT2 #(
		.INIT('h8)
	) name5398 (
		\wishbone_bd_ram_mem0_reg[202][1]/P0001 ,
		_w12870_,
		_w15910_
	);
	LUT2 #(
		.INIT('h8)
	) name5399 (
		\wishbone_bd_ram_mem0_reg[224][1]/P0001 ,
		_w12902_,
		_w15911_
	);
	LUT2 #(
		.INIT('h8)
	) name5400 (
		\wishbone_bd_ram_mem0_reg[30][1]/P0001 ,
		_w13104_,
		_w15912_
	);
	LUT2 #(
		.INIT('h8)
	) name5401 (
		\wishbone_bd_ram_mem0_reg[237][1]/P0001 ,
		_w12990_,
		_w15913_
	);
	LUT2 #(
		.INIT('h8)
	) name5402 (
		\wishbone_bd_ram_mem0_reg[234][1]/P0001 ,
		_w13214_,
		_w15914_
	);
	LUT2 #(
		.INIT('h8)
	) name5403 (
		\wishbone_bd_ram_mem0_reg[86][1]/P0001 ,
		_w12735_,
		_w15915_
	);
	LUT2 #(
		.INIT('h8)
	) name5404 (
		\wishbone_bd_ram_mem0_reg[118][1]/P0001 ,
		_w12830_,
		_w15916_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		\wishbone_bd_ram_mem0_reg[99][1]/P0001 ,
		_w13038_,
		_w15917_
	);
	LUT2 #(
		.INIT('h8)
	) name5406 (
		\wishbone_bd_ram_mem0_reg[206][1]/P0001 ,
		_w12954_,
		_w15918_
	);
	LUT2 #(
		.INIT('h8)
	) name5407 (
		\wishbone_bd_ram_mem0_reg[49][1]/P0001 ,
		_w12994_,
		_w15919_
	);
	LUT2 #(
		.INIT('h8)
	) name5408 (
		\wishbone_bd_ram_mem0_reg[153][1]/P0001 ,
		_w12890_,
		_w15920_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\wishbone_bd_ram_mem0_reg[77][1]/P0001 ,
		_w12982_,
		_w15921_
	);
	LUT2 #(
		.INIT('h8)
	) name5410 (
		\wishbone_bd_ram_mem0_reg[172][1]/P0001 ,
		_w12944_,
		_w15922_
	);
	LUT2 #(
		.INIT('h8)
	) name5411 (
		\wishbone_bd_ram_mem0_reg[98][1]/P0001 ,
		_w12816_,
		_w15923_
	);
	LUT2 #(
		.INIT('h8)
	) name5412 (
		\wishbone_bd_ram_mem0_reg[203][1]/P0001 ,
		_w13158_,
		_w15924_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		\wishbone_bd_ram_mem0_reg[253][1]/P0001 ,
		_w13100_,
		_w15925_
	);
	LUT2 #(
		.INIT('h8)
	) name5414 (
		\wishbone_bd_ram_mem0_reg[156][1]/P0001 ,
		_w13190_,
		_w15926_
	);
	LUT2 #(
		.INIT('h8)
	) name5415 (
		\wishbone_bd_ram_mem0_reg[192][1]/P0001 ,
		_w12938_,
		_w15927_
	);
	LUT2 #(
		.INIT('h8)
	) name5416 (
		\wishbone_bd_ram_mem0_reg[0][1]/P0001 ,
		_w12717_,
		_w15928_
	);
	LUT2 #(
		.INIT('h8)
	) name5417 (
		\wishbone_bd_ram_mem0_reg[195][1]/P0001 ,
		_w13144_,
		_w15929_
	);
	LUT2 #(
		.INIT('h8)
	) name5418 (
		\wishbone_bd_ram_mem0_reg[178][1]/P0001 ,
		_w12886_,
		_w15930_
	);
	LUT2 #(
		.INIT('h8)
	) name5419 (
		\wishbone_bd_ram_mem0_reg[246][1]/P0001 ,
		_w13076_,
		_w15931_
	);
	LUT2 #(
		.INIT('h8)
	) name5420 (
		\wishbone_bd_ram_mem0_reg[179][1]/P0001 ,
		_w13050_,
		_w15932_
	);
	LUT2 #(
		.INIT('h8)
	) name5421 (
		\wishbone_bd_ram_mem0_reg[189][1]/P0001 ,
		_w13042_,
		_w15933_
	);
	LUT2 #(
		.INIT('h8)
	) name5422 (
		\wishbone_bd_ram_mem0_reg[183][1]/P0001 ,
		_w12787_,
		_w15934_
	);
	LUT2 #(
		.INIT('h8)
	) name5423 (
		\wishbone_bd_ram_mem0_reg[15][1]/P0001 ,
		_w13210_,
		_w15935_
	);
	LUT2 #(
		.INIT('h8)
	) name5424 (
		\wishbone_bd_ram_mem0_reg[39][1]/P0001 ,
		_w13018_,
		_w15936_
	);
	LUT2 #(
		.INIT('h8)
	) name5425 (
		\wishbone_bd_ram_mem0_reg[186][1]/P0001 ,
		_w12783_,
		_w15937_
	);
	LUT2 #(
		.INIT('h8)
	) name5426 (
		\wishbone_bd_ram_mem0_reg[138][1]/P0001 ,
		_w12958_,
		_w15938_
	);
	LUT2 #(
		.INIT('h8)
	) name5427 (
		\wishbone_bd_ram_mem0_reg[92][1]/P0001 ,
		_w13010_,
		_w15939_
	);
	LUT2 #(
		.INIT('h8)
	) name5428 (
		\wishbone_bd_ram_mem0_reg[37][1]/P0001 ,
		_w13102_,
		_w15940_
	);
	LUT2 #(
		.INIT('h8)
	) name5429 (
		\wishbone_bd_ram_mem0_reg[82][1]/P0001 ,
		_w12942_,
		_w15941_
	);
	LUT2 #(
		.INIT('h8)
	) name5430 (
		\wishbone_bd_ram_mem0_reg[117][1]/P0001 ,
		_w12715_,
		_w15942_
	);
	LUT2 #(
		.INIT('h8)
	) name5431 (
		\wishbone_bd_ram_mem0_reg[240][1]/P0001 ,
		_w12864_,
		_w15943_
	);
	LUT2 #(
		.INIT('h8)
	) name5432 (
		\wishbone_bd_ram_mem0_reg[32][1]/P0001 ,
		_w13120_,
		_w15944_
	);
	LUT2 #(
		.INIT('h8)
	) name5433 (
		\wishbone_bd_ram_mem0_reg[106][1]/P0001 ,
		_w12713_,
		_w15945_
	);
	LUT2 #(
		.INIT('h8)
	) name5434 (
		\wishbone_bd_ram_mem0_reg[185][1]/P0001 ,
		_w12940_,
		_w15946_
	);
	LUT2 #(
		.INIT('h8)
	) name5435 (
		\wishbone_bd_ram_mem0_reg[20][1]/P0001 ,
		_w13174_,
		_w15947_
	);
	LUT2 #(
		.INIT('h8)
	) name5436 (
		\wishbone_bd_ram_mem0_reg[36][1]/P0001 ,
		_w12800_,
		_w15948_
	);
	LUT2 #(
		.INIT('h8)
	) name5437 (
		\wishbone_bd_ram_mem0_reg[28][1]/P0001 ,
		_w13170_,
		_w15949_
	);
	LUT2 #(
		.INIT('h8)
	) name5438 (
		\wishbone_bd_ram_mem0_reg[101][1]/P0001 ,
		_w13192_,
		_w15950_
	);
	LUT2 #(
		.INIT('h8)
	) name5439 (
		\wishbone_bd_ram_mem0_reg[173][1]/P0001 ,
		_w12854_,
		_w15951_
	);
	LUT2 #(
		.INIT('h8)
	) name5440 (
		\wishbone_bd_ram_mem0_reg[136][1]/P0001 ,
		_w13064_,
		_w15952_
	);
	LUT2 #(
		.INIT('h8)
	) name5441 (
		\wishbone_bd_ram_mem0_reg[9][1]/P0001 ,
		_w12808_,
		_w15953_
	);
	LUT2 #(
		.INIT('h8)
	) name5442 (
		\wishbone_bd_ram_mem0_reg[131][1]/P0001 ,
		_w12852_,
		_w15954_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w15699_,
		_w15700_,
		_w15955_
	);
	LUT2 #(
		.INIT('h1)
	) name5444 (
		_w15701_,
		_w15702_,
		_w15956_
	);
	LUT2 #(
		.INIT('h1)
	) name5445 (
		_w15703_,
		_w15704_,
		_w15957_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w15705_,
		_w15706_,
		_w15958_
	);
	LUT2 #(
		.INIT('h1)
	) name5447 (
		_w15707_,
		_w15708_,
		_w15959_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		_w15709_,
		_w15710_,
		_w15960_
	);
	LUT2 #(
		.INIT('h1)
	) name5449 (
		_w15711_,
		_w15712_,
		_w15961_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		_w15713_,
		_w15714_,
		_w15962_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		_w15715_,
		_w15716_,
		_w15963_
	);
	LUT2 #(
		.INIT('h1)
	) name5452 (
		_w15717_,
		_w15718_,
		_w15964_
	);
	LUT2 #(
		.INIT('h1)
	) name5453 (
		_w15719_,
		_w15720_,
		_w15965_
	);
	LUT2 #(
		.INIT('h1)
	) name5454 (
		_w15721_,
		_w15722_,
		_w15966_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w15723_,
		_w15724_,
		_w15967_
	);
	LUT2 #(
		.INIT('h1)
	) name5456 (
		_w15725_,
		_w15726_,
		_w15968_
	);
	LUT2 #(
		.INIT('h1)
	) name5457 (
		_w15727_,
		_w15728_,
		_w15969_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w15729_,
		_w15730_,
		_w15970_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		_w15731_,
		_w15732_,
		_w15971_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		_w15733_,
		_w15734_,
		_w15972_
	);
	LUT2 #(
		.INIT('h1)
	) name5461 (
		_w15735_,
		_w15736_,
		_w15973_
	);
	LUT2 #(
		.INIT('h1)
	) name5462 (
		_w15737_,
		_w15738_,
		_w15974_
	);
	LUT2 #(
		.INIT('h1)
	) name5463 (
		_w15739_,
		_w15740_,
		_w15975_
	);
	LUT2 #(
		.INIT('h1)
	) name5464 (
		_w15741_,
		_w15742_,
		_w15976_
	);
	LUT2 #(
		.INIT('h1)
	) name5465 (
		_w15743_,
		_w15744_,
		_w15977_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		_w15745_,
		_w15746_,
		_w15978_
	);
	LUT2 #(
		.INIT('h1)
	) name5467 (
		_w15747_,
		_w15748_,
		_w15979_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		_w15749_,
		_w15750_,
		_w15980_
	);
	LUT2 #(
		.INIT('h1)
	) name5469 (
		_w15751_,
		_w15752_,
		_w15981_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w15753_,
		_w15754_,
		_w15982_
	);
	LUT2 #(
		.INIT('h1)
	) name5471 (
		_w15755_,
		_w15756_,
		_w15983_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w15757_,
		_w15758_,
		_w15984_
	);
	LUT2 #(
		.INIT('h1)
	) name5473 (
		_w15759_,
		_w15760_,
		_w15985_
	);
	LUT2 #(
		.INIT('h1)
	) name5474 (
		_w15761_,
		_w15762_,
		_w15986_
	);
	LUT2 #(
		.INIT('h1)
	) name5475 (
		_w15763_,
		_w15764_,
		_w15987_
	);
	LUT2 #(
		.INIT('h1)
	) name5476 (
		_w15765_,
		_w15766_,
		_w15988_
	);
	LUT2 #(
		.INIT('h1)
	) name5477 (
		_w15767_,
		_w15768_,
		_w15989_
	);
	LUT2 #(
		.INIT('h1)
	) name5478 (
		_w15769_,
		_w15770_,
		_w15990_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		_w15771_,
		_w15772_,
		_w15991_
	);
	LUT2 #(
		.INIT('h1)
	) name5480 (
		_w15773_,
		_w15774_,
		_w15992_
	);
	LUT2 #(
		.INIT('h1)
	) name5481 (
		_w15775_,
		_w15776_,
		_w15993_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w15777_,
		_w15778_,
		_w15994_
	);
	LUT2 #(
		.INIT('h1)
	) name5483 (
		_w15779_,
		_w15780_,
		_w15995_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		_w15781_,
		_w15782_,
		_w15996_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w15783_,
		_w15784_,
		_w15997_
	);
	LUT2 #(
		.INIT('h1)
	) name5486 (
		_w15785_,
		_w15786_,
		_w15998_
	);
	LUT2 #(
		.INIT('h1)
	) name5487 (
		_w15787_,
		_w15788_,
		_w15999_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		_w15789_,
		_w15790_,
		_w16000_
	);
	LUT2 #(
		.INIT('h1)
	) name5489 (
		_w15791_,
		_w15792_,
		_w16001_
	);
	LUT2 #(
		.INIT('h1)
	) name5490 (
		_w15793_,
		_w15794_,
		_w16002_
	);
	LUT2 #(
		.INIT('h1)
	) name5491 (
		_w15795_,
		_w15796_,
		_w16003_
	);
	LUT2 #(
		.INIT('h1)
	) name5492 (
		_w15797_,
		_w15798_,
		_w16004_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w15799_,
		_w15800_,
		_w16005_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		_w15801_,
		_w15802_,
		_w16006_
	);
	LUT2 #(
		.INIT('h1)
	) name5495 (
		_w15803_,
		_w15804_,
		_w16007_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w15805_,
		_w15806_,
		_w16008_
	);
	LUT2 #(
		.INIT('h1)
	) name5497 (
		_w15807_,
		_w15808_,
		_w16009_
	);
	LUT2 #(
		.INIT('h1)
	) name5498 (
		_w15809_,
		_w15810_,
		_w16010_
	);
	LUT2 #(
		.INIT('h1)
	) name5499 (
		_w15811_,
		_w15812_,
		_w16011_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w15813_,
		_w15814_,
		_w16012_
	);
	LUT2 #(
		.INIT('h1)
	) name5501 (
		_w15815_,
		_w15816_,
		_w16013_
	);
	LUT2 #(
		.INIT('h1)
	) name5502 (
		_w15817_,
		_w15818_,
		_w16014_
	);
	LUT2 #(
		.INIT('h1)
	) name5503 (
		_w15819_,
		_w15820_,
		_w16015_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		_w15821_,
		_w15822_,
		_w16016_
	);
	LUT2 #(
		.INIT('h1)
	) name5505 (
		_w15823_,
		_w15824_,
		_w16017_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w15825_,
		_w15826_,
		_w16018_
	);
	LUT2 #(
		.INIT('h1)
	) name5507 (
		_w15827_,
		_w15828_,
		_w16019_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		_w15829_,
		_w15830_,
		_w16020_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		_w15831_,
		_w15832_,
		_w16021_
	);
	LUT2 #(
		.INIT('h1)
	) name5510 (
		_w15833_,
		_w15834_,
		_w16022_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w15835_,
		_w15836_,
		_w16023_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		_w15837_,
		_w15838_,
		_w16024_
	);
	LUT2 #(
		.INIT('h1)
	) name5513 (
		_w15839_,
		_w15840_,
		_w16025_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		_w15841_,
		_w15842_,
		_w16026_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w15843_,
		_w15844_,
		_w16027_
	);
	LUT2 #(
		.INIT('h1)
	) name5516 (
		_w15845_,
		_w15846_,
		_w16028_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w15847_,
		_w15848_,
		_w16029_
	);
	LUT2 #(
		.INIT('h1)
	) name5518 (
		_w15849_,
		_w15850_,
		_w16030_
	);
	LUT2 #(
		.INIT('h1)
	) name5519 (
		_w15851_,
		_w15852_,
		_w16031_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		_w15853_,
		_w15854_,
		_w16032_
	);
	LUT2 #(
		.INIT('h1)
	) name5521 (
		_w15855_,
		_w15856_,
		_w16033_
	);
	LUT2 #(
		.INIT('h1)
	) name5522 (
		_w15857_,
		_w15858_,
		_w16034_
	);
	LUT2 #(
		.INIT('h1)
	) name5523 (
		_w15859_,
		_w15860_,
		_w16035_
	);
	LUT2 #(
		.INIT('h1)
	) name5524 (
		_w15861_,
		_w15862_,
		_w16036_
	);
	LUT2 #(
		.INIT('h1)
	) name5525 (
		_w15863_,
		_w15864_,
		_w16037_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w15865_,
		_w15866_,
		_w16038_
	);
	LUT2 #(
		.INIT('h1)
	) name5527 (
		_w15867_,
		_w15868_,
		_w16039_
	);
	LUT2 #(
		.INIT('h1)
	) name5528 (
		_w15869_,
		_w15870_,
		_w16040_
	);
	LUT2 #(
		.INIT('h1)
	) name5529 (
		_w15871_,
		_w15872_,
		_w16041_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w15873_,
		_w15874_,
		_w16042_
	);
	LUT2 #(
		.INIT('h1)
	) name5531 (
		_w15875_,
		_w15876_,
		_w16043_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w15877_,
		_w15878_,
		_w16044_
	);
	LUT2 #(
		.INIT('h1)
	) name5533 (
		_w15879_,
		_w15880_,
		_w16045_
	);
	LUT2 #(
		.INIT('h1)
	) name5534 (
		_w15881_,
		_w15882_,
		_w16046_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w15883_,
		_w15884_,
		_w16047_
	);
	LUT2 #(
		.INIT('h1)
	) name5536 (
		_w15885_,
		_w15886_,
		_w16048_
	);
	LUT2 #(
		.INIT('h1)
	) name5537 (
		_w15887_,
		_w15888_,
		_w16049_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		_w15889_,
		_w15890_,
		_w16050_
	);
	LUT2 #(
		.INIT('h1)
	) name5539 (
		_w15891_,
		_w15892_,
		_w16051_
	);
	LUT2 #(
		.INIT('h1)
	) name5540 (
		_w15893_,
		_w15894_,
		_w16052_
	);
	LUT2 #(
		.INIT('h1)
	) name5541 (
		_w15895_,
		_w15896_,
		_w16053_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		_w15897_,
		_w15898_,
		_w16054_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		_w15899_,
		_w15900_,
		_w16055_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		_w15901_,
		_w15902_,
		_w16056_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w15903_,
		_w15904_,
		_w16057_
	);
	LUT2 #(
		.INIT('h1)
	) name5546 (
		_w15905_,
		_w15906_,
		_w16058_
	);
	LUT2 #(
		.INIT('h1)
	) name5547 (
		_w15907_,
		_w15908_,
		_w16059_
	);
	LUT2 #(
		.INIT('h1)
	) name5548 (
		_w15909_,
		_w15910_,
		_w16060_
	);
	LUT2 #(
		.INIT('h1)
	) name5549 (
		_w15911_,
		_w15912_,
		_w16061_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w15913_,
		_w15914_,
		_w16062_
	);
	LUT2 #(
		.INIT('h1)
	) name5551 (
		_w15915_,
		_w15916_,
		_w16063_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w15917_,
		_w15918_,
		_w16064_
	);
	LUT2 #(
		.INIT('h1)
	) name5553 (
		_w15919_,
		_w15920_,
		_w16065_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		_w15921_,
		_w15922_,
		_w16066_
	);
	LUT2 #(
		.INIT('h1)
	) name5555 (
		_w15923_,
		_w15924_,
		_w16067_
	);
	LUT2 #(
		.INIT('h1)
	) name5556 (
		_w15925_,
		_w15926_,
		_w16068_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		_w15927_,
		_w15928_,
		_w16069_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w15929_,
		_w15930_,
		_w16070_
	);
	LUT2 #(
		.INIT('h1)
	) name5559 (
		_w15931_,
		_w15932_,
		_w16071_
	);
	LUT2 #(
		.INIT('h1)
	) name5560 (
		_w15933_,
		_w15934_,
		_w16072_
	);
	LUT2 #(
		.INIT('h1)
	) name5561 (
		_w15935_,
		_w15936_,
		_w16073_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		_w15937_,
		_w15938_,
		_w16074_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		_w15939_,
		_w15940_,
		_w16075_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		_w15941_,
		_w15942_,
		_w16076_
	);
	LUT2 #(
		.INIT('h1)
	) name5565 (
		_w15943_,
		_w15944_,
		_w16077_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w15945_,
		_w15946_,
		_w16078_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		_w15947_,
		_w15948_,
		_w16079_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		_w15949_,
		_w15950_,
		_w16080_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w15951_,
		_w15952_,
		_w16081_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		_w15953_,
		_w15954_,
		_w16082_
	);
	LUT2 #(
		.INIT('h8)
	) name5571 (
		_w16081_,
		_w16082_,
		_w16083_
	);
	LUT2 #(
		.INIT('h8)
	) name5572 (
		_w16079_,
		_w16080_,
		_w16084_
	);
	LUT2 #(
		.INIT('h8)
	) name5573 (
		_w16077_,
		_w16078_,
		_w16085_
	);
	LUT2 #(
		.INIT('h8)
	) name5574 (
		_w16075_,
		_w16076_,
		_w16086_
	);
	LUT2 #(
		.INIT('h8)
	) name5575 (
		_w16073_,
		_w16074_,
		_w16087_
	);
	LUT2 #(
		.INIT('h8)
	) name5576 (
		_w16071_,
		_w16072_,
		_w16088_
	);
	LUT2 #(
		.INIT('h8)
	) name5577 (
		_w16069_,
		_w16070_,
		_w16089_
	);
	LUT2 #(
		.INIT('h8)
	) name5578 (
		_w16067_,
		_w16068_,
		_w16090_
	);
	LUT2 #(
		.INIT('h8)
	) name5579 (
		_w16065_,
		_w16066_,
		_w16091_
	);
	LUT2 #(
		.INIT('h8)
	) name5580 (
		_w16063_,
		_w16064_,
		_w16092_
	);
	LUT2 #(
		.INIT('h8)
	) name5581 (
		_w16061_,
		_w16062_,
		_w16093_
	);
	LUT2 #(
		.INIT('h8)
	) name5582 (
		_w16059_,
		_w16060_,
		_w16094_
	);
	LUT2 #(
		.INIT('h8)
	) name5583 (
		_w16057_,
		_w16058_,
		_w16095_
	);
	LUT2 #(
		.INIT('h8)
	) name5584 (
		_w16055_,
		_w16056_,
		_w16096_
	);
	LUT2 #(
		.INIT('h8)
	) name5585 (
		_w16053_,
		_w16054_,
		_w16097_
	);
	LUT2 #(
		.INIT('h8)
	) name5586 (
		_w16051_,
		_w16052_,
		_w16098_
	);
	LUT2 #(
		.INIT('h8)
	) name5587 (
		_w16049_,
		_w16050_,
		_w16099_
	);
	LUT2 #(
		.INIT('h8)
	) name5588 (
		_w16047_,
		_w16048_,
		_w16100_
	);
	LUT2 #(
		.INIT('h8)
	) name5589 (
		_w16045_,
		_w16046_,
		_w16101_
	);
	LUT2 #(
		.INIT('h8)
	) name5590 (
		_w16043_,
		_w16044_,
		_w16102_
	);
	LUT2 #(
		.INIT('h8)
	) name5591 (
		_w16041_,
		_w16042_,
		_w16103_
	);
	LUT2 #(
		.INIT('h8)
	) name5592 (
		_w16039_,
		_w16040_,
		_w16104_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w16037_,
		_w16038_,
		_w16105_
	);
	LUT2 #(
		.INIT('h8)
	) name5594 (
		_w16035_,
		_w16036_,
		_w16106_
	);
	LUT2 #(
		.INIT('h8)
	) name5595 (
		_w16033_,
		_w16034_,
		_w16107_
	);
	LUT2 #(
		.INIT('h8)
	) name5596 (
		_w16031_,
		_w16032_,
		_w16108_
	);
	LUT2 #(
		.INIT('h8)
	) name5597 (
		_w16029_,
		_w16030_,
		_w16109_
	);
	LUT2 #(
		.INIT('h8)
	) name5598 (
		_w16027_,
		_w16028_,
		_w16110_
	);
	LUT2 #(
		.INIT('h8)
	) name5599 (
		_w16025_,
		_w16026_,
		_w16111_
	);
	LUT2 #(
		.INIT('h8)
	) name5600 (
		_w16023_,
		_w16024_,
		_w16112_
	);
	LUT2 #(
		.INIT('h8)
	) name5601 (
		_w16021_,
		_w16022_,
		_w16113_
	);
	LUT2 #(
		.INIT('h8)
	) name5602 (
		_w16019_,
		_w16020_,
		_w16114_
	);
	LUT2 #(
		.INIT('h8)
	) name5603 (
		_w16017_,
		_w16018_,
		_w16115_
	);
	LUT2 #(
		.INIT('h8)
	) name5604 (
		_w16015_,
		_w16016_,
		_w16116_
	);
	LUT2 #(
		.INIT('h8)
	) name5605 (
		_w16013_,
		_w16014_,
		_w16117_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		_w16011_,
		_w16012_,
		_w16118_
	);
	LUT2 #(
		.INIT('h8)
	) name5607 (
		_w16009_,
		_w16010_,
		_w16119_
	);
	LUT2 #(
		.INIT('h8)
	) name5608 (
		_w16007_,
		_w16008_,
		_w16120_
	);
	LUT2 #(
		.INIT('h8)
	) name5609 (
		_w16005_,
		_w16006_,
		_w16121_
	);
	LUT2 #(
		.INIT('h8)
	) name5610 (
		_w16003_,
		_w16004_,
		_w16122_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		_w16001_,
		_w16002_,
		_w16123_
	);
	LUT2 #(
		.INIT('h8)
	) name5612 (
		_w15999_,
		_w16000_,
		_w16124_
	);
	LUT2 #(
		.INIT('h8)
	) name5613 (
		_w15997_,
		_w15998_,
		_w16125_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		_w15995_,
		_w15996_,
		_w16126_
	);
	LUT2 #(
		.INIT('h8)
	) name5615 (
		_w15993_,
		_w15994_,
		_w16127_
	);
	LUT2 #(
		.INIT('h8)
	) name5616 (
		_w15991_,
		_w15992_,
		_w16128_
	);
	LUT2 #(
		.INIT('h8)
	) name5617 (
		_w15989_,
		_w15990_,
		_w16129_
	);
	LUT2 #(
		.INIT('h8)
	) name5618 (
		_w15987_,
		_w15988_,
		_w16130_
	);
	LUT2 #(
		.INIT('h8)
	) name5619 (
		_w15985_,
		_w15986_,
		_w16131_
	);
	LUT2 #(
		.INIT('h8)
	) name5620 (
		_w15983_,
		_w15984_,
		_w16132_
	);
	LUT2 #(
		.INIT('h8)
	) name5621 (
		_w15981_,
		_w15982_,
		_w16133_
	);
	LUT2 #(
		.INIT('h8)
	) name5622 (
		_w15979_,
		_w15980_,
		_w16134_
	);
	LUT2 #(
		.INIT('h8)
	) name5623 (
		_w15977_,
		_w15978_,
		_w16135_
	);
	LUT2 #(
		.INIT('h8)
	) name5624 (
		_w15975_,
		_w15976_,
		_w16136_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		_w15973_,
		_w15974_,
		_w16137_
	);
	LUT2 #(
		.INIT('h8)
	) name5626 (
		_w15971_,
		_w15972_,
		_w16138_
	);
	LUT2 #(
		.INIT('h8)
	) name5627 (
		_w15969_,
		_w15970_,
		_w16139_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w15967_,
		_w15968_,
		_w16140_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		_w15965_,
		_w15966_,
		_w16141_
	);
	LUT2 #(
		.INIT('h8)
	) name5630 (
		_w15963_,
		_w15964_,
		_w16142_
	);
	LUT2 #(
		.INIT('h8)
	) name5631 (
		_w15961_,
		_w15962_,
		_w16143_
	);
	LUT2 #(
		.INIT('h8)
	) name5632 (
		_w15959_,
		_w15960_,
		_w16144_
	);
	LUT2 #(
		.INIT('h8)
	) name5633 (
		_w15957_,
		_w15958_,
		_w16145_
	);
	LUT2 #(
		.INIT('h8)
	) name5634 (
		_w15955_,
		_w15956_,
		_w16146_
	);
	LUT2 #(
		.INIT('h8)
	) name5635 (
		_w16145_,
		_w16146_,
		_w16147_
	);
	LUT2 #(
		.INIT('h8)
	) name5636 (
		_w16143_,
		_w16144_,
		_w16148_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		_w16141_,
		_w16142_,
		_w16149_
	);
	LUT2 #(
		.INIT('h8)
	) name5638 (
		_w16139_,
		_w16140_,
		_w16150_
	);
	LUT2 #(
		.INIT('h8)
	) name5639 (
		_w16137_,
		_w16138_,
		_w16151_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		_w16135_,
		_w16136_,
		_w16152_
	);
	LUT2 #(
		.INIT('h8)
	) name5641 (
		_w16133_,
		_w16134_,
		_w16153_
	);
	LUT2 #(
		.INIT('h8)
	) name5642 (
		_w16131_,
		_w16132_,
		_w16154_
	);
	LUT2 #(
		.INIT('h8)
	) name5643 (
		_w16129_,
		_w16130_,
		_w16155_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		_w16127_,
		_w16128_,
		_w16156_
	);
	LUT2 #(
		.INIT('h8)
	) name5645 (
		_w16125_,
		_w16126_,
		_w16157_
	);
	LUT2 #(
		.INIT('h8)
	) name5646 (
		_w16123_,
		_w16124_,
		_w16158_
	);
	LUT2 #(
		.INIT('h8)
	) name5647 (
		_w16121_,
		_w16122_,
		_w16159_
	);
	LUT2 #(
		.INIT('h8)
	) name5648 (
		_w16119_,
		_w16120_,
		_w16160_
	);
	LUT2 #(
		.INIT('h8)
	) name5649 (
		_w16117_,
		_w16118_,
		_w16161_
	);
	LUT2 #(
		.INIT('h8)
	) name5650 (
		_w16115_,
		_w16116_,
		_w16162_
	);
	LUT2 #(
		.INIT('h8)
	) name5651 (
		_w16113_,
		_w16114_,
		_w16163_
	);
	LUT2 #(
		.INIT('h8)
	) name5652 (
		_w16111_,
		_w16112_,
		_w16164_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		_w16109_,
		_w16110_,
		_w16165_
	);
	LUT2 #(
		.INIT('h8)
	) name5654 (
		_w16107_,
		_w16108_,
		_w16166_
	);
	LUT2 #(
		.INIT('h8)
	) name5655 (
		_w16105_,
		_w16106_,
		_w16167_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		_w16103_,
		_w16104_,
		_w16168_
	);
	LUT2 #(
		.INIT('h8)
	) name5657 (
		_w16101_,
		_w16102_,
		_w16169_
	);
	LUT2 #(
		.INIT('h8)
	) name5658 (
		_w16099_,
		_w16100_,
		_w16170_
	);
	LUT2 #(
		.INIT('h8)
	) name5659 (
		_w16097_,
		_w16098_,
		_w16171_
	);
	LUT2 #(
		.INIT('h8)
	) name5660 (
		_w16095_,
		_w16096_,
		_w16172_
	);
	LUT2 #(
		.INIT('h8)
	) name5661 (
		_w16093_,
		_w16094_,
		_w16173_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		_w16091_,
		_w16092_,
		_w16174_
	);
	LUT2 #(
		.INIT('h8)
	) name5663 (
		_w16089_,
		_w16090_,
		_w16175_
	);
	LUT2 #(
		.INIT('h8)
	) name5664 (
		_w16087_,
		_w16088_,
		_w16176_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		_w16085_,
		_w16086_,
		_w16177_
	);
	LUT2 #(
		.INIT('h8)
	) name5666 (
		_w16083_,
		_w16084_,
		_w16178_
	);
	LUT2 #(
		.INIT('h8)
	) name5667 (
		_w16177_,
		_w16178_,
		_w16179_
	);
	LUT2 #(
		.INIT('h8)
	) name5668 (
		_w16175_,
		_w16176_,
		_w16180_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		_w16173_,
		_w16174_,
		_w16181_
	);
	LUT2 #(
		.INIT('h8)
	) name5670 (
		_w16171_,
		_w16172_,
		_w16182_
	);
	LUT2 #(
		.INIT('h8)
	) name5671 (
		_w16169_,
		_w16170_,
		_w16183_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		_w16167_,
		_w16168_,
		_w16184_
	);
	LUT2 #(
		.INIT('h8)
	) name5673 (
		_w16165_,
		_w16166_,
		_w16185_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		_w16163_,
		_w16164_,
		_w16186_
	);
	LUT2 #(
		.INIT('h8)
	) name5675 (
		_w16161_,
		_w16162_,
		_w16187_
	);
	LUT2 #(
		.INIT('h8)
	) name5676 (
		_w16159_,
		_w16160_,
		_w16188_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		_w16157_,
		_w16158_,
		_w16189_
	);
	LUT2 #(
		.INIT('h8)
	) name5678 (
		_w16155_,
		_w16156_,
		_w16190_
	);
	LUT2 #(
		.INIT('h8)
	) name5679 (
		_w16153_,
		_w16154_,
		_w16191_
	);
	LUT2 #(
		.INIT('h8)
	) name5680 (
		_w16151_,
		_w16152_,
		_w16192_
	);
	LUT2 #(
		.INIT('h8)
	) name5681 (
		_w16149_,
		_w16150_,
		_w16193_
	);
	LUT2 #(
		.INIT('h8)
	) name5682 (
		_w16147_,
		_w16148_,
		_w16194_
	);
	LUT2 #(
		.INIT('h8)
	) name5683 (
		_w16193_,
		_w16194_,
		_w16195_
	);
	LUT2 #(
		.INIT('h8)
	) name5684 (
		_w16191_,
		_w16192_,
		_w16196_
	);
	LUT2 #(
		.INIT('h8)
	) name5685 (
		_w16189_,
		_w16190_,
		_w16197_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w16187_,
		_w16188_,
		_w16198_
	);
	LUT2 #(
		.INIT('h8)
	) name5687 (
		_w16185_,
		_w16186_,
		_w16199_
	);
	LUT2 #(
		.INIT('h8)
	) name5688 (
		_w16183_,
		_w16184_,
		_w16200_
	);
	LUT2 #(
		.INIT('h8)
	) name5689 (
		_w16181_,
		_w16182_,
		_w16201_
	);
	LUT2 #(
		.INIT('h8)
	) name5690 (
		_w16179_,
		_w16180_,
		_w16202_
	);
	LUT2 #(
		.INIT('h8)
	) name5691 (
		_w16201_,
		_w16202_,
		_w16203_
	);
	LUT2 #(
		.INIT('h8)
	) name5692 (
		_w16199_,
		_w16200_,
		_w16204_
	);
	LUT2 #(
		.INIT('h8)
	) name5693 (
		_w16197_,
		_w16198_,
		_w16205_
	);
	LUT2 #(
		.INIT('h8)
	) name5694 (
		_w16195_,
		_w16196_,
		_w16206_
	);
	LUT2 #(
		.INIT('h8)
	) name5695 (
		_w16205_,
		_w16206_,
		_w16207_
	);
	LUT2 #(
		.INIT('h8)
	) name5696 (
		_w16203_,
		_w16204_,
		_w16208_
	);
	LUT2 #(
		.INIT('h8)
	) name5697 (
		_w16207_,
		_w16208_,
		_w16209_
	);
	LUT2 #(
		.INIT('h1)
	) name5698 (
		wb_rst_i_pad,
		_w16209_,
		_w16210_
	);
	LUT2 #(
		.INIT('h2)
	) name5699 (
		_w15696_,
		_w16210_,
		_w16211_
	);
	LUT2 #(
		.INIT('h1)
	) name5700 (
		_w15697_,
		_w15698_,
		_w16212_
	);
	LUT2 #(
		.INIT('h4)
	) name5701 (
		_w16211_,
		_w16212_,
		_w16213_
	);
	LUT2 #(
		.INIT('h2)
	) name5702 (
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w11818_,
		_w16214_
	);
	LUT2 #(
		.INIT('h4)
	) name5703 (
		\rxethmac1_crcrx_Crc_reg[21]/NET0131 ,
		_w11818_,
		_w16215_
	);
	LUT2 #(
		.INIT('h2)
	) name5704 (
		_w10580_,
		_w16214_,
		_w16216_
	);
	LUT2 #(
		.INIT('h4)
	) name5705 (
		_w16215_,
		_w16216_,
		_w16217_
	);
	LUT2 #(
		.INIT('h2)
	) name5706 (
		\txethmac1_txcrc_Crc_reg[4]/NET0131 ,
		_w12472_,
		_w16218_
	);
	LUT2 #(
		.INIT('h4)
	) name5707 (
		\txethmac1_txcrc_Crc_reg[4]/NET0131 ,
		_w12472_,
		_w16219_
	);
	LUT2 #(
		.INIT('h2)
	) name5708 (
		_w11181_,
		_w16218_,
		_w16220_
	);
	LUT2 #(
		.INIT('h4)
	) name5709 (
		_w16219_,
		_w16220_,
		_w16221_
	);
	LUT2 #(
		.INIT('h8)
	) name5710 (
		\m_wb_adr_o[18]_pad ,
		_w12636_,
		_w16222_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		\m_wb_adr_o[17]_pad ,
		_w12592_,
		_w16223_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		\m_wb_adr_o[18]_pad ,
		_w16223_,
		_w16224_
	);
	LUT2 #(
		.INIT('h1)
	) name5713 (
		_w12594_,
		_w14591_,
		_w16225_
	);
	LUT2 #(
		.INIT('h4)
	) name5714 (
		_w16224_,
		_w16225_,
		_w16226_
	);
	LUT2 #(
		.INIT('h8)
	) name5715 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		_w12634_,
		_w16227_
	);
	LUT2 #(
		.INIT('h8)
	) name5716 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		_w12577_,
		_w16228_
	);
	LUT2 #(
		.INIT('h1)
	) name5717 (
		_w16222_,
		_w16227_,
		_w16229_
	);
	LUT2 #(
		.INIT('h4)
	) name5718 (
		_w16228_,
		_w16229_,
		_w16230_
	);
	LUT2 #(
		.INIT('h4)
	) name5719 (
		_w16226_,
		_w16230_,
		_w16231_
	);
	LUT2 #(
		.INIT('h8)
	) name5720 (
		\wishbone_bd_ram_mem2_reg[177][20]/P0001 ,
		_w12996_,
		_w16232_
	);
	LUT2 #(
		.INIT('h8)
	) name5721 (
		\wishbone_bd_ram_mem2_reg[166][20]/P0001 ,
		_w13040_,
		_w16233_
	);
	LUT2 #(
		.INIT('h8)
	) name5722 (
		\wishbone_bd_ram_mem2_reg[149][20]/P0001 ,
		_w12741_,
		_w16234_
	);
	LUT2 #(
		.INIT('h8)
	) name5723 (
		\wishbone_bd_ram_mem2_reg[121][20]/P0001 ,
		_w13078_,
		_w16235_
	);
	LUT2 #(
		.INIT('h8)
	) name5724 (
		\wishbone_bd_ram_mem2_reg[203][20]/P0001 ,
		_w13158_,
		_w16236_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		\wishbone_bd_ram_mem2_reg[118][20]/P0001 ,
		_w12830_,
		_w16237_
	);
	LUT2 #(
		.INIT('h8)
	) name5726 (
		\wishbone_bd_ram_mem2_reg[231][20]/P0001 ,
		_w12856_,
		_w16238_
	);
	LUT2 #(
		.INIT('h8)
	) name5727 (
		\wishbone_bd_ram_mem2_reg[15][20]/P0001 ,
		_w13210_,
		_w16239_
	);
	LUT2 #(
		.INIT('h8)
	) name5728 (
		\wishbone_bd_ram_mem2_reg[64][20]/P0001 ,
		_w12976_,
		_w16240_
	);
	LUT2 #(
		.INIT('h8)
	) name5729 (
		\wishbone_bd_ram_mem2_reg[225][20]/P0001 ,
		_w13092_,
		_w16241_
	);
	LUT2 #(
		.INIT('h8)
	) name5730 (
		\wishbone_bd_ram_mem2_reg[85][20]/P0001 ,
		_w13216_,
		_w16242_
	);
	LUT2 #(
		.INIT('h8)
	) name5731 (
		\wishbone_bd_ram_mem2_reg[237][20]/P0001 ,
		_w12990_,
		_w16243_
	);
	LUT2 #(
		.INIT('h8)
	) name5732 (
		\wishbone_bd_ram_mem2_reg[37][20]/P0001 ,
		_w13102_,
		_w16244_
	);
	LUT2 #(
		.INIT('h8)
	) name5733 (
		\wishbone_bd_ram_mem2_reg[234][20]/P0001 ,
		_w13214_,
		_w16245_
	);
	LUT2 #(
		.INIT('h8)
	) name5734 (
		\wishbone_bd_ram_mem2_reg[20][20]/P0001 ,
		_w13174_,
		_w16246_
	);
	LUT2 #(
		.INIT('h8)
	) name5735 (
		\wishbone_bd_ram_mem2_reg[147][20]/P0001 ,
		_w13146_,
		_w16247_
	);
	LUT2 #(
		.INIT('h8)
	) name5736 (
		\wishbone_bd_ram_mem2_reg[56][20]/P0001 ,
		_w12778_,
		_w16248_
	);
	LUT2 #(
		.INIT('h8)
	) name5737 (
		\wishbone_bd_ram_mem2_reg[100][20]/P0001 ,
		_w12960_,
		_w16249_
	);
	LUT2 #(
		.INIT('h8)
	) name5738 (
		\wishbone_bd_ram_mem2_reg[127][20]/P0001 ,
		_w13164_,
		_w16250_
	);
	LUT2 #(
		.INIT('h8)
	) name5739 (
		\wishbone_bd_ram_mem2_reg[144][20]/P0001 ,
		_w12756_,
		_w16251_
	);
	LUT2 #(
		.INIT('h8)
	) name5740 (
		\wishbone_bd_ram_mem2_reg[120][20]/P0001 ,
		_w12707_,
		_w16252_
	);
	LUT2 #(
		.INIT('h8)
	) name5741 (
		\wishbone_bd_ram_mem2_reg[239][20]/P0001 ,
		_w12862_,
		_w16253_
	);
	LUT2 #(
		.INIT('h8)
	) name5742 (
		\wishbone_bd_ram_mem2_reg[16][20]/P0001 ,
		_w13140_,
		_w16254_
	);
	LUT2 #(
		.INIT('h8)
	) name5743 (
		\wishbone_bd_ram_mem2_reg[79][20]/P0001 ,
		_w13212_,
		_w16255_
	);
	LUT2 #(
		.INIT('h8)
	) name5744 (
		\wishbone_bd_ram_mem2_reg[76][20]/P0001 ,
		_w13184_,
		_w16256_
	);
	LUT2 #(
		.INIT('h8)
	) name5745 (
		\wishbone_bd_ram_mem2_reg[39][20]/P0001 ,
		_w13018_,
		_w16257_
	);
	LUT2 #(
		.INIT('h8)
	) name5746 (
		\wishbone_bd_ram_mem2_reg[145][20]/P0001 ,
		_w13106_,
		_w16258_
	);
	LUT2 #(
		.INIT('h8)
	) name5747 (
		\wishbone_bd_ram_mem2_reg[111][20]/P0001 ,
		_w12744_,
		_w16259_
	);
	LUT2 #(
		.INIT('h8)
	) name5748 (
		\wishbone_bd_ram_mem2_reg[206][20]/P0001 ,
		_w12954_,
		_w16260_
	);
	LUT2 #(
		.INIT('h8)
	) name5749 (
		\wishbone_bd_ram_mem2_reg[169][20]/P0001 ,
		_w12722_,
		_w16261_
	);
	LUT2 #(
		.INIT('h8)
	) name5750 (
		\wishbone_bd_ram_mem2_reg[250][20]/P0001 ,
		_w13128_,
		_w16262_
	);
	LUT2 #(
		.INIT('h8)
	) name5751 (
		\wishbone_bd_ram_mem2_reg[38][20]/P0001 ,
		_w13182_,
		_w16263_
	);
	LUT2 #(
		.INIT('h8)
	) name5752 (
		\wishbone_bd_ram_mem2_reg[115][20]/P0001 ,
		_w13112_,
		_w16264_
	);
	LUT2 #(
		.INIT('h8)
	) name5753 (
		\wishbone_bd_ram_mem2_reg[154][20]/P0001 ,
		_w12962_,
		_w16265_
	);
	LUT2 #(
		.INIT('h8)
	) name5754 (
		\wishbone_bd_ram_mem2_reg[105][20]/P0001 ,
		_w12751_,
		_w16266_
	);
	LUT2 #(
		.INIT('h8)
	) name5755 (
		\wishbone_bd_ram_mem2_reg[152][20]/P0001 ,
		_w12966_,
		_w16267_
	);
	LUT2 #(
		.INIT('h8)
	) name5756 (
		\wishbone_bd_ram_mem2_reg[57][20]/P0001 ,
		_w13116_,
		_w16268_
	);
	LUT2 #(
		.INIT('h8)
	) name5757 (
		\wishbone_bd_ram_mem2_reg[101][20]/P0001 ,
		_w13192_,
		_w16269_
	);
	LUT2 #(
		.INIT('h8)
	) name5758 (
		\wishbone_bd_ram_mem2_reg[70][20]/P0001 ,
		_w12840_,
		_w16270_
	);
	LUT2 #(
		.INIT('h8)
	) name5759 (
		\wishbone_bd_ram_mem2_reg[150][20]/P0001 ,
		_w13136_,
		_w16271_
	);
	LUT2 #(
		.INIT('h8)
	) name5760 (
		\wishbone_bd_ram_mem2_reg[173][20]/P0001 ,
		_w12854_,
		_w16272_
	);
	LUT2 #(
		.INIT('h8)
	) name5761 (
		\wishbone_bd_ram_mem2_reg[142][20]/P0001 ,
		_w12928_,
		_w16273_
	);
	LUT2 #(
		.INIT('h8)
	) name5762 (
		\wishbone_bd_ram_mem2_reg[106][20]/P0001 ,
		_w12713_,
		_w16274_
	);
	LUT2 #(
		.INIT('h8)
	) name5763 (
		\wishbone_bd_ram_mem2_reg[148][20]/P0001 ,
		_w13000_,
		_w16275_
	);
	LUT2 #(
		.INIT('h8)
	) name5764 (
		\wishbone_bd_ram_mem2_reg[21][20]/P0001 ,
		_w12906_,
		_w16276_
	);
	LUT2 #(
		.INIT('h8)
	) name5765 (
		\wishbone_bd_ram_mem2_reg[201][20]/P0001 ,
		_w12822_,
		_w16277_
	);
	LUT2 #(
		.INIT('h8)
	) name5766 (
		\wishbone_bd_ram_mem2_reg[190][20]/P0001 ,
		_w12858_,
		_w16278_
	);
	LUT2 #(
		.INIT('h8)
	) name5767 (
		\wishbone_bd_ram_mem2_reg[22][20]/P0001 ,
		_w13110_,
		_w16279_
	);
	LUT2 #(
		.INIT('h8)
	) name5768 (
		\wishbone_bd_ram_mem2_reg[114][20]/P0001 ,
		_w13202_,
		_w16280_
	);
	LUT2 #(
		.INIT('h8)
	) name5769 (
		\wishbone_bd_ram_mem2_reg[168][20]/P0001 ,
		_w13208_,
		_w16281_
	);
	LUT2 #(
		.INIT('h8)
	) name5770 (
		\wishbone_bd_ram_mem2_reg[96][20]/P0001 ,
		_w12912_,
		_w16282_
	);
	LUT2 #(
		.INIT('h8)
	) name5771 (
		\wishbone_bd_ram_mem2_reg[247][20]/P0001 ,
		_w12818_,
		_w16283_
	);
	LUT2 #(
		.INIT('h8)
	) name5772 (
		\wishbone_bd_ram_mem2_reg[124][20]/P0001 ,
		_w13058_,
		_w16284_
	);
	LUT2 #(
		.INIT('h8)
	) name5773 (
		\wishbone_bd_ram_mem2_reg[71][20]/P0001 ,
		_w12798_,
		_w16285_
	);
	LUT2 #(
		.INIT('h8)
	) name5774 (
		\wishbone_bd_ram_mem2_reg[223][20]/P0001 ,
		_w12838_,
		_w16286_
	);
	LUT2 #(
		.INIT('h8)
	) name5775 (
		\wishbone_bd_ram_mem2_reg[242][20]/P0001 ,
		_w12932_,
		_w16287_
	);
	LUT2 #(
		.INIT('h8)
	) name5776 (
		\wishbone_bd_ram_mem2_reg[160][20]/P0001 ,
		_w12872_,
		_w16288_
	);
	LUT2 #(
		.INIT('h8)
	) name5777 (
		\wishbone_bd_ram_mem2_reg[92][20]/P0001 ,
		_w13010_,
		_w16289_
	);
	LUT2 #(
		.INIT('h8)
	) name5778 (
		\wishbone_bd_ram_mem2_reg[210][20]/P0001 ,
		_w12924_,
		_w16290_
	);
	LUT2 #(
		.INIT('h8)
	) name5779 (
		\wishbone_bd_ram_mem2_reg[254][20]/P0001 ,
		_w12892_,
		_w16291_
	);
	LUT2 #(
		.INIT('h8)
	) name5780 (
		\wishbone_bd_ram_mem2_reg[198][20]/P0001 ,
		_w12832_,
		_w16292_
	);
	LUT2 #(
		.INIT('h8)
	) name5781 (
		\wishbone_bd_ram_mem2_reg[128][20]/P0001 ,
		_w12793_,
		_w16293_
	);
	LUT2 #(
		.INIT('h8)
	) name5782 (
		\wishbone_bd_ram_mem2_reg[112][20]/P0001 ,
		_w12733_,
		_w16294_
	);
	LUT2 #(
		.INIT('h8)
	) name5783 (
		\wishbone_bd_ram_mem2_reg[44][20]/P0001 ,
		_w12896_,
		_w16295_
	);
	LUT2 #(
		.INIT('h8)
	) name5784 (
		\wishbone_bd_ram_mem2_reg[53][20]/P0001 ,
		_w13020_,
		_w16296_
	);
	LUT2 #(
		.INIT('h8)
	) name5785 (
		\wishbone_bd_ram_mem2_reg[164][20]/P0001 ,
		_w12876_,
		_w16297_
	);
	LUT2 #(
		.INIT('h8)
	) name5786 (
		\wishbone_bd_ram_mem2_reg[215][20]/P0001 ,
		_w12974_,
		_w16298_
	);
	LUT2 #(
		.INIT('h8)
	) name5787 (
		\wishbone_bd_ram_mem2_reg[4][20]/P0001 ,
		_w12666_,
		_w16299_
	);
	LUT2 #(
		.INIT('h8)
	) name5788 (
		\wishbone_bd_ram_mem2_reg[9][20]/P0001 ,
		_w12808_,
		_w16300_
	);
	LUT2 #(
		.INIT('h8)
	) name5789 (
		\wishbone_bd_ram_mem2_reg[135][20]/P0001 ,
		_w13124_,
		_w16301_
	);
	LUT2 #(
		.INIT('h8)
	) name5790 (
		\wishbone_bd_ram_mem2_reg[0][20]/P0001 ,
		_w12717_,
		_w16302_
	);
	LUT2 #(
		.INIT('h8)
	) name5791 (
		\wishbone_bd_ram_mem2_reg[19][20]/P0001 ,
		_w13012_,
		_w16303_
	);
	LUT2 #(
		.INIT('h8)
	) name5792 (
		\wishbone_bd_ram_mem2_reg[211][20]/P0001 ,
		_w13166_,
		_w16304_
	);
	LUT2 #(
		.INIT('h8)
	) name5793 (
		\wishbone_bd_ram_mem2_reg[235][20]/P0001 ,
		_w12696_,
		_w16305_
	);
	LUT2 #(
		.INIT('h8)
	) name5794 (
		\wishbone_bd_ram_mem2_reg[119][20]/P0001 ,
		_w13048_,
		_w16306_
	);
	LUT2 #(
		.INIT('h8)
	) name5795 (
		\wishbone_bd_ram_mem2_reg[10][20]/P0001 ,
		_w13172_,
		_w16307_
	);
	LUT2 #(
		.INIT('h8)
	) name5796 (
		\wishbone_bd_ram_mem2_reg[65][20]/P0001 ,
		_w13176_,
		_w16308_
	);
	LUT2 #(
		.INIT('h8)
	) name5797 (
		\wishbone_bd_ram_mem2_reg[165][20]/P0001 ,
		_w13044_,
		_w16309_
	);
	LUT2 #(
		.INIT('h8)
	) name5798 (
		\wishbone_bd_ram_mem2_reg[134][20]/P0001 ,
		_w12763_,
		_w16310_
	);
	LUT2 #(
		.INIT('h8)
	) name5799 (
		\wishbone_bd_ram_mem2_reg[146][20]/P0001 ,
		_w13060_,
		_w16311_
	);
	LUT2 #(
		.INIT('h8)
	) name5800 (
		\wishbone_bd_ram_mem2_reg[99][20]/P0001 ,
		_w13038_,
		_w16312_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		\wishbone_bd_ram_mem2_reg[133][20]/P0001 ,
		_w12761_,
		_w16313_
	);
	LUT2 #(
		.INIT('h8)
	) name5802 (
		\wishbone_bd_ram_mem2_reg[43][20]/P0001 ,
		_w13200_,
		_w16314_
	);
	LUT2 #(
		.INIT('h8)
	) name5803 (
		\wishbone_bd_ram_mem2_reg[34][20]/P0001 ,
		_w12930_,
		_w16315_
	);
	LUT2 #(
		.INIT('h8)
	) name5804 (
		\wishbone_bd_ram_mem2_reg[67][20]/P0001 ,
		_w13134_,
		_w16316_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		\wishbone_bd_ram_mem2_reg[113][20]/P0001 ,
		_w13026_,
		_w16317_
	);
	LUT2 #(
		.INIT('h8)
	) name5806 (
		\wishbone_bd_ram_mem2_reg[140][20]/P0001 ,
		_w12894_,
		_w16318_
	);
	LUT2 #(
		.INIT('h8)
	) name5807 (
		\wishbone_bd_ram_mem2_reg[245][20]/P0001 ,
		_w13022_,
		_w16319_
	);
	LUT2 #(
		.INIT('h8)
	) name5808 (
		\wishbone_bd_ram_mem2_reg[87][20]/P0001 ,
		_w13154_,
		_w16320_
	);
	LUT2 #(
		.INIT('h8)
	) name5809 (
		\wishbone_bd_ram_mem2_reg[194][20]/P0001 ,
		_w12772_,
		_w16321_
	);
	LUT2 #(
		.INIT('h8)
	) name5810 (
		\wishbone_bd_ram_mem2_reg[32][20]/P0001 ,
		_w13120_,
		_w16322_
	);
	LUT2 #(
		.INIT('h8)
	) name5811 (
		\wishbone_bd_ram_mem2_reg[29][20]/P0001 ,
		_w12952_,
		_w16323_
	);
	LUT2 #(
		.INIT('h8)
	) name5812 (
		\wishbone_bd_ram_mem2_reg[252][20]/P0001 ,
		_w13080_,
		_w16324_
	);
	LUT2 #(
		.INIT('h8)
	) name5813 (
		\wishbone_bd_ram_mem2_reg[3][20]/P0001 ,
		_w12866_,
		_w16325_
	);
	LUT2 #(
		.INIT('h8)
	) name5814 (
		\wishbone_bd_ram_mem2_reg[180][20]/P0001 ,
		_w12791_,
		_w16326_
	);
	LUT2 #(
		.INIT('h8)
	) name5815 (
		\wishbone_bd_ram_mem2_reg[83][20]/P0001 ,
		_w12916_,
		_w16327_
	);
	LUT2 #(
		.INIT('h8)
	) name5816 (
		\wishbone_bd_ram_mem2_reg[41][20]/P0001 ,
		_w13052_,
		_w16328_
	);
	LUT2 #(
		.INIT('h8)
	) name5817 (
		\wishbone_bd_ram_mem2_reg[33][20]/P0001 ,
		_w12980_,
		_w16329_
	);
	LUT2 #(
		.INIT('h8)
	) name5818 (
		\wishbone_bd_ram_mem2_reg[30][20]/P0001 ,
		_w13104_,
		_w16330_
	);
	LUT2 #(
		.INIT('h8)
	) name5819 (
		\wishbone_bd_ram_mem2_reg[5][20]/P0001 ,
		_w12878_,
		_w16331_
	);
	LUT2 #(
		.INIT('h8)
	) name5820 (
		\wishbone_bd_ram_mem2_reg[158][20]/P0001 ,
		_w12898_,
		_w16332_
	);
	LUT2 #(
		.INIT('h8)
	) name5821 (
		\wishbone_bd_ram_mem2_reg[8][20]/P0001 ,
		_w12920_,
		_w16333_
	);
	LUT2 #(
		.INIT('h8)
	) name5822 (
		\wishbone_bd_ram_mem2_reg[89][20]/P0001 ,
		_w12964_,
		_w16334_
	);
	LUT2 #(
		.INIT('h8)
	) name5823 (
		\wishbone_bd_ram_mem2_reg[204][20]/P0001 ,
		_w13162_,
		_w16335_
	);
	LUT2 #(
		.INIT('h8)
	) name5824 (
		\wishbone_bd_ram_mem2_reg[82][20]/P0001 ,
		_w12942_,
		_w16336_
	);
	LUT2 #(
		.INIT('h8)
	) name5825 (
		\wishbone_bd_ram_mem2_reg[202][20]/P0001 ,
		_w12870_,
		_w16337_
	);
	LUT2 #(
		.INIT('h8)
	) name5826 (
		\wishbone_bd_ram_mem2_reg[18][20]/P0001 ,
		_w12679_,
		_w16338_
	);
	LUT2 #(
		.INIT('h8)
	) name5827 (
		\wishbone_bd_ram_mem2_reg[108][20]/P0001 ,
		_w13156_,
		_w16339_
	);
	LUT2 #(
		.INIT('h8)
	) name5828 (
		\wishbone_bd_ram_mem2_reg[219][20]/P0001 ,
		_w12806_,
		_w16340_
	);
	LUT2 #(
		.INIT('h8)
	) name5829 (
		\wishbone_bd_ram_mem2_reg[189][20]/P0001 ,
		_w13042_,
		_w16341_
	);
	LUT2 #(
		.INIT('h8)
	) name5830 (
		\wishbone_bd_ram_mem2_reg[217][20]/P0001 ,
		_w13188_,
		_w16342_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		\wishbone_bd_ram_mem2_reg[26][20]/P0001 ,
		_w12699_,
		_w16343_
	);
	LUT2 #(
		.INIT('h8)
	) name5832 (
		\wishbone_bd_ram_mem2_reg[157][20]/P0001 ,
		_w12926_,
		_w16344_
	);
	LUT2 #(
		.INIT('h8)
	) name5833 (
		\wishbone_bd_ram_mem2_reg[90][20]/P0001 ,
		_w12978_,
		_w16345_
	);
	LUT2 #(
		.INIT('h8)
	) name5834 (
		\wishbone_bd_ram_mem2_reg[45][20]/P0001 ,
		_w12908_,
		_w16346_
	);
	LUT2 #(
		.INIT('h8)
	) name5835 (
		\wishbone_bd_ram_mem2_reg[125][20]/P0001 ,
		_w12956_,
		_w16347_
	);
	LUT2 #(
		.INIT('h8)
	) name5836 (
		\wishbone_bd_ram_mem2_reg[40][20]/P0001 ,
		_w13132_,
		_w16348_
	);
	LUT2 #(
		.INIT('h8)
	) name5837 (
		\wishbone_bd_ram_mem2_reg[229][20]/P0001 ,
		_w12711_,
		_w16349_
	);
	LUT2 #(
		.INIT('h8)
	) name5838 (
		\wishbone_bd_ram_mem2_reg[73][20]/P0001 ,
		_w12918_,
		_w16350_
	);
	LUT2 #(
		.INIT('h8)
	) name5839 (
		\wishbone_bd_ram_mem2_reg[236][20]/P0001 ,
		_w12731_,
		_w16351_
	);
	LUT2 #(
		.INIT('h8)
	) name5840 (
		\wishbone_bd_ram_mem2_reg[222][20]/P0001 ,
		_w13094_,
		_w16352_
	);
	LUT2 #(
		.INIT('h8)
	) name5841 (
		\wishbone_bd_ram_mem2_reg[137][20]/P0001 ,
		_w13168_,
		_w16353_
	);
	LUT2 #(
		.INIT('h8)
	) name5842 (
		\wishbone_bd_ram_mem2_reg[126][20]/P0001 ,
		_w13218_,
		_w16354_
	);
	LUT2 #(
		.INIT('h8)
	) name5843 (
		\wishbone_bd_ram_mem2_reg[109][20]/P0001 ,
		_w12888_,
		_w16355_
	);
	LUT2 #(
		.INIT('h8)
	) name5844 (
		\wishbone_bd_ram_mem2_reg[244][20]/P0001 ,
		_w12747_,
		_w16356_
	);
	LUT2 #(
		.INIT('h8)
	) name5845 (
		\wishbone_bd_ram_mem2_reg[193][20]/P0001 ,
		_w13056_,
		_w16357_
	);
	LUT2 #(
		.INIT('h8)
	) name5846 (
		\wishbone_bd_ram_mem2_reg[172][20]/P0001 ,
		_w12944_,
		_w16358_
	);
	LUT2 #(
		.INIT('h8)
	) name5847 (
		\wishbone_bd_ram_mem2_reg[116][20]/P0001 ,
		_w12998_,
		_w16359_
	);
	LUT2 #(
		.INIT('h8)
	) name5848 (
		\wishbone_bd_ram_mem2_reg[192][20]/P0001 ,
		_w12938_,
		_w16360_
	);
	LUT2 #(
		.INIT('h8)
	) name5849 (
		\wishbone_bd_ram_mem2_reg[232][20]/P0001 ,
		_w12758_,
		_w16361_
	);
	LUT2 #(
		.INIT('h8)
	) name5850 (
		\wishbone_bd_ram_mem2_reg[11][20]/P0001 ,
		_w13194_,
		_w16362_
	);
	LUT2 #(
		.INIT('h8)
	) name5851 (
		\wishbone_bd_ram_mem2_reg[213][20]/P0001 ,
		_w13002_,
		_w16363_
	);
	LUT2 #(
		.INIT('h8)
	) name5852 (
		\wishbone_bd_ram_mem2_reg[61][20]/P0001 ,
		_w12725_,
		_w16364_
	);
	LUT2 #(
		.INIT('h8)
	) name5853 (
		\wishbone_bd_ram_mem2_reg[6][20]/P0001 ,
		_w12968_,
		_w16365_
	);
	LUT2 #(
		.INIT('h8)
	) name5854 (
		\wishbone_bd_ram_mem2_reg[191][20]/P0001 ,
		_w13034_,
		_w16366_
	);
	LUT2 #(
		.INIT('h8)
	) name5855 (
		\wishbone_bd_ram_mem2_reg[17][20]/P0001 ,
		_w12848_,
		_w16367_
	);
	LUT2 #(
		.INIT('h8)
	) name5856 (
		\wishbone_bd_ram_mem2_reg[199][20]/P0001 ,
		_w12768_,
		_w16368_
	);
	LUT2 #(
		.INIT('h8)
	) name5857 (
		\wishbone_bd_ram_mem2_reg[78][20]/P0001 ,
		_w12874_,
		_w16369_
	);
	LUT2 #(
		.INIT('h8)
	) name5858 (
		\wishbone_bd_ram_mem2_reg[251][20]/P0001 ,
		_w13054_,
		_w16370_
	);
	LUT2 #(
		.INIT('h8)
	) name5859 (
		\wishbone_bd_ram_mem2_reg[48][20]/P0001 ,
		_w12970_,
		_w16371_
	);
	LUT2 #(
		.INIT('h8)
	) name5860 (
		\wishbone_bd_ram_mem2_reg[224][20]/P0001 ,
		_w12902_,
		_w16372_
	);
	LUT2 #(
		.INIT('h8)
	) name5861 (
		\wishbone_bd_ram_mem2_reg[138][20]/P0001 ,
		_w12958_,
		_w16373_
	);
	LUT2 #(
		.INIT('h8)
	) name5862 (
		\wishbone_bd_ram_mem2_reg[221][20]/P0001 ,
		_w12802_,
		_w16374_
	);
	LUT2 #(
		.INIT('h8)
	) name5863 (
		\wishbone_bd_ram_mem2_reg[174][20]/P0001 ,
		_w12972_,
		_w16375_
	);
	LUT2 #(
		.INIT('h8)
	) name5864 (
		\wishbone_bd_ram_mem2_reg[68][20]/P0001 ,
		_w12946_,
		_w16376_
	);
	LUT2 #(
		.INIT('h8)
	) name5865 (
		\wishbone_bd_ram_mem2_reg[248][20]/P0001 ,
		_w12789_,
		_w16377_
	);
	LUT2 #(
		.INIT('h8)
	) name5866 (
		\wishbone_bd_ram_mem2_reg[230][20]/P0001 ,
		_w13036_,
		_w16378_
	);
	LUT2 #(
		.INIT('h8)
	) name5867 (
		\wishbone_bd_ram_mem2_reg[35][20]/P0001 ,
		_w12703_,
		_w16379_
	);
	LUT2 #(
		.INIT('h8)
	) name5868 (
		\wishbone_bd_ram_mem2_reg[209][20]/P0001 ,
		_w13152_,
		_w16380_
	);
	LUT2 #(
		.INIT('h8)
	) name5869 (
		\wishbone_bd_ram_mem2_reg[228][20]/P0001 ,
		_w12765_,
		_w16381_
	);
	LUT2 #(
		.INIT('h8)
	) name5870 (
		\wishbone_bd_ram_mem2_reg[246][20]/P0001 ,
		_w13076_,
		_w16382_
	);
	LUT2 #(
		.INIT('h8)
	) name5871 (
		\wishbone_bd_ram_mem2_reg[81][20]/P0001 ,
		_w12950_,
		_w16383_
	);
	LUT2 #(
		.INIT('h8)
	) name5872 (
		\wishbone_bd_ram_mem2_reg[216][20]/P0001 ,
		_w13028_,
		_w16384_
	);
	LUT2 #(
		.INIT('h8)
	) name5873 (
		\wishbone_bd_ram_mem2_reg[2][20]/P0001 ,
		_w13088_,
		_w16385_
	);
	LUT2 #(
		.INIT('h8)
	) name5874 (
		\wishbone_bd_ram_mem2_reg[178][20]/P0001 ,
		_w12886_,
		_w16386_
	);
	LUT2 #(
		.INIT('h8)
	) name5875 (
		\wishbone_bd_ram_mem2_reg[12][20]/P0001 ,
		_w13118_,
		_w16387_
	);
	LUT2 #(
		.INIT('h8)
	) name5876 (
		\wishbone_bd_ram_mem2_reg[176][20]/P0001 ,
		_w12868_,
		_w16388_
	);
	LUT2 #(
		.INIT('h8)
	) name5877 (
		\wishbone_bd_ram_mem2_reg[59][20]/P0001 ,
		_w12780_,
		_w16389_
	);
	LUT2 #(
		.INIT('h8)
	) name5878 (
		\wishbone_bd_ram_mem2_reg[226][20]/P0001 ,
		_w13138_,
		_w16390_
	);
	LUT2 #(
		.INIT('h8)
	) name5879 (
		\wishbone_bd_ram_mem2_reg[143][20]/P0001 ,
		_w12922_,
		_w16391_
	);
	LUT2 #(
		.INIT('h8)
	) name5880 (
		\wishbone_bd_ram_mem2_reg[93][20]/P0001 ,
		_w13016_,
		_w16392_
	);
	LUT2 #(
		.INIT('h8)
	) name5881 (
		\wishbone_bd_ram_mem2_reg[86][20]/P0001 ,
		_w12735_,
		_w16393_
	);
	LUT2 #(
		.INIT('h8)
	) name5882 (
		\wishbone_bd_ram_mem2_reg[63][20]/P0001 ,
		_w12850_,
		_w16394_
	);
	LUT2 #(
		.INIT('h8)
	) name5883 (
		\wishbone_bd_ram_mem2_reg[77][20]/P0001 ,
		_w12982_,
		_w16395_
	);
	LUT2 #(
		.INIT('h8)
	) name5884 (
		\wishbone_bd_ram_mem2_reg[98][20]/P0001 ,
		_w12816_,
		_w16396_
	);
	LUT2 #(
		.INIT('h8)
	) name5885 (
		\wishbone_bd_ram_mem2_reg[123][20]/P0001 ,
		_w13114_,
		_w16397_
	);
	LUT2 #(
		.INIT('h8)
	) name5886 (
		\wishbone_bd_ram_mem2_reg[171][20]/P0001 ,
		_w12910_,
		_w16398_
	);
	LUT2 #(
		.INIT('h8)
	) name5887 (
		\wishbone_bd_ram_mem2_reg[131][20]/P0001 ,
		_w12852_,
		_w16399_
	);
	LUT2 #(
		.INIT('h8)
	) name5888 (
		\wishbone_bd_ram_mem2_reg[74][20]/P0001 ,
		_w12812_,
		_w16400_
	);
	LUT2 #(
		.INIT('h8)
	) name5889 (
		\wishbone_bd_ram_mem2_reg[136][20]/P0001 ,
		_w13064_,
		_w16401_
	);
	LUT2 #(
		.INIT('h8)
	) name5890 (
		\wishbone_bd_ram_mem2_reg[182][20]/P0001 ,
		_w12820_,
		_w16402_
	);
	LUT2 #(
		.INIT('h8)
	) name5891 (
		\wishbone_bd_ram_mem2_reg[153][20]/P0001 ,
		_w12890_,
		_w16403_
	);
	LUT2 #(
		.INIT('h8)
	) name5892 (
		\wishbone_bd_ram_mem2_reg[227][20]/P0001 ,
		_w12936_,
		_w16404_
	);
	LUT2 #(
		.INIT('h8)
	) name5893 (
		\wishbone_bd_ram_mem2_reg[122][20]/P0001 ,
		_w13130_,
		_w16405_
	);
	LUT2 #(
		.INIT('h8)
	) name5894 (
		\wishbone_bd_ram_mem2_reg[167][20]/P0001 ,
		_w12986_,
		_w16406_
	);
	LUT2 #(
		.INIT('h8)
	) name5895 (
		\wishbone_bd_ram_mem2_reg[132][20]/P0001 ,
		_w12992_,
		_w16407_
	);
	LUT2 #(
		.INIT('h8)
	) name5896 (
		\wishbone_bd_ram_mem2_reg[58][20]/P0001 ,
		_w13070_,
		_w16408_
	);
	LUT2 #(
		.INIT('h8)
	) name5897 (
		\wishbone_bd_ram_mem2_reg[208][20]/P0001 ,
		_w13032_,
		_w16409_
	);
	LUT2 #(
		.INIT('h8)
	) name5898 (
		\wishbone_bd_ram_mem2_reg[187][20]/P0001 ,
		_w13196_,
		_w16410_
	);
	LUT2 #(
		.INIT('h8)
	) name5899 (
		\wishbone_bd_ram_mem2_reg[13][20]/P0001 ,
		_w13178_,
		_w16411_
	);
	LUT2 #(
		.INIT('h8)
	) name5900 (
		\wishbone_bd_ram_mem2_reg[52][20]/P0001 ,
		_w13082_,
		_w16412_
	);
	LUT2 #(
		.INIT('h8)
	) name5901 (
		\wishbone_bd_ram_mem2_reg[175][20]/P0001 ,
		_w13126_,
		_w16413_
	);
	LUT2 #(
		.INIT('h8)
	) name5902 (
		\wishbone_bd_ram_mem2_reg[156][20]/P0001 ,
		_w13190_,
		_w16414_
	);
	LUT2 #(
		.INIT('h8)
	) name5903 (
		\wishbone_bd_ram_mem2_reg[241][20]/P0001 ,
		_w13006_,
		_w16415_
	);
	LUT2 #(
		.INIT('h8)
	) name5904 (
		\wishbone_bd_ram_mem2_reg[159][20]/P0001 ,
		_w12774_,
		_w16416_
	);
	LUT2 #(
		.INIT('h8)
	) name5905 (
		\wishbone_bd_ram_mem2_reg[220][20]/P0001 ,
		_w13066_,
		_w16417_
	);
	LUT2 #(
		.INIT('h8)
	) name5906 (
		\wishbone_bd_ram_mem2_reg[218][20]/P0001 ,
		_w13206_,
		_w16418_
	);
	LUT2 #(
		.INIT('h8)
	) name5907 (
		\wishbone_bd_ram_mem2_reg[104][20]/P0001 ,
		_w13148_,
		_w16419_
	);
	LUT2 #(
		.INIT('h8)
	) name5908 (
		\wishbone_bd_ram_mem2_reg[183][20]/P0001 ,
		_w12787_,
		_w16420_
	);
	LUT2 #(
		.INIT('h8)
	) name5909 (
		\wishbone_bd_ram_mem2_reg[55][20]/P0001 ,
		_w12785_,
		_w16421_
	);
	LUT2 #(
		.INIT('h8)
	) name5910 (
		\wishbone_bd_ram_mem2_reg[50][20]/P0001 ,
		_w13150_,
		_w16422_
	);
	LUT2 #(
		.INIT('h8)
	) name5911 (
		\wishbone_bd_ram_mem2_reg[155][20]/P0001 ,
		_w13122_,
		_w16423_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		\wishbone_bd_ram_mem2_reg[184][20]/P0001 ,
		_w13062_,
		_w16424_
	);
	LUT2 #(
		.INIT('h8)
	) name5913 (
		\wishbone_bd_ram_mem2_reg[110][20]/P0001 ,
		_w13046_,
		_w16425_
	);
	LUT2 #(
		.INIT('h8)
	) name5914 (
		\wishbone_bd_ram_mem2_reg[28][20]/P0001 ,
		_w13170_,
		_w16426_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		\wishbone_bd_ram_mem2_reg[91][20]/P0001 ,
		_w13074_,
		_w16427_
	);
	LUT2 #(
		.INIT('h8)
	) name5916 (
		\wishbone_bd_ram_mem2_reg[240][20]/P0001 ,
		_w12864_,
		_w16428_
	);
	LUT2 #(
		.INIT('h8)
	) name5917 (
		\wishbone_bd_ram_mem2_reg[243][20]/P0001 ,
		_w12804_,
		_w16429_
	);
	LUT2 #(
		.INIT('h8)
	) name5918 (
		\wishbone_bd_ram_mem2_reg[24][20]/P0001 ,
		_w13084_,
		_w16430_
	);
	LUT2 #(
		.INIT('h8)
	) name5919 (
		\wishbone_bd_ram_mem2_reg[103][20]/P0001 ,
		_w12846_,
		_w16431_
	);
	LUT2 #(
		.INIT('h8)
	) name5920 (
		\wishbone_bd_ram_mem2_reg[7][20]/P0001 ,
		_w12728_,
		_w16432_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		\wishbone_bd_ram_mem2_reg[97][20]/P0001 ,
		_w13096_,
		_w16433_
	);
	LUT2 #(
		.INIT('h8)
	) name5922 (
		\wishbone_bd_ram_mem2_reg[31][20]/P0001 ,
		_w13198_,
		_w16434_
	);
	LUT2 #(
		.INIT('h8)
	) name5923 (
		\wishbone_bd_ram_mem2_reg[54][20]/P0001 ,
		_w12770_,
		_w16435_
	);
	LUT2 #(
		.INIT('h8)
	) name5924 (
		\wishbone_bd_ram_mem2_reg[27][20]/P0001 ,
		_w12880_,
		_w16436_
	);
	LUT2 #(
		.INIT('h8)
	) name5925 (
		\wishbone_bd_ram_mem2_reg[170][20]/P0001 ,
		_w13030_,
		_w16437_
	);
	LUT2 #(
		.INIT('h8)
	) name5926 (
		\wishbone_bd_ram_mem2_reg[195][20]/P0001 ,
		_w13144_,
		_w16438_
	);
	LUT2 #(
		.INIT('h8)
	) name5927 (
		\wishbone_bd_ram_mem2_reg[233][20]/P0001 ,
		_w12836_,
		_w16439_
	);
	LUT2 #(
		.INIT('h8)
	) name5928 (
		\wishbone_bd_ram_mem2_reg[185][20]/P0001 ,
		_w12940_,
		_w16440_
	);
	LUT2 #(
		.INIT('h8)
	) name5929 (
		\wishbone_bd_ram_mem2_reg[1][20]/P0001 ,
		_w13014_,
		_w16441_
	);
	LUT2 #(
		.INIT('h8)
	) name5930 (
		\wishbone_bd_ram_mem2_reg[23][20]/P0001 ,
		_w13008_,
		_w16442_
	);
	LUT2 #(
		.INIT('h8)
	) name5931 (
		\wishbone_bd_ram_mem2_reg[129][20]/P0001 ,
		_w12776_,
		_w16443_
	);
	LUT2 #(
		.INIT('h8)
	) name5932 (
		\wishbone_bd_ram_mem2_reg[84][20]/P0001 ,
		_w12934_,
		_w16444_
	);
	LUT2 #(
		.INIT('h8)
	) name5933 (
		\wishbone_bd_ram_mem2_reg[102][20]/P0001 ,
		_w12685_,
		_w16445_
	);
	LUT2 #(
		.INIT('h8)
	) name5934 (
		\wishbone_bd_ram_mem2_reg[139][20]/P0001 ,
		_w12814_,
		_w16446_
	);
	LUT2 #(
		.INIT('h8)
	) name5935 (
		\wishbone_bd_ram_mem2_reg[66][20]/P0001 ,
		_w12824_,
		_w16447_
	);
	LUT2 #(
		.INIT('h8)
	) name5936 (
		\wishbone_bd_ram_mem2_reg[205][20]/P0001 ,
		_w13068_,
		_w16448_
	);
	LUT2 #(
		.INIT('h8)
	) name5937 (
		\wishbone_bd_ram_mem2_reg[130][20]/P0001 ,
		_w12914_,
		_w16449_
	);
	LUT2 #(
		.INIT('h8)
	) name5938 (
		\wishbone_bd_ram_mem2_reg[163][20]/P0001 ,
		_w12882_,
		_w16450_
	);
	LUT2 #(
		.INIT('h8)
	) name5939 (
		\wishbone_bd_ram_mem2_reg[253][20]/P0001 ,
		_w13100_,
		_w16451_
	);
	LUT2 #(
		.INIT('h8)
	) name5940 (
		\wishbone_bd_ram_mem2_reg[69][20]/P0001 ,
		_w12738_,
		_w16452_
	);
	LUT2 #(
		.INIT('h8)
	) name5941 (
		\wishbone_bd_ram_mem2_reg[197][20]/P0001 ,
		_w12834_,
		_w16453_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		\wishbone_bd_ram_mem2_reg[72][20]/P0001 ,
		_w12810_,
		_w16454_
	);
	LUT2 #(
		.INIT('h8)
	) name5943 (
		\wishbone_bd_ram_mem2_reg[94][20]/P0001 ,
		_w13186_,
		_w16455_
	);
	LUT2 #(
		.INIT('h8)
	) name5944 (
		\wishbone_bd_ram_mem2_reg[60][20]/P0001 ,
		_w13204_,
		_w16456_
	);
	LUT2 #(
		.INIT('h8)
	) name5945 (
		\wishbone_bd_ram_mem2_reg[255][20]/P0001 ,
		_w13072_,
		_w16457_
	);
	LUT2 #(
		.INIT('h8)
	) name5946 (
		\wishbone_bd_ram_mem2_reg[249][20]/P0001 ,
		_w12900_,
		_w16458_
	);
	LUT2 #(
		.INIT('h8)
	) name5947 (
		\wishbone_bd_ram_mem2_reg[42][20]/P0001 ,
		_w12842_,
		_w16459_
	);
	LUT2 #(
		.INIT('h8)
	) name5948 (
		\wishbone_bd_ram_mem2_reg[179][20]/P0001 ,
		_w13050_,
		_w16460_
	);
	LUT2 #(
		.INIT('h8)
	) name5949 (
		\wishbone_bd_ram_mem2_reg[49][20]/P0001 ,
		_w12994_,
		_w16461_
	);
	LUT2 #(
		.INIT('h8)
	) name5950 (
		\wishbone_bd_ram_mem2_reg[117][20]/P0001 ,
		_w12715_,
		_w16462_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		\wishbone_bd_ram_mem2_reg[162][20]/P0001 ,
		_w13098_,
		_w16463_
	);
	LUT2 #(
		.INIT('h8)
	) name5952 (
		\wishbone_bd_ram_mem2_reg[186][20]/P0001 ,
		_w12783_,
		_w16464_
	);
	LUT2 #(
		.INIT('h8)
	) name5953 (
		\wishbone_bd_ram_mem2_reg[47][20]/P0001 ,
		_w12904_,
		_w16465_
	);
	LUT2 #(
		.INIT('h8)
	) name5954 (
		\wishbone_bd_ram_mem2_reg[151][20]/P0001 ,
		_w13142_,
		_w16466_
	);
	LUT2 #(
		.INIT('h8)
	) name5955 (
		\wishbone_bd_ram_mem2_reg[95][20]/P0001 ,
		_w12844_,
		_w16467_
	);
	LUT2 #(
		.INIT('h8)
	) name5956 (
		\wishbone_bd_ram_mem2_reg[214][20]/P0001 ,
		_w12984_,
		_w16468_
	);
	LUT2 #(
		.INIT('h8)
	) name5957 (
		\wishbone_bd_ram_mem2_reg[107][20]/P0001 ,
		_w12749_,
		_w16469_
	);
	LUT2 #(
		.INIT('h8)
	) name5958 (
		\wishbone_bd_ram_mem2_reg[188][20]/P0001 ,
		_w12948_,
		_w16470_
	);
	LUT2 #(
		.INIT('h8)
	) name5959 (
		\wishbone_bd_ram_mem2_reg[25][20]/P0001 ,
		_w13108_,
		_w16471_
	);
	LUT2 #(
		.INIT('h8)
	) name5960 (
		\wishbone_bd_ram_mem2_reg[75][20]/P0001 ,
		_w12826_,
		_w16472_
	);
	LUT2 #(
		.INIT('h8)
	) name5961 (
		\wishbone_bd_ram_mem2_reg[161][20]/P0001 ,
		_w12754_,
		_w16473_
	);
	LUT2 #(
		.INIT('h8)
	) name5962 (
		\wishbone_bd_ram_mem2_reg[36][20]/P0001 ,
		_w12800_,
		_w16474_
	);
	LUT2 #(
		.INIT('h8)
	) name5963 (
		\wishbone_bd_ram_mem2_reg[51][20]/P0001 ,
		_w13024_,
		_w16475_
	);
	LUT2 #(
		.INIT('h8)
	) name5964 (
		\wishbone_bd_ram_mem2_reg[46][20]/P0001 ,
		_w12884_,
		_w16476_
	);
	LUT2 #(
		.INIT('h8)
	) name5965 (
		\wishbone_bd_ram_mem2_reg[207][20]/P0001 ,
		_w13180_,
		_w16477_
	);
	LUT2 #(
		.INIT('h8)
	) name5966 (
		\wishbone_bd_ram_mem2_reg[212][20]/P0001 ,
		_w12796_,
		_w16478_
	);
	LUT2 #(
		.INIT('h8)
	) name5967 (
		\wishbone_bd_ram_mem2_reg[62][20]/P0001 ,
		_w12673_,
		_w16479_
	);
	LUT2 #(
		.INIT('h8)
	) name5968 (
		\wishbone_bd_ram_mem2_reg[88][20]/P0001 ,
		_w12860_,
		_w16480_
	);
	LUT2 #(
		.INIT('h8)
	) name5969 (
		\wishbone_bd_ram_mem2_reg[196][20]/P0001 ,
		_w13090_,
		_w16481_
	);
	LUT2 #(
		.INIT('h8)
	) name5970 (
		\wishbone_bd_ram_mem2_reg[238][20]/P0001 ,
		_w13160_,
		_w16482_
	);
	LUT2 #(
		.INIT('h8)
	) name5971 (
		\wishbone_bd_ram_mem2_reg[181][20]/P0001 ,
		_w12828_,
		_w16483_
	);
	LUT2 #(
		.INIT('h8)
	) name5972 (
		\wishbone_bd_ram_mem2_reg[80][20]/P0001 ,
		_w12689_,
		_w16484_
	);
	LUT2 #(
		.INIT('h8)
	) name5973 (
		\wishbone_bd_ram_mem2_reg[14][20]/P0001 ,
		_w13086_,
		_w16485_
	);
	LUT2 #(
		.INIT('h8)
	) name5974 (
		\wishbone_bd_ram_mem2_reg[200][20]/P0001 ,
		_w12988_,
		_w16486_
	);
	LUT2 #(
		.INIT('h8)
	) name5975 (
		\wishbone_bd_ram_mem2_reg[141][20]/P0001 ,
		_w13004_,
		_w16487_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		_w16232_,
		_w16233_,
		_w16488_
	);
	LUT2 #(
		.INIT('h1)
	) name5977 (
		_w16234_,
		_w16235_,
		_w16489_
	);
	LUT2 #(
		.INIT('h1)
	) name5978 (
		_w16236_,
		_w16237_,
		_w16490_
	);
	LUT2 #(
		.INIT('h1)
	) name5979 (
		_w16238_,
		_w16239_,
		_w16491_
	);
	LUT2 #(
		.INIT('h1)
	) name5980 (
		_w16240_,
		_w16241_,
		_w16492_
	);
	LUT2 #(
		.INIT('h1)
	) name5981 (
		_w16242_,
		_w16243_,
		_w16493_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w16244_,
		_w16245_,
		_w16494_
	);
	LUT2 #(
		.INIT('h1)
	) name5983 (
		_w16246_,
		_w16247_,
		_w16495_
	);
	LUT2 #(
		.INIT('h1)
	) name5984 (
		_w16248_,
		_w16249_,
		_w16496_
	);
	LUT2 #(
		.INIT('h1)
	) name5985 (
		_w16250_,
		_w16251_,
		_w16497_
	);
	LUT2 #(
		.INIT('h1)
	) name5986 (
		_w16252_,
		_w16253_,
		_w16498_
	);
	LUT2 #(
		.INIT('h1)
	) name5987 (
		_w16254_,
		_w16255_,
		_w16499_
	);
	LUT2 #(
		.INIT('h1)
	) name5988 (
		_w16256_,
		_w16257_,
		_w16500_
	);
	LUT2 #(
		.INIT('h1)
	) name5989 (
		_w16258_,
		_w16259_,
		_w16501_
	);
	LUT2 #(
		.INIT('h1)
	) name5990 (
		_w16260_,
		_w16261_,
		_w16502_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w16262_,
		_w16263_,
		_w16503_
	);
	LUT2 #(
		.INIT('h1)
	) name5992 (
		_w16264_,
		_w16265_,
		_w16504_
	);
	LUT2 #(
		.INIT('h1)
	) name5993 (
		_w16266_,
		_w16267_,
		_w16505_
	);
	LUT2 #(
		.INIT('h1)
	) name5994 (
		_w16268_,
		_w16269_,
		_w16506_
	);
	LUT2 #(
		.INIT('h1)
	) name5995 (
		_w16270_,
		_w16271_,
		_w16507_
	);
	LUT2 #(
		.INIT('h1)
	) name5996 (
		_w16272_,
		_w16273_,
		_w16508_
	);
	LUT2 #(
		.INIT('h1)
	) name5997 (
		_w16274_,
		_w16275_,
		_w16509_
	);
	LUT2 #(
		.INIT('h1)
	) name5998 (
		_w16276_,
		_w16277_,
		_w16510_
	);
	LUT2 #(
		.INIT('h1)
	) name5999 (
		_w16278_,
		_w16279_,
		_w16511_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w16280_,
		_w16281_,
		_w16512_
	);
	LUT2 #(
		.INIT('h1)
	) name6001 (
		_w16282_,
		_w16283_,
		_w16513_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w16284_,
		_w16285_,
		_w16514_
	);
	LUT2 #(
		.INIT('h1)
	) name6003 (
		_w16286_,
		_w16287_,
		_w16515_
	);
	LUT2 #(
		.INIT('h1)
	) name6004 (
		_w16288_,
		_w16289_,
		_w16516_
	);
	LUT2 #(
		.INIT('h1)
	) name6005 (
		_w16290_,
		_w16291_,
		_w16517_
	);
	LUT2 #(
		.INIT('h1)
	) name6006 (
		_w16292_,
		_w16293_,
		_w16518_
	);
	LUT2 #(
		.INIT('h1)
	) name6007 (
		_w16294_,
		_w16295_,
		_w16519_
	);
	LUT2 #(
		.INIT('h1)
	) name6008 (
		_w16296_,
		_w16297_,
		_w16520_
	);
	LUT2 #(
		.INIT('h1)
	) name6009 (
		_w16298_,
		_w16299_,
		_w16521_
	);
	LUT2 #(
		.INIT('h1)
	) name6010 (
		_w16300_,
		_w16301_,
		_w16522_
	);
	LUT2 #(
		.INIT('h1)
	) name6011 (
		_w16302_,
		_w16303_,
		_w16523_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		_w16304_,
		_w16305_,
		_w16524_
	);
	LUT2 #(
		.INIT('h1)
	) name6013 (
		_w16306_,
		_w16307_,
		_w16525_
	);
	LUT2 #(
		.INIT('h1)
	) name6014 (
		_w16308_,
		_w16309_,
		_w16526_
	);
	LUT2 #(
		.INIT('h1)
	) name6015 (
		_w16310_,
		_w16311_,
		_w16527_
	);
	LUT2 #(
		.INIT('h1)
	) name6016 (
		_w16312_,
		_w16313_,
		_w16528_
	);
	LUT2 #(
		.INIT('h1)
	) name6017 (
		_w16314_,
		_w16315_,
		_w16529_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w16316_,
		_w16317_,
		_w16530_
	);
	LUT2 #(
		.INIT('h1)
	) name6019 (
		_w16318_,
		_w16319_,
		_w16531_
	);
	LUT2 #(
		.INIT('h1)
	) name6020 (
		_w16320_,
		_w16321_,
		_w16532_
	);
	LUT2 #(
		.INIT('h1)
	) name6021 (
		_w16322_,
		_w16323_,
		_w16533_
	);
	LUT2 #(
		.INIT('h1)
	) name6022 (
		_w16324_,
		_w16325_,
		_w16534_
	);
	LUT2 #(
		.INIT('h1)
	) name6023 (
		_w16326_,
		_w16327_,
		_w16535_
	);
	LUT2 #(
		.INIT('h1)
	) name6024 (
		_w16328_,
		_w16329_,
		_w16536_
	);
	LUT2 #(
		.INIT('h1)
	) name6025 (
		_w16330_,
		_w16331_,
		_w16537_
	);
	LUT2 #(
		.INIT('h1)
	) name6026 (
		_w16332_,
		_w16333_,
		_w16538_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		_w16334_,
		_w16335_,
		_w16539_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w16336_,
		_w16337_,
		_w16540_
	);
	LUT2 #(
		.INIT('h1)
	) name6029 (
		_w16338_,
		_w16339_,
		_w16541_
	);
	LUT2 #(
		.INIT('h1)
	) name6030 (
		_w16340_,
		_w16341_,
		_w16542_
	);
	LUT2 #(
		.INIT('h1)
	) name6031 (
		_w16342_,
		_w16343_,
		_w16543_
	);
	LUT2 #(
		.INIT('h1)
	) name6032 (
		_w16344_,
		_w16345_,
		_w16544_
	);
	LUT2 #(
		.INIT('h1)
	) name6033 (
		_w16346_,
		_w16347_,
		_w16545_
	);
	LUT2 #(
		.INIT('h1)
	) name6034 (
		_w16348_,
		_w16349_,
		_w16546_
	);
	LUT2 #(
		.INIT('h1)
	) name6035 (
		_w16350_,
		_w16351_,
		_w16547_
	);
	LUT2 #(
		.INIT('h1)
	) name6036 (
		_w16352_,
		_w16353_,
		_w16548_
	);
	LUT2 #(
		.INIT('h1)
	) name6037 (
		_w16354_,
		_w16355_,
		_w16549_
	);
	LUT2 #(
		.INIT('h1)
	) name6038 (
		_w16356_,
		_w16357_,
		_w16550_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w16358_,
		_w16359_,
		_w16551_
	);
	LUT2 #(
		.INIT('h1)
	) name6040 (
		_w16360_,
		_w16361_,
		_w16552_
	);
	LUT2 #(
		.INIT('h1)
	) name6041 (
		_w16362_,
		_w16363_,
		_w16553_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w16364_,
		_w16365_,
		_w16554_
	);
	LUT2 #(
		.INIT('h1)
	) name6043 (
		_w16366_,
		_w16367_,
		_w16555_
	);
	LUT2 #(
		.INIT('h1)
	) name6044 (
		_w16368_,
		_w16369_,
		_w16556_
	);
	LUT2 #(
		.INIT('h1)
	) name6045 (
		_w16370_,
		_w16371_,
		_w16557_
	);
	LUT2 #(
		.INIT('h1)
	) name6046 (
		_w16372_,
		_w16373_,
		_w16558_
	);
	LUT2 #(
		.INIT('h1)
	) name6047 (
		_w16374_,
		_w16375_,
		_w16559_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		_w16376_,
		_w16377_,
		_w16560_
	);
	LUT2 #(
		.INIT('h1)
	) name6049 (
		_w16378_,
		_w16379_,
		_w16561_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w16380_,
		_w16381_,
		_w16562_
	);
	LUT2 #(
		.INIT('h1)
	) name6051 (
		_w16382_,
		_w16383_,
		_w16563_
	);
	LUT2 #(
		.INIT('h1)
	) name6052 (
		_w16384_,
		_w16385_,
		_w16564_
	);
	LUT2 #(
		.INIT('h1)
	) name6053 (
		_w16386_,
		_w16387_,
		_w16565_
	);
	LUT2 #(
		.INIT('h1)
	) name6054 (
		_w16388_,
		_w16389_,
		_w16566_
	);
	LUT2 #(
		.INIT('h1)
	) name6055 (
		_w16390_,
		_w16391_,
		_w16567_
	);
	LUT2 #(
		.INIT('h1)
	) name6056 (
		_w16392_,
		_w16393_,
		_w16568_
	);
	LUT2 #(
		.INIT('h1)
	) name6057 (
		_w16394_,
		_w16395_,
		_w16569_
	);
	LUT2 #(
		.INIT('h1)
	) name6058 (
		_w16396_,
		_w16397_,
		_w16570_
	);
	LUT2 #(
		.INIT('h1)
	) name6059 (
		_w16398_,
		_w16399_,
		_w16571_
	);
	LUT2 #(
		.INIT('h1)
	) name6060 (
		_w16400_,
		_w16401_,
		_w16572_
	);
	LUT2 #(
		.INIT('h1)
	) name6061 (
		_w16402_,
		_w16403_,
		_w16573_
	);
	LUT2 #(
		.INIT('h1)
	) name6062 (
		_w16404_,
		_w16405_,
		_w16574_
	);
	LUT2 #(
		.INIT('h1)
	) name6063 (
		_w16406_,
		_w16407_,
		_w16575_
	);
	LUT2 #(
		.INIT('h1)
	) name6064 (
		_w16408_,
		_w16409_,
		_w16576_
	);
	LUT2 #(
		.INIT('h1)
	) name6065 (
		_w16410_,
		_w16411_,
		_w16577_
	);
	LUT2 #(
		.INIT('h1)
	) name6066 (
		_w16412_,
		_w16413_,
		_w16578_
	);
	LUT2 #(
		.INIT('h1)
	) name6067 (
		_w16414_,
		_w16415_,
		_w16579_
	);
	LUT2 #(
		.INIT('h1)
	) name6068 (
		_w16416_,
		_w16417_,
		_w16580_
	);
	LUT2 #(
		.INIT('h1)
	) name6069 (
		_w16418_,
		_w16419_,
		_w16581_
	);
	LUT2 #(
		.INIT('h1)
	) name6070 (
		_w16420_,
		_w16421_,
		_w16582_
	);
	LUT2 #(
		.INIT('h1)
	) name6071 (
		_w16422_,
		_w16423_,
		_w16583_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w16424_,
		_w16425_,
		_w16584_
	);
	LUT2 #(
		.INIT('h1)
	) name6073 (
		_w16426_,
		_w16427_,
		_w16585_
	);
	LUT2 #(
		.INIT('h1)
	) name6074 (
		_w16428_,
		_w16429_,
		_w16586_
	);
	LUT2 #(
		.INIT('h1)
	) name6075 (
		_w16430_,
		_w16431_,
		_w16587_
	);
	LUT2 #(
		.INIT('h1)
	) name6076 (
		_w16432_,
		_w16433_,
		_w16588_
	);
	LUT2 #(
		.INIT('h1)
	) name6077 (
		_w16434_,
		_w16435_,
		_w16589_
	);
	LUT2 #(
		.INIT('h1)
	) name6078 (
		_w16436_,
		_w16437_,
		_w16590_
	);
	LUT2 #(
		.INIT('h1)
	) name6079 (
		_w16438_,
		_w16439_,
		_w16591_
	);
	LUT2 #(
		.INIT('h1)
	) name6080 (
		_w16440_,
		_w16441_,
		_w16592_
	);
	LUT2 #(
		.INIT('h1)
	) name6081 (
		_w16442_,
		_w16443_,
		_w16593_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		_w16444_,
		_w16445_,
		_w16594_
	);
	LUT2 #(
		.INIT('h1)
	) name6083 (
		_w16446_,
		_w16447_,
		_w16595_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		_w16448_,
		_w16449_,
		_w16596_
	);
	LUT2 #(
		.INIT('h1)
	) name6085 (
		_w16450_,
		_w16451_,
		_w16597_
	);
	LUT2 #(
		.INIT('h1)
	) name6086 (
		_w16452_,
		_w16453_,
		_w16598_
	);
	LUT2 #(
		.INIT('h1)
	) name6087 (
		_w16454_,
		_w16455_,
		_w16599_
	);
	LUT2 #(
		.INIT('h1)
	) name6088 (
		_w16456_,
		_w16457_,
		_w16600_
	);
	LUT2 #(
		.INIT('h1)
	) name6089 (
		_w16458_,
		_w16459_,
		_w16601_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		_w16460_,
		_w16461_,
		_w16602_
	);
	LUT2 #(
		.INIT('h1)
	) name6091 (
		_w16462_,
		_w16463_,
		_w16603_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w16464_,
		_w16465_,
		_w16604_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		_w16466_,
		_w16467_,
		_w16605_
	);
	LUT2 #(
		.INIT('h1)
	) name6094 (
		_w16468_,
		_w16469_,
		_w16606_
	);
	LUT2 #(
		.INIT('h1)
	) name6095 (
		_w16470_,
		_w16471_,
		_w16607_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		_w16472_,
		_w16473_,
		_w16608_
	);
	LUT2 #(
		.INIT('h1)
	) name6097 (
		_w16474_,
		_w16475_,
		_w16609_
	);
	LUT2 #(
		.INIT('h1)
	) name6098 (
		_w16476_,
		_w16477_,
		_w16610_
	);
	LUT2 #(
		.INIT('h1)
	) name6099 (
		_w16478_,
		_w16479_,
		_w16611_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		_w16480_,
		_w16481_,
		_w16612_
	);
	LUT2 #(
		.INIT('h1)
	) name6101 (
		_w16482_,
		_w16483_,
		_w16613_
	);
	LUT2 #(
		.INIT('h1)
	) name6102 (
		_w16484_,
		_w16485_,
		_w16614_
	);
	LUT2 #(
		.INIT('h1)
	) name6103 (
		_w16486_,
		_w16487_,
		_w16615_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		_w16614_,
		_w16615_,
		_w16616_
	);
	LUT2 #(
		.INIT('h8)
	) name6105 (
		_w16612_,
		_w16613_,
		_w16617_
	);
	LUT2 #(
		.INIT('h8)
	) name6106 (
		_w16610_,
		_w16611_,
		_w16618_
	);
	LUT2 #(
		.INIT('h8)
	) name6107 (
		_w16608_,
		_w16609_,
		_w16619_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		_w16606_,
		_w16607_,
		_w16620_
	);
	LUT2 #(
		.INIT('h8)
	) name6109 (
		_w16604_,
		_w16605_,
		_w16621_
	);
	LUT2 #(
		.INIT('h8)
	) name6110 (
		_w16602_,
		_w16603_,
		_w16622_
	);
	LUT2 #(
		.INIT('h8)
	) name6111 (
		_w16600_,
		_w16601_,
		_w16623_
	);
	LUT2 #(
		.INIT('h8)
	) name6112 (
		_w16598_,
		_w16599_,
		_w16624_
	);
	LUT2 #(
		.INIT('h8)
	) name6113 (
		_w16596_,
		_w16597_,
		_w16625_
	);
	LUT2 #(
		.INIT('h8)
	) name6114 (
		_w16594_,
		_w16595_,
		_w16626_
	);
	LUT2 #(
		.INIT('h8)
	) name6115 (
		_w16592_,
		_w16593_,
		_w16627_
	);
	LUT2 #(
		.INIT('h8)
	) name6116 (
		_w16590_,
		_w16591_,
		_w16628_
	);
	LUT2 #(
		.INIT('h8)
	) name6117 (
		_w16588_,
		_w16589_,
		_w16629_
	);
	LUT2 #(
		.INIT('h8)
	) name6118 (
		_w16586_,
		_w16587_,
		_w16630_
	);
	LUT2 #(
		.INIT('h8)
	) name6119 (
		_w16584_,
		_w16585_,
		_w16631_
	);
	LUT2 #(
		.INIT('h8)
	) name6120 (
		_w16582_,
		_w16583_,
		_w16632_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		_w16580_,
		_w16581_,
		_w16633_
	);
	LUT2 #(
		.INIT('h8)
	) name6122 (
		_w16578_,
		_w16579_,
		_w16634_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		_w16576_,
		_w16577_,
		_w16635_
	);
	LUT2 #(
		.INIT('h8)
	) name6124 (
		_w16574_,
		_w16575_,
		_w16636_
	);
	LUT2 #(
		.INIT('h8)
	) name6125 (
		_w16572_,
		_w16573_,
		_w16637_
	);
	LUT2 #(
		.INIT('h8)
	) name6126 (
		_w16570_,
		_w16571_,
		_w16638_
	);
	LUT2 #(
		.INIT('h8)
	) name6127 (
		_w16568_,
		_w16569_,
		_w16639_
	);
	LUT2 #(
		.INIT('h8)
	) name6128 (
		_w16566_,
		_w16567_,
		_w16640_
	);
	LUT2 #(
		.INIT('h8)
	) name6129 (
		_w16564_,
		_w16565_,
		_w16641_
	);
	LUT2 #(
		.INIT('h8)
	) name6130 (
		_w16562_,
		_w16563_,
		_w16642_
	);
	LUT2 #(
		.INIT('h8)
	) name6131 (
		_w16560_,
		_w16561_,
		_w16643_
	);
	LUT2 #(
		.INIT('h8)
	) name6132 (
		_w16558_,
		_w16559_,
		_w16644_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		_w16556_,
		_w16557_,
		_w16645_
	);
	LUT2 #(
		.INIT('h8)
	) name6134 (
		_w16554_,
		_w16555_,
		_w16646_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		_w16552_,
		_w16553_,
		_w16647_
	);
	LUT2 #(
		.INIT('h8)
	) name6136 (
		_w16550_,
		_w16551_,
		_w16648_
	);
	LUT2 #(
		.INIT('h8)
	) name6137 (
		_w16548_,
		_w16549_,
		_w16649_
	);
	LUT2 #(
		.INIT('h8)
	) name6138 (
		_w16546_,
		_w16547_,
		_w16650_
	);
	LUT2 #(
		.INIT('h8)
	) name6139 (
		_w16544_,
		_w16545_,
		_w16651_
	);
	LUT2 #(
		.INIT('h8)
	) name6140 (
		_w16542_,
		_w16543_,
		_w16652_
	);
	LUT2 #(
		.INIT('h8)
	) name6141 (
		_w16540_,
		_w16541_,
		_w16653_
	);
	LUT2 #(
		.INIT('h8)
	) name6142 (
		_w16538_,
		_w16539_,
		_w16654_
	);
	LUT2 #(
		.INIT('h8)
	) name6143 (
		_w16536_,
		_w16537_,
		_w16655_
	);
	LUT2 #(
		.INIT('h8)
	) name6144 (
		_w16534_,
		_w16535_,
		_w16656_
	);
	LUT2 #(
		.INIT('h8)
	) name6145 (
		_w16532_,
		_w16533_,
		_w16657_
	);
	LUT2 #(
		.INIT('h8)
	) name6146 (
		_w16530_,
		_w16531_,
		_w16658_
	);
	LUT2 #(
		.INIT('h8)
	) name6147 (
		_w16528_,
		_w16529_,
		_w16659_
	);
	LUT2 #(
		.INIT('h8)
	) name6148 (
		_w16526_,
		_w16527_,
		_w16660_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		_w16524_,
		_w16525_,
		_w16661_
	);
	LUT2 #(
		.INIT('h8)
	) name6150 (
		_w16522_,
		_w16523_,
		_w16662_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		_w16520_,
		_w16521_,
		_w16663_
	);
	LUT2 #(
		.INIT('h8)
	) name6152 (
		_w16518_,
		_w16519_,
		_w16664_
	);
	LUT2 #(
		.INIT('h8)
	) name6153 (
		_w16516_,
		_w16517_,
		_w16665_
	);
	LUT2 #(
		.INIT('h8)
	) name6154 (
		_w16514_,
		_w16515_,
		_w16666_
	);
	LUT2 #(
		.INIT('h8)
	) name6155 (
		_w16512_,
		_w16513_,
		_w16667_
	);
	LUT2 #(
		.INIT('h8)
	) name6156 (
		_w16510_,
		_w16511_,
		_w16668_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		_w16508_,
		_w16509_,
		_w16669_
	);
	LUT2 #(
		.INIT('h8)
	) name6158 (
		_w16506_,
		_w16507_,
		_w16670_
	);
	LUT2 #(
		.INIT('h8)
	) name6159 (
		_w16504_,
		_w16505_,
		_w16671_
	);
	LUT2 #(
		.INIT('h8)
	) name6160 (
		_w16502_,
		_w16503_,
		_w16672_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		_w16500_,
		_w16501_,
		_w16673_
	);
	LUT2 #(
		.INIT('h8)
	) name6162 (
		_w16498_,
		_w16499_,
		_w16674_
	);
	LUT2 #(
		.INIT('h8)
	) name6163 (
		_w16496_,
		_w16497_,
		_w16675_
	);
	LUT2 #(
		.INIT('h8)
	) name6164 (
		_w16494_,
		_w16495_,
		_w16676_
	);
	LUT2 #(
		.INIT('h8)
	) name6165 (
		_w16492_,
		_w16493_,
		_w16677_
	);
	LUT2 #(
		.INIT('h8)
	) name6166 (
		_w16490_,
		_w16491_,
		_w16678_
	);
	LUT2 #(
		.INIT('h8)
	) name6167 (
		_w16488_,
		_w16489_,
		_w16679_
	);
	LUT2 #(
		.INIT('h8)
	) name6168 (
		_w16678_,
		_w16679_,
		_w16680_
	);
	LUT2 #(
		.INIT('h8)
	) name6169 (
		_w16676_,
		_w16677_,
		_w16681_
	);
	LUT2 #(
		.INIT('h8)
	) name6170 (
		_w16674_,
		_w16675_,
		_w16682_
	);
	LUT2 #(
		.INIT('h8)
	) name6171 (
		_w16672_,
		_w16673_,
		_w16683_
	);
	LUT2 #(
		.INIT('h8)
	) name6172 (
		_w16670_,
		_w16671_,
		_w16684_
	);
	LUT2 #(
		.INIT('h8)
	) name6173 (
		_w16668_,
		_w16669_,
		_w16685_
	);
	LUT2 #(
		.INIT('h8)
	) name6174 (
		_w16666_,
		_w16667_,
		_w16686_
	);
	LUT2 #(
		.INIT('h8)
	) name6175 (
		_w16664_,
		_w16665_,
		_w16687_
	);
	LUT2 #(
		.INIT('h8)
	) name6176 (
		_w16662_,
		_w16663_,
		_w16688_
	);
	LUT2 #(
		.INIT('h8)
	) name6177 (
		_w16660_,
		_w16661_,
		_w16689_
	);
	LUT2 #(
		.INIT('h8)
	) name6178 (
		_w16658_,
		_w16659_,
		_w16690_
	);
	LUT2 #(
		.INIT('h8)
	) name6179 (
		_w16656_,
		_w16657_,
		_w16691_
	);
	LUT2 #(
		.INIT('h8)
	) name6180 (
		_w16654_,
		_w16655_,
		_w16692_
	);
	LUT2 #(
		.INIT('h8)
	) name6181 (
		_w16652_,
		_w16653_,
		_w16693_
	);
	LUT2 #(
		.INIT('h8)
	) name6182 (
		_w16650_,
		_w16651_,
		_w16694_
	);
	LUT2 #(
		.INIT('h8)
	) name6183 (
		_w16648_,
		_w16649_,
		_w16695_
	);
	LUT2 #(
		.INIT('h8)
	) name6184 (
		_w16646_,
		_w16647_,
		_w16696_
	);
	LUT2 #(
		.INIT('h8)
	) name6185 (
		_w16644_,
		_w16645_,
		_w16697_
	);
	LUT2 #(
		.INIT('h8)
	) name6186 (
		_w16642_,
		_w16643_,
		_w16698_
	);
	LUT2 #(
		.INIT('h8)
	) name6187 (
		_w16640_,
		_w16641_,
		_w16699_
	);
	LUT2 #(
		.INIT('h8)
	) name6188 (
		_w16638_,
		_w16639_,
		_w16700_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		_w16636_,
		_w16637_,
		_w16701_
	);
	LUT2 #(
		.INIT('h8)
	) name6190 (
		_w16634_,
		_w16635_,
		_w16702_
	);
	LUT2 #(
		.INIT('h8)
	) name6191 (
		_w16632_,
		_w16633_,
		_w16703_
	);
	LUT2 #(
		.INIT('h8)
	) name6192 (
		_w16630_,
		_w16631_,
		_w16704_
	);
	LUT2 #(
		.INIT('h8)
	) name6193 (
		_w16628_,
		_w16629_,
		_w16705_
	);
	LUT2 #(
		.INIT('h8)
	) name6194 (
		_w16626_,
		_w16627_,
		_w16706_
	);
	LUT2 #(
		.INIT('h8)
	) name6195 (
		_w16624_,
		_w16625_,
		_w16707_
	);
	LUT2 #(
		.INIT('h8)
	) name6196 (
		_w16622_,
		_w16623_,
		_w16708_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		_w16620_,
		_w16621_,
		_w16709_
	);
	LUT2 #(
		.INIT('h8)
	) name6198 (
		_w16618_,
		_w16619_,
		_w16710_
	);
	LUT2 #(
		.INIT('h8)
	) name6199 (
		_w16616_,
		_w16617_,
		_w16711_
	);
	LUT2 #(
		.INIT('h8)
	) name6200 (
		_w16710_,
		_w16711_,
		_w16712_
	);
	LUT2 #(
		.INIT('h8)
	) name6201 (
		_w16708_,
		_w16709_,
		_w16713_
	);
	LUT2 #(
		.INIT('h8)
	) name6202 (
		_w16706_,
		_w16707_,
		_w16714_
	);
	LUT2 #(
		.INIT('h8)
	) name6203 (
		_w16704_,
		_w16705_,
		_w16715_
	);
	LUT2 #(
		.INIT('h8)
	) name6204 (
		_w16702_,
		_w16703_,
		_w16716_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		_w16700_,
		_w16701_,
		_w16717_
	);
	LUT2 #(
		.INIT('h8)
	) name6206 (
		_w16698_,
		_w16699_,
		_w16718_
	);
	LUT2 #(
		.INIT('h8)
	) name6207 (
		_w16696_,
		_w16697_,
		_w16719_
	);
	LUT2 #(
		.INIT('h8)
	) name6208 (
		_w16694_,
		_w16695_,
		_w16720_
	);
	LUT2 #(
		.INIT('h8)
	) name6209 (
		_w16692_,
		_w16693_,
		_w16721_
	);
	LUT2 #(
		.INIT('h8)
	) name6210 (
		_w16690_,
		_w16691_,
		_w16722_
	);
	LUT2 #(
		.INIT('h8)
	) name6211 (
		_w16688_,
		_w16689_,
		_w16723_
	);
	LUT2 #(
		.INIT('h8)
	) name6212 (
		_w16686_,
		_w16687_,
		_w16724_
	);
	LUT2 #(
		.INIT('h8)
	) name6213 (
		_w16684_,
		_w16685_,
		_w16725_
	);
	LUT2 #(
		.INIT('h8)
	) name6214 (
		_w16682_,
		_w16683_,
		_w16726_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		_w16680_,
		_w16681_,
		_w16727_
	);
	LUT2 #(
		.INIT('h8)
	) name6216 (
		_w16726_,
		_w16727_,
		_w16728_
	);
	LUT2 #(
		.INIT('h8)
	) name6217 (
		_w16724_,
		_w16725_,
		_w16729_
	);
	LUT2 #(
		.INIT('h8)
	) name6218 (
		_w16722_,
		_w16723_,
		_w16730_
	);
	LUT2 #(
		.INIT('h8)
	) name6219 (
		_w16720_,
		_w16721_,
		_w16731_
	);
	LUT2 #(
		.INIT('h8)
	) name6220 (
		_w16718_,
		_w16719_,
		_w16732_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		_w16716_,
		_w16717_,
		_w16733_
	);
	LUT2 #(
		.INIT('h8)
	) name6222 (
		_w16714_,
		_w16715_,
		_w16734_
	);
	LUT2 #(
		.INIT('h8)
	) name6223 (
		_w16712_,
		_w16713_,
		_w16735_
	);
	LUT2 #(
		.INIT('h8)
	) name6224 (
		_w16734_,
		_w16735_,
		_w16736_
	);
	LUT2 #(
		.INIT('h8)
	) name6225 (
		_w16732_,
		_w16733_,
		_w16737_
	);
	LUT2 #(
		.INIT('h8)
	) name6226 (
		_w16730_,
		_w16731_,
		_w16738_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		_w16728_,
		_w16729_,
		_w16739_
	);
	LUT2 #(
		.INIT('h8)
	) name6228 (
		_w16738_,
		_w16739_,
		_w16740_
	);
	LUT2 #(
		.INIT('h8)
	) name6229 (
		_w16736_,
		_w16737_,
		_w16741_
	);
	LUT2 #(
		.INIT('h8)
	) name6230 (
		_w16740_,
		_w16741_,
		_w16742_
	);
	LUT2 #(
		.INIT('h1)
	) name6231 (
		wb_rst_i_pad,
		_w16742_,
		_w16743_
	);
	LUT2 #(
		.INIT('h8)
	) name6232 (
		_w12656_,
		_w16743_,
		_w16744_
	);
	LUT2 #(
		.INIT('h2)
	) name6233 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w12657_,
		_w16745_
	);
	LUT2 #(
		.INIT('h2)
	) name6234 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w13480_,
		_w16746_
	);
	LUT2 #(
		.INIT('h1)
	) name6235 (
		_w13481_,
		_w16746_,
		_w16747_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w16748_
	);
	LUT2 #(
		.INIT('h4)
	) name6237 (
		_w16747_,
		_w16748_,
		_w16749_
	);
	LUT2 #(
		.INIT('h4)
	) name6238 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w16750_
	);
	LUT2 #(
		.INIT('h4)
	) name6239 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w13480_,
		_w16751_
	);
	LUT2 #(
		.INIT('h2)
	) name6240 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w16751_,
		_w16752_
	);
	LUT2 #(
		.INIT('h4)
	) name6241 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w13481_,
		_w16753_
	);
	LUT2 #(
		.INIT('h1)
	) name6242 (
		_w16752_,
		_w16753_,
		_w16754_
	);
	LUT2 #(
		.INIT('h2)
	) name6243 (
		_w16750_,
		_w16754_,
		_w16755_
	);
	LUT2 #(
		.INIT('h2)
	) name6244 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w16756_
	);
	LUT2 #(
		.INIT('h8)
	) name6245 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w16757_
	);
	LUT2 #(
		.INIT('h2)
	) name6246 (
		_w16747_,
		_w16757_,
		_w16758_
	);
	LUT2 #(
		.INIT('h4)
	) name6247 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w16757_,
		_w16759_
	);
	LUT2 #(
		.INIT('h2)
	) name6248 (
		_w16756_,
		_w16759_,
		_w16760_
	);
	LUT2 #(
		.INIT('h4)
	) name6249 (
		_w16758_,
		_w16760_,
		_w16761_
	);
	LUT2 #(
		.INIT('h8)
	) name6250 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w16762_
	);
	LUT2 #(
		.INIT('h1)
	) name6251 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w16763_
	);
	LUT2 #(
		.INIT('h8)
	) name6252 (
		_w13480_,
		_w16763_,
		_w16764_
	);
	LUT2 #(
		.INIT('h2)
	) name6253 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w16764_,
		_w16765_
	);
	LUT2 #(
		.INIT('h8)
	) name6254 (
		_w13481_,
		_w16763_,
		_w16766_
	);
	LUT2 #(
		.INIT('h1)
	) name6255 (
		_w16765_,
		_w16766_,
		_w16767_
	);
	LUT2 #(
		.INIT('h2)
	) name6256 (
		_w16762_,
		_w16767_,
		_w16768_
	);
	LUT2 #(
		.INIT('h1)
	) name6257 (
		_w16749_,
		_w16755_,
		_w16769_
	);
	LUT2 #(
		.INIT('h1)
	) name6258 (
		_w16761_,
		_w16768_,
		_w16770_
	);
	LUT2 #(
		.INIT('h8)
	) name6259 (
		_w16769_,
		_w16770_,
		_w16771_
	);
	LUT2 #(
		.INIT('h2)
	) name6260 (
		_w13500_,
		_w16771_,
		_w16772_
	);
	LUT2 #(
		.INIT('h1)
	) name6261 (
		_w16745_,
		_w16772_,
		_w16773_
	);
	LUT2 #(
		.INIT('h1)
	) name6262 (
		_w12656_,
		_w16773_,
		_w16774_
	);
	LUT2 #(
		.INIT('h1)
	) name6263 (
		_w16744_,
		_w16774_,
		_w16775_
	);
	LUT2 #(
		.INIT('h8)
	) name6264 (
		\wishbone_bd_ram_mem3_reg[89][26]/P0001 ,
		_w12964_,
		_w16776_
	);
	LUT2 #(
		.INIT('h8)
	) name6265 (
		\wishbone_bd_ram_mem3_reg[77][26]/P0001 ,
		_w12982_,
		_w16777_
	);
	LUT2 #(
		.INIT('h8)
	) name6266 (
		\wishbone_bd_ram_mem3_reg[166][26]/P0001 ,
		_w13040_,
		_w16778_
	);
	LUT2 #(
		.INIT('h8)
	) name6267 (
		\wishbone_bd_ram_mem3_reg[107][26]/P0001 ,
		_w12749_,
		_w16779_
	);
	LUT2 #(
		.INIT('h8)
	) name6268 (
		\wishbone_bd_ram_mem3_reg[47][26]/P0001 ,
		_w12904_,
		_w16780_
	);
	LUT2 #(
		.INIT('h8)
	) name6269 (
		\wishbone_bd_ram_mem3_reg[113][26]/P0001 ,
		_w13026_,
		_w16781_
	);
	LUT2 #(
		.INIT('h8)
	) name6270 (
		\wishbone_bd_ram_mem3_reg[131][26]/P0001 ,
		_w12852_,
		_w16782_
	);
	LUT2 #(
		.INIT('h8)
	) name6271 (
		\wishbone_bd_ram_mem3_reg[19][26]/P0001 ,
		_w13012_,
		_w16783_
	);
	LUT2 #(
		.INIT('h8)
	) name6272 (
		\wishbone_bd_ram_mem3_reg[102][26]/P0001 ,
		_w12685_,
		_w16784_
	);
	LUT2 #(
		.INIT('h8)
	) name6273 (
		\wishbone_bd_ram_mem3_reg[233][26]/P0001 ,
		_w12836_,
		_w16785_
	);
	LUT2 #(
		.INIT('h8)
	) name6274 (
		\wishbone_bd_ram_mem3_reg[255][26]/P0001 ,
		_w13072_,
		_w16786_
	);
	LUT2 #(
		.INIT('h8)
	) name6275 (
		\wishbone_bd_ram_mem3_reg[155][26]/P0001 ,
		_w13122_,
		_w16787_
	);
	LUT2 #(
		.INIT('h8)
	) name6276 (
		\wishbone_bd_ram_mem3_reg[43][26]/P0001 ,
		_w13200_,
		_w16788_
	);
	LUT2 #(
		.INIT('h8)
	) name6277 (
		\wishbone_bd_ram_mem3_reg[132][26]/P0001 ,
		_w12992_,
		_w16789_
	);
	LUT2 #(
		.INIT('h8)
	) name6278 (
		\wishbone_bd_ram_mem3_reg[62][26]/P0001 ,
		_w12673_,
		_w16790_
	);
	LUT2 #(
		.INIT('h8)
	) name6279 (
		\wishbone_bd_ram_mem3_reg[48][26]/P0001 ,
		_w12970_,
		_w16791_
	);
	LUT2 #(
		.INIT('h8)
	) name6280 (
		\wishbone_bd_ram_mem3_reg[231][26]/P0001 ,
		_w12856_,
		_w16792_
	);
	LUT2 #(
		.INIT('h8)
	) name6281 (
		\wishbone_bd_ram_mem3_reg[176][26]/P0001 ,
		_w12868_,
		_w16793_
	);
	LUT2 #(
		.INIT('h8)
	) name6282 (
		\wishbone_bd_ram_mem3_reg[50][26]/P0001 ,
		_w13150_,
		_w16794_
	);
	LUT2 #(
		.INIT('h8)
	) name6283 (
		\wishbone_bd_ram_mem3_reg[153][26]/P0001 ,
		_w12890_,
		_w16795_
	);
	LUT2 #(
		.INIT('h8)
	) name6284 (
		\wishbone_bd_ram_mem3_reg[16][26]/P0001 ,
		_w13140_,
		_w16796_
	);
	LUT2 #(
		.INIT('h8)
	) name6285 (
		\wishbone_bd_ram_mem3_reg[81][26]/P0001 ,
		_w12950_,
		_w16797_
	);
	LUT2 #(
		.INIT('h8)
	) name6286 (
		\wishbone_bd_ram_mem3_reg[140][26]/P0001 ,
		_w12894_,
		_w16798_
	);
	LUT2 #(
		.INIT('h8)
	) name6287 (
		\wishbone_bd_ram_mem3_reg[98][26]/P0001 ,
		_w12816_,
		_w16799_
	);
	LUT2 #(
		.INIT('h8)
	) name6288 (
		\wishbone_bd_ram_mem3_reg[133][26]/P0001 ,
		_w12761_,
		_w16800_
	);
	LUT2 #(
		.INIT('h8)
	) name6289 (
		\wishbone_bd_ram_mem3_reg[1][26]/P0001 ,
		_w13014_,
		_w16801_
	);
	LUT2 #(
		.INIT('h8)
	) name6290 (
		\wishbone_bd_ram_mem3_reg[223][26]/P0001 ,
		_w12838_,
		_w16802_
	);
	LUT2 #(
		.INIT('h8)
	) name6291 (
		\wishbone_bd_ram_mem3_reg[137][26]/P0001 ,
		_w13168_,
		_w16803_
	);
	LUT2 #(
		.INIT('h8)
	) name6292 (
		\wishbone_bd_ram_mem3_reg[105][26]/P0001 ,
		_w12751_,
		_w16804_
	);
	LUT2 #(
		.INIT('h8)
	) name6293 (
		\wishbone_bd_ram_mem3_reg[92][26]/P0001 ,
		_w13010_,
		_w16805_
	);
	LUT2 #(
		.INIT('h8)
	) name6294 (
		\wishbone_bd_ram_mem3_reg[193][26]/P0001 ,
		_w13056_,
		_w16806_
	);
	LUT2 #(
		.INIT('h8)
	) name6295 (
		\wishbone_bd_ram_mem3_reg[203][26]/P0001 ,
		_w13158_,
		_w16807_
	);
	LUT2 #(
		.INIT('h8)
	) name6296 (
		\wishbone_bd_ram_mem3_reg[136][26]/P0001 ,
		_w13064_,
		_w16808_
	);
	LUT2 #(
		.INIT('h8)
	) name6297 (
		\wishbone_bd_ram_mem3_reg[216][26]/P0001 ,
		_w13028_,
		_w16809_
	);
	LUT2 #(
		.INIT('h8)
	) name6298 (
		\wishbone_bd_ram_mem3_reg[97][26]/P0001 ,
		_w13096_,
		_w16810_
	);
	LUT2 #(
		.INIT('h8)
	) name6299 (
		\wishbone_bd_ram_mem3_reg[53][26]/P0001 ,
		_w13020_,
		_w16811_
	);
	LUT2 #(
		.INIT('h8)
	) name6300 (
		\wishbone_bd_ram_mem3_reg[60][26]/P0001 ,
		_w13204_,
		_w16812_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		\wishbone_bd_ram_mem3_reg[100][26]/P0001 ,
		_w12960_,
		_w16813_
	);
	LUT2 #(
		.INIT('h8)
	) name6302 (
		\wishbone_bd_ram_mem3_reg[83][26]/P0001 ,
		_w12916_,
		_w16814_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		\wishbone_bd_ram_mem3_reg[169][26]/P0001 ,
		_w12722_,
		_w16815_
	);
	LUT2 #(
		.INIT('h8)
	) name6304 (
		\wishbone_bd_ram_mem3_reg[114][26]/P0001 ,
		_w13202_,
		_w16816_
	);
	LUT2 #(
		.INIT('h8)
	) name6305 (
		\wishbone_bd_ram_mem3_reg[251][26]/P0001 ,
		_w13054_,
		_w16817_
	);
	LUT2 #(
		.INIT('h8)
	) name6306 (
		\wishbone_bd_ram_mem3_reg[3][26]/P0001 ,
		_w12866_,
		_w16818_
	);
	LUT2 #(
		.INIT('h8)
	) name6307 (
		\wishbone_bd_ram_mem3_reg[49][26]/P0001 ,
		_w12994_,
		_w16819_
	);
	LUT2 #(
		.INIT('h8)
	) name6308 (
		\wishbone_bd_ram_mem3_reg[220][26]/P0001 ,
		_w13066_,
		_w16820_
	);
	LUT2 #(
		.INIT('h8)
	) name6309 (
		\wishbone_bd_ram_mem3_reg[82][26]/P0001 ,
		_w12942_,
		_w16821_
	);
	LUT2 #(
		.INIT('h8)
	) name6310 (
		\wishbone_bd_ram_mem3_reg[196][26]/P0001 ,
		_w13090_,
		_w16822_
	);
	LUT2 #(
		.INIT('h8)
	) name6311 (
		\wishbone_bd_ram_mem3_reg[226][26]/P0001 ,
		_w13138_,
		_w16823_
	);
	LUT2 #(
		.INIT('h8)
	) name6312 (
		\wishbone_bd_ram_mem3_reg[192][26]/P0001 ,
		_w12938_,
		_w16824_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		\wishbone_bd_ram_mem3_reg[225][26]/P0001 ,
		_w13092_,
		_w16825_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		\wishbone_bd_ram_mem3_reg[88][26]/P0001 ,
		_w12860_,
		_w16826_
	);
	LUT2 #(
		.INIT('h8)
	) name6315 (
		\wishbone_bd_ram_mem3_reg[148][26]/P0001 ,
		_w13000_,
		_w16827_
	);
	LUT2 #(
		.INIT('h8)
	) name6316 (
		\wishbone_bd_ram_mem3_reg[250][26]/P0001 ,
		_w13128_,
		_w16828_
	);
	LUT2 #(
		.INIT('h8)
	) name6317 (
		\wishbone_bd_ram_mem3_reg[124][26]/P0001 ,
		_w13058_,
		_w16829_
	);
	LUT2 #(
		.INIT('h8)
	) name6318 (
		\wishbone_bd_ram_mem3_reg[78][26]/P0001 ,
		_w12874_,
		_w16830_
	);
	LUT2 #(
		.INIT('h8)
	) name6319 (
		\wishbone_bd_ram_mem3_reg[191][26]/P0001 ,
		_w13034_,
		_w16831_
	);
	LUT2 #(
		.INIT('h8)
	) name6320 (
		\wishbone_bd_ram_mem3_reg[171][26]/P0001 ,
		_w12910_,
		_w16832_
	);
	LUT2 #(
		.INIT('h8)
	) name6321 (
		\wishbone_bd_ram_mem3_reg[214][26]/P0001 ,
		_w12984_,
		_w16833_
	);
	LUT2 #(
		.INIT('h8)
	) name6322 (
		\wishbone_bd_ram_mem3_reg[93][26]/P0001 ,
		_w13016_,
		_w16834_
	);
	LUT2 #(
		.INIT('h8)
	) name6323 (
		\wishbone_bd_ram_mem3_reg[152][26]/P0001 ,
		_w12966_,
		_w16835_
	);
	LUT2 #(
		.INIT('h8)
	) name6324 (
		\wishbone_bd_ram_mem3_reg[227][26]/P0001 ,
		_w12936_,
		_w16836_
	);
	LUT2 #(
		.INIT('h8)
	) name6325 (
		\wishbone_bd_ram_mem3_reg[180][26]/P0001 ,
		_w12791_,
		_w16837_
	);
	LUT2 #(
		.INIT('h8)
	) name6326 (
		\wishbone_bd_ram_mem3_reg[202][26]/P0001 ,
		_w12870_,
		_w16838_
	);
	LUT2 #(
		.INIT('h8)
	) name6327 (
		\wishbone_bd_ram_mem3_reg[200][26]/P0001 ,
		_w12988_,
		_w16839_
	);
	LUT2 #(
		.INIT('h8)
	) name6328 (
		\wishbone_bd_ram_mem3_reg[248][26]/P0001 ,
		_w12789_,
		_w16840_
	);
	LUT2 #(
		.INIT('h8)
	) name6329 (
		\wishbone_bd_ram_mem3_reg[209][26]/P0001 ,
		_w13152_,
		_w16841_
	);
	LUT2 #(
		.INIT('h8)
	) name6330 (
		\wishbone_bd_ram_mem3_reg[15][26]/P0001 ,
		_w13210_,
		_w16842_
	);
	LUT2 #(
		.INIT('h8)
	) name6331 (
		\wishbone_bd_ram_mem3_reg[247][26]/P0001 ,
		_w12818_,
		_w16843_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		\wishbone_bd_ram_mem3_reg[90][26]/P0001 ,
		_w12978_,
		_w16844_
	);
	LUT2 #(
		.INIT('h8)
	) name6333 (
		\wishbone_bd_ram_mem3_reg[143][26]/P0001 ,
		_w12922_,
		_w16845_
	);
	LUT2 #(
		.INIT('h8)
	) name6334 (
		\wishbone_bd_ram_mem3_reg[160][26]/P0001 ,
		_w12872_,
		_w16846_
	);
	LUT2 #(
		.INIT('h8)
	) name6335 (
		\wishbone_bd_ram_mem3_reg[75][26]/P0001 ,
		_w12826_,
		_w16847_
	);
	LUT2 #(
		.INIT('h8)
	) name6336 (
		\wishbone_bd_ram_mem3_reg[67][26]/P0001 ,
		_w13134_,
		_w16848_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		\wishbone_bd_ram_mem3_reg[242][26]/P0001 ,
		_w12932_,
		_w16849_
	);
	LUT2 #(
		.INIT('h8)
	) name6338 (
		\wishbone_bd_ram_mem3_reg[120][26]/P0001 ,
		_w12707_,
		_w16850_
	);
	LUT2 #(
		.INIT('h8)
	) name6339 (
		\wishbone_bd_ram_mem3_reg[178][26]/P0001 ,
		_w12886_,
		_w16851_
	);
	LUT2 #(
		.INIT('h8)
	) name6340 (
		\wishbone_bd_ram_mem3_reg[125][26]/P0001 ,
		_w12956_,
		_w16852_
	);
	LUT2 #(
		.INIT('h8)
	) name6341 (
		\wishbone_bd_ram_mem3_reg[217][26]/P0001 ,
		_w13188_,
		_w16853_
	);
	LUT2 #(
		.INIT('h8)
	) name6342 (
		\wishbone_bd_ram_mem3_reg[215][26]/P0001 ,
		_w12974_,
		_w16854_
	);
	LUT2 #(
		.INIT('h8)
	) name6343 (
		\wishbone_bd_ram_mem3_reg[65][26]/P0001 ,
		_w13176_,
		_w16855_
	);
	LUT2 #(
		.INIT('h8)
	) name6344 (
		\wishbone_bd_ram_mem3_reg[36][26]/P0001 ,
		_w12800_,
		_w16856_
	);
	LUT2 #(
		.INIT('h8)
	) name6345 (
		\wishbone_bd_ram_mem3_reg[159][26]/P0001 ,
		_w12774_,
		_w16857_
	);
	LUT2 #(
		.INIT('h8)
	) name6346 (
		\wishbone_bd_ram_mem3_reg[64][26]/P0001 ,
		_w12976_,
		_w16858_
	);
	LUT2 #(
		.INIT('h8)
	) name6347 (
		\wishbone_bd_ram_mem3_reg[204][26]/P0001 ,
		_w13162_,
		_w16859_
	);
	LUT2 #(
		.INIT('h8)
	) name6348 (
		\wishbone_bd_ram_mem3_reg[57][26]/P0001 ,
		_w13116_,
		_w16860_
	);
	LUT2 #(
		.INIT('h8)
	) name6349 (
		\wishbone_bd_ram_mem3_reg[185][26]/P0001 ,
		_w12940_,
		_w16861_
	);
	LUT2 #(
		.INIT('h8)
	) name6350 (
		\wishbone_bd_ram_mem3_reg[189][26]/P0001 ,
		_w13042_,
		_w16862_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		\wishbone_bd_ram_mem3_reg[55][26]/P0001 ,
		_w12785_,
		_w16863_
	);
	LUT2 #(
		.INIT('h8)
	) name6352 (
		\wishbone_bd_ram_mem3_reg[63][26]/P0001 ,
		_w12850_,
		_w16864_
	);
	LUT2 #(
		.INIT('h8)
	) name6353 (
		\wishbone_bd_ram_mem3_reg[207][26]/P0001 ,
		_w13180_,
		_w16865_
	);
	LUT2 #(
		.INIT('h8)
	) name6354 (
		\wishbone_bd_ram_mem3_reg[254][26]/P0001 ,
		_w12892_,
		_w16866_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		\wishbone_bd_ram_mem3_reg[119][26]/P0001 ,
		_w13048_,
		_w16867_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		\wishbone_bd_ram_mem3_reg[201][26]/P0001 ,
		_w12822_,
		_w16868_
	);
	LUT2 #(
		.INIT('h8)
	) name6357 (
		\wishbone_bd_ram_mem3_reg[127][26]/P0001 ,
		_w13164_,
		_w16869_
	);
	LUT2 #(
		.INIT('h8)
	) name6358 (
		\wishbone_bd_ram_mem3_reg[86][26]/P0001 ,
		_w12735_,
		_w16870_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		\wishbone_bd_ram_mem3_reg[111][26]/P0001 ,
		_w12744_,
		_w16871_
	);
	LUT2 #(
		.INIT('h8)
	) name6360 (
		\wishbone_bd_ram_mem3_reg[112][26]/P0001 ,
		_w12733_,
		_w16872_
	);
	LUT2 #(
		.INIT('h8)
	) name6361 (
		\wishbone_bd_ram_mem3_reg[108][26]/P0001 ,
		_w13156_,
		_w16873_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		\wishbone_bd_ram_mem3_reg[135][26]/P0001 ,
		_w13124_,
		_w16874_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		\wishbone_bd_ram_mem3_reg[12][26]/P0001 ,
		_w13118_,
		_w16875_
	);
	LUT2 #(
		.INIT('h8)
	) name6364 (
		\wishbone_bd_ram_mem3_reg[76][26]/P0001 ,
		_w13184_,
		_w16876_
	);
	LUT2 #(
		.INIT('h8)
	) name6365 (
		\wishbone_bd_ram_mem3_reg[157][26]/P0001 ,
		_w12926_,
		_w16877_
	);
	LUT2 #(
		.INIT('h8)
	) name6366 (
		\wishbone_bd_ram_mem3_reg[145][26]/P0001 ,
		_w13106_,
		_w16878_
	);
	LUT2 #(
		.INIT('h8)
	) name6367 (
		\wishbone_bd_ram_mem3_reg[104][26]/P0001 ,
		_w13148_,
		_w16879_
	);
	LUT2 #(
		.INIT('h8)
	) name6368 (
		\wishbone_bd_ram_mem3_reg[11][26]/P0001 ,
		_w13194_,
		_w16880_
	);
	LUT2 #(
		.INIT('h8)
	) name6369 (
		\wishbone_bd_ram_mem3_reg[41][26]/P0001 ,
		_w13052_,
		_w16881_
	);
	LUT2 #(
		.INIT('h8)
	) name6370 (
		\wishbone_bd_ram_mem3_reg[40][26]/P0001 ,
		_w13132_,
		_w16882_
	);
	LUT2 #(
		.INIT('h8)
	) name6371 (
		\wishbone_bd_ram_mem3_reg[151][26]/P0001 ,
		_w13142_,
		_w16883_
	);
	LUT2 #(
		.INIT('h8)
	) name6372 (
		\wishbone_bd_ram_mem3_reg[10][26]/P0001 ,
		_w13172_,
		_w16884_
	);
	LUT2 #(
		.INIT('h8)
	) name6373 (
		\wishbone_bd_ram_mem3_reg[29][26]/P0001 ,
		_w12952_,
		_w16885_
	);
	LUT2 #(
		.INIT('h8)
	) name6374 (
		\wishbone_bd_ram_mem3_reg[87][26]/P0001 ,
		_w13154_,
		_w16886_
	);
	LUT2 #(
		.INIT('h8)
	) name6375 (
		\wishbone_bd_ram_mem3_reg[141][26]/P0001 ,
		_w13004_,
		_w16887_
	);
	LUT2 #(
		.INIT('h8)
	) name6376 (
		\wishbone_bd_ram_mem3_reg[205][26]/P0001 ,
		_w13068_,
		_w16888_
	);
	LUT2 #(
		.INIT('h8)
	) name6377 (
		\wishbone_bd_ram_mem3_reg[26][26]/P0001 ,
		_w12699_,
		_w16889_
	);
	LUT2 #(
		.INIT('h8)
	) name6378 (
		\wishbone_bd_ram_mem3_reg[229][26]/P0001 ,
		_w12711_,
		_w16890_
	);
	LUT2 #(
		.INIT('h8)
	) name6379 (
		\wishbone_bd_ram_mem3_reg[146][26]/P0001 ,
		_w13060_,
		_w16891_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		\wishbone_bd_ram_mem3_reg[212][26]/P0001 ,
		_w12796_,
		_w16892_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		\wishbone_bd_ram_mem3_reg[54][26]/P0001 ,
		_w12770_,
		_w16893_
	);
	LUT2 #(
		.INIT('h8)
	) name6382 (
		\wishbone_bd_ram_mem3_reg[228][26]/P0001 ,
		_w12765_,
		_w16894_
	);
	LUT2 #(
		.INIT('h8)
	) name6383 (
		\wishbone_bd_ram_mem3_reg[18][26]/P0001 ,
		_w12679_,
		_w16895_
	);
	LUT2 #(
		.INIT('h8)
	) name6384 (
		\wishbone_bd_ram_mem3_reg[239][26]/P0001 ,
		_w12862_,
		_w16896_
	);
	LUT2 #(
		.INIT('h8)
	) name6385 (
		\wishbone_bd_ram_mem3_reg[206][26]/P0001 ,
		_w12954_,
		_w16897_
	);
	LUT2 #(
		.INIT('h8)
	) name6386 (
		\wishbone_bd_ram_mem3_reg[56][26]/P0001 ,
		_w12778_,
		_w16898_
	);
	LUT2 #(
		.INIT('h8)
	) name6387 (
		\wishbone_bd_ram_mem3_reg[253][26]/P0001 ,
		_w13100_,
		_w16899_
	);
	LUT2 #(
		.INIT('h8)
	) name6388 (
		\wishbone_bd_ram_mem3_reg[182][26]/P0001 ,
		_w12820_,
		_w16900_
	);
	LUT2 #(
		.INIT('h8)
	) name6389 (
		\wishbone_bd_ram_mem3_reg[188][26]/P0001 ,
		_w12948_,
		_w16901_
	);
	LUT2 #(
		.INIT('h8)
	) name6390 (
		\wishbone_bd_ram_mem3_reg[32][26]/P0001 ,
		_w13120_,
		_w16902_
	);
	LUT2 #(
		.INIT('h8)
	) name6391 (
		\wishbone_bd_ram_mem3_reg[138][26]/P0001 ,
		_w12958_,
		_w16903_
	);
	LUT2 #(
		.INIT('h8)
	) name6392 (
		\wishbone_bd_ram_mem3_reg[156][26]/P0001 ,
		_w13190_,
		_w16904_
	);
	LUT2 #(
		.INIT('h8)
	) name6393 (
		\wishbone_bd_ram_mem3_reg[208][26]/P0001 ,
		_w13032_,
		_w16905_
	);
	LUT2 #(
		.INIT('h8)
	) name6394 (
		\wishbone_bd_ram_mem3_reg[28][26]/P0001 ,
		_w13170_,
		_w16906_
	);
	LUT2 #(
		.INIT('h8)
	) name6395 (
		\wishbone_bd_ram_mem3_reg[7][26]/P0001 ,
		_w12728_,
		_w16907_
	);
	LUT2 #(
		.INIT('h8)
	) name6396 (
		\wishbone_bd_ram_mem3_reg[27][26]/P0001 ,
		_w12880_,
		_w16908_
	);
	LUT2 #(
		.INIT('h8)
	) name6397 (
		\wishbone_bd_ram_mem3_reg[147][26]/P0001 ,
		_w13146_,
		_w16909_
	);
	LUT2 #(
		.INIT('h8)
	) name6398 (
		\wishbone_bd_ram_mem3_reg[80][26]/P0001 ,
		_w12689_,
		_w16910_
	);
	LUT2 #(
		.INIT('h8)
	) name6399 (
		\wishbone_bd_ram_mem3_reg[103][26]/P0001 ,
		_w12846_,
		_w16911_
	);
	LUT2 #(
		.INIT('h8)
	) name6400 (
		\wishbone_bd_ram_mem3_reg[30][26]/P0001 ,
		_w13104_,
		_w16912_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		\wishbone_bd_ram_mem3_reg[20][26]/P0001 ,
		_w13174_,
		_w16913_
	);
	LUT2 #(
		.INIT('h8)
	) name6402 (
		\wishbone_bd_ram_mem3_reg[252][26]/P0001 ,
		_w13080_,
		_w16914_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		\wishbone_bd_ram_mem3_reg[71][26]/P0001 ,
		_w12798_,
		_w16915_
	);
	LUT2 #(
		.INIT('h8)
	) name6404 (
		\wishbone_bd_ram_mem3_reg[177][26]/P0001 ,
		_w12996_,
		_w16916_
	);
	LUT2 #(
		.INIT('h8)
	) name6405 (
		\wishbone_bd_ram_mem3_reg[139][26]/P0001 ,
		_w12814_,
		_w16917_
	);
	LUT2 #(
		.INIT('h8)
	) name6406 (
		\wishbone_bd_ram_mem3_reg[165][26]/P0001 ,
		_w13044_,
		_w16918_
	);
	LUT2 #(
		.INIT('h8)
	) name6407 (
		\wishbone_bd_ram_mem3_reg[128][26]/P0001 ,
		_w12793_,
		_w16919_
	);
	LUT2 #(
		.INIT('h8)
	) name6408 (
		\wishbone_bd_ram_mem3_reg[96][26]/P0001 ,
		_w12912_,
		_w16920_
	);
	LUT2 #(
		.INIT('h8)
	) name6409 (
		\wishbone_bd_ram_mem3_reg[59][26]/P0001 ,
		_w12780_,
		_w16921_
	);
	LUT2 #(
		.INIT('h8)
	) name6410 (
		\wishbone_bd_ram_mem3_reg[161][26]/P0001 ,
		_w12754_,
		_w16922_
	);
	LUT2 #(
		.INIT('h8)
	) name6411 (
		\wishbone_bd_ram_mem3_reg[221][26]/P0001 ,
		_w12802_,
		_w16923_
	);
	LUT2 #(
		.INIT('h8)
	) name6412 (
		\wishbone_bd_ram_mem3_reg[84][26]/P0001 ,
		_w12934_,
		_w16924_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		\wishbone_bd_ram_mem3_reg[186][26]/P0001 ,
		_w12783_,
		_w16925_
	);
	LUT2 #(
		.INIT('h8)
	) name6414 (
		\wishbone_bd_ram_mem3_reg[99][26]/P0001 ,
		_w13038_,
		_w16926_
	);
	LUT2 #(
		.INIT('h8)
	) name6415 (
		\wishbone_bd_ram_mem3_reg[123][26]/P0001 ,
		_w13114_,
		_w16927_
	);
	LUT2 #(
		.INIT('h8)
	) name6416 (
		\wishbone_bd_ram_mem3_reg[70][26]/P0001 ,
		_w12840_,
		_w16928_
	);
	LUT2 #(
		.INIT('h8)
	) name6417 (
		\wishbone_bd_ram_mem3_reg[9][26]/P0001 ,
		_w12808_,
		_w16929_
	);
	LUT2 #(
		.INIT('h8)
	) name6418 (
		\wishbone_bd_ram_mem3_reg[51][26]/P0001 ,
		_w13024_,
		_w16930_
	);
	LUT2 #(
		.INIT('h8)
	) name6419 (
		\wishbone_bd_ram_mem3_reg[72][26]/P0001 ,
		_w12810_,
		_w16931_
	);
	LUT2 #(
		.INIT('h8)
	) name6420 (
		\wishbone_bd_ram_mem3_reg[129][26]/P0001 ,
		_w12776_,
		_w16932_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		\wishbone_bd_ram_mem3_reg[237][26]/P0001 ,
		_w12990_,
		_w16933_
	);
	LUT2 #(
		.INIT('h8)
	) name6422 (
		\wishbone_bd_ram_mem3_reg[22][26]/P0001 ,
		_w13110_,
		_w16934_
	);
	LUT2 #(
		.INIT('h8)
	) name6423 (
		\wishbone_bd_ram_mem3_reg[199][26]/P0001 ,
		_w12768_,
		_w16935_
	);
	LUT2 #(
		.INIT('h8)
	) name6424 (
		\wishbone_bd_ram_mem3_reg[194][26]/P0001 ,
		_w12772_,
		_w16936_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		\wishbone_bd_ram_mem3_reg[179][26]/P0001 ,
		_w13050_,
		_w16937_
	);
	LUT2 #(
		.INIT('h8)
	) name6426 (
		\wishbone_bd_ram_mem3_reg[6][26]/P0001 ,
		_w12968_,
		_w16938_
	);
	LUT2 #(
		.INIT('h8)
	) name6427 (
		\wishbone_bd_ram_mem3_reg[173][26]/P0001 ,
		_w12854_,
		_w16939_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		\wishbone_bd_ram_mem3_reg[34][26]/P0001 ,
		_w12930_,
		_w16940_
	);
	LUT2 #(
		.INIT('h8)
	) name6429 (
		\wishbone_bd_ram_mem3_reg[134][26]/P0001 ,
		_w12763_,
		_w16941_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		\wishbone_bd_ram_mem3_reg[121][26]/P0001 ,
		_w13078_,
		_w16942_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		\wishbone_bd_ram_mem3_reg[21][26]/P0001 ,
		_w12906_,
		_w16943_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		\wishbone_bd_ram_mem3_reg[101][26]/P0001 ,
		_w13192_,
		_w16944_
	);
	LUT2 #(
		.INIT('h8)
	) name6433 (
		\wishbone_bd_ram_mem3_reg[198][26]/P0001 ,
		_w12832_,
		_w16945_
	);
	LUT2 #(
		.INIT('h8)
	) name6434 (
		\wishbone_bd_ram_mem3_reg[144][26]/P0001 ,
		_w12756_,
		_w16946_
	);
	LUT2 #(
		.INIT('h8)
	) name6435 (
		\wishbone_bd_ram_mem3_reg[170][26]/P0001 ,
		_w13030_,
		_w16947_
	);
	LUT2 #(
		.INIT('h8)
	) name6436 (
		\wishbone_bd_ram_mem3_reg[115][26]/P0001 ,
		_w13112_,
		_w16948_
	);
	LUT2 #(
		.INIT('h8)
	) name6437 (
		\wishbone_bd_ram_mem3_reg[181][26]/P0001 ,
		_w12828_,
		_w16949_
	);
	LUT2 #(
		.INIT('h8)
	) name6438 (
		\wishbone_bd_ram_mem3_reg[234][26]/P0001 ,
		_w13214_,
		_w16950_
	);
	LUT2 #(
		.INIT('h8)
	) name6439 (
		\wishbone_bd_ram_mem3_reg[158][26]/P0001 ,
		_w12898_,
		_w16951_
	);
	LUT2 #(
		.INIT('h8)
	) name6440 (
		\wishbone_bd_ram_mem3_reg[79][26]/P0001 ,
		_w13212_,
		_w16952_
	);
	LUT2 #(
		.INIT('h8)
	) name6441 (
		\wishbone_bd_ram_mem3_reg[232][26]/P0001 ,
		_w12758_,
		_w16953_
	);
	LUT2 #(
		.INIT('h8)
	) name6442 (
		\wishbone_bd_ram_mem3_reg[122][26]/P0001 ,
		_w13130_,
		_w16954_
	);
	LUT2 #(
		.INIT('h8)
	) name6443 (
		\wishbone_bd_ram_mem3_reg[197][26]/P0001 ,
		_w12834_,
		_w16955_
	);
	LUT2 #(
		.INIT('h8)
	) name6444 (
		\wishbone_bd_ram_mem3_reg[236][26]/P0001 ,
		_w12731_,
		_w16956_
	);
	LUT2 #(
		.INIT('h8)
	) name6445 (
		\wishbone_bd_ram_mem3_reg[5][26]/P0001 ,
		_w12878_,
		_w16957_
	);
	LUT2 #(
		.INIT('h8)
	) name6446 (
		\wishbone_bd_ram_mem3_reg[106][26]/P0001 ,
		_w12713_,
		_w16958_
	);
	LUT2 #(
		.INIT('h8)
	) name6447 (
		\wishbone_bd_ram_mem3_reg[184][26]/P0001 ,
		_w13062_,
		_w16959_
	);
	LUT2 #(
		.INIT('h8)
	) name6448 (
		\wishbone_bd_ram_mem3_reg[245][26]/P0001 ,
		_w13022_,
		_w16960_
	);
	LUT2 #(
		.INIT('h8)
	) name6449 (
		\wishbone_bd_ram_mem3_reg[164][26]/P0001 ,
		_w12876_,
		_w16961_
	);
	LUT2 #(
		.INIT('h8)
	) name6450 (
		\wishbone_bd_ram_mem3_reg[246][26]/P0001 ,
		_w13076_,
		_w16962_
	);
	LUT2 #(
		.INIT('h8)
	) name6451 (
		\wishbone_bd_ram_mem3_reg[95][26]/P0001 ,
		_w12844_,
		_w16963_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		\wishbone_bd_ram_mem3_reg[85][26]/P0001 ,
		_w13216_,
		_w16964_
	);
	LUT2 #(
		.INIT('h8)
	) name6453 (
		\wishbone_bd_ram_mem3_reg[46][26]/P0001 ,
		_w12884_,
		_w16965_
	);
	LUT2 #(
		.INIT('h8)
	) name6454 (
		\wishbone_bd_ram_mem3_reg[44][26]/P0001 ,
		_w12896_,
		_w16966_
	);
	LUT2 #(
		.INIT('h8)
	) name6455 (
		\wishbone_bd_ram_mem3_reg[35][26]/P0001 ,
		_w12703_,
		_w16967_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		\wishbone_bd_ram_mem3_reg[219][26]/P0001 ,
		_w12806_,
		_w16968_
	);
	LUT2 #(
		.INIT('h8)
	) name6457 (
		\wishbone_bd_ram_mem3_reg[45][26]/P0001 ,
		_w12908_,
		_w16969_
	);
	LUT2 #(
		.INIT('h8)
	) name6458 (
		\wishbone_bd_ram_mem3_reg[94][26]/P0001 ,
		_w13186_,
		_w16970_
	);
	LUT2 #(
		.INIT('h8)
	) name6459 (
		\wishbone_bd_ram_mem3_reg[222][26]/P0001 ,
		_w13094_,
		_w16971_
	);
	LUT2 #(
		.INIT('h8)
	) name6460 (
		\wishbone_bd_ram_mem3_reg[241][26]/P0001 ,
		_w13006_,
		_w16972_
	);
	LUT2 #(
		.INIT('h8)
	) name6461 (
		\wishbone_bd_ram_mem3_reg[42][26]/P0001 ,
		_w12842_,
		_w16973_
	);
	LUT2 #(
		.INIT('h8)
	) name6462 (
		\wishbone_bd_ram_mem3_reg[17][26]/P0001 ,
		_w12848_,
		_w16974_
	);
	LUT2 #(
		.INIT('h8)
	) name6463 (
		\wishbone_bd_ram_mem3_reg[38][26]/P0001 ,
		_w13182_,
		_w16975_
	);
	LUT2 #(
		.INIT('h8)
	) name6464 (
		\wishbone_bd_ram_mem3_reg[167][26]/P0001 ,
		_w12986_,
		_w16976_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		\wishbone_bd_ram_mem3_reg[14][26]/P0001 ,
		_w13086_,
		_w16977_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		\wishbone_bd_ram_mem3_reg[25][26]/P0001 ,
		_w13108_,
		_w16978_
	);
	LUT2 #(
		.INIT('h8)
	) name6467 (
		\wishbone_bd_ram_mem3_reg[31][26]/P0001 ,
		_w13198_,
		_w16979_
	);
	LUT2 #(
		.INIT('h8)
	) name6468 (
		\wishbone_bd_ram_mem3_reg[68][26]/P0001 ,
		_w12946_,
		_w16980_
	);
	LUT2 #(
		.INIT('h8)
	) name6469 (
		\wishbone_bd_ram_mem3_reg[58][26]/P0001 ,
		_w13070_,
		_w16981_
	);
	LUT2 #(
		.INIT('h8)
	) name6470 (
		\wishbone_bd_ram_mem3_reg[91][26]/P0001 ,
		_w13074_,
		_w16982_
	);
	LUT2 #(
		.INIT('h8)
	) name6471 (
		\wishbone_bd_ram_mem3_reg[74][26]/P0001 ,
		_w12812_,
		_w16983_
	);
	LUT2 #(
		.INIT('h8)
	) name6472 (
		\wishbone_bd_ram_mem3_reg[118][26]/P0001 ,
		_w12830_,
		_w16984_
	);
	LUT2 #(
		.INIT('h8)
	) name6473 (
		\wishbone_bd_ram_mem3_reg[37][26]/P0001 ,
		_w13102_,
		_w16985_
	);
	LUT2 #(
		.INIT('h8)
	) name6474 (
		\wishbone_bd_ram_mem3_reg[190][26]/P0001 ,
		_w12858_,
		_w16986_
	);
	LUT2 #(
		.INIT('h8)
	) name6475 (
		\wishbone_bd_ram_mem3_reg[210][26]/P0001 ,
		_w12924_,
		_w16987_
	);
	LUT2 #(
		.INIT('h8)
	) name6476 (
		\wishbone_bd_ram_mem3_reg[39][26]/P0001 ,
		_w13018_,
		_w16988_
	);
	LUT2 #(
		.INIT('h8)
	) name6477 (
		\wishbone_bd_ram_mem3_reg[244][26]/P0001 ,
		_w12747_,
		_w16989_
	);
	LUT2 #(
		.INIT('h8)
	) name6478 (
		\wishbone_bd_ram_mem3_reg[23][26]/P0001 ,
		_w13008_,
		_w16990_
	);
	LUT2 #(
		.INIT('h8)
	) name6479 (
		\wishbone_bd_ram_mem3_reg[238][26]/P0001 ,
		_w13160_,
		_w16991_
	);
	LUT2 #(
		.INIT('h8)
	) name6480 (
		\wishbone_bd_ram_mem3_reg[61][26]/P0001 ,
		_w12725_,
		_w16992_
	);
	LUT2 #(
		.INIT('h8)
	) name6481 (
		\wishbone_bd_ram_mem3_reg[52][26]/P0001 ,
		_w13082_,
		_w16993_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		\wishbone_bd_ram_mem3_reg[162][26]/P0001 ,
		_w13098_,
		_w16994_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		\wishbone_bd_ram_mem3_reg[109][26]/P0001 ,
		_w12888_,
		_w16995_
	);
	LUT2 #(
		.INIT('h8)
	) name6484 (
		\wishbone_bd_ram_mem3_reg[130][26]/P0001 ,
		_w12914_,
		_w16996_
	);
	LUT2 #(
		.INIT('h8)
	) name6485 (
		\wishbone_bd_ram_mem3_reg[13][26]/P0001 ,
		_w13178_,
		_w16997_
	);
	LUT2 #(
		.INIT('h8)
	) name6486 (
		\wishbone_bd_ram_mem3_reg[224][26]/P0001 ,
		_w12902_,
		_w16998_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		\wishbone_bd_ram_mem3_reg[117][26]/P0001 ,
		_w12715_,
		_w16999_
	);
	LUT2 #(
		.INIT('h8)
	) name6488 (
		\wishbone_bd_ram_mem3_reg[174][26]/P0001 ,
		_w12972_,
		_w17000_
	);
	LUT2 #(
		.INIT('h8)
	) name6489 (
		\wishbone_bd_ram_mem3_reg[211][26]/P0001 ,
		_w13166_,
		_w17001_
	);
	LUT2 #(
		.INIT('h8)
	) name6490 (
		\wishbone_bd_ram_mem3_reg[195][26]/P0001 ,
		_w13144_,
		_w17002_
	);
	LUT2 #(
		.INIT('h8)
	) name6491 (
		\wishbone_bd_ram_mem3_reg[243][26]/P0001 ,
		_w12804_,
		_w17003_
	);
	LUT2 #(
		.INIT('h8)
	) name6492 (
		\wishbone_bd_ram_mem3_reg[183][26]/P0001 ,
		_w12787_,
		_w17004_
	);
	LUT2 #(
		.INIT('h8)
	) name6493 (
		\wishbone_bd_ram_mem3_reg[126][26]/P0001 ,
		_w13218_,
		_w17005_
	);
	LUT2 #(
		.INIT('h8)
	) name6494 (
		\wishbone_bd_ram_mem3_reg[142][26]/P0001 ,
		_w12928_,
		_w17006_
	);
	LUT2 #(
		.INIT('h8)
	) name6495 (
		\wishbone_bd_ram_mem3_reg[172][26]/P0001 ,
		_w12944_,
		_w17007_
	);
	LUT2 #(
		.INIT('h8)
	) name6496 (
		\wishbone_bd_ram_mem3_reg[73][26]/P0001 ,
		_w12918_,
		_w17008_
	);
	LUT2 #(
		.INIT('h8)
	) name6497 (
		\wishbone_bd_ram_mem3_reg[24][26]/P0001 ,
		_w13084_,
		_w17009_
	);
	LUT2 #(
		.INIT('h8)
	) name6498 (
		\wishbone_bd_ram_mem3_reg[33][26]/P0001 ,
		_w12980_,
		_w17010_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		\wishbone_bd_ram_mem3_reg[8][26]/P0001 ,
		_w12920_,
		_w17011_
	);
	LUT2 #(
		.INIT('h8)
	) name6500 (
		\wishbone_bd_ram_mem3_reg[240][26]/P0001 ,
		_w12864_,
		_w17012_
	);
	LUT2 #(
		.INIT('h8)
	) name6501 (
		\wishbone_bd_ram_mem3_reg[69][26]/P0001 ,
		_w12738_,
		_w17013_
	);
	LUT2 #(
		.INIT('h8)
	) name6502 (
		\wishbone_bd_ram_mem3_reg[154][26]/P0001 ,
		_w12962_,
		_w17014_
	);
	LUT2 #(
		.INIT('h8)
	) name6503 (
		\wishbone_bd_ram_mem3_reg[110][26]/P0001 ,
		_w13046_,
		_w17015_
	);
	LUT2 #(
		.INIT('h8)
	) name6504 (
		\wishbone_bd_ram_mem3_reg[249][26]/P0001 ,
		_w12900_,
		_w17016_
	);
	LUT2 #(
		.INIT('h8)
	) name6505 (
		\wishbone_bd_ram_mem3_reg[230][26]/P0001 ,
		_w13036_,
		_w17017_
	);
	LUT2 #(
		.INIT('h8)
	) name6506 (
		\wishbone_bd_ram_mem3_reg[163][26]/P0001 ,
		_w12882_,
		_w17018_
	);
	LUT2 #(
		.INIT('h8)
	) name6507 (
		\wishbone_bd_ram_mem3_reg[66][26]/P0001 ,
		_w12824_,
		_w17019_
	);
	LUT2 #(
		.INIT('h8)
	) name6508 (
		\wishbone_bd_ram_mem3_reg[213][26]/P0001 ,
		_w13002_,
		_w17020_
	);
	LUT2 #(
		.INIT('h8)
	) name6509 (
		\wishbone_bd_ram_mem3_reg[168][26]/P0001 ,
		_w13208_,
		_w17021_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		\wishbone_bd_ram_mem3_reg[0][26]/P0001 ,
		_w12717_,
		_w17022_
	);
	LUT2 #(
		.INIT('h8)
	) name6511 (
		\wishbone_bd_ram_mem3_reg[175][26]/P0001 ,
		_w13126_,
		_w17023_
	);
	LUT2 #(
		.INIT('h8)
	) name6512 (
		\wishbone_bd_ram_mem3_reg[4][26]/P0001 ,
		_w12666_,
		_w17024_
	);
	LUT2 #(
		.INIT('h8)
	) name6513 (
		\wishbone_bd_ram_mem3_reg[116][26]/P0001 ,
		_w12998_,
		_w17025_
	);
	LUT2 #(
		.INIT('h8)
	) name6514 (
		\wishbone_bd_ram_mem3_reg[150][26]/P0001 ,
		_w13136_,
		_w17026_
	);
	LUT2 #(
		.INIT('h8)
	) name6515 (
		\wishbone_bd_ram_mem3_reg[187][26]/P0001 ,
		_w13196_,
		_w17027_
	);
	LUT2 #(
		.INIT('h8)
	) name6516 (
		\wishbone_bd_ram_mem3_reg[2][26]/P0001 ,
		_w13088_,
		_w17028_
	);
	LUT2 #(
		.INIT('h8)
	) name6517 (
		\wishbone_bd_ram_mem3_reg[218][26]/P0001 ,
		_w13206_,
		_w17029_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		\wishbone_bd_ram_mem3_reg[149][26]/P0001 ,
		_w12741_,
		_w17030_
	);
	LUT2 #(
		.INIT('h8)
	) name6519 (
		\wishbone_bd_ram_mem3_reg[235][26]/P0001 ,
		_w12696_,
		_w17031_
	);
	LUT2 #(
		.INIT('h1)
	) name6520 (
		_w16776_,
		_w16777_,
		_w17032_
	);
	LUT2 #(
		.INIT('h1)
	) name6521 (
		_w16778_,
		_w16779_,
		_w17033_
	);
	LUT2 #(
		.INIT('h1)
	) name6522 (
		_w16780_,
		_w16781_,
		_w17034_
	);
	LUT2 #(
		.INIT('h1)
	) name6523 (
		_w16782_,
		_w16783_,
		_w17035_
	);
	LUT2 #(
		.INIT('h1)
	) name6524 (
		_w16784_,
		_w16785_,
		_w17036_
	);
	LUT2 #(
		.INIT('h1)
	) name6525 (
		_w16786_,
		_w16787_,
		_w17037_
	);
	LUT2 #(
		.INIT('h1)
	) name6526 (
		_w16788_,
		_w16789_,
		_w17038_
	);
	LUT2 #(
		.INIT('h1)
	) name6527 (
		_w16790_,
		_w16791_,
		_w17039_
	);
	LUT2 #(
		.INIT('h1)
	) name6528 (
		_w16792_,
		_w16793_,
		_w17040_
	);
	LUT2 #(
		.INIT('h1)
	) name6529 (
		_w16794_,
		_w16795_,
		_w17041_
	);
	LUT2 #(
		.INIT('h1)
	) name6530 (
		_w16796_,
		_w16797_,
		_w17042_
	);
	LUT2 #(
		.INIT('h1)
	) name6531 (
		_w16798_,
		_w16799_,
		_w17043_
	);
	LUT2 #(
		.INIT('h1)
	) name6532 (
		_w16800_,
		_w16801_,
		_w17044_
	);
	LUT2 #(
		.INIT('h1)
	) name6533 (
		_w16802_,
		_w16803_,
		_w17045_
	);
	LUT2 #(
		.INIT('h1)
	) name6534 (
		_w16804_,
		_w16805_,
		_w17046_
	);
	LUT2 #(
		.INIT('h1)
	) name6535 (
		_w16806_,
		_w16807_,
		_w17047_
	);
	LUT2 #(
		.INIT('h1)
	) name6536 (
		_w16808_,
		_w16809_,
		_w17048_
	);
	LUT2 #(
		.INIT('h1)
	) name6537 (
		_w16810_,
		_w16811_,
		_w17049_
	);
	LUT2 #(
		.INIT('h1)
	) name6538 (
		_w16812_,
		_w16813_,
		_w17050_
	);
	LUT2 #(
		.INIT('h1)
	) name6539 (
		_w16814_,
		_w16815_,
		_w17051_
	);
	LUT2 #(
		.INIT('h1)
	) name6540 (
		_w16816_,
		_w16817_,
		_w17052_
	);
	LUT2 #(
		.INIT('h1)
	) name6541 (
		_w16818_,
		_w16819_,
		_w17053_
	);
	LUT2 #(
		.INIT('h1)
	) name6542 (
		_w16820_,
		_w16821_,
		_w17054_
	);
	LUT2 #(
		.INIT('h1)
	) name6543 (
		_w16822_,
		_w16823_,
		_w17055_
	);
	LUT2 #(
		.INIT('h1)
	) name6544 (
		_w16824_,
		_w16825_,
		_w17056_
	);
	LUT2 #(
		.INIT('h1)
	) name6545 (
		_w16826_,
		_w16827_,
		_w17057_
	);
	LUT2 #(
		.INIT('h1)
	) name6546 (
		_w16828_,
		_w16829_,
		_w17058_
	);
	LUT2 #(
		.INIT('h1)
	) name6547 (
		_w16830_,
		_w16831_,
		_w17059_
	);
	LUT2 #(
		.INIT('h1)
	) name6548 (
		_w16832_,
		_w16833_,
		_w17060_
	);
	LUT2 #(
		.INIT('h1)
	) name6549 (
		_w16834_,
		_w16835_,
		_w17061_
	);
	LUT2 #(
		.INIT('h1)
	) name6550 (
		_w16836_,
		_w16837_,
		_w17062_
	);
	LUT2 #(
		.INIT('h1)
	) name6551 (
		_w16838_,
		_w16839_,
		_w17063_
	);
	LUT2 #(
		.INIT('h1)
	) name6552 (
		_w16840_,
		_w16841_,
		_w17064_
	);
	LUT2 #(
		.INIT('h1)
	) name6553 (
		_w16842_,
		_w16843_,
		_w17065_
	);
	LUT2 #(
		.INIT('h1)
	) name6554 (
		_w16844_,
		_w16845_,
		_w17066_
	);
	LUT2 #(
		.INIT('h1)
	) name6555 (
		_w16846_,
		_w16847_,
		_w17067_
	);
	LUT2 #(
		.INIT('h1)
	) name6556 (
		_w16848_,
		_w16849_,
		_w17068_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		_w16850_,
		_w16851_,
		_w17069_
	);
	LUT2 #(
		.INIT('h1)
	) name6558 (
		_w16852_,
		_w16853_,
		_w17070_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		_w16854_,
		_w16855_,
		_w17071_
	);
	LUT2 #(
		.INIT('h1)
	) name6560 (
		_w16856_,
		_w16857_,
		_w17072_
	);
	LUT2 #(
		.INIT('h1)
	) name6561 (
		_w16858_,
		_w16859_,
		_w17073_
	);
	LUT2 #(
		.INIT('h1)
	) name6562 (
		_w16860_,
		_w16861_,
		_w17074_
	);
	LUT2 #(
		.INIT('h1)
	) name6563 (
		_w16862_,
		_w16863_,
		_w17075_
	);
	LUT2 #(
		.INIT('h1)
	) name6564 (
		_w16864_,
		_w16865_,
		_w17076_
	);
	LUT2 #(
		.INIT('h1)
	) name6565 (
		_w16866_,
		_w16867_,
		_w17077_
	);
	LUT2 #(
		.INIT('h1)
	) name6566 (
		_w16868_,
		_w16869_,
		_w17078_
	);
	LUT2 #(
		.INIT('h1)
	) name6567 (
		_w16870_,
		_w16871_,
		_w17079_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		_w16872_,
		_w16873_,
		_w17080_
	);
	LUT2 #(
		.INIT('h1)
	) name6569 (
		_w16874_,
		_w16875_,
		_w17081_
	);
	LUT2 #(
		.INIT('h1)
	) name6570 (
		_w16876_,
		_w16877_,
		_w17082_
	);
	LUT2 #(
		.INIT('h1)
	) name6571 (
		_w16878_,
		_w16879_,
		_w17083_
	);
	LUT2 #(
		.INIT('h1)
	) name6572 (
		_w16880_,
		_w16881_,
		_w17084_
	);
	LUT2 #(
		.INIT('h1)
	) name6573 (
		_w16882_,
		_w16883_,
		_w17085_
	);
	LUT2 #(
		.INIT('h1)
	) name6574 (
		_w16884_,
		_w16885_,
		_w17086_
	);
	LUT2 #(
		.INIT('h1)
	) name6575 (
		_w16886_,
		_w16887_,
		_w17087_
	);
	LUT2 #(
		.INIT('h1)
	) name6576 (
		_w16888_,
		_w16889_,
		_w17088_
	);
	LUT2 #(
		.INIT('h1)
	) name6577 (
		_w16890_,
		_w16891_,
		_w17089_
	);
	LUT2 #(
		.INIT('h1)
	) name6578 (
		_w16892_,
		_w16893_,
		_w17090_
	);
	LUT2 #(
		.INIT('h1)
	) name6579 (
		_w16894_,
		_w16895_,
		_w17091_
	);
	LUT2 #(
		.INIT('h1)
	) name6580 (
		_w16896_,
		_w16897_,
		_w17092_
	);
	LUT2 #(
		.INIT('h1)
	) name6581 (
		_w16898_,
		_w16899_,
		_w17093_
	);
	LUT2 #(
		.INIT('h1)
	) name6582 (
		_w16900_,
		_w16901_,
		_w17094_
	);
	LUT2 #(
		.INIT('h1)
	) name6583 (
		_w16902_,
		_w16903_,
		_w17095_
	);
	LUT2 #(
		.INIT('h1)
	) name6584 (
		_w16904_,
		_w16905_,
		_w17096_
	);
	LUT2 #(
		.INIT('h1)
	) name6585 (
		_w16906_,
		_w16907_,
		_w17097_
	);
	LUT2 #(
		.INIT('h1)
	) name6586 (
		_w16908_,
		_w16909_,
		_w17098_
	);
	LUT2 #(
		.INIT('h1)
	) name6587 (
		_w16910_,
		_w16911_,
		_w17099_
	);
	LUT2 #(
		.INIT('h1)
	) name6588 (
		_w16912_,
		_w16913_,
		_w17100_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w16914_,
		_w16915_,
		_w17101_
	);
	LUT2 #(
		.INIT('h1)
	) name6590 (
		_w16916_,
		_w16917_,
		_w17102_
	);
	LUT2 #(
		.INIT('h1)
	) name6591 (
		_w16918_,
		_w16919_,
		_w17103_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		_w16920_,
		_w16921_,
		_w17104_
	);
	LUT2 #(
		.INIT('h1)
	) name6593 (
		_w16922_,
		_w16923_,
		_w17105_
	);
	LUT2 #(
		.INIT('h1)
	) name6594 (
		_w16924_,
		_w16925_,
		_w17106_
	);
	LUT2 #(
		.INIT('h1)
	) name6595 (
		_w16926_,
		_w16927_,
		_w17107_
	);
	LUT2 #(
		.INIT('h1)
	) name6596 (
		_w16928_,
		_w16929_,
		_w17108_
	);
	LUT2 #(
		.INIT('h1)
	) name6597 (
		_w16930_,
		_w16931_,
		_w17109_
	);
	LUT2 #(
		.INIT('h1)
	) name6598 (
		_w16932_,
		_w16933_,
		_w17110_
	);
	LUT2 #(
		.INIT('h1)
	) name6599 (
		_w16934_,
		_w16935_,
		_w17111_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w16936_,
		_w16937_,
		_w17112_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		_w16938_,
		_w16939_,
		_w17113_
	);
	LUT2 #(
		.INIT('h1)
	) name6602 (
		_w16940_,
		_w16941_,
		_w17114_
	);
	LUT2 #(
		.INIT('h1)
	) name6603 (
		_w16942_,
		_w16943_,
		_w17115_
	);
	LUT2 #(
		.INIT('h1)
	) name6604 (
		_w16944_,
		_w16945_,
		_w17116_
	);
	LUT2 #(
		.INIT('h1)
	) name6605 (
		_w16946_,
		_w16947_,
		_w17117_
	);
	LUT2 #(
		.INIT('h1)
	) name6606 (
		_w16948_,
		_w16949_,
		_w17118_
	);
	LUT2 #(
		.INIT('h1)
	) name6607 (
		_w16950_,
		_w16951_,
		_w17119_
	);
	LUT2 #(
		.INIT('h1)
	) name6608 (
		_w16952_,
		_w16953_,
		_w17120_
	);
	LUT2 #(
		.INIT('h1)
	) name6609 (
		_w16954_,
		_w16955_,
		_w17121_
	);
	LUT2 #(
		.INIT('h1)
	) name6610 (
		_w16956_,
		_w16957_,
		_w17122_
	);
	LUT2 #(
		.INIT('h1)
	) name6611 (
		_w16958_,
		_w16959_,
		_w17123_
	);
	LUT2 #(
		.INIT('h1)
	) name6612 (
		_w16960_,
		_w16961_,
		_w17124_
	);
	LUT2 #(
		.INIT('h1)
	) name6613 (
		_w16962_,
		_w16963_,
		_w17125_
	);
	LUT2 #(
		.INIT('h1)
	) name6614 (
		_w16964_,
		_w16965_,
		_w17126_
	);
	LUT2 #(
		.INIT('h1)
	) name6615 (
		_w16966_,
		_w16967_,
		_w17127_
	);
	LUT2 #(
		.INIT('h1)
	) name6616 (
		_w16968_,
		_w16969_,
		_w17128_
	);
	LUT2 #(
		.INIT('h1)
	) name6617 (
		_w16970_,
		_w16971_,
		_w17129_
	);
	LUT2 #(
		.INIT('h1)
	) name6618 (
		_w16972_,
		_w16973_,
		_w17130_
	);
	LUT2 #(
		.INIT('h1)
	) name6619 (
		_w16974_,
		_w16975_,
		_w17131_
	);
	LUT2 #(
		.INIT('h1)
	) name6620 (
		_w16976_,
		_w16977_,
		_w17132_
	);
	LUT2 #(
		.INIT('h1)
	) name6621 (
		_w16978_,
		_w16979_,
		_w17133_
	);
	LUT2 #(
		.INIT('h1)
	) name6622 (
		_w16980_,
		_w16981_,
		_w17134_
	);
	LUT2 #(
		.INIT('h1)
	) name6623 (
		_w16982_,
		_w16983_,
		_w17135_
	);
	LUT2 #(
		.INIT('h1)
	) name6624 (
		_w16984_,
		_w16985_,
		_w17136_
	);
	LUT2 #(
		.INIT('h1)
	) name6625 (
		_w16986_,
		_w16987_,
		_w17137_
	);
	LUT2 #(
		.INIT('h1)
	) name6626 (
		_w16988_,
		_w16989_,
		_w17138_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		_w16990_,
		_w16991_,
		_w17139_
	);
	LUT2 #(
		.INIT('h1)
	) name6628 (
		_w16992_,
		_w16993_,
		_w17140_
	);
	LUT2 #(
		.INIT('h1)
	) name6629 (
		_w16994_,
		_w16995_,
		_w17141_
	);
	LUT2 #(
		.INIT('h1)
	) name6630 (
		_w16996_,
		_w16997_,
		_w17142_
	);
	LUT2 #(
		.INIT('h1)
	) name6631 (
		_w16998_,
		_w16999_,
		_w17143_
	);
	LUT2 #(
		.INIT('h1)
	) name6632 (
		_w17000_,
		_w17001_,
		_w17144_
	);
	LUT2 #(
		.INIT('h1)
	) name6633 (
		_w17002_,
		_w17003_,
		_w17145_
	);
	LUT2 #(
		.INIT('h1)
	) name6634 (
		_w17004_,
		_w17005_,
		_w17146_
	);
	LUT2 #(
		.INIT('h1)
	) name6635 (
		_w17006_,
		_w17007_,
		_w17147_
	);
	LUT2 #(
		.INIT('h1)
	) name6636 (
		_w17008_,
		_w17009_,
		_w17148_
	);
	LUT2 #(
		.INIT('h1)
	) name6637 (
		_w17010_,
		_w17011_,
		_w17149_
	);
	LUT2 #(
		.INIT('h1)
	) name6638 (
		_w17012_,
		_w17013_,
		_w17150_
	);
	LUT2 #(
		.INIT('h1)
	) name6639 (
		_w17014_,
		_w17015_,
		_w17151_
	);
	LUT2 #(
		.INIT('h1)
	) name6640 (
		_w17016_,
		_w17017_,
		_w17152_
	);
	LUT2 #(
		.INIT('h1)
	) name6641 (
		_w17018_,
		_w17019_,
		_w17153_
	);
	LUT2 #(
		.INIT('h1)
	) name6642 (
		_w17020_,
		_w17021_,
		_w17154_
	);
	LUT2 #(
		.INIT('h1)
	) name6643 (
		_w17022_,
		_w17023_,
		_w17155_
	);
	LUT2 #(
		.INIT('h1)
	) name6644 (
		_w17024_,
		_w17025_,
		_w17156_
	);
	LUT2 #(
		.INIT('h1)
	) name6645 (
		_w17026_,
		_w17027_,
		_w17157_
	);
	LUT2 #(
		.INIT('h1)
	) name6646 (
		_w17028_,
		_w17029_,
		_w17158_
	);
	LUT2 #(
		.INIT('h1)
	) name6647 (
		_w17030_,
		_w17031_,
		_w17159_
	);
	LUT2 #(
		.INIT('h8)
	) name6648 (
		_w17158_,
		_w17159_,
		_w17160_
	);
	LUT2 #(
		.INIT('h8)
	) name6649 (
		_w17156_,
		_w17157_,
		_w17161_
	);
	LUT2 #(
		.INIT('h8)
	) name6650 (
		_w17154_,
		_w17155_,
		_w17162_
	);
	LUT2 #(
		.INIT('h8)
	) name6651 (
		_w17152_,
		_w17153_,
		_w17163_
	);
	LUT2 #(
		.INIT('h8)
	) name6652 (
		_w17150_,
		_w17151_,
		_w17164_
	);
	LUT2 #(
		.INIT('h8)
	) name6653 (
		_w17148_,
		_w17149_,
		_w17165_
	);
	LUT2 #(
		.INIT('h8)
	) name6654 (
		_w17146_,
		_w17147_,
		_w17166_
	);
	LUT2 #(
		.INIT('h8)
	) name6655 (
		_w17144_,
		_w17145_,
		_w17167_
	);
	LUT2 #(
		.INIT('h8)
	) name6656 (
		_w17142_,
		_w17143_,
		_w17168_
	);
	LUT2 #(
		.INIT('h8)
	) name6657 (
		_w17140_,
		_w17141_,
		_w17169_
	);
	LUT2 #(
		.INIT('h8)
	) name6658 (
		_w17138_,
		_w17139_,
		_w17170_
	);
	LUT2 #(
		.INIT('h8)
	) name6659 (
		_w17136_,
		_w17137_,
		_w17171_
	);
	LUT2 #(
		.INIT('h8)
	) name6660 (
		_w17134_,
		_w17135_,
		_w17172_
	);
	LUT2 #(
		.INIT('h8)
	) name6661 (
		_w17132_,
		_w17133_,
		_w17173_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		_w17130_,
		_w17131_,
		_w17174_
	);
	LUT2 #(
		.INIT('h8)
	) name6663 (
		_w17128_,
		_w17129_,
		_w17175_
	);
	LUT2 #(
		.INIT('h8)
	) name6664 (
		_w17126_,
		_w17127_,
		_w17176_
	);
	LUT2 #(
		.INIT('h8)
	) name6665 (
		_w17124_,
		_w17125_,
		_w17177_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		_w17122_,
		_w17123_,
		_w17178_
	);
	LUT2 #(
		.INIT('h8)
	) name6667 (
		_w17120_,
		_w17121_,
		_w17179_
	);
	LUT2 #(
		.INIT('h8)
	) name6668 (
		_w17118_,
		_w17119_,
		_w17180_
	);
	LUT2 #(
		.INIT('h8)
	) name6669 (
		_w17116_,
		_w17117_,
		_w17181_
	);
	LUT2 #(
		.INIT('h8)
	) name6670 (
		_w17114_,
		_w17115_,
		_w17182_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		_w17112_,
		_w17113_,
		_w17183_
	);
	LUT2 #(
		.INIT('h8)
	) name6672 (
		_w17110_,
		_w17111_,
		_w17184_
	);
	LUT2 #(
		.INIT('h8)
	) name6673 (
		_w17108_,
		_w17109_,
		_w17185_
	);
	LUT2 #(
		.INIT('h8)
	) name6674 (
		_w17106_,
		_w17107_,
		_w17186_
	);
	LUT2 #(
		.INIT('h8)
	) name6675 (
		_w17104_,
		_w17105_,
		_w17187_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		_w17102_,
		_w17103_,
		_w17188_
	);
	LUT2 #(
		.INIT('h8)
	) name6677 (
		_w17100_,
		_w17101_,
		_w17189_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		_w17098_,
		_w17099_,
		_w17190_
	);
	LUT2 #(
		.INIT('h8)
	) name6679 (
		_w17096_,
		_w17097_,
		_w17191_
	);
	LUT2 #(
		.INIT('h8)
	) name6680 (
		_w17094_,
		_w17095_,
		_w17192_
	);
	LUT2 #(
		.INIT('h8)
	) name6681 (
		_w17092_,
		_w17093_,
		_w17193_
	);
	LUT2 #(
		.INIT('h8)
	) name6682 (
		_w17090_,
		_w17091_,
		_w17194_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		_w17088_,
		_w17089_,
		_w17195_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		_w17086_,
		_w17087_,
		_w17196_
	);
	LUT2 #(
		.INIT('h8)
	) name6685 (
		_w17084_,
		_w17085_,
		_w17197_
	);
	LUT2 #(
		.INIT('h8)
	) name6686 (
		_w17082_,
		_w17083_,
		_w17198_
	);
	LUT2 #(
		.INIT('h8)
	) name6687 (
		_w17080_,
		_w17081_,
		_w17199_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		_w17078_,
		_w17079_,
		_w17200_
	);
	LUT2 #(
		.INIT('h8)
	) name6689 (
		_w17076_,
		_w17077_,
		_w17201_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		_w17074_,
		_w17075_,
		_w17202_
	);
	LUT2 #(
		.INIT('h8)
	) name6691 (
		_w17072_,
		_w17073_,
		_w17203_
	);
	LUT2 #(
		.INIT('h8)
	) name6692 (
		_w17070_,
		_w17071_,
		_w17204_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		_w17068_,
		_w17069_,
		_w17205_
	);
	LUT2 #(
		.INIT('h8)
	) name6694 (
		_w17066_,
		_w17067_,
		_w17206_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		_w17064_,
		_w17065_,
		_w17207_
	);
	LUT2 #(
		.INIT('h8)
	) name6696 (
		_w17062_,
		_w17063_,
		_w17208_
	);
	LUT2 #(
		.INIT('h8)
	) name6697 (
		_w17060_,
		_w17061_,
		_w17209_
	);
	LUT2 #(
		.INIT('h8)
	) name6698 (
		_w17058_,
		_w17059_,
		_w17210_
	);
	LUT2 #(
		.INIT('h8)
	) name6699 (
		_w17056_,
		_w17057_,
		_w17211_
	);
	LUT2 #(
		.INIT('h8)
	) name6700 (
		_w17054_,
		_w17055_,
		_w17212_
	);
	LUT2 #(
		.INIT('h8)
	) name6701 (
		_w17052_,
		_w17053_,
		_w17213_
	);
	LUT2 #(
		.INIT('h8)
	) name6702 (
		_w17050_,
		_w17051_,
		_w17214_
	);
	LUT2 #(
		.INIT('h8)
	) name6703 (
		_w17048_,
		_w17049_,
		_w17215_
	);
	LUT2 #(
		.INIT('h8)
	) name6704 (
		_w17046_,
		_w17047_,
		_w17216_
	);
	LUT2 #(
		.INIT('h8)
	) name6705 (
		_w17044_,
		_w17045_,
		_w17217_
	);
	LUT2 #(
		.INIT('h8)
	) name6706 (
		_w17042_,
		_w17043_,
		_w17218_
	);
	LUT2 #(
		.INIT('h8)
	) name6707 (
		_w17040_,
		_w17041_,
		_w17219_
	);
	LUT2 #(
		.INIT('h8)
	) name6708 (
		_w17038_,
		_w17039_,
		_w17220_
	);
	LUT2 #(
		.INIT('h8)
	) name6709 (
		_w17036_,
		_w17037_,
		_w17221_
	);
	LUT2 #(
		.INIT('h8)
	) name6710 (
		_w17034_,
		_w17035_,
		_w17222_
	);
	LUT2 #(
		.INIT('h8)
	) name6711 (
		_w17032_,
		_w17033_,
		_w17223_
	);
	LUT2 #(
		.INIT('h8)
	) name6712 (
		_w17222_,
		_w17223_,
		_w17224_
	);
	LUT2 #(
		.INIT('h8)
	) name6713 (
		_w17220_,
		_w17221_,
		_w17225_
	);
	LUT2 #(
		.INIT('h8)
	) name6714 (
		_w17218_,
		_w17219_,
		_w17226_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		_w17216_,
		_w17217_,
		_w17227_
	);
	LUT2 #(
		.INIT('h8)
	) name6716 (
		_w17214_,
		_w17215_,
		_w17228_
	);
	LUT2 #(
		.INIT('h8)
	) name6717 (
		_w17212_,
		_w17213_,
		_w17229_
	);
	LUT2 #(
		.INIT('h8)
	) name6718 (
		_w17210_,
		_w17211_,
		_w17230_
	);
	LUT2 #(
		.INIT('h8)
	) name6719 (
		_w17208_,
		_w17209_,
		_w17231_
	);
	LUT2 #(
		.INIT('h8)
	) name6720 (
		_w17206_,
		_w17207_,
		_w17232_
	);
	LUT2 #(
		.INIT('h8)
	) name6721 (
		_w17204_,
		_w17205_,
		_w17233_
	);
	LUT2 #(
		.INIT('h8)
	) name6722 (
		_w17202_,
		_w17203_,
		_w17234_
	);
	LUT2 #(
		.INIT('h8)
	) name6723 (
		_w17200_,
		_w17201_,
		_w17235_
	);
	LUT2 #(
		.INIT('h8)
	) name6724 (
		_w17198_,
		_w17199_,
		_w17236_
	);
	LUT2 #(
		.INIT('h8)
	) name6725 (
		_w17196_,
		_w17197_,
		_w17237_
	);
	LUT2 #(
		.INIT('h8)
	) name6726 (
		_w17194_,
		_w17195_,
		_w17238_
	);
	LUT2 #(
		.INIT('h8)
	) name6727 (
		_w17192_,
		_w17193_,
		_w17239_
	);
	LUT2 #(
		.INIT('h8)
	) name6728 (
		_w17190_,
		_w17191_,
		_w17240_
	);
	LUT2 #(
		.INIT('h8)
	) name6729 (
		_w17188_,
		_w17189_,
		_w17241_
	);
	LUT2 #(
		.INIT('h8)
	) name6730 (
		_w17186_,
		_w17187_,
		_w17242_
	);
	LUT2 #(
		.INIT('h8)
	) name6731 (
		_w17184_,
		_w17185_,
		_w17243_
	);
	LUT2 #(
		.INIT('h8)
	) name6732 (
		_w17182_,
		_w17183_,
		_w17244_
	);
	LUT2 #(
		.INIT('h8)
	) name6733 (
		_w17180_,
		_w17181_,
		_w17245_
	);
	LUT2 #(
		.INIT('h8)
	) name6734 (
		_w17178_,
		_w17179_,
		_w17246_
	);
	LUT2 #(
		.INIT('h8)
	) name6735 (
		_w17176_,
		_w17177_,
		_w17247_
	);
	LUT2 #(
		.INIT('h8)
	) name6736 (
		_w17174_,
		_w17175_,
		_w17248_
	);
	LUT2 #(
		.INIT('h8)
	) name6737 (
		_w17172_,
		_w17173_,
		_w17249_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		_w17170_,
		_w17171_,
		_w17250_
	);
	LUT2 #(
		.INIT('h8)
	) name6739 (
		_w17168_,
		_w17169_,
		_w17251_
	);
	LUT2 #(
		.INIT('h8)
	) name6740 (
		_w17166_,
		_w17167_,
		_w17252_
	);
	LUT2 #(
		.INIT('h8)
	) name6741 (
		_w17164_,
		_w17165_,
		_w17253_
	);
	LUT2 #(
		.INIT('h8)
	) name6742 (
		_w17162_,
		_w17163_,
		_w17254_
	);
	LUT2 #(
		.INIT('h8)
	) name6743 (
		_w17160_,
		_w17161_,
		_w17255_
	);
	LUT2 #(
		.INIT('h8)
	) name6744 (
		_w17254_,
		_w17255_,
		_w17256_
	);
	LUT2 #(
		.INIT('h8)
	) name6745 (
		_w17252_,
		_w17253_,
		_w17257_
	);
	LUT2 #(
		.INIT('h8)
	) name6746 (
		_w17250_,
		_w17251_,
		_w17258_
	);
	LUT2 #(
		.INIT('h8)
	) name6747 (
		_w17248_,
		_w17249_,
		_w17259_
	);
	LUT2 #(
		.INIT('h8)
	) name6748 (
		_w17246_,
		_w17247_,
		_w17260_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		_w17244_,
		_w17245_,
		_w17261_
	);
	LUT2 #(
		.INIT('h8)
	) name6750 (
		_w17242_,
		_w17243_,
		_w17262_
	);
	LUT2 #(
		.INIT('h8)
	) name6751 (
		_w17240_,
		_w17241_,
		_w17263_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		_w17238_,
		_w17239_,
		_w17264_
	);
	LUT2 #(
		.INIT('h8)
	) name6753 (
		_w17236_,
		_w17237_,
		_w17265_
	);
	LUT2 #(
		.INIT('h8)
	) name6754 (
		_w17234_,
		_w17235_,
		_w17266_
	);
	LUT2 #(
		.INIT('h8)
	) name6755 (
		_w17232_,
		_w17233_,
		_w17267_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		_w17230_,
		_w17231_,
		_w17268_
	);
	LUT2 #(
		.INIT('h8)
	) name6757 (
		_w17228_,
		_w17229_,
		_w17269_
	);
	LUT2 #(
		.INIT('h8)
	) name6758 (
		_w17226_,
		_w17227_,
		_w17270_
	);
	LUT2 #(
		.INIT('h8)
	) name6759 (
		_w17224_,
		_w17225_,
		_w17271_
	);
	LUT2 #(
		.INIT('h8)
	) name6760 (
		_w17270_,
		_w17271_,
		_w17272_
	);
	LUT2 #(
		.INIT('h8)
	) name6761 (
		_w17268_,
		_w17269_,
		_w17273_
	);
	LUT2 #(
		.INIT('h8)
	) name6762 (
		_w17266_,
		_w17267_,
		_w17274_
	);
	LUT2 #(
		.INIT('h8)
	) name6763 (
		_w17264_,
		_w17265_,
		_w17275_
	);
	LUT2 #(
		.INIT('h8)
	) name6764 (
		_w17262_,
		_w17263_,
		_w17276_
	);
	LUT2 #(
		.INIT('h8)
	) name6765 (
		_w17260_,
		_w17261_,
		_w17277_
	);
	LUT2 #(
		.INIT('h8)
	) name6766 (
		_w17258_,
		_w17259_,
		_w17278_
	);
	LUT2 #(
		.INIT('h8)
	) name6767 (
		_w17256_,
		_w17257_,
		_w17279_
	);
	LUT2 #(
		.INIT('h8)
	) name6768 (
		_w17278_,
		_w17279_,
		_w17280_
	);
	LUT2 #(
		.INIT('h8)
	) name6769 (
		_w17276_,
		_w17277_,
		_w17281_
	);
	LUT2 #(
		.INIT('h8)
	) name6770 (
		_w17274_,
		_w17275_,
		_w17282_
	);
	LUT2 #(
		.INIT('h8)
	) name6771 (
		_w17272_,
		_w17273_,
		_w17283_
	);
	LUT2 #(
		.INIT('h8)
	) name6772 (
		_w17282_,
		_w17283_,
		_w17284_
	);
	LUT2 #(
		.INIT('h8)
	) name6773 (
		_w17280_,
		_w17281_,
		_w17285_
	);
	LUT2 #(
		.INIT('h8)
	) name6774 (
		_w17284_,
		_w17285_,
		_w17286_
	);
	LUT2 #(
		.INIT('h1)
	) name6775 (
		wb_rst_i_pad,
		_w17286_,
		_w17287_
	);
	LUT2 #(
		.INIT('h8)
	) name6776 (
		_w12656_,
		_w17287_,
		_w17288_
	);
	LUT2 #(
		.INIT('h2)
	) name6777 (
		_w12657_,
		_w13489_,
		_w17289_
	);
	LUT2 #(
		.INIT('h8)
	) name6778 (
		_w13484_,
		_w17289_,
		_w17290_
	);
	LUT2 #(
		.INIT('h1)
	) name6779 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		_w17290_,
		_w17291_
	);
	LUT2 #(
		.INIT('h2)
	) name6780 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		_w13489_,
		_w17292_
	);
	LUT2 #(
		.INIT('h1)
	) name6781 (
		_w13498_,
		_w17292_,
		_w17293_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		_w12657_,
		_w13484_,
		_w17294_
	);
	LUT2 #(
		.INIT('h4)
	) name6783 (
		_w17293_,
		_w17294_,
		_w17295_
	);
	LUT2 #(
		.INIT('h1)
	) name6784 (
		_w12656_,
		_w17291_,
		_w17296_
	);
	LUT2 #(
		.INIT('h4)
	) name6785 (
		_w17295_,
		_w17296_,
		_w17297_
	);
	LUT2 #(
		.INIT('h1)
	) name6786 (
		_w17288_,
		_w17297_,
		_w17298_
	);
	LUT2 #(
		.INIT('h8)
	) name6787 (
		\wishbone_bd_ram_mem3_reg[17][25]/P0001 ,
		_w12848_,
		_w17299_
	);
	LUT2 #(
		.INIT('h8)
	) name6788 (
		\wishbone_bd_ram_mem3_reg[235][25]/P0001 ,
		_w12696_,
		_w17300_
	);
	LUT2 #(
		.INIT('h8)
	) name6789 (
		\wishbone_bd_ram_mem3_reg[141][25]/P0001 ,
		_w13004_,
		_w17301_
	);
	LUT2 #(
		.INIT('h8)
	) name6790 (
		\wishbone_bd_ram_mem3_reg[49][25]/P0001 ,
		_w12994_,
		_w17302_
	);
	LUT2 #(
		.INIT('h8)
	) name6791 (
		\wishbone_bd_ram_mem3_reg[57][25]/P0001 ,
		_w13116_,
		_w17303_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		\wishbone_bd_ram_mem3_reg[179][25]/P0001 ,
		_w13050_,
		_w17304_
	);
	LUT2 #(
		.INIT('h8)
	) name6793 (
		\wishbone_bd_ram_mem3_reg[160][25]/P0001 ,
		_w12872_,
		_w17305_
	);
	LUT2 #(
		.INIT('h8)
	) name6794 (
		\wishbone_bd_ram_mem3_reg[169][25]/P0001 ,
		_w12722_,
		_w17306_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		\wishbone_bd_ram_mem3_reg[13][25]/P0001 ,
		_w13178_,
		_w17307_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		\wishbone_bd_ram_mem3_reg[214][25]/P0001 ,
		_w12984_,
		_w17308_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		\wishbone_bd_ram_mem3_reg[156][25]/P0001 ,
		_w13190_,
		_w17309_
	);
	LUT2 #(
		.INIT('h8)
	) name6798 (
		\wishbone_bd_ram_mem3_reg[167][25]/P0001 ,
		_w12986_,
		_w17310_
	);
	LUT2 #(
		.INIT('h8)
	) name6799 (
		\wishbone_bd_ram_mem3_reg[12][25]/P0001 ,
		_w13118_,
		_w17311_
	);
	LUT2 #(
		.INIT('h8)
	) name6800 (
		\wishbone_bd_ram_mem3_reg[237][25]/P0001 ,
		_w12990_,
		_w17312_
	);
	LUT2 #(
		.INIT('h8)
	) name6801 (
		\wishbone_bd_ram_mem3_reg[68][25]/P0001 ,
		_w12946_,
		_w17313_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		\wishbone_bd_ram_mem3_reg[19][25]/P0001 ,
		_w13012_,
		_w17314_
	);
	LUT2 #(
		.INIT('h8)
	) name6803 (
		\wishbone_bd_ram_mem3_reg[130][25]/P0001 ,
		_w12914_,
		_w17315_
	);
	LUT2 #(
		.INIT('h8)
	) name6804 (
		\wishbone_bd_ram_mem3_reg[124][25]/P0001 ,
		_w13058_,
		_w17316_
	);
	LUT2 #(
		.INIT('h8)
	) name6805 (
		\wishbone_bd_ram_mem3_reg[0][25]/P0001 ,
		_w12717_,
		_w17317_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		\wishbone_bd_ram_mem3_reg[5][25]/P0001 ,
		_w12878_,
		_w17318_
	);
	LUT2 #(
		.INIT('h8)
	) name6807 (
		\wishbone_bd_ram_mem3_reg[38][25]/P0001 ,
		_w13182_,
		_w17319_
	);
	LUT2 #(
		.INIT('h8)
	) name6808 (
		\wishbone_bd_ram_mem3_reg[229][25]/P0001 ,
		_w12711_,
		_w17320_
	);
	LUT2 #(
		.INIT('h8)
	) name6809 (
		\wishbone_bd_ram_mem3_reg[126][25]/P0001 ,
		_w13218_,
		_w17321_
	);
	LUT2 #(
		.INIT('h8)
	) name6810 (
		\wishbone_bd_ram_mem3_reg[86][25]/P0001 ,
		_w12735_,
		_w17322_
	);
	LUT2 #(
		.INIT('h8)
	) name6811 (
		\wishbone_bd_ram_mem3_reg[152][25]/P0001 ,
		_w12966_,
		_w17323_
	);
	LUT2 #(
		.INIT('h8)
	) name6812 (
		\wishbone_bd_ram_mem3_reg[230][25]/P0001 ,
		_w13036_,
		_w17324_
	);
	LUT2 #(
		.INIT('h8)
	) name6813 (
		\wishbone_bd_ram_mem3_reg[164][25]/P0001 ,
		_w12876_,
		_w17325_
	);
	LUT2 #(
		.INIT('h8)
	) name6814 (
		\wishbone_bd_ram_mem3_reg[109][25]/P0001 ,
		_w12888_,
		_w17326_
	);
	LUT2 #(
		.INIT('h8)
	) name6815 (
		\wishbone_bd_ram_mem3_reg[195][25]/P0001 ,
		_w13144_,
		_w17327_
	);
	LUT2 #(
		.INIT('h8)
	) name6816 (
		\wishbone_bd_ram_mem3_reg[251][25]/P0001 ,
		_w13054_,
		_w17328_
	);
	LUT2 #(
		.INIT('h8)
	) name6817 (
		\wishbone_bd_ram_mem3_reg[159][25]/P0001 ,
		_w12774_,
		_w17329_
	);
	LUT2 #(
		.INIT('h8)
	) name6818 (
		\wishbone_bd_ram_mem3_reg[199][25]/P0001 ,
		_w12768_,
		_w17330_
	);
	LUT2 #(
		.INIT('h8)
	) name6819 (
		\wishbone_bd_ram_mem3_reg[63][25]/P0001 ,
		_w12850_,
		_w17331_
	);
	LUT2 #(
		.INIT('h8)
	) name6820 (
		\wishbone_bd_ram_mem3_reg[201][25]/P0001 ,
		_w12822_,
		_w17332_
	);
	LUT2 #(
		.INIT('h8)
	) name6821 (
		\wishbone_bd_ram_mem3_reg[76][25]/P0001 ,
		_w13184_,
		_w17333_
	);
	LUT2 #(
		.INIT('h8)
	) name6822 (
		\wishbone_bd_ram_mem3_reg[134][25]/P0001 ,
		_w12763_,
		_w17334_
	);
	LUT2 #(
		.INIT('h8)
	) name6823 (
		\wishbone_bd_ram_mem3_reg[43][25]/P0001 ,
		_w13200_,
		_w17335_
	);
	LUT2 #(
		.INIT('h8)
	) name6824 (
		\wishbone_bd_ram_mem3_reg[48][25]/P0001 ,
		_w12970_,
		_w17336_
	);
	LUT2 #(
		.INIT('h8)
	) name6825 (
		\wishbone_bd_ram_mem3_reg[75][25]/P0001 ,
		_w12826_,
		_w17337_
	);
	LUT2 #(
		.INIT('h8)
	) name6826 (
		\wishbone_bd_ram_mem3_reg[142][25]/P0001 ,
		_w12928_,
		_w17338_
	);
	LUT2 #(
		.INIT('h8)
	) name6827 (
		\wishbone_bd_ram_mem3_reg[236][25]/P0001 ,
		_w12731_,
		_w17339_
	);
	LUT2 #(
		.INIT('h8)
	) name6828 (
		\wishbone_bd_ram_mem3_reg[238][25]/P0001 ,
		_w13160_,
		_w17340_
	);
	LUT2 #(
		.INIT('h8)
	) name6829 (
		\wishbone_bd_ram_mem3_reg[174][25]/P0001 ,
		_w12972_,
		_w17341_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		\wishbone_bd_ram_mem3_reg[62][25]/P0001 ,
		_w12673_,
		_w17342_
	);
	LUT2 #(
		.INIT('h8)
	) name6831 (
		\wishbone_bd_ram_mem3_reg[224][25]/P0001 ,
		_w12902_,
		_w17343_
	);
	LUT2 #(
		.INIT('h8)
	) name6832 (
		\wishbone_bd_ram_mem3_reg[35][25]/P0001 ,
		_w12703_,
		_w17344_
	);
	LUT2 #(
		.INIT('h8)
	) name6833 (
		\wishbone_bd_ram_mem3_reg[31][25]/P0001 ,
		_w13198_,
		_w17345_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		\wishbone_bd_ram_mem3_reg[187][25]/P0001 ,
		_w13196_,
		_w17346_
	);
	LUT2 #(
		.INIT('h8)
	) name6835 (
		\wishbone_bd_ram_mem3_reg[161][25]/P0001 ,
		_w12754_,
		_w17347_
	);
	LUT2 #(
		.INIT('h8)
	) name6836 (
		\wishbone_bd_ram_mem3_reg[184][25]/P0001 ,
		_w13062_,
		_w17348_
	);
	LUT2 #(
		.INIT('h8)
	) name6837 (
		\wishbone_bd_ram_mem3_reg[89][25]/P0001 ,
		_w12964_,
		_w17349_
	);
	LUT2 #(
		.INIT('h8)
	) name6838 (
		\wishbone_bd_ram_mem3_reg[26][25]/P0001 ,
		_w12699_,
		_w17350_
	);
	LUT2 #(
		.INIT('h8)
	) name6839 (
		\wishbone_bd_ram_mem3_reg[225][25]/P0001 ,
		_w13092_,
		_w17351_
	);
	LUT2 #(
		.INIT('h8)
	) name6840 (
		\wishbone_bd_ram_mem3_reg[22][25]/P0001 ,
		_w13110_,
		_w17352_
	);
	LUT2 #(
		.INIT('h8)
	) name6841 (
		\wishbone_bd_ram_mem3_reg[203][25]/P0001 ,
		_w13158_,
		_w17353_
	);
	LUT2 #(
		.INIT('h8)
	) name6842 (
		\wishbone_bd_ram_mem3_reg[209][25]/P0001 ,
		_w13152_,
		_w17354_
	);
	LUT2 #(
		.INIT('h8)
	) name6843 (
		\wishbone_bd_ram_mem3_reg[192][25]/P0001 ,
		_w12938_,
		_w17355_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		\wishbone_bd_ram_mem3_reg[215][25]/P0001 ,
		_w12974_,
		_w17356_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		\wishbone_bd_ram_mem3_reg[137][25]/P0001 ,
		_w13168_,
		_w17357_
	);
	LUT2 #(
		.INIT('h8)
	) name6846 (
		\wishbone_bd_ram_mem3_reg[117][25]/P0001 ,
		_w12715_,
		_w17358_
	);
	LUT2 #(
		.INIT('h8)
	) name6847 (
		\wishbone_bd_ram_mem3_reg[240][25]/P0001 ,
		_w12864_,
		_w17359_
	);
	LUT2 #(
		.INIT('h8)
	) name6848 (
		\wishbone_bd_ram_mem3_reg[84][25]/P0001 ,
		_w12934_,
		_w17360_
	);
	LUT2 #(
		.INIT('h8)
	) name6849 (
		\wishbone_bd_ram_mem3_reg[198][25]/P0001 ,
		_w12832_,
		_w17361_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		\wishbone_bd_ram_mem3_reg[197][25]/P0001 ,
		_w12834_,
		_w17362_
	);
	LUT2 #(
		.INIT('h8)
	) name6851 (
		\wishbone_bd_ram_mem3_reg[213][25]/P0001 ,
		_w13002_,
		_w17363_
	);
	LUT2 #(
		.INIT('h8)
	) name6852 (
		\wishbone_bd_ram_mem3_reg[90][25]/P0001 ,
		_w12978_,
		_w17364_
	);
	LUT2 #(
		.INIT('h8)
	) name6853 (
		\wishbone_bd_ram_mem3_reg[110][25]/P0001 ,
		_w13046_,
		_w17365_
	);
	LUT2 #(
		.INIT('h8)
	) name6854 (
		\wishbone_bd_ram_mem3_reg[243][25]/P0001 ,
		_w12804_,
		_w17366_
	);
	LUT2 #(
		.INIT('h8)
	) name6855 (
		\wishbone_bd_ram_mem3_reg[61][25]/P0001 ,
		_w12725_,
		_w17367_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		\wishbone_bd_ram_mem3_reg[98][25]/P0001 ,
		_w12816_,
		_w17368_
	);
	LUT2 #(
		.INIT('h8)
	) name6857 (
		\wishbone_bd_ram_mem3_reg[79][25]/P0001 ,
		_w13212_,
		_w17369_
	);
	LUT2 #(
		.INIT('h8)
	) name6858 (
		\wishbone_bd_ram_mem3_reg[202][25]/P0001 ,
		_w12870_,
		_w17370_
	);
	LUT2 #(
		.INIT('h8)
	) name6859 (
		\wishbone_bd_ram_mem3_reg[1][25]/P0001 ,
		_w13014_,
		_w17371_
	);
	LUT2 #(
		.INIT('h8)
	) name6860 (
		\wishbone_bd_ram_mem3_reg[220][25]/P0001 ,
		_w13066_,
		_w17372_
	);
	LUT2 #(
		.INIT('h8)
	) name6861 (
		\wishbone_bd_ram_mem3_reg[64][25]/P0001 ,
		_w12976_,
		_w17373_
	);
	LUT2 #(
		.INIT('h8)
	) name6862 (
		\wishbone_bd_ram_mem3_reg[190][25]/P0001 ,
		_w12858_,
		_w17374_
	);
	LUT2 #(
		.INIT('h8)
	) name6863 (
		\wishbone_bd_ram_mem3_reg[153][25]/P0001 ,
		_w12890_,
		_w17375_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		\wishbone_bd_ram_mem3_reg[94][25]/P0001 ,
		_w13186_,
		_w17376_
	);
	LUT2 #(
		.INIT('h8)
	) name6865 (
		\wishbone_bd_ram_mem3_reg[122][25]/P0001 ,
		_w13130_,
		_w17377_
	);
	LUT2 #(
		.INIT('h8)
	) name6866 (
		\wishbone_bd_ram_mem3_reg[144][25]/P0001 ,
		_w12756_,
		_w17378_
	);
	LUT2 #(
		.INIT('h8)
	) name6867 (
		\wishbone_bd_ram_mem3_reg[222][25]/P0001 ,
		_w13094_,
		_w17379_
	);
	LUT2 #(
		.INIT('h8)
	) name6868 (
		\wishbone_bd_ram_mem3_reg[172][25]/P0001 ,
		_w12944_,
		_w17380_
	);
	LUT2 #(
		.INIT('h8)
	) name6869 (
		\wishbone_bd_ram_mem3_reg[85][25]/P0001 ,
		_w13216_,
		_w17381_
	);
	LUT2 #(
		.INIT('h8)
	) name6870 (
		\wishbone_bd_ram_mem3_reg[242][25]/P0001 ,
		_w12932_,
		_w17382_
	);
	LUT2 #(
		.INIT('h8)
	) name6871 (
		\wishbone_bd_ram_mem3_reg[157][25]/P0001 ,
		_w12926_,
		_w17383_
	);
	LUT2 #(
		.INIT('h8)
	) name6872 (
		\wishbone_bd_ram_mem3_reg[183][25]/P0001 ,
		_w12787_,
		_w17384_
	);
	LUT2 #(
		.INIT('h8)
	) name6873 (
		\wishbone_bd_ram_mem3_reg[24][25]/P0001 ,
		_w13084_,
		_w17385_
	);
	LUT2 #(
		.INIT('h8)
	) name6874 (
		\wishbone_bd_ram_mem3_reg[51][25]/P0001 ,
		_w13024_,
		_w17386_
	);
	LUT2 #(
		.INIT('h8)
	) name6875 (
		\wishbone_bd_ram_mem3_reg[234][25]/P0001 ,
		_w13214_,
		_w17387_
	);
	LUT2 #(
		.INIT('h8)
	) name6876 (
		\wishbone_bd_ram_mem3_reg[105][25]/P0001 ,
		_w12751_,
		_w17388_
	);
	LUT2 #(
		.INIT('h8)
	) name6877 (
		\wishbone_bd_ram_mem3_reg[253][25]/P0001 ,
		_w13100_,
		_w17389_
	);
	LUT2 #(
		.INIT('h8)
	) name6878 (
		\wishbone_bd_ram_mem3_reg[108][25]/P0001 ,
		_w13156_,
		_w17390_
	);
	LUT2 #(
		.INIT('h8)
	) name6879 (
		\wishbone_bd_ram_mem3_reg[217][25]/P0001 ,
		_w13188_,
		_w17391_
	);
	LUT2 #(
		.INIT('h8)
	) name6880 (
		\wishbone_bd_ram_mem3_reg[140][25]/P0001 ,
		_w12894_,
		_w17392_
	);
	LUT2 #(
		.INIT('h8)
	) name6881 (
		\wishbone_bd_ram_mem3_reg[34][25]/P0001 ,
		_w12930_,
		_w17393_
	);
	LUT2 #(
		.INIT('h8)
	) name6882 (
		\wishbone_bd_ram_mem3_reg[93][25]/P0001 ,
		_w13016_,
		_w17394_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		\wishbone_bd_ram_mem3_reg[100][25]/P0001 ,
		_w12960_,
		_w17395_
	);
	LUT2 #(
		.INIT('h8)
	) name6884 (
		\wishbone_bd_ram_mem3_reg[60][25]/P0001 ,
		_w13204_,
		_w17396_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		\wishbone_bd_ram_mem3_reg[39][25]/P0001 ,
		_w13018_,
		_w17397_
	);
	LUT2 #(
		.INIT('h8)
	) name6886 (
		\wishbone_bd_ram_mem3_reg[166][25]/P0001 ,
		_w13040_,
		_w17398_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		\wishbone_bd_ram_mem3_reg[59][25]/P0001 ,
		_w12780_,
		_w17399_
	);
	LUT2 #(
		.INIT('h8)
	) name6888 (
		\wishbone_bd_ram_mem3_reg[128][25]/P0001 ,
		_w12793_,
		_w17400_
	);
	LUT2 #(
		.INIT('h8)
	) name6889 (
		\wishbone_bd_ram_mem3_reg[47][25]/P0001 ,
		_w12904_,
		_w17401_
	);
	LUT2 #(
		.INIT('h8)
	) name6890 (
		\wishbone_bd_ram_mem3_reg[177][25]/P0001 ,
		_w12996_,
		_w17402_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		\wishbone_bd_ram_mem3_reg[36][25]/P0001 ,
		_w12800_,
		_w17403_
	);
	LUT2 #(
		.INIT('h8)
	) name6892 (
		\wishbone_bd_ram_mem3_reg[55][25]/P0001 ,
		_w12785_,
		_w17404_
	);
	LUT2 #(
		.INIT('h8)
	) name6893 (
		\wishbone_bd_ram_mem3_reg[106][25]/P0001 ,
		_w12713_,
		_w17405_
	);
	LUT2 #(
		.INIT('h8)
	) name6894 (
		\wishbone_bd_ram_mem3_reg[143][25]/P0001 ,
		_w12922_,
		_w17406_
	);
	LUT2 #(
		.INIT('h8)
	) name6895 (
		\wishbone_bd_ram_mem3_reg[176][25]/P0001 ,
		_w12868_,
		_w17407_
	);
	LUT2 #(
		.INIT('h8)
	) name6896 (
		\wishbone_bd_ram_mem3_reg[3][25]/P0001 ,
		_w12866_,
		_w17408_
	);
	LUT2 #(
		.INIT('h8)
	) name6897 (
		\wishbone_bd_ram_mem3_reg[81][25]/P0001 ,
		_w12950_,
		_w17409_
	);
	LUT2 #(
		.INIT('h8)
	) name6898 (
		\wishbone_bd_ram_mem3_reg[77][25]/P0001 ,
		_w12982_,
		_w17410_
	);
	LUT2 #(
		.INIT('h8)
	) name6899 (
		\wishbone_bd_ram_mem3_reg[211][25]/P0001 ,
		_w13166_,
		_w17411_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		\wishbone_bd_ram_mem3_reg[149][25]/P0001 ,
		_w12741_,
		_w17412_
	);
	LUT2 #(
		.INIT('h8)
	) name6901 (
		\wishbone_bd_ram_mem3_reg[227][25]/P0001 ,
		_w12936_,
		_w17413_
	);
	LUT2 #(
		.INIT('h8)
	) name6902 (
		\wishbone_bd_ram_mem3_reg[96][25]/P0001 ,
		_w12912_,
		_w17414_
	);
	LUT2 #(
		.INIT('h8)
	) name6903 (
		\wishbone_bd_ram_mem3_reg[127][25]/P0001 ,
		_w13164_,
		_w17415_
	);
	LUT2 #(
		.INIT('h8)
	) name6904 (
		\wishbone_bd_ram_mem3_reg[101][25]/P0001 ,
		_w13192_,
		_w17416_
	);
	LUT2 #(
		.INIT('h8)
	) name6905 (
		\wishbone_bd_ram_mem3_reg[154][25]/P0001 ,
		_w12962_,
		_w17417_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		\wishbone_bd_ram_mem3_reg[50][25]/P0001 ,
		_w13150_,
		_w17418_
	);
	LUT2 #(
		.INIT('h8)
	) name6907 (
		\wishbone_bd_ram_mem3_reg[165][25]/P0001 ,
		_w13044_,
		_w17419_
	);
	LUT2 #(
		.INIT('h8)
	) name6908 (
		\wishbone_bd_ram_mem3_reg[252][25]/P0001 ,
		_w13080_,
		_w17420_
	);
	LUT2 #(
		.INIT('h8)
	) name6909 (
		\wishbone_bd_ram_mem3_reg[29][25]/P0001 ,
		_w12952_,
		_w17421_
	);
	LUT2 #(
		.INIT('h8)
	) name6910 (
		\wishbone_bd_ram_mem3_reg[205][25]/P0001 ,
		_w13068_,
		_w17422_
	);
	LUT2 #(
		.INIT('h8)
	) name6911 (
		\wishbone_bd_ram_mem3_reg[52][25]/P0001 ,
		_w13082_,
		_w17423_
	);
	LUT2 #(
		.INIT('h8)
	) name6912 (
		\wishbone_bd_ram_mem3_reg[196][25]/P0001 ,
		_w13090_,
		_w17424_
	);
	LUT2 #(
		.INIT('h8)
	) name6913 (
		\wishbone_bd_ram_mem3_reg[74][25]/P0001 ,
		_w12812_,
		_w17425_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		\wishbone_bd_ram_mem3_reg[112][25]/P0001 ,
		_w12733_,
		_w17426_
	);
	LUT2 #(
		.INIT('h8)
	) name6915 (
		\wishbone_bd_ram_mem3_reg[125][25]/P0001 ,
		_w12956_,
		_w17427_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		\wishbone_bd_ram_mem3_reg[44][25]/P0001 ,
		_w12896_,
		_w17428_
	);
	LUT2 #(
		.INIT('h8)
	) name6917 (
		\wishbone_bd_ram_mem3_reg[70][25]/P0001 ,
		_w12840_,
		_w17429_
	);
	LUT2 #(
		.INIT('h8)
	) name6918 (
		\wishbone_bd_ram_mem3_reg[206][25]/P0001 ,
		_w12954_,
		_w17430_
	);
	LUT2 #(
		.INIT('h8)
	) name6919 (
		\wishbone_bd_ram_mem3_reg[145][25]/P0001 ,
		_w13106_,
		_w17431_
	);
	LUT2 #(
		.INIT('h8)
	) name6920 (
		\wishbone_bd_ram_mem3_reg[11][25]/P0001 ,
		_w13194_,
		_w17432_
	);
	LUT2 #(
		.INIT('h8)
	) name6921 (
		\wishbone_bd_ram_mem3_reg[21][25]/P0001 ,
		_w12906_,
		_w17433_
	);
	LUT2 #(
		.INIT('h8)
	) name6922 (
		\wishbone_bd_ram_mem3_reg[121][25]/P0001 ,
		_w13078_,
		_w17434_
	);
	LUT2 #(
		.INIT('h8)
	) name6923 (
		\wishbone_bd_ram_mem3_reg[4][25]/P0001 ,
		_w12666_,
		_w17435_
	);
	LUT2 #(
		.INIT('h8)
	) name6924 (
		\wishbone_bd_ram_mem3_reg[33][25]/P0001 ,
		_w12980_,
		_w17436_
	);
	LUT2 #(
		.INIT('h8)
	) name6925 (
		\wishbone_bd_ram_mem3_reg[221][25]/P0001 ,
		_w12802_,
		_w17437_
	);
	LUT2 #(
		.INIT('h8)
	) name6926 (
		\wishbone_bd_ram_mem3_reg[168][25]/P0001 ,
		_w13208_,
		_w17438_
	);
	LUT2 #(
		.INIT('h8)
	) name6927 (
		\wishbone_bd_ram_mem3_reg[170][25]/P0001 ,
		_w13030_,
		_w17439_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		\wishbone_bd_ram_mem3_reg[71][25]/P0001 ,
		_w12798_,
		_w17440_
	);
	LUT2 #(
		.INIT('h8)
	) name6929 (
		\wishbone_bd_ram_mem3_reg[186][25]/P0001 ,
		_w12783_,
		_w17441_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		\wishbone_bd_ram_mem3_reg[37][25]/P0001 ,
		_w13102_,
		_w17442_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		\wishbone_bd_ram_mem3_reg[80][25]/P0001 ,
		_w12689_,
		_w17443_
	);
	LUT2 #(
		.INIT('h8)
	) name6932 (
		\wishbone_bd_ram_mem3_reg[116][25]/P0001 ,
		_w12998_,
		_w17444_
	);
	LUT2 #(
		.INIT('h8)
	) name6933 (
		\wishbone_bd_ram_mem3_reg[131][25]/P0001 ,
		_w12852_,
		_w17445_
	);
	LUT2 #(
		.INIT('h8)
	) name6934 (
		\wishbone_bd_ram_mem3_reg[249][25]/P0001 ,
		_w12900_,
		_w17446_
	);
	LUT2 #(
		.INIT('h8)
	) name6935 (
		\wishbone_bd_ram_mem3_reg[78][25]/P0001 ,
		_w12874_,
		_w17447_
	);
	LUT2 #(
		.INIT('h8)
	) name6936 (
		\wishbone_bd_ram_mem3_reg[162][25]/P0001 ,
		_w13098_,
		_w17448_
	);
	LUT2 #(
		.INIT('h8)
	) name6937 (
		\wishbone_bd_ram_mem3_reg[138][25]/P0001 ,
		_w12958_,
		_w17449_
	);
	LUT2 #(
		.INIT('h8)
	) name6938 (
		\wishbone_bd_ram_mem3_reg[41][25]/P0001 ,
		_w13052_,
		_w17450_
	);
	LUT2 #(
		.INIT('h8)
	) name6939 (
		\wishbone_bd_ram_mem3_reg[73][25]/P0001 ,
		_w12918_,
		_w17451_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		\wishbone_bd_ram_mem3_reg[58][25]/P0001 ,
		_w13070_,
		_w17452_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		\wishbone_bd_ram_mem3_reg[7][25]/P0001 ,
		_w12728_,
		_w17453_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		\wishbone_bd_ram_mem3_reg[151][25]/P0001 ,
		_w13142_,
		_w17454_
	);
	LUT2 #(
		.INIT('h8)
	) name6943 (
		\wishbone_bd_ram_mem3_reg[147][25]/P0001 ,
		_w13146_,
		_w17455_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		\wishbone_bd_ram_mem3_reg[133][25]/P0001 ,
		_w12761_,
		_w17456_
	);
	LUT2 #(
		.INIT('h8)
	) name6945 (
		\wishbone_bd_ram_mem3_reg[97][25]/P0001 ,
		_w13096_,
		_w17457_
	);
	LUT2 #(
		.INIT('h8)
	) name6946 (
		\wishbone_bd_ram_mem3_reg[114][25]/P0001 ,
		_w13202_,
		_w17458_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		\wishbone_bd_ram_mem3_reg[250][25]/P0001 ,
		_w13128_,
		_w17459_
	);
	LUT2 #(
		.INIT('h8)
	) name6948 (
		\wishbone_bd_ram_mem3_reg[244][25]/P0001 ,
		_w12747_,
		_w17460_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		\wishbone_bd_ram_mem3_reg[232][25]/P0001 ,
		_w12758_,
		_w17461_
	);
	LUT2 #(
		.INIT('h8)
	) name6950 (
		\wishbone_bd_ram_mem3_reg[175][25]/P0001 ,
		_w13126_,
		_w17462_
	);
	LUT2 #(
		.INIT('h8)
	) name6951 (
		\wishbone_bd_ram_mem3_reg[42][25]/P0001 ,
		_w12842_,
		_w17463_
	);
	LUT2 #(
		.INIT('h8)
	) name6952 (
		\wishbone_bd_ram_mem3_reg[163][25]/P0001 ,
		_w12882_,
		_w17464_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		\wishbone_bd_ram_mem3_reg[231][25]/P0001 ,
		_w12856_,
		_w17465_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		\wishbone_bd_ram_mem3_reg[16][25]/P0001 ,
		_w13140_,
		_w17466_
	);
	LUT2 #(
		.INIT('h8)
	) name6955 (
		\wishbone_bd_ram_mem3_reg[218][25]/P0001 ,
		_w13206_,
		_w17467_
	);
	LUT2 #(
		.INIT('h8)
	) name6956 (
		\wishbone_bd_ram_mem3_reg[111][25]/P0001 ,
		_w12744_,
		_w17468_
	);
	LUT2 #(
		.INIT('h8)
	) name6957 (
		\wishbone_bd_ram_mem3_reg[189][25]/P0001 ,
		_w13042_,
		_w17469_
	);
	LUT2 #(
		.INIT('h8)
	) name6958 (
		\wishbone_bd_ram_mem3_reg[191][25]/P0001 ,
		_w13034_,
		_w17470_
	);
	LUT2 #(
		.INIT('h8)
	) name6959 (
		\wishbone_bd_ram_mem3_reg[32][25]/P0001 ,
		_w13120_,
		_w17471_
	);
	LUT2 #(
		.INIT('h8)
	) name6960 (
		\wishbone_bd_ram_mem3_reg[194][25]/P0001 ,
		_w12772_,
		_w17472_
	);
	LUT2 #(
		.INIT('h8)
	) name6961 (
		\wishbone_bd_ram_mem3_reg[241][25]/P0001 ,
		_w13006_,
		_w17473_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		\wishbone_bd_ram_mem3_reg[53][25]/P0001 ,
		_w13020_,
		_w17474_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		\wishbone_bd_ram_mem3_reg[72][25]/P0001 ,
		_w12810_,
		_w17475_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		\wishbone_bd_ram_mem3_reg[182][25]/P0001 ,
		_w12820_,
		_w17476_
	);
	LUT2 #(
		.INIT('h8)
	) name6965 (
		\wishbone_bd_ram_mem3_reg[136][25]/P0001 ,
		_w13064_,
		_w17477_
	);
	LUT2 #(
		.INIT('h8)
	) name6966 (
		\wishbone_bd_ram_mem3_reg[185][25]/P0001 ,
		_w12940_,
		_w17478_
	);
	LUT2 #(
		.INIT('h8)
	) name6967 (
		\wishbone_bd_ram_mem3_reg[247][25]/P0001 ,
		_w12818_,
		_w17479_
	);
	LUT2 #(
		.INIT('h8)
	) name6968 (
		\wishbone_bd_ram_mem3_reg[103][25]/P0001 ,
		_w12846_,
		_w17480_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		\wishbone_bd_ram_mem3_reg[223][25]/P0001 ,
		_w12838_,
		_w17481_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		\wishbone_bd_ram_mem3_reg[228][25]/P0001 ,
		_w12765_,
		_w17482_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		\wishbone_bd_ram_mem3_reg[254][25]/P0001 ,
		_w12892_,
		_w17483_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		\wishbone_bd_ram_mem3_reg[146][25]/P0001 ,
		_w13060_,
		_w17484_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		\wishbone_bd_ram_mem3_reg[233][25]/P0001 ,
		_w12836_,
		_w17485_
	);
	LUT2 #(
		.INIT('h8)
	) name6974 (
		\wishbone_bd_ram_mem3_reg[69][25]/P0001 ,
		_w12738_,
		_w17486_
	);
	LUT2 #(
		.INIT('h8)
	) name6975 (
		\wishbone_bd_ram_mem3_reg[8][25]/P0001 ,
		_w12920_,
		_w17487_
	);
	LUT2 #(
		.INIT('h8)
	) name6976 (
		\wishbone_bd_ram_mem3_reg[219][25]/P0001 ,
		_w12806_,
		_w17488_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		\wishbone_bd_ram_mem3_reg[180][25]/P0001 ,
		_w12791_,
		_w17489_
	);
	LUT2 #(
		.INIT('h8)
	) name6978 (
		\wishbone_bd_ram_mem3_reg[23][25]/P0001 ,
		_w13008_,
		_w17490_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		\wishbone_bd_ram_mem3_reg[239][25]/P0001 ,
		_w12862_,
		_w17491_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		\wishbone_bd_ram_mem3_reg[46][25]/P0001 ,
		_w12884_,
		_w17492_
	);
	LUT2 #(
		.INIT('h8)
	) name6981 (
		\wishbone_bd_ram_mem3_reg[99][25]/P0001 ,
		_w13038_,
		_w17493_
	);
	LUT2 #(
		.INIT('h8)
	) name6982 (
		\wishbone_bd_ram_mem3_reg[54][25]/P0001 ,
		_w12770_,
		_w17494_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		\wishbone_bd_ram_mem3_reg[208][25]/P0001 ,
		_w13032_,
		_w17495_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		\wishbone_bd_ram_mem3_reg[66][25]/P0001 ,
		_w12824_,
		_w17496_
	);
	LUT2 #(
		.INIT('h8)
	) name6985 (
		\wishbone_bd_ram_mem3_reg[30][25]/P0001 ,
		_w13104_,
		_w17497_
	);
	LUT2 #(
		.INIT('h8)
	) name6986 (
		\wishbone_bd_ram_mem3_reg[40][25]/P0001 ,
		_w13132_,
		_w17498_
	);
	LUT2 #(
		.INIT('h8)
	) name6987 (
		\wishbone_bd_ram_mem3_reg[83][25]/P0001 ,
		_w12916_,
		_w17499_
	);
	LUT2 #(
		.INIT('h8)
	) name6988 (
		\wishbone_bd_ram_mem3_reg[139][25]/P0001 ,
		_w12814_,
		_w17500_
	);
	LUT2 #(
		.INIT('h8)
	) name6989 (
		\wishbone_bd_ram_mem3_reg[115][25]/P0001 ,
		_w13112_,
		_w17501_
	);
	LUT2 #(
		.INIT('h8)
	) name6990 (
		\wishbone_bd_ram_mem3_reg[158][25]/P0001 ,
		_w12898_,
		_w17502_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		\wishbone_bd_ram_mem3_reg[9][25]/P0001 ,
		_w12808_,
		_w17503_
	);
	LUT2 #(
		.INIT('h8)
	) name6992 (
		\wishbone_bd_ram_mem3_reg[65][25]/P0001 ,
		_w13176_,
		_w17504_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		\wishbone_bd_ram_mem3_reg[25][25]/P0001 ,
		_w13108_,
		_w17505_
	);
	LUT2 #(
		.INIT('h8)
	) name6994 (
		\wishbone_bd_ram_mem3_reg[6][25]/P0001 ,
		_w12968_,
		_w17506_
	);
	LUT2 #(
		.INIT('h8)
	) name6995 (
		\wishbone_bd_ram_mem3_reg[135][25]/P0001 ,
		_w13124_,
		_w17507_
	);
	LUT2 #(
		.INIT('h8)
	) name6996 (
		\wishbone_bd_ram_mem3_reg[2][25]/P0001 ,
		_w13088_,
		_w17508_
	);
	LUT2 #(
		.INIT('h8)
	) name6997 (
		\wishbone_bd_ram_mem3_reg[248][25]/P0001 ,
		_w12789_,
		_w17509_
	);
	LUT2 #(
		.INIT('h8)
	) name6998 (
		\wishbone_bd_ram_mem3_reg[87][25]/P0001 ,
		_w13154_,
		_w17510_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		\wishbone_bd_ram_mem3_reg[171][25]/P0001 ,
		_w12910_,
		_w17511_
	);
	LUT2 #(
		.INIT('h8)
	) name7000 (
		\wishbone_bd_ram_mem3_reg[255][25]/P0001 ,
		_w13072_,
		_w17512_
	);
	LUT2 #(
		.INIT('h8)
	) name7001 (
		\wishbone_bd_ram_mem3_reg[45][25]/P0001 ,
		_w12908_,
		_w17513_
	);
	LUT2 #(
		.INIT('h8)
	) name7002 (
		\wishbone_bd_ram_mem3_reg[226][25]/P0001 ,
		_w13138_,
		_w17514_
	);
	LUT2 #(
		.INIT('h8)
	) name7003 (
		\wishbone_bd_ram_mem3_reg[119][25]/P0001 ,
		_w13048_,
		_w17515_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		\wishbone_bd_ram_mem3_reg[88][25]/P0001 ,
		_w12860_,
		_w17516_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		\wishbone_bd_ram_mem3_reg[82][25]/P0001 ,
		_w12942_,
		_w17517_
	);
	LUT2 #(
		.INIT('h8)
	) name7006 (
		\wishbone_bd_ram_mem3_reg[155][25]/P0001 ,
		_w13122_,
		_w17518_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		\wishbone_bd_ram_mem3_reg[148][25]/P0001 ,
		_w13000_,
		_w17519_
	);
	LUT2 #(
		.INIT('h8)
	) name7008 (
		\wishbone_bd_ram_mem3_reg[95][25]/P0001 ,
		_w12844_,
		_w17520_
	);
	LUT2 #(
		.INIT('h8)
	) name7009 (
		\wishbone_bd_ram_mem3_reg[113][25]/P0001 ,
		_w13026_,
		_w17521_
	);
	LUT2 #(
		.INIT('h8)
	) name7010 (
		\wishbone_bd_ram_mem3_reg[150][25]/P0001 ,
		_w13136_,
		_w17522_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		\wishbone_bd_ram_mem3_reg[102][25]/P0001 ,
		_w12685_,
		_w17523_
	);
	LUT2 #(
		.INIT('h8)
	) name7012 (
		\wishbone_bd_ram_mem3_reg[173][25]/P0001 ,
		_w12854_,
		_w17524_
	);
	LUT2 #(
		.INIT('h8)
	) name7013 (
		\wishbone_bd_ram_mem3_reg[216][25]/P0001 ,
		_w13028_,
		_w17525_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		\wishbone_bd_ram_mem3_reg[246][25]/P0001 ,
		_w13076_,
		_w17526_
	);
	LUT2 #(
		.INIT('h8)
	) name7015 (
		\wishbone_bd_ram_mem3_reg[104][25]/P0001 ,
		_w13148_,
		_w17527_
	);
	LUT2 #(
		.INIT('h8)
	) name7016 (
		\wishbone_bd_ram_mem3_reg[212][25]/P0001 ,
		_w12796_,
		_w17528_
	);
	LUT2 #(
		.INIT('h8)
	) name7017 (
		\wishbone_bd_ram_mem3_reg[92][25]/P0001 ,
		_w13010_,
		_w17529_
	);
	LUT2 #(
		.INIT('h8)
	) name7018 (
		\wishbone_bd_ram_mem3_reg[91][25]/P0001 ,
		_w13074_,
		_w17530_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		\wishbone_bd_ram_mem3_reg[188][25]/P0001 ,
		_w12948_,
		_w17531_
	);
	LUT2 #(
		.INIT('h8)
	) name7020 (
		\wishbone_bd_ram_mem3_reg[107][25]/P0001 ,
		_w12749_,
		_w17532_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		\wishbone_bd_ram_mem3_reg[18][25]/P0001 ,
		_w12679_,
		_w17533_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		\wishbone_bd_ram_mem3_reg[120][25]/P0001 ,
		_w12707_,
		_w17534_
	);
	LUT2 #(
		.INIT('h8)
	) name7023 (
		\wishbone_bd_ram_mem3_reg[245][25]/P0001 ,
		_w13022_,
		_w17535_
	);
	LUT2 #(
		.INIT('h8)
	) name7024 (
		\wishbone_bd_ram_mem3_reg[56][25]/P0001 ,
		_w12778_,
		_w17536_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		\wishbone_bd_ram_mem3_reg[15][25]/P0001 ,
		_w13210_,
		_w17537_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		\wishbone_bd_ram_mem3_reg[132][25]/P0001 ,
		_w12992_,
		_w17538_
	);
	LUT2 #(
		.INIT('h8)
	) name7027 (
		\wishbone_bd_ram_mem3_reg[181][25]/P0001 ,
		_w12828_,
		_w17539_
	);
	LUT2 #(
		.INIT('h8)
	) name7028 (
		\wishbone_bd_ram_mem3_reg[193][25]/P0001 ,
		_w13056_,
		_w17540_
	);
	LUT2 #(
		.INIT('h8)
	) name7029 (
		\wishbone_bd_ram_mem3_reg[28][25]/P0001 ,
		_w13170_,
		_w17541_
	);
	LUT2 #(
		.INIT('h8)
	) name7030 (
		\wishbone_bd_ram_mem3_reg[210][25]/P0001 ,
		_w12924_,
		_w17542_
	);
	LUT2 #(
		.INIT('h8)
	) name7031 (
		\wishbone_bd_ram_mem3_reg[178][25]/P0001 ,
		_w12886_,
		_w17543_
	);
	LUT2 #(
		.INIT('h8)
	) name7032 (
		\wishbone_bd_ram_mem3_reg[14][25]/P0001 ,
		_w13086_,
		_w17544_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		\wishbone_bd_ram_mem3_reg[204][25]/P0001 ,
		_w13162_,
		_w17545_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		\wishbone_bd_ram_mem3_reg[118][25]/P0001 ,
		_w12830_,
		_w17546_
	);
	LUT2 #(
		.INIT('h8)
	) name7035 (
		\wishbone_bd_ram_mem3_reg[67][25]/P0001 ,
		_w13134_,
		_w17547_
	);
	LUT2 #(
		.INIT('h8)
	) name7036 (
		\wishbone_bd_ram_mem3_reg[10][25]/P0001 ,
		_w13172_,
		_w17548_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		\wishbone_bd_ram_mem3_reg[123][25]/P0001 ,
		_w13114_,
		_w17549_
	);
	LUT2 #(
		.INIT('h8)
	) name7038 (
		\wishbone_bd_ram_mem3_reg[207][25]/P0001 ,
		_w13180_,
		_w17550_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		\wishbone_bd_ram_mem3_reg[27][25]/P0001 ,
		_w12880_,
		_w17551_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		\wishbone_bd_ram_mem3_reg[129][25]/P0001 ,
		_w12776_,
		_w17552_
	);
	LUT2 #(
		.INIT('h8)
	) name7041 (
		\wishbone_bd_ram_mem3_reg[20][25]/P0001 ,
		_w13174_,
		_w17553_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		\wishbone_bd_ram_mem3_reg[200][25]/P0001 ,
		_w12988_,
		_w17554_
	);
	LUT2 #(
		.INIT('h1)
	) name7043 (
		_w17299_,
		_w17300_,
		_w17555_
	);
	LUT2 #(
		.INIT('h1)
	) name7044 (
		_w17301_,
		_w17302_,
		_w17556_
	);
	LUT2 #(
		.INIT('h1)
	) name7045 (
		_w17303_,
		_w17304_,
		_w17557_
	);
	LUT2 #(
		.INIT('h1)
	) name7046 (
		_w17305_,
		_w17306_,
		_w17558_
	);
	LUT2 #(
		.INIT('h1)
	) name7047 (
		_w17307_,
		_w17308_,
		_w17559_
	);
	LUT2 #(
		.INIT('h1)
	) name7048 (
		_w17309_,
		_w17310_,
		_w17560_
	);
	LUT2 #(
		.INIT('h1)
	) name7049 (
		_w17311_,
		_w17312_,
		_w17561_
	);
	LUT2 #(
		.INIT('h1)
	) name7050 (
		_w17313_,
		_w17314_,
		_w17562_
	);
	LUT2 #(
		.INIT('h1)
	) name7051 (
		_w17315_,
		_w17316_,
		_w17563_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		_w17317_,
		_w17318_,
		_w17564_
	);
	LUT2 #(
		.INIT('h1)
	) name7053 (
		_w17319_,
		_w17320_,
		_w17565_
	);
	LUT2 #(
		.INIT('h1)
	) name7054 (
		_w17321_,
		_w17322_,
		_w17566_
	);
	LUT2 #(
		.INIT('h1)
	) name7055 (
		_w17323_,
		_w17324_,
		_w17567_
	);
	LUT2 #(
		.INIT('h1)
	) name7056 (
		_w17325_,
		_w17326_,
		_w17568_
	);
	LUT2 #(
		.INIT('h1)
	) name7057 (
		_w17327_,
		_w17328_,
		_w17569_
	);
	LUT2 #(
		.INIT('h1)
	) name7058 (
		_w17329_,
		_w17330_,
		_w17570_
	);
	LUT2 #(
		.INIT('h1)
	) name7059 (
		_w17331_,
		_w17332_,
		_w17571_
	);
	LUT2 #(
		.INIT('h1)
	) name7060 (
		_w17333_,
		_w17334_,
		_w17572_
	);
	LUT2 #(
		.INIT('h1)
	) name7061 (
		_w17335_,
		_w17336_,
		_w17573_
	);
	LUT2 #(
		.INIT('h1)
	) name7062 (
		_w17337_,
		_w17338_,
		_w17574_
	);
	LUT2 #(
		.INIT('h1)
	) name7063 (
		_w17339_,
		_w17340_,
		_w17575_
	);
	LUT2 #(
		.INIT('h1)
	) name7064 (
		_w17341_,
		_w17342_,
		_w17576_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w17343_,
		_w17344_,
		_w17577_
	);
	LUT2 #(
		.INIT('h1)
	) name7066 (
		_w17345_,
		_w17346_,
		_w17578_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		_w17347_,
		_w17348_,
		_w17579_
	);
	LUT2 #(
		.INIT('h1)
	) name7068 (
		_w17349_,
		_w17350_,
		_w17580_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w17351_,
		_w17352_,
		_w17581_
	);
	LUT2 #(
		.INIT('h1)
	) name7070 (
		_w17353_,
		_w17354_,
		_w17582_
	);
	LUT2 #(
		.INIT('h1)
	) name7071 (
		_w17355_,
		_w17356_,
		_w17583_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		_w17357_,
		_w17358_,
		_w17584_
	);
	LUT2 #(
		.INIT('h1)
	) name7073 (
		_w17359_,
		_w17360_,
		_w17585_
	);
	LUT2 #(
		.INIT('h1)
	) name7074 (
		_w17361_,
		_w17362_,
		_w17586_
	);
	LUT2 #(
		.INIT('h1)
	) name7075 (
		_w17363_,
		_w17364_,
		_w17587_
	);
	LUT2 #(
		.INIT('h1)
	) name7076 (
		_w17365_,
		_w17366_,
		_w17588_
	);
	LUT2 #(
		.INIT('h1)
	) name7077 (
		_w17367_,
		_w17368_,
		_w17589_
	);
	LUT2 #(
		.INIT('h1)
	) name7078 (
		_w17369_,
		_w17370_,
		_w17590_
	);
	LUT2 #(
		.INIT('h1)
	) name7079 (
		_w17371_,
		_w17372_,
		_w17591_
	);
	LUT2 #(
		.INIT('h1)
	) name7080 (
		_w17373_,
		_w17374_,
		_w17592_
	);
	LUT2 #(
		.INIT('h1)
	) name7081 (
		_w17375_,
		_w17376_,
		_w17593_
	);
	LUT2 #(
		.INIT('h1)
	) name7082 (
		_w17377_,
		_w17378_,
		_w17594_
	);
	LUT2 #(
		.INIT('h1)
	) name7083 (
		_w17379_,
		_w17380_,
		_w17595_
	);
	LUT2 #(
		.INIT('h1)
	) name7084 (
		_w17381_,
		_w17382_,
		_w17596_
	);
	LUT2 #(
		.INIT('h1)
	) name7085 (
		_w17383_,
		_w17384_,
		_w17597_
	);
	LUT2 #(
		.INIT('h1)
	) name7086 (
		_w17385_,
		_w17386_,
		_w17598_
	);
	LUT2 #(
		.INIT('h1)
	) name7087 (
		_w17387_,
		_w17388_,
		_w17599_
	);
	LUT2 #(
		.INIT('h1)
	) name7088 (
		_w17389_,
		_w17390_,
		_w17600_
	);
	LUT2 #(
		.INIT('h1)
	) name7089 (
		_w17391_,
		_w17392_,
		_w17601_
	);
	LUT2 #(
		.INIT('h1)
	) name7090 (
		_w17393_,
		_w17394_,
		_w17602_
	);
	LUT2 #(
		.INIT('h1)
	) name7091 (
		_w17395_,
		_w17396_,
		_w17603_
	);
	LUT2 #(
		.INIT('h1)
	) name7092 (
		_w17397_,
		_w17398_,
		_w17604_
	);
	LUT2 #(
		.INIT('h1)
	) name7093 (
		_w17399_,
		_w17400_,
		_w17605_
	);
	LUT2 #(
		.INIT('h1)
	) name7094 (
		_w17401_,
		_w17402_,
		_w17606_
	);
	LUT2 #(
		.INIT('h1)
	) name7095 (
		_w17403_,
		_w17404_,
		_w17607_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w17405_,
		_w17406_,
		_w17608_
	);
	LUT2 #(
		.INIT('h1)
	) name7097 (
		_w17407_,
		_w17408_,
		_w17609_
	);
	LUT2 #(
		.INIT('h1)
	) name7098 (
		_w17409_,
		_w17410_,
		_w17610_
	);
	LUT2 #(
		.INIT('h1)
	) name7099 (
		_w17411_,
		_w17412_,
		_w17611_
	);
	LUT2 #(
		.INIT('h1)
	) name7100 (
		_w17413_,
		_w17414_,
		_w17612_
	);
	LUT2 #(
		.INIT('h1)
	) name7101 (
		_w17415_,
		_w17416_,
		_w17613_
	);
	LUT2 #(
		.INIT('h1)
	) name7102 (
		_w17417_,
		_w17418_,
		_w17614_
	);
	LUT2 #(
		.INIT('h1)
	) name7103 (
		_w17419_,
		_w17420_,
		_w17615_
	);
	LUT2 #(
		.INIT('h1)
	) name7104 (
		_w17421_,
		_w17422_,
		_w17616_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w17423_,
		_w17424_,
		_w17617_
	);
	LUT2 #(
		.INIT('h1)
	) name7106 (
		_w17425_,
		_w17426_,
		_w17618_
	);
	LUT2 #(
		.INIT('h1)
	) name7107 (
		_w17427_,
		_w17428_,
		_w17619_
	);
	LUT2 #(
		.INIT('h1)
	) name7108 (
		_w17429_,
		_w17430_,
		_w17620_
	);
	LUT2 #(
		.INIT('h1)
	) name7109 (
		_w17431_,
		_w17432_,
		_w17621_
	);
	LUT2 #(
		.INIT('h1)
	) name7110 (
		_w17433_,
		_w17434_,
		_w17622_
	);
	LUT2 #(
		.INIT('h1)
	) name7111 (
		_w17435_,
		_w17436_,
		_w17623_
	);
	LUT2 #(
		.INIT('h1)
	) name7112 (
		_w17437_,
		_w17438_,
		_w17624_
	);
	LUT2 #(
		.INIT('h1)
	) name7113 (
		_w17439_,
		_w17440_,
		_w17625_
	);
	LUT2 #(
		.INIT('h1)
	) name7114 (
		_w17441_,
		_w17442_,
		_w17626_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		_w17443_,
		_w17444_,
		_w17627_
	);
	LUT2 #(
		.INIT('h1)
	) name7116 (
		_w17445_,
		_w17446_,
		_w17628_
	);
	LUT2 #(
		.INIT('h1)
	) name7117 (
		_w17447_,
		_w17448_,
		_w17629_
	);
	LUT2 #(
		.INIT('h1)
	) name7118 (
		_w17449_,
		_w17450_,
		_w17630_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w17451_,
		_w17452_,
		_w17631_
	);
	LUT2 #(
		.INIT('h1)
	) name7120 (
		_w17453_,
		_w17454_,
		_w17632_
	);
	LUT2 #(
		.INIT('h1)
	) name7121 (
		_w17455_,
		_w17456_,
		_w17633_
	);
	LUT2 #(
		.INIT('h1)
	) name7122 (
		_w17457_,
		_w17458_,
		_w17634_
	);
	LUT2 #(
		.INIT('h1)
	) name7123 (
		_w17459_,
		_w17460_,
		_w17635_
	);
	LUT2 #(
		.INIT('h1)
	) name7124 (
		_w17461_,
		_w17462_,
		_w17636_
	);
	LUT2 #(
		.INIT('h1)
	) name7125 (
		_w17463_,
		_w17464_,
		_w17637_
	);
	LUT2 #(
		.INIT('h1)
	) name7126 (
		_w17465_,
		_w17466_,
		_w17638_
	);
	LUT2 #(
		.INIT('h1)
	) name7127 (
		_w17467_,
		_w17468_,
		_w17639_
	);
	LUT2 #(
		.INIT('h1)
	) name7128 (
		_w17469_,
		_w17470_,
		_w17640_
	);
	LUT2 #(
		.INIT('h1)
	) name7129 (
		_w17471_,
		_w17472_,
		_w17641_
	);
	LUT2 #(
		.INIT('h1)
	) name7130 (
		_w17473_,
		_w17474_,
		_w17642_
	);
	LUT2 #(
		.INIT('h1)
	) name7131 (
		_w17475_,
		_w17476_,
		_w17643_
	);
	LUT2 #(
		.INIT('h1)
	) name7132 (
		_w17477_,
		_w17478_,
		_w17644_
	);
	LUT2 #(
		.INIT('h1)
	) name7133 (
		_w17479_,
		_w17480_,
		_w17645_
	);
	LUT2 #(
		.INIT('h1)
	) name7134 (
		_w17481_,
		_w17482_,
		_w17646_
	);
	LUT2 #(
		.INIT('h1)
	) name7135 (
		_w17483_,
		_w17484_,
		_w17647_
	);
	LUT2 #(
		.INIT('h1)
	) name7136 (
		_w17485_,
		_w17486_,
		_w17648_
	);
	LUT2 #(
		.INIT('h1)
	) name7137 (
		_w17487_,
		_w17488_,
		_w17649_
	);
	LUT2 #(
		.INIT('h1)
	) name7138 (
		_w17489_,
		_w17490_,
		_w17650_
	);
	LUT2 #(
		.INIT('h1)
	) name7139 (
		_w17491_,
		_w17492_,
		_w17651_
	);
	LUT2 #(
		.INIT('h1)
	) name7140 (
		_w17493_,
		_w17494_,
		_w17652_
	);
	LUT2 #(
		.INIT('h1)
	) name7141 (
		_w17495_,
		_w17496_,
		_w17653_
	);
	LUT2 #(
		.INIT('h1)
	) name7142 (
		_w17497_,
		_w17498_,
		_w17654_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w17499_,
		_w17500_,
		_w17655_
	);
	LUT2 #(
		.INIT('h1)
	) name7144 (
		_w17501_,
		_w17502_,
		_w17656_
	);
	LUT2 #(
		.INIT('h1)
	) name7145 (
		_w17503_,
		_w17504_,
		_w17657_
	);
	LUT2 #(
		.INIT('h1)
	) name7146 (
		_w17505_,
		_w17506_,
		_w17658_
	);
	LUT2 #(
		.INIT('h1)
	) name7147 (
		_w17507_,
		_w17508_,
		_w17659_
	);
	LUT2 #(
		.INIT('h1)
	) name7148 (
		_w17509_,
		_w17510_,
		_w17660_
	);
	LUT2 #(
		.INIT('h1)
	) name7149 (
		_w17511_,
		_w17512_,
		_w17661_
	);
	LUT2 #(
		.INIT('h1)
	) name7150 (
		_w17513_,
		_w17514_,
		_w17662_
	);
	LUT2 #(
		.INIT('h1)
	) name7151 (
		_w17515_,
		_w17516_,
		_w17663_
	);
	LUT2 #(
		.INIT('h1)
	) name7152 (
		_w17517_,
		_w17518_,
		_w17664_
	);
	LUT2 #(
		.INIT('h1)
	) name7153 (
		_w17519_,
		_w17520_,
		_w17665_
	);
	LUT2 #(
		.INIT('h1)
	) name7154 (
		_w17521_,
		_w17522_,
		_w17666_
	);
	LUT2 #(
		.INIT('h1)
	) name7155 (
		_w17523_,
		_w17524_,
		_w17667_
	);
	LUT2 #(
		.INIT('h1)
	) name7156 (
		_w17525_,
		_w17526_,
		_w17668_
	);
	LUT2 #(
		.INIT('h1)
	) name7157 (
		_w17527_,
		_w17528_,
		_w17669_
	);
	LUT2 #(
		.INIT('h1)
	) name7158 (
		_w17529_,
		_w17530_,
		_w17670_
	);
	LUT2 #(
		.INIT('h1)
	) name7159 (
		_w17531_,
		_w17532_,
		_w17671_
	);
	LUT2 #(
		.INIT('h1)
	) name7160 (
		_w17533_,
		_w17534_,
		_w17672_
	);
	LUT2 #(
		.INIT('h1)
	) name7161 (
		_w17535_,
		_w17536_,
		_w17673_
	);
	LUT2 #(
		.INIT('h1)
	) name7162 (
		_w17537_,
		_w17538_,
		_w17674_
	);
	LUT2 #(
		.INIT('h1)
	) name7163 (
		_w17539_,
		_w17540_,
		_w17675_
	);
	LUT2 #(
		.INIT('h1)
	) name7164 (
		_w17541_,
		_w17542_,
		_w17676_
	);
	LUT2 #(
		.INIT('h1)
	) name7165 (
		_w17543_,
		_w17544_,
		_w17677_
	);
	LUT2 #(
		.INIT('h1)
	) name7166 (
		_w17545_,
		_w17546_,
		_w17678_
	);
	LUT2 #(
		.INIT('h1)
	) name7167 (
		_w17547_,
		_w17548_,
		_w17679_
	);
	LUT2 #(
		.INIT('h1)
	) name7168 (
		_w17549_,
		_w17550_,
		_w17680_
	);
	LUT2 #(
		.INIT('h1)
	) name7169 (
		_w17551_,
		_w17552_,
		_w17681_
	);
	LUT2 #(
		.INIT('h1)
	) name7170 (
		_w17553_,
		_w17554_,
		_w17682_
	);
	LUT2 #(
		.INIT('h8)
	) name7171 (
		_w17681_,
		_w17682_,
		_w17683_
	);
	LUT2 #(
		.INIT('h8)
	) name7172 (
		_w17679_,
		_w17680_,
		_w17684_
	);
	LUT2 #(
		.INIT('h8)
	) name7173 (
		_w17677_,
		_w17678_,
		_w17685_
	);
	LUT2 #(
		.INIT('h8)
	) name7174 (
		_w17675_,
		_w17676_,
		_w17686_
	);
	LUT2 #(
		.INIT('h8)
	) name7175 (
		_w17673_,
		_w17674_,
		_w17687_
	);
	LUT2 #(
		.INIT('h8)
	) name7176 (
		_w17671_,
		_w17672_,
		_w17688_
	);
	LUT2 #(
		.INIT('h8)
	) name7177 (
		_w17669_,
		_w17670_,
		_w17689_
	);
	LUT2 #(
		.INIT('h8)
	) name7178 (
		_w17667_,
		_w17668_,
		_w17690_
	);
	LUT2 #(
		.INIT('h8)
	) name7179 (
		_w17665_,
		_w17666_,
		_w17691_
	);
	LUT2 #(
		.INIT('h8)
	) name7180 (
		_w17663_,
		_w17664_,
		_w17692_
	);
	LUT2 #(
		.INIT('h8)
	) name7181 (
		_w17661_,
		_w17662_,
		_w17693_
	);
	LUT2 #(
		.INIT('h8)
	) name7182 (
		_w17659_,
		_w17660_,
		_w17694_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		_w17657_,
		_w17658_,
		_w17695_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		_w17655_,
		_w17656_,
		_w17696_
	);
	LUT2 #(
		.INIT('h8)
	) name7185 (
		_w17653_,
		_w17654_,
		_w17697_
	);
	LUT2 #(
		.INIT('h8)
	) name7186 (
		_w17651_,
		_w17652_,
		_w17698_
	);
	LUT2 #(
		.INIT('h8)
	) name7187 (
		_w17649_,
		_w17650_,
		_w17699_
	);
	LUT2 #(
		.INIT('h8)
	) name7188 (
		_w17647_,
		_w17648_,
		_w17700_
	);
	LUT2 #(
		.INIT('h8)
	) name7189 (
		_w17645_,
		_w17646_,
		_w17701_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		_w17643_,
		_w17644_,
		_w17702_
	);
	LUT2 #(
		.INIT('h8)
	) name7191 (
		_w17641_,
		_w17642_,
		_w17703_
	);
	LUT2 #(
		.INIT('h8)
	) name7192 (
		_w17639_,
		_w17640_,
		_w17704_
	);
	LUT2 #(
		.INIT('h8)
	) name7193 (
		_w17637_,
		_w17638_,
		_w17705_
	);
	LUT2 #(
		.INIT('h8)
	) name7194 (
		_w17635_,
		_w17636_,
		_w17706_
	);
	LUT2 #(
		.INIT('h8)
	) name7195 (
		_w17633_,
		_w17634_,
		_w17707_
	);
	LUT2 #(
		.INIT('h8)
	) name7196 (
		_w17631_,
		_w17632_,
		_w17708_
	);
	LUT2 #(
		.INIT('h8)
	) name7197 (
		_w17629_,
		_w17630_,
		_w17709_
	);
	LUT2 #(
		.INIT('h8)
	) name7198 (
		_w17627_,
		_w17628_,
		_w17710_
	);
	LUT2 #(
		.INIT('h8)
	) name7199 (
		_w17625_,
		_w17626_,
		_w17711_
	);
	LUT2 #(
		.INIT('h8)
	) name7200 (
		_w17623_,
		_w17624_,
		_w17712_
	);
	LUT2 #(
		.INIT('h8)
	) name7201 (
		_w17621_,
		_w17622_,
		_w17713_
	);
	LUT2 #(
		.INIT('h8)
	) name7202 (
		_w17619_,
		_w17620_,
		_w17714_
	);
	LUT2 #(
		.INIT('h8)
	) name7203 (
		_w17617_,
		_w17618_,
		_w17715_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		_w17615_,
		_w17616_,
		_w17716_
	);
	LUT2 #(
		.INIT('h8)
	) name7205 (
		_w17613_,
		_w17614_,
		_w17717_
	);
	LUT2 #(
		.INIT('h8)
	) name7206 (
		_w17611_,
		_w17612_,
		_w17718_
	);
	LUT2 #(
		.INIT('h8)
	) name7207 (
		_w17609_,
		_w17610_,
		_w17719_
	);
	LUT2 #(
		.INIT('h8)
	) name7208 (
		_w17607_,
		_w17608_,
		_w17720_
	);
	LUT2 #(
		.INIT('h8)
	) name7209 (
		_w17605_,
		_w17606_,
		_w17721_
	);
	LUT2 #(
		.INIT('h8)
	) name7210 (
		_w17603_,
		_w17604_,
		_w17722_
	);
	LUT2 #(
		.INIT('h8)
	) name7211 (
		_w17601_,
		_w17602_,
		_w17723_
	);
	LUT2 #(
		.INIT('h8)
	) name7212 (
		_w17599_,
		_w17600_,
		_w17724_
	);
	LUT2 #(
		.INIT('h8)
	) name7213 (
		_w17597_,
		_w17598_,
		_w17725_
	);
	LUT2 #(
		.INIT('h8)
	) name7214 (
		_w17595_,
		_w17596_,
		_w17726_
	);
	LUT2 #(
		.INIT('h8)
	) name7215 (
		_w17593_,
		_w17594_,
		_w17727_
	);
	LUT2 #(
		.INIT('h8)
	) name7216 (
		_w17591_,
		_w17592_,
		_w17728_
	);
	LUT2 #(
		.INIT('h8)
	) name7217 (
		_w17589_,
		_w17590_,
		_w17729_
	);
	LUT2 #(
		.INIT('h8)
	) name7218 (
		_w17587_,
		_w17588_,
		_w17730_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		_w17585_,
		_w17586_,
		_w17731_
	);
	LUT2 #(
		.INIT('h8)
	) name7220 (
		_w17583_,
		_w17584_,
		_w17732_
	);
	LUT2 #(
		.INIT('h8)
	) name7221 (
		_w17581_,
		_w17582_,
		_w17733_
	);
	LUT2 #(
		.INIT('h8)
	) name7222 (
		_w17579_,
		_w17580_,
		_w17734_
	);
	LUT2 #(
		.INIT('h8)
	) name7223 (
		_w17577_,
		_w17578_,
		_w17735_
	);
	LUT2 #(
		.INIT('h8)
	) name7224 (
		_w17575_,
		_w17576_,
		_w17736_
	);
	LUT2 #(
		.INIT('h8)
	) name7225 (
		_w17573_,
		_w17574_,
		_w17737_
	);
	LUT2 #(
		.INIT('h8)
	) name7226 (
		_w17571_,
		_w17572_,
		_w17738_
	);
	LUT2 #(
		.INIT('h8)
	) name7227 (
		_w17569_,
		_w17570_,
		_w17739_
	);
	LUT2 #(
		.INIT('h8)
	) name7228 (
		_w17567_,
		_w17568_,
		_w17740_
	);
	LUT2 #(
		.INIT('h8)
	) name7229 (
		_w17565_,
		_w17566_,
		_w17741_
	);
	LUT2 #(
		.INIT('h8)
	) name7230 (
		_w17563_,
		_w17564_,
		_w17742_
	);
	LUT2 #(
		.INIT('h8)
	) name7231 (
		_w17561_,
		_w17562_,
		_w17743_
	);
	LUT2 #(
		.INIT('h8)
	) name7232 (
		_w17559_,
		_w17560_,
		_w17744_
	);
	LUT2 #(
		.INIT('h8)
	) name7233 (
		_w17557_,
		_w17558_,
		_w17745_
	);
	LUT2 #(
		.INIT('h8)
	) name7234 (
		_w17555_,
		_w17556_,
		_w17746_
	);
	LUT2 #(
		.INIT('h8)
	) name7235 (
		_w17745_,
		_w17746_,
		_w17747_
	);
	LUT2 #(
		.INIT('h8)
	) name7236 (
		_w17743_,
		_w17744_,
		_w17748_
	);
	LUT2 #(
		.INIT('h8)
	) name7237 (
		_w17741_,
		_w17742_,
		_w17749_
	);
	LUT2 #(
		.INIT('h8)
	) name7238 (
		_w17739_,
		_w17740_,
		_w17750_
	);
	LUT2 #(
		.INIT('h8)
	) name7239 (
		_w17737_,
		_w17738_,
		_w17751_
	);
	LUT2 #(
		.INIT('h8)
	) name7240 (
		_w17735_,
		_w17736_,
		_w17752_
	);
	LUT2 #(
		.INIT('h8)
	) name7241 (
		_w17733_,
		_w17734_,
		_w17753_
	);
	LUT2 #(
		.INIT('h8)
	) name7242 (
		_w17731_,
		_w17732_,
		_w17754_
	);
	LUT2 #(
		.INIT('h8)
	) name7243 (
		_w17729_,
		_w17730_,
		_w17755_
	);
	LUT2 #(
		.INIT('h8)
	) name7244 (
		_w17727_,
		_w17728_,
		_w17756_
	);
	LUT2 #(
		.INIT('h8)
	) name7245 (
		_w17725_,
		_w17726_,
		_w17757_
	);
	LUT2 #(
		.INIT('h8)
	) name7246 (
		_w17723_,
		_w17724_,
		_w17758_
	);
	LUT2 #(
		.INIT('h8)
	) name7247 (
		_w17721_,
		_w17722_,
		_w17759_
	);
	LUT2 #(
		.INIT('h8)
	) name7248 (
		_w17719_,
		_w17720_,
		_w17760_
	);
	LUT2 #(
		.INIT('h8)
	) name7249 (
		_w17717_,
		_w17718_,
		_w17761_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		_w17715_,
		_w17716_,
		_w17762_
	);
	LUT2 #(
		.INIT('h8)
	) name7251 (
		_w17713_,
		_w17714_,
		_w17763_
	);
	LUT2 #(
		.INIT('h8)
	) name7252 (
		_w17711_,
		_w17712_,
		_w17764_
	);
	LUT2 #(
		.INIT('h8)
	) name7253 (
		_w17709_,
		_w17710_,
		_w17765_
	);
	LUT2 #(
		.INIT('h8)
	) name7254 (
		_w17707_,
		_w17708_,
		_w17766_
	);
	LUT2 #(
		.INIT('h8)
	) name7255 (
		_w17705_,
		_w17706_,
		_w17767_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		_w17703_,
		_w17704_,
		_w17768_
	);
	LUT2 #(
		.INIT('h8)
	) name7257 (
		_w17701_,
		_w17702_,
		_w17769_
	);
	LUT2 #(
		.INIT('h8)
	) name7258 (
		_w17699_,
		_w17700_,
		_w17770_
	);
	LUT2 #(
		.INIT('h8)
	) name7259 (
		_w17697_,
		_w17698_,
		_w17771_
	);
	LUT2 #(
		.INIT('h8)
	) name7260 (
		_w17695_,
		_w17696_,
		_w17772_
	);
	LUT2 #(
		.INIT('h8)
	) name7261 (
		_w17693_,
		_w17694_,
		_w17773_
	);
	LUT2 #(
		.INIT('h8)
	) name7262 (
		_w17691_,
		_w17692_,
		_w17774_
	);
	LUT2 #(
		.INIT('h8)
	) name7263 (
		_w17689_,
		_w17690_,
		_w17775_
	);
	LUT2 #(
		.INIT('h8)
	) name7264 (
		_w17687_,
		_w17688_,
		_w17776_
	);
	LUT2 #(
		.INIT('h8)
	) name7265 (
		_w17685_,
		_w17686_,
		_w17777_
	);
	LUT2 #(
		.INIT('h8)
	) name7266 (
		_w17683_,
		_w17684_,
		_w17778_
	);
	LUT2 #(
		.INIT('h8)
	) name7267 (
		_w17777_,
		_w17778_,
		_w17779_
	);
	LUT2 #(
		.INIT('h8)
	) name7268 (
		_w17775_,
		_w17776_,
		_w17780_
	);
	LUT2 #(
		.INIT('h8)
	) name7269 (
		_w17773_,
		_w17774_,
		_w17781_
	);
	LUT2 #(
		.INIT('h8)
	) name7270 (
		_w17771_,
		_w17772_,
		_w17782_
	);
	LUT2 #(
		.INIT('h8)
	) name7271 (
		_w17769_,
		_w17770_,
		_w17783_
	);
	LUT2 #(
		.INIT('h8)
	) name7272 (
		_w17767_,
		_w17768_,
		_w17784_
	);
	LUT2 #(
		.INIT('h8)
	) name7273 (
		_w17765_,
		_w17766_,
		_w17785_
	);
	LUT2 #(
		.INIT('h8)
	) name7274 (
		_w17763_,
		_w17764_,
		_w17786_
	);
	LUT2 #(
		.INIT('h8)
	) name7275 (
		_w17761_,
		_w17762_,
		_w17787_
	);
	LUT2 #(
		.INIT('h8)
	) name7276 (
		_w17759_,
		_w17760_,
		_w17788_
	);
	LUT2 #(
		.INIT('h8)
	) name7277 (
		_w17757_,
		_w17758_,
		_w17789_
	);
	LUT2 #(
		.INIT('h8)
	) name7278 (
		_w17755_,
		_w17756_,
		_w17790_
	);
	LUT2 #(
		.INIT('h8)
	) name7279 (
		_w17753_,
		_w17754_,
		_w17791_
	);
	LUT2 #(
		.INIT('h8)
	) name7280 (
		_w17751_,
		_w17752_,
		_w17792_
	);
	LUT2 #(
		.INIT('h8)
	) name7281 (
		_w17749_,
		_w17750_,
		_w17793_
	);
	LUT2 #(
		.INIT('h8)
	) name7282 (
		_w17747_,
		_w17748_,
		_w17794_
	);
	LUT2 #(
		.INIT('h8)
	) name7283 (
		_w17793_,
		_w17794_,
		_w17795_
	);
	LUT2 #(
		.INIT('h8)
	) name7284 (
		_w17791_,
		_w17792_,
		_w17796_
	);
	LUT2 #(
		.INIT('h8)
	) name7285 (
		_w17789_,
		_w17790_,
		_w17797_
	);
	LUT2 #(
		.INIT('h8)
	) name7286 (
		_w17787_,
		_w17788_,
		_w17798_
	);
	LUT2 #(
		.INIT('h8)
	) name7287 (
		_w17785_,
		_w17786_,
		_w17799_
	);
	LUT2 #(
		.INIT('h8)
	) name7288 (
		_w17783_,
		_w17784_,
		_w17800_
	);
	LUT2 #(
		.INIT('h8)
	) name7289 (
		_w17781_,
		_w17782_,
		_w17801_
	);
	LUT2 #(
		.INIT('h8)
	) name7290 (
		_w17779_,
		_w17780_,
		_w17802_
	);
	LUT2 #(
		.INIT('h8)
	) name7291 (
		_w17801_,
		_w17802_,
		_w17803_
	);
	LUT2 #(
		.INIT('h8)
	) name7292 (
		_w17799_,
		_w17800_,
		_w17804_
	);
	LUT2 #(
		.INIT('h8)
	) name7293 (
		_w17797_,
		_w17798_,
		_w17805_
	);
	LUT2 #(
		.INIT('h8)
	) name7294 (
		_w17795_,
		_w17796_,
		_w17806_
	);
	LUT2 #(
		.INIT('h8)
	) name7295 (
		_w17805_,
		_w17806_,
		_w17807_
	);
	LUT2 #(
		.INIT('h8)
	) name7296 (
		_w17803_,
		_w17804_,
		_w17808_
	);
	LUT2 #(
		.INIT('h8)
	) name7297 (
		_w17807_,
		_w17808_,
		_w17809_
	);
	LUT2 #(
		.INIT('h1)
	) name7298 (
		wb_rst_i_pad,
		_w17809_,
		_w17810_
	);
	LUT2 #(
		.INIT('h8)
	) name7299 (
		_w12656_,
		_w17810_,
		_w17811_
	);
	LUT2 #(
		.INIT('h8)
	) name7300 (
		_w13483_,
		_w17289_,
		_w17812_
	);
	LUT2 #(
		.INIT('h8)
	) name7301 (
		_w13478_,
		_w17812_,
		_w17813_
	);
	LUT2 #(
		.INIT('h2)
	) name7302 (
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w17813_,
		_w17814_
	);
	LUT2 #(
		.INIT('h1)
	) name7303 (
		_w13484_,
		_w17814_,
		_w17815_
	);
	LUT2 #(
		.INIT('h1)
	) name7304 (
		\wishbone_TxLength_reg[9]/NET0131 ,
		_w17289_,
		_w17816_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w12656_,
		_w13499_,
		_w17817_
	);
	LUT2 #(
		.INIT('h1)
	) name7306 (
		_w12658_,
		_w17817_,
		_w17818_
	);
	LUT2 #(
		.INIT('h1)
	) name7307 (
		_w17816_,
		_w17818_,
		_w17819_
	);
	LUT2 #(
		.INIT('h4)
	) name7308 (
		_w17815_,
		_w17819_,
		_w17820_
	);
	LUT2 #(
		.INIT('h1)
	) name7309 (
		_w17811_,
		_w17820_,
		_w17821_
	);
	LUT2 #(
		.INIT('h8)
	) name7310 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		_w15147_,
		_w17822_
	);
	LUT2 #(
		.INIT('h4)
	) name7311 (
		_w15147_,
		_w15150_,
		_w17823_
	);
	LUT2 #(
		.INIT('h1)
	) name7312 (
		_w15149_,
		_w17823_,
		_w17824_
	);
	LUT2 #(
		.INIT('h2)
	) name7313 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w17824_,
		_w17825_
	);
	LUT2 #(
		.INIT('h1)
	) name7314 (
		_w17822_,
		_w17825_,
		_w17826_
	);
	LUT2 #(
		.INIT('h8)
	) name7315 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w15147_,
		_w17827_
	);
	LUT2 #(
		.INIT('h2)
	) name7316 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w17824_,
		_w17828_
	);
	LUT2 #(
		.INIT('h1)
	) name7317 (
		_w17827_,
		_w17828_,
		_w17829_
	);
	LUT2 #(
		.INIT('h8)
	) name7318 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		_w15147_,
		_w17830_
	);
	LUT2 #(
		.INIT('h2)
	) name7319 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w17824_,
		_w17831_
	);
	LUT2 #(
		.INIT('h1)
	) name7320 (
		_w17830_,
		_w17831_,
		_w17832_
	);
	LUT2 #(
		.INIT('h8)
	) name7321 (
		\wishbone_RxDataLatched2_reg[3]/NET0131 ,
		_w15147_,
		_w17833_
	);
	LUT2 #(
		.INIT('h2)
	) name7322 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w17824_,
		_w17834_
	);
	LUT2 #(
		.INIT('h1)
	) name7323 (
		_w17833_,
		_w17834_,
		_w17835_
	);
	LUT2 #(
		.INIT('h8)
	) name7324 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		_w15147_,
		_w17836_
	);
	LUT2 #(
		.INIT('h2)
	) name7325 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w17824_,
		_w17837_
	);
	LUT2 #(
		.INIT('h1)
	) name7326 (
		_w17836_,
		_w17837_,
		_w17838_
	);
	LUT2 #(
		.INIT('h8)
	) name7327 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w15147_,
		_w17839_
	);
	LUT2 #(
		.INIT('h2)
	) name7328 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w17824_,
		_w17840_
	);
	LUT2 #(
		.INIT('h1)
	) name7329 (
		_w17839_,
		_w17840_,
		_w17841_
	);
	LUT2 #(
		.INIT('h8)
	) name7330 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		_w15147_,
		_w17842_
	);
	LUT2 #(
		.INIT('h2)
	) name7331 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w17824_,
		_w17843_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		_w17842_,
		_w17843_,
		_w17844_
	);
	LUT2 #(
		.INIT('h8)
	) name7333 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w15147_,
		_w17845_
	);
	LUT2 #(
		.INIT('h2)
	) name7334 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w17824_,
		_w17846_
	);
	LUT2 #(
		.INIT('h1)
	) name7335 (
		_w17845_,
		_w17846_,
		_w17847_
	);
	LUT2 #(
		.INIT('h8)
	) name7336 (
		_w14536_,
		_w15696_,
		_w17848_
	);
	LUT2 #(
		.INIT('h8)
	) name7337 (
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		_w15698_,
		_w17849_
	);
	LUT2 #(
		.INIT('h8)
	) name7338 (
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w17849_,
		_w17850_
	);
	LUT2 #(
		.INIT('h8)
	) name7339 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		_w17850_,
		_w17851_
	);
	LUT2 #(
		.INIT('h8)
	) name7340 (
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w17851_,
		_w17852_
	);
	LUT2 #(
		.INIT('h8)
	) name7341 (
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w17852_,
		_w17853_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		_w17853_,
		_w17854_
	);
	LUT2 #(
		.INIT('h8)
	) name7343 (
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w17855_
	);
	LUT2 #(
		.INIT('h8)
	) name7344 (
		_w17854_,
		_w17855_,
		_w17856_
	);
	LUT2 #(
		.INIT('h8)
	) name7345 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		_w17856_,
		_w17857_
	);
	LUT2 #(
		.INIT('h8)
	) name7346 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		_w17857_,
		_w17858_
	);
	LUT2 #(
		.INIT('h8)
	) name7347 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w17859_
	);
	LUT2 #(
		.INIT('h8)
	) name7348 (
		_w17858_,
		_w17859_,
		_w17860_
	);
	LUT2 #(
		.INIT('h8)
	) name7349 (
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w17860_,
		_w17861_
	);
	LUT2 #(
		.INIT('h8)
	) name7350 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w17861_,
		_w17862_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w17863_
	);
	LUT2 #(
		.INIT('h8)
	) name7352 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w17864_
	);
	LUT2 #(
		.INIT('h8)
	) name7353 (
		_w17863_,
		_w17864_,
		_w17865_
	);
	LUT2 #(
		.INIT('h8)
	) name7354 (
		_w17862_,
		_w17865_,
		_w17866_
	);
	LUT2 #(
		.INIT('h8)
	) name7355 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w17866_,
		_w17867_
	);
	LUT2 #(
		.INIT('h8)
	) name7356 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w17868_
	);
	LUT2 #(
		.INIT('h8)
	) name7357 (
		_w17867_,
		_w17868_,
		_w17869_
	);
	LUT2 #(
		.INIT('h8)
	) name7358 (
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w17869_,
		_w17870_
	);
	LUT2 #(
		.INIT('h8)
	) name7359 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w17870_,
		_w17871_
	);
	LUT2 #(
		.INIT('h8)
	) name7360 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		_w17871_,
		_w17872_
	);
	LUT2 #(
		.INIT('h8)
	) name7361 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w17873_
	);
	LUT2 #(
		.INIT('h8)
	) name7362 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w17873_,
		_w17874_
	);
	LUT2 #(
		.INIT('h8)
	) name7363 (
		_w17872_,
		_w17874_,
		_w17875_
	);
	LUT2 #(
		.INIT('h8)
	) name7364 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w17875_,
		_w17876_
	);
	LUT2 #(
		.INIT('h1)
	) name7365 (
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w17876_,
		_w17877_
	);
	LUT2 #(
		.INIT('h8)
	) name7366 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		\wishbone_RxPointerMSB_reg[30]/NET0131 ,
		_w17878_
	);
	LUT2 #(
		.INIT('h8)
	) name7367 (
		_w17875_,
		_w17878_,
		_w17879_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w15696_,
		_w17879_,
		_w17880_
	);
	LUT2 #(
		.INIT('h4)
	) name7369 (
		_w17877_,
		_w17880_,
		_w17881_
	);
	LUT2 #(
		.INIT('h1)
	) name7370 (
		_w17848_,
		_w17881_,
		_w17882_
	);
	LUT2 #(
		.INIT('h8)
	) name7371 (
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w12655_,
		_w17883_
	);
	LUT2 #(
		.INIT('h8)
	) name7372 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w17884_
	);
	LUT2 #(
		.INIT('h4)
	) name7373 (
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w17885_
	);
	LUT2 #(
		.INIT('h8)
	) name7374 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w17885_,
		_w17886_
	);
	LUT2 #(
		.INIT('h8)
	) name7375 (
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w17886_,
		_w17887_
	);
	LUT2 #(
		.INIT('h8)
	) name7376 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		_w17887_,
		_w17888_
	);
	LUT2 #(
		.INIT('h8)
	) name7377 (
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w17888_,
		_w17889_
	);
	LUT2 #(
		.INIT('h8)
	) name7378 (
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w17889_,
		_w17890_
	);
	LUT2 #(
		.INIT('h8)
	) name7379 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		_w17890_,
		_w17891_
	);
	LUT2 #(
		.INIT('h8)
	) name7380 (
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w17891_,
		_w17892_
	);
	LUT2 #(
		.INIT('h8)
	) name7381 (
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w17892_,
		_w17893_
	);
	LUT2 #(
		.INIT('h8)
	) name7382 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		_w17893_,
		_w17894_
	);
	LUT2 #(
		.INIT('h8)
	) name7383 (
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w17894_,
		_w17895_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w17895_,
		_w17896_
	);
	LUT2 #(
		.INIT('h8)
	) name7385 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w17897_
	);
	LUT2 #(
		.INIT('h8)
	) name7386 (
		_w17896_,
		_w17897_,
		_w17898_
	);
	LUT2 #(
		.INIT('h8)
	) name7387 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w17899_
	);
	LUT2 #(
		.INIT('h8)
	) name7388 (
		_w17898_,
		_w17899_,
		_w17900_
	);
	LUT2 #(
		.INIT('h8)
	) name7389 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w17900_,
		_w17901_
	);
	LUT2 #(
		.INIT('h8)
	) name7390 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		_w17901_,
		_w17902_
	);
	LUT2 #(
		.INIT('h8)
	) name7391 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w17903_
	);
	LUT2 #(
		.INIT('h8)
	) name7392 (
		_w17902_,
		_w17903_,
		_w17904_
	);
	LUT2 #(
		.INIT('h8)
	) name7393 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w17905_
	);
	LUT2 #(
		.INIT('h8)
	) name7394 (
		_w17904_,
		_w17905_,
		_w17906_
	);
	LUT2 #(
		.INIT('h8)
	) name7395 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w17907_
	);
	LUT2 #(
		.INIT('h8)
	) name7396 (
		_w17906_,
		_w17907_,
		_w17908_
	);
	LUT2 #(
		.INIT('h8)
	) name7397 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w17909_
	);
	LUT2 #(
		.INIT('h8)
	) name7398 (
		_w17908_,
		_w17909_,
		_w17910_
	);
	LUT2 #(
		.INIT('h8)
	) name7399 (
		_w17884_,
		_w17910_,
		_w17911_
	);
	LUT2 #(
		.INIT('h8)
	) name7400 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w17912_
	);
	LUT2 #(
		.INIT('h1)
	) name7401 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w17913_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w17912_,
		_w17913_,
		_w17914_
	);
	LUT2 #(
		.INIT('h2)
	) name7403 (
		_w17911_,
		_w17914_,
		_w17915_
	);
	LUT2 #(
		.INIT('h1)
	) name7404 (
		\wishbone_TxPointerMSB_reg[30]/NET0131 ,
		_w17911_,
		_w17916_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		_w17915_,
		_w17916_,
		_w17917_
	);
	LUT2 #(
		.INIT('h1)
	) name7406 (
		_w17883_,
		_w17917_,
		_w17918_
	);
	LUT2 #(
		.INIT('h4)
	) name7407 (
		_w14536_,
		_w17883_,
		_w17919_
	);
	LUT2 #(
		.INIT('h1)
	) name7408 (
		_w17918_,
		_w17919_,
		_w17920_
	);
	LUT2 #(
		.INIT('h8)
	) name7409 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w15147_,
		_w17921_
	);
	LUT2 #(
		.INIT('h2)
	) name7410 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w17922_
	);
	LUT2 #(
		.INIT('h8)
	) name7411 (
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w17922_,
		_w17923_
	);
	LUT2 #(
		.INIT('h1)
	) name7412 (
		_w15147_,
		_w17923_,
		_w17924_
	);
	LUT2 #(
		.INIT('h8)
	) name7413 (
		\wishbone_RxDataLatched1_reg[16]/NET0131 ,
		_w17924_,
		_w17925_
	);
	LUT2 #(
		.INIT('h1)
	) name7414 (
		_w17921_,
		_w17925_,
		_w17926_
	);
	LUT2 #(
		.INIT('h8)
	) name7415 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		_w15147_,
		_w17927_
	);
	LUT2 #(
		.INIT('h8)
	) name7416 (
		\wishbone_RxDataLatched1_reg[17]/NET0131 ,
		_w17924_,
		_w17928_
	);
	LUT2 #(
		.INIT('h1)
	) name7417 (
		_w17927_,
		_w17928_,
		_w17929_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		_w15147_,
		_w17930_
	);
	LUT2 #(
		.INIT('h8)
	) name7419 (
		\wishbone_RxDataLatched1_reg[18]/NET0131 ,
		_w17924_,
		_w17931_
	);
	LUT2 #(
		.INIT('h1)
	) name7420 (
		_w17930_,
		_w17931_,
		_w17932_
	);
	LUT2 #(
		.INIT('h8)
	) name7421 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w15147_,
		_w17933_
	);
	LUT2 #(
		.INIT('h8)
	) name7422 (
		\wishbone_RxDataLatched1_reg[19]/NET0131 ,
		_w17924_,
		_w17934_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		_w17933_,
		_w17934_,
		_w17935_
	);
	LUT2 #(
		.INIT('h8)
	) name7424 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		_w15147_,
		_w17936_
	);
	LUT2 #(
		.INIT('h8)
	) name7425 (
		\wishbone_RxDataLatched1_reg[20]/NET0131 ,
		_w17924_,
		_w17937_
	);
	LUT2 #(
		.INIT('h1)
	) name7426 (
		_w17936_,
		_w17937_,
		_w17938_
	);
	LUT2 #(
		.INIT('h8)
	) name7427 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w15147_,
		_w17939_
	);
	LUT2 #(
		.INIT('h8)
	) name7428 (
		\wishbone_RxDataLatched1_reg[21]/NET0131 ,
		_w17924_,
		_w17940_
	);
	LUT2 #(
		.INIT('h1)
	) name7429 (
		_w17939_,
		_w17940_,
		_w17941_
	);
	LUT2 #(
		.INIT('h8)
	) name7430 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w15147_,
		_w17942_
	);
	LUT2 #(
		.INIT('h8)
	) name7431 (
		\wishbone_RxDataLatched1_reg[22]/NET0131 ,
		_w17924_,
		_w17943_
	);
	LUT2 #(
		.INIT('h1)
	) name7432 (
		_w17942_,
		_w17943_,
		_w17944_
	);
	LUT2 #(
		.INIT('h8)
	) name7433 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w15147_,
		_w17945_
	);
	LUT2 #(
		.INIT('h8)
	) name7434 (
		\wishbone_RxDataLatched1_reg[23]/NET0131 ,
		_w17924_,
		_w17946_
	);
	LUT2 #(
		.INIT('h1)
	) name7435 (
		_w17945_,
		_w17946_,
		_w17947_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		_w12577_,
		_w17948_
	);
	LUT2 #(
		.INIT('h8)
	) name7437 (
		\m_wb_adr_o[13]_pad ,
		_w12588_,
		_w17949_
	);
	LUT2 #(
		.INIT('h4)
	) name7438 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w12608_,
		_w17950_
	);
	LUT2 #(
		.INIT('h2)
	) name7439 (
		_w12621_,
		_w17950_,
		_w17951_
	);
	LUT2 #(
		.INIT('h1)
	) name7440 (
		_w12623_,
		_w17951_,
		_w17952_
	);
	LUT2 #(
		.INIT('h1)
	) name7441 (
		\m_wb_adr_o[13]_pad ,
		_w12588_,
		_w17953_
	);
	LUT2 #(
		.INIT('h1)
	) name7442 (
		_w17949_,
		_w17952_,
		_w17954_
	);
	LUT2 #(
		.INIT('h4)
	) name7443 (
		_w17953_,
		_w17954_,
		_w17955_
	);
	LUT2 #(
		.INIT('h8)
	) name7444 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w12634_,
		_w17956_
	);
	LUT2 #(
		.INIT('h8)
	) name7445 (
		\m_wb_adr_o[13]_pad ,
		_w12636_,
		_w17957_
	);
	LUT2 #(
		.INIT('h1)
	) name7446 (
		_w17948_,
		_w17956_,
		_w17958_
	);
	LUT2 #(
		.INIT('h4)
	) name7447 (
		_w17957_,
		_w17958_,
		_w17959_
	);
	LUT2 #(
		.INIT('h4)
	) name7448 (
		_w17955_,
		_w17959_,
		_w17960_
	);
	LUT2 #(
		.INIT('h1)
	) name7449 (
		\m_wb_adr_o[14]_pad ,
		_w17949_,
		_w17961_
	);
	LUT2 #(
		.INIT('h1)
	) name7450 (
		_w12590_,
		_w17961_,
		_w17962_
	);
	LUT2 #(
		.INIT('h4)
	) name7451 (
		_w14591_,
		_w17962_,
		_w17963_
	);
	LUT2 #(
		.INIT('h8)
	) name7452 (
		\m_wb_adr_o[14]_pad ,
		_w12636_,
		_w17964_
	);
	LUT2 #(
		.INIT('h2)
	) name7453 (
		_w12576_,
		_w17962_,
		_w17965_
	);
	LUT2 #(
		.INIT('h2)
	) name7454 (
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w12573_,
		_w17966_
	);
	LUT2 #(
		.INIT('h4)
	) name7455 (
		_w17965_,
		_w17966_,
		_w17967_
	);
	LUT2 #(
		.INIT('h2)
	) name7456 (
		_w12633_,
		_w17962_,
		_w17968_
	);
	LUT2 #(
		.INIT('h2)
	) name7457 (
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w12632_,
		_w17969_
	);
	LUT2 #(
		.INIT('h4)
	) name7458 (
		_w17968_,
		_w17969_,
		_w17970_
	);
	LUT2 #(
		.INIT('h1)
	) name7459 (
		_w17963_,
		_w17964_,
		_w17971_
	);
	LUT2 #(
		.INIT('h4)
	) name7460 (
		_w17967_,
		_w17971_,
		_w17972_
	);
	LUT2 #(
		.INIT('h4)
	) name7461 (
		_w17970_,
		_w17972_,
		_w17973_
	);
	LUT2 #(
		.INIT('h8)
	) name7462 (
		\m_wb_adr_o[8]_pad ,
		_w12636_,
		_w17974_
	);
	LUT2 #(
		.INIT('h8)
	) name7463 (
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w12577_,
		_w17975_
	);
	LUT2 #(
		.INIT('h8)
	) name7464 (
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w12634_,
		_w17976_
	);
	LUT2 #(
		.INIT('h1)
	) name7465 (
		\m_wb_adr_o[8]_pad ,
		_w12583_,
		_w17977_
	);
	LUT2 #(
		.INIT('h1)
	) name7466 (
		_w12584_,
		_w17977_,
		_w17978_
	);
	LUT2 #(
		.INIT('h4)
	) name7467 (
		_w14591_,
		_w17978_,
		_w17979_
	);
	LUT2 #(
		.INIT('h1)
	) name7468 (
		_w17974_,
		_w17976_,
		_w17980_
	);
	LUT2 #(
		.INIT('h1)
	) name7469 (
		_w17975_,
		_w17979_,
		_w17981_
	);
	LUT2 #(
		.INIT('h8)
	) name7470 (
		_w17980_,
		_w17981_,
		_w17982_
	);
	LUT2 #(
		.INIT('h8)
	) name7471 (
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w12577_,
		_w17983_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		\m_wb_adr_o[11]_pad ,
		_w12586_,
		_w17984_
	);
	LUT2 #(
		.INIT('h4)
	) name7473 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		_w12608_,
		_w17985_
	);
	LUT2 #(
		.INIT('h2)
	) name7474 (
		_w12621_,
		_w17985_,
		_w17986_
	);
	LUT2 #(
		.INIT('h1)
	) name7475 (
		_w12623_,
		_w17986_,
		_w17987_
	);
	LUT2 #(
		.INIT('h1)
	) name7476 (
		_w12587_,
		_w17984_,
		_w17988_
	);
	LUT2 #(
		.INIT('h4)
	) name7477 (
		_w17987_,
		_w17988_,
		_w17989_
	);
	LUT2 #(
		.INIT('h8)
	) name7478 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		_w12634_,
		_w17990_
	);
	LUT2 #(
		.INIT('h8)
	) name7479 (
		\m_wb_adr_o[11]_pad ,
		_w12636_,
		_w17991_
	);
	LUT2 #(
		.INIT('h1)
	) name7480 (
		_w17983_,
		_w17990_,
		_w17992_
	);
	LUT2 #(
		.INIT('h4)
	) name7481 (
		_w17991_,
		_w17992_,
		_w17993_
	);
	LUT2 #(
		.INIT('h4)
	) name7482 (
		_w17989_,
		_w17993_,
		_w17994_
	);
	LUT2 #(
		.INIT('h8)
	) name7483 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w12577_,
		_w17995_
	);
	LUT2 #(
		.INIT('h1)
	) name7484 (
		\m_wb_adr_o[15]_pad ,
		_w12590_,
		_w17996_
	);
	LUT2 #(
		.INIT('h8)
	) name7485 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w12561_,
		_w17997_
	);
	LUT2 #(
		.INIT('h2)
	) name7486 (
		_w14591_,
		_w17997_,
		_w17998_
	);
	LUT2 #(
		.INIT('h1)
	) name7487 (
		_w12591_,
		_w17998_,
		_w17999_
	);
	LUT2 #(
		.INIT('h4)
	) name7488 (
		_w17996_,
		_w17999_,
		_w18000_
	);
	LUT2 #(
		.INIT('h8)
	) name7489 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w12634_,
		_w18001_
	);
	LUT2 #(
		.INIT('h8)
	) name7490 (
		\m_wb_adr_o[15]_pad ,
		_w12636_,
		_w18002_
	);
	LUT2 #(
		.INIT('h1)
	) name7491 (
		_w17995_,
		_w18001_,
		_w18003_
	);
	LUT2 #(
		.INIT('h4)
	) name7492 (
		_w18002_,
		_w18003_,
		_w18004_
	);
	LUT2 #(
		.INIT('h4)
	) name7493 (
		_w18000_,
		_w18004_,
		_w18005_
	);
	LUT2 #(
		.INIT('h8)
	) name7494 (
		\m_wb_adr_o[4]_pad ,
		_w12636_,
		_w18006_
	);
	LUT2 #(
		.INIT('h8)
	) name7495 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		_w12577_,
		_w18007_
	);
	LUT2 #(
		.INIT('h8)
	) name7496 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		_w12634_,
		_w18008_
	);
	LUT2 #(
		.INIT('h1)
	) name7497 (
		\m_wb_adr_o[4]_pad ,
		_w12579_,
		_w18009_
	);
	LUT2 #(
		.INIT('h1)
	) name7498 (
		_w12580_,
		_w18009_,
		_w18010_
	);
	LUT2 #(
		.INIT('h4)
	) name7499 (
		_w14591_,
		_w18010_,
		_w18011_
	);
	LUT2 #(
		.INIT('h1)
	) name7500 (
		_w18006_,
		_w18008_,
		_w18012_
	);
	LUT2 #(
		.INIT('h1)
	) name7501 (
		_w18007_,
		_w18011_,
		_w18013_
	);
	LUT2 #(
		.INIT('h8)
	) name7502 (
		_w18012_,
		_w18013_,
		_w18014_
	);
	LUT2 #(
		.INIT('h8)
	) name7503 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w12577_,
		_w18015_
	);
	LUT2 #(
		.INIT('h1)
	) name7504 (
		\m_wb_adr_o[27]_pad ,
		_w12602_,
		_w18016_
	);
	LUT2 #(
		.INIT('h8)
	) name7505 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w12561_,
		_w18017_
	);
	LUT2 #(
		.INIT('h2)
	) name7506 (
		_w14591_,
		_w18017_,
		_w18018_
	);
	LUT2 #(
		.INIT('h8)
	) name7507 (
		\m_wb_adr_o[27]_pad ,
		_w12602_,
		_w18019_
	);
	LUT2 #(
		.INIT('h1)
	) name7508 (
		_w18016_,
		_w18018_,
		_w18020_
	);
	LUT2 #(
		.INIT('h4)
	) name7509 (
		_w18019_,
		_w18020_,
		_w18021_
	);
	LUT2 #(
		.INIT('h8)
	) name7510 (
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w12634_,
		_w18022_
	);
	LUT2 #(
		.INIT('h8)
	) name7511 (
		\m_wb_adr_o[27]_pad ,
		_w12636_,
		_w18023_
	);
	LUT2 #(
		.INIT('h1)
	) name7512 (
		_w18015_,
		_w18022_,
		_w18024_
	);
	LUT2 #(
		.INIT('h4)
	) name7513 (
		_w18023_,
		_w18024_,
		_w18025_
	);
	LUT2 #(
		.INIT('h4)
	) name7514 (
		_w18021_,
		_w18025_,
		_w18026_
	);
	LUT2 #(
		.INIT('h8)
	) name7515 (
		\m_wb_adr_o[31]_pad ,
		_w12636_,
		_w18027_
	);
	LUT2 #(
		.INIT('h8)
	) name7516 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w12634_,
		_w18028_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		\wishbone_TxPointerMSB_reg[31]/NET0131 ,
		_w12577_,
		_w18029_
	);
	LUT2 #(
		.INIT('h4)
	) name7518 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w12608_,
		_w18030_
	);
	LUT2 #(
		.INIT('h2)
	) name7519 (
		_w12621_,
		_w18030_,
		_w18031_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		_w12623_,
		_w18031_,
		_w18032_
	);
	LUT2 #(
		.INIT('h1)
	) name7521 (
		\m_wb_adr_o[31]_pad ,
		_w12606_,
		_w18033_
	);
	LUT2 #(
		.INIT('h8)
	) name7522 (
		\m_wb_adr_o[31]_pad ,
		_w12606_,
		_w18034_
	);
	LUT2 #(
		.INIT('h1)
	) name7523 (
		_w18032_,
		_w18033_,
		_w18035_
	);
	LUT2 #(
		.INIT('h4)
	) name7524 (
		_w18034_,
		_w18035_,
		_w18036_
	);
	LUT2 #(
		.INIT('h1)
	) name7525 (
		_w18027_,
		_w18028_,
		_w18037_
	);
	LUT2 #(
		.INIT('h4)
	) name7526 (
		_w18029_,
		_w18037_,
		_w18038_
	);
	LUT2 #(
		.INIT('h4)
	) name7527 (
		_w18036_,
		_w18038_,
		_w18039_
	);
	LUT2 #(
		.INIT('h4)
	) name7528 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w12641_,
		_w18040_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w18040_,
		_w18041_
	);
	LUT2 #(
		.INIT('h4)
	) name7530 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w18042_
	);
	LUT2 #(
		.INIT('h8)
	) name7531 (
		_w11908_,
		_w18042_,
		_w18043_
	);
	LUT2 #(
		.INIT('h8)
	) name7532 (
		_w11836_,
		_w18043_,
		_w18044_
	);
	LUT2 #(
		.INIT('h8)
	) name7533 (
		_w12641_,
		_w18044_,
		_w18045_
	);
	LUT2 #(
		.INIT('h1)
	) name7534 (
		_w18041_,
		_w18045_,
		_w18046_
	);
	LUT2 #(
		.INIT('h2)
	) name7535 (
		\maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 ,
		_w18046_,
		_w18047_
	);
	LUT2 #(
		.INIT('h8)
	) name7536 (
		_w11831_,
		_w11832_,
		_w18048_
	);
	LUT2 #(
		.INIT('h8)
	) name7537 (
		_w18042_,
		_w18048_,
		_w18049_
	);
	LUT2 #(
		.INIT('h8)
	) name7538 (
		_w11872_,
		_w18049_,
		_w18050_
	);
	LUT2 #(
		.INIT('h8)
	) name7539 (
		_w12641_,
		_w18050_,
		_w18051_
	);
	LUT2 #(
		.INIT('h1)
	) name7540 (
		_w18047_,
		_w18051_,
		_w18052_
	);
	LUT2 #(
		.INIT('h8)
	) name7541 (
		\wishbone_bd_ram_mem2_reg[211][18]/P0001 ,
		_w13166_,
		_w18053_
	);
	LUT2 #(
		.INIT('h8)
	) name7542 (
		\wishbone_bd_ram_mem2_reg[200][18]/P0001 ,
		_w12988_,
		_w18054_
	);
	LUT2 #(
		.INIT('h8)
	) name7543 (
		\wishbone_bd_ram_mem2_reg[96][18]/P0001 ,
		_w12912_,
		_w18055_
	);
	LUT2 #(
		.INIT('h8)
	) name7544 (
		\wishbone_bd_ram_mem2_reg[5][18]/P0001 ,
		_w12878_,
		_w18056_
	);
	LUT2 #(
		.INIT('h8)
	) name7545 (
		\wishbone_bd_ram_mem2_reg[156][18]/P0001 ,
		_w13190_,
		_w18057_
	);
	LUT2 #(
		.INIT('h8)
	) name7546 (
		\wishbone_bd_ram_mem2_reg[37][18]/P0001 ,
		_w13102_,
		_w18058_
	);
	LUT2 #(
		.INIT('h8)
	) name7547 (
		\wishbone_bd_ram_mem2_reg[88][18]/P0001 ,
		_w12860_,
		_w18059_
	);
	LUT2 #(
		.INIT('h8)
	) name7548 (
		\wishbone_bd_ram_mem2_reg[252][18]/P0001 ,
		_w13080_,
		_w18060_
	);
	LUT2 #(
		.INIT('h8)
	) name7549 (
		\wishbone_bd_ram_mem2_reg[95][18]/P0001 ,
		_w12844_,
		_w18061_
	);
	LUT2 #(
		.INIT('h8)
	) name7550 (
		\wishbone_bd_ram_mem2_reg[101][18]/P0001 ,
		_w13192_,
		_w18062_
	);
	LUT2 #(
		.INIT('h8)
	) name7551 (
		\wishbone_bd_ram_mem2_reg[89][18]/P0001 ,
		_w12964_,
		_w18063_
	);
	LUT2 #(
		.INIT('h8)
	) name7552 (
		\wishbone_bd_ram_mem2_reg[172][18]/P0001 ,
		_w12944_,
		_w18064_
	);
	LUT2 #(
		.INIT('h8)
	) name7553 (
		\wishbone_bd_ram_mem2_reg[68][18]/P0001 ,
		_w12946_,
		_w18065_
	);
	LUT2 #(
		.INIT('h8)
	) name7554 (
		\wishbone_bd_ram_mem2_reg[76][18]/P0001 ,
		_w13184_,
		_w18066_
	);
	LUT2 #(
		.INIT('h8)
	) name7555 (
		\wishbone_bd_ram_mem2_reg[125][18]/P0001 ,
		_w12956_,
		_w18067_
	);
	LUT2 #(
		.INIT('h8)
	) name7556 (
		\wishbone_bd_ram_mem2_reg[163][18]/P0001 ,
		_w12882_,
		_w18068_
	);
	LUT2 #(
		.INIT('h8)
	) name7557 (
		\wishbone_bd_ram_mem2_reg[113][18]/P0001 ,
		_w13026_,
		_w18069_
	);
	LUT2 #(
		.INIT('h8)
	) name7558 (
		\wishbone_bd_ram_mem2_reg[134][18]/P0001 ,
		_w12763_,
		_w18070_
	);
	LUT2 #(
		.INIT('h8)
	) name7559 (
		\wishbone_bd_ram_mem2_reg[47][18]/P0001 ,
		_w12904_,
		_w18071_
	);
	LUT2 #(
		.INIT('h8)
	) name7560 (
		\wishbone_bd_ram_mem2_reg[153][18]/P0001 ,
		_w12890_,
		_w18072_
	);
	LUT2 #(
		.INIT('h8)
	) name7561 (
		\wishbone_bd_ram_mem2_reg[16][18]/P0001 ,
		_w13140_,
		_w18073_
	);
	LUT2 #(
		.INIT('h8)
	) name7562 (
		\wishbone_bd_ram_mem2_reg[167][18]/P0001 ,
		_w12986_,
		_w18074_
	);
	LUT2 #(
		.INIT('h8)
	) name7563 (
		\wishbone_bd_ram_mem2_reg[120][18]/P0001 ,
		_w12707_,
		_w18075_
	);
	LUT2 #(
		.INIT('h8)
	) name7564 (
		\wishbone_bd_ram_mem2_reg[247][18]/P0001 ,
		_w12818_,
		_w18076_
	);
	LUT2 #(
		.INIT('h8)
	) name7565 (
		\wishbone_bd_ram_mem2_reg[75][18]/P0001 ,
		_w12826_,
		_w18077_
	);
	LUT2 #(
		.INIT('h8)
	) name7566 (
		\wishbone_bd_ram_mem2_reg[39][18]/P0001 ,
		_w13018_,
		_w18078_
	);
	LUT2 #(
		.INIT('h8)
	) name7567 (
		\wishbone_bd_ram_mem2_reg[2][18]/P0001 ,
		_w13088_,
		_w18079_
	);
	LUT2 #(
		.INIT('h8)
	) name7568 (
		\wishbone_bd_ram_mem2_reg[111][18]/P0001 ,
		_w12744_,
		_w18080_
	);
	LUT2 #(
		.INIT('h8)
	) name7569 (
		\wishbone_bd_ram_mem2_reg[216][18]/P0001 ,
		_w13028_,
		_w18081_
	);
	LUT2 #(
		.INIT('h8)
	) name7570 (
		\wishbone_bd_ram_mem2_reg[238][18]/P0001 ,
		_w13160_,
		_w18082_
	);
	LUT2 #(
		.INIT('h8)
	) name7571 (
		\wishbone_bd_ram_mem2_reg[87][18]/P0001 ,
		_w13154_,
		_w18083_
	);
	LUT2 #(
		.INIT('h8)
	) name7572 (
		\wishbone_bd_ram_mem2_reg[38][18]/P0001 ,
		_w13182_,
		_w18084_
	);
	LUT2 #(
		.INIT('h8)
	) name7573 (
		\wishbone_bd_ram_mem2_reg[232][18]/P0001 ,
		_w12758_,
		_w18085_
	);
	LUT2 #(
		.INIT('h8)
	) name7574 (
		\wishbone_bd_ram_mem2_reg[70][18]/P0001 ,
		_w12840_,
		_w18086_
	);
	LUT2 #(
		.INIT('h8)
	) name7575 (
		\wishbone_bd_ram_mem2_reg[59][18]/P0001 ,
		_w12780_,
		_w18087_
	);
	LUT2 #(
		.INIT('h8)
	) name7576 (
		\wishbone_bd_ram_mem2_reg[169][18]/P0001 ,
		_w12722_,
		_w18088_
	);
	LUT2 #(
		.INIT('h8)
	) name7577 (
		\wishbone_bd_ram_mem2_reg[20][18]/P0001 ,
		_w13174_,
		_w18089_
	);
	LUT2 #(
		.INIT('h8)
	) name7578 (
		\wishbone_bd_ram_mem2_reg[123][18]/P0001 ,
		_w13114_,
		_w18090_
	);
	LUT2 #(
		.INIT('h8)
	) name7579 (
		\wishbone_bd_ram_mem2_reg[122][18]/P0001 ,
		_w13130_,
		_w18091_
	);
	LUT2 #(
		.INIT('h8)
	) name7580 (
		\wishbone_bd_ram_mem2_reg[162][18]/P0001 ,
		_w13098_,
		_w18092_
	);
	LUT2 #(
		.INIT('h8)
	) name7581 (
		\wishbone_bd_ram_mem2_reg[34][18]/P0001 ,
		_w12930_,
		_w18093_
	);
	LUT2 #(
		.INIT('h8)
	) name7582 (
		\wishbone_bd_ram_mem2_reg[207][18]/P0001 ,
		_w13180_,
		_w18094_
	);
	LUT2 #(
		.INIT('h8)
	) name7583 (
		\wishbone_bd_ram_mem2_reg[127][18]/P0001 ,
		_w13164_,
		_w18095_
	);
	LUT2 #(
		.INIT('h8)
	) name7584 (
		\wishbone_bd_ram_mem2_reg[166][18]/P0001 ,
		_w13040_,
		_w18096_
	);
	LUT2 #(
		.INIT('h8)
	) name7585 (
		\wishbone_bd_ram_mem2_reg[149][18]/P0001 ,
		_w12741_,
		_w18097_
	);
	LUT2 #(
		.INIT('h8)
	) name7586 (
		\wishbone_bd_ram_mem2_reg[100][18]/P0001 ,
		_w12960_,
		_w18098_
	);
	LUT2 #(
		.INIT('h8)
	) name7587 (
		\wishbone_bd_ram_mem2_reg[226][18]/P0001 ,
		_w13138_,
		_w18099_
	);
	LUT2 #(
		.INIT('h8)
	) name7588 (
		\wishbone_bd_ram_mem2_reg[196][18]/P0001 ,
		_w13090_,
		_w18100_
	);
	LUT2 #(
		.INIT('h8)
	) name7589 (
		\wishbone_bd_ram_mem2_reg[114][18]/P0001 ,
		_w13202_,
		_w18101_
	);
	LUT2 #(
		.INIT('h8)
	) name7590 (
		\wishbone_bd_ram_mem2_reg[91][18]/P0001 ,
		_w13074_,
		_w18102_
	);
	LUT2 #(
		.INIT('h8)
	) name7591 (
		\wishbone_bd_ram_mem2_reg[151][18]/P0001 ,
		_w13142_,
		_w18103_
	);
	LUT2 #(
		.INIT('h8)
	) name7592 (
		\wishbone_bd_ram_mem2_reg[244][18]/P0001 ,
		_w12747_,
		_w18104_
	);
	LUT2 #(
		.INIT('h8)
	) name7593 (
		\wishbone_bd_ram_mem2_reg[41][18]/P0001 ,
		_w13052_,
		_w18105_
	);
	LUT2 #(
		.INIT('h8)
	) name7594 (
		\wishbone_bd_ram_mem2_reg[97][18]/P0001 ,
		_w13096_,
		_w18106_
	);
	LUT2 #(
		.INIT('h8)
	) name7595 (
		\wishbone_bd_ram_mem2_reg[160][18]/P0001 ,
		_w12872_,
		_w18107_
	);
	LUT2 #(
		.INIT('h8)
	) name7596 (
		\wishbone_bd_ram_mem2_reg[0][18]/P0001 ,
		_w12717_,
		_w18108_
	);
	LUT2 #(
		.INIT('h8)
	) name7597 (
		\wishbone_bd_ram_mem2_reg[9][18]/P0001 ,
		_w12808_,
		_w18109_
	);
	LUT2 #(
		.INIT('h8)
	) name7598 (
		\wishbone_bd_ram_mem2_reg[25][18]/P0001 ,
		_w13108_,
		_w18110_
	);
	LUT2 #(
		.INIT('h8)
	) name7599 (
		\wishbone_bd_ram_mem2_reg[201][18]/P0001 ,
		_w12822_,
		_w18111_
	);
	LUT2 #(
		.INIT('h8)
	) name7600 (
		\wishbone_bd_ram_mem2_reg[250][18]/P0001 ,
		_w13128_,
		_w18112_
	);
	LUT2 #(
		.INIT('h8)
	) name7601 (
		\wishbone_bd_ram_mem2_reg[208][18]/P0001 ,
		_w13032_,
		_w18113_
	);
	LUT2 #(
		.INIT('h8)
	) name7602 (
		\wishbone_bd_ram_mem2_reg[121][18]/P0001 ,
		_w13078_,
		_w18114_
	);
	LUT2 #(
		.INIT('h8)
	) name7603 (
		\wishbone_bd_ram_mem2_reg[187][18]/P0001 ,
		_w13196_,
		_w18115_
	);
	LUT2 #(
		.INIT('h8)
	) name7604 (
		\wishbone_bd_ram_mem2_reg[131][18]/P0001 ,
		_w12852_,
		_w18116_
	);
	LUT2 #(
		.INIT('h8)
	) name7605 (
		\wishbone_bd_ram_mem2_reg[14][18]/P0001 ,
		_w13086_,
		_w18117_
	);
	LUT2 #(
		.INIT('h8)
	) name7606 (
		\wishbone_bd_ram_mem2_reg[61][18]/P0001 ,
		_w12725_,
		_w18118_
	);
	LUT2 #(
		.INIT('h8)
	) name7607 (
		\wishbone_bd_ram_mem2_reg[234][18]/P0001 ,
		_w13214_,
		_w18119_
	);
	LUT2 #(
		.INIT('h8)
	) name7608 (
		\wishbone_bd_ram_mem2_reg[4][18]/P0001 ,
		_w12666_,
		_w18120_
	);
	LUT2 #(
		.INIT('h8)
	) name7609 (
		\wishbone_bd_ram_mem2_reg[40][18]/P0001 ,
		_w13132_,
		_w18121_
	);
	LUT2 #(
		.INIT('h8)
	) name7610 (
		\wishbone_bd_ram_mem2_reg[42][18]/P0001 ,
		_w12842_,
		_w18122_
	);
	LUT2 #(
		.INIT('h8)
	) name7611 (
		\wishbone_bd_ram_mem2_reg[179][18]/P0001 ,
		_w13050_,
		_w18123_
	);
	LUT2 #(
		.INIT('h8)
	) name7612 (
		\wishbone_bd_ram_mem2_reg[210][18]/P0001 ,
		_w12924_,
		_w18124_
	);
	LUT2 #(
		.INIT('h8)
	) name7613 (
		\wishbone_bd_ram_mem2_reg[146][18]/P0001 ,
		_w13060_,
		_w18125_
	);
	LUT2 #(
		.INIT('h8)
	) name7614 (
		\wishbone_bd_ram_mem2_reg[65][18]/P0001 ,
		_w13176_,
		_w18126_
	);
	LUT2 #(
		.INIT('h8)
	) name7615 (
		\wishbone_bd_ram_mem2_reg[13][18]/P0001 ,
		_w13178_,
		_w18127_
	);
	LUT2 #(
		.INIT('h8)
	) name7616 (
		\wishbone_bd_ram_mem2_reg[10][18]/P0001 ,
		_w13172_,
		_w18128_
	);
	LUT2 #(
		.INIT('h8)
	) name7617 (
		\wishbone_bd_ram_mem2_reg[80][18]/P0001 ,
		_w12689_,
		_w18129_
	);
	LUT2 #(
		.INIT('h8)
	) name7618 (
		\wishbone_bd_ram_mem2_reg[99][18]/P0001 ,
		_w13038_,
		_w18130_
	);
	LUT2 #(
		.INIT('h8)
	) name7619 (
		\wishbone_bd_ram_mem2_reg[159][18]/P0001 ,
		_w12774_,
		_w18131_
	);
	LUT2 #(
		.INIT('h8)
	) name7620 (
		\wishbone_bd_ram_mem2_reg[107][18]/P0001 ,
		_w12749_,
		_w18132_
	);
	LUT2 #(
		.INIT('h8)
	) name7621 (
		\wishbone_bd_ram_mem2_reg[221][18]/P0001 ,
		_w12802_,
		_w18133_
	);
	LUT2 #(
		.INIT('h8)
	) name7622 (
		\wishbone_bd_ram_mem2_reg[55][18]/P0001 ,
		_w12785_,
		_w18134_
	);
	LUT2 #(
		.INIT('h8)
	) name7623 (
		\wishbone_bd_ram_mem2_reg[102][18]/P0001 ,
		_w12685_,
		_w18135_
	);
	LUT2 #(
		.INIT('h8)
	) name7624 (
		\wishbone_bd_ram_mem2_reg[157][18]/P0001 ,
		_w12926_,
		_w18136_
	);
	LUT2 #(
		.INIT('h8)
	) name7625 (
		\wishbone_bd_ram_mem2_reg[85][18]/P0001 ,
		_w13216_,
		_w18137_
	);
	LUT2 #(
		.INIT('h8)
	) name7626 (
		\wishbone_bd_ram_mem2_reg[106][18]/P0001 ,
		_w12713_,
		_w18138_
	);
	LUT2 #(
		.INIT('h8)
	) name7627 (
		\wishbone_bd_ram_mem2_reg[197][18]/P0001 ,
		_w12834_,
		_w18139_
	);
	LUT2 #(
		.INIT('h8)
	) name7628 (
		\wishbone_bd_ram_mem2_reg[176][18]/P0001 ,
		_w12868_,
		_w18140_
	);
	LUT2 #(
		.INIT('h8)
	) name7629 (
		\wishbone_bd_ram_mem2_reg[6][18]/P0001 ,
		_w12968_,
		_w18141_
	);
	LUT2 #(
		.INIT('h8)
	) name7630 (
		\wishbone_bd_ram_mem2_reg[222][18]/P0001 ,
		_w13094_,
		_w18142_
	);
	LUT2 #(
		.INIT('h8)
	) name7631 (
		\wishbone_bd_ram_mem2_reg[32][18]/P0001 ,
		_w13120_,
		_w18143_
	);
	LUT2 #(
		.INIT('h8)
	) name7632 (
		\wishbone_bd_ram_mem2_reg[119][18]/P0001 ,
		_w13048_,
		_w18144_
	);
	LUT2 #(
		.INIT('h8)
	) name7633 (
		\wishbone_bd_ram_mem2_reg[7][18]/P0001 ,
		_w12728_,
		_w18145_
	);
	LUT2 #(
		.INIT('h8)
	) name7634 (
		\wishbone_bd_ram_mem2_reg[3][18]/P0001 ,
		_w12866_,
		_w18146_
	);
	LUT2 #(
		.INIT('h8)
	) name7635 (
		\wishbone_bd_ram_mem2_reg[191][18]/P0001 ,
		_w13034_,
		_w18147_
	);
	LUT2 #(
		.INIT('h8)
	) name7636 (
		\wishbone_bd_ram_mem2_reg[254][18]/P0001 ,
		_w12892_,
		_w18148_
	);
	LUT2 #(
		.INIT('h8)
	) name7637 (
		\wishbone_bd_ram_mem2_reg[48][18]/P0001 ,
		_w12970_,
		_w18149_
	);
	LUT2 #(
		.INIT('h8)
	) name7638 (
		\wishbone_bd_ram_mem2_reg[43][18]/P0001 ,
		_w13200_,
		_w18150_
	);
	LUT2 #(
		.INIT('h8)
	) name7639 (
		\wishbone_bd_ram_mem2_reg[230][18]/P0001 ,
		_w13036_,
		_w18151_
	);
	LUT2 #(
		.INIT('h8)
	) name7640 (
		\wishbone_bd_ram_mem2_reg[242][18]/P0001 ,
		_w12932_,
		_w18152_
	);
	LUT2 #(
		.INIT('h8)
	) name7641 (
		\wishbone_bd_ram_mem2_reg[195][18]/P0001 ,
		_w13144_,
		_w18153_
	);
	LUT2 #(
		.INIT('h8)
	) name7642 (
		\wishbone_bd_ram_mem2_reg[103][18]/P0001 ,
		_w12846_,
		_w18154_
	);
	LUT2 #(
		.INIT('h8)
	) name7643 (
		\wishbone_bd_ram_mem2_reg[86][18]/P0001 ,
		_w12735_,
		_w18155_
	);
	LUT2 #(
		.INIT('h8)
	) name7644 (
		\wishbone_bd_ram_mem2_reg[170][18]/P0001 ,
		_w13030_,
		_w18156_
	);
	LUT2 #(
		.INIT('h8)
	) name7645 (
		\wishbone_bd_ram_mem2_reg[251][18]/P0001 ,
		_w13054_,
		_w18157_
	);
	LUT2 #(
		.INIT('h8)
	) name7646 (
		\wishbone_bd_ram_mem2_reg[206][18]/P0001 ,
		_w12954_,
		_w18158_
	);
	LUT2 #(
		.INIT('h8)
	) name7647 (
		\wishbone_bd_ram_mem2_reg[224][18]/P0001 ,
		_w12902_,
		_w18159_
	);
	LUT2 #(
		.INIT('h8)
	) name7648 (
		\wishbone_bd_ram_mem2_reg[185][18]/P0001 ,
		_w12940_,
		_w18160_
	);
	LUT2 #(
		.INIT('h8)
	) name7649 (
		\wishbone_bd_ram_mem2_reg[178][18]/P0001 ,
		_w12886_,
		_w18161_
	);
	LUT2 #(
		.INIT('h8)
	) name7650 (
		\wishbone_bd_ram_mem2_reg[29][18]/P0001 ,
		_w12952_,
		_w18162_
	);
	LUT2 #(
		.INIT('h8)
	) name7651 (
		\wishbone_bd_ram_mem2_reg[229][18]/P0001 ,
		_w12711_,
		_w18163_
	);
	LUT2 #(
		.INIT('h8)
	) name7652 (
		\wishbone_bd_ram_mem2_reg[130][18]/P0001 ,
		_w12914_,
		_w18164_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		\wishbone_bd_ram_mem2_reg[79][18]/P0001 ,
		_w13212_,
		_w18165_
	);
	LUT2 #(
		.INIT('h8)
	) name7654 (
		\wishbone_bd_ram_mem2_reg[90][18]/P0001 ,
		_w12978_,
		_w18166_
	);
	LUT2 #(
		.INIT('h8)
	) name7655 (
		\wishbone_bd_ram_mem2_reg[45][18]/P0001 ,
		_w12908_,
		_w18167_
	);
	LUT2 #(
		.INIT('h8)
	) name7656 (
		\wishbone_bd_ram_mem2_reg[128][18]/P0001 ,
		_w12793_,
		_w18168_
	);
	LUT2 #(
		.INIT('h8)
	) name7657 (
		\wishbone_bd_ram_mem2_reg[12][18]/P0001 ,
		_w13118_,
		_w18169_
	);
	LUT2 #(
		.INIT('h8)
	) name7658 (
		\wishbone_bd_ram_mem2_reg[184][18]/P0001 ,
		_w13062_,
		_w18170_
	);
	LUT2 #(
		.INIT('h8)
	) name7659 (
		\wishbone_bd_ram_mem2_reg[82][18]/P0001 ,
		_w12942_,
		_w18171_
	);
	LUT2 #(
		.INIT('h8)
	) name7660 (
		\wishbone_bd_ram_mem2_reg[174][18]/P0001 ,
		_w12972_,
		_w18172_
	);
	LUT2 #(
		.INIT('h8)
	) name7661 (
		\wishbone_bd_ram_mem2_reg[11][18]/P0001 ,
		_w13194_,
		_w18173_
	);
	LUT2 #(
		.INIT('h8)
	) name7662 (
		\wishbone_bd_ram_mem2_reg[218][18]/P0001 ,
		_w13206_,
		_w18174_
	);
	LUT2 #(
		.INIT('h8)
	) name7663 (
		\wishbone_bd_ram_mem2_reg[126][18]/P0001 ,
		_w13218_,
		_w18175_
	);
	LUT2 #(
		.INIT('h8)
	) name7664 (
		\wishbone_bd_ram_mem2_reg[115][18]/P0001 ,
		_w13112_,
		_w18176_
	);
	LUT2 #(
		.INIT('h8)
	) name7665 (
		\wishbone_bd_ram_mem2_reg[84][18]/P0001 ,
		_w12934_,
		_w18177_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		\wishbone_bd_ram_mem2_reg[193][18]/P0001 ,
		_w13056_,
		_w18178_
	);
	LUT2 #(
		.INIT('h8)
	) name7667 (
		\wishbone_bd_ram_mem2_reg[241][18]/P0001 ,
		_w13006_,
		_w18179_
	);
	LUT2 #(
		.INIT('h8)
	) name7668 (
		\wishbone_bd_ram_mem2_reg[138][18]/P0001 ,
		_w12958_,
		_w18180_
	);
	LUT2 #(
		.INIT('h8)
	) name7669 (
		\wishbone_bd_ram_mem2_reg[231][18]/P0001 ,
		_w12856_,
		_w18181_
	);
	LUT2 #(
		.INIT('h8)
	) name7670 (
		\wishbone_bd_ram_mem2_reg[136][18]/P0001 ,
		_w13064_,
		_w18182_
	);
	LUT2 #(
		.INIT('h8)
	) name7671 (
		\wishbone_bd_ram_mem2_reg[225][18]/P0001 ,
		_w13092_,
		_w18183_
	);
	LUT2 #(
		.INIT('h8)
	) name7672 (
		\wishbone_bd_ram_mem2_reg[81][18]/P0001 ,
		_w12950_,
		_w18184_
	);
	LUT2 #(
		.INIT('h8)
	) name7673 (
		\wishbone_bd_ram_mem2_reg[220][18]/P0001 ,
		_w13066_,
		_w18185_
	);
	LUT2 #(
		.INIT('h8)
	) name7674 (
		\wishbone_bd_ram_mem2_reg[51][18]/P0001 ,
		_w13024_,
		_w18186_
	);
	LUT2 #(
		.INIT('h8)
	) name7675 (
		\wishbone_bd_ram_mem2_reg[60][18]/P0001 ,
		_w13204_,
		_w18187_
	);
	LUT2 #(
		.INIT('h8)
	) name7676 (
		\wishbone_bd_ram_mem2_reg[148][18]/P0001 ,
		_w13000_,
		_w18188_
	);
	LUT2 #(
		.INIT('h8)
	) name7677 (
		\wishbone_bd_ram_mem2_reg[243][18]/P0001 ,
		_w12804_,
		_w18189_
	);
	LUT2 #(
		.INIT('h8)
	) name7678 (
		\wishbone_bd_ram_mem2_reg[236][18]/P0001 ,
		_w12731_,
		_w18190_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		\wishbone_bd_ram_mem2_reg[73][18]/P0001 ,
		_w12918_,
		_w18191_
	);
	LUT2 #(
		.INIT('h8)
	) name7680 (
		\wishbone_bd_ram_mem2_reg[124][18]/P0001 ,
		_w13058_,
		_w18192_
	);
	LUT2 #(
		.INIT('h8)
	) name7681 (
		\wishbone_bd_ram_mem2_reg[26][18]/P0001 ,
		_w12699_,
		_w18193_
	);
	LUT2 #(
		.INIT('h8)
	) name7682 (
		\wishbone_bd_ram_mem2_reg[22][18]/P0001 ,
		_w13110_,
		_w18194_
	);
	LUT2 #(
		.INIT('h8)
	) name7683 (
		\wishbone_bd_ram_mem2_reg[92][18]/P0001 ,
		_w13010_,
		_w18195_
	);
	LUT2 #(
		.INIT('h8)
	) name7684 (
		\wishbone_bd_ram_mem2_reg[175][18]/P0001 ,
		_w13126_,
		_w18196_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		\wishbone_bd_ram_mem2_reg[144][18]/P0001 ,
		_w12756_,
		_w18197_
	);
	LUT2 #(
		.INIT('h8)
	) name7686 (
		\wishbone_bd_ram_mem2_reg[248][18]/P0001 ,
		_w12789_,
		_w18198_
	);
	LUT2 #(
		.INIT('h8)
	) name7687 (
		\wishbone_bd_ram_mem2_reg[135][18]/P0001 ,
		_w13124_,
		_w18199_
	);
	LUT2 #(
		.INIT('h8)
	) name7688 (
		\wishbone_bd_ram_mem2_reg[150][18]/P0001 ,
		_w13136_,
		_w18200_
	);
	LUT2 #(
		.INIT('h8)
	) name7689 (
		\wishbone_bd_ram_mem2_reg[203][18]/P0001 ,
		_w13158_,
		_w18201_
	);
	LUT2 #(
		.INIT('h8)
	) name7690 (
		\wishbone_bd_ram_mem2_reg[129][18]/P0001 ,
		_w12776_,
		_w18202_
	);
	LUT2 #(
		.INIT('h8)
	) name7691 (
		\wishbone_bd_ram_mem2_reg[246][18]/P0001 ,
		_w13076_,
		_w18203_
	);
	LUT2 #(
		.INIT('h8)
	) name7692 (
		\wishbone_bd_ram_mem2_reg[245][18]/P0001 ,
		_w13022_,
		_w18204_
	);
	LUT2 #(
		.INIT('h8)
	) name7693 (
		\wishbone_bd_ram_mem2_reg[35][18]/P0001 ,
		_w12703_,
		_w18205_
	);
	LUT2 #(
		.INIT('h8)
	) name7694 (
		\wishbone_bd_ram_mem2_reg[255][18]/P0001 ,
		_w13072_,
		_w18206_
	);
	LUT2 #(
		.INIT('h8)
	) name7695 (
		\wishbone_bd_ram_mem2_reg[54][18]/P0001 ,
		_w12770_,
		_w18207_
	);
	LUT2 #(
		.INIT('h8)
	) name7696 (
		\wishbone_bd_ram_mem2_reg[180][18]/P0001 ,
		_w12791_,
		_w18208_
	);
	LUT2 #(
		.INIT('h8)
	) name7697 (
		\wishbone_bd_ram_mem2_reg[215][18]/P0001 ,
		_w12974_,
		_w18209_
	);
	LUT2 #(
		.INIT('h8)
	) name7698 (
		\wishbone_bd_ram_mem2_reg[181][18]/P0001 ,
		_w12828_,
		_w18210_
	);
	LUT2 #(
		.INIT('h8)
	) name7699 (
		\wishbone_bd_ram_mem2_reg[190][18]/P0001 ,
		_w12858_,
		_w18211_
	);
	LUT2 #(
		.INIT('h8)
	) name7700 (
		\wishbone_bd_ram_mem2_reg[161][18]/P0001 ,
		_w12754_,
		_w18212_
	);
	LUT2 #(
		.INIT('h8)
	) name7701 (
		\wishbone_bd_ram_mem2_reg[213][18]/P0001 ,
		_w13002_,
		_w18213_
	);
	LUT2 #(
		.INIT('h8)
	) name7702 (
		\wishbone_bd_ram_mem2_reg[212][18]/P0001 ,
		_w12796_,
		_w18214_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		\wishbone_bd_ram_mem2_reg[63][18]/P0001 ,
		_w12850_,
		_w18215_
	);
	LUT2 #(
		.INIT('h8)
	) name7704 (
		\wishbone_bd_ram_mem2_reg[17][18]/P0001 ,
		_w12848_,
		_w18216_
	);
	LUT2 #(
		.INIT('h8)
	) name7705 (
		\wishbone_bd_ram_mem2_reg[98][18]/P0001 ,
		_w12816_,
		_w18217_
	);
	LUT2 #(
		.INIT('h8)
	) name7706 (
		\wishbone_bd_ram_mem2_reg[228][18]/P0001 ,
		_w12765_,
		_w18218_
	);
	LUT2 #(
		.INIT('h8)
	) name7707 (
		\wishbone_bd_ram_mem2_reg[69][18]/P0001 ,
		_w12738_,
		_w18219_
	);
	LUT2 #(
		.INIT('h8)
	) name7708 (
		\wishbone_bd_ram_mem2_reg[44][18]/P0001 ,
		_w12896_,
		_w18220_
	);
	LUT2 #(
		.INIT('h8)
	) name7709 (
		\wishbone_bd_ram_mem2_reg[168][18]/P0001 ,
		_w13208_,
		_w18221_
	);
	LUT2 #(
		.INIT('h8)
	) name7710 (
		\wishbone_bd_ram_mem2_reg[109][18]/P0001 ,
		_w12888_,
		_w18222_
	);
	LUT2 #(
		.INIT('h8)
	) name7711 (
		\wishbone_bd_ram_mem2_reg[182][18]/P0001 ,
		_w12820_,
		_w18223_
	);
	LUT2 #(
		.INIT('h8)
	) name7712 (
		\wishbone_bd_ram_mem2_reg[58][18]/P0001 ,
		_w13070_,
		_w18224_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		\wishbone_bd_ram_mem2_reg[253][18]/P0001 ,
		_w13100_,
		_w18225_
	);
	LUT2 #(
		.INIT('h8)
	) name7714 (
		\wishbone_bd_ram_mem2_reg[147][18]/P0001 ,
		_w13146_,
		_w18226_
	);
	LUT2 #(
		.INIT('h8)
	) name7715 (
		\wishbone_bd_ram_mem2_reg[28][18]/P0001 ,
		_w13170_,
		_w18227_
	);
	LUT2 #(
		.INIT('h8)
	) name7716 (
		\wishbone_bd_ram_mem2_reg[15][18]/P0001 ,
		_w13210_,
		_w18228_
	);
	LUT2 #(
		.INIT('h8)
	) name7717 (
		\wishbone_bd_ram_mem2_reg[118][18]/P0001 ,
		_w12830_,
		_w18229_
	);
	LUT2 #(
		.INIT('h8)
	) name7718 (
		\wishbone_bd_ram_mem2_reg[227][18]/P0001 ,
		_w12936_,
		_w18230_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		\wishbone_bd_ram_mem2_reg[112][18]/P0001 ,
		_w12733_,
		_w18231_
	);
	LUT2 #(
		.INIT('h8)
	) name7720 (
		\wishbone_bd_ram_mem2_reg[189][18]/P0001 ,
		_w13042_,
		_w18232_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		\wishbone_bd_ram_mem2_reg[141][18]/P0001 ,
		_w13004_,
		_w18233_
	);
	LUT2 #(
		.INIT('h8)
	) name7722 (
		\wishbone_bd_ram_mem2_reg[171][18]/P0001 ,
		_w12910_,
		_w18234_
	);
	LUT2 #(
		.INIT('h8)
	) name7723 (
		\wishbone_bd_ram_mem2_reg[164][18]/P0001 ,
		_w12876_,
		_w18235_
	);
	LUT2 #(
		.INIT('h8)
	) name7724 (
		\wishbone_bd_ram_mem2_reg[237][18]/P0001 ,
		_w12990_,
		_w18236_
	);
	LUT2 #(
		.INIT('h8)
	) name7725 (
		\wishbone_bd_ram_mem2_reg[142][18]/P0001 ,
		_w12928_,
		_w18237_
	);
	LUT2 #(
		.INIT('h8)
	) name7726 (
		\wishbone_bd_ram_mem2_reg[77][18]/P0001 ,
		_w12982_,
		_w18238_
	);
	LUT2 #(
		.INIT('h8)
	) name7727 (
		\wishbone_bd_ram_mem2_reg[83][18]/P0001 ,
		_w12916_,
		_w18239_
	);
	LUT2 #(
		.INIT('h8)
	) name7728 (
		\wishbone_bd_ram_mem2_reg[56][18]/P0001 ,
		_w12778_,
		_w18240_
	);
	LUT2 #(
		.INIT('h8)
	) name7729 (
		\wishbone_bd_ram_mem2_reg[223][18]/P0001 ,
		_w12838_,
		_w18241_
	);
	LUT2 #(
		.INIT('h8)
	) name7730 (
		\wishbone_bd_ram_mem2_reg[249][18]/P0001 ,
		_w12900_,
		_w18242_
	);
	LUT2 #(
		.INIT('h8)
	) name7731 (
		\wishbone_bd_ram_mem2_reg[173][18]/P0001 ,
		_w12854_,
		_w18243_
	);
	LUT2 #(
		.INIT('h8)
	) name7732 (
		\wishbone_bd_ram_mem2_reg[66][18]/P0001 ,
		_w12824_,
		_w18244_
	);
	LUT2 #(
		.INIT('h8)
	) name7733 (
		\wishbone_bd_ram_mem2_reg[165][18]/P0001 ,
		_w13044_,
		_w18245_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		\wishbone_bd_ram_mem2_reg[105][18]/P0001 ,
		_w12751_,
		_w18246_
	);
	LUT2 #(
		.INIT('h8)
	) name7735 (
		\wishbone_bd_ram_mem2_reg[46][18]/P0001 ,
		_w12884_,
		_w18247_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		\wishbone_bd_ram_mem2_reg[93][18]/P0001 ,
		_w13016_,
		_w18248_
	);
	LUT2 #(
		.INIT('h8)
	) name7737 (
		\wishbone_bd_ram_mem2_reg[240][18]/P0001 ,
		_w12864_,
		_w18249_
	);
	LUT2 #(
		.INIT('h8)
	) name7738 (
		\wishbone_bd_ram_mem2_reg[143][18]/P0001 ,
		_w12922_,
		_w18250_
	);
	LUT2 #(
		.INIT('h8)
	) name7739 (
		\wishbone_bd_ram_mem2_reg[24][18]/P0001 ,
		_w13084_,
		_w18251_
	);
	LUT2 #(
		.INIT('h8)
	) name7740 (
		\wishbone_bd_ram_mem2_reg[104][18]/P0001 ,
		_w13148_,
		_w18252_
	);
	LUT2 #(
		.INIT('h8)
	) name7741 (
		\wishbone_bd_ram_mem2_reg[194][18]/P0001 ,
		_w12772_,
		_w18253_
	);
	LUT2 #(
		.INIT('h8)
	) name7742 (
		\wishbone_bd_ram_mem2_reg[71][18]/P0001 ,
		_w12798_,
		_w18254_
	);
	LUT2 #(
		.INIT('h8)
	) name7743 (
		\wishbone_bd_ram_mem2_reg[31][18]/P0001 ,
		_w13198_,
		_w18255_
	);
	LUT2 #(
		.INIT('h8)
	) name7744 (
		\wishbone_bd_ram_mem2_reg[53][18]/P0001 ,
		_w13020_,
		_w18256_
	);
	LUT2 #(
		.INIT('h8)
	) name7745 (
		\wishbone_bd_ram_mem2_reg[209][18]/P0001 ,
		_w13152_,
		_w18257_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		\wishbone_bd_ram_mem2_reg[21][18]/P0001 ,
		_w12906_,
		_w18258_
	);
	LUT2 #(
		.INIT('h8)
	) name7747 (
		\wishbone_bd_ram_mem2_reg[233][18]/P0001 ,
		_w12836_,
		_w18259_
	);
	LUT2 #(
		.INIT('h8)
	) name7748 (
		\wishbone_bd_ram_mem2_reg[186][18]/P0001 ,
		_w12783_,
		_w18260_
	);
	LUT2 #(
		.INIT('h8)
	) name7749 (
		\wishbone_bd_ram_mem2_reg[108][18]/P0001 ,
		_w13156_,
		_w18261_
	);
	LUT2 #(
		.INIT('h8)
	) name7750 (
		\wishbone_bd_ram_mem2_reg[50][18]/P0001 ,
		_w13150_,
		_w18262_
	);
	LUT2 #(
		.INIT('h8)
	) name7751 (
		\wishbone_bd_ram_mem2_reg[139][18]/P0001 ,
		_w12814_,
		_w18263_
	);
	LUT2 #(
		.INIT('h8)
	) name7752 (
		\wishbone_bd_ram_mem2_reg[132][18]/P0001 ,
		_w12992_,
		_w18264_
	);
	LUT2 #(
		.INIT('h8)
	) name7753 (
		\wishbone_bd_ram_mem2_reg[1][18]/P0001 ,
		_w13014_,
		_w18265_
	);
	LUT2 #(
		.INIT('h8)
	) name7754 (
		\wishbone_bd_ram_mem2_reg[33][18]/P0001 ,
		_w12980_,
		_w18266_
	);
	LUT2 #(
		.INIT('h8)
	) name7755 (
		\wishbone_bd_ram_mem2_reg[23][18]/P0001 ,
		_w13008_,
		_w18267_
	);
	LUT2 #(
		.INIT('h8)
	) name7756 (
		\wishbone_bd_ram_mem2_reg[155][18]/P0001 ,
		_w13122_,
		_w18268_
	);
	LUT2 #(
		.INIT('h8)
	) name7757 (
		\wishbone_bd_ram_mem2_reg[205][18]/P0001 ,
		_w13068_,
		_w18269_
	);
	LUT2 #(
		.INIT('h8)
	) name7758 (
		\wishbone_bd_ram_mem2_reg[18][18]/P0001 ,
		_w12679_,
		_w18270_
	);
	LUT2 #(
		.INIT('h8)
	) name7759 (
		\wishbone_bd_ram_mem2_reg[188][18]/P0001 ,
		_w12948_,
		_w18271_
	);
	LUT2 #(
		.INIT('h8)
	) name7760 (
		\wishbone_bd_ram_mem2_reg[198][18]/P0001 ,
		_w12832_,
		_w18272_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		\wishbone_bd_ram_mem2_reg[72][18]/P0001 ,
		_w12810_,
		_w18273_
	);
	LUT2 #(
		.INIT('h8)
	) name7762 (
		\wishbone_bd_ram_mem2_reg[140][18]/P0001 ,
		_w12894_,
		_w18274_
	);
	LUT2 #(
		.INIT('h8)
	) name7763 (
		\wishbone_bd_ram_mem2_reg[67][18]/P0001 ,
		_w13134_,
		_w18275_
	);
	LUT2 #(
		.INIT('h8)
	) name7764 (
		\wishbone_bd_ram_mem2_reg[94][18]/P0001 ,
		_w13186_,
		_w18276_
	);
	LUT2 #(
		.INIT('h8)
	) name7765 (
		\wishbone_bd_ram_mem2_reg[62][18]/P0001 ,
		_w12673_,
		_w18277_
	);
	LUT2 #(
		.INIT('h8)
	) name7766 (
		\wishbone_bd_ram_mem2_reg[57][18]/P0001 ,
		_w13116_,
		_w18278_
	);
	LUT2 #(
		.INIT('h8)
	) name7767 (
		\wishbone_bd_ram_mem2_reg[117][18]/P0001 ,
		_w12715_,
		_w18279_
	);
	LUT2 #(
		.INIT('h8)
	) name7768 (
		\wishbone_bd_ram_mem2_reg[30][18]/P0001 ,
		_w13104_,
		_w18280_
	);
	LUT2 #(
		.INIT('h8)
	) name7769 (
		\wishbone_bd_ram_mem2_reg[145][18]/P0001 ,
		_w13106_,
		_w18281_
	);
	LUT2 #(
		.INIT('h8)
	) name7770 (
		\wishbone_bd_ram_mem2_reg[8][18]/P0001 ,
		_w12920_,
		_w18282_
	);
	LUT2 #(
		.INIT('h8)
	) name7771 (
		\wishbone_bd_ram_mem2_reg[133][18]/P0001 ,
		_w12761_,
		_w18283_
	);
	LUT2 #(
		.INIT('h8)
	) name7772 (
		\wishbone_bd_ram_mem2_reg[202][18]/P0001 ,
		_w12870_,
		_w18284_
	);
	LUT2 #(
		.INIT('h8)
	) name7773 (
		\wishbone_bd_ram_mem2_reg[158][18]/P0001 ,
		_w12898_,
		_w18285_
	);
	LUT2 #(
		.INIT('h8)
	) name7774 (
		\wishbone_bd_ram_mem2_reg[49][18]/P0001 ,
		_w12994_,
		_w18286_
	);
	LUT2 #(
		.INIT('h8)
	) name7775 (
		\wishbone_bd_ram_mem2_reg[204][18]/P0001 ,
		_w13162_,
		_w18287_
	);
	LUT2 #(
		.INIT('h8)
	) name7776 (
		\wishbone_bd_ram_mem2_reg[64][18]/P0001 ,
		_w12976_,
		_w18288_
	);
	LUT2 #(
		.INIT('h8)
	) name7777 (
		\wishbone_bd_ram_mem2_reg[137][18]/P0001 ,
		_w13168_,
		_w18289_
	);
	LUT2 #(
		.INIT('h8)
	) name7778 (
		\wishbone_bd_ram_mem2_reg[177][18]/P0001 ,
		_w12996_,
		_w18290_
	);
	LUT2 #(
		.INIT('h8)
	) name7779 (
		\wishbone_bd_ram_mem2_reg[154][18]/P0001 ,
		_w12962_,
		_w18291_
	);
	LUT2 #(
		.INIT('h8)
	) name7780 (
		\wishbone_bd_ram_mem2_reg[152][18]/P0001 ,
		_w12966_,
		_w18292_
	);
	LUT2 #(
		.INIT('h8)
	) name7781 (
		\wishbone_bd_ram_mem2_reg[74][18]/P0001 ,
		_w12812_,
		_w18293_
	);
	LUT2 #(
		.INIT('h8)
	) name7782 (
		\wishbone_bd_ram_mem2_reg[199][18]/P0001 ,
		_w12768_,
		_w18294_
	);
	LUT2 #(
		.INIT('h8)
	) name7783 (
		\wishbone_bd_ram_mem2_reg[217][18]/P0001 ,
		_w13188_,
		_w18295_
	);
	LUT2 #(
		.INIT('h8)
	) name7784 (
		\wishbone_bd_ram_mem2_reg[214][18]/P0001 ,
		_w12984_,
		_w18296_
	);
	LUT2 #(
		.INIT('h8)
	) name7785 (
		\wishbone_bd_ram_mem2_reg[19][18]/P0001 ,
		_w13012_,
		_w18297_
	);
	LUT2 #(
		.INIT('h8)
	) name7786 (
		\wishbone_bd_ram_mem2_reg[239][18]/P0001 ,
		_w12862_,
		_w18298_
	);
	LUT2 #(
		.INIT('h8)
	) name7787 (
		\wishbone_bd_ram_mem2_reg[78][18]/P0001 ,
		_w12874_,
		_w18299_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		\wishbone_bd_ram_mem2_reg[52][18]/P0001 ,
		_w13082_,
		_w18300_
	);
	LUT2 #(
		.INIT('h8)
	) name7789 (
		\wishbone_bd_ram_mem2_reg[192][18]/P0001 ,
		_w12938_,
		_w18301_
	);
	LUT2 #(
		.INIT('h8)
	) name7790 (
		\wishbone_bd_ram_mem2_reg[116][18]/P0001 ,
		_w12998_,
		_w18302_
	);
	LUT2 #(
		.INIT('h8)
	) name7791 (
		\wishbone_bd_ram_mem2_reg[36][18]/P0001 ,
		_w12800_,
		_w18303_
	);
	LUT2 #(
		.INIT('h8)
	) name7792 (
		\wishbone_bd_ram_mem2_reg[219][18]/P0001 ,
		_w12806_,
		_w18304_
	);
	LUT2 #(
		.INIT('h8)
	) name7793 (
		\wishbone_bd_ram_mem2_reg[235][18]/P0001 ,
		_w12696_,
		_w18305_
	);
	LUT2 #(
		.INIT('h8)
	) name7794 (
		\wishbone_bd_ram_mem2_reg[110][18]/P0001 ,
		_w13046_,
		_w18306_
	);
	LUT2 #(
		.INIT('h8)
	) name7795 (
		\wishbone_bd_ram_mem2_reg[27][18]/P0001 ,
		_w12880_,
		_w18307_
	);
	LUT2 #(
		.INIT('h8)
	) name7796 (
		\wishbone_bd_ram_mem2_reg[183][18]/P0001 ,
		_w12787_,
		_w18308_
	);
	LUT2 #(
		.INIT('h1)
	) name7797 (
		_w18053_,
		_w18054_,
		_w18309_
	);
	LUT2 #(
		.INIT('h1)
	) name7798 (
		_w18055_,
		_w18056_,
		_w18310_
	);
	LUT2 #(
		.INIT('h1)
	) name7799 (
		_w18057_,
		_w18058_,
		_w18311_
	);
	LUT2 #(
		.INIT('h1)
	) name7800 (
		_w18059_,
		_w18060_,
		_w18312_
	);
	LUT2 #(
		.INIT('h1)
	) name7801 (
		_w18061_,
		_w18062_,
		_w18313_
	);
	LUT2 #(
		.INIT('h1)
	) name7802 (
		_w18063_,
		_w18064_,
		_w18314_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w18065_,
		_w18066_,
		_w18315_
	);
	LUT2 #(
		.INIT('h1)
	) name7804 (
		_w18067_,
		_w18068_,
		_w18316_
	);
	LUT2 #(
		.INIT('h1)
	) name7805 (
		_w18069_,
		_w18070_,
		_w18317_
	);
	LUT2 #(
		.INIT('h1)
	) name7806 (
		_w18071_,
		_w18072_,
		_w18318_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w18073_,
		_w18074_,
		_w18319_
	);
	LUT2 #(
		.INIT('h1)
	) name7808 (
		_w18075_,
		_w18076_,
		_w18320_
	);
	LUT2 #(
		.INIT('h1)
	) name7809 (
		_w18077_,
		_w18078_,
		_w18321_
	);
	LUT2 #(
		.INIT('h1)
	) name7810 (
		_w18079_,
		_w18080_,
		_w18322_
	);
	LUT2 #(
		.INIT('h1)
	) name7811 (
		_w18081_,
		_w18082_,
		_w18323_
	);
	LUT2 #(
		.INIT('h1)
	) name7812 (
		_w18083_,
		_w18084_,
		_w18324_
	);
	LUT2 #(
		.INIT('h1)
	) name7813 (
		_w18085_,
		_w18086_,
		_w18325_
	);
	LUT2 #(
		.INIT('h1)
	) name7814 (
		_w18087_,
		_w18088_,
		_w18326_
	);
	LUT2 #(
		.INIT('h1)
	) name7815 (
		_w18089_,
		_w18090_,
		_w18327_
	);
	LUT2 #(
		.INIT('h1)
	) name7816 (
		_w18091_,
		_w18092_,
		_w18328_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w18093_,
		_w18094_,
		_w18329_
	);
	LUT2 #(
		.INIT('h1)
	) name7818 (
		_w18095_,
		_w18096_,
		_w18330_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		_w18097_,
		_w18098_,
		_w18331_
	);
	LUT2 #(
		.INIT('h1)
	) name7820 (
		_w18099_,
		_w18100_,
		_w18332_
	);
	LUT2 #(
		.INIT('h1)
	) name7821 (
		_w18101_,
		_w18102_,
		_w18333_
	);
	LUT2 #(
		.INIT('h1)
	) name7822 (
		_w18103_,
		_w18104_,
		_w18334_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w18105_,
		_w18106_,
		_w18335_
	);
	LUT2 #(
		.INIT('h1)
	) name7824 (
		_w18107_,
		_w18108_,
		_w18336_
	);
	LUT2 #(
		.INIT('h1)
	) name7825 (
		_w18109_,
		_w18110_,
		_w18337_
	);
	LUT2 #(
		.INIT('h1)
	) name7826 (
		_w18111_,
		_w18112_,
		_w18338_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w18113_,
		_w18114_,
		_w18339_
	);
	LUT2 #(
		.INIT('h1)
	) name7828 (
		_w18115_,
		_w18116_,
		_w18340_
	);
	LUT2 #(
		.INIT('h1)
	) name7829 (
		_w18117_,
		_w18118_,
		_w18341_
	);
	LUT2 #(
		.INIT('h1)
	) name7830 (
		_w18119_,
		_w18120_,
		_w18342_
	);
	LUT2 #(
		.INIT('h1)
	) name7831 (
		_w18121_,
		_w18122_,
		_w18343_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		_w18123_,
		_w18124_,
		_w18344_
	);
	LUT2 #(
		.INIT('h1)
	) name7833 (
		_w18125_,
		_w18126_,
		_w18345_
	);
	LUT2 #(
		.INIT('h1)
	) name7834 (
		_w18127_,
		_w18128_,
		_w18346_
	);
	LUT2 #(
		.INIT('h1)
	) name7835 (
		_w18129_,
		_w18130_,
		_w18347_
	);
	LUT2 #(
		.INIT('h1)
	) name7836 (
		_w18131_,
		_w18132_,
		_w18348_
	);
	LUT2 #(
		.INIT('h1)
	) name7837 (
		_w18133_,
		_w18134_,
		_w18349_
	);
	LUT2 #(
		.INIT('h1)
	) name7838 (
		_w18135_,
		_w18136_,
		_w18350_
	);
	LUT2 #(
		.INIT('h1)
	) name7839 (
		_w18137_,
		_w18138_,
		_w18351_
	);
	LUT2 #(
		.INIT('h1)
	) name7840 (
		_w18139_,
		_w18140_,
		_w18352_
	);
	LUT2 #(
		.INIT('h1)
	) name7841 (
		_w18141_,
		_w18142_,
		_w18353_
	);
	LUT2 #(
		.INIT('h1)
	) name7842 (
		_w18143_,
		_w18144_,
		_w18354_
	);
	LUT2 #(
		.INIT('h1)
	) name7843 (
		_w18145_,
		_w18146_,
		_w18355_
	);
	LUT2 #(
		.INIT('h1)
	) name7844 (
		_w18147_,
		_w18148_,
		_w18356_
	);
	LUT2 #(
		.INIT('h1)
	) name7845 (
		_w18149_,
		_w18150_,
		_w18357_
	);
	LUT2 #(
		.INIT('h1)
	) name7846 (
		_w18151_,
		_w18152_,
		_w18358_
	);
	LUT2 #(
		.INIT('h1)
	) name7847 (
		_w18153_,
		_w18154_,
		_w18359_
	);
	LUT2 #(
		.INIT('h1)
	) name7848 (
		_w18155_,
		_w18156_,
		_w18360_
	);
	LUT2 #(
		.INIT('h1)
	) name7849 (
		_w18157_,
		_w18158_,
		_w18361_
	);
	LUT2 #(
		.INIT('h1)
	) name7850 (
		_w18159_,
		_w18160_,
		_w18362_
	);
	LUT2 #(
		.INIT('h1)
	) name7851 (
		_w18161_,
		_w18162_,
		_w18363_
	);
	LUT2 #(
		.INIT('h1)
	) name7852 (
		_w18163_,
		_w18164_,
		_w18364_
	);
	LUT2 #(
		.INIT('h1)
	) name7853 (
		_w18165_,
		_w18166_,
		_w18365_
	);
	LUT2 #(
		.INIT('h1)
	) name7854 (
		_w18167_,
		_w18168_,
		_w18366_
	);
	LUT2 #(
		.INIT('h1)
	) name7855 (
		_w18169_,
		_w18170_,
		_w18367_
	);
	LUT2 #(
		.INIT('h1)
	) name7856 (
		_w18171_,
		_w18172_,
		_w18368_
	);
	LUT2 #(
		.INIT('h1)
	) name7857 (
		_w18173_,
		_w18174_,
		_w18369_
	);
	LUT2 #(
		.INIT('h1)
	) name7858 (
		_w18175_,
		_w18176_,
		_w18370_
	);
	LUT2 #(
		.INIT('h1)
	) name7859 (
		_w18177_,
		_w18178_,
		_w18371_
	);
	LUT2 #(
		.INIT('h1)
	) name7860 (
		_w18179_,
		_w18180_,
		_w18372_
	);
	LUT2 #(
		.INIT('h1)
	) name7861 (
		_w18181_,
		_w18182_,
		_w18373_
	);
	LUT2 #(
		.INIT('h1)
	) name7862 (
		_w18183_,
		_w18184_,
		_w18374_
	);
	LUT2 #(
		.INIT('h1)
	) name7863 (
		_w18185_,
		_w18186_,
		_w18375_
	);
	LUT2 #(
		.INIT('h1)
	) name7864 (
		_w18187_,
		_w18188_,
		_w18376_
	);
	LUT2 #(
		.INIT('h1)
	) name7865 (
		_w18189_,
		_w18190_,
		_w18377_
	);
	LUT2 #(
		.INIT('h1)
	) name7866 (
		_w18191_,
		_w18192_,
		_w18378_
	);
	LUT2 #(
		.INIT('h1)
	) name7867 (
		_w18193_,
		_w18194_,
		_w18379_
	);
	LUT2 #(
		.INIT('h1)
	) name7868 (
		_w18195_,
		_w18196_,
		_w18380_
	);
	LUT2 #(
		.INIT('h1)
	) name7869 (
		_w18197_,
		_w18198_,
		_w18381_
	);
	LUT2 #(
		.INIT('h1)
	) name7870 (
		_w18199_,
		_w18200_,
		_w18382_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w18201_,
		_w18202_,
		_w18383_
	);
	LUT2 #(
		.INIT('h1)
	) name7872 (
		_w18203_,
		_w18204_,
		_w18384_
	);
	LUT2 #(
		.INIT('h1)
	) name7873 (
		_w18205_,
		_w18206_,
		_w18385_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		_w18207_,
		_w18208_,
		_w18386_
	);
	LUT2 #(
		.INIT('h1)
	) name7875 (
		_w18209_,
		_w18210_,
		_w18387_
	);
	LUT2 #(
		.INIT('h1)
	) name7876 (
		_w18211_,
		_w18212_,
		_w18388_
	);
	LUT2 #(
		.INIT('h1)
	) name7877 (
		_w18213_,
		_w18214_,
		_w18389_
	);
	LUT2 #(
		.INIT('h1)
	) name7878 (
		_w18215_,
		_w18216_,
		_w18390_
	);
	LUT2 #(
		.INIT('h1)
	) name7879 (
		_w18217_,
		_w18218_,
		_w18391_
	);
	LUT2 #(
		.INIT('h1)
	) name7880 (
		_w18219_,
		_w18220_,
		_w18392_
	);
	LUT2 #(
		.INIT('h1)
	) name7881 (
		_w18221_,
		_w18222_,
		_w18393_
	);
	LUT2 #(
		.INIT('h1)
	) name7882 (
		_w18223_,
		_w18224_,
		_w18394_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		_w18225_,
		_w18226_,
		_w18395_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w18227_,
		_w18228_,
		_w18396_
	);
	LUT2 #(
		.INIT('h1)
	) name7885 (
		_w18229_,
		_w18230_,
		_w18397_
	);
	LUT2 #(
		.INIT('h1)
	) name7886 (
		_w18231_,
		_w18232_,
		_w18398_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w18233_,
		_w18234_,
		_w18399_
	);
	LUT2 #(
		.INIT('h1)
	) name7888 (
		_w18235_,
		_w18236_,
		_w18400_
	);
	LUT2 #(
		.INIT('h1)
	) name7889 (
		_w18237_,
		_w18238_,
		_w18401_
	);
	LUT2 #(
		.INIT('h1)
	) name7890 (
		_w18239_,
		_w18240_,
		_w18402_
	);
	LUT2 #(
		.INIT('h1)
	) name7891 (
		_w18241_,
		_w18242_,
		_w18403_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		_w18243_,
		_w18244_,
		_w18404_
	);
	LUT2 #(
		.INIT('h1)
	) name7893 (
		_w18245_,
		_w18246_,
		_w18405_
	);
	LUT2 #(
		.INIT('h1)
	) name7894 (
		_w18247_,
		_w18248_,
		_w18406_
	);
	LUT2 #(
		.INIT('h1)
	) name7895 (
		_w18249_,
		_w18250_,
		_w18407_
	);
	LUT2 #(
		.INIT('h1)
	) name7896 (
		_w18251_,
		_w18252_,
		_w18408_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		_w18253_,
		_w18254_,
		_w18409_
	);
	LUT2 #(
		.INIT('h1)
	) name7898 (
		_w18255_,
		_w18256_,
		_w18410_
	);
	LUT2 #(
		.INIT('h1)
	) name7899 (
		_w18257_,
		_w18258_,
		_w18411_
	);
	LUT2 #(
		.INIT('h1)
	) name7900 (
		_w18259_,
		_w18260_,
		_w18412_
	);
	LUT2 #(
		.INIT('h1)
	) name7901 (
		_w18261_,
		_w18262_,
		_w18413_
	);
	LUT2 #(
		.INIT('h1)
	) name7902 (
		_w18263_,
		_w18264_,
		_w18414_
	);
	LUT2 #(
		.INIT('h1)
	) name7903 (
		_w18265_,
		_w18266_,
		_w18415_
	);
	LUT2 #(
		.INIT('h1)
	) name7904 (
		_w18267_,
		_w18268_,
		_w18416_
	);
	LUT2 #(
		.INIT('h1)
	) name7905 (
		_w18269_,
		_w18270_,
		_w18417_
	);
	LUT2 #(
		.INIT('h1)
	) name7906 (
		_w18271_,
		_w18272_,
		_w18418_
	);
	LUT2 #(
		.INIT('h1)
	) name7907 (
		_w18273_,
		_w18274_,
		_w18419_
	);
	LUT2 #(
		.INIT('h1)
	) name7908 (
		_w18275_,
		_w18276_,
		_w18420_
	);
	LUT2 #(
		.INIT('h1)
	) name7909 (
		_w18277_,
		_w18278_,
		_w18421_
	);
	LUT2 #(
		.INIT('h1)
	) name7910 (
		_w18279_,
		_w18280_,
		_w18422_
	);
	LUT2 #(
		.INIT('h1)
	) name7911 (
		_w18281_,
		_w18282_,
		_w18423_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w18283_,
		_w18284_,
		_w18424_
	);
	LUT2 #(
		.INIT('h1)
	) name7913 (
		_w18285_,
		_w18286_,
		_w18425_
	);
	LUT2 #(
		.INIT('h1)
	) name7914 (
		_w18287_,
		_w18288_,
		_w18426_
	);
	LUT2 #(
		.INIT('h1)
	) name7915 (
		_w18289_,
		_w18290_,
		_w18427_
	);
	LUT2 #(
		.INIT('h1)
	) name7916 (
		_w18291_,
		_w18292_,
		_w18428_
	);
	LUT2 #(
		.INIT('h1)
	) name7917 (
		_w18293_,
		_w18294_,
		_w18429_
	);
	LUT2 #(
		.INIT('h1)
	) name7918 (
		_w18295_,
		_w18296_,
		_w18430_
	);
	LUT2 #(
		.INIT('h1)
	) name7919 (
		_w18297_,
		_w18298_,
		_w18431_
	);
	LUT2 #(
		.INIT('h1)
	) name7920 (
		_w18299_,
		_w18300_,
		_w18432_
	);
	LUT2 #(
		.INIT('h1)
	) name7921 (
		_w18301_,
		_w18302_,
		_w18433_
	);
	LUT2 #(
		.INIT('h1)
	) name7922 (
		_w18303_,
		_w18304_,
		_w18434_
	);
	LUT2 #(
		.INIT('h1)
	) name7923 (
		_w18305_,
		_w18306_,
		_w18435_
	);
	LUT2 #(
		.INIT('h1)
	) name7924 (
		_w18307_,
		_w18308_,
		_w18436_
	);
	LUT2 #(
		.INIT('h8)
	) name7925 (
		_w18435_,
		_w18436_,
		_w18437_
	);
	LUT2 #(
		.INIT('h8)
	) name7926 (
		_w18433_,
		_w18434_,
		_w18438_
	);
	LUT2 #(
		.INIT('h8)
	) name7927 (
		_w18431_,
		_w18432_,
		_w18439_
	);
	LUT2 #(
		.INIT('h8)
	) name7928 (
		_w18429_,
		_w18430_,
		_w18440_
	);
	LUT2 #(
		.INIT('h8)
	) name7929 (
		_w18427_,
		_w18428_,
		_w18441_
	);
	LUT2 #(
		.INIT('h8)
	) name7930 (
		_w18425_,
		_w18426_,
		_w18442_
	);
	LUT2 #(
		.INIT('h8)
	) name7931 (
		_w18423_,
		_w18424_,
		_w18443_
	);
	LUT2 #(
		.INIT('h8)
	) name7932 (
		_w18421_,
		_w18422_,
		_w18444_
	);
	LUT2 #(
		.INIT('h8)
	) name7933 (
		_w18419_,
		_w18420_,
		_w18445_
	);
	LUT2 #(
		.INIT('h8)
	) name7934 (
		_w18417_,
		_w18418_,
		_w18446_
	);
	LUT2 #(
		.INIT('h8)
	) name7935 (
		_w18415_,
		_w18416_,
		_w18447_
	);
	LUT2 #(
		.INIT('h8)
	) name7936 (
		_w18413_,
		_w18414_,
		_w18448_
	);
	LUT2 #(
		.INIT('h8)
	) name7937 (
		_w18411_,
		_w18412_,
		_w18449_
	);
	LUT2 #(
		.INIT('h8)
	) name7938 (
		_w18409_,
		_w18410_,
		_w18450_
	);
	LUT2 #(
		.INIT('h8)
	) name7939 (
		_w18407_,
		_w18408_,
		_w18451_
	);
	LUT2 #(
		.INIT('h8)
	) name7940 (
		_w18405_,
		_w18406_,
		_w18452_
	);
	LUT2 #(
		.INIT('h8)
	) name7941 (
		_w18403_,
		_w18404_,
		_w18453_
	);
	LUT2 #(
		.INIT('h8)
	) name7942 (
		_w18401_,
		_w18402_,
		_w18454_
	);
	LUT2 #(
		.INIT('h8)
	) name7943 (
		_w18399_,
		_w18400_,
		_w18455_
	);
	LUT2 #(
		.INIT('h8)
	) name7944 (
		_w18397_,
		_w18398_,
		_w18456_
	);
	LUT2 #(
		.INIT('h8)
	) name7945 (
		_w18395_,
		_w18396_,
		_w18457_
	);
	LUT2 #(
		.INIT('h8)
	) name7946 (
		_w18393_,
		_w18394_,
		_w18458_
	);
	LUT2 #(
		.INIT('h8)
	) name7947 (
		_w18391_,
		_w18392_,
		_w18459_
	);
	LUT2 #(
		.INIT('h8)
	) name7948 (
		_w18389_,
		_w18390_,
		_w18460_
	);
	LUT2 #(
		.INIT('h8)
	) name7949 (
		_w18387_,
		_w18388_,
		_w18461_
	);
	LUT2 #(
		.INIT('h8)
	) name7950 (
		_w18385_,
		_w18386_,
		_w18462_
	);
	LUT2 #(
		.INIT('h8)
	) name7951 (
		_w18383_,
		_w18384_,
		_w18463_
	);
	LUT2 #(
		.INIT('h8)
	) name7952 (
		_w18381_,
		_w18382_,
		_w18464_
	);
	LUT2 #(
		.INIT('h8)
	) name7953 (
		_w18379_,
		_w18380_,
		_w18465_
	);
	LUT2 #(
		.INIT('h8)
	) name7954 (
		_w18377_,
		_w18378_,
		_w18466_
	);
	LUT2 #(
		.INIT('h8)
	) name7955 (
		_w18375_,
		_w18376_,
		_w18467_
	);
	LUT2 #(
		.INIT('h8)
	) name7956 (
		_w18373_,
		_w18374_,
		_w18468_
	);
	LUT2 #(
		.INIT('h8)
	) name7957 (
		_w18371_,
		_w18372_,
		_w18469_
	);
	LUT2 #(
		.INIT('h8)
	) name7958 (
		_w18369_,
		_w18370_,
		_w18470_
	);
	LUT2 #(
		.INIT('h8)
	) name7959 (
		_w18367_,
		_w18368_,
		_w18471_
	);
	LUT2 #(
		.INIT('h8)
	) name7960 (
		_w18365_,
		_w18366_,
		_w18472_
	);
	LUT2 #(
		.INIT('h8)
	) name7961 (
		_w18363_,
		_w18364_,
		_w18473_
	);
	LUT2 #(
		.INIT('h8)
	) name7962 (
		_w18361_,
		_w18362_,
		_w18474_
	);
	LUT2 #(
		.INIT('h8)
	) name7963 (
		_w18359_,
		_w18360_,
		_w18475_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		_w18357_,
		_w18358_,
		_w18476_
	);
	LUT2 #(
		.INIT('h8)
	) name7965 (
		_w18355_,
		_w18356_,
		_w18477_
	);
	LUT2 #(
		.INIT('h8)
	) name7966 (
		_w18353_,
		_w18354_,
		_w18478_
	);
	LUT2 #(
		.INIT('h8)
	) name7967 (
		_w18351_,
		_w18352_,
		_w18479_
	);
	LUT2 #(
		.INIT('h8)
	) name7968 (
		_w18349_,
		_w18350_,
		_w18480_
	);
	LUT2 #(
		.INIT('h8)
	) name7969 (
		_w18347_,
		_w18348_,
		_w18481_
	);
	LUT2 #(
		.INIT('h8)
	) name7970 (
		_w18345_,
		_w18346_,
		_w18482_
	);
	LUT2 #(
		.INIT('h8)
	) name7971 (
		_w18343_,
		_w18344_,
		_w18483_
	);
	LUT2 #(
		.INIT('h8)
	) name7972 (
		_w18341_,
		_w18342_,
		_w18484_
	);
	LUT2 #(
		.INIT('h8)
	) name7973 (
		_w18339_,
		_w18340_,
		_w18485_
	);
	LUT2 #(
		.INIT('h8)
	) name7974 (
		_w18337_,
		_w18338_,
		_w18486_
	);
	LUT2 #(
		.INIT('h8)
	) name7975 (
		_w18335_,
		_w18336_,
		_w18487_
	);
	LUT2 #(
		.INIT('h8)
	) name7976 (
		_w18333_,
		_w18334_,
		_w18488_
	);
	LUT2 #(
		.INIT('h8)
	) name7977 (
		_w18331_,
		_w18332_,
		_w18489_
	);
	LUT2 #(
		.INIT('h8)
	) name7978 (
		_w18329_,
		_w18330_,
		_w18490_
	);
	LUT2 #(
		.INIT('h8)
	) name7979 (
		_w18327_,
		_w18328_,
		_w18491_
	);
	LUT2 #(
		.INIT('h8)
	) name7980 (
		_w18325_,
		_w18326_,
		_w18492_
	);
	LUT2 #(
		.INIT('h8)
	) name7981 (
		_w18323_,
		_w18324_,
		_w18493_
	);
	LUT2 #(
		.INIT('h8)
	) name7982 (
		_w18321_,
		_w18322_,
		_w18494_
	);
	LUT2 #(
		.INIT('h8)
	) name7983 (
		_w18319_,
		_w18320_,
		_w18495_
	);
	LUT2 #(
		.INIT('h8)
	) name7984 (
		_w18317_,
		_w18318_,
		_w18496_
	);
	LUT2 #(
		.INIT('h8)
	) name7985 (
		_w18315_,
		_w18316_,
		_w18497_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		_w18313_,
		_w18314_,
		_w18498_
	);
	LUT2 #(
		.INIT('h8)
	) name7987 (
		_w18311_,
		_w18312_,
		_w18499_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		_w18309_,
		_w18310_,
		_w18500_
	);
	LUT2 #(
		.INIT('h8)
	) name7989 (
		_w18499_,
		_w18500_,
		_w18501_
	);
	LUT2 #(
		.INIT('h8)
	) name7990 (
		_w18497_,
		_w18498_,
		_w18502_
	);
	LUT2 #(
		.INIT('h8)
	) name7991 (
		_w18495_,
		_w18496_,
		_w18503_
	);
	LUT2 #(
		.INIT('h8)
	) name7992 (
		_w18493_,
		_w18494_,
		_w18504_
	);
	LUT2 #(
		.INIT('h8)
	) name7993 (
		_w18491_,
		_w18492_,
		_w18505_
	);
	LUT2 #(
		.INIT('h8)
	) name7994 (
		_w18489_,
		_w18490_,
		_w18506_
	);
	LUT2 #(
		.INIT('h8)
	) name7995 (
		_w18487_,
		_w18488_,
		_w18507_
	);
	LUT2 #(
		.INIT('h8)
	) name7996 (
		_w18485_,
		_w18486_,
		_w18508_
	);
	LUT2 #(
		.INIT('h8)
	) name7997 (
		_w18483_,
		_w18484_,
		_w18509_
	);
	LUT2 #(
		.INIT('h8)
	) name7998 (
		_w18481_,
		_w18482_,
		_w18510_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		_w18479_,
		_w18480_,
		_w18511_
	);
	LUT2 #(
		.INIT('h8)
	) name8000 (
		_w18477_,
		_w18478_,
		_w18512_
	);
	LUT2 #(
		.INIT('h8)
	) name8001 (
		_w18475_,
		_w18476_,
		_w18513_
	);
	LUT2 #(
		.INIT('h8)
	) name8002 (
		_w18473_,
		_w18474_,
		_w18514_
	);
	LUT2 #(
		.INIT('h8)
	) name8003 (
		_w18471_,
		_w18472_,
		_w18515_
	);
	LUT2 #(
		.INIT('h8)
	) name8004 (
		_w18469_,
		_w18470_,
		_w18516_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		_w18467_,
		_w18468_,
		_w18517_
	);
	LUT2 #(
		.INIT('h8)
	) name8006 (
		_w18465_,
		_w18466_,
		_w18518_
	);
	LUT2 #(
		.INIT('h8)
	) name8007 (
		_w18463_,
		_w18464_,
		_w18519_
	);
	LUT2 #(
		.INIT('h8)
	) name8008 (
		_w18461_,
		_w18462_,
		_w18520_
	);
	LUT2 #(
		.INIT('h8)
	) name8009 (
		_w18459_,
		_w18460_,
		_w18521_
	);
	LUT2 #(
		.INIT('h8)
	) name8010 (
		_w18457_,
		_w18458_,
		_w18522_
	);
	LUT2 #(
		.INIT('h8)
	) name8011 (
		_w18455_,
		_w18456_,
		_w18523_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		_w18453_,
		_w18454_,
		_w18524_
	);
	LUT2 #(
		.INIT('h8)
	) name8013 (
		_w18451_,
		_w18452_,
		_w18525_
	);
	LUT2 #(
		.INIT('h8)
	) name8014 (
		_w18449_,
		_w18450_,
		_w18526_
	);
	LUT2 #(
		.INIT('h8)
	) name8015 (
		_w18447_,
		_w18448_,
		_w18527_
	);
	LUT2 #(
		.INIT('h8)
	) name8016 (
		_w18445_,
		_w18446_,
		_w18528_
	);
	LUT2 #(
		.INIT('h8)
	) name8017 (
		_w18443_,
		_w18444_,
		_w18529_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		_w18441_,
		_w18442_,
		_w18530_
	);
	LUT2 #(
		.INIT('h8)
	) name8019 (
		_w18439_,
		_w18440_,
		_w18531_
	);
	LUT2 #(
		.INIT('h8)
	) name8020 (
		_w18437_,
		_w18438_,
		_w18532_
	);
	LUT2 #(
		.INIT('h8)
	) name8021 (
		_w18531_,
		_w18532_,
		_w18533_
	);
	LUT2 #(
		.INIT('h8)
	) name8022 (
		_w18529_,
		_w18530_,
		_w18534_
	);
	LUT2 #(
		.INIT('h8)
	) name8023 (
		_w18527_,
		_w18528_,
		_w18535_
	);
	LUT2 #(
		.INIT('h8)
	) name8024 (
		_w18525_,
		_w18526_,
		_w18536_
	);
	LUT2 #(
		.INIT('h8)
	) name8025 (
		_w18523_,
		_w18524_,
		_w18537_
	);
	LUT2 #(
		.INIT('h8)
	) name8026 (
		_w18521_,
		_w18522_,
		_w18538_
	);
	LUT2 #(
		.INIT('h8)
	) name8027 (
		_w18519_,
		_w18520_,
		_w18539_
	);
	LUT2 #(
		.INIT('h8)
	) name8028 (
		_w18517_,
		_w18518_,
		_w18540_
	);
	LUT2 #(
		.INIT('h8)
	) name8029 (
		_w18515_,
		_w18516_,
		_w18541_
	);
	LUT2 #(
		.INIT('h8)
	) name8030 (
		_w18513_,
		_w18514_,
		_w18542_
	);
	LUT2 #(
		.INIT('h8)
	) name8031 (
		_w18511_,
		_w18512_,
		_w18543_
	);
	LUT2 #(
		.INIT('h8)
	) name8032 (
		_w18509_,
		_w18510_,
		_w18544_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		_w18507_,
		_w18508_,
		_w18545_
	);
	LUT2 #(
		.INIT('h8)
	) name8034 (
		_w18505_,
		_w18506_,
		_w18546_
	);
	LUT2 #(
		.INIT('h8)
	) name8035 (
		_w18503_,
		_w18504_,
		_w18547_
	);
	LUT2 #(
		.INIT('h8)
	) name8036 (
		_w18501_,
		_w18502_,
		_w18548_
	);
	LUT2 #(
		.INIT('h8)
	) name8037 (
		_w18547_,
		_w18548_,
		_w18549_
	);
	LUT2 #(
		.INIT('h8)
	) name8038 (
		_w18545_,
		_w18546_,
		_w18550_
	);
	LUT2 #(
		.INIT('h8)
	) name8039 (
		_w18543_,
		_w18544_,
		_w18551_
	);
	LUT2 #(
		.INIT('h8)
	) name8040 (
		_w18541_,
		_w18542_,
		_w18552_
	);
	LUT2 #(
		.INIT('h8)
	) name8041 (
		_w18539_,
		_w18540_,
		_w18553_
	);
	LUT2 #(
		.INIT('h8)
	) name8042 (
		_w18537_,
		_w18538_,
		_w18554_
	);
	LUT2 #(
		.INIT('h8)
	) name8043 (
		_w18535_,
		_w18536_,
		_w18555_
	);
	LUT2 #(
		.INIT('h8)
	) name8044 (
		_w18533_,
		_w18534_,
		_w18556_
	);
	LUT2 #(
		.INIT('h8)
	) name8045 (
		_w18555_,
		_w18556_,
		_w18557_
	);
	LUT2 #(
		.INIT('h8)
	) name8046 (
		_w18553_,
		_w18554_,
		_w18558_
	);
	LUT2 #(
		.INIT('h8)
	) name8047 (
		_w18551_,
		_w18552_,
		_w18559_
	);
	LUT2 #(
		.INIT('h8)
	) name8048 (
		_w18549_,
		_w18550_,
		_w18560_
	);
	LUT2 #(
		.INIT('h8)
	) name8049 (
		_w18559_,
		_w18560_,
		_w18561_
	);
	LUT2 #(
		.INIT('h8)
	) name8050 (
		_w18557_,
		_w18558_,
		_w18562_
	);
	LUT2 #(
		.INIT('h8)
	) name8051 (
		_w18561_,
		_w18562_,
		_w18563_
	);
	LUT2 #(
		.INIT('h1)
	) name8052 (
		wb_rst_i_pad,
		_w18563_,
		_w18564_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		_w12656_,
		_w18564_,
		_w18565_
	);
	LUT2 #(
		.INIT('h1)
	) name8054 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w17289_,
		_w18566_
	);
	LUT2 #(
		.INIT('h8)
	) name8055 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w17289_,
		_w18567_
	);
	LUT2 #(
		.INIT('h8)
	) name8056 (
		_w12657_,
		_w13499_,
		_w18568_
	);
	LUT2 #(
		.INIT('h1)
	) name8057 (
		_w12656_,
		_w18568_,
		_w18569_
	);
	LUT2 #(
		.INIT('h1)
	) name8058 (
		_w18566_,
		_w18567_,
		_w18570_
	);
	LUT2 #(
		.INIT('h8)
	) name8059 (
		_w18569_,
		_w18570_,
		_w18571_
	);
	LUT2 #(
		.INIT('h1)
	) name8060 (
		_w18565_,
		_w18571_,
		_w18572_
	);
	LUT2 #(
		.INIT('h2)
	) name8061 (
		_w10580_,
		_w11743_,
		_w18573_
	);
	LUT2 #(
		.INIT('h1)
	) name8062 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w18574_
	);
	LUT2 #(
		.INIT('h1)
	) name8063 (
		_w13485_,
		_w18574_,
		_w18575_
	);
	LUT2 #(
		.INIT('h8)
	) name8064 (
		_w13501_,
		_w18575_,
		_w18576_
	);
	LUT2 #(
		.INIT('h8)
	) name8065 (
		\wishbone_bd_ram_mem2_reg[24][16]/P0001 ,
		_w13084_,
		_w18577_
	);
	LUT2 #(
		.INIT('h8)
	) name8066 (
		\wishbone_bd_ram_mem2_reg[108][16]/P0001 ,
		_w13156_,
		_w18578_
	);
	LUT2 #(
		.INIT('h8)
	) name8067 (
		\wishbone_bd_ram_mem2_reg[77][16]/P0001 ,
		_w12982_,
		_w18579_
	);
	LUT2 #(
		.INIT('h8)
	) name8068 (
		\wishbone_bd_ram_mem2_reg[147][16]/P0001 ,
		_w13146_,
		_w18580_
	);
	LUT2 #(
		.INIT('h8)
	) name8069 (
		\wishbone_bd_ram_mem2_reg[126][16]/P0001 ,
		_w13218_,
		_w18581_
	);
	LUT2 #(
		.INIT('h8)
	) name8070 (
		\wishbone_bd_ram_mem2_reg[235][16]/P0001 ,
		_w12696_,
		_w18582_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		\wishbone_bd_ram_mem2_reg[32][16]/P0001 ,
		_w13120_,
		_w18583_
	);
	LUT2 #(
		.INIT('h8)
	) name8072 (
		\wishbone_bd_ram_mem2_reg[185][16]/P0001 ,
		_w12940_,
		_w18584_
	);
	LUT2 #(
		.INIT('h8)
	) name8073 (
		\wishbone_bd_ram_mem2_reg[148][16]/P0001 ,
		_w13000_,
		_w18585_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		\wishbone_bd_ram_mem2_reg[117][16]/P0001 ,
		_w12715_,
		_w18586_
	);
	LUT2 #(
		.INIT('h8)
	) name8075 (
		\wishbone_bd_ram_mem2_reg[59][16]/P0001 ,
		_w12780_,
		_w18587_
	);
	LUT2 #(
		.INIT('h8)
	) name8076 (
		\wishbone_bd_ram_mem2_reg[160][16]/P0001 ,
		_w12872_,
		_w18588_
	);
	LUT2 #(
		.INIT('h8)
	) name8077 (
		\wishbone_bd_ram_mem2_reg[219][16]/P0001 ,
		_w12806_,
		_w18589_
	);
	LUT2 #(
		.INIT('h8)
	) name8078 (
		\wishbone_bd_ram_mem2_reg[47][16]/P0001 ,
		_w12904_,
		_w18590_
	);
	LUT2 #(
		.INIT('h8)
	) name8079 (
		\wishbone_bd_ram_mem2_reg[30][16]/P0001 ,
		_w13104_,
		_w18591_
	);
	LUT2 #(
		.INIT('h8)
	) name8080 (
		\wishbone_bd_ram_mem2_reg[7][16]/P0001 ,
		_w12728_,
		_w18592_
	);
	LUT2 #(
		.INIT('h8)
	) name8081 (
		\wishbone_bd_ram_mem2_reg[74][16]/P0001 ,
		_w12812_,
		_w18593_
	);
	LUT2 #(
		.INIT('h8)
	) name8082 (
		\wishbone_bd_ram_mem2_reg[116][16]/P0001 ,
		_w12998_,
		_w18594_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		\wishbone_bd_ram_mem2_reg[101][16]/P0001 ,
		_w13192_,
		_w18595_
	);
	LUT2 #(
		.INIT('h8)
	) name8084 (
		\wishbone_bd_ram_mem2_reg[58][16]/P0001 ,
		_w13070_,
		_w18596_
	);
	LUT2 #(
		.INIT('h8)
	) name8085 (
		\wishbone_bd_ram_mem2_reg[182][16]/P0001 ,
		_w12820_,
		_w18597_
	);
	LUT2 #(
		.INIT('h8)
	) name8086 (
		\wishbone_bd_ram_mem2_reg[42][16]/P0001 ,
		_w12842_,
		_w18598_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		\wishbone_bd_ram_mem2_reg[23][16]/P0001 ,
		_w13008_,
		_w18599_
	);
	LUT2 #(
		.INIT('h8)
	) name8088 (
		\wishbone_bd_ram_mem2_reg[213][16]/P0001 ,
		_w13002_,
		_w18600_
	);
	LUT2 #(
		.INIT('h8)
	) name8089 (
		\wishbone_bd_ram_mem2_reg[218][16]/P0001 ,
		_w13206_,
		_w18601_
	);
	LUT2 #(
		.INIT('h8)
	) name8090 (
		\wishbone_bd_ram_mem2_reg[10][16]/P0001 ,
		_w13172_,
		_w18602_
	);
	LUT2 #(
		.INIT('h8)
	) name8091 (
		\wishbone_bd_ram_mem2_reg[75][16]/P0001 ,
		_w12826_,
		_w18603_
	);
	LUT2 #(
		.INIT('h8)
	) name8092 (
		\wishbone_bd_ram_mem2_reg[184][16]/P0001 ,
		_w13062_,
		_w18604_
	);
	LUT2 #(
		.INIT('h8)
	) name8093 (
		\wishbone_bd_ram_mem2_reg[196][16]/P0001 ,
		_w13090_,
		_w18605_
	);
	LUT2 #(
		.INIT('h8)
	) name8094 (
		\wishbone_bd_ram_mem2_reg[1][16]/P0001 ,
		_w13014_,
		_w18606_
	);
	LUT2 #(
		.INIT('h8)
	) name8095 (
		\wishbone_bd_ram_mem2_reg[17][16]/P0001 ,
		_w12848_,
		_w18607_
	);
	LUT2 #(
		.INIT('h8)
	) name8096 (
		\wishbone_bd_ram_mem2_reg[2][16]/P0001 ,
		_w13088_,
		_w18608_
	);
	LUT2 #(
		.INIT('h8)
	) name8097 (
		\wishbone_bd_ram_mem2_reg[191][16]/P0001 ,
		_w13034_,
		_w18609_
	);
	LUT2 #(
		.INIT('h8)
	) name8098 (
		\wishbone_bd_ram_mem2_reg[80][16]/P0001 ,
		_w12689_,
		_w18610_
	);
	LUT2 #(
		.INIT('h8)
	) name8099 (
		\wishbone_bd_ram_mem2_reg[214][16]/P0001 ,
		_w12984_,
		_w18611_
	);
	LUT2 #(
		.INIT('h8)
	) name8100 (
		\wishbone_bd_ram_mem2_reg[194][16]/P0001 ,
		_w12772_,
		_w18612_
	);
	LUT2 #(
		.INIT('h8)
	) name8101 (
		\wishbone_bd_ram_mem2_reg[62][16]/P0001 ,
		_w12673_,
		_w18613_
	);
	LUT2 #(
		.INIT('h8)
	) name8102 (
		\wishbone_bd_ram_mem2_reg[21][16]/P0001 ,
		_w12906_,
		_w18614_
	);
	LUT2 #(
		.INIT('h8)
	) name8103 (
		\wishbone_bd_ram_mem2_reg[67][16]/P0001 ,
		_w13134_,
		_w18615_
	);
	LUT2 #(
		.INIT('h8)
	) name8104 (
		\wishbone_bd_ram_mem2_reg[159][16]/P0001 ,
		_w12774_,
		_w18616_
	);
	LUT2 #(
		.INIT('h8)
	) name8105 (
		\wishbone_bd_ram_mem2_reg[231][16]/P0001 ,
		_w12856_,
		_w18617_
	);
	LUT2 #(
		.INIT('h8)
	) name8106 (
		\wishbone_bd_ram_mem2_reg[183][16]/P0001 ,
		_w12787_,
		_w18618_
	);
	LUT2 #(
		.INIT('h8)
	) name8107 (
		\wishbone_bd_ram_mem2_reg[112][16]/P0001 ,
		_w12733_,
		_w18619_
	);
	LUT2 #(
		.INIT('h8)
	) name8108 (
		\wishbone_bd_ram_mem2_reg[88][16]/P0001 ,
		_w12860_,
		_w18620_
	);
	LUT2 #(
		.INIT('h8)
	) name8109 (
		\wishbone_bd_ram_mem2_reg[246][16]/P0001 ,
		_w13076_,
		_w18621_
	);
	LUT2 #(
		.INIT('h8)
	) name8110 (
		\wishbone_bd_ram_mem2_reg[151][16]/P0001 ,
		_w13142_,
		_w18622_
	);
	LUT2 #(
		.INIT('h8)
	) name8111 (
		\wishbone_bd_ram_mem2_reg[172][16]/P0001 ,
		_w12944_,
		_w18623_
	);
	LUT2 #(
		.INIT('h8)
	) name8112 (
		\wishbone_bd_ram_mem2_reg[86][16]/P0001 ,
		_w12735_,
		_w18624_
	);
	LUT2 #(
		.INIT('h8)
	) name8113 (
		\wishbone_bd_ram_mem2_reg[134][16]/P0001 ,
		_w12763_,
		_w18625_
	);
	LUT2 #(
		.INIT('h8)
	) name8114 (
		\wishbone_bd_ram_mem2_reg[234][16]/P0001 ,
		_w13214_,
		_w18626_
	);
	LUT2 #(
		.INIT('h8)
	) name8115 (
		\wishbone_bd_ram_mem2_reg[203][16]/P0001 ,
		_w13158_,
		_w18627_
	);
	LUT2 #(
		.INIT('h8)
	) name8116 (
		\wishbone_bd_ram_mem2_reg[49][16]/P0001 ,
		_w12994_,
		_w18628_
	);
	LUT2 #(
		.INIT('h8)
	) name8117 (
		\wishbone_bd_ram_mem2_reg[124][16]/P0001 ,
		_w13058_,
		_w18629_
	);
	LUT2 #(
		.INIT('h8)
	) name8118 (
		\wishbone_bd_ram_mem2_reg[57][16]/P0001 ,
		_w13116_,
		_w18630_
	);
	LUT2 #(
		.INIT('h8)
	) name8119 (
		\wishbone_bd_ram_mem2_reg[45][16]/P0001 ,
		_w12908_,
		_w18631_
	);
	LUT2 #(
		.INIT('h8)
	) name8120 (
		\wishbone_bd_ram_mem2_reg[190][16]/P0001 ,
		_w12858_,
		_w18632_
	);
	LUT2 #(
		.INIT('h8)
	) name8121 (
		\wishbone_bd_ram_mem2_reg[200][16]/P0001 ,
		_w12988_,
		_w18633_
	);
	LUT2 #(
		.INIT('h8)
	) name8122 (
		\wishbone_bd_ram_mem2_reg[44][16]/P0001 ,
		_w12896_,
		_w18634_
	);
	LUT2 #(
		.INIT('h8)
	) name8123 (
		\wishbone_bd_ram_mem2_reg[96][16]/P0001 ,
		_w12912_,
		_w18635_
	);
	LUT2 #(
		.INIT('h8)
	) name8124 (
		\wishbone_bd_ram_mem2_reg[38][16]/P0001 ,
		_w13182_,
		_w18636_
	);
	LUT2 #(
		.INIT('h8)
	) name8125 (
		\wishbone_bd_ram_mem2_reg[36][16]/P0001 ,
		_w12800_,
		_w18637_
	);
	LUT2 #(
		.INIT('h8)
	) name8126 (
		\wishbone_bd_ram_mem2_reg[150][16]/P0001 ,
		_w13136_,
		_w18638_
	);
	LUT2 #(
		.INIT('h8)
	) name8127 (
		\wishbone_bd_ram_mem2_reg[115][16]/P0001 ,
		_w13112_,
		_w18639_
	);
	LUT2 #(
		.INIT('h8)
	) name8128 (
		\wishbone_bd_ram_mem2_reg[163][16]/P0001 ,
		_w12882_,
		_w18640_
	);
	LUT2 #(
		.INIT('h8)
	) name8129 (
		\wishbone_bd_ram_mem2_reg[221][16]/P0001 ,
		_w12802_,
		_w18641_
	);
	LUT2 #(
		.INIT('h8)
	) name8130 (
		\wishbone_bd_ram_mem2_reg[0][16]/P0001 ,
		_w12717_,
		_w18642_
	);
	LUT2 #(
		.INIT('h8)
	) name8131 (
		\wishbone_bd_ram_mem2_reg[8][16]/P0001 ,
		_w12920_,
		_w18643_
	);
	LUT2 #(
		.INIT('h8)
	) name8132 (
		\wishbone_bd_ram_mem2_reg[100][16]/P0001 ,
		_w12960_,
		_w18644_
	);
	LUT2 #(
		.INIT('h8)
	) name8133 (
		\wishbone_bd_ram_mem2_reg[204][16]/P0001 ,
		_w13162_,
		_w18645_
	);
	LUT2 #(
		.INIT('h8)
	) name8134 (
		\wishbone_bd_ram_mem2_reg[120][16]/P0001 ,
		_w12707_,
		_w18646_
	);
	LUT2 #(
		.INIT('h8)
	) name8135 (
		\wishbone_bd_ram_mem2_reg[79][16]/P0001 ,
		_w13212_,
		_w18647_
	);
	LUT2 #(
		.INIT('h8)
	) name8136 (
		\wishbone_bd_ram_mem2_reg[6][16]/P0001 ,
		_w12968_,
		_w18648_
	);
	LUT2 #(
		.INIT('h8)
	) name8137 (
		\wishbone_bd_ram_mem2_reg[122][16]/P0001 ,
		_w13130_,
		_w18649_
	);
	LUT2 #(
		.INIT('h8)
	) name8138 (
		\wishbone_bd_ram_mem2_reg[33][16]/P0001 ,
		_w12980_,
		_w18650_
	);
	LUT2 #(
		.INIT('h8)
	) name8139 (
		\wishbone_bd_ram_mem2_reg[91][16]/P0001 ,
		_w13074_,
		_w18651_
	);
	LUT2 #(
		.INIT('h8)
	) name8140 (
		\wishbone_bd_ram_mem2_reg[161][16]/P0001 ,
		_w12754_,
		_w18652_
	);
	LUT2 #(
		.INIT('h8)
	) name8141 (
		\wishbone_bd_ram_mem2_reg[164][16]/P0001 ,
		_w12876_,
		_w18653_
	);
	LUT2 #(
		.INIT('h8)
	) name8142 (
		\wishbone_bd_ram_mem2_reg[188][16]/P0001 ,
		_w12948_,
		_w18654_
	);
	LUT2 #(
		.INIT('h8)
	) name8143 (
		\wishbone_bd_ram_mem2_reg[241][16]/P0001 ,
		_w13006_,
		_w18655_
	);
	LUT2 #(
		.INIT('h8)
	) name8144 (
		\wishbone_bd_ram_mem2_reg[197][16]/P0001 ,
		_w12834_,
		_w18656_
	);
	LUT2 #(
		.INIT('h8)
	) name8145 (
		\wishbone_bd_ram_mem2_reg[220][16]/P0001 ,
		_w13066_,
		_w18657_
	);
	LUT2 #(
		.INIT('h8)
	) name8146 (
		\wishbone_bd_ram_mem2_reg[118][16]/P0001 ,
		_w12830_,
		_w18658_
	);
	LUT2 #(
		.INIT('h8)
	) name8147 (
		\wishbone_bd_ram_mem2_reg[138][16]/P0001 ,
		_w12958_,
		_w18659_
	);
	LUT2 #(
		.INIT('h8)
	) name8148 (
		\wishbone_bd_ram_mem2_reg[127][16]/P0001 ,
		_w13164_,
		_w18660_
	);
	LUT2 #(
		.INIT('h8)
	) name8149 (
		\wishbone_bd_ram_mem2_reg[128][16]/P0001 ,
		_w12793_,
		_w18661_
	);
	LUT2 #(
		.INIT('h8)
	) name8150 (
		\wishbone_bd_ram_mem2_reg[55][16]/P0001 ,
		_w12785_,
		_w18662_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		\wishbone_bd_ram_mem2_reg[34][16]/P0001 ,
		_w12930_,
		_w18663_
	);
	LUT2 #(
		.INIT('h8)
	) name8152 (
		\wishbone_bd_ram_mem2_reg[125][16]/P0001 ,
		_w12956_,
		_w18664_
	);
	LUT2 #(
		.INIT('h8)
	) name8153 (
		\wishbone_bd_ram_mem2_reg[137][16]/P0001 ,
		_w13168_,
		_w18665_
	);
	LUT2 #(
		.INIT('h8)
	) name8154 (
		\wishbone_bd_ram_mem2_reg[20][16]/P0001 ,
		_w13174_,
		_w18666_
	);
	LUT2 #(
		.INIT('h8)
	) name8155 (
		\wishbone_bd_ram_mem2_reg[31][16]/P0001 ,
		_w13198_,
		_w18667_
	);
	LUT2 #(
		.INIT('h8)
	) name8156 (
		\wishbone_bd_ram_mem2_reg[237][16]/P0001 ,
		_w12990_,
		_w18668_
	);
	LUT2 #(
		.INIT('h8)
	) name8157 (
		\wishbone_bd_ram_mem2_reg[103][16]/P0001 ,
		_w12846_,
		_w18669_
	);
	LUT2 #(
		.INIT('h8)
	) name8158 (
		\wishbone_bd_ram_mem2_reg[69][16]/P0001 ,
		_w12738_,
		_w18670_
	);
	LUT2 #(
		.INIT('h8)
	) name8159 (
		\wishbone_bd_ram_mem2_reg[254][16]/P0001 ,
		_w12892_,
		_w18671_
	);
	LUT2 #(
		.INIT('h8)
	) name8160 (
		\wishbone_bd_ram_mem2_reg[39][16]/P0001 ,
		_w13018_,
		_w18672_
	);
	LUT2 #(
		.INIT('h8)
	) name8161 (
		\wishbone_bd_ram_mem2_reg[202][16]/P0001 ,
		_w12870_,
		_w18673_
	);
	LUT2 #(
		.INIT('h8)
	) name8162 (
		\wishbone_bd_ram_mem2_reg[99][16]/P0001 ,
		_w13038_,
		_w18674_
	);
	LUT2 #(
		.INIT('h8)
	) name8163 (
		\wishbone_bd_ram_mem2_reg[13][16]/P0001 ,
		_w13178_,
		_w18675_
	);
	LUT2 #(
		.INIT('h8)
	) name8164 (
		\wishbone_bd_ram_mem2_reg[193][16]/P0001 ,
		_w13056_,
		_w18676_
	);
	LUT2 #(
		.INIT('h8)
	) name8165 (
		\wishbone_bd_ram_mem2_reg[121][16]/P0001 ,
		_w13078_,
		_w18677_
	);
	LUT2 #(
		.INIT('h8)
	) name8166 (
		\wishbone_bd_ram_mem2_reg[102][16]/P0001 ,
		_w12685_,
		_w18678_
	);
	LUT2 #(
		.INIT('h8)
	) name8167 (
		\wishbone_bd_ram_mem2_reg[93][16]/P0001 ,
		_w13016_,
		_w18679_
	);
	LUT2 #(
		.INIT('h8)
	) name8168 (
		\wishbone_bd_ram_mem2_reg[158][16]/P0001 ,
		_w12898_,
		_w18680_
	);
	LUT2 #(
		.INIT('h8)
	) name8169 (
		\wishbone_bd_ram_mem2_reg[28][16]/P0001 ,
		_w13170_,
		_w18681_
	);
	LUT2 #(
		.INIT('h8)
	) name8170 (
		\wishbone_bd_ram_mem2_reg[105][16]/P0001 ,
		_w12751_,
		_w18682_
	);
	LUT2 #(
		.INIT('h8)
	) name8171 (
		\wishbone_bd_ram_mem2_reg[252][16]/P0001 ,
		_w13080_,
		_w18683_
	);
	LUT2 #(
		.INIT('h8)
	) name8172 (
		\wishbone_bd_ram_mem2_reg[149][16]/P0001 ,
		_w12741_,
		_w18684_
	);
	LUT2 #(
		.INIT('h8)
	) name8173 (
		\wishbone_bd_ram_mem2_reg[229][16]/P0001 ,
		_w12711_,
		_w18685_
	);
	LUT2 #(
		.INIT('h8)
	) name8174 (
		\wishbone_bd_ram_mem2_reg[206][16]/P0001 ,
		_w12954_,
		_w18686_
	);
	LUT2 #(
		.INIT('h8)
	) name8175 (
		\wishbone_bd_ram_mem2_reg[239][16]/P0001 ,
		_w12862_,
		_w18687_
	);
	LUT2 #(
		.INIT('h8)
	) name8176 (
		\wishbone_bd_ram_mem2_reg[48][16]/P0001 ,
		_w12970_,
		_w18688_
	);
	LUT2 #(
		.INIT('h8)
	) name8177 (
		\wishbone_bd_ram_mem2_reg[244][16]/P0001 ,
		_w12747_,
		_w18689_
	);
	LUT2 #(
		.INIT('h8)
	) name8178 (
		\wishbone_bd_ram_mem2_reg[129][16]/P0001 ,
		_w12776_,
		_w18690_
	);
	LUT2 #(
		.INIT('h8)
	) name8179 (
		\wishbone_bd_ram_mem2_reg[242][16]/P0001 ,
		_w12932_,
		_w18691_
	);
	LUT2 #(
		.INIT('h8)
	) name8180 (
		\wishbone_bd_ram_mem2_reg[11][16]/P0001 ,
		_w13194_,
		_w18692_
	);
	LUT2 #(
		.INIT('h8)
	) name8181 (
		\wishbone_bd_ram_mem2_reg[170][16]/P0001 ,
		_w13030_,
		_w18693_
	);
	LUT2 #(
		.INIT('h8)
	) name8182 (
		\wishbone_bd_ram_mem2_reg[71][16]/P0001 ,
		_w12798_,
		_w18694_
	);
	LUT2 #(
		.INIT('h8)
	) name8183 (
		\wishbone_bd_ram_mem2_reg[52][16]/P0001 ,
		_w13082_,
		_w18695_
	);
	LUT2 #(
		.INIT('h8)
	) name8184 (
		\wishbone_bd_ram_mem2_reg[40][16]/P0001 ,
		_w13132_,
		_w18696_
	);
	LUT2 #(
		.INIT('h8)
	) name8185 (
		\wishbone_bd_ram_mem2_reg[19][16]/P0001 ,
		_w13012_,
		_w18697_
	);
	LUT2 #(
		.INIT('h8)
	) name8186 (
		\wishbone_bd_ram_mem2_reg[247][16]/P0001 ,
		_w12818_,
		_w18698_
	);
	LUT2 #(
		.INIT('h8)
	) name8187 (
		\wishbone_bd_ram_mem2_reg[192][16]/P0001 ,
		_w12938_,
		_w18699_
	);
	LUT2 #(
		.INIT('h8)
	) name8188 (
		\wishbone_bd_ram_mem2_reg[81][16]/P0001 ,
		_w12950_,
		_w18700_
	);
	LUT2 #(
		.INIT('h8)
	) name8189 (
		\wishbone_bd_ram_mem2_reg[41][16]/P0001 ,
		_w13052_,
		_w18701_
	);
	LUT2 #(
		.INIT('h8)
	) name8190 (
		\wishbone_bd_ram_mem2_reg[240][16]/P0001 ,
		_w12864_,
		_w18702_
	);
	LUT2 #(
		.INIT('h8)
	) name8191 (
		\wishbone_bd_ram_mem2_reg[143][16]/P0001 ,
		_w12922_,
		_w18703_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		\wishbone_bd_ram_mem2_reg[139][16]/P0001 ,
		_w12814_,
		_w18704_
	);
	LUT2 #(
		.INIT('h8)
	) name8193 (
		\wishbone_bd_ram_mem2_reg[180][16]/P0001 ,
		_w12791_,
		_w18705_
	);
	LUT2 #(
		.INIT('h8)
	) name8194 (
		\wishbone_bd_ram_mem2_reg[167][16]/P0001 ,
		_w12986_,
		_w18706_
	);
	LUT2 #(
		.INIT('h8)
	) name8195 (
		\wishbone_bd_ram_mem2_reg[113][16]/P0001 ,
		_w13026_,
		_w18707_
	);
	LUT2 #(
		.INIT('h8)
	) name8196 (
		\wishbone_bd_ram_mem2_reg[95][16]/P0001 ,
		_w12844_,
		_w18708_
	);
	LUT2 #(
		.INIT('h8)
	) name8197 (
		\wishbone_bd_ram_mem2_reg[225][16]/P0001 ,
		_w13092_,
		_w18709_
	);
	LUT2 #(
		.INIT('h8)
	) name8198 (
		\wishbone_bd_ram_mem2_reg[135][16]/P0001 ,
		_w13124_,
		_w18710_
	);
	LUT2 #(
		.INIT('h8)
	) name8199 (
		\wishbone_bd_ram_mem2_reg[199][16]/P0001 ,
		_w12768_,
		_w18711_
	);
	LUT2 #(
		.INIT('h8)
	) name8200 (
		\wishbone_bd_ram_mem2_reg[186][16]/P0001 ,
		_w12783_,
		_w18712_
	);
	LUT2 #(
		.INIT('h8)
	) name8201 (
		\wishbone_bd_ram_mem2_reg[60][16]/P0001 ,
		_w13204_,
		_w18713_
	);
	LUT2 #(
		.INIT('h8)
	) name8202 (
		\wishbone_bd_ram_mem2_reg[35][16]/P0001 ,
		_w12703_,
		_w18714_
	);
	LUT2 #(
		.INIT('h8)
	) name8203 (
		\wishbone_bd_ram_mem2_reg[89][16]/P0001 ,
		_w12964_,
		_w18715_
	);
	LUT2 #(
		.INIT('h8)
	) name8204 (
		\wishbone_bd_ram_mem2_reg[165][16]/P0001 ,
		_w13044_,
		_w18716_
	);
	LUT2 #(
		.INIT('h8)
	) name8205 (
		\wishbone_bd_ram_mem2_reg[26][16]/P0001 ,
		_w12699_,
		_w18717_
	);
	LUT2 #(
		.INIT('h8)
	) name8206 (
		\wishbone_bd_ram_mem2_reg[250][16]/P0001 ,
		_w13128_,
		_w18718_
	);
	LUT2 #(
		.INIT('h8)
	) name8207 (
		\wishbone_bd_ram_mem2_reg[82][16]/P0001 ,
		_w12942_,
		_w18719_
	);
	LUT2 #(
		.INIT('h8)
	) name8208 (
		\wishbone_bd_ram_mem2_reg[248][16]/P0001 ,
		_w12789_,
		_w18720_
	);
	LUT2 #(
		.INIT('h8)
	) name8209 (
		\wishbone_bd_ram_mem2_reg[15][16]/P0001 ,
		_w13210_,
		_w18721_
	);
	LUT2 #(
		.INIT('h8)
	) name8210 (
		\wishbone_bd_ram_mem2_reg[230][16]/P0001 ,
		_w13036_,
		_w18722_
	);
	LUT2 #(
		.INIT('h8)
	) name8211 (
		\wishbone_bd_ram_mem2_reg[189][16]/P0001 ,
		_w13042_,
		_w18723_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		\wishbone_bd_ram_mem2_reg[243][16]/P0001 ,
		_w12804_,
		_w18724_
	);
	LUT2 #(
		.INIT('h8)
	) name8213 (
		\wishbone_bd_ram_mem2_reg[65][16]/P0001 ,
		_w13176_,
		_w18725_
	);
	LUT2 #(
		.INIT('h8)
	) name8214 (
		\wishbone_bd_ram_mem2_reg[207][16]/P0001 ,
		_w13180_,
		_w18726_
	);
	LUT2 #(
		.INIT('h8)
	) name8215 (
		\wishbone_bd_ram_mem2_reg[142][16]/P0001 ,
		_w12928_,
		_w18727_
	);
	LUT2 #(
		.INIT('h8)
	) name8216 (
		\wishbone_bd_ram_mem2_reg[181][16]/P0001 ,
		_w12828_,
		_w18728_
	);
	LUT2 #(
		.INIT('h8)
	) name8217 (
		\wishbone_bd_ram_mem2_reg[249][16]/P0001 ,
		_w12900_,
		_w18729_
	);
	LUT2 #(
		.INIT('h8)
	) name8218 (
		\wishbone_bd_ram_mem2_reg[110][16]/P0001 ,
		_w13046_,
		_w18730_
	);
	LUT2 #(
		.INIT('h8)
	) name8219 (
		\wishbone_bd_ram_mem2_reg[63][16]/P0001 ,
		_w12850_,
		_w18731_
	);
	LUT2 #(
		.INIT('h8)
	) name8220 (
		\wishbone_bd_ram_mem2_reg[104][16]/P0001 ,
		_w13148_,
		_w18732_
	);
	LUT2 #(
		.INIT('h8)
	) name8221 (
		\wishbone_bd_ram_mem2_reg[25][16]/P0001 ,
		_w13108_,
		_w18733_
	);
	LUT2 #(
		.INIT('h8)
	) name8222 (
		\wishbone_bd_ram_mem2_reg[97][16]/P0001 ,
		_w13096_,
		_w18734_
	);
	LUT2 #(
		.INIT('h8)
	) name8223 (
		\wishbone_bd_ram_mem2_reg[251][16]/P0001 ,
		_w13054_,
		_w18735_
	);
	LUT2 #(
		.INIT('h8)
	) name8224 (
		\wishbone_bd_ram_mem2_reg[61][16]/P0001 ,
		_w12725_,
		_w18736_
	);
	LUT2 #(
		.INIT('h8)
	) name8225 (
		\wishbone_bd_ram_mem2_reg[209][16]/P0001 ,
		_w13152_,
		_w18737_
	);
	LUT2 #(
		.INIT('h8)
	) name8226 (
		\wishbone_bd_ram_mem2_reg[178][16]/P0001 ,
		_w12886_,
		_w18738_
	);
	LUT2 #(
		.INIT('h8)
	) name8227 (
		\wishbone_bd_ram_mem2_reg[205][16]/P0001 ,
		_w13068_,
		_w18739_
	);
	LUT2 #(
		.INIT('h8)
	) name8228 (
		\wishbone_bd_ram_mem2_reg[141][16]/P0001 ,
		_w13004_,
		_w18740_
	);
	LUT2 #(
		.INIT('h8)
	) name8229 (
		\wishbone_bd_ram_mem2_reg[76][16]/P0001 ,
		_w13184_,
		_w18741_
	);
	LUT2 #(
		.INIT('h8)
	) name8230 (
		\wishbone_bd_ram_mem2_reg[106][16]/P0001 ,
		_w12713_,
		_w18742_
	);
	LUT2 #(
		.INIT('h8)
	) name8231 (
		\wishbone_bd_ram_mem2_reg[228][16]/P0001 ,
		_w12765_,
		_w18743_
	);
	LUT2 #(
		.INIT('h8)
	) name8232 (
		\wishbone_bd_ram_mem2_reg[169][16]/P0001 ,
		_w12722_,
		_w18744_
	);
	LUT2 #(
		.INIT('h8)
	) name8233 (
		\wishbone_bd_ram_mem2_reg[195][16]/P0001 ,
		_w13144_,
		_w18745_
	);
	LUT2 #(
		.INIT('h8)
	) name8234 (
		\wishbone_bd_ram_mem2_reg[119][16]/P0001 ,
		_w13048_,
		_w18746_
	);
	LUT2 #(
		.INIT('h8)
	) name8235 (
		\wishbone_bd_ram_mem2_reg[171][16]/P0001 ,
		_w12910_,
		_w18747_
	);
	LUT2 #(
		.INIT('h8)
	) name8236 (
		\wishbone_bd_ram_mem2_reg[226][16]/P0001 ,
		_w13138_,
		_w18748_
	);
	LUT2 #(
		.INIT('h8)
	) name8237 (
		\wishbone_bd_ram_mem2_reg[140][16]/P0001 ,
		_w12894_,
		_w18749_
	);
	LUT2 #(
		.INIT('h8)
	) name8238 (
		\wishbone_bd_ram_mem2_reg[56][16]/P0001 ,
		_w12778_,
		_w18750_
	);
	LUT2 #(
		.INIT('h8)
	) name8239 (
		\wishbone_bd_ram_mem2_reg[175][16]/P0001 ,
		_w13126_,
		_w18751_
	);
	LUT2 #(
		.INIT('h8)
	) name8240 (
		\wishbone_bd_ram_mem2_reg[46][16]/P0001 ,
		_w12884_,
		_w18752_
	);
	LUT2 #(
		.INIT('h8)
	) name8241 (
		\wishbone_bd_ram_mem2_reg[92][16]/P0001 ,
		_w13010_,
		_w18753_
	);
	LUT2 #(
		.INIT('h8)
	) name8242 (
		\wishbone_bd_ram_mem2_reg[227][16]/P0001 ,
		_w12936_,
		_w18754_
	);
	LUT2 #(
		.INIT('h8)
	) name8243 (
		\wishbone_bd_ram_mem2_reg[245][16]/P0001 ,
		_w13022_,
		_w18755_
	);
	LUT2 #(
		.INIT('h8)
	) name8244 (
		\wishbone_bd_ram_mem2_reg[111][16]/P0001 ,
		_w12744_,
		_w18756_
	);
	LUT2 #(
		.INIT('h8)
	) name8245 (
		\wishbone_bd_ram_mem2_reg[201][16]/P0001 ,
		_w12822_,
		_w18757_
	);
	LUT2 #(
		.INIT('h8)
	) name8246 (
		\wishbone_bd_ram_mem2_reg[208][16]/P0001 ,
		_w13032_,
		_w18758_
	);
	LUT2 #(
		.INIT('h8)
	) name8247 (
		\wishbone_bd_ram_mem2_reg[29][16]/P0001 ,
		_w12952_,
		_w18759_
	);
	LUT2 #(
		.INIT('h8)
	) name8248 (
		\wishbone_bd_ram_mem2_reg[132][16]/P0001 ,
		_w12992_,
		_w18760_
	);
	LUT2 #(
		.INIT('h8)
	) name8249 (
		\wishbone_bd_ram_mem2_reg[212][16]/P0001 ,
		_w12796_,
		_w18761_
	);
	LUT2 #(
		.INIT('h8)
	) name8250 (
		\wishbone_bd_ram_mem2_reg[173][16]/P0001 ,
		_w12854_,
		_w18762_
	);
	LUT2 #(
		.INIT('h8)
	) name8251 (
		\wishbone_bd_ram_mem2_reg[43][16]/P0001 ,
		_w13200_,
		_w18763_
	);
	LUT2 #(
		.INIT('h8)
	) name8252 (
		\wishbone_bd_ram_mem2_reg[233][16]/P0001 ,
		_w12836_,
		_w18764_
	);
	LUT2 #(
		.INIT('h8)
	) name8253 (
		\wishbone_bd_ram_mem2_reg[12][16]/P0001 ,
		_w13118_,
		_w18765_
	);
	LUT2 #(
		.INIT('h8)
	) name8254 (
		\wishbone_bd_ram_mem2_reg[90][16]/P0001 ,
		_w12978_,
		_w18766_
	);
	LUT2 #(
		.INIT('h8)
	) name8255 (
		\wishbone_bd_ram_mem2_reg[85][16]/P0001 ,
		_w13216_,
		_w18767_
	);
	LUT2 #(
		.INIT('h8)
	) name8256 (
		\wishbone_bd_ram_mem2_reg[87][16]/P0001 ,
		_w13154_,
		_w18768_
	);
	LUT2 #(
		.INIT('h8)
	) name8257 (
		\wishbone_bd_ram_mem2_reg[22][16]/P0001 ,
		_w13110_,
		_w18769_
	);
	LUT2 #(
		.INIT('h8)
	) name8258 (
		\wishbone_bd_ram_mem2_reg[236][16]/P0001 ,
		_w12731_,
		_w18770_
	);
	LUT2 #(
		.INIT('h8)
	) name8259 (
		\wishbone_bd_ram_mem2_reg[255][16]/P0001 ,
		_w13072_,
		_w18771_
	);
	LUT2 #(
		.INIT('h8)
	) name8260 (
		\wishbone_bd_ram_mem2_reg[211][16]/P0001 ,
		_w13166_,
		_w18772_
	);
	LUT2 #(
		.INIT('h8)
	) name8261 (
		\wishbone_bd_ram_mem2_reg[50][16]/P0001 ,
		_w13150_,
		_w18773_
	);
	LUT2 #(
		.INIT('h8)
	) name8262 (
		\wishbone_bd_ram_mem2_reg[162][16]/P0001 ,
		_w13098_,
		_w18774_
	);
	LUT2 #(
		.INIT('h8)
	) name8263 (
		\wishbone_bd_ram_mem2_reg[157][16]/P0001 ,
		_w12926_,
		_w18775_
	);
	LUT2 #(
		.INIT('h8)
	) name8264 (
		\wishbone_bd_ram_mem2_reg[253][16]/P0001 ,
		_w13100_,
		_w18776_
	);
	LUT2 #(
		.INIT('h8)
	) name8265 (
		\wishbone_bd_ram_mem2_reg[156][16]/P0001 ,
		_w13190_,
		_w18777_
	);
	LUT2 #(
		.INIT('h8)
	) name8266 (
		\wishbone_bd_ram_mem2_reg[166][16]/P0001 ,
		_w13040_,
		_w18778_
	);
	LUT2 #(
		.INIT('h8)
	) name8267 (
		\wishbone_bd_ram_mem2_reg[53][16]/P0001 ,
		_w13020_,
		_w18779_
	);
	LUT2 #(
		.INIT('h8)
	) name8268 (
		\wishbone_bd_ram_mem2_reg[123][16]/P0001 ,
		_w13114_,
		_w18780_
	);
	LUT2 #(
		.INIT('h8)
	) name8269 (
		\wishbone_bd_ram_mem2_reg[72][16]/P0001 ,
		_w12810_,
		_w18781_
	);
	LUT2 #(
		.INIT('h8)
	) name8270 (
		\wishbone_bd_ram_mem2_reg[174][16]/P0001 ,
		_w12972_,
		_w18782_
	);
	LUT2 #(
		.INIT('h8)
	) name8271 (
		\wishbone_bd_ram_mem2_reg[27][16]/P0001 ,
		_w12880_,
		_w18783_
	);
	LUT2 #(
		.INIT('h8)
	) name8272 (
		\wishbone_bd_ram_mem2_reg[154][16]/P0001 ,
		_w12962_,
		_w18784_
	);
	LUT2 #(
		.INIT('h8)
	) name8273 (
		\wishbone_bd_ram_mem2_reg[18][16]/P0001 ,
		_w12679_,
		_w18785_
	);
	LUT2 #(
		.INIT('h8)
	) name8274 (
		\wishbone_bd_ram_mem2_reg[136][16]/P0001 ,
		_w13064_,
		_w18786_
	);
	LUT2 #(
		.INIT('h8)
	) name8275 (
		\wishbone_bd_ram_mem2_reg[152][16]/P0001 ,
		_w12966_,
		_w18787_
	);
	LUT2 #(
		.INIT('h8)
	) name8276 (
		\wishbone_bd_ram_mem2_reg[146][16]/P0001 ,
		_w13060_,
		_w18788_
	);
	LUT2 #(
		.INIT('h8)
	) name8277 (
		\wishbone_bd_ram_mem2_reg[3][16]/P0001 ,
		_w12866_,
		_w18789_
	);
	LUT2 #(
		.INIT('h8)
	) name8278 (
		\wishbone_bd_ram_mem2_reg[98][16]/P0001 ,
		_w12816_,
		_w18790_
	);
	LUT2 #(
		.INIT('h8)
	) name8279 (
		\wishbone_bd_ram_mem2_reg[168][16]/P0001 ,
		_w13208_,
		_w18791_
	);
	LUT2 #(
		.INIT('h8)
	) name8280 (
		\wishbone_bd_ram_mem2_reg[64][16]/P0001 ,
		_w12976_,
		_w18792_
	);
	LUT2 #(
		.INIT('h8)
	) name8281 (
		\wishbone_bd_ram_mem2_reg[215][16]/P0001 ,
		_w12974_,
		_w18793_
	);
	LUT2 #(
		.INIT('h8)
	) name8282 (
		\wishbone_bd_ram_mem2_reg[176][16]/P0001 ,
		_w12868_,
		_w18794_
	);
	LUT2 #(
		.INIT('h8)
	) name8283 (
		\wishbone_bd_ram_mem2_reg[37][16]/P0001 ,
		_w13102_,
		_w18795_
	);
	LUT2 #(
		.INIT('h8)
	) name8284 (
		\wishbone_bd_ram_mem2_reg[54][16]/P0001 ,
		_w12770_,
		_w18796_
	);
	LUT2 #(
		.INIT('h8)
	) name8285 (
		\wishbone_bd_ram_mem2_reg[51][16]/P0001 ,
		_w13024_,
		_w18797_
	);
	LUT2 #(
		.INIT('h8)
	) name8286 (
		\wishbone_bd_ram_mem2_reg[223][16]/P0001 ,
		_w12838_,
		_w18798_
	);
	LUT2 #(
		.INIT('h8)
	) name8287 (
		\wishbone_bd_ram_mem2_reg[9][16]/P0001 ,
		_w12808_,
		_w18799_
	);
	LUT2 #(
		.INIT('h8)
	) name8288 (
		\wishbone_bd_ram_mem2_reg[70][16]/P0001 ,
		_w12840_,
		_w18800_
	);
	LUT2 #(
		.INIT('h8)
	) name8289 (
		\wishbone_bd_ram_mem2_reg[222][16]/P0001 ,
		_w13094_,
		_w18801_
	);
	LUT2 #(
		.INIT('h8)
	) name8290 (
		\wishbone_bd_ram_mem2_reg[155][16]/P0001 ,
		_w13122_,
		_w18802_
	);
	LUT2 #(
		.INIT('h8)
	) name8291 (
		\wishbone_bd_ram_mem2_reg[78][16]/P0001 ,
		_w12874_,
		_w18803_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		\wishbone_bd_ram_mem2_reg[177][16]/P0001 ,
		_w12996_,
		_w18804_
	);
	LUT2 #(
		.INIT('h8)
	) name8293 (
		\wishbone_bd_ram_mem2_reg[187][16]/P0001 ,
		_w13196_,
		_w18805_
	);
	LUT2 #(
		.INIT('h8)
	) name8294 (
		\wishbone_bd_ram_mem2_reg[68][16]/P0001 ,
		_w12946_,
		_w18806_
	);
	LUT2 #(
		.INIT('h8)
	) name8295 (
		\wishbone_bd_ram_mem2_reg[66][16]/P0001 ,
		_w12824_,
		_w18807_
	);
	LUT2 #(
		.INIT('h8)
	) name8296 (
		\wishbone_bd_ram_mem2_reg[14][16]/P0001 ,
		_w13086_,
		_w18808_
	);
	LUT2 #(
		.INIT('h8)
	) name8297 (
		\wishbone_bd_ram_mem2_reg[232][16]/P0001 ,
		_w12758_,
		_w18809_
	);
	LUT2 #(
		.INIT('h8)
	) name8298 (
		\wishbone_bd_ram_mem2_reg[16][16]/P0001 ,
		_w13140_,
		_w18810_
	);
	LUT2 #(
		.INIT('h8)
	) name8299 (
		\wishbone_bd_ram_mem2_reg[109][16]/P0001 ,
		_w12888_,
		_w18811_
	);
	LUT2 #(
		.INIT('h8)
	) name8300 (
		\wishbone_bd_ram_mem2_reg[216][16]/P0001 ,
		_w13028_,
		_w18812_
	);
	LUT2 #(
		.INIT('h8)
	) name8301 (
		\wishbone_bd_ram_mem2_reg[238][16]/P0001 ,
		_w13160_,
		_w18813_
	);
	LUT2 #(
		.INIT('h8)
	) name8302 (
		\wishbone_bd_ram_mem2_reg[5][16]/P0001 ,
		_w12878_,
		_w18814_
	);
	LUT2 #(
		.INIT('h8)
	) name8303 (
		\wishbone_bd_ram_mem2_reg[133][16]/P0001 ,
		_w12761_,
		_w18815_
	);
	LUT2 #(
		.INIT('h8)
	) name8304 (
		\wishbone_bd_ram_mem2_reg[114][16]/P0001 ,
		_w13202_,
		_w18816_
	);
	LUT2 #(
		.INIT('h8)
	) name8305 (
		\wishbone_bd_ram_mem2_reg[84][16]/P0001 ,
		_w12934_,
		_w18817_
	);
	LUT2 #(
		.INIT('h8)
	) name8306 (
		\wishbone_bd_ram_mem2_reg[83][16]/P0001 ,
		_w12916_,
		_w18818_
	);
	LUT2 #(
		.INIT('h8)
	) name8307 (
		\wishbone_bd_ram_mem2_reg[179][16]/P0001 ,
		_w13050_,
		_w18819_
	);
	LUT2 #(
		.INIT('h8)
	) name8308 (
		\wishbone_bd_ram_mem2_reg[130][16]/P0001 ,
		_w12914_,
		_w18820_
	);
	LUT2 #(
		.INIT('h8)
	) name8309 (
		\wishbone_bd_ram_mem2_reg[4][16]/P0001 ,
		_w12666_,
		_w18821_
	);
	LUT2 #(
		.INIT('h8)
	) name8310 (
		\wishbone_bd_ram_mem2_reg[224][16]/P0001 ,
		_w12902_,
		_w18822_
	);
	LUT2 #(
		.INIT('h8)
	) name8311 (
		\wishbone_bd_ram_mem2_reg[107][16]/P0001 ,
		_w12749_,
		_w18823_
	);
	LUT2 #(
		.INIT('h8)
	) name8312 (
		\wishbone_bd_ram_mem2_reg[145][16]/P0001 ,
		_w13106_,
		_w18824_
	);
	LUT2 #(
		.INIT('h8)
	) name8313 (
		\wishbone_bd_ram_mem2_reg[210][16]/P0001 ,
		_w12924_,
		_w18825_
	);
	LUT2 #(
		.INIT('h8)
	) name8314 (
		\wishbone_bd_ram_mem2_reg[198][16]/P0001 ,
		_w12832_,
		_w18826_
	);
	LUT2 #(
		.INIT('h8)
	) name8315 (
		\wishbone_bd_ram_mem2_reg[153][16]/P0001 ,
		_w12890_,
		_w18827_
	);
	LUT2 #(
		.INIT('h8)
	) name8316 (
		\wishbone_bd_ram_mem2_reg[131][16]/P0001 ,
		_w12852_,
		_w18828_
	);
	LUT2 #(
		.INIT('h8)
	) name8317 (
		\wishbone_bd_ram_mem2_reg[94][16]/P0001 ,
		_w13186_,
		_w18829_
	);
	LUT2 #(
		.INIT('h8)
	) name8318 (
		\wishbone_bd_ram_mem2_reg[217][16]/P0001 ,
		_w13188_,
		_w18830_
	);
	LUT2 #(
		.INIT('h8)
	) name8319 (
		\wishbone_bd_ram_mem2_reg[144][16]/P0001 ,
		_w12756_,
		_w18831_
	);
	LUT2 #(
		.INIT('h8)
	) name8320 (
		\wishbone_bd_ram_mem2_reg[73][16]/P0001 ,
		_w12918_,
		_w18832_
	);
	LUT2 #(
		.INIT('h1)
	) name8321 (
		_w18577_,
		_w18578_,
		_w18833_
	);
	LUT2 #(
		.INIT('h1)
	) name8322 (
		_w18579_,
		_w18580_,
		_w18834_
	);
	LUT2 #(
		.INIT('h1)
	) name8323 (
		_w18581_,
		_w18582_,
		_w18835_
	);
	LUT2 #(
		.INIT('h1)
	) name8324 (
		_w18583_,
		_w18584_,
		_w18836_
	);
	LUT2 #(
		.INIT('h1)
	) name8325 (
		_w18585_,
		_w18586_,
		_w18837_
	);
	LUT2 #(
		.INIT('h1)
	) name8326 (
		_w18587_,
		_w18588_,
		_w18838_
	);
	LUT2 #(
		.INIT('h1)
	) name8327 (
		_w18589_,
		_w18590_,
		_w18839_
	);
	LUT2 #(
		.INIT('h1)
	) name8328 (
		_w18591_,
		_w18592_,
		_w18840_
	);
	LUT2 #(
		.INIT('h1)
	) name8329 (
		_w18593_,
		_w18594_,
		_w18841_
	);
	LUT2 #(
		.INIT('h1)
	) name8330 (
		_w18595_,
		_w18596_,
		_w18842_
	);
	LUT2 #(
		.INIT('h1)
	) name8331 (
		_w18597_,
		_w18598_,
		_w18843_
	);
	LUT2 #(
		.INIT('h1)
	) name8332 (
		_w18599_,
		_w18600_,
		_w18844_
	);
	LUT2 #(
		.INIT('h1)
	) name8333 (
		_w18601_,
		_w18602_,
		_w18845_
	);
	LUT2 #(
		.INIT('h1)
	) name8334 (
		_w18603_,
		_w18604_,
		_w18846_
	);
	LUT2 #(
		.INIT('h1)
	) name8335 (
		_w18605_,
		_w18606_,
		_w18847_
	);
	LUT2 #(
		.INIT('h1)
	) name8336 (
		_w18607_,
		_w18608_,
		_w18848_
	);
	LUT2 #(
		.INIT('h1)
	) name8337 (
		_w18609_,
		_w18610_,
		_w18849_
	);
	LUT2 #(
		.INIT('h1)
	) name8338 (
		_w18611_,
		_w18612_,
		_w18850_
	);
	LUT2 #(
		.INIT('h1)
	) name8339 (
		_w18613_,
		_w18614_,
		_w18851_
	);
	LUT2 #(
		.INIT('h1)
	) name8340 (
		_w18615_,
		_w18616_,
		_w18852_
	);
	LUT2 #(
		.INIT('h1)
	) name8341 (
		_w18617_,
		_w18618_,
		_w18853_
	);
	LUT2 #(
		.INIT('h1)
	) name8342 (
		_w18619_,
		_w18620_,
		_w18854_
	);
	LUT2 #(
		.INIT('h1)
	) name8343 (
		_w18621_,
		_w18622_,
		_w18855_
	);
	LUT2 #(
		.INIT('h1)
	) name8344 (
		_w18623_,
		_w18624_,
		_w18856_
	);
	LUT2 #(
		.INIT('h1)
	) name8345 (
		_w18625_,
		_w18626_,
		_w18857_
	);
	LUT2 #(
		.INIT('h1)
	) name8346 (
		_w18627_,
		_w18628_,
		_w18858_
	);
	LUT2 #(
		.INIT('h1)
	) name8347 (
		_w18629_,
		_w18630_,
		_w18859_
	);
	LUT2 #(
		.INIT('h1)
	) name8348 (
		_w18631_,
		_w18632_,
		_w18860_
	);
	LUT2 #(
		.INIT('h1)
	) name8349 (
		_w18633_,
		_w18634_,
		_w18861_
	);
	LUT2 #(
		.INIT('h1)
	) name8350 (
		_w18635_,
		_w18636_,
		_w18862_
	);
	LUT2 #(
		.INIT('h1)
	) name8351 (
		_w18637_,
		_w18638_,
		_w18863_
	);
	LUT2 #(
		.INIT('h1)
	) name8352 (
		_w18639_,
		_w18640_,
		_w18864_
	);
	LUT2 #(
		.INIT('h1)
	) name8353 (
		_w18641_,
		_w18642_,
		_w18865_
	);
	LUT2 #(
		.INIT('h1)
	) name8354 (
		_w18643_,
		_w18644_,
		_w18866_
	);
	LUT2 #(
		.INIT('h1)
	) name8355 (
		_w18645_,
		_w18646_,
		_w18867_
	);
	LUT2 #(
		.INIT('h1)
	) name8356 (
		_w18647_,
		_w18648_,
		_w18868_
	);
	LUT2 #(
		.INIT('h1)
	) name8357 (
		_w18649_,
		_w18650_,
		_w18869_
	);
	LUT2 #(
		.INIT('h1)
	) name8358 (
		_w18651_,
		_w18652_,
		_w18870_
	);
	LUT2 #(
		.INIT('h1)
	) name8359 (
		_w18653_,
		_w18654_,
		_w18871_
	);
	LUT2 #(
		.INIT('h1)
	) name8360 (
		_w18655_,
		_w18656_,
		_w18872_
	);
	LUT2 #(
		.INIT('h1)
	) name8361 (
		_w18657_,
		_w18658_,
		_w18873_
	);
	LUT2 #(
		.INIT('h1)
	) name8362 (
		_w18659_,
		_w18660_,
		_w18874_
	);
	LUT2 #(
		.INIT('h1)
	) name8363 (
		_w18661_,
		_w18662_,
		_w18875_
	);
	LUT2 #(
		.INIT('h1)
	) name8364 (
		_w18663_,
		_w18664_,
		_w18876_
	);
	LUT2 #(
		.INIT('h1)
	) name8365 (
		_w18665_,
		_w18666_,
		_w18877_
	);
	LUT2 #(
		.INIT('h1)
	) name8366 (
		_w18667_,
		_w18668_,
		_w18878_
	);
	LUT2 #(
		.INIT('h1)
	) name8367 (
		_w18669_,
		_w18670_,
		_w18879_
	);
	LUT2 #(
		.INIT('h1)
	) name8368 (
		_w18671_,
		_w18672_,
		_w18880_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w18673_,
		_w18674_,
		_w18881_
	);
	LUT2 #(
		.INIT('h1)
	) name8370 (
		_w18675_,
		_w18676_,
		_w18882_
	);
	LUT2 #(
		.INIT('h1)
	) name8371 (
		_w18677_,
		_w18678_,
		_w18883_
	);
	LUT2 #(
		.INIT('h1)
	) name8372 (
		_w18679_,
		_w18680_,
		_w18884_
	);
	LUT2 #(
		.INIT('h1)
	) name8373 (
		_w18681_,
		_w18682_,
		_w18885_
	);
	LUT2 #(
		.INIT('h1)
	) name8374 (
		_w18683_,
		_w18684_,
		_w18886_
	);
	LUT2 #(
		.INIT('h1)
	) name8375 (
		_w18685_,
		_w18686_,
		_w18887_
	);
	LUT2 #(
		.INIT('h1)
	) name8376 (
		_w18687_,
		_w18688_,
		_w18888_
	);
	LUT2 #(
		.INIT('h1)
	) name8377 (
		_w18689_,
		_w18690_,
		_w18889_
	);
	LUT2 #(
		.INIT('h1)
	) name8378 (
		_w18691_,
		_w18692_,
		_w18890_
	);
	LUT2 #(
		.INIT('h1)
	) name8379 (
		_w18693_,
		_w18694_,
		_w18891_
	);
	LUT2 #(
		.INIT('h1)
	) name8380 (
		_w18695_,
		_w18696_,
		_w18892_
	);
	LUT2 #(
		.INIT('h1)
	) name8381 (
		_w18697_,
		_w18698_,
		_w18893_
	);
	LUT2 #(
		.INIT('h1)
	) name8382 (
		_w18699_,
		_w18700_,
		_w18894_
	);
	LUT2 #(
		.INIT('h1)
	) name8383 (
		_w18701_,
		_w18702_,
		_w18895_
	);
	LUT2 #(
		.INIT('h1)
	) name8384 (
		_w18703_,
		_w18704_,
		_w18896_
	);
	LUT2 #(
		.INIT('h1)
	) name8385 (
		_w18705_,
		_w18706_,
		_w18897_
	);
	LUT2 #(
		.INIT('h1)
	) name8386 (
		_w18707_,
		_w18708_,
		_w18898_
	);
	LUT2 #(
		.INIT('h1)
	) name8387 (
		_w18709_,
		_w18710_,
		_w18899_
	);
	LUT2 #(
		.INIT('h1)
	) name8388 (
		_w18711_,
		_w18712_,
		_w18900_
	);
	LUT2 #(
		.INIT('h1)
	) name8389 (
		_w18713_,
		_w18714_,
		_w18901_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w18715_,
		_w18716_,
		_w18902_
	);
	LUT2 #(
		.INIT('h1)
	) name8391 (
		_w18717_,
		_w18718_,
		_w18903_
	);
	LUT2 #(
		.INIT('h1)
	) name8392 (
		_w18719_,
		_w18720_,
		_w18904_
	);
	LUT2 #(
		.INIT('h1)
	) name8393 (
		_w18721_,
		_w18722_,
		_w18905_
	);
	LUT2 #(
		.INIT('h1)
	) name8394 (
		_w18723_,
		_w18724_,
		_w18906_
	);
	LUT2 #(
		.INIT('h1)
	) name8395 (
		_w18725_,
		_w18726_,
		_w18907_
	);
	LUT2 #(
		.INIT('h1)
	) name8396 (
		_w18727_,
		_w18728_,
		_w18908_
	);
	LUT2 #(
		.INIT('h1)
	) name8397 (
		_w18729_,
		_w18730_,
		_w18909_
	);
	LUT2 #(
		.INIT('h1)
	) name8398 (
		_w18731_,
		_w18732_,
		_w18910_
	);
	LUT2 #(
		.INIT('h1)
	) name8399 (
		_w18733_,
		_w18734_,
		_w18911_
	);
	LUT2 #(
		.INIT('h1)
	) name8400 (
		_w18735_,
		_w18736_,
		_w18912_
	);
	LUT2 #(
		.INIT('h1)
	) name8401 (
		_w18737_,
		_w18738_,
		_w18913_
	);
	LUT2 #(
		.INIT('h1)
	) name8402 (
		_w18739_,
		_w18740_,
		_w18914_
	);
	LUT2 #(
		.INIT('h1)
	) name8403 (
		_w18741_,
		_w18742_,
		_w18915_
	);
	LUT2 #(
		.INIT('h1)
	) name8404 (
		_w18743_,
		_w18744_,
		_w18916_
	);
	LUT2 #(
		.INIT('h1)
	) name8405 (
		_w18745_,
		_w18746_,
		_w18917_
	);
	LUT2 #(
		.INIT('h1)
	) name8406 (
		_w18747_,
		_w18748_,
		_w18918_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		_w18749_,
		_w18750_,
		_w18919_
	);
	LUT2 #(
		.INIT('h1)
	) name8408 (
		_w18751_,
		_w18752_,
		_w18920_
	);
	LUT2 #(
		.INIT('h1)
	) name8409 (
		_w18753_,
		_w18754_,
		_w18921_
	);
	LUT2 #(
		.INIT('h1)
	) name8410 (
		_w18755_,
		_w18756_,
		_w18922_
	);
	LUT2 #(
		.INIT('h1)
	) name8411 (
		_w18757_,
		_w18758_,
		_w18923_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		_w18759_,
		_w18760_,
		_w18924_
	);
	LUT2 #(
		.INIT('h1)
	) name8413 (
		_w18761_,
		_w18762_,
		_w18925_
	);
	LUT2 #(
		.INIT('h1)
	) name8414 (
		_w18763_,
		_w18764_,
		_w18926_
	);
	LUT2 #(
		.INIT('h1)
	) name8415 (
		_w18765_,
		_w18766_,
		_w18927_
	);
	LUT2 #(
		.INIT('h1)
	) name8416 (
		_w18767_,
		_w18768_,
		_w18928_
	);
	LUT2 #(
		.INIT('h1)
	) name8417 (
		_w18769_,
		_w18770_,
		_w18929_
	);
	LUT2 #(
		.INIT('h1)
	) name8418 (
		_w18771_,
		_w18772_,
		_w18930_
	);
	LUT2 #(
		.INIT('h1)
	) name8419 (
		_w18773_,
		_w18774_,
		_w18931_
	);
	LUT2 #(
		.INIT('h1)
	) name8420 (
		_w18775_,
		_w18776_,
		_w18932_
	);
	LUT2 #(
		.INIT('h1)
	) name8421 (
		_w18777_,
		_w18778_,
		_w18933_
	);
	LUT2 #(
		.INIT('h1)
	) name8422 (
		_w18779_,
		_w18780_,
		_w18934_
	);
	LUT2 #(
		.INIT('h1)
	) name8423 (
		_w18781_,
		_w18782_,
		_w18935_
	);
	LUT2 #(
		.INIT('h1)
	) name8424 (
		_w18783_,
		_w18784_,
		_w18936_
	);
	LUT2 #(
		.INIT('h1)
	) name8425 (
		_w18785_,
		_w18786_,
		_w18937_
	);
	LUT2 #(
		.INIT('h1)
	) name8426 (
		_w18787_,
		_w18788_,
		_w18938_
	);
	LUT2 #(
		.INIT('h1)
	) name8427 (
		_w18789_,
		_w18790_,
		_w18939_
	);
	LUT2 #(
		.INIT('h1)
	) name8428 (
		_w18791_,
		_w18792_,
		_w18940_
	);
	LUT2 #(
		.INIT('h1)
	) name8429 (
		_w18793_,
		_w18794_,
		_w18941_
	);
	LUT2 #(
		.INIT('h1)
	) name8430 (
		_w18795_,
		_w18796_,
		_w18942_
	);
	LUT2 #(
		.INIT('h1)
	) name8431 (
		_w18797_,
		_w18798_,
		_w18943_
	);
	LUT2 #(
		.INIT('h1)
	) name8432 (
		_w18799_,
		_w18800_,
		_w18944_
	);
	LUT2 #(
		.INIT('h1)
	) name8433 (
		_w18801_,
		_w18802_,
		_w18945_
	);
	LUT2 #(
		.INIT('h1)
	) name8434 (
		_w18803_,
		_w18804_,
		_w18946_
	);
	LUT2 #(
		.INIT('h1)
	) name8435 (
		_w18805_,
		_w18806_,
		_w18947_
	);
	LUT2 #(
		.INIT('h1)
	) name8436 (
		_w18807_,
		_w18808_,
		_w18948_
	);
	LUT2 #(
		.INIT('h1)
	) name8437 (
		_w18809_,
		_w18810_,
		_w18949_
	);
	LUT2 #(
		.INIT('h1)
	) name8438 (
		_w18811_,
		_w18812_,
		_w18950_
	);
	LUT2 #(
		.INIT('h1)
	) name8439 (
		_w18813_,
		_w18814_,
		_w18951_
	);
	LUT2 #(
		.INIT('h1)
	) name8440 (
		_w18815_,
		_w18816_,
		_w18952_
	);
	LUT2 #(
		.INIT('h1)
	) name8441 (
		_w18817_,
		_w18818_,
		_w18953_
	);
	LUT2 #(
		.INIT('h1)
	) name8442 (
		_w18819_,
		_w18820_,
		_w18954_
	);
	LUT2 #(
		.INIT('h1)
	) name8443 (
		_w18821_,
		_w18822_,
		_w18955_
	);
	LUT2 #(
		.INIT('h1)
	) name8444 (
		_w18823_,
		_w18824_,
		_w18956_
	);
	LUT2 #(
		.INIT('h1)
	) name8445 (
		_w18825_,
		_w18826_,
		_w18957_
	);
	LUT2 #(
		.INIT('h1)
	) name8446 (
		_w18827_,
		_w18828_,
		_w18958_
	);
	LUT2 #(
		.INIT('h1)
	) name8447 (
		_w18829_,
		_w18830_,
		_w18959_
	);
	LUT2 #(
		.INIT('h1)
	) name8448 (
		_w18831_,
		_w18832_,
		_w18960_
	);
	LUT2 #(
		.INIT('h8)
	) name8449 (
		_w18959_,
		_w18960_,
		_w18961_
	);
	LUT2 #(
		.INIT('h8)
	) name8450 (
		_w18957_,
		_w18958_,
		_w18962_
	);
	LUT2 #(
		.INIT('h8)
	) name8451 (
		_w18955_,
		_w18956_,
		_w18963_
	);
	LUT2 #(
		.INIT('h8)
	) name8452 (
		_w18953_,
		_w18954_,
		_w18964_
	);
	LUT2 #(
		.INIT('h8)
	) name8453 (
		_w18951_,
		_w18952_,
		_w18965_
	);
	LUT2 #(
		.INIT('h8)
	) name8454 (
		_w18949_,
		_w18950_,
		_w18966_
	);
	LUT2 #(
		.INIT('h8)
	) name8455 (
		_w18947_,
		_w18948_,
		_w18967_
	);
	LUT2 #(
		.INIT('h8)
	) name8456 (
		_w18945_,
		_w18946_,
		_w18968_
	);
	LUT2 #(
		.INIT('h8)
	) name8457 (
		_w18943_,
		_w18944_,
		_w18969_
	);
	LUT2 #(
		.INIT('h8)
	) name8458 (
		_w18941_,
		_w18942_,
		_w18970_
	);
	LUT2 #(
		.INIT('h8)
	) name8459 (
		_w18939_,
		_w18940_,
		_w18971_
	);
	LUT2 #(
		.INIT('h8)
	) name8460 (
		_w18937_,
		_w18938_,
		_w18972_
	);
	LUT2 #(
		.INIT('h8)
	) name8461 (
		_w18935_,
		_w18936_,
		_w18973_
	);
	LUT2 #(
		.INIT('h8)
	) name8462 (
		_w18933_,
		_w18934_,
		_w18974_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		_w18931_,
		_w18932_,
		_w18975_
	);
	LUT2 #(
		.INIT('h8)
	) name8464 (
		_w18929_,
		_w18930_,
		_w18976_
	);
	LUT2 #(
		.INIT('h8)
	) name8465 (
		_w18927_,
		_w18928_,
		_w18977_
	);
	LUT2 #(
		.INIT('h8)
	) name8466 (
		_w18925_,
		_w18926_,
		_w18978_
	);
	LUT2 #(
		.INIT('h8)
	) name8467 (
		_w18923_,
		_w18924_,
		_w18979_
	);
	LUT2 #(
		.INIT('h8)
	) name8468 (
		_w18921_,
		_w18922_,
		_w18980_
	);
	LUT2 #(
		.INIT('h8)
	) name8469 (
		_w18919_,
		_w18920_,
		_w18981_
	);
	LUT2 #(
		.INIT('h8)
	) name8470 (
		_w18917_,
		_w18918_,
		_w18982_
	);
	LUT2 #(
		.INIT('h8)
	) name8471 (
		_w18915_,
		_w18916_,
		_w18983_
	);
	LUT2 #(
		.INIT('h8)
	) name8472 (
		_w18913_,
		_w18914_,
		_w18984_
	);
	LUT2 #(
		.INIT('h8)
	) name8473 (
		_w18911_,
		_w18912_,
		_w18985_
	);
	LUT2 #(
		.INIT('h8)
	) name8474 (
		_w18909_,
		_w18910_,
		_w18986_
	);
	LUT2 #(
		.INIT('h8)
	) name8475 (
		_w18907_,
		_w18908_,
		_w18987_
	);
	LUT2 #(
		.INIT('h8)
	) name8476 (
		_w18905_,
		_w18906_,
		_w18988_
	);
	LUT2 #(
		.INIT('h8)
	) name8477 (
		_w18903_,
		_w18904_,
		_w18989_
	);
	LUT2 #(
		.INIT('h8)
	) name8478 (
		_w18901_,
		_w18902_,
		_w18990_
	);
	LUT2 #(
		.INIT('h8)
	) name8479 (
		_w18899_,
		_w18900_,
		_w18991_
	);
	LUT2 #(
		.INIT('h8)
	) name8480 (
		_w18897_,
		_w18898_,
		_w18992_
	);
	LUT2 #(
		.INIT('h8)
	) name8481 (
		_w18895_,
		_w18896_,
		_w18993_
	);
	LUT2 #(
		.INIT('h8)
	) name8482 (
		_w18893_,
		_w18894_,
		_w18994_
	);
	LUT2 #(
		.INIT('h8)
	) name8483 (
		_w18891_,
		_w18892_,
		_w18995_
	);
	LUT2 #(
		.INIT('h8)
	) name8484 (
		_w18889_,
		_w18890_,
		_w18996_
	);
	LUT2 #(
		.INIT('h8)
	) name8485 (
		_w18887_,
		_w18888_,
		_w18997_
	);
	LUT2 #(
		.INIT('h8)
	) name8486 (
		_w18885_,
		_w18886_,
		_w18998_
	);
	LUT2 #(
		.INIT('h8)
	) name8487 (
		_w18883_,
		_w18884_,
		_w18999_
	);
	LUT2 #(
		.INIT('h8)
	) name8488 (
		_w18881_,
		_w18882_,
		_w19000_
	);
	LUT2 #(
		.INIT('h8)
	) name8489 (
		_w18879_,
		_w18880_,
		_w19001_
	);
	LUT2 #(
		.INIT('h8)
	) name8490 (
		_w18877_,
		_w18878_,
		_w19002_
	);
	LUT2 #(
		.INIT('h8)
	) name8491 (
		_w18875_,
		_w18876_,
		_w19003_
	);
	LUT2 #(
		.INIT('h8)
	) name8492 (
		_w18873_,
		_w18874_,
		_w19004_
	);
	LUT2 #(
		.INIT('h8)
	) name8493 (
		_w18871_,
		_w18872_,
		_w19005_
	);
	LUT2 #(
		.INIT('h8)
	) name8494 (
		_w18869_,
		_w18870_,
		_w19006_
	);
	LUT2 #(
		.INIT('h8)
	) name8495 (
		_w18867_,
		_w18868_,
		_w19007_
	);
	LUT2 #(
		.INIT('h8)
	) name8496 (
		_w18865_,
		_w18866_,
		_w19008_
	);
	LUT2 #(
		.INIT('h8)
	) name8497 (
		_w18863_,
		_w18864_,
		_w19009_
	);
	LUT2 #(
		.INIT('h8)
	) name8498 (
		_w18861_,
		_w18862_,
		_w19010_
	);
	LUT2 #(
		.INIT('h8)
	) name8499 (
		_w18859_,
		_w18860_,
		_w19011_
	);
	LUT2 #(
		.INIT('h8)
	) name8500 (
		_w18857_,
		_w18858_,
		_w19012_
	);
	LUT2 #(
		.INIT('h8)
	) name8501 (
		_w18855_,
		_w18856_,
		_w19013_
	);
	LUT2 #(
		.INIT('h8)
	) name8502 (
		_w18853_,
		_w18854_,
		_w19014_
	);
	LUT2 #(
		.INIT('h8)
	) name8503 (
		_w18851_,
		_w18852_,
		_w19015_
	);
	LUT2 #(
		.INIT('h8)
	) name8504 (
		_w18849_,
		_w18850_,
		_w19016_
	);
	LUT2 #(
		.INIT('h8)
	) name8505 (
		_w18847_,
		_w18848_,
		_w19017_
	);
	LUT2 #(
		.INIT('h8)
	) name8506 (
		_w18845_,
		_w18846_,
		_w19018_
	);
	LUT2 #(
		.INIT('h8)
	) name8507 (
		_w18843_,
		_w18844_,
		_w19019_
	);
	LUT2 #(
		.INIT('h8)
	) name8508 (
		_w18841_,
		_w18842_,
		_w19020_
	);
	LUT2 #(
		.INIT('h8)
	) name8509 (
		_w18839_,
		_w18840_,
		_w19021_
	);
	LUT2 #(
		.INIT('h8)
	) name8510 (
		_w18837_,
		_w18838_,
		_w19022_
	);
	LUT2 #(
		.INIT('h8)
	) name8511 (
		_w18835_,
		_w18836_,
		_w19023_
	);
	LUT2 #(
		.INIT('h8)
	) name8512 (
		_w18833_,
		_w18834_,
		_w19024_
	);
	LUT2 #(
		.INIT('h8)
	) name8513 (
		_w19023_,
		_w19024_,
		_w19025_
	);
	LUT2 #(
		.INIT('h8)
	) name8514 (
		_w19021_,
		_w19022_,
		_w19026_
	);
	LUT2 #(
		.INIT('h8)
	) name8515 (
		_w19019_,
		_w19020_,
		_w19027_
	);
	LUT2 #(
		.INIT('h8)
	) name8516 (
		_w19017_,
		_w19018_,
		_w19028_
	);
	LUT2 #(
		.INIT('h8)
	) name8517 (
		_w19015_,
		_w19016_,
		_w19029_
	);
	LUT2 #(
		.INIT('h8)
	) name8518 (
		_w19013_,
		_w19014_,
		_w19030_
	);
	LUT2 #(
		.INIT('h8)
	) name8519 (
		_w19011_,
		_w19012_,
		_w19031_
	);
	LUT2 #(
		.INIT('h8)
	) name8520 (
		_w19009_,
		_w19010_,
		_w19032_
	);
	LUT2 #(
		.INIT('h8)
	) name8521 (
		_w19007_,
		_w19008_,
		_w19033_
	);
	LUT2 #(
		.INIT('h8)
	) name8522 (
		_w19005_,
		_w19006_,
		_w19034_
	);
	LUT2 #(
		.INIT('h8)
	) name8523 (
		_w19003_,
		_w19004_,
		_w19035_
	);
	LUT2 #(
		.INIT('h8)
	) name8524 (
		_w19001_,
		_w19002_,
		_w19036_
	);
	LUT2 #(
		.INIT('h8)
	) name8525 (
		_w18999_,
		_w19000_,
		_w19037_
	);
	LUT2 #(
		.INIT('h8)
	) name8526 (
		_w18997_,
		_w18998_,
		_w19038_
	);
	LUT2 #(
		.INIT('h8)
	) name8527 (
		_w18995_,
		_w18996_,
		_w19039_
	);
	LUT2 #(
		.INIT('h8)
	) name8528 (
		_w18993_,
		_w18994_,
		_w19040_
	);
	LUT2 #(
		.INIT('h8)
	) name8529 (
		_w18991_,
		_w18992_,
		_w19041_
	);
	LUT2 #(
		.INIT('h8)
	) name8530 (
		_w18989_,
		_w18990_,
		_w19042_
	);
	LUT2 #(
		.INIT('h8)
	) name8531 (
		_w18987_,
		_w18988_,
		_w19043_
	);
	LUT2 #(
		.INIT('h8)
	) name8532 (
		_w18985_,
		_w18986_,
		_w19044_
	);
	LUT2 #(
		.INIT('h8)
	) name8533 (
		_w18983_,
		_w18984_,
		_w19045_
	);
	LUT2 #(
		.INIT('h8)
	) name8534 (
		_w18981_,
		_w18982_,
		_w19046_
	);
	LUT2 #(
		.INIT('h8)
	) name8535 (
		_w18979_,
		_w18980_,
		_w19047_
	);
	LUT2 #(
		.INIT('h8)
	) name8536 (
		_w18977_,
		_w18978_,
		_w19048_
	);
	LUT2 #(
		.INIT('h8)
	) name8537 (
		_w18975_,
		_w18976_,
		_w19049_
	);
	LUT2 #(
		.INIT('h8)
	) name8538 (
		_w18973_,
		_w18974_,
		_w19050_
	);
	LUT2 #(
		.INIT('h8)
	) name8539 (
		_w18971_,
		_w18972_,
		_w19051_
	);
	LUT2 #(
		.INIT('h8)
	) name8540 (
		_w18969_,
		_w18970_,
		_w19052_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		_w18967_,
		_w18968_,
		_w19053_
	);
	LUT2 #(
		.INIT('h8)
	) name8542 (
		_w18965_,
		_w18966_,
		_w19054_
	);
	LUT2 #(
		.INIT('h8)
	) name8543 (
		_w18963_,
		_w18964_,
		_w19055_
	);
	LUT2 #(
		.INIT('h8)
	) name8544 (
		_w18961_,
		_w18962_,
		_w19056_
	);
	LUT2 #(
		.INIT('h8)
	) name8545 (
		_w19055_,
		_w19056_,
		_w19057_
	);
	LUT2 #(
		.INIT('h8)
	) name8546 (
		_w19053_,
		_w19054_,
		_w19058_
	);
	LUT2 #(
		.INIT('h8)
	) name8547 (
		_w19051_,
		_w19052_,
		_w19059_
	);
	LUT2 #(
		.INIT('h8)
	) name8548 (
		_w19049_,
		_w19050_,
		_w19060_
	);
	LUT2 #(
		.INIT('h8)
	) name8549 (
		_w19047_,
		_w19048_,
		_w19061_
	);
	LUT2 #(
		.INIT('h8)
	) name8550 (
		_w19045_,
		_w19046_,
		_w19062_
	);
	LUT2 #(
		.INIT('h8)
	) name8551 (
		_w19043_,
		_w19044_,
		_w19063_
	);
	LUT2 #(
		.INIT('h8)
	) name8552 (
		_w19041_,
		_w19042_,
		_w19064_
	);
	LUT2 #(
		.INIT('h8)
	) name8553 (
		_w19039_,
		_w19040_,
		_w19065_
	);
	LUT2 #(
		.INIT('h8)
	) name8554 (
		_w19037_,
		_w19038_,
		_w19066_
	);
	LUT2 #(
		.INIT('h8)
	) name8555 (
		_w19035_,
		_w19036_,
		_w19067_
	);
	LUT2 #(
		.INIT('h8)
	) name8556 (
		_w19033_,
		_w19034_,
		_w19068_
	);
	LUT2 #(
		.INIT('h8)
	) name8557 (
		_w19031_,
		_w19032_,
		_w19069_
	);
	LUT2 #(
		.INIT('h8)
	) name8558 (
		_w19029_,
		_w19030_,
		_w19070_
	);
	LUT2 #(
		.INIT('h8)
	) name8559 (
		_w19027_,
		_w19028_,
		_w19071_
	);
	LUT2 #(
		.INIT('h8)
	) name8560 (
		_w19025_,
		_w19026_,
		_w19072_
	);
	LUT2 #(
		.INIT('h8)
	) name8561 (
		_w19071_,
		_w19072_,
		_w19073_
	);
	LUT2 #(
		.INIT('h8)
	) name8562 (
		_w19069_,
		_w19070_,
		_w19074_
	);
	LUT2 #(
		.INIT('h8)
	) name8563 (
		_w19067_,
		_w19068_,
		_w19075_
	);
	LUT2 #(
		.INIT('h8)
	) name8564 (
		_w19065_,
		_w19066_,
		_w19076_
	);
	LUT2 #(
		.INIT('h8)
	) name8565 (
		_w19063_,
		_w19064_,
		_w19077_
	);
	LUT2 #(
		.INIT('h8)
	) name8566 (
		_w19061_,
		_w19062_,
		_w19078_
	);
	LUT2 #(
		.INIT('h8)
	) name8567 (
		_w19059_,
		_w19060_,
		_w19079_
	);
	LUT2 #(
		.INIT('h8)
	) name8568 (
		_w19057_,
		_w19058_,
		_w19080_
	);
	LUT2 #(
		.INIT('h8)
	) name8569 (
		_w19079_,
		_w19080_,
		_w19081_
	);
	LUT2 #(
		.INIT('h8)
	) name8570 (
		_w19077_,
		_w19078_,
		_w19082_
	);
	LUT2 #(
		.INIT('h8)
	) name8571 (
		_w19075_,
		_w19076_,
		_w19083_
	);
	LUT2 #(
		.INIT('h8)
	) name8572 (
		_w19073_,
		_w19074_,
		_w19084_
	);
	LUT2 #(
		.INIT('h8)
	) name8573 (
		_w19083_,
		_w19084_,
		_w19085_
	);
	LUT2 #(
		.INIT('h8)
	) name8574 (
		_w19081_,
		_w19082_,
		_w19086_
	);
	LUT2 #(
		.INIT('h8)
	) name8575 (
		_w19085_,
		_w19086_,
		_w19087_
	);
	LUT2 #(
		.INIT('h1)
	) name8576 (
		wb_rst_i_pad,
		_w19087_,
		_w19088_
	);
	LUT2 #(
		.INIT('h8)
	) name8577 (
		_w12656_,
		_w19088_,
		_w19089_
	);
	LUT2 #(
		.INIT('h8)
	) name8578 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		_w12658_,
		_w19090_
	);
	LUT2 #(
		.INIT('h1)
	) name8579 (
		_w18576_,
		_w19090_,
		_w19091_
	);
	LUT2 #(
		.INIT('h4)
	) name8580 (
		_w19089_,
		_w19091_,
		_w19092_
	);
	LUT2 #(
		.INIT('h8)
	) name8581 (
		\wishbone_bd_ram_mem3_reg[67][31]/P0001 ,
		_w13134_,
		_w19093_
	);
	LUT2 #(
		.INIT('h8)
	) name8582 (
		\wishbone_bd_ram_mem3_reg[38][31]/P0001 ,
		_w13182_,
		_w19094_
	);
	LUT2 #(
		.INIT('h8)
	) name8583 (
		\wishbone_bd_ram_mem3_reg[58][31]/P0001 ,
		_w13070_,
		_w19095_
	);
	LUT2 #(
		.INIT('h8)
	) name8584 (
		\wishbone_bd_ram_mem3_reg[143][31]/P0001 ,
		_w12922_,
		_w19096_
	);
	LUT2 #(
		.INIT('h8)
	) name8585 (
		\wishbone_bd_ram_mem3_reg[157][31]/P0001 ,
		_w12926_,
		_w19097_
	);
	LUT2 #(
		.INIT('h8)
	) name8586 (
		\wishbone_bd_ram_mem3_reg[244][31]/P0001 ,
		_w12747_,
		_w19098_
	);
	LUT2 #(
		.INIT('h8)
	) name8587 (
		\wishbone_bd_ram_mem3_reg[84][31]/P0001 ,
		_w12934_,
		_w19099_
	);
	LUT2 #(
		.INIT('h8)
	) name8588 (
		\wishbone_bd_ram_mem3_reg[109][31]/P0001 ,
		_w12888_,
		_w19100_
	);
	LUT2 #(
		.INIT('h8)
	) name8589 (
		\wishbone_bd_ram_mem3_reg[192][31]/P0001 ,
		_w12938_,
		_w19101_
	);
	LUT2 #(
		.INIT('h8)
	) name8590 (
		\wishbone_bd_ram_mem3_reg[190][31]/P0001 ,
		_w12858_,
		_w19102_
	);
	LUT2 #(
		.INIT('h8)
	) name8591 (
		\wishbone_bd_ram_mem3_reg[242][31]/P0001 ,
		_w12932_,
		_w19103_
	);
	LUT2 #(
		.INIT('h8)
	) name8592 (
		\wishbone_bd_ram_mem3_reg[87][31]/P0001 ,
		_w13154_,
		_w19104_
	);
	LUT2 #(
		.INIT('h8)
	) name8593 (
		\wishbone_bd_ram_mem3_reg[43][31]/P0001 ,
		_w13200_,
		_w19105_
	);
	LUT2 #(
		.INIT('h8)
	) name8594 (
		\wishbone_bd_ram_mem3_reg[133][31]/P0001 ,
		_w12761_,
		_w19106_
	);
	LUT2 #(
		.INIT('h8)
	) name8595 (
		\wishbone_bd_ram_mem3_reg[161][31]/P0001 ,
		_w12754_,
		_w19107_
	);
	LUT2 #(
		.INIT('h8)
	) name8596 (
		\wishbone_bd_ram_mem3_reg[48][31]/P0001 ,
		_w12970_,
		_w19108_
	);
	LUT2 #(
		.INIT('h8)
	) name8597 (
		\wishbone_bd_ram_mem3_reg[113][31]/P0001 ,
		_w13026_,
		_w19109_
	);
	LUT2 #(
		.INIT('h8)
	) name8598 (
		\wishbone_bd_ram_mem3_reg[94][31]/P0001 ,
		_w13186_,
		_w19110_
	);
	LUT2 #(
		.INIT('h8)
	) name8599 (
		\wishbone_bd_ram_mem3_reg[47][31]/P0001 ,
		_w12904_,
		_w19111_
	);
	LUT2 #(
		.INIT('h8)
	) name8600 (
		\wishbone_bd_ram_mem3_reg[37][31]/P0001 ,
		_w13102_,
		_w19112_
	);
	LUT2 #(
		.INIT('h8)
	) name8601 (
		\wishbone_bd_ram_mem3_reg[160][31]/P0001 ,
		_w12872_,
		_w19113_
	);
	LUT2 #(
		.INIT('h8)
	) name8602 (
		\wishbone_bd_ram_mem3_reg[234][31]/P0001 ,
		_w13214_,
		_w19114_
	);
	LUT2 #(
		.INIT('h8)
	) name8603 (
		\wishbone_bd_ram_mem3_reg[183][31]/P0001 ,
		_w12787_,
		_w19115_
	);
	LUT2 #(
		.INIT('h8)
	) name8604 (
		\wishbone_bd_ram_mem3_reg[182][31]/P0001 ,
		_w12820_,
		_w19116_
	);
	LUT2 #(
		.INIT('h8)
	) name8605 (
		\wishbone_bd_ram_mem3_reg[228][31]/P0001 ,
		_w12765_,
		_w19117_
	);
	LUT2 #(
		.INIT('h8)
	) name8606 (
		\wishbone_bd_ram_mem3_reg[118][31]/P0001 ,
		_w12830_,
		_w19118_
	);
	LUT2 #(
		.INIT('h8)
	) name8607 (
		\wishbone_bd_ram_mem3_reg[230][31]/P0001 ,
		_w13036_,
		_w19119_
	);
	LUT2 #(
		.INIT('h8)
	) name8608 (
		\wishbone_bd_ram_mem3_reg[202][31]/P0001 ,
		_w12870_,
		_w19120_
	);
	LUT2 #(
		.INIT('h8)
	) name8609 (
		\wishbone_bd_ram_mem3_reg[105][31]/P0001 ,
		_w12751_,
		_w19121_
	);
	LUT2 #(
		.INIT('h8)
	) name8610 (
		\wishbone_bd_ram_mem3_reg[45][31]/P0001 ,
		_w12908_,
		_w19122_
	);
	LUT2 #(
		.INIT('h8)
	) name8611 (
		\wishbone_bd_ram_mem3_reg[172][31]/P0001 ,
		_w12944_,
		_w19123_
	);
	LUT2 #(
		.INIT('h8)
	) name8612 (
		\wishbone_bd_ram_mem3_reg[200][31]/P0001 ,
		_w12988_,
		_w19124_
	);
	LUT2 #(
		.INIT('h8)
	) name8613 (
		\wishbone_bd_ram_mem3_reg[9][31]/P0001 ,
		_w12808_,
		_w19125_
	);
	LUT2 #(
		.INIT('h8)
	) name8614 (
		\wishbone_bd_ram_mem3_reg[217][31]/P0001 ,
		_w13188_,
		_w19126_
	);
	LUT2 #(
		.INIT('h8)
	) name8615 (
		\wishbone_bd_ram_mem3_reg[32][31]/P0001 ,
		_w13120_,
		_w19127_
	);
	LUT2 #(
		.INIT('h8)
	) name8616 (
		\wishbone_bd_ram_mem3_reg[53][31]/P0001 ,
		_w13020_,
		_w19128_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		\wishbone_bd_ram_mem3_reg[135][31]/P0001 ,
		_w13124_,
		_w19129_
	);
	LUT2 #(
		.INIT('h8)
	) name8618 (
		\wishbone_bd_ram_mem3_reg[136][31]/P0001 ,
		_w13064_,
		_w19130_
	);
	LUT2 #(
		.INIT('h8)
	) name8619 (
		\wishbone_bd_ram_mem3_reg[97][31]/P0001 ,
		_w13096_,
		_w19131_
	);
	LUT2 #(
		.INIT('h8)
	) name8620 (
		\wishbone_bd_ram_mem3_reg[70][31]/P0001 ,
		_w12840_,
		_w19132_
	);
	LUT2 #(
		.INIT('h8)
	) name8621 (
		\wishbone_bd_ram_mem3_reg[205][31]/P0001 ,
		_w13068_,
		_w19133_
	);
	LUT2 #(
		.INIT('h8)
	) name8622 (
		\wishbone_bd_ram_mem3_reg[215][31]/P0001 ,
		_w12974_,
		_w19134_
	);
	LUT2 #(
		.INIT('h8)
	) name8623 (
		\wishbone_bd_ram_mem3_reg[98][31]/P0001 ,
		_w12816_,
		_w19135_
	);
	LUT2 #(
		.INIT('h8)
	) name8624 (
		\wishbone_bd_ram_mem3_reg[49][31]/P0001 ,
		_w12994_,
		_w19136_
	);
	LUT2 #(
		.INIT('h8)
	) name8625 (
		\wishbone_bd_ram_mem3_reg[204][31]/P0001 ,
		_w13162_,
		_w19137_
	);
	LUT2 #(
		.INIT('h8)
	) name8626 (
		\wishbone_bd_ram_mem3_reg[81][31]/P0001 ,
		_w12950_,
		_w19138_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		\wishbone_bd_ram_mem3_reg[159][31]/P0001 ,
		_w12774_,
		_w19139_
	);
	LUT2 #(
		.INIT('h8)
	) name8628 (
		\wishbone_bd_ram_mem3_reg[233][31]/P0001 ,
		_w12836_,
		_w19140_
	);
	LUT2 #(
		.INIT('h8)
	) name8629 (
		\wishbone_bd_ram_mem3_reg[203][31]/P0001 ,
		_w13158_,
		_w19141_
	);
	LUT2 #(
		.INIT('h8)
	) name8630 (
		\wishbone_bd_ram_mem3_reg[252][31]/P0001 ,
		_w13080_,
		_w19142_
	);
	LUT2 #(
		.INIT('h8)
	) name8631 (
		\wishbone_bd_ram_mem3_reg[3][31]/P0001 ,
		_w12866_,
		_w19143_
	);
	LUT2 #(
		.INIT('h8)
	) name8632 (
		\wishbone_bd_ram_mem3_reg[149][31]/P0001 ,
		_w12741_,
		_w19144_
	);
	LUT2 #(
		.INIT('h8)
	) name8633 (
		\wishbone_bd_ram_mem3_reg[41][31]/P0001 ,
		_w13052_,
		_w19145_
	);
	LUT2 #(
		.INIT('h8)
	) name8634 (
		\wishbone_bd_ram_mem3_reg[241][31]/P0001 ,
		_w13006_,
		_w19146_
	);
	LUT2 #(
		.INIT('h8)
	) name8635 (
		\wishbone_bd_ram_mem3_reg[171][31]/P0001 ,
		_w12910_,
		_w19147_
	);
	LUT2 #(
		.INIT('h8)
	) name8636 (
		\wishbone_bd_ram_mem3_reg[197][31]/P0001 ,
		_w12834_,
		_w19148_
	);
	LUT2 #(
		.INIT('h8)
	) name8637 (
		\wishbone_bd_ram_mem3_reg[174][31]/P0001 ,
		_w12972_,
		_w19149_
	);
	LUT2 #(
		.INIT('h8)
	) name8638 (
		\wishbone_bd_ram_mem3_reg[248][31]/P0001 ,
		_w12789_,
		_w19150_
	);
	LUT2 #(
		.INIT('h8)
	) name8639 (
		\wishbone_bd_ram_mem3_reg[168][31]/P0001 ,
		_w13208_,
		_w19151_
	);
	LUT2 #(
		.INIT('h8)
	) name8640 (
		\wishbone_bd_ram_mem3_reg[150][31]/P0001 ,
		_w13136_,
		_w19152_
	);
	LUT2 #(
		.INIT('h8)
	) name8641 (
		\wishbone_bd_ram_mem3_reg[191][31]/P0001 ,
		_w13034_,
		_w19153_
	);
	LUT2 #(
		.INIT('h8)
	) name8642 (
		\wishbone_bd_ram_mem3_reg[29][31]/P0001 ,
		_w12952_,
		_w19154_
	);
	LUT2 #(
		.INIT('h8)
	) name8643 (
		\wishbone_bd_ram_mem3_reg[188][31]/P0001 ,
		_w12948_,
		_w19155_
	);
	LUT2 #(
		.INIT('h8)
	) name8644 (
		\wishbone_bd_ram_mem3_reg[127][31]/P0001 ,
		_w13164_,
		_w19156_
	);
	LUT2 #(
		.INIT('h8)
	) name8645 (
		\wishbone_bd_ram_mem3_reg[240][31]/P0001 ,
		_w12864_,
		_w19157_
	);
	LUT2 #(
		.INIT('h8)
	) name8646 (
		\wishbone_bd_ram_mem3_reg[185][31]/P0001 ,
		_w12940_,
		_w19158_
	);
	LUT2 #(
		.INIT('h8)
	) name8647 (
		\wishbone_bd_ram_mem3_reg[15][31]/P0001 ,
		_w13210_,
		_w19159_
	);
	LUT2 #(
		.INIT('h8)
	) name8648 (
		\wishbone_bd_ram_mem3_reg[17][31]/P0001 ,
		_w12848_,
		_w19160_
	);
	LUT2 #(
		.INIT('h8)
	) name8649 (
		\wishbone_bd_ram_mem3_reg[89][31]/P0001 ,
		_w12964_,
		_w19161_
	);
	LUT2 #(
		.INIT('h8)
	) name8650 (
		\wishbone_bd_ram_mem3_reg[186][31]/P0001 ,
		_w12783_,
		_w19162_
	);
	LUT2 #(
		.INIT('h8)
	) name8651 (
		\wishbone_bd_ram_mem3_reg[13][31]/P0001 ,
		_w13178_,
		_w19163_
	);
	LUT2 #(
		.INIT('h8)
	) name8652 (
		\wishbone_bd_ram_mem3_reg[93][31]/P0001 ,
		_w13016_,
		_w19164_
	);
	LUT2 #(
		.INIT('h8)
	) name8653 (
		\wishbone_bd_ram_mem3_reg[69][31]/P0001 ,
		_w12738_,
		_w19165_
	);
	LUT2 #(
		.INIT('h8)
	) name8654 (
		\wishbone_bd_ram_mem3_reg[179][31]/P0001 ,
		_w13050_,
		_w19166_
	);
	LUT2 #(
		.INIT('h8)
	) name8655 (
		\wishbone_bd_ram_mem3_reg[107][31]/P0001 ,
		_w12749_,
		_w19167_
	);
	LUT2 #(
		.INIT('h8)
	) name8656 (
		\wishbone_bd_ram_mem3_reg[254][31]/P0001 ,
		_w12892_,
		_w19168_
	);
	LUT2 #(
		.INIT('h8)
	) name8657 (
		\wishbone_bd_ram_mem3_reg[121][31]/P0001 ,
		_w13078_,
		_w19169_
	);
	LUT2 #(
		.INIT('h8)
	) name8658 (
		\wishbone_bd_ram_mem3_reg[187][31]/P0001 ,
		_w13196_,
		_w19170_
	);
	LUT2 #(
		.INIT('h8)
	) name8659 (
		\wishbone_bd_ram_mem3_reg[245][31]/P0001 ,
		_w13022_,
		_w19171_
	);
	LUT2 #(
		.INIT('h8)
	) name8660 (
		\wishbone_bd_ram_mem3_reg[72][31]/P0001 ,
		_w12810_,
		_w19172_
	);
	LUT2 #(
		.INIT('h8)
	) name8661 (
		\wishbone_bd_ram_mem3_reg[184][31]/P0001 ,
		_w13062_,
		_w19173_
	);
	LUT2 #(
		.INIT('h8)
	) name8662 (
		\wishbone_bd_ram_mem3_reg[139][31]/P0001 ,
		_w12814_,
		_w19174_
	);
	LUT2 #(
		.INIT('h8)
	) name8663 (
		\wishbone_bd_ram_mem3_reg[39][31]/P0001 ,
		_w13018_,
		_w19175_
	);
	LUT2 #(
		.INIT('h8)
	) name8664 (
		\wishbone_bd_ram_mem3_reg[220][31]/P0001 ,
		_w13066_,
		_w19176_
	);
	LUT2 #(
		.INIT('h8)
	) name8665 (
		\wishbone_bd_ram_mem3_reg[128][31]/P0001 ,
		_w12793_,
		_w19177_
	);
	LUT2 #(
		.INIT('h8)
	) name8666 (
		\wishbone_bd_ram_mem3_reg[68][31]/P0001 ,
		_w12946_,
		_w19178_
	);
	LUT2 #(
		.INIT('h8)
	) name8667 (
		\wishbone_bd_ram_mem3_reg[52][31]/P0001 ,
		_w13082_,
		_w19179_
	);
	LUT2 #(
		.INIT('h8)
	) name8668 (
		\wishbone_bd_ram_mem3_reg[7][31]/P0001 ,
		_w12728_,
		_w19180_
	);
	LUT2 #(
		.INIT('h8)
	) name8669 (
		\wishbone_bd_ram_mem3_reg[66][31]/P0001 ,
		_w12824_,
		_w19181_
	);
	LUT2 #(
		.INIT('h8)
	) name8670 (
		\wishbone_bd_ram_mem3_reg[227][31]/P0001 ,
		_w12936_,
		_w19182_
	);
	LUT2 #(
		.INIT('h8)
	) name8671 (
		\wishbone_bd_ram_mem3_reg[25][31]/P0001 ,
		_w13108_,
		_w19183_
	);
	LUT2 #(
		.INIT('h8)
	) name8672 (
		\wishbone_bd_ram_mem3_reg[180][31]/P0001 ,
		_w12791_,
		_w19184_
	);
	LUT2 #(
		.INIT('h8)
	) name8673 (
		\wishbone_bd_ram_mem3_reg[226][31]/P0001 ,
		_w13138_,
		_w19185_
	);
	LUT2 #(
		.INIT('h8)
	) name8674 (
		\wishbone_bd_ram_mem3_reg[247][31]/P0001 ,
		_w12818_,
		_w19186_
	);
	LUT2 #(
		.INIT('h8)
	) name8675 (
		\wishbone_bd_ram_mem3_reg[85][31]/P0001 ,
		_w13216_,
		_w19187_
	);
	LUT2 #(
		.INIT('h8)
	) name8676 (
		\wishbone_bd_ram_mem3_reg[193][31]/P0001 ,
		_w13056_,
		_w19188_
	);
	LUT2 #(
		.INIT('h8)
	) name8677 (
		\wishbone_bd_ram_mem3_reg[216][31]/P0001 ,
		_w13028_,
		_w19189_
	);
	LUT2 #(
		.INIT('h8)
	) name8678 (
		\wishbone_bd_ram_mem3_reg[170][31]/P0001 ,
		_w13030_,
		_w19190_
	);
	LUT2 #(
		.INIT('h8)
	) name8679 (
		\wishbone_bd_ram_mem3_reg[28][31]/P0001 ,
		_w13170_,
		_w19191_
	);
	LUT2 #(
		.INIT('h8)
	) name8680 (
		\wishbone_bd_ram_mem3_reg[42][31]/P0001 ,
		_w12842_,
		_w19192_
	);
	LUT2 #(
		.INIT('h8)
	) name8681 (
		\wishbone_bd_ram_mem3_reg[82][31]/P0001 ,
		_w12942_,
		_w19193_
	);
	LUT2 #(
		.INIT('h8)
	) name8682 (
		\wishbone_bd_ram_mem3_reg[103][31]/P0001 ,
		_w12846_,
		_w19194_
	);
	LUT2 #(
		.INIT('h8)
	) name8683 (
		\wishbone_bd_ram_mem3_reg[145][31]/P0001 ,
		_w13106_,
		_w19195_
	);
	LUT2 #(
		.INIT('h8)
	) name8684 (
		\wishbone_bd_ram_mem3_reg[104][31]/P0001 ,
		_w13148_,
		_w19196_
	);
	LUT2 #(
		.INIT('h8)
	) name8685 (
		\wishbone_bd_ram_mem3_reg[55][31]/P0001 ,
		_w12785_,
		_w19197_
	);
	LUT2 #(
		.INIT('h8)
	) name8686 (
		\wishbone_bd_ram_mem3_reg[51][31]/P0001 ,
		_w13024_,
		_w19198_
	);
	LUT2 #(
		.INIT('h8)
	) name8687 (
		\wishbone_bd_ram_mem3_reg[30][31]/P0001 ,
		_w13104_,
		_w19199_
	);
	LUT2 #(
		.INIT('h8)
	) name8688 (
		\wishbone_bd_ram_mem3_reg[144][31]/P0001 ,
		_w12756_,
		_w19200_
	);
	LUT2 #(
		.INIT('h8)
	) name8689 (
		\wishbone_bd_ram_mem3_reg[111][31]/P0001 ,
		_w12744_,
		_w19201_
	);
	LUT2 #(
		.INIT('h8)
	) name8690 (
		\wishbone_bd_ram_mem3_reg[60][31]/P0001 ,
		_w13204_,
		_w19202_
	);
	LUT2 #(
		.INIT('h8)
	) name8691 (
		\wishbone_bd_ram_mem3_reg[71][31]/P0001 ,
		_w12798_,
		_w19203_
	);
	LUT2 #(
		.INIT('h8)
	) name8692 (
		\wishbone_bd_ram_mem3_reg[119][31]/P0001 ,
		_w13048_,
		_w19204_
	);
	LUT2 #(
		.INIT('h8)
	) name8693 (
		\wishbone_bd_ram_mem3_reg[173][31]/P0001 ,
		_w12854_,
		_w19205_
	);
	LUT2 #(
		.INIT('h8)
	) name8694 (
		\wishbone_bd_ram_mem3_reg[57][31]/P0001 ,
		_w13116_,
		_w19206_
	);
	LUT2 #(
		.INIT('h8)
	) name8695 (
		\wishbone_bd_ram_mem3_reg[238][31]/P0001 ,
		_w13160_,
		_w19207_
	);
	LUT2 #(
		.INIT('h8)
	) name8696 (
		\wishbone_bd_ram_mem3_reg[189][31]/P0001 ,
		_w13042_,
		_w19208_
	);
	LUT2 #(
		.INIT('h8)
	) name8697 (
		\wishbone_bd_ram_mem3_reg[235][31]/P0001 ,
		_w12696_,
		_w19209_
	);
	LUT2 #(
		.INIT('h8)
	) name8698 (
		\wishbone_bd_ram_mem3_reg[218][31]/P0001 ,
		_w13206_,
		_w19210_
	);
	LUT2 #(
		.INIT('h8)
	) name8699 (
		\wishbone_bd_ram_mem3_reg[132][31]/P0001 ,
		_w12992_,
		_w19211_
	);
	LUT2 #(
		.INIT('h8)
	) name8700 (
		\wishbone_bd_ram_mem3_reg[0][31]/P0001 ,
		_w12717_,
		_w19212_
	);
	LUT2 #(
		.INIT('h8)
	) name8701 (
		\wishbone_bd_ram_mem3_reg[232][31]/P0001 ,
		_w12758_,
		_w19213_
	);
	LUT2 #(
		.INIT('h8)
	) name8702 (
		\wishbone_bd_ram_mem3_reg[221][31]/P0001 ,
		_w12802_,
		_w19214_
	);
	LUT2 #(
		.INIT('h8)
	) name8703 (
		\wishbone_bd_ram_mem3_reg[34][31]/P0001 ,
		_w12930_,
		_w19215_
	);
	LUT2 #(
		.INIT('h8)
	) name8704 (
		\wishbone_bd_ram_mem3_reg[239][31]/P0001 ,
		_w12862_,
		_w19216_
	);
	LUT2 #(
		.INIT('h8)
	) name8705 (
		\wishbone_bd_ram_mem3_reg[88][31]/P0001 ,
		_w12860_,
		_w19217_
	);
	LUT2 #(
		.INIT('h8)
	) name8706 (
		\wishbone_bd_ram_mem3_reg[14][31]/P0001 ,
		_w13086_,
		_w19218_
	);
	LUT2 #(
		.INIT('h8)
	) name8707 (
		\wishbone_bd_ram_mem3_reg[155][31]/P0001 ,
		_w13122_,
		_w19219_
	);
	LUT2 #(
		.INIT('h8)
	) name8708 (
		\wishbone_bd_ram_mem3_reg[210][31]/P0001 ,
		_w12924_,
		_w19220_
	);
	LUT2 #(
		.INIT('h8)
	) name8709 (
		\wishbone_bd_ram_mem3_reg[153][31]/P0001 ,
		_w12890_,
		_w19221_
	);
	LUT2 #(
		.INIT('h8)
	) name8710 (
		\wishbone_bd_ram_mem3_reg[134][31]/P0001 ,
		_w12763_,
		_w19222_
	);
	LUT2 #(
		.INIT('h8)
	) name8711 (
		\wishbone_bd_ram_mem3_reg[23][31]/P0001 ,
		_w13008_,
		_w19223_
	);
	LUT2 #(
		.INIT('h8)
	) name8712 (
		\wishbone_bd_ram_mem3_reg[11][31]/P0001 ,
		_w13194_,
		_w19224_
	);
	LUT2 #(
		.INIT('h8)
	) name8713 (
		\wishbone_bd_ram_mem3_reg[156][31]/P0001 ,
		_w13190_,
		_w19225_
	);
	LUT2 #(
		.INIT('h8)
	) name8714 (
		\wishbone_bd_ram_mem3_reg[36][31]/P0001 ,
		_w12800_,
		_w19226_
	);
	LUT2 #(
		.INIT('h8)
	) name8715 (
		\wishbone_bd_ram_mem3_reg[78][31]/P0001 ,
		_w12874_,
		_w19227_
	);
	LUT2 #(
		.INIT('h8)
	) name8716 (
		\wishbone_bd_ram_mem3_reg[231][31]/P0001 ,
		_w12856_,
		_w19228_
	);
	LUT2 #(
		.INIT('h8)
	) name8717 (
		\wishbone_bd_ram_mem3_reg[142][31]/P0001 ,
		_w12928_,
		_w19229_
	);
	LUT2 #(
		.INIT('h8)
	) name8718 (
		\wishbone_bd_ram_mem3_reg[20][31]/P0001 ,
		_w13174_,
		_w19230_
	);
	LUT2 #(
		.INIT('h8)
	) name8719 (
		\wishbone_bd_ram_mem3_reg[194][31]/P0001 ,
		_w12772_,
		_w19231_
	);
	LUT2 #(
		.INIT('h8)
	) name8720 (
		\wishbone_bd_ram_mem3_reg[63][31]/P0001 ,
		_w12850_,
		_w19232_
	);
	LUT2 #(
		.INIT('h8)
	) name8721 (
		\wishbone_bd_ram_mem3_reg[243][31]/P0001 ,
		_w12804_,
		_w19233_
	);
	LUT2 #(
		.INIT('h8)
	) name8722 (
		\wishbone_bd_ram_mem3_reg[158][31]/P0001 ,
		_w12898_,
		_w19234_
	);
	LUT2 #(
		.INIT('h8)
	) name8723 (
		\wishbone_bd_ram_mem3_reg[162][31]/P0001 ,
		_w13098_,
		_w19235_
	);
	LUT2 #(
		.INIT('h8)
	) name8724 (
		\wishbone_bd_ram_mem3_reg[26][31]/P0001 ,
		_w12699_,
		_w19236_
	);
	LUT2 #(
		.INIT('h8)
	) name8725 (
		\wishbone_bd_ram_mem3_reg[108][31]/P0001 ,
		_w13156_,
		_w19237_
	);
	LUT2 #(
		.INIT('h8)
	) name8726 (
		\wishbone_bd_ram_mem3_reg[137][31]/P0001 ,
		_w13168_,
		_w19238_
	);
	LUT2 #(
		.INIT('h8)
	) name8727 (
		\wishbone_bd_ram_mem3_reg[62][31]/P0001 ,
		_w12673_,
		_w19239_
	);
	LUT2 #(
		.INIT('h8)
	) name8728 (
		\wishbone_bd_ram_mem3_reg[206][31]/P0001 ,
		_w12954_,
		_w19240_
	);
	LUT2 #(
		.INIT('h8)
	) name8729 (
		\wishbone_bd_ram_mem3_reg[64][31]/P0001 ,
		_w12976_,
		_w19241_
	);
	LUT2 #(
		.INIT('h8)
	) name8730 (
		\wishbone_bd_ram_mem3_reg[196][31]/P0001 ,
		_w13090_,
		_w19242_
	);
	LUT2 #(
		.INIT('h8)
	) name8731 (
		\wishbone_bd_ram_mem3_reg[59][31]/P0001 ,
		_w12780_,
		_w19243_
	);
	LUT2 #(
		.INIT('h8)
	) name8732 (
		\wishbone_bd_ram_mem3_reg[123][31]/P0001 ,
		_w13114_,
		_w19244_
	);
	LUT2 #(
		.INIT('h8)
	) name8733 (
		\wishbone_bd_ram_mem3_reg[31][31]/P0001 ,
		_w13198_,
		_w19245_
	);
	LUT2 #(
		.INIT('h8)
	) name8734 (
		\wishbone_bd_ram_mem3_reg[16][31]/P0001 ,
		_w13140_,
		_w19246_
	);
	LUT2 #(
		.INIT('h8)
	) name8735 (
		\wishbone_bd_ram_mem3_reg[54][31]/P0001 ,
		_w12770_,
		_w19247_
	);
	LUT2 #(
		.INIT('h8)
	) name8736 (
		\wishbone_bd_ram_mem3_reg[86][31]/P0001 ,
		_w12735_,
		_w19248_
	);
	LUT2 #(
		.INIT('h8)
	) name8737 (
		\wishbone_bd_ram_mem3_reg[117][31]/P0001 ,
		_w12715_,
		_w19249_
	);
	LUT2 #(
		.INIT('h8)
	) name8738 (
		\wishbone_bd_ram_mem3_reg[181][31]/P0001 ,
		_w12828_,
		_w19250_
	);
	LUT2 #(
		.INIT('h8)
	) name8739 (
		\wishbone_bd_ram_mem3_reg[46][31]/P0001 ,
		_w12884_,
		_w19251_
	);
	LUT2 #(
		.INIT('h8)
	) name8740 (
		\wishbone_bd_ram_mem3_reg[201][31]/P0001 ,
		_w12822_,
		_w19252_
	);
	LUT2 #(
		.INIT('h8)
	) name8741 (
		\wishbone_bd_ram_mem3_reg[225][31]/P0001 ,
		_w13092_,
		_w19253_
	);
	LUT2 #(
		.INIT('h8)
	) name8742 (
		\wishbone_bd_ram_mem3_reg[255][31]/P0001 ,
		_w13072_,
		_w19254_
	);
	LUT2 #(
		.INIT('h8)
	) name8743 (
		\wishbone_bd_ram_mem3_reg[122][31]/P0001 ,
		_w13130_,
		_w19255_
	);
	LUT2 #(
		.INIT('h8)
	) name8744 (
		\wishbone_bd_ram_mem3_reg[126][31]/P0001 ,
		_w13218_,
		_w19256_
	);
	LUT2 #(
		.INIT('h8)
	) name8745 (
		\wishbone_bd_ram_mem3_reg[151][31]/P0001 ,
		_w13142_,
		_w19257_
	);
	LUT2 #(
		.INIT('h8)
	) name8746 (
		\wishbone_bd_ram_mem3_reg[208][31]/P0001 ,
		_w13032_,
		_w19258_
	);
	LUT2 #(
		.INIT('h8)
	) name8747 (
		\wishbone_bd_ram_mem3_reg[130][31]/P0001 ,
		_w12914_,
		_w19259_
	);
	LUT2 #(
		.INIT('h8)
	) name8748 (
		\wishbone_bd_ram_mem3_reg[102][31]/P0001 ,
		_w12685_,
		_w19260_
	);
	LUT2 #(
		.INIT('h8)
	) name8749 (
		\wishbone_bd_ram_mem3_reg[129][31]/P0001 ,
		_w12776_,
		_w19261_
	);
	LUT2 #(
		.INIT('h8)
	) name8750 (
		\wishbone_bd_ram_mem3_reg[146][31]/P0001 ,
		_w13060_,
		_w19262_
	);
	LUT2 #(
		.INIT('h8)
	) name8751 (
		\wishbone_bd_ram_mem3_reg[8][31]/P0001 ,
		_w12920_,
		_w19263_
	);
	LUT2 #(
		.INIT('h8)
	) name8752 (
		\wishbone_bd_ram_mem3_reg[209][31]/P0001 ,
		_w13152_,
		_w19264_
	);
	LUT2 #(
		.INIT('h8)
	) name8753 (
		\wishbone_bd_ram_mem3_reg[141][31]/P0001 ,
		_w13004_,
		_w19265_
	);
	LUT2 #(
		.INIT('h8)
	) name8754 (
		\wishbone_bd_ram_mem3_reg[250][31]/P0001 ,
		_w13128_,
		_w19266_
	);
	LUT2 #(
		.INIT('h8)
	) name8755 (
		\wishbone_bd_ram_mem3_reg[176][31]/P0001 ,
		_w12868_,
		_w19267_
	);
	LUT2 #(
		.INIT('h8)
	) name8756 (
		\wishbone_bd_ram_mem3_reg[198][31]/P0001 ,
		_w12832_,
		_w19268_
	);
	LUT2 #(
		.INIT('h8)
	) name8757 (
		\wishbone_bd_ram_mem3_reg[95][31]/P0001 ,
		_w12844_,
		_w19269_
	);
	LUT2 #(
		.INIT('h8)
	) name8758 (
		\wishbone_bd_ram_mem3_reg[195][31]/P0001 ,
		_w13144_,
		_w19270_
	);
	LUT2 #(
		.INIT('h8)
	) name8759 (
		\wishbone_bd_ram_mem3_reg[99][31]/P0001 ,
		_w13038_,
		_w19271_
	);
	LUT2 #(
		.INIT('h8)
	) name8760 (
		\wishbone_bd_ram_mem3_reg[211][31]/P0001 ,
		_w13166_,
		_w19272_
	);
	LUT2 #(
		.INIT('h8)
	) name8761 (
		\wishbone_bd_ram_mem3_reg[212][31]/P0001 ,
		_w12796_,
		_w19273_
	);
	LUT2 #(
		.INIT('h8)
	) name8762 (
		\wishbone_bd_ram_mem3_reg[5][31]/P0001 ,
		_w12878_,
		_w19274_
	);
	LUT2 #(
		.INIT('h8)
	) name8763 (
		\wishbone_bd_ram_mem3_reg[106][31]/P0001 ,
		_w12713_,
		_w19275_
	);
	LUT2 #(
		.INIT('h8)
	) name8764 (
		\wishbone_bd_ram_mem3_reg[154][31]/P0001 ,
		_w12962_,
		_w19276_
	);
	LUT2 #(
		.INIT('h8)
	) name8765 (
		\wishbone_bd_ram_mem3_reg[213][31]/P0001 ,
		_w13002_,
		_w19277_
	);
	LUT2 #(
		.INIT('h8)
	) name8766 (
		\wishbone_bd_ram_mem3_reg[96][31]/P0001 ,
		_w12912_,
		_w19278_
	);
	LUT2 #(
		.INIT('h8)
	) name8767 (
		\wishbone_bd_ram_mem3_reg[214][31]/P0001 ,
		_w12984_,
		_w19279_
	);
	LUT2 #(
		.INIT('h8)
	) name8768 (
		\wishbone_bd_ram_mem3_reg[4][31]/P0001 ,
		_w12666_,
		_w19280_
	);
	LUT2 #(
		.INIT('h8)
	) name8769 (
		\wishbone_bd_ram_mem3_reg[65][31]/P0001 ,
		_w13176_,
		_w19281_
	);
	LUT2 #(
		.INIT('h8)
	) name8770 (
		\wishbone_bd_ram_mem3_reg[115][31]/P0001 ,
		_w13112_,
		_w19282_
	);
	LUT2 #(
		.INIT('h8)
	) name8771 (
		\wishbone_bd_ram_mem3_reg[79][31]/P0001 ,
		_w13212_,
		_w19283_
	);
	LUT2 #(
		.INIT('h8)
	) name8772 (
		\wishbone_bd_ram_mem3_reg[124][31]/P0001 ,
		_w13058_,
		_w19284_
	);
	LUT2 #(
		.INIT('h8)
	) name8773 (
		\wishbone_bd_ram_mem3_reg[219][31]/P0001 ,
		_w12806_,
		_w19285_
	);
	LUT2 #(
		.INIT('h8)
	) name8774 (
		\wishbone_bd_ram_mem3_reg[169][31]/P0001 ,
		_w12722_,
		_w19286_
	);
	LUT2 #(
		.INIT('h8)
	) name8775 (
		\wishbone_bd_ram_mem3_reg[91][31]/P0001 ,
		_w13074_,
		_w19287_
	);
	LUT2 #(
		.INIT('h8)
	) name8776 (
		\wishbone_bd_ram_mem3_reg[222][31]/P0001 ,
		_w13094_,
		_w19288_
	);
	LUT2 #(
		.INIT('h8)
	) name8777 (
		\wishbone_bd_ram_mem3_reg[229][31]/P0001 ,
		_w12711_,
		_w19289_
	);
	LUT2 #(
		.INIT('h8)
	) name8778 (
		\wishbone_bd_ram_mem3_reg[12][31]/P0001 ,
		_w13118_,
		_w19290_
	);
	LUT2 #(
		.INIT('h8)
	) name8779 (
		\wishbone_bd_ram_mem3_reg[21][31]/P0001 ,
		_w12906_,
		_w19291_
	);
	LUT2 #(
		.INIT('h8)
	) name8780 (
		\wishbone_bd_ram_mem3_reg[166][31]/P0001 ,
		_w13040_,
		_w19292_
	);
	LUT2 #(
		.INIT('h8)
	) name8781 (
		\wishbone_bd_ram_mem3_reg[22][31]/P0001 ,
		_w13110_,
		_w19293_
	);
	LUT2 #(
		.INIT('h8)
	) name8782 (
		\wishbone_bd_ram_mem3_reg[6][31]/P0001 ,
		_w12968_,
		_w19294_
	);
	LUT2 #(
		.INIT('h8)
	) name8783 (
		\wishbone_bd_ram_mem3_reg[35][31]/P0001 ,
		_w12703_,
		_w19295_
	);
	LUT2 #(
		.INIT('h8)
	) name8784 (
		\wishbone_bd_ram_mem3_reg[165][31]/P0001 ,
		_w13044_,
		_w19296_
	);
	LUT2 #(
		.INIT('h8)
	) name8785 (
		\wishbone_bd_ram_mem3_reg[77][31]/P0001 ,
		_w12982_,
		_w19297_
	);
	LUT2 #(
		.INIT('h8)
	) name8786 (
		\wishbone_bd_ram_mem3_reg[24][31]/P0001 ,
		_w13084_,
		_w19298_
	);
	LUT2 #(
		.INIT('h8)
	) name8787 (
		\wishbone_bd_ram_mem3_reg[74][31]/P0001 ,
		_w12812_,
		_w19299_
	);
	LUT2 #(
		.INIT('h8)
	) name8788 (
		\wishbone_bd_ram_mem3_reg[76][31]/P0001 ,
		_w13184_,
		_w19300_
	);
	LUT2 #(
		.INIT('h8)
	) name8789 (
		\wishbone_bd_ram_mem3_reg[61][31]/P0001 ,
		_w12725_,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name8790 (
		\wishbone_bd_ram_mem3_reg[27][31]/P0001 ,
		_w12880_,
		_w19302_
	);
	LUT2 #(
		.INIT('h8)
	) name8791 (
		\wishbone_bd_ram_mem3_reg[207][31]/P0001 ,
		_w13180_,
		_w19303_
	);
	LUT2 #(
		.INIT('h8)
	) name8792 (
		\wishbone_bd_ram_mem3_reg[116][31]/P0001 ,
		_w12998_,
		_w19304_
	);
	LUT2 #(
		.INIT('h8)
	) name8793 (
		\wishbone_bd_ram_mem3_reg[44][31]/P0001 ,
		_w12896_,
		_w19305_
	);
	LUT2 #(
		.INIT('h8)
	) name8794 (
		\wishbone_bd_ram_mem3_reg[33][31]/P0001 ,
		_w12980_,
		_w19306_
	);
	LUT2 #(
		.INIT('h8)
	) name8795 (
		\wishbone_bd_ram_mem3_reg[167][31]/P0001 ,
		_w12986_,
		_w19307_
	);
	LUT2 #(
		.INIT('h8)
	) name8796 (
		\wishbone_bd_ram_mem3_reg[178][31]/P0001 ,
		_w12886_,
		_w19308_
	);
	LUT2 #(
		.INIT('h8)
	) name8797 (
		\wishbone_bd_ram_mem3_reg[56][31]/P0001 ,
		_w12778_,
		_w19309_
	);
	LUT2 #(
		.INIT('h8)
	) name8798 (
		\wishbone_bd_ram_mem3_reg[120][31]/P0001 ,
		_w12707_,
		_w19310_
	);
	LUT2 #(
		.INIT('h8)
	) name8799 (
		\wishbone_bd_ram_mem3_reg[112][31]/P0001 ,
		_w12733_,
		_w19311_
	);
	LUT2 #(
		.INIT('h8)
	) name8800 (
		\wishbone_bd_ram_mem3_reg[19][31]/P0001 ,
		_w13012_,
		_w19312_
	);
	LUT2 #(
		.INIT('h8)
	) name8801 (
		\wishbone_bd_ram_mem3_reg[125][31]/P0001 ,
		_w12956_,
		_w19313_
	);
	LUT2 #(
		.INIT('h8)
	) name8802 (
		\wishbone_bd_ram_mem3_reg[40][31]/P0001 ,
		_w13132_,
		_w19314_
	);
	LUT2 #(
		.INIT('h8)
	) name8803 (
		\wishbone_bd_ram_mem3_reg[224][31]/P0001 ,
		_w12902_,
		_w19315_
	);
	LUT2 #(
		.INIT('h8)
	) name8804 (
		\wishbone_bd_ram_mem3_reg[101][31]/P0001 ,
		_w13192_,
		_w19316_
	);
	LUT2 #(
		.INIT('h8)
	) name8805 (
		\wishbone_bd_ram_mem3_reg[90][31]/P0001 ,
		_w12978_,
		_w19317_
	);
	LUT2 #(
		.INIT('h8)
	) name8806 (
		\wishbone_bd_ram_mem3_reg[140][31]/P0001 ,
		_w12894_,
		_w19318_
	);
	LUT2 #(
		.INIT('h8)
	) name8807 (
		\wishbone_bd_ram_mem3_reg[253][31]/P0001 ,
		_w13100_,
		_w19319_
	);
	LUT2 #(
		.INIT('h8)
	) name8808 (
		\wishbone_bd_ram_mem3_reg[223][31]/P0001 ,
		_w12838_,
		_w19320_
	);
	LUT2 #(
		.INIT('h8)
	) name8809 (
		\wishbone_bd_ram_mem3_reg[199][31]/P0001 ,
		_w12768_,
		_w19321_
	);
	LUT2 #(
		.INIT('h8)
	) name8810 (
		\wishbone_bd_ram_mem3_reg[114][31]/P0001 ,
		_w13202_,
		_w19322_
	);
	LUT2 #(
		.INIT('h8)
	) name8811 (
		\wishbone_bd_ram_mem3_reg[138][31]/P0001 ,
		_w12958_,
		_w19323_
	);
	LUT2 #(
		.INIT('h8)
	) name8812 (
		\wishbone_bd_ram_mem3_reg[10][31]/P0001 ,
		_w13172_,
		_w19324_
	);
	LUT2 #(
		.INIT('h8)
	) name8813 (
		\wishbone_bd_ram_mem3_reg[75][31]/P0001 ,
		_w12826_,
		_w19325_
	);
	LUT2 #(
		.INIT('h8)
	) name8814 (
		\wishbone_bd_ram_mem3_reg[164][31]/P0001 ,
		_w12876_,
		_w19326_
	);
	LUT2 #(
		.INIT('h8)
	) name8815 (
		\wishbone_bd_ram_mem3_reg[50][31]/P0001 ,
		_w13150_,
		_w19327_
	);
	LUT2 #(
		.INIT('h8)
	) name8816 (
		\wishbone_bd_ram_mem3_reg[1][31]/P0001 ,
		_w13014_,
		_w19328_
	);
	LUT2 #(
		.INIT('h8)
	) name8817 (
		\wishbone_bd_ram_mem3_reg[246][31]/P0001 ,
		_w13076_,
		_w19329_
	);
	LUT2 #(
		.INIT('h8)
	) name8818 (
		\wishbone_bd_ram_mem3_reg[80][31]/P0001 ,
		_w12689_,
		_w19330_
	);
	LUT2 #(
		.INIT('h8)
	) name8819 (
		\wishbone_bd_ram_mem3_reg[147][31]/P0001 ,
		_w13146_,
		_w19331_
	);
	LUT2 #(
		.INIT('h8)
	) name8820 (
		\wishbone_bd_ram_mem3_reg[237][31]/P0001 ,
		_w12990_,
		_w19332_
	);
	LUT2 #(
		.INIT('h8)
	) name8821 (
		\wishbone_bd_ram_mem3_reg[249][31]/P0001 ,
		_w12900_,
		_w19333_
	);
	LUT2 #(
		.INIT('h8)
	) name8822 (
		\wishbone_bd_ram_mem3_reg[177][31]/P0001 ,
		_w12996_,
		_w19334_
	);
	LUT2 #(
		.INIT('h8)
	) name8823 (
		\wishbone_bd_ram_mem3_reg[92][31]/P0001 ,
		_w13010_,
		_w19335_
	);
	LUT2 #(
		.INIT('h8)
	) name8824 (
		\wishbone_bd_ram_mem3_reg[83][31]/P0001 ,
		_w12916_,
		_w19336_
	);
	LUT2 #(
		.INIT('h8)
	) name8825 (
		\wishbone_bd_ram_mem3_reg[251][31]/P0001 ,
		_w13054_,
		_w19337_
	);
	LUT2 #(
		.INIT('h8)
	) name8826 (
		\wishbone_bd_ram_mem3_reg[73][31]/P0001 ,
		_w12918_,
		_w19338_
	);
	LUT2 #(
		.INIT('h8)
	) name8827 (
		\wishbone_bd_ram_mem3_reg[2][31]/P0001 ,
		_w13088_,
		_w19339_
	);
	LUT2 #(
		.INIT('h8)
	) name8828 (
		\wishbone_bd_ram_mem3_reg[236][31]/P0001 ,
		_w12731_,
		_w19340_
	);
	LUT2 #(
		.INIT('h8)
	) name8829 (
		\wishbone_bd_ram_mem3_reg[131][31]/P0001 ,
		_w12852_,
		_w19341_
	);
	LUT2 #(
		.INIT('h8)
	) name8830 (
		\wishbone_bd_ram_mem3_reg[100][31]/P0001 ,
		_w12960_,
		_w19342_
	);
	LUT2 #(
		.INIT('h8)
	) name8831 (
		\wishbone_bd_ram_mem3_reg[152][31]/P0001 ,
		_w12966_,
		_w19343_
	);
	LUT2 #(
		.INIT('h8)
	) name8832 (
		\wishbone_bd_ram_mem3_reg[163][31]/P0001 ,
		_w12882_,
		_w19344_
	);
	LUT2 #(
		.INIT('h8)
	) name8833 (
		\wishbone_bd_ram_mem3_reg[18][31]/P0001 ,
		_w12679_,
		_w19345_
	);
	LUT2 #(
		.INIT('h8)
	) name8834 (
		\wishbone_bd_ram_mem3_reg[110][31]/P0001 ,
		_w13046_,
		_w19346_
	);
	LUT2 #(
		.INIT('h8)
	) name8835 (
		\wishbone_bd_ram_mem3_reg[148][31]/P0001 ,
		_w13000_,
		_w19347_
	);
	LUT2 #(
		.INIT('h8)
	) name8836 (
		\wishbone_bd_ram_mem3_reg[175][31]/P0001 ,
		_w13126_,
		_w19348_
	);
	LUT2 #(
		.INIT('h1)
	) name8837 (
		_w19093_,
		_w19094_,
		_w19349_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		_w19095_,
		_w19096_,
		_w19350_
	);
	LUT2 #(
		.INIT('h1)
	) name8839 (
		_w19097_,
		_w19098_,
		_w19351_
	);
	LUT2 #(
		.INIT('h1)
	) name8840 (
		_w19099_,
		_w19100_,
		_w19352_
	);
	LUT2 #(
		.INIT('h1)
	) name8841 (
		_w19101_,
		_w19102_,
		_w19353_
	);
	LUT2 #(
		.INIT('h1)
	) name8842 (
		_w19103_,
		_w19104_,
		_w19354_
	);
	LUT2 #(
		.INIT('h1)
	) name8843 (
		_w19105_,
		_w19106_,
		_w19355_
	);
	LUT2 #(
		.INIT('h1)
	) name8844 (
		_w19107_,
		_w19108_,
		_w19356_
	);
	LUT2 #(
		.INIT('h1)
	) name8845 (
		_w19109_,
		_w19110_,
		_w19357_
	);
	LUT2 #(
		.INIT('h1)
	) name8846 (
		_w19111_,
		_w19112_,
		_w19358_
	);
	LUT2 #(
		.INIT('h1)
	) name8847 (
		_w19113_,
		_w19114_,
		_w19359_
	);
	LUT2 #(
		.INIT('h1)
	) name8848 (
		_w19115_,
		_w19116_,
		_w19360_
	);
	LUT2 #(
		.INIT('h1)
	) name8849 (
		_w19117_,
		_w19118_,
		_w19361_
	);
	LUT2 #(
		.INIT('h1)
	) name8850 (
		_w19119_,
		_w19120_,
		_w19362_
	);
	LUT2 #(
		.INIT('h1)
	) name8851 (
		_w19121_,
		_w19122_,
		_w19363_
	);
	LUT2 #(
		.INIT('h1)
	) name8852 (
		_w19123_,
		_w19124_,
		_w19364_
	);
	LUT2 #(
		.INIT('h1)
	) name8853 (
		_w19125_,
		_w19126_,
		_w19365_
	);
	LUT2 #(
		.INIT('h1)
	) name8854 (
		_w19127_,
		_w19128_,
		_w19366_
	);
	LUT2 #(
		.INIT('h1)
	) name8855 (
		_w19129_,
		_w19130_,
		_w19367_
	);
	LUT2 #(
		.INIT('h1)
	) name8856 (
		_w19131_,
		_w19132_,
		_w19368_
	);
	LUT2 #(
		.INIT('h1)
	) name8857 (
		_w19133_,
		_w19134_,
		_w19369_
	);
	LUT2 #(
		.INIT('h1)
	) name8858 (
		_w19135_,
		_w19136_,
		_w19370_
	);
	LUT2 #(
		.INIT('h1)
	) name8859 (
		_w19137_,
		_w19138_,
		_w19371_
	);
	LUT2 #(
		.INIT('h1)
	) name8860 (
		_w19139_,
		_w19140_,
		_w19372_
	);
	LUT2 #(
		.INIT('h1)
	) name8861 (
		_w19141_,
		_w19142_,
		_w19373_
	);
	LUT2 #(
		.INIT('h1)
	) name8862 (
		_w19143_,
		_w19144_,
		_w19374_
	);
	LUT2 #(
		.INIT('h1)
	) name8863 (
		_w19145_,
		_w19146_,
		_w19375_
	);
	LUT2 #(
		.INIT('h1)
	) name8864 (
		_w19147_,
		_w19148_,
		_w19376_
	);
	LUT2 #(
		.INIT('h1)
	) name8865 (
		_w19149_,
		_w19150_,
		_w19377_
	);
	LUT2 #(
		.INIT('h1)
	) name8866 (
		_w19151_,
		_w19152_,
		_w19378_
	);
	LUT2 #(
		.INIT('h1)
	) name8867 (
		_w19153_,
		_w19154_,
		_w19379_
	);
	LUT2 #(
		.INIT('h1)
	) name8868 (
		_w19155_,
		_w19156_,
		_w19380_
	);
	LUT2 #(
		.INIT('h1)
	) name8869 (
		_w19157_,
		_w19158_,
		_w19381_
	);
	LUT2 #(
		.INIT('h1)
	) name8870 (
		_w19159_,
		_w19160_,
		_w19382_
	);
	LUT2 #(
		.INIT('h1)
	) name8871 (
		_w19161_,
		_w19162_,
		_w19383_
	);
	LUT2 #(
		.INIT('h1)
	) name8872 (
		_w19163_,
		_w19164_,
		_w19384_
	);
	LUT2 #(
		.INIT('h1)
	) name8873 (
		_w19165_,
		_w19166_,
		_w19385_
	);
	LUT2 #(
		.INIT('h1)
	) name8874 (
		_w19167_,
		_w19168_,
		_w19386_
	);
	LUT2 #(
		.INIT('h1)
	) name8875 (
		_w19169_,
		_w19170_,
		_w19387_
	);
	LUT2 #(
		.INIT('h1)
	) name8876 (
		_w19171_,
		_w19172_,
		_w19388_
	);
	LUT2 #(
		.INIT('h1)
	) name8877 (
		_w19173_,
		_w19174_,
		_w19389_
	);
	LUT2 #(
		.INIT('h1)
	) name8878 (
		_w19175_,
		_w19176_,
		_w19390_
	);
	LUT2 #(
		.INIT('h1)
	) name8879 (
		_w19177_,
		_w19178_,
		_w19391_
	);
	LUT2 #(
		.INIT('h1)
	) name8880 (
		_w19179_,
		_w19180_,
		_w19392_
	);
	LUT2 #(
		.INIT('h1)
	) name8881 (
		_w19181_,
		_w19182_,
		_w19393_
	);
	LUT2 #(
		.INIT('h1)
	) name8882 (
		_w19183_,
		_w19184_,
		_w19394_
	);
	LUT2 #(
		.INIT('h1)
	) name8883 (
		_w19185_,
		_w19186_,
		_w19395_
	);
	LUT2 #(
		.INIT('h1)
	) name8884 (
		_w19187_,
		_w19188_,
		_w19396_
	);
	LUT2 #(
		.INIT('h1)
	) name8885 (
		_w19189_,
		_w19190_,
		_w19397_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w19191_,
		_w19192_,
		_w19398_
	);
	LUT2 #(
		.INIT('h1)
	) name8887 (
		_w19193_,
		_w19194_,
		_w19399_
	);
	LUT2 #(
		.INIT('h1)
	) name8888 (
		_w19195_,
		_w19196_,
		_w19400_
	);
	LUT2 #(
		.INIT('h1)
	) name8889 (
		_w19197_,
		_w19198_,
		_w19401_
	);
	LUT2 #(
		.INIT('h1)
	) name8890 (
		_w19199_,
		_w19200_,
		_w19402_
	);
	LUT2 #(
		.INIT('h1)
	) name8891 (
		_w19201_,
		_w19202_,
		_w19403_
	);
	LUT2 #(
		.INIT('h1)
	) name8892 (
		_w19203_,
		_w19204_,
		_w19404_
	);
	LUT2 #(
		.INIT('h1)
	) name8893 (
		_w19205_,
		_w19206_,
		_w19405_
	);
	LUT2 #(
		.INIT('h1)
	) name8894 (
		_w19207_,
		_w19208_,
		_w19406_
	);
	LUT2 #(
		.INIT('h1)
	) name8895 (
		_w19209_,
		_w19210_,
		_w19407_
	);
	LUT2 #(
		.INIT('h1)
	) name8896 (
		_w19211_,
		_w19212_,
		_w19408_
	);
	LUT2 #(
		.INIT('h1)
	) name8897 (
		_w19213_,
		_w19214_,
		_w19409_
	);
	LUT2 #(
		.INIT('h1)
	) name8898 (
		_w19215_,
		_w19216_,
		_w19410_
	);
	LUT2 #(
		.INIT('h1)
	) name8899 (
		_w19217_,
		_w19218_,
		_w19411_
	);
	LUT2 #(
		.INIT('h1)
	) name8900 (
		_w19219_,
		_w19220_,
		_w19412_
	);
	LUT2 #(
		.INIT('h1)
	) name8901 (
		_w19221_,
		_w19222_,
		_w19413_
	);
	LUT2 #(
		.INIT('h1)
	) name8902 (
		_w19223_,
		_w19224_,
		_w19414_
	);
	LUT2 #(
		.INIT('h1)
	) name8903 (
		_w19225_,
		_w19226_,
		_w19415_
	);
	LUT2 #(
		.INIT('h1)
	) name8904 (
		_w19227_,
		_w19228_,
		_w19416_
	);
	LUT2 #(
		.INIT('h1)
	) name8905 (
		_w19229_,
		_w19230_,
		_w19417_
	);
	LUT2 #(
		.INIT('h1)
	) name8906 (
		_w19231_,
		_w19232_,
		_w19418_
	);
	LUT2 #(
		.INIT('h1)
	) name8907 (
		_w19233_,
		_w19234_,
		_w19419_
	);
	LUT2 #(
		.INIT('h1)
	) name8908 (
		_w19235_,
		_w19236_,
		_w19420_
	);
	LUT2 #(
		.INIT('h1)
	) name8909 (
		_w19237_,
		_w19238_,
		_w19421_
	);
	LUT2 #(
		.INIT('h1)
	) name8910 (
		_w19239_,
		_w19240_,
		_w19422_
	);
	LUT2 #(
		.INIT('h1)
	) name8911 (
		_w19241_,
		_w19242_,
		_w19423_
	);
	LUT2 #(
		.INIT('h1)
	) name8912 (
		_w19243_,
		_w19244_,
		_w19424_
	);
	LUT2 #(
		.INIT('h1)
	) name8913 (
		_w19245_,
		_w19246_,
		_w19425_
	);
	LUT2 #(
		.INIT('h1)
	) name8914 (
		_w19247_,
		_w19248_,
		_w19426_
	);
	LUT2 #(
		.INIT('h1)
	) name8915 (
		_w19249_,
		_w19250_,
		_w19427_
	);
	LUT2 #(
		.INIT('h1)
	) name8916 (
		_w19251_,
		_w19252_,
		_w19428_
	);
	LUT2 #(
		.INIT('h1)
	) name8917 (
		_w19253_,
		_w19254_,
		_w19429_
	);
	LUT2 #(
		.INIT('h1)
	) name8918 (
		_w19255_,
		_w19256_,
		_w19430_
	);
	LUT2 #(
		.INIT('h1)
	) name8919 (
		_w19257_,
		_w19258_,
		_w19431_
	);
	LUT2 #(
		.INIT('h1)
	) name8920 (
		_w19259_,
		_w19260_,
		_w19432_
	);
	LUT2 #(
		.INIT('h1)
	) name8921 (
		_w19261_,
		_w19262_,
		_w19433_
	);
	LUT2 #(
		.INIT('h1)
	) name8922 (
		_w19263_,
		_w19264_,
		_w19434_
	);
	LUT2 #(
		.INIT('h1)
	) name8923 (
		_w19265_,
		_w19266_,
		_w19435_
	);
	LUT2 #(
		.INIT('h1)
	) name8924 (
		_w19267_,
		_w19268_,
		_w19436_
	);
	LUT2 #(
		.INIT('h1)
	) name8925 (
		_w19269_,
		_w19270_,
		_w19437_
	);
	LUT2 #(
		.INIT('h1)
	) name8926 (
		_w19271_,
		_w19272_,
		_w19438_
	);
	LUT2 #(
		.INIT('h1)
	) name8927 (
		_w19273_,
		_w19274_,
		_w19439_
	);
	LUT2 #(
		.INIT('h1)
	) name8928 (
		_w19275_,
		_w19276_,
		_w19440_
	);
	LUT2 #(
		.INIT('h1)
	) name8929 (
		_w19277_,
		_w19278_,
		_w19441_
	);
	LUT2 #(
		.INIT('h1)
	) name8930 (
		_w19279_,
		_w19280_,
		_w19442_
	);
	LUT2 #(
		.INIT('h1)
	) name8931 (
		_w19281_,
		_w19282_,
		_w19443_
	);
	LUT2 #(
		.INIT('h1)
	) name8932 (
		_w19283_,
		_w19284_,
		_w19444_
	);
	LUT2 #(
		.INIT('h1)
	) name8933 (
		_w19285_,
		_w19286_,
		_w19445_
	);
	LUT2 #(
		.INIT('h1)
	) name8934 (
		_w19287_,
		_w19288_,
		_w19446_
	);
	LUT2 #(
		.INIT('h1)
	) name8935 (
		_w19289_,
		_w19290_,
		_w19447_
	);
	LUT2 #(
		.INIT('h1)
	) name8936 (
		_w19291_,
		_w19292_,
		_w19448_
	);
	LUT2 #(
		.INIT('h1)
	) name8937 (
		_w19293_,
		_w19294_,
		_w19449_
	);
	LUT2 #(
		.INIT('h1)
	) name8938 (
		_w19295_,
		_w19296_,
		_w19450_
	);
	LUT2 #(
		.INIT('h1)
	) name8939 (
		_w19297_,
		_w19298_,
		_w19451_
	);
	LUT2 #(
		.INIT('h1)
	) name8940 (
		_w19299_,
		_w19300_,
		_w19452_
	);
	LUT2 #(
		.INIT('h1)
	) name8941 (
		_w19301_,
		_w19302_,
		_w19453_
	);
	LUT2 #(
		.INIT('h1)
	) name8942 (
		_w19303_,
		_w19304_,
		_w19454_
	);
	LUT2 #(
		.INIT('h1)
	) name8943 (
		_w19305_,
		_w19306_,
		_w19455_
	);
	LUT2 #(
		.INIT('h1)
	) name8944 (
		_w19307_,
		_w19308_,
		_w19456_
	);
	LUT2 #(
		.INIT('h1)
	) name8945 (
		_w19309_,
		_w19310_,
		_w19457_
	);
	LUT2 #(
		.INIT('h1)
	) name8946 (
		_w19311_,
		_w19312_,
		_w19458_
	);
	LUT2 #(
		.INIT('h1)
	) name8947 (
		_w19313_,
		_w19314_,
		_w19459_
	);
	LUT2 #(
		.INIT('h1)
	) name8948 (
		_w19315_,
		_w19316_,
		_w19460_
	);
	LUT2 #(
		.INIT('h1)
	) name8949 (
		_w19317_,
		_w19318_,
		_w19461_
	);
	LUT2 #(
		.INIT('h1)
	) name8950 (
		_w19319_,
		_w19320_,
		_w19462_
	);
	LUT2 #(
		.INIT('h1)
	) name8951 (
		_w19321_,
		_w19322_,
		_w19463_
	);
	LUT2 #(
		.INIT('h1)
	) name8952 (
		_w19323_,
		_w19324_,
		_w19464_
	);
	LUT2 #(
		.INIT('h1)
	) name8953 (
		_w19325_,
		_w19326_,
		_w19465_
	);
	LUT2 #(
		.INIT('h1)
	) name8954 (
		_w19327_,
		_w19328_,
		_w19466_
	);
	LUT2 #(
		.INIT('h1)
	) name8955 (
		_w19329_,
		_w19330_,
		_w19467_
	);
	LUT2 #(
		.INIT('h1)
	) name8956 (
		_w19331_,
		_w19332_,
		_w19468_
	);
	LUT2 #(
		.INIT('h1)
	) name8957 (
		_w19333_,
		_w19334_,
		_w19469_
	);
	LUT2 #(
		.INIT('h1)
	) name8958 (
		_w19335_,
		_w19336_,
		_w19470_
	);
	LUT2 #(
		.INIT('h1)
	) name8959 (
		_w19337_,
		_w19338_,
		_w19471_
	);
	LUT2 #(
		.INIT('h1)
	) name8960 (
		_w19339_,
		_w19340_,
		_w19472_
	);
	LUT2 #(
		.INIT('h1)
	) name8961 (
		_w19341_,
		_w19342_,
		_w19473_
	);
	LUT2 #(
		.INIT('h1)
	) name8962 (
		_w19343_,
		_w19344_,
		_w19474_
	);
	LUT2 #(
		.INIT('h1)
	) name8963 (
		_w19345_,
		_w19346_,
		_w19475_
	);
	LUT2 #(
		.INIT('h1)
	) name8964 (
		_w19347_,
		_w19348_,
		_w19476_
	);
	LUT2 #(
		.INIT('h8)
	) name8965 (
		_w19475_,
		_w19476_,
		_w19477_
	);
	LUT2 #(
		.INIT('h8)
	) name8966 (
		_w19473_,
		_w19474_,
		_w19478_
	);
	LUT2 #(
		.INIT('h8)
	) name8967 (
		_w19471_,
		_w19472_,
		_w19479_
	);
	LUT2 #(
		.INIT('h8)
	) name8968 (
		_w19469_,
		_w19470_,
		_w19480_
	);
	LUT2 #(
		.INIT('h8)
	) name8969 (
		_w19467_,
		_w19468_,
		_w19481_
	);
	LUT2 #(
		.INIT('h8)
	) name8970 (
		_w19465_,
		_w19466_,
		_w19482_
	);
	LUT2 #(
		.INIT('h8)
	) name8971 (
		_w19463_,
		_w19464_,
		_w19483_
	);
	LUT2 #(
		.INIT('h8)
	) name8972 (
		_w19461_,
		_w19462_,
		_w19484_
	);
	LUT2 #(
		.INIT('h8)
	) name8973 (
		_w19459_,
		_w19460_,
		_w19485_
	);
	LUT2 #(
		.INIT('h8)
	) name8974 (
		_w19457_,
		_w19458_,
		_w19486_
	);
	LUT2 #(
		.INIT('h8)
	) name8975 (
		_w19455_,
		_w19456_,
		_w19487_
	);
	LUT2 #(
		.INIT('h8)
	) name8976 (
		_w19453_,
		_w19454_,
		_w19488_
	);
	LUT2 #(
		.INIT('h8)
	) name8977 (
		_w19451_,
		_w19452_,
		_w19489_
	);
	LUT2 #(
		.INIT('h8)
	) name8978 (
		_w19449_,
		_w19450_,
		_w19490_
	);
	LUT2 #(
		.INIT('h8)
	) name8979 (
		_w19447_,
		_w19448_,
		_w19491_
	);
	LUT2 #(
		.INIT('h8)
	) name8980 (
		_w19445_,
		_w19446_,
		_w19492_
	);
	LUT2 #(
		.INIT('h8)
	) name8981 (
		_w19443_,
		_w19444_,
		_w19493_
	);
	LUT2 #(
		.INIT('h8)
	) name8982 (
		_w19441_,
		_w19442_,
		_w19494_
	);
	LUT2 #(
		.INIT('h8)
	) name8983 (
		_w19439_,
		_w19440_,
		_w19495_
	);
	LUT2 #(
		.INIT('h8)
	) name8984 (
		_w19437_,
		_w19438_,
		_w19496_
	);
	LUT2 #(
		.INIT('h8)
	) name8985 (
		_w19435_,
		_w19436_,
		_w19497_
	);
	LUT2 #(
		.INIT('h8)
	) name8986 (
		_w19433_,
		_w19434_,
		_w19498_
	);
	LUT2 #(
		.INIT('h8)
	) name8987 (
		_w19431_,
		_w19432_,
		_w19499_
	);
	LUT2 #(
		.INIT('h8)
	) name8988 (
		_w19429_,
		_w19430_,
		_w19500_
	);
	LUT2 #(
		.INIT('h8)
	) name8989 (
		_w19427_,
		_w19428_,
		_w19501_
	);
	LUT2 #(
		.INIT('h8)
	) name8990 (
		_w19425_,
		_w19426_,
		_w19502_
	);
	LUT2 #(
		.INIT('h8)
	) name8991 (
		_w19423_,
		_w19424_,
		_w19503_
	);
	LUT2 #(
		.INIT('h8)
	) name8992 (
		_w19421_,
		_w19422_,
		_w19504_
	);
	LUT2 #(
		.INIT('h8)
	) name8993 (
		_w19419_,
		_w19420_,
		_w19505_
	);
	LUT2 #(
		.INIT('h8)
	) name8994 (
		_w19417_,
		_w19418_,
		_w19506_
	);
	LUT2 #(
		.INIT('h8)
	) name8995 (
		_w19415_,
		_w19416_,
		_w19507_
	);
	LUT2 #(
		.INIT('h8)
	) name8996 (
		_w19413_,
		_w19414_,
		_w19508_
	);
	LUT2 #(
		.INIT('h8)
	) name8997 (
		_w19411_,
		_w19412_,
		_w19509_
	);
	LUT2 #(
		.INIT('h8)
	) name8998 (
		_w19409_,
		_w19410_,
		_w19510_
	);
	LUT2 #(
		.INIT('h8)
	) name8999 (
		_w19407_,
		_w19408_,
		_w19511_
	);
	LUT2 #(
		.INIT('h8)
	) name9000 (
		_w19405_,
		_w19406_,
		_w19512_
	);
	LUT2 #(
		.INIT('h8)
	) name9001 (
		_w19403_,
		_w19404_,
		_w19513_
	);
	LUT2 #(
		.INIT('h8)
	) name9002 (
		_w19401_,
		_w19402_,
		_w19514_
	);
	LUT2 #(
		.INIT('h8)
	) name9003 (
		_w19399_,
		_w19400_,
		_w19515_
	);
	LUT2 #(
		.INIT('h8)
	) name9004 (
		_w19397_,
		_w19398_,
		_w19516_
	);
	LUT2 #(
		.INIT('h8)
	) name9005 (
		_w19395_,
		_w19396_,
		_w19517_
	);
	LUT2 #(
		.INIT('h8)
	) name9006 (
		_w19393_,
		_w19394_,
		_w19518_
	);
	LUT2 #(
		.INIT('h8)
	) name9007 (
		_w19391_,
		_w19392_,
		_w19519_
	);
	LUT2 #(
		.INIT('h8)
	) name9008 (
		_w19389_,
		_w19390_,
		_w19520_
	);
	LUT2 #(
		.INIT('h8)
	) name9009 (
		_w19387_,
		_w19388_,
		_w19521_
	);
	LUT2 #(
		.INIT('h8)
	) name9010 (
		_w19385_,
		_w19386_,
		_w19522_
	);
	LUT2 #(
		.INIT('h8)
	) name9011 (
		_w19383_,
		_w19384_,
		_w19523_
	);
	LUT2 #(
		.INIT('h8)
	) name9012 (
		_w19381_,
		_w19382_,
		_w19524_
	);
	LUT2 #(
		.INIT('h8)
	) name9013 (
		_w19379_,
		_w19380_,
		_w19525_
	);
	LUT2 #(
		.INIT('h8)
	) name9014 (
		_w19377_,
		_w19378_,
		_w19526_
	);
	LUT2 #(
		.INIT('h8)
	) name9015 (
		_w19375_,
		_w19376_,
		_w19527_
	);
	LUT2 #(
		.INIT('h8)
	) name9016 (
		_w19373_,
		_w19374_,
		_w19528_
	);
	LUT2 #(
		.INIT('h8)
	) name9017 (
		_w19371_,
		_w19372_,
		_w19529_
	);
	LUT2 #(
		.INIT('h8)
	) name9018 (
		_w19369_,
		_w19370_,
		_w19530_
	);
	LUT2 #(
		.INIT('h8)
	) name9019 (
		_w19367_,
		_w19368_,
		_w19531_
	);
	LUT2 #(
		.INIT('h8)
	) name9020 (
		_w19365_,
		_w19366_,
		_w19532_
	);
	LUT2 #(
		.INIT('h8)
	) name9021 (
		_w19363_,
		_w19364_,
		_w19533_
	);
	LUT2 #(
		.INIT('h8)
	) name9022 (
		_w19361_,
		_w19362_,
		_w19534_
	);
	LUT2 #(
		.INIT('h8)
	) name9023 (
		_w19359_,
		_w19360_,
		_w19535_
	);
	LUT2 #(
		.INIT('h8)
	) name9024 (
		_w19357_,
		_w19358_,
		_w19536_
	);
	LUT2 #(
		.INIT('h8)
	) name9025 (
		_w19355_,
		_w19356_,
		_w19537_
	);
	LUT2 #(
		.INIT('h8)
	) name9026 (
		_w19353_,
		_w19354_,
		_w19538_
	);
	LUT2 #(
		.INIT('h8)
	) name9027 (
		_w19351_,
		_w19352_,
		_w19539_
	);
	LUT2 #(
		.INIT('h8)
	) name9028 (
		_w19349_,
		_w19350_,
		_w19540_
	);
	LUT2 #(
		.INIT('h8)
	) name9029 (
		_w19539_,
		_w19540_,
		_w19541_
	);
	LUT2 #(
		.INIT('h8)
	) name9030 (
		_w19537_,
		_w19538_,
		_w19542_
	);
	LUT2 #(
		.INIT('h8)
	) name9031 (
		_w19535_,
		_w19536_,
		_w19543_
	);
	LUT2 #(
		.INIT('h8)
	) name9032 (
		_w19533_,
		_w19534_,
		_w19544_
	);
	LUT2 #(
		.INIT('h8)
	) name9033 (
		_w19531_,
		_w19532_,
		_w19545_
	);
	LUT2 #(
		.INIT('h8)
	) name9034 (
		_w19529_,
		_w19530_,
		_w19546_
	);
	LUT2 #(
		.INIT('h8)
	) name9035 (
		_w19527_,
		_w19528_,
		_w19547_
	);
	LUT2 #(
		.INIT('h8)
	) name9036 (
		_w19525_,
		_w19526_,
		_w19548_
	);
	LUT2 #(
		.INIT('h8)
	) name9037 (
		_w19523_,
		_w19524_,
		_w19549_
	);
	LUT2 #(
		.INIT('h8)
	) name9038 (
		_w19521_,
		_w19522_,
		_w19550_
	);
	LUT2 #(
		.INIT('h8)
	) name9039 (
		_w19519_,
		_w19520_,
		_w19551_
	);
	LUT2 #(
		.INIT('h8)
	) name9040 (
		_w19517_,
		_w19518_,
		_w19552_
	);
	LUT2 #(
		.INIT('h8)
	) name9041 (
		_w19515_,
		_w19516_,
		_w19553_
	);
	LUT2 #(
		.INIT('h8)
	) name9042 (
		_w19513_,
		_w19514_,
		_w19554_
	);
	LUT2 #(
		.INIT('h8)
	) name9043 (
		_w19511_,
		_w19512_,
		_w19555_
	);
	LUT2 #(
		.INIT('h8)
	) name9044 (
		_w19509_,
		_w19510_,
		_w19556_
	);
	LUT2 #(
		.INIT('h8)
	) name9045 (
		_w19507_,
		_w19508_,
		_w19557_
	);
	LUT2 #(
		.INIT('h8)
	) name9046 (
		_w19505_,
		_w19506_,
		_w19558_
	);
	LUT2 #(
		.INIT('h8)
	) name9047 (
		_w19503_,
		_w19504_,
		_w19559_
	);
	LUT2 #(
		.INIT('h8)
	) name9048 (
		_w19501_,
		_w19502_,
		_w19560_
	);
	LUT2 #(
		.INIT('h8)
	) name9049 (
		_w19499_,
		_w19500_,
		_w19561_
	);
	LUT2 #(
		.INIT('h8)
	) name9050 (
		_w19497_,
		_w19498_,
		_w19562_
	);
	LUT2 #(
		.INIT('h8)
	) name9051 (
		_w19495_,
		_w19496_,
		_w19563_
	);
	LUT2 #(
		.INIT('h8)
	) name9052 (
		_w19493_,
		_w19494_,
		_w19564_
	);
	LUT2 #(
		.INIT('h8)
	) name9053 (
		_w19491_,
		_w19492_,
		_w19565_
	);
	LUT2 #(
		.INIT('h8)
	) name9054 (
		_w19489_,
		_w19490_,
		_w19566_
	);
	LUT2 #(
		.INIT('h8)
	) name9055 (
		_w19487_,
		_w19488_,
		_w19567_
	);
	LUT2 #(
		.INIT('h8)
	) name9056 (
		_w19485_,
		_w19486_,
		_w19568_
	);
	LUT2 #(
		.INIT('h8)
	) name9057 (
		_w19483_,
		_w19484_,
		_w19569_
	);
	LUT2 #(
		.INIT('h8)
	) name9058 (
		_w19481_,
		_w19482_,
		_w19570_
	);
	LUT2 #(
		.INIT('h8)
	) name9059 (
		_w19479_,
		_w19480_,
		_w19571_
	);
	LUT2 #(
		.INIT('h8)
	) name9060 (
		_w19477_,
		_w19478_,
		_w19572_
	);
	LUT2 #(
		.INIT('h8)
	) name9061 (
		_w19571_,
		_w19572_,
		_w19573_
	);
	LUT2 #(
		.INIT('h8)
	) name9062 (
		_w19569_,
		_w19570_,
		_w19574_
	);
	LUT2 #(
		.INIT('h8)
	) name9063 (
		_w19567_,
		_w19568_,
		_w19575_
	);
	LUT2 #(
		.INIT('h8)
	) name9064 (
		_w19565_,
		_w19566_,
		_w19576_
	);
	LUT2 #(
		.INIT('h8)
	) name9065 (
		_w19563_,
		_w19564_,
		_w19577_
	);
	LUT2 #(
		.INIT('h8)
	) name9066 (
		_w19561_,
		_w19562_,
		_w19578_
	);
	LUT2 #(
		.INIT('h8)
	) name9067 (
		_w19559_,
		_w19560_,
		_w19579_
	);
	LUT2 #(
		.INIT('h8)
	) name9068 (
		_w19557_,
		_w19558_,
		_w19580_
	);
	LUT2 #(
		.INIT('h8)
	) name9069 (
		_w19555_,
		_w19556_,
		_w19581_
	);
	LUT2 #(
		.INIT('h8)
	) name9070 (
		_w19553_,
		_w19554_,
		_w19582_
	);
	LUT2 #(
		.INIT('h8)
	) name9071 (
		_w19551_,
		_w19552_,
		_w19583_
	);
	LUT2 #(
		.INIT('h8)
	) name9072 (
		_w19549_,
		_w19550_,
		_w19584_
	);
	LUT2 #(
		.INIT('h8)
	) name9073 (
		_w19547_,
		_w19548_,
		_w19585_
	);
	LUT2 #(
		.INIT('h8)
	) name9074 (
		_w19545_,
		_w19546_,
		_w19586_
	);
	LUT2 #(
		.INIT('h8)
	) name9075 (
		_w19543_,
		_w19544_,
		_w19587_
	);
	LUT2 #(
		.INIT('h8)
	) name9076 (
		_w19541_,
		_w19542_,
		_w19588_
	);
	LUT2 #(
		.INIT('h8)
	) name9077 (
		_w19587_,
		_w19588_,
		_w19589_
	);
	LUT2 #(
		.INIT('h8)
	) name9078 (
		_w19585_,
		_w19586_,
		_w19590_
	);
	LUT2 #(
		.INIT('h8)
	) name9079 (
		_w19583_,
		_w19584_,
		_w19591_
	);
	LUT2 #(
		.INIT('h8)
	) name9080 (
		_w19581_,
		_w19582_,
		_w19592_
	);
	LUT2 #(
		.INIT('h8)
	) name9081 (
		_w19579_,
		_w19580_,
		_w19593_
	);
	LUT2 #(
		.INIT('h8)
	) name9082 (
		_w19577_,
		_w19578_,
		_w19594_
	);
	LUT2 #(
		.INIT('h8)
	) name9083 (
		_w19575_,
		_w19576_,
		_w19595_
	);
	LUT2 #(
		.INIT('h8)
	) name9084 (
		_w19573_,
		_w19574_,
		_w19596_
	);
	LUT2 #(
		.INIT('h8)
	) name9085 (
		_w19595_,
		_w19596_,
		_w19597_
	);
	LUT2 #(
		.INIT('h8)
	) name9086 (
		_w19593_,
		_w19594_,
		_w19598_
	);
	LUT2 #(
		.INIT('h8)
	) name9087 (
		_w19591_,
		_w19592_,
		_w19599_
	);
	LUT2 #(
		.INIT('h8)
	) name9088 (
		_w19589_,
		_w19590_,
		_w19600_
	);
	LUT2 #(
		.INIT('h8)
	) name9089 (
		_w19599_,
		_w19600_,
		_w19601_
	);
	LUT2 #(
		.INIT('h8)
	) name9090 (
		_w19597_,
		_w19598_,
		_w19602_
	);
	LUT2 #(
		.INIT('h8)
	) name9091 (
		_w19601_,
		_w19602_,
		_w19603_
	);
	LUT2 #(
		.INIT('h1)
	) name9092 (
		wb_rst_i_pad,
		_w19603_,
		_w19604_
	);
	LUT2 #(
		.INIT('h2)
	) name9093 (
		_w12656_,
		_w19604_,
		_w19605_
	);
	LUT2 #(
		.INIT('h8)
	) name9094 (
		_w13497_,
		_w17290_,
		_w19606_
	);
	LUT2 #(
		.INIT('h2)
	) name9095 (
		\wishbone_TxLength_reg[15]/NET0131 ,
		_w19606_,
		_w19607_
	);
	LUT2 #(
		.INIT('h1)
	) name9096 (
		_w12656_,
		_w19607_,
		_w19608_
	);
	LUT2 #(
		.INIT('h1)
	) name9097 (
		_w19605_,
		_w19608_,
		_w19609_
	);
	LUT2 #(
		.INIT('h1)
	) name9098 (
		_w13486_,
		_w13487_,
		_w19610_
	);
	LUT2 #(
		.INIT('h8)
	) name9099 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19610_,
		_w19611_
	);
	LUT2 #(
		.INIT('h1)
	) name9100 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w19610_,
		_w19612_
	);
	LUT2 #(
		.INIT('h1)
	) name9101 (
		_w19611_,
		_w19612_,
		_w19613_
	);
	LUT2 #(
		.INIT('h8)
	) name9102 (
		_w13501_,
		_w19613_,
		_w19614_
	);
	LUT2 #(
		.INIT('h8)
	) name9103 (
		\wishbone_bd_ram_mem2_reg[26][17]/P0001 ,
		_w12699_,
		_w19615_
	);
	LUT2 #(
		.INIT('h8)
	) name9104 (
		\wishbone_bd_ram_mem2_reg[125][17]/P0001 ,
		_w12956_,
		_w19616_
	);
	LUT2 #(
		.INIT('h8)
	) name9105 (
		\wishbone_bd_ram_mem2_reg[89][17]/P0001 ,
		_w12964_,
		_w19617_
	);
	LUT2 #(
		.INIT('h8)
	) name9106 (
		\wishbone_bd_ram_mem2_reg[136][17]/P0001 ,
		_w13064_,
		_w19618_
	);
	LUT2 #(
		.INIT('h8)
	) name9107 (
		\wishbone_bd_ram_mem2_reg[145][17]/P0001 ,
		_w13106_,
		_w19619_
	);
	LUT2 #(
		.INIT('h8)
	) name9108 (
		\wishbone_bd_ram_mem2_reg[61][17]/P0001 ,
		_w12725_,
		_w19620_
	);
	LUT2 #(
		.INIT('h8)
	) name9109 (
		\wishbone_bd_ram_mem2_reg[55][17]/P0001 ,
		_w12785_,
		_w19621_
	);
	LUT2 #(
		.INIT('h8)
	) name9110 (
		\wishbone_bd_ram_mem2_reg[242][17]/P0001 ,
		_w12932_,
		_w19622_
	);
	LUT2 #(
		.INIT('h8)
	) name9111 (
		\wishbone_bd_ram_mem2_reg[30][17]/P0001 ,
		_w13104_,
		_w19623_
	);
	LUT2 #(
		.INIT('h8)
	) name9112 (
		\wishbone_bd_ram_mem2_reg[70][17]/P0001 ,
		_w12840_,
		_w19624_
	);
	LUT2 #(
		.INIT('h8)
	) name9113 (
		\wishbone_bd_ram_mem2_reg[46][17]/P0001 ,
		_w12884_,
		_w19625_
	);
	LUT2 #(
		.INIT('h8)
	) name9114 (
		\wishbone_bd_ram_mem2_reg[131][17]/P0001 ,
		_w12852_,
		_w19626_
	);
	LUT2 #(
		.INIT('h8)
	) name9115 (
		\wishbone_bd_ram_mem2_reg[167][17]/P0001 ,
		_w12986_,
		_w19627_
	);
	LUT2 #(
		.INIT('h8)
	) name9116 (
		\wishbone_bd_ram_mem2_reg[42][17]/P0001 ,
		_w12842_,
		_w19628_
	);
	LUT2 #(
		.INIT('h8)
	) name9117 (
		\wishbone_bd_ram_mem2_reg[27][17]/P0001 ,
		_w12880_,
		_w19629_
	);
	LUT2 #(
		.INIT('h8)
	) name9118 (
		\wishbone_bd_ram_mem2_reg[87][17]/P0001 ,
		_w13154_,
		_w19630_
	);
	LUT2 #(
		.INIT('h8)
	) name9119 (
		\wishbone_bd_ram_mem2_reg[147][17]/P0001 ,
		_w13146_,
		_w19631_
	);
	LUT2 #(
		.INIT('h8)
	) name9120 (
		\wishbone_bd_ram_mem2_reg[14][17]/P0001 ,
		_w13086_,
		_w19632_
	);
	LUT2 #(
		.INIT('h8)
	) name9121 (
		\wishbone_bd_ram_mem2_reg[48][17]/P0001 ,
		_w12970_,
		_w19633_
	);
	LUT2 #(
		.INIT('h8)
	) name9122 (
		\wishbone_bd_ram_mem2_reg[175][17]/P0001 ,
		_w13126_,
		_w19634_
	);
	LUT2 #(
		.INIT('h8)
	) name9123 (
		\wishbone_bd_ram_mem2_reg[130][17]/P0001 ,
		_w12914_,
		_w19635_
	);
	LUT2 #(
		.INIT('h8)
	) name9124 (
		\wishbone_bd_ram_mem2_reg[192][17]/P0001 ,
		_w12938_,
		_w19636_
	);
	LUT2 #(
		.INIT('h8)
	) name9125 (
		\wishbone_bd_ram_mem2_reg[218][17]/P0001 ,
		_w13206_,
		_w19637_
	);
	LUT2 #(
		.INIT('h8)
	) name9126 (
		\wishbone_bd_ram_mem2_reg[181][17]/P0001 ,
		_w12828_,
		_w19638_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		\wishbone_bd_ram_mem2_reg[226][17]/P0001 ,
		_w13138_,
		_w19639_
	);
	LUT2 #(
		.INIT('h8)
	) name9128 (
		\wishbone_bd_ram_mem2_reg[249][17]/P0001 ,
		_w12900_,
		_w19640_
	);
	LUT2 #(
		.INIT('h8)
	) name9129 (
		\wishbone_bd_ram_mem2_reg[25][17]/P0001 ,
		_w13108_,
		_w19641_
	);
	LUT2 #(
		.INIT('h8)
	) name9130 (
		\wishbone_bd_ram_mem2_reg[227][17]/P0001 ,
		_w12936_,
		_w19642_
	);
	LUT2 #(
		.INIT('h8)
	) name9131 (
		\wishbone_bd_ram_mem2_reg[250][17]/P0001 ,
		_w13128_,
		_w19643_
	);
	LUT2 #(
		.INIT('h8)
	) name9132 (
		\wishbone_bd_ram_mem2_reg[174][17]/P0001 ,
		_w12972_,
		_w19644_
	);
	LUT2 #(
		.INIT('h8)
	) name9133 (
		\wishbone_bd_ram_mem2_reg[223][17]/P0001 ,
		_w12838_,
		_w19645_
	);
	LUT2 #(
		.INIT('h8)
	) name9134 (
		\wishbone_bd_ram_mem2_reg[77][17]/P0001 ,
		_w12982_,
		_w19646_
	);
	LUT2 #(
		.INIT('h8)
	) name9135 (
		\wishbone_bd_ram_mem2_reg[185][17]/P0001 ,
		_w12940_,
		_w19647_
	);
	LUT2 #(
		.INIT('h8)
	) name9136 (
		\wishbone_bd_ram_mem2_reg[21][17]/P0001 ,
		_w12906_,
		_w19648_
	);
	LUT2 #(
		.INIT('h8)
	) name9137 (
		\wishbone_bd_ram_mem2_reg[73][17]/P0001 ,
		_w12918_,
		_w19649_
	);
	LUT2 #(
		.INIT('h8)
	) name9138 (
		\wishbone_bd_ram_mem2_reg[219][17]/P0001 ,
		_w12806_,
		_w19650_
	);
	LUT2 #(
		.INIT('h8)
	) name9139 (
		\wishbone_bd_ram_mem2_reg[98][17]/P0001 ,
		_w12816_,
		_w19651_
	);
	LUT2 #(
		.INIT('h8)
	) name9140 (
		\wishbone_bd_ram_mem2_reg[236][17]/P0001 ,
		_w12731_,
		_w19652_
	);
	LUT2 #(
		.INIT('h8)
	) name9141 (
		\wishbone_bd_ram_mem2_reg[37][17]/P0001 ,
		_w13102_,
		_w19653_
	);
	LUT2 #(
		.INIT('h8)
	) name9142 (
		\wishbone_bd_ram_mem2_reg[66][17]/P0001 ,
		_w12824_,
		_w19654_
	);
	LUT2 #(
		.INIT('h8)
	) name9143 (
		\wishbone_bd_ram_mem2_reg[16][17]/P0001 ,
		_w13140_,
		_w19655_
	);
	LUT2 #(
		.INIT('h8)
	) name9144 (
		\wishbone_bd_ram_mem2_reg[126][17]/P0001 ,
		_w13218_,
		_w19656_
	);
	LUT2 #(
		.INIT('h8)
	) name9145 (
		\wishbone_bd_ram_mem2_reg[228][17]/P0001 ,
		_w12765_,
		_w19657_
	);
	LUT2 #(
		.INIT('h8)
	) name9146 (
		\wishbone_bd_ram_mem2_reg[80][17]/P0001 ,
		_w12689_,
		_w19658_
	);
	LUT2 #(
		.INIT('h8)
	) name9147 (
		\wishbone_bd_ram_mem2_reg[129][17]/P0001 ,
		_w12776_,
		_w19659_
	);
	LUT2 #(
		.INIT('h8)
	) name9148 (
		\wishbone_bd_ram_mem2_reg[62][17]/P0001 ,
		_w12673_,
		_w19660_
	);
	LUT2 #(
		.INIT('h8)
	) name9149 (
		\wishbone_bd_ram_mem2_reg[82][17]/P0001 ,
		_w12942_,
		_w19661_
	);
	LUT2 #(
		.INIT('h8)
	) name9150 (
		\wishbone_bd_ram_mem2_reg[156][17]/P0001 ,
		_w13190_,
		_w19662_
	);
	LUT2 #(
		.INIT('h8)
	) name9151 (
		\wishbone_bd_ram_mem2_reg[111][17]/P0001 ,
		_w12744_,
		_w19663_
	);
	LUT2 #(
		.INIT('h8)
	) name9152 (
		\wishbone_bd_ram_mem2_reg[152][17]/P0001 ,
		_w12966_,
		_w19664_
	);
	LUT2 #(
		.INIT('h8)
	) name9153 (
		\wishbone_bd_ram_mem2_reg[177][17]/P0001 ,
		_w12996_,
		_w19665_
	);
	LUT2 #(
		.INIT('h8)
	) name9154 (
		\wishbone_bd_ram_mem2_reg[52][17]/P0001 ,
		_w13082_,
		_w19666_
	);
	LUT2 #(
		.INIT('h8)
	) name9155 (
		\wishbone_bd_ram_mem2_reg[158][17]/P0001 ,
		_w12898_,
		_w19667_
	);
	LUT2 #(
		.INIT('h8)
	) name9156 (
		\wishbone_bd_ram_mem2_reg[43][17]/P0001 ,
		_w13200_,
		_w19668_
	);
	LUT2 #(
		.INIT('h8)
	) name9157 (
		\wishbone_bd_ram_mem2_reg[11][17]/P0001 ,
		_w13194_,
		_w19669_
	);
	LUT2 #(
		.INIT('h8)
	) name9158 (
		\wishbone_bd_ram_mem2_reg[178][17]/P0001 ,
		_w12886_,
		_w19670_
	);
	LUT2 #(
		.INIT('h8)
	) name9159 (
		\wishbone_bd_ram_mem2_reg[67][17]/P0001 ,
		_w13134_,
		_w19671_
	);
	LUT2 #(
		.INIT('h8)
	) name9160 (
		\wishbone_bd_ram_mem2_reg[0][17]/P0001 ,
		_w12717_,
		_w19672_
	);
	LUT2 #(
		.INIT('h8)
	) name9161 (
		\wishbone_bd_ram_mem2_reg[72][17]/P0001 ,
		_w12810_,
		_w19673_
	);
	LUT2 #(
		.INIT('h8)
	) name9162 (
		\wishbone_bd_ram_mem2_reg[2][17]/P0001 ,
		_w13088_,
		_w19674_
	);
	LUT2 #(
		.INIT('h8)
	) name9163 (
		\wishbone_bd_ram_mem2_reg[139][17]/P0001 ,
		_w12814_,
		_w19675_
	);
	LUT2 #(
		.INIT('h8)
	) name9164 (
		\wishbone_bd_ram_mem2_reg[116][17]/P0001 ,
		_w12998_,
		_w19676_
	);
	LUT2 #(
		.INIT('h8)
	) name9165 (
		\wishbone_bd_ram_mem2_reg[36][17]/P0001 ,
		_w12800_,
		_w19677_
	);
	LUT2 #(
		.INIT('h8)
	) name9166 (
		\wishbone_bd_ram_mem2_reg[201][17]/P0001 ,
		_w12822_,
		_w19678_
	);
	LUT2 #(
		.INIT('h8)
	) name9167 (
		\wishbone_bd_ram_mem2_reg[22][17]/P0001 ,
		_w13110_,
		_w19679_
	);
	LUT2 #(
		.INIT('h8)
	) name9168 (
		\wishbone_bd_ram_mem2_reg[84][17]/P0001 ,
		_w12934_,
		_w19680_
	);
	LUT2 #(
		.INIT('h8)
	) name9169 (
		\wishbone_bd_ram_mem2_reg[60][17]/P0001 ,
		_w13204_,
		_w19681_
	);
	LUT2 #(
		.INIT('h8)
	) name9170 (
		\wishbone_bd_ram_mem2_reg[10][17]/P0001 ,
		_w13172_,
		_w19682_
	);
	LUT2 #(
		.INIT('h8)
	) name9171 (
		\wishbone_bd_ram_mem2_reg[143][17]/P0001 ,
		_w12922_,
		_w19683_
	);
	LUT2 #(
		.INIT('h8)
	) name9172 (
		\wishbone_bd_ram_mem2_reg[102][17]/P0001 ,
		_w12685_,
		_w19684_
	);
	LUT2 #(
		.INIT('h8)
	) name9173 (
		\wishbone_bd_ram_mem2_reg[90][17]/P0001 ,
		_w12978_,
		_w19685_
	);
	LUT2 #(
		.INIT('h8)
	) name9174 (
		\wishbone_bd_ram_mem2_reg[176][17]/P0001 ,
		_w12868_,
		_w19686_
	);
	LUT2 #(
		.INIT('h8)
	) name9175 (
		\wishbone_bd_ram_mem2_reg[19][17]/P0001 ,
		_w13012_,
		_w19687_
	);
	LUT2 #(
		.INIT('h8)
	) name9176 (
		\wishbone_bd_ram_mem2_reg[243][17]/P0001 ,
		_w12804_,
		_w19688_
	);
	LUT2 #(
		.INIT('h8)
	) name9177 (
		\wishbone_bd_ram_mem2_reg[122][17]/P0001 ,
		_w13130_,
		_w19689_
	);
	LUT2 #(
		.INIT('h8)
	) name9178 (
		\wishbone_bd_ram_mem2_reg[34][17]/P0001 ,
		_w12930_,
		_w19690_
	);
	LUT2 #(
		.INIT('h8)
	) name9179 (
		\wishbone_bd_ram_mem2_reg[9][17]/P0001 ,
		_w12808_,
		_w19691_
	);
	LUT2 #(
		.INIT('h8)
	) name9180 (
		\wishbone_bd_ram_mem2_reg[234][17]/P0001 ,
		_w13214_,
		_w19692_
	);
	LUT2 #(
		.INIT('h8)
	) name9181 (
		\wishbone_bd_ram_mem2_reg[168][17]/P0001 ,
		_w13208_,
		_w19693_
	);
	LUT2 #(
		.INIT('h8)
	) name9182 (
		\wishbone_bd_ram_mem2_reg[231][17]/P0001 ,
		_w12856_,
		_w19694_
	);
	LUT2 #(
		.INIT('h8)
	) name9183 (
		\wishbone_bd_ram_mem2_reg[13][17]/P0001 ,
		_w13178_,
		_w19695_
	);
	LUT2 #(
		.INIT('h8)
	) name9184 (
		\wishbone_bd_ram_mem2_reg[12][17]/P0001 ,
		_w13118_,
		_w19696_
	);
	LUT2 #(
		.INIT('h8)
	) name9185 (
		\wishbone_bd_ram_mem2_reg[51][17]/P0001 ,
		_w13024_,
		_w19697_
	);
	LUT2 #(
		.INIT('h8)
	) name9186 (
		\wishbone_bd_ram_mem2_reg[183][17]/P0001 ,
		_w12787_,
		_w19698_
	);
	LUT2 #(
		.INIT('h8)
	) name9187 (
		\wishbone_bd_ram_mem2_reg[173][17]/P0001 ,
		_w12854_,
		_w19699_
	);
	LUT2 #(
		.INIT('h8)
	) name9188 (
		\wishbone_bd_ram_mem2_reg[105][17]/P0001 ,
		_w12751_,
		_w19700_
	);
	LUT2 #(
		.INIT('h8)
	) name9189 (
		\wishbone_bd_ram_mem2_reg[212][17]/P0001 ,
		_w12796_,
		_w19701_
	);
	LUT2 #(
		.INIT('h8)
	) name9190 (
		\wishbone_bd_ram_mem2_reg[209][17]/P0001 ,
		_w13152_,
		_w19702_
	);
	LUT2 #(
		.INIT('h8)
	) name9191 (
		\wishbone_bd_ram_mem2_reg[213][17]/P0001 ,
		_w13002_,
		_w19703_
	);
	LUT2 #(
		.INIT('h8)
	) name9192 (
		\wishbone_bd_ram_mem2_reg[166][17]/P0001 ,
		_w13040_,
		_w19704_
	);
	LUT2 #(
		.INIT('h8)
	) name9193 (
		\wishbone_bd_ram_mem2_reg[117][17]/P0001 ,
		_w12715_,
		_w19705_
	);
	LUT2 #(
		.INIT('h8)
	) name9194 (
		\wishbone_bd_ram_mem2_reg[23][17]/P0001 ,
		_w13008_,
		_w19706_
	);
	LUT2 #(
		.INIT('h8)
	) name9195 (
		\wishbone_bd_ram_mem2_reg[161][17]/P0001 ,
		_w12754_,
		_w19707_
	);
	LUT2 #(
		.INIT('h8)
	) name9196 (
		\wishbone_bd_ram_mem2_reg[33][17]/P0001 ,
		_w12980_,
		_w19708_
	);
	LUT2 #(
		.INIT('h8)
	) name9197 (
		\wishbone_bd_ram_mem2_reg[76][17]/P0001 ,
		_w13184_,
		_w19709_
	);
	LUT2 #(
		.INIT('h8)
	) name9198 (
		\wishbone_bd_ram_mem2_reg[57][17]/P0001 ,
		_w13116_,
		_w19710_
	);
	LUT2 #(
		.INIT('h8)
	) name9199 (
		\wishbone_bd_ram_mem2_reg[134][17]/P0001 ,
		_w12763_,
		_w19711_
	);
	LUT2 #(
		.INIT('h8)
	) name9200 (
		\wishbone_bd_ram_mem2_reg[93][17]/P0001 ,
		_w13016_,
		_w19712_
	);
	LUT2 #(
		.INIT('h8)
	) name9201 (
		\wishbone_bd_ram_mem2_reg[56][17]/P0001 ,
		_w12778_,
		_w19713_
	);
	LUT2 #(
		.INIT('h8)
	) name9202 (
		\wishbone_bd_ram_mem2_reg[133][17]/P0001 ,
		_w12761_,
		_w19714_
	);
	LUT2 #(
		.INIT('h8)
	) name9203 (
		\wishbone_bd_ram_mem2_reg[49][17]/P0001 ,
		_w12994_,
		_w19715_
	);
	LUT2 #(
		.INIT('h8)
	) name9204 (
		\wishbone_bd_ram_mem2_reg[107][17]/P0001 ,
		_w12749_,
		_w19716_
	);
	LUT2 #(
		.INIT('h8)
	) name9205 (
		\wishbone_bd_ram_mem2_reg[184][17]/P0001 ,
		_w13062_,
		_w19717_
	);
	LUT2 #(
		.INIT('h8)
	) name9206 (
		\wishbone_bd_ram_mem2_reg[97][17]/P0001 ,
		_w13096_,
		_w19718_
	);
	LUT2 #(
		.INIT('h8)
	) name9207 (
		\wishbone_bd_ram_mem2_reg[45][17]/P0001 ,
		_w12908_,
		_w19719_
	);
	LUT2 #(
		.INIT('h8)
	) name9208 (
		\wishbone_bd_ram_mem2_reg[233][17]/P0001 ,
		_w12836_,
		_w19720_
	);
	LUT2 #(
		.INIT('h8)
	) name9209 (
		\wishbone_bd_ram_mem2_reg[162][17]/P0001 ,
		_w13098_,
		_w19721_
	);
	LUT2 #(
		.INIT('h8)
	) name9210 (
		\wishbone_bd_ram_mem2_reg[29][17]/P0001 ,
		_w12952_,
		_w19722_
	);
	LUT2 #(
		.INIT('h8)
	) name9211 (
		\wishbone_bd_ram_mem2_reg[195][17]/P0001 ,
		_w13144_,
		_w19723_
	);
	LUT2 #(
		.INIT('h8)
	) name9212 (
		\wishbone_bd_ram_mem2_reg[198][17]/P0001 ,
		_w12832_,
		_w19724_
	);
	LUT2 #(
		.INIT('h8)
	) name9213 (
		\wishbone_bd_ram_mem2_reg[240][17]/P0001 ,
		_w12864_,
		_w19725_
	);
	LUT2 #(
		.INIT('h8)
	) name9214 (
		\wishbone_bd_ram_mem2_reg[210][17]/P0001 ,
		_w12924_,
		_w19726_
	);
	LUT2 #(
		.INIT('h8)
	) name9215 (
		\wishbone_bd_ram_mem2_reg[119][17]/P0001 ,
		_w13048_,
		_w19727_
	);
	LUT2 #(
		.INIT('h8)
	) name9216 (
		\wishbone_bd_ram_mem2_reg[214][17]/P0001 ,
		_w12984_,
		_w19728_
	);
	LUT2 #(
		.INIT('h8)
	) name9217 (
		\wishbone_bd_ram_mem2_reg[96][17]/P0001 ,
		_w12912_,
		_w19729_
	);
	LUT2 #(
		.INIT('h8)
	) name9218 (
		\wishbone_bd_ram_mem2_reg[92][17]/P0001 ,
		_w13010_,
		_w19730_
	);
	LUT2 #(
		.INIT('h8)
	) name9219 (
		\wishbone_bd_ram_mem2_reg[146][17]/P0001 ,
		_w13060_,
		_w19731_
	);
	LUT2 #(
		.INIT('h8)
	) name9220 (
		\wishbone_bd_ram_mem2_reg[15][17]/P0001 ,
		_w13210_,
		_w19732_
	);
	LUT2 #(
		.INIT('h8)
	) name9221 (
		\wishbone_bd_ram_mem2_reg[44][17]/P0001 ,
		_w12896_,
		_w19733_
	);
	LUT2 #(
		.INIT('h8)
	) name9222 (
		\wishbone_bd_ram_mem2_reg[64][17]/P0001 ,
		_w12976_,
		_w19734_
	);
	LUT2 #(
		.INIT('h8)
	) name9223 (
		\wishbone_bd_ram_mem2_reg[63][17]/P0001 ,
		_w12850_,
		_w19735_
	);
	LUT2 #(
		.INIT('h8)
	) name9224 (
		\wishbone_bd_ram_mem2_reg[69][17]/P0001 ,
		_w12738_,
		_w19736_
	);
	LUT2 #(
		.INIT('h8)
	) name9225 (
		\wishbone_bd_ram_mem2_reg[85][17]/P0001 ,
		_w13216_,
		_w19737_
	);
	LUT2 #(
		.INIT('h8)
	) name9226 (
		\wishbone_bd_ram_mem2_reg[229][17]/P0001 ,
		_w12711_,
		_w19738_
	);
	LUT2 #(
		.INIT('h8)
	) name9227 (
		\wishbone_bd_ram_mem2_reg[253][17]/P0001 ,
		_w13100_,
		_w19739_
	);
	LUT2 #(
		.INIT('h8)
	) name9228 (
		\wishbone_bd_ram_mem2_reg[132][17]/P0001 ,
		_w12992_,
		_w19740_
	);
	LUT2 #(
		.INIT('h8)
	) name9229 (
		\wishbone_bd_ram_mem2_reg[149][17]/P0001 ,
		_w12741_,
		_w19741_
	);
	LUT2 #(
		.INIT('h8)
	) name9230 (
		\wishbone_bd_ram_mem2_reg[124][17]/P0001 ,
		_w13058_,
		_w19742_
	);
	LUT2 #(
		.INIT('h8)
	) name9231 (
		\wishbone_bd_ram_mem2_reg[205][17]/P0001 ,
		_w13068_,
		_w19743_
	);
	LUT2 #(
		.INIT('h8)
	) name9232 (
		\wishbone_bd_ram_mem2_reg[155][17]/P0001 ,
		_w13122_,
		_w19744_
	);
	LUT2 #(
		.INIT('h8)
	) name9233 (
		\wishbone_bd_ram_mem2_reg[230][17]/P0001 ,
		_w13036_,
		_w19745_
	);
	LUT2 #(
		.INIT('h8)
	) name9234 (
		\wishbone_bd_ram_mem2_reg[20][17]/P0001 ,
		_w13174_,
		_w19746_
	);
	LUT2 #(
		.INIT('h8)
	) name9235 (
		\wishbone_bd_ram_mem2_reg[172][17]/P0001 ,
		_w12944_,
		_w19747_
	);
	LUT2 #(
		.INIT('h8)
	) name9236 (
		\wishbone_bd_ram_mem2_reg[153][17]/P0001 ,
		_w12890_,
		_w19748_
	);
	LUT2 #(
		.INIT('h8)
	) name9237 (
		\wishbone_bd_ram_mem2_reg[220][17]/P0001 ,
		_w13066_,
		_w19749_
	);
	LUT2 #(
		.INIT('h8)
	) name9238 (
		\wishbone_bd_ram_mem2_reg[112][17]/P0001 ,
		_w12733_,
		_w19750_
	);
	LUT2 #(
		.INIT('h8)
	) name9239 (
		\wishbone_bd_ram_mem2_reg[3][17]/P0001 ,
		_w12866_,
		_w19751_
	);
	LUT2 #(
		.INIT('h8)
	) name9240 (
		\wishbone_bd_ram_mem2_reg[245][17]/P0001 ,
		_w13022_,
		_w19752_
	);
	LUT2 #(
		.INIT('h8)
	) name9241 (
		\wishbone_bd_ram_mem2_reg[118][17]/P0001 ,
		_w12830_,
		_w19753_
	);
	LUT2 #(
		.INIT('h8)
	) name9242 (
		\wishbone_bd_ram_mem2_reg[28][17]/P0001 ,
		_w13170_,
		_w19754_
	);
	LUT2 #(
		.INIT('h8)
	) name9243 (
		\wishbone_bd_ram_mem2_reg[58][17]/P0001 ,
		_w13070_,
		_w19755_
	);
	LUT2 #(
		.INIT('h8)
	) name9244 (
		\wishbone_bd_ram_mem2_reg[138][17]/P0001 ,
		_w12958_,
		_w19756_
	);
	LUT2 #(
		.INIT('h8)
	) name9245 (
		\wishbone_bd_ram_mem2_reg[35][17]/P0001 ,
		_w12703_,
		_w19757_
	);
	LUT2 #(
		.INIT('h8)
	) name9246 (
		\wishbone_bd_ram_mem2_reg[222][17]/P0001 ,
		_w13094_,
		_w19758_
	);
	LUT2 #(
		.INIT('h8)
	) name9247 (
		\wishbone_bd_ram_mem2_reg[165][17]/P0001 ,
		_w13044_,
		_w19759_
	);
	LUT2 #(
		.INIT('h8)
	) name9248 (
		\wishbone_bd_ram_mem2_reg[1][17]/P0001 ,
		_w13014_,
		_w19760_
	);
	LUT2 #(
		.INIT('h8)
	) name9249 (
		\wishbone_bd_ram_mem2_reg[244][17]/P0001 ,
		_w12747_,
		_w19761_
	);
	LUT2 #(
		.INIT('h8)
	) name9250 (
		\wishbone_bd_ram_mem2_reg[247][17]/P0001 ,
		_w12818_,
		_w19762_
	);
	LUT2 #(
		.INIT('h8)
	) name9251 (
		\wishbone_bd_ram_mem2_reg[200][17]/P0001 ,
		_w12988_,
		_w19763_
	);
	LUT2 #(
		.INIT('h8)
	) name9252 (
		\wishbone_bd_ram_mem2_reg[248][17]/P0001 ,
		_w12789_,
		_w19764_
	);
	LUT2 #(
		.INIT('h8)
	) name9253 (
		\wishbone_bd_ram_mem2_reg[31][17]/P0001 ,
		_w13198_,
		_w19765_
	);
	LUT2 #(
		.INIT('h8)
	) name9254 (
		\wishbone_bd_ram_mem2_reg[232][17]/P0001 ,
		_w12758_,
		_w19766_
	);
	LUT2 #(
		.INIT('h8)
	) name9255 (
		\wishbone_bd_ram_mem2_reg[163][17]/P0001 ,
		_w12882_,
		_w19767_
	);
	LUT2 #(
		.INIT('h8)
	) name9256 (
		\wishbone_bd_ram_mem2_reg[208][17]/P0001 ,
		_w13032_,
		_w19768_
	);
	LUT2 #(
		.INIT('h8)
	) name9257 (
		\wishbone_bd_ram_mem2_reg[101][17]/P0001 ,
		_w13192_,
		_w19769_
	);
	LUT2 #(
		.INIT('h8)
	) name9258 (
		\wishbone_bd_ram_mem2_reg[211][17]/P0001 ,
		_w13166_,
		_w19770_
	);
	LUT2 #(
		.INIT('h8)
	) name9259 (
		\wishbone_bd_ram_mem2_reg[239][17]/P0001 ,
		_w12862_,
		_w19771_
	);
	LUT2 #(
		.INIT('h8)
	) name9260 (
		\wishbone_bd_ram_mem2_reg[123][17]/P0001 ,
		_w13114_,
		_w19772_
	);
	LUT2 #(
		.INIT('h8)
	) name9261 (
		\wishbone_bd_ram_mem2_reg[99][17]/P0001 ,
		_w13038_,
		_w19773_
	);
	LUT2 #(
		.INIT('h8)
	) name9262 (
		\wishbone_bd_ram_mem2_reg[86][17]/P0001 ,
		_w12735_,
		_w19774_
	);
	LUT2 #(
		.INIT('h8)
	) name9263 (
		\wishbone_bd_ram_mem2_reg[78][17]/P0001 ,
		_w12874_,
		_w19775_
	);
	LUT2 #(
		.INIT('h8)
	) name9264 (
		\wishbone_bd_ram_mem2_reg[207][17]/P0001 ,
		_w13180_,
		_w19776_
	);
	LUT2 #(
		.INIT('h8)
	) name9265 (
		\wishbone_bd_ram_mem2_reg[128][17]/P0001 ,
		_w12793_,
		_w19777_
	);
	LUT2 #(
		.INIT('h8)
	) name9266 (
		\wishbone_bd_ram_mem2_reg[24][17]/P0001 ,
		_w13084_,
		_w19778_
	);
	LUT2 #(
		.INIT('h8)
	) name9267 (
		\wishbone_bd_ram_mem2_reg[41][17]/P0001 ,
		_w13052_,
		_w19779_
	);
	LUT2 #(
		.INIT('h8)
	) name9268 (
		\wishbone_bd_ram_mem2_reg[160][17]/P0001 ,
		_w12872_,
		_w19780_
	);
	LUT2 #(
		.INIT('h8)
	) name9269 (
		\wishbone_bd_ram_mem2_reg[217][17]/P0001 ,
		_w13188_,
		_w19781_
	);
	LUT2 #(
		.INIT('h8)
	) name9270 (
		\wishbone_bd_ram_mem2_reg[142][17]/P0001 ,
		_w12928_,
		_w19782_
	);
	LUT2 #(
		.INIT('h8)
	) name9271 (
		\wishbone_bd_ram_mem2_reg[32][17]/P0001 ,
		_w13120_,
		_w19783_
	);
	LUT2 #(
		.INIT('h8)
	) name9272 (
		\wishbone_bd_ram_mem2_reg[50][17]/P0001 ,
		_w13150_,
		_w19784_
	);
	LUT2 #(
		.INIT('h8)
	) name9273 (
		\wishbone_bd_ram_mem2_reg[148][17]/P0001 ,
		_w13000_,
		_w19785_
	);
	LUT2 #(
		.INIT('h8)
	) name9274 (
		\wishbone_bd_ram_mem2_reg[237][17]/P0001 ,
		_w12990_,
		_w19786_
	);
	LUT2 #(
		.INIT('h8)
	) name9275 (
		\wishbone_bd_ram_mem2_reg[127][17]/P0001 ,
		_w13164_,
		_w19787_
	);
	LUT2 #(
		.INIT('h8)
	) name9276 (
		\wishbone_bd_ram_mem2_reg[40][17]/P0001 ,
		_w13132_,
		_w19788_
	);
	LUT2 #(
		.INIT('h8)
	) name9277 (
		\wishbone_bd_ram_mem2_reg[151][17]/P0001 ,
		_w13142_,
		_w19789_
	);
	LUT2 #(
		.INIT('h8)
	) name9278 (
		\wishbone_bd_ram_mem2_reg[71][17]/P0001 ,
		_w12798_,
		_w19790_
	);
	LUT2 #(
		.INIT('h8)
	) name9279 (
		\wishbone_bd_ram_mem2_reg[91][17]/P0001 ,
		_w13074_,
		_w19791_
	);
	LUT2 #(
		.INIT('h8)
	) name9280 (
		\wishbone_bd_ram_mem2_reg[221][17]/P0001 ,
		_w12802_,
		_w19792_
	);
	LUT2 #(
		.INIT('h8)
	) name9281 (
		\wishbone_bd_ram_mem2_reg[206][17]/P0001 ,
		_w12954_,
		_w19793_
	);
	LUT2 #(
		.INIT('h8)
	) name9282 (
		\wishbone_bd_ram_mem2_reg[194][17]/P0001 ,
		_w12772_,
		_w19794_
	);
	LUT2 #(
		.INIT('h8)
	) name9283 (
		\wishbone_bd_ram_mem2_reg[187][17]/P0001 ,
		_w13196_,
		_w19795_
	);
	LUT2 #(
		.INIT('h8)
	) name9284 (
		\wishbone_bd_ram_mem2_reg[137][17]/P0001 ,
		_w13168_,
		_w19796_
	);
	LUT2 #(
		.INIT('h8)
	) name9285 (
		\wishbone_bd_ram_mem2_reg[8][17]/P0001 ,
		_w12920_,
		_w19797_
	);
	LUT2 #(
		.INIT('h8)
	) name9286 (
		\wishbone_bd_ram_mem2_reg[53][17]/P0001 ,
		_w13020_,
		_w19798_
	);
	LUT2 #(
		.INIT('h8)
	) name9287 (
		\wishbone_bd_ram_mem2_reg[113][17]/P0001 ,
		_w13026_,
		_w19799_
	);
	LUT2 #(
		.INIT('h8)
	) name9288 (
		\wishbone_bd_ram_mem2_reg[65][17]/P0001 ,
		_w13176_,
		_w19800_
	);
	LUT2 #(
		.INIT('h8)
	) name9289 (
		\wishbone_bd_ram_mem2_reg[180][17]/P0001 ,
		_w12791_,
		_w19801_
	);
	LUT2 #(
		.INIT('h8)
	) name9290 (
		\wishbone_bd_ram_mem2_reg[193][17]/P0001 ,
		_w13056_,
		_w19802_
	);
	LUT2 #(
		.INIT('h8)
	) name9291 (
		\wishbone_bd_ram_mem2_reg[39][17]/P0001 ,
		_w13018_,
		_w19803_
	);
	LUT2 #(
		.INIT('h8)
	) name9292 (
		\wishbone_bd_ram_mem2_reg[144][17]/P0001 ,
		_w12756_,
		_w19804_
	);
	LUT2 #(
		.INIT('h8)
	) name9293 (
		\wishbone_bd_ram_mem2_reg[47][17]/P0001 ,
		_w12904_,
		_w19805_
	);
	LUT2 #(
		.INIT('h8)
	) name9294 (
		\wishbone_bd_ram_mem2_reg[251][17]/P0001 ,
		_w13054_,
		_w19806_
	);
	LUT2 #(
		.INIT('h8)
	) name9295 (
		\wishbone_bd_ram_mem2_reg[59][17]/P0001 ,
		_w12780_,
		_w19807_
	);
	LUT2 #(
		.INIT('h8)
	) name9296 (
		\wishbone_bd_ram_mem2_reg[204][17]/P0001 ,
		_w13162_,
		_w19808_
	);
	LUT2 #(
		.INIT('h8)
	) name9297 (
		\wishbone_bd_ram_mem2_reg[88][17]/P0001 ,
		_w12860_,
		_w19809_
	);
	LUT2 #(
		.INIT('h8)
	) name9298 (
		\wishbone_bd_ram_mem2_reg[182][17]/P0001 ,
		_w12820_,
		_w19810_
	);
	LUT2 #(
		.INIT('h8)
	) name9299 (
		\wishbone_bd_ram_mem2_reg[189][17]/P0001 ,
		_w13042_,
		_w19811_
	);
	LUT2 #(
		.INIT('h8)
	) name9300 (
		\wishbone_bd_ram_mem2_reg[75][17]/P0001 ,
		_w12826_,
		_w19812_
	);
	LUT2 #(
		.INIT('h8)
	) name9301 (
		\wishbone_bd_ram_mem2_reg[197][17]/P0001 ,
		_w12834_,
		_w19813_
	);
	LUT2 #(
		.INIT('h8)
	) name9302 (
		\wishbone_bd_ram_mem2_reg[254][17]/P0001 ,
		_w12892_,
		_w19814_
	);
	LUT2 #(
		.INIT('h8)
	) name9303 (
		\wishbone_bd_ram_mem2_reg[199][17]/P0001 ,
		_w12768_,
		_w19815_
	);
	LUT2 #(
		.INIT('h8)
	) name9304 (
		\wishbone_bd_ram_mem2_reg[141][17]/P0001 ,
		_w13004_,
		_w19816_
	);
	LUT2 #(
		.INIT('h8)
	) name9305 (
		\wishbone_bd_ram_mem2_reg[159][17]/P0001 ,
		_w12774_,
		_w19817_
	);
	LUT2 #(
		.INIT('h8)
	) name9306 (
		\wishbone_bd_ram_mem2_reg[169][17]/P0001 ,
		_w12722_,
		_w19818_
	);
	LUT2 #(
		.INIT('h8)
	) name9307 (
		\wishbone_bd_ram_mem2_reg[17][17]/P0001 ,
		_w12848_,
		_w19819_
	);
	LUT2 #(
		.INIT('h8)
	) name9308 (
		\wishbone_bd_ram_mem2_reg[103][17]/P0001 ,
		_w12846_,
		_w19820_
	);
	LUT2 #(
		.INIT('h8)
	) name9309 (
		\wishbone_bd_ram_mem2_reg[120][17]/P0001 ,
		_w12707_,
		_w19821_
	);
	LUT2 #(
		.INIT('h8)
	) name9310 (
		\wishbone_bd_ram_mem2_reg[190][17]/P0001 ,
		_w12858_,
		_w19822_
	);
	LUT2 #(
		.INIT('h8)
	) name9311 (
		\wishbone_bd_ram_mem2_reg[104][17]/P0001 ,
		_w13148_,
		_w19823_
	);
	LUT2 #(
		.INIT('h8)
	) name9312 (
		\wishbone_bd_ram_mem2_reg[154][17]/P0001 ,
		_w12962_,
		_w19824_
	);
	LUT2 #(
		.INIT('h8)
	) name9313 (
		\wishbone_bd_ram_mem2_reg[115][17]/P0001 ,
		_w13112_,
		_w19825_
	);
	LUT2 #(
		.INIT('h8)
	) name9314 (
		\wishbone_bd_ram_mem2_reg[108][17]/P0001 ,
		_w13156_,
		_w19826_
	);
	LUT2 #(
		.INIT('h8)
	) name9315 (
		\wishbone_bd_ram_mem2_reg[224][17]/P0001 ,
		_w12902_,
		_w19827_
	);
	LUT2 #(
		.INIT('h8)
	) name9316 (
		\wishbone_bd_ram_mem2_reg[179][17]/P0001 ,
		_w13050_,
		_w19828_
	);
	LUT2 #(
		.INIT('h8)
	) name9317 (
		\wishbone_bd_ram_mem2_reg[54][17]/P0001 ,
		_w12770_,
		_w19829_
	);
	LUT2 #(
		.INIT('h8)
	) name9318 (
		\wishbone_bd_ram_mem2_reg[5][17]/P0001 ,
		_w12878_,
		_w19830_
	);
	LUT2 #(
		.INIT('h8)
	) name9319 (
		\wishbone_bd_ram_mem2_reg[202][17]/P0001 ,
		_w12870_,
		_w19831_
	);
	LUT2 #(
		.INIT('h8)
	) name9320 (
		\wishbone_bd_ram_mem2_reg[110][17]/P0001 ,
		_w13046_,
		_w19832_
	);
	LUT2 #(
		.INIT('h8)
	) name9321 (
		\wishbone_bd_ram_mem2_reg[135][17]/P0001 ,
		_w13124_,
		_w19833_
	);
	LUT2 #(
		.INIT('h8)
	) name9322 (
		\wishbone_bd_ram_mem2_reg[109][17]/P0001 ,
		_w12888_,
		_w19834_
	);
	LUT2 #(
		.INIT('h8)
	) name9323 (
		\wishbone_bd_ram_mem2_reg[196][17]/P0001 ,
		_w13090_,
		_w19835_
	);
	LUT2 #(
		.INIT('h8)
	) name9324 (
		\wishbone_bd_ram_mem2_reg[114][17]/P0001 ,
		_w13202_,
		_w19836_
	);
	LUT2 #(
		.INIT('h8)
	) name9325 (
		\wishbone_bd_ram_mem2_reg[38][17]/P0001 ,
		_w13182_,
		_w19837_
	);
	LUT2 #(
		.INIT('h8)
	) name9326 (
		\wishbone_bd_ram_mem2_reg[215][17]/P0001 ,
		_w12974_,
		_w19838_
	);
	LUT2 #(
		.INIT('h8)
	) name9327 (
		\wishbone_bd_ram_mem2_reg[216][17]/P0001 ,
		_w13028_,
		_w19839_
	);
	LUT2 #(
		.INIT('h8)
	) name9328 (
		\wishbone_bd_ram_mem2_reg[225][17]/P0001 ,
		_w13092_,
		_w19840_
	);
	LUT2 #(
		.INIT('h8)
	) name9329 (
		\wishbone_bd_ram_mem2_reg[203][17]/P0001 ,
		_w13158_,
		_w19841_
	);
	LUT2 #(
		.INIT('h8)
	) name9330 (
		\wishbone_bd_ram_mem2_reg[4][17]/P0001 ,
		_w12666_,
		_w19842_
	);
	LUT2 #(
		.INIT('h8)
	) name9331 (
		\wishbone_bd_ram_mem2_reg[252][17]/P0001 ,
		_w13080_,
		_w19843_
	);
	LUT2 #(
		.INIT('h8)
	) name9332 (
		\wishbone_bd_ram_mem2_reg[191][17]/P0001 ,
		_w13034_,
		_w19844_
	);
	LUT2 #(
		.INIT('h8)
	) name9333 (
		\wishbone_bd_ram_mem2_reg[7][17]/P0001 ,
		_w12728_,
		_w19845_
	);
	LUT2 #(
		.INIT('h8)
	) name9334 (
		\wishbone_bd_ram_mem2_reg[100][17]/P0001 ,
		_w12960_,
		_w19846_
	);
	LUT2 #(
		.INIT('h8)
	) name9335 (
		\wishbone_bd_ram_mem2_reg[6][17]/P0001 ,
		_w12968_,
		_w19847_
	);
	LUT2 #(
		.INIT('h8)
	) name9336 (
		\wishbone_bd_ram_mem2_reg[157][17]/P0001 ,
		_w12926_,
		_w19848_
	);
	LUT2 #(
		.INIT('h8)
	) name9337 (
		\wishbone_bd_ram_mem2_reg[241][17]/P0001 ,
		_w13006_,
		_w19849_
	);
	LUT2 #(
		.INIT('h8)
	) name9338 (
		\wishbone_bd_ram_mem2_reg[186][17]/P0001 ,
		_w12783_,
		_w19850_
	);
	LUT2 #(
		.INIT('h8)
	) name9339 (
		\wishbone_bd_ram_mem2_reg[74][17]/P0001 ,
		_w12812_,
		_w19851_
	);
	LUT2 #(
		.INIT('h8)
	) name9340 (
		\wishbone_bd_ram_mem2_reg[164][17]/P0001 ,
		_w12876_,
		_w19852_
	);
	LUT2 #(
		.INIT('h8)
	) name9341 (
		\wishbone_bd_ram_mem2_reg[83][17]/P0001 ,
		_w12916_,
		_w19853_
	);
	LUT2 #(
		.INIT('h8)
	) name9342 (
		\wishbone_bd_ram_mem2_reg[121][17]/P0001 ,
		_w13078_,
		_w19854_
	);
	LUT2 #(
		.INIT('h8)
	) name9343 (
		\wishbone_bd_ram_mem2_reg[235][17]/P0001 ,
		_w12696_,
		_w19855_
	);
	LUT2 #(
		.INIT('h8)
	) name9344 (
		\wishbone_bd_ram_mem2_reg[94][17]/P0001 ,
		_w13186_,
		_w19856_
	);
	LUT2 #(
		.INIT('h8)
	) name9345 (
		\wishbone_bd_ram_mem2_reg[106][17]/P0001 ,
		_w12713_,
		_w19857_
	);
	LUT2 #(
		.INIT('h8)
	) name9346 (
		\wishbone_bd_ram_mem2_reg[79][17]/P0001 ,
		_w13212_,
		_w19858_
	);
	LUT2 #(
		.INIT('h8)
	) name9347 (
		\wishbone_bd_ram_mem2_reg[18][17]/P0001 ,
		_w12679_,
		_w19859_
	);
	LUT2 #(
		.INIT('h8)
	) name9348 (
		\wishbone_bd_ram_mem2_reg[68][17]/P0001 ,
		_w12946_,
		_w19860_
	);
	LUT2 #(
		.INIT('h8)
	) name9349 (
		\wishbone_bd_ram_mem2_reg[95][17]/P0001 ,
		_w12844_,
		_w19861_
	);
	LUT2 #(
		.INIT('h8)
	) name9350 (
		\wishbone_bd_ram_mem2_reg[170][17]/P0001 ,
		_w13030_,
		_w19862_
	);
	LUT2 #(
		.INIT('h8)
	) name9351 (
		\wishbone_bd_ram_mem2_reg[246][17]/P0001 ,
		_w13076_,
		_w19863_
	);
	LUT2 #(
		.INIT('h8)
	) name9352 (
		\wishbone_bd_ram_mem2_reg[150][17]/P0001 ,
		_w13136_,
		_w19864_
	);
	LUT2 #(
		.INIT('h8)
	) name9353 (
		\wishbone_bd_ram_mem2_reg[140][17]/P0001 ,
		_w12894_,
		_w19865_
	);
	LUT2 #(
		.INIT('h8)
	) name9354 (
		\wishbone_bd_ram_mem2_reg[255][17]/P0001 ,
		_w13072_,
		_w19866_
	);
	LUT2 #(
		.INIT('h8)
	) name9355 (
		\wishbone_bd_ram_mem2_reg[188][17]/P0001 ,
		_w12948_,
		_w19867_
	);
	LUT2 #(
		.INIT('h8)
	) name9356 (
		\wishbone_bd_ram_mem2_reg[81][17]/P0001 ,
		_w12950_,
		_w19868_
	);
	LUT2 #(
		.INIT('h8)
	) name9357 (
		\wishbone_bd_ram_mem2_reg[171][17]/P0001 ,
		_w12910_,
		_w19869_
	);
	LUT2 #(
		.INIT('h8)
	) name9358 (
		\wishbone_bd_ram_mem2_reg[238][17]/P0001 ,
		_w13160_,
		_w19870_
	);
	LUT2 #(
		.INIT('h1)
	) name9359 (
		_w19615_,
		_w19616_,
		_w19871_
	);
	LUT2 #(
		.INIT('h1)
	) name9360 (
		_w19617_,
		_w19618_,
		_w19872_
	);
	LUT2 #(
		.INIT('h1)
	) name9361 (
		_w19619_,
		_w19620_,
		_w19873_
	);
	LUT2 #(
		.INIT('h1)
	) name9362 (
		_w19621_,
		_w19622_,
		_w19874_
	);
	LUT2 #(
		.INIT('h1)
	) name9363 (
		_w19623_,
		_w19624_,
		_w19875_
	);
	LUT2 #(
		.INIT('h1)
	) name9364 (
		_w19625_,
		_w19626_,
		_w19876_
	);
	LUT2 #(
		.INIT('h1)
	) name9365 (
		_w19627_,
		_w19628_,
		_w19877_
	);
	LUT2 #(
		.INIT('h1)
	) name9366 (
		_w19629_,
		_w19630_,
		_w19878_
	);
	LUT2 #(
		.INIT('h1)
	) name9367 (
		_w19631_,
		_w19632_,
		_w19879_
	);
	LUT2 #(
		.INIT('h1)
	) name9368 (
		_w19633_,
		_w19634_,
		_w19880_
	);
	LUT2 #(
		.INIT('h1)
	) name9369 (
		_w19635_,
		_w19636_,
		_w19881_
	);
	LUT2 #(
		.INIT('h1)
	) name9370 (
		_w19637_,
		_w19638_,
		_w19882_
	);
	LUT2 #(
		.INIT('h1)
	) name9371 (
		_w19639_,
		_w19640_,
		_w19883_
	);
	LUT2 #(
		.INIT('h1)
	) name9372 (
		_w19641_,
		_w19642_,
		_w19884_
	);
	LUT2 #(
		.INIT('h1)
	) name9373 (
		_w19643_,
		_w19644_,
		_w19885_
	);
	LUT2 #(
		.INIT('h1)
	) name9374 (
		_w19645_,
		_w19646_,
		_w19886_
	);
	LUT2 #(
		.INIT('h1)
	) name9375 (
		_w19647_,
		_w19648_,
		_w19887_
	);
	LUT2 #(
		.INIT('h1)
	) name9376 (
		_w19649_,
		_w19650_,
		_w19888_
	);
	LUT2 #(
		.INIT('h1)
	) name9377 (
		_w19651_,
		_w19652_,
		_w19889_
	);
	LUT2 #(
		.INIT('h1)
	) name9378 (
		_w19653_,
		_w19654_,
		_w19890_
	);
	LUT2 #(
		.INIT('h1)
	) name9379 (
		_w19655_,
		_w19656_,
		_w19891_
	);
	LUT2 #(
		.INIT('h1)
	) name9380 (
		_w19657_,
		_w19658_,
		_w19892_
	);
	LUT2 #(
		.INIT('h1)
	) name9381 (
		_w19659_,
		_w19660_,
		_w19893_
	);
	LUT2 #(
		.INIT('h1)
	) name9382 (
		_w19661_,
		_w19662_,
		_w19894_
	);
	LUT2 #(
		.INIT('h1)
	) name9383 (
		_w19663_,
		_w19664_,
		_w19895_
	);
	LUT2 #(
		.INIT('h1)
	) name9384 (
		_w19665_,
		_w19666_,
		_w19896_
	);
	LUT2 #(
		.INIT('h1)
	) name9385 (
		_w19667_,
		_w19668_,
		_w19897_
	);
	LUT2 #(
		.INIT('h1)
	) name9386 (
		_w19669_,
		_w19670_,
		_w19898_
	);
	LUT2 #(
		.INIT('h1)
	) name9387 (
		_w19671_,
		_w19672_,
		_w19899_
	);
	LUT2 #(
		.INIT('h1)
	) name9388 (
		_w19673_,
		_w19674_,
		_w19900_
	);
	LUT2 #(
		.INIT('h1)
	) name9389 (
		_w19675_,
		_w19676_,
		_w19901_
	);
	LUT2 #(
		.INIT('h1)
	) name9390 (
		_w19677_,
		_w19678_,
		_w19902_
	);
	LUT2 #(
		.INIT('h1)
	) name9391 (
		_w19679_,
		_w19680_,
		_w19903_
	);
	LUT2 #(
		.INIT('h1)
	) name9392 (
		_w19681_,
		_w19682_,
		_w19904_
	);
	LUT2 #(
		.INIT('h1)
	) name9393 (
		_w19683_,
		_w19684_,
		_w19905_
	);
	LUT2 #(
		.INIT('h1)
	) name9394 (
		_w19685_,
		_w19686_,
		_w19906_
	);
	LUT2 #(
		.INIT('h1)
	) name9395 (
		_w19687_,
		_w19688_,
		_w19907_
	);
	LUT2 #(
		.INIT('h1)
	) name9396 (
		_w19689_,
		_w19690_,
		_w19908_
	);
	LUT2 #(
		.INIT('h1)
	) name9397 (
		_w19691_,
		_w19692_,
		_w19909_
	);
	LUT2 #(
		.INIT('h1)
	) name9398 (
		_w19693_,
		_w19694_,
		_w19910_
	);
	LUT2 #(
		.INIT('h1)
	) name9399 (
		_w19695_,
		_w19696_,
		_w19911_
	);
	LUT2 #(
		.INIT('h1)
	) name9400 (
		_w19697_,
		_w19698_,
		_w19912_
	);
	LUT2 #(
		.INIT('h1)
	) name9401 (
		_w19699_,
		_w19700_,
		_w19913_
	);
	LUT2 #(
		.INIT('h1)
	) name9402 (
		_w19701_,
		_w19702_,
		_w19914_
	);
	LUT2 #(
		.INIT('h1)
	) name9403 (
		_w19703_,
		_w19704_,
		_w19915_
	);
	LUT2 #(
		.INIT('h1)
	) name9404 (
		_w19705_,
		_w19706_,
		_w19916_
	);
	LUT2 #(
		.INIT('h1)
	) name9405 (
		_w19707_,
		_w19708_,
		_w19917_
	);
	LUT2 #(
		.INIT('h1)
	) name9406 (
		_w19709_,
		_w19710_,
		_w19918_
	);
	LUT2 #(
		.INIT('h1)
	) name9407 (
		_w19711_,
		_w19712_,
		_w19919_
	);
	LUT2 #(
		.INIT('h1)
	) name9408 (
		_w19713_,
		_w19714_,
		_w19920_
	);
	LUT2 #(
		.INIT('h1)
	) name9409 (
		_w19715_,
		_w19716_,
		_w19921_
	);
	LUT2 #(
		.INIT('h1)
	) name9410 (
		_w19717_,
		_w19718_,
		_w19922_
	);
	LUT2 #(
		.INIT('h1)
	) name9411 (
		_w19719_,
		_w19720_,
		_w19923_
	);
	LUT2 #(
		.INIT('h1)
	) name9412 (
		_w19721_,
		_w19722_,
		_w19924_
	);
	LUT2 #(
		.INIT('h1)
	) name9413 (
		_w19723_,
		_w19724_,
		_w19925_
	);
	LUT2 #(
		.INIT('h1)
	) name9414 (
		_w19725_,
		_w19726_,
		_w19926_
	);
	LUT2 #(
		.INIT('h1)
	) name9415 (
		_w19727_,
		_w19728_,
		_w19927_
	);
	LUT2 #(
		.INIT('h1)
	) name9416 (
		_w19729_,
		_w19730_,
		_w19928_
	);
	LUT2 #(
		.INIT('h1)
	) name9417 (
		_w19731_,
		_w19732_,
		_w19929_
	);
	LUT2 #(
		.INIT('h1)
	) name9418 (
		_w19733_,
		_w19734_,
		_w19930_
	);
	LUT2 #(
		.INIT('h1)
	) name9419 (
		_w19735_,
		_w19736_,
		_w19931_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		_w19737_,
		_w19738_,
		_w19932_
	);
	LUT2 #(
		.INIT('h1)
	) name9421 (
		_w19739_,
		_w19740_,
		_w19933_
	);
	LUT2 #(
		.INIT('h1)
	) name9422 (
		_w19741_,
		_w19742_,
		_w19934_
	);
	LUT2 #(
		.INIT('h1)
	) name9423 (
		_w19743_,
		_w19744_,
		_w19935_
	);
	LUT2 #(
		.INIT('h1)
	) name9424 (
		_w19745_,
		_w19746_,
		_w19936_
	);
	LUT2 #(
		.INIT('h1)
	) name9425 (
		_w19747_,
		_w19748_,
		_w19937_
	);
	LUT2 #(
		.INIT('h1)
	) name9426 (
		_w19749_,
		_w19750_,
		_w19938_
	);
	LUT2 #(
		.INIT('h1)
	) name9427 (
		_w19751_,
		_w19752_,
		_w19939_
	);
	LUT2 #(
		.INIT('h1)
	) name9428 (
		_w19753_,
		_w19754_,
		_w19940_
	);
	LUT2 #(
		.INIT('h1)
	) name9429 (
		_w19755_,
		_w19756_,
		_w19941_
	);
	LUT2 #(
		.INIT('h1)
	) name9430 (
		_w19757_,
		_w19758_,
		_w19942_
	);
	LUT2 #(
		.INIT('h1)
	) name9431 (
		_w19759_,
		_w19760_,
		_w19943_
	);
	LUT2 #(
		.INIT('h1)
	) name9432 (
		_w19761_,
		_w19762_,
		_w19944_
	);
	LUT2 #(
		.INIT('h1)
	) name9433 (
		_w19763_,
		_w19764_,
		_w19945_
	);
	LUT2 #(
		.INIT('h1)
	) name9434 (
		_w19765_,
		_w19766_,
		_w19946_
	);
	LUT2 #(
		.INIT('h1)
	) name9435 (
		_w19767_,
		_w19768_,
		_w19947_
	);
	LUT2 #(
		.INIT('h1)
	) name9436 (
		_w19769_,
		_w19770_,
		_w19948_
	);
	LUT2 #(
		.INIT('h1)
	) name9437 (
		_w19771_,
		_w19772_,
		_w19949_
	);
	LUT2 #(
		.INIT('h1)
	) name9438 (
		_w19773_,
		_w19774_,
		_w19950_
	);
	LUT2 #(
		.INIT('h1)
	) name9439 (
		_w19775_,
		_w19776_,
		_w19951_
	);
	LUT2 #(
		.INIT('h1)
	) name9440 (
		_w19777_,
		_w19778_,
		_w19952_
	);
	LUT2 #(
		.INIT('h1)
	) name9441 (
		_w19779_,
		_w19780_,
		_w19953_
	);
	LUT2 #(
		.INIT('h1)
	) name9442 (
		_w19781_,
		_w19782_,
		_w19954_
	);
	LUT2 #(
		.INIT('h1)
	) name9443 (
		_w19783_,
		_w19784_,
		_w19955_
	);
	LUT2 #(
		.INIT('h1)
	) name9444 (
		_w19785_,
		_w19786_,
		_w19956_
	);
	LUT2 #(
		.INIT('h1)
	) name9445 (
		_w19787_,
		_w19788_,
		_w19957_
	);
	LUT2 #(
		.INIT('h1)
	) name9446 (
		_w19789_,
		_w19790_,
		_w19958_
	);
	LUT2 #(
		.INIT('h1)
	) name9447 (
		_w19791_,
		_w19792_,
		_w19959_
	);
	LUT2 #(
		.INIT('h1)
	) name9448 (
		_w19793_,
		_w19794_,
		_w19960_
	);
	LUT2 #(
		.INIT('h1)
	) name9449 (
		_w19795_,
		_w19796_,
		_w19961_
	);
	LUT2 #(
		.INIT('h1)
	) name9450 (
		_w19797_,
		_w19798_,
		_w19962_
	);
	LUT2 #(
		.INIT('h1)
	) name9451 (
		_w19799_,
		_w19800_,
		_w19963_
	);
	LUT2 #(
		.INIT('h1)
	) name9452 (
		_w19801_,
		_w19802_,
		_w19964_
	);
	LUT2 #(
		.INIT('h1)
	) name9453 (
		_w19803_,
		_w19804_,
		_w19965_
	);
	LUT2 #(
		.INIT('h1)
	) name9454 (
		_w19805_,
		_w19806_,
		_w19966_
	);
	LUT2 #(
		.INIT('h1)
	) name9455 (
		_w19807_,
		_w19808_,
		_w19967_
	);
	LUT2 #(
		.INIT('h1)
	) name9456 (
		_w19809_,
		_w19810_,
		_w19968_
	);
	LUT2 #(
		.INIT('h1)
	) name9457 (
		_w19811_,
		_w19812_,
		_w19969_
	);
	LUT2 #(
		.INIT('h1)
	) name9458 (
		_w19813_,
		_w19814_,
		_w19970_
	);
	LUT2 #(
		.INIT('h1)
	) name9459 (
		_w19815_,
		_w19816_,
		_w19971_
	);
	LUT2 #(
		.INIT('h1)
	) name9460 (
		_w19817_,
		_w19818_,
		_w19972_
	);
	LUT2 #(
		.INIT('h1)
	) name9461 (
		_w19819_,
		_w19820_,
		_w19973_
	);
	LUT2 #(
		.INIT('h1)
	) name9462 (
		_w19821_,
		_w19822_,
		_w19974_
	);
	LUT2 #(
		.INIT('h1)
	) name9463 (
		_w19823_,
		_w19824_,
		_w19975_
	);
	LUT2 #(
		.INIT('h1)
	) name9464 (
		_w19825_,
		_w19826_,
		_w19976_
	);
	LUT2 #(
		.INIT('h1)
	) name9465 (
		_w19827_,
		_w19828_,
		_w19977_
	);
	LUT2 #(
		.INIT('h1)
	) name9466 (
		_w19829_,
		_w19830_,
		_w19978_
	);
	LUT2 #(
		.INIT('h1)
	) name9467 (
		_w19831_,
		_w19832_,
		_w19979_
	);
	LUT2 #(
		.INIT('h1)
	) name9468 (
		_w19833_,
		_w19834_,
		_w19980_
	);
	LUT2 #(
		.INIT('h1)
	) name9469 (
		_w19835_,
		_w19836_,
		_w19981_
	);
	LUT2 #(
		.INIT('h1)
	) name9470 (
		_w19837_,
		_w19838_,
		_w19982_
	);
	LUT2 #(
		.INIT('h1)
	) name9471 (
		_w19839_,
		_w19840_,
		_w19983_
	);
	LUT2 #(
		.INIT('h1)
	) name9472 (
		_w19841_,
		_w19842_,
		_w19984_
	);
	LUT2 #(
		.INIT('h1)
	) name9473 (
		_w19843_,
		_w19844_,
		_w19985_
	);
	LUT2 #(
		.INIT('h1)
	) name9474 (
		_w19845_,
		_w19846_,
		_w19986_
	);
	LUT2 #(
		.INIT('h1)
	) name9475 (
		_w19847_,
		_w19848_,
		_w19987_
	);
	LUT2 #(
		.INIT('h1)
	) name9476 (
		_w19849_,
		_w19850_,
		_w19988_
	);
	LUT2 #(
		.INIT('h1)
	) name9477 (
		_w19851_,
		_w19852_,
		_w19989_
	);
	LUT2 #(
		.INIT('h1)
	) name9478 (
		_w19853_,
		_w19854_,
		_w19990_
	);
	LUT2 #(
		.INIT('h1)
	) name9479 (
		_w19855_,
		_w19856_,
		_w19991_
	);
	LUT2 #(
		.INIT('h1)
	) name9480 (
		_w19857_,
		_w19858_,
		_w19992_
	);
	LUT2 #(
		.INIT('h1)
	) name9481 (
		_w19859_,
		_w19860_,
		_w19993_
	);
	LUT2 #(
		.INIT('h1)
	) name9482 (
		_w19861_,
		_w19862_,
		_w19994_
	);
	LUT2 #(
		.INIT('h1)
	) name9483 (
		_w19863_,
		_w19864_,
		_w19995_
	);
	LUT2 #(
		.INIT('h1)
	) name9484 (
		_w19865_,
		_w19866_,
		_w19996_
	);
	LUT2 #(
		.INIT('h1)
	) name9485 (
		_w19867_,
		_w19868_,
		_w19997_
	);
	LUT2 #(
		.INIT('h1)
	) name9486 (
		_w19869_,
		_w19870_,
		_w19998_
	);
	LUT2 #(
		.INIT('h8)
	) name9487 (
		_w19997_,
		_w19998_,
		_w19999_
	);
	LUT2 #(
		.INIT('h8)
	) name9488 (
		_w19995_,
		_w19996_,
		_w20000_
	);
	LUT2 #(
		.INIT('h8)
	) name9489 (
		_w19993_,
		_w19994_,
		_w20001_
	);
	LUT2 #(
		.INIT('h8)
	) name9490 (
		_w19991_,
		_w19992_,
		_w20002_
	);
	LUT2 #(
		.INIT('h8)
	) name9491 (
		_w19989_,
		_w19990_,
		_w20003_
	);
	LUT2 #(
		.INIT('h8)
	) name9492 (
		_w19987_,
		_w19988_,
		_w20004_
	);
	LUT2 #(
		.INIT('h8)
	) name9493 (
		_w19985_,
		_w19986_,
		_w20005_
	);
	LUT2 #(
		.INIT('h8)
	) name9494 (
		_w19983_,
		_w19984_,
		_w20006_
	);
	LUT2 #(
		.INIT('h8)
	) name9495 (
		_w19981_,
		_w19982_,
		_w20007_
	);
	LUT2 #(
		.INIT('h8)
	) name9496 (
		_w19979_,
		_w19980_,
		_w20008_
	);
	LUT2 #(
		.INIT('h8)
	) name9497 (
		_w19977_,
		_w19978_,
		_w20009_
	);
	LUT2 #(
		.INIT('h8)
	) name9498 (
		_w19975_,
		_w19976_,
		_w20010_
	);
	LUT2 #(
		.INIT('h8)
	) name9499 (
		_w19973_,
		_w19974_,
		_w20011_
	);
	LUT2 #(
		.INIT('h8)
	) name9500 (
		_w19971_,
		_w19972_,
		_w20012_
	);
	LUT2 #(
		.INIT('h8)
	) name9501 (
		_w19969_,
		_w19970_,
		_w20013_
	);
	LUT2 #(
		.INIT('h8)
	) name9502 (
		_w19967_,
		_w19968_,
		_w20014_
	);
	LUT2 #(
		.INIT('h8)
	) name9503 (
		_w19965_,
		_w19966_,
		_w20015_
	);
	LUT2 #(
		.INIT('h8)
	) name9504 (
		_w19963_,
		_w19964_,
		_w20016_
	);
	LUT2 #(
		.INIT('h8)
	) name9505 (
		_w19961_,
		_w19962_,
		_w20017_
	);
	LUT2 #(
		.INIT('h8)
	) name9506 (
		_w19959_,
		_w19960_,
		_w20018_
	);
	LUT2 #(
		.INIT('h8)
	) name9507 (
		_w19957_,
		_w19958_,
		_w20019_
	);
	LUT2 #(
		.INIT('h8)
	) name9508 (
		_w19955_,
		_w19956_,
		_w20020_
	);
	LUT2 #(
		.INIT('h8)
	) name9509 (
		_w19953_,
		_w19954_,
		_w20021_
	);
	LUT2 #(
		.INIT('h8)
	) name9510 (
		_w19951_,
		_w19952_,
		_w20022_
	);
	LUT2 #(
		.INIT('h8)
	) name9511 (
		_w19949_,
		_w19950_,
		_w20023_
	);
	LUT2 #(
		.INIT('h8)
	) name9512 (
		_w19947_,
		_w19948_,
		_w20024_
	);
	LUT2 #(
		.INIT('h8)
	) name9513 (
		_w19945_,
		_w19946_,
		_w20025_
	);
	LUT2 #(
		.INIT('h8)
	) name9514 (
		_w19943_,
		_w19944_,
		_w20026_
	);
	LUT2 #(
		.INIT('h8)
	) name9515 (
		_w19941_,
		_w19942_,
		_w20027_
	);
	LUT2 #(
		.INIT('h8)
	) name9516 (
		_w19939_,
		_w19940_,
		_w20028_
	);
	LUT2 #(
		.INIT('h8)
	) name9517 (
		_w19937_,
		_w19938_,
		_w20029_
	);
	LUT2 #(
		.INIT('h8)
	) name9518 (
		_w19935_,
		_w19936_,
		_w20030_
	);
	LUT2 #(
		.INIT('h8)
	) name9519 (
		_w19933_,
		_w19934_,
		_w20031_
	);
	LUT2 #(
		.INIT('h8)
	) name9520 (
		_w19931_,
		_w19932_,
		_w20032_
	);
	LUT2 #(
		.INIT('h8)
	) name9521 (
		_w19929_,
		_w19930_,
		_w20033_
	);
	LUT2 #(
		.INIT('h8)
	) name9522 (
		_w19927_,
		_w19928_,
		_w20034_
	);
	LUT2 #(
		.INIT('h8)
	) name9523 (
		_w19925_,
		_w19926_,
		_w20035_
	);
	LUT2 #(
		.INIT('h8)
	) name9524 (
		_w19923_,
		_w19924_,
		_w20036_
	);
	LUT2 #(
		.INIT('h8)
	) name9525 (
		_w19921_,
		_w19922_,
		_w20037_
	);
	LUT2 #(
		.INIT('h8)
	) name9526 (
		_w19919_,
		_w19920_,
		_w20038_
	);
	LUT2 #(
		.INIT('h8)
	) name9527 (
		_w19917_,
		_w19918_,
		_w20039_
	);
	LUT2 #(
		.INIT('h8)
	) name9528 (
		_w19915_,
		_w19916_,
		_w20040_
	);
	LUT2 #(
		.INIT('h8)
	) name9529 (
		_w19913_,
		_w19914_,
		_w20041_
	);
	LUT2 #(
		.INIT('h8)
	) name9530 (
		_w19911_,
		_w19912_,
		_w20042_
	);
	LUT2 #(
		.INIT('h8)
	) name9531 (
		_w19909_,
		_w19910_,
		_w20043_
	);
	LUT2 #(
		.INIT('h8)
	) name9532 (
		_w19907_,
		_w19908_,
		_w20044_
	);
	LUT2 #(
		.INIT('h8)
	) name9533 (
		_w19905_,
		_w19906_,
		_w20045_
	);
	LUT2 #(
		.INIT('h8)
	) name9534 (
		_w19903_,
		_w19904_,
		_w20046_
	);
	LUT2 #(
		.INIT('h8)
	) name9535 (
		_w19901_,
		_w19902_,
		_w20047_
	);
	LUT2 #(
		.INIT('h8)
	) name9536 (
		_w19899_,
		_w19900_,
		_w20048_
	);
	LUT2 #(
		.INIT('h8)
	) name9537 (
		_w19897_,
		_w19898_,
		_w20049_
	);
	LUT2 #(
		.INIT('h8)
	) name9538 (
		_w19895_,
		_w19896_,
		_w20050_
	);
	LUT2 #(
		.INIT('h8)
	) name9539 (
		_w19893_,
		_w19894_,
		_w20051_
	);
	LUT2 #(
		.INIT('h8)
	) name9540 (
		_w19891_,
		_w19892_,
		_w20052_
	);
	LUT2 #(
		.INIT('h8)
	) name9541 (
		_w19889_,
		_w19890_,
		_w20053_
	);
	LUT2 #(
		.INIT('h8)
	) name9542 (
		_w19887_,
		_w19888_,
		_w20054_
	);
	LUT2 #(
		.INIT('h8)
	) name9543 (
		_w19885_,
		_w19886_,
		_w20055_
	);
	LUT2 #(
		.INIT('h8)
	) name9544 (
		_w19883_,
		_w19884_,
		_w20056_
	);
	LUT2 #(
		.INIT('h8)
	) name9545 (
		_w19881_,
		_w19882_,
		_w20057_
	);
	LUT2 #(
		.INIT('h8)
	) name9546 (
		_w19879_,
		_w19880_,
		_w20058_
	);
	LUT2 #(
		.INIT('h8)
	) name9547 (
		_w19877_,
		_w19878_,
		_w20059_
	);
	LUT2 #(
		.INIT('h8)
	) name9548 (
		_w19875_,
		_w19876_,
		_w20060_
	);
	LUT2 #(
		.INIT('h8)
	) name9549 (
		_w19873_,
		_w19874_,
		_w20061_
	);
	LUT2 #(
		.INIT('h8)
	) name9550 (
		_w19871_,
		_w19872_,
		_w20062_
	);
	LUT2 #(
		.INIT('h8)
	) name9551 (
		_w20061_,
		_w20062_,
		_w20063_
	);
	LUT2 #(
		.INIT('h8)
	) name9552 (
		_w20059_,
		_w20060_,
		_w20064_
	);
	LUT2 #(
		.INIT('h8)
	) name9553 (
		_w20057_,
		_w20058_,
		_w20065_
	);
	LUT2 #(
		.INIT('h8)
	) name9554 (
		_w20055_,
		_w20056_,
		_w20066_
	);
	LUT2 #(
		.INIT('h8)
	) name9555 (
		_w20053_,
		_w20054_,
		_w20067_
	);
	LUT2 #(
		.INIT('h8)
	) name9556 (
		_w20051_,
		_w20052_,
		_w20068_
	);
	LUT2 #(
		.INIT('h8)
	) name9557 (
		_w20049_,
		_w20050_,
		_w20069_
	);
	LUT2 #(
		.INIT('h8)
	) name9558 (
		_w20047_,
		_w20048_,
		_w20070_
	);
	LUT2 #(
		.INIT('h8)
	) name9559 (
		_w20045_,
		_w20046_,
		_w20071_
	);
	LUT2 #(
		.INIT('h8)
	) name9560 (
		_w20043_,
		_w20044_,
		_w20072_
	);
	LUT2 #(
		.INIT('h8)
	) name9561 (
		_w20041_,
		_w20042_,
		_w20073_
	);
	LUT2 #(
		.INIT('h8)
	) name9562 (
		_w20039_,
		_w20040_,
		_w20074_
	);
	LUT2 #(
		.INIT('h8)
	) name9563 (
		_w20037_,
		_w20038_,
		_w20075_
	);
	LUT2 #(
		.INIT('h8)
	) name9564 (
		_w20035_,
		_w20036_,
		_w20076_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		_w20033_,
		_w20034_,
		_w20077_
	);
	LUT2 #(
		.INIT('h8)
	) name9566 (
		_w20031_,
		_w20032_,
		_w20078_
	);
	LUT2 #(
		.INIT('h8)
	) name9567 (
		_w20029_,
		_w20030_,
		_w20079_
	);
	LUT2 #(
		.INIT('h8)
	) name9568 (
		_w20027_,
		_w20028_,
		_w20080_
	);
	LUT2 #(
		.INIT('h8)
	) name9569 (
		_w20025_,
		_w20026_,
		_w20081_
	);
	LUT2 #(
		.INIT('h8)
	) name9570 (
		_w20023_,
		_w20024_,
		_w20082_
	);
	LUT2 #(
		.INIT('h8)
	) name9571 (
		_w20021_,
		_w20022_,
		_w20083_
	);
	LUT2 #(
		.INIT('h8)
	) name9572 (
		_w20019_,
		_w20020_,
		_w20084_
	);
	LUT2 #(
		.INIT('h8)
	) name9573 (
		_w20017_,
		_w20018_,
		_w20085_
	);
	LUT2 #(
		.INIT('h8)
	) name9574 (
		_w20015_,
		_w20016_,
		_w20086_
	);
	LUT2 #(
		.INIT('h8)
	) name9575 (
		_w20013_,
		_w20014_,
		_w20087_
	);
	LUT2 #(
		.INIT('h8)
	) name9576 (
		_w20011_,
		_w20012_,
		_w20088_
	);
	LUT2 #(
		.INIT('h8)
	) name9577 (
		_w20009_,
		_w20010_,
		_w20089_
	);
	LUT2 #(
		.INIT('h8)
	) name9578 (
		_w20007_,
		_w20008_,
		_w20090_
	);
	LUT2 #(
		.INIT('h8)
	) name9579 (
		_w20005_,
		_w20006_,
		_w20091_
	);
	LUT2 #(
		.INIT('h8)
	) name9580 (
		_w20003_,
		_w20004_,
		_w20092_
	);
	LUT2 #(
		.INIT('h8)
	) name9581 (
		_w20001_,
		_w20002_,
		_w20093_
	);
	LUT2 #(
		.INIT('h8)
	) name9582 (
		_w19999_,
		_w20000_,
		_w20094_
	);
	LUT2 #(
		.INIT('h8)
	) name9583 (
		_w20093_,
		_w20094_,
		_w20095_
	);
	LUT2 #(
		.INIT('h8)
	) name9584 (
		_w20091_,
		_w20092_,
		_w20096_
	);
	LUT2 #(
		.INIT('h8)
	) name9585 (
		_w20089_,
		_w20090_,
		_w20097_
	);
	LUT2 #(
		.INIT('h8)
	) name9586 (
		_w20087_,
		_w20088_,
		_w20098_
	);
	LUT2 #(
		.INIT('h8)
	) name9587 (
		_w20085_,
		_w20086_,
		_w20099_
	);
	LUT2 #(
		.INIT('h8)
	) name9588 (
		_w20083_,
		_w20084_,
		_w20100_
	);
	LUT2 #(
		.INIT('h8)
	) name9589 (
		_w20081_,
		_w20082_,
		_w20101_
	);
	LUT2 #(
		.INIT('h8)
	) name9590 (
		_w20079_,
		_w20080_,
		_w20102_
	);
	LUT2 #(
		.INIT('h8)
	) name9591 (
		_w20077_,
		_w20078_,
		_w20103_
	);
	LUT2 #(
		.INIT('h8)
	) name9592 (
		_w20075_,
		_w20076_,
		_w20104_
	);
	LUT2 #(
		.INIT('h8)
	) name9593 (
		_w20073_,
		_w20074_,
		_w20105_
	);
	LUT2 #(
		.INIT('h8)
	) name9594 (
		_w20071_,
		_w20072_,
		_w20106_
	);
	LUT2 #(
		.INIT('h8)
	) name9595 (
		_w20069_,
		_w20070_,
		_w20107_
	);
	LUT2 #(
		.INIT('h8)
	) name9596 (
		_w20067_,
		_w20068_,
		_w20108_
	);
	LUT2 #(
		.INIT('h8)
	) name9597 (
		_w20065_,
		_w20066_,
		_w20109_
	);
	LUT2 #(
		.INIT('h8)
	) name9598 (
		_w20063_,
		_w20064_,
		_w20110_
	);
	LUT2 #(
		.INIT('h8)
	) name9599 (
		_w20109_,
		_w20110_,
		_w20111_
	);
	LUT2 #(
		.INIT('h8)
	) name9600 (
		_w20107_,
		_w20108_,
		_w20112_
	);
	LUT2 #(
		.INIT('h8)
	) name9601 (
		_w20105_,
		_w20106_,
		_w20113_
	);
	LUT2 #(
		.INIT('h8)
	) name9602 (
		_w20103_,
		_w20104_,
		_w20114_
	);
	LUT2 #(
		.INIT('h8)
	) name9603 (
		_w20101_,
		_w20102_,
		_w20115_
	);
	LUT2 #(
		.INIT('h8)
	) name9604 (
		_w20099_,
		_w20100_,
		_w20116_
	);
	LUT2 #(
		.INIT('h8)
	) name9605 (
		_w20097_,
		_w20098_,
		_w20117_
	);
	LUT2 #(
		.INIT('h8)
	) name9606 (
		_w20095_,
		_w20096_,
		_w20118_
	);
	LUT2 #(
		.INIT('h8)
	) name9607 (
		_w20117_,
		_w20118_,
		_w20119_
	);
	LUT2 #(
		.INIT('h8)
	) name9608 (
		_w20115_,
		_w20116_,
		_w20120_
	);
	LUT2 #(
		.INIT('h8)
	) name9609 (
		_w20113_,
		_w20114_,
		_w20121_
	);
	LUT2 #(
		.INIT('h8)
	) name9610 (
		_w20111_,
		_w20112_,
		_w20122_
	);
	LUT2 #(
		.INIT('h8)
	) name9611 (
		_w20121_,
		_w20122_,
		_w20123_
	);
	LUT2 #(
		.INIT('h8)
	) name9612 (
		_w20119_,
		_w20120_,
		_w20124_
	);
	LUT2 #(
		.INIT('h8)
	) name9613 (
		_w20123_,
		_w20124_,
		_w20125_
	);
	LUT2 #(
		.INIT('h1)
	) name9614 (
		wb_rst_i_pad,
		_w20125_,
		_w20126_
	);
	LUT2 #(
		.INIT('h8)
	) name9615 (
		_w12656_,
		_w20126_,
		_w20127_
	);
	LUT2 #(
		.INIT('h8)
	) name9616 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w12658_,
		_w20128_
	);
	LUT2 #(
		.INIT('h1)
	) name9617 (
		_w19614_,
		_w20128_,
		_w20129_
	);
	LUT2 #(
		.INIT('h4)
	) name9618 (
		_w20127_,
		_w20129_,
		_w20130_
	);
	LUT2 #(
		.INIT('h1)
	) name9619 (
		\txethmac1_txcounters1_ByteCnt_reg[11]/NET0131 ,
		_w14577_,
		_w20131_
	);
	LUT2 #(
		.INIT('h4)
	) name9620 (
		_w14578_,
		_w14582_,
		_w20132_
	);
	LUT2 #(
		.INIT('h4)
	) name9621 (
		_w20131_,
		_w20132_,
		_w20133_
	);
	LUT2 #(
		.INIT('h2)
	) name9622 (
		\txethmac1_txcrc_Crc_reg[5]/NET0131 ,
		_w11422_,
		_w20134_
	);
	LUT2 #(
		.INIT('h4)
	) name9623 (
		\txethmac1_txcrc_Crc_reg[5]/NET0131 ,
		_w11422_,
		_w20135_
	);
	LUT2 #(
		.INIT('h2)
	) name9624 (
		_w11181_,
		_w20134_,
		_w20136_
	);
	LUT2 #(
		.INIT('h4)
	) name9625 (
		_w20135_,
		_w20136_,
		_w20137_
	);
	LUT2 #(
		.INIT('h8)
	) name9626 (
		\m_wb_adr_o[12]_pad ,
		_w12636_,
		_w20138_
	);
	LUT2 #(
		.INIT('h1)
	) name9627 (
		\m_wb_adr_o[12]_pad ,
		_w12587_,
		_w20139_
	);
	LUT2 #(
		.INIT('h4)
	) name9628 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w12608_,
		_w20140_
	);
	LUT2 #(
		.INIT('h2)
	) name9629 (
		_w12621_,
		_w20140_,
		_w20141_
	);
	LUT2 #(
		.INIT('h1)
	) name9630 (
		_w12623_,
		_w20141_,
		_w20142_
	);
	LUT2 #(
		.INIT('h1)
	) name9631 (
		_w12588_,
		_w20142_,
		_w20143_
	);
	LUT2 #(
		.INIT('h4)
	) name9632 (
		_w20139_,
		_w20143_,
		_w20144_
	);
	LUT2 #(
		.INIT('h8)
	) name9633 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w12634_,
		_w20145_
	);
	LUT2 #(
		.INIT('h8)
	) name9634 (
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w12577_,
		_w20146_
	);
	LUT2 #(
		.INIT('h1)
	) name9635 (
		_w20138_,
		_w20145_,
		_w20147_
	);
	LUT2 #(
		.INIT('h4)
	) name9636 (
		_w20146_,
		_w20147_,
		_w20148_
	);
	LUT2 #(
		.INIT('h4)
	) name9637 (
		_w20144_,
		_w20148_,
		_w20149_
	);
	LUT2 #(
		.INIT('h8)
	) name9638 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w12577_,
		_w20150_
	);
	LUT2 #(
		.INIT('h1)
	) name9639 (
		\m_wb_adr_o[16]_pad ,
		_w12591_,
		_w20151_
	);
	LUT2 #(
		.INIT('h4)
	) name9640 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w12575_,
		_w20152_
	);
	LUT2 #(
		.INIT('h2)
	) name9641 (
		_w12561_,
		_w20152_,
		_w20153_
	);
	LUT2 #(
		.INIT('h1)
	) name9642 (
		_w14590_,
		_w20153_,
		_w20154_
	);
	LUT2 #(
		.INIT('h1)
	) name9643 (
		_w12592_,
		_w20154_,
		_w20155_
	);
	LUT2 #(
		.INIT('h4)
	) name9644 (
		_w20151_,
		_w20155_,
		_w20156_
	);
	LUT2 #(
		.INIT('h8)
	) name9645 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w12634_,
		_w20157_
	);
	LUT2 #(
		.INIT('h8)
	) name9646 (
		\m_wb_adr_o[16]_pad ,
		_w12636_,
		_w20158_
	);
	LUT2 #(
		.INIT('h1)
	) name9647 (
		_w20150_,
		_w20157_,
		_w20159_
	);
	LUT2 #(
		.INIT('h4)
	) name9648 (
		_w20158_,
		_w20159_,
		_w20160_
	);
	LUT2 #(
		.INIT('h4)
	) name9649 (
		_w20156_,
		_w20160_,
		_w20161_
	);
	LUT2 #(
		.INIT('h8)
	) name9650 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w12577_,
		_w20162_
	);
	LUT2 #(
		.INIT('h1)
	) name9651 (
		\m_wb_adr_o[17]_pad ,
		_w12592_,
		_w20163_
	);
	LUT2 #(
		.INIT('h4)
	) name9652 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w12575_,
		_w20164_
	);
	LUT2 #(
		.INIT('h2)
	) name9653 (
		_w12561_,
		_w20164_,
		_w20165_
	);
	LUT2 #(
		.INIT('h1)
	) name9654 (
		_w14590_,
		_w20165_,
		_w20166_
	);
	LUT2 #(
		.INIT('h1)
	) name9655 (
		_w16223_,
		_w20166_,
		_w20167_
	);
	LUT2 #(
		.INIT('h4)
	) name9656 (
		_w20163_,
		_w20167_,
		_w20168_
	);
	LUT2 #(
		.INIT('h8)
	) name9657 (
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w12634_,
		_w20169_
	);
	LUT2 #(
		.INIT('h8)
	) name9658 (
		\m_wb_adr_o[17]_pad ,
		_w12636_,
		_w20170_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		_w20162_,
		_w20169_,
		_w20171_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w20170_,
		_w20171_,
		_w20172_
	);
	LUT2 #(
		.INIT('h4)
	) name9661 (
		_w20168_,
		_w20172_,
		_w20173_
	);
	LUT2 #(
		.INIT('h8)
	) name9662 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w12577_,
		_w20174_
	);
	LUT2 #(
		.INIT('h1)
	) name9663 (
		\m_wb_adr_o[19]_pad ,
		_w12594_,
		_w20175_
	);
	LUT2 #(
		.INIT('h4)
	) name9664 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w12575_,
		_w20176_
	);
	LUT2 #(
		.INIT('h2)
	) name9665 (
		_w12561_,
		_w20176_,
		_w20177_
	);
	LUT2 #(
		.INIT('h1)
	) name9666 (
		_w14590_,
		_w20177_,
		_w20178_
	);
	LUT2 #(
		.INIT('h1)
	) name9667 (
		_w12595_,
		_w20178_,
		_w20179_
	);
	LUT2 #(
		.INIT('h4)
	) name9668 (
		_w20175_,
		_w20179_,
		_w20180_
	);
	LUT2 #(
		.INIT('h8)
	) name9669 (
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w12634_,
		_w20181_
	);
	LUT2 #(
		.INIT('h8)
	) name9670 (
		\m_wb_adr_o[19]_pad ,
		_w12636_,
		_w20182_
	);
	LUT2 #(
		.INIT('h1)
	) name9671 (
		_w20174_,
		_w20181_,
		_w20183_
	);
	LUT2 #(
		.INIT('h4)
	) name9672 (
		_w20182_,
		_w20183_,
		_w20184_
	);
	LUT2 #(
		.INIT('h4)
	) name9673 (
		_w20180_,
		_w20184_,
		_w20185_
	);
	LUT2 #(
		.INIT('h8)
	) name9674 (
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w12577_,
		_w20186_
	);
	LUT2 #(
		.INIT('h1)
	) name9675 (
		\m_wb_adr_o[20]_pad ,
		_w12595_,
		_w20187_
	);
	LUT2 #(
		.INIT('h4)
	) name9676 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w12608_,
		_w20188_
	);
	LUT2 #(
		.INIT('h2)
	) name9677 (
		_w12621_,
		_w20188_,
		_w20189_
	);
	LUT2 #(
		.INIT('h1)
	) name9678 (
		_w12623_,
		_w20189_,
		_w20190_
	);
	LUT2 #(
		.INIT('h1)
	) name9679 (
		_w12596_,
		_w20190_,
		_w20191_
	);
	LUT2 #(
		.INIT('h4)
	) name9680 (
		_w20187_,
		_w20191_,
		_w20192_
	);
	LUT2 #(
		.INIT('h8)
	) name9681 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w12634_,
		_w20193_
	);
	LUT2 #(
		.INIT('h8)
	) name9682 (
		\m_wb_adr_o[20]_pad ,
		_w12636_,
		_w20194_
	);
	LUT2 #(
		.INIT('h1)
	) name9683 (
		_w20186_,
		_w20193_,
		_w20195_
	);
	LUT2 #(
		.INIT('h4)
	) name9684 (
		_w20194_,
		_w20195_,
		_w20196_
	);
	LUT2 #(
		.INIT('h4)
	) name9685 (
		_w20192_,
		_w20196_,
		_w20197_
	);
	LUT2 #(
		.INIT('h8)
	) name9686 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w12577_,
		_w20198_
	);
	LUT2 #(
		.INIT('h1)
	) name9687 (
		\m_wb_adr_o[21]_pad ,
		_w12596_,
		_w20199_
	);
	LUT2 #(
		.INIT('h4)
	) name9688 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w12575_,
		_w20200_
	);
	LUT2 #(
		.INIT('h2)
	) name9689 (
		_w12561_,
		_w20200_,
		_w20201_
	);
	LUT2 #(
		.INIT('h1)
	) name9690 (
		_w14590_,
		_w20201_,
		_w20202_
	);
	LUT2 #(
		.INIT('h1)
	) name9691 (
		_w12597_,
		_w20202_,
		_w20203_
	);
	LUT2 #(
		.INIT('h4)
	) name9692 (
		_w20199_,
		_w20203_,
		_w20204_
	);
	LUT2 #(
		.INIT('h8)
	) name9693 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		_w12634_,
		_w20205_
	);
	LUT2 #(
		.INIT('h8)
	) name9694 (
		\m_wb_adr_o[21]_pad ,
		_w12636_,
		_w20206_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		_w20198_,
		_w20205_,
		_w20207_
	);
	LUT2 #(
		.INIT('h4)
	) name9696 (
		_w20206_,
		_w20207_,
		_w20208_
	);
	LUT2 #(
		.INIT('h4)
	) name9697 (
		_w20204_,
		_w20208_,
		_w20209_
	);
	LUT2 #(
		.INIT('h8)
	) name9698 (
		\m_wb_adr_o[3]_pad ,
		_w12636_,
		_w20210_
	);
	LUT2 #(
		.INIT('h8)
	) name9699 (
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w12577_,
		_w20211_
	);
	LUT2 #(
		.INIT('h8)
	) name9700 (
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w12634_,
		_w20212_
	);
	LUT2 #(
		.INIT('h1)
	) name9701 (
		\m_wb_adr_o[2]_pad ,
		\m_wb_adr_o[3]_pad ,
		_w20213_
	);
	LUT2 #(
		.INIT('h1)
	) name9702 (
		_w12579_,
		_w20213_,
		_w20214_
	);
	LUT2 #(
		.INIT('h4)
	) name9703 (
		_w14591_,
		_w20214_,
		_w20215_
	);
	LUT2 #(
		.INIT('h1)
	) name9704 (
		_w20210_,
		_w20212_,
		_w20216_
	);
	LUT2 #(
		.INIT('h1)
	) name9705 (
		_w20211_,
		_w20215_,
		_w20217_
	);
	LUT2 #(
		.INIT('h8)
	) name9706 (
		_w20216_,
		_w20217_,
		_w20218_
	);
	LUT2 #(
		.INIT('h8)
	) name9707 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w12577_,
		_w20219_
	);
	LUT2 #(
		.INIT('h1)
	) name9708 (
		\m_wb_adr_o[22]_pad ,
		_w12597_,
		_w20220_
	);
	LUT2 #(
		.INIT('h4)
	) name9709 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w12575_,
		_w20221_
	);
	LUT2 #(
		.INIT('h2)
	) name9710 (
		_w12561_,
		_w20221_,
		_w20222_
	);
	LUT2 #(
		.INIT('h1)
	) name9711 (
		_w14590_,
		_w20222_,
		_w20223_
	);
	LUT2 #(
		.INIT('h8)
	) name9712 (
		\m_wb_adr_o[22]_pad ,
		_w12597_,
		_w20224_
	);
	LUT2 #(
		.INIT('h1)
	) name9713 (
		_w20220_,
		_w20223_,
		_w20225_
	);
	LUT2 #(
		.INIT('h4)
	) name9714 (
		_w20224_,
		_w20225_,
		_w20226_
	);
	LUT2 #(
		.INIT('h8)
	) name9715 (
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w12634_,
		_w20227_
	);
	LUT2 #(
		.INIT('h8)
	) name9716 (
		\m_wb_adr_o[22]_pad ,
		_w12636_,
		_w20228_
	);
	LUT2 #(
		.INIT('h1)
	) name9717 (
		_w20219_,
		_w20227_,
		_w20229_
	);
	LUT2 #(
		.INIT('h4)
	) name9718 (
		_w20228_,
		_w20229_,
		_w20230_
	);
	LUT2 #(
		.INIT('h4)
	) name9719 (
		_w20226_,
		_w20230_,
		_w20231_
	);
	LUT2 #(
		.INIT('h8)
	) name9720 (
		\m_wb_adr_o[23]_pad ,
		_w12636_,
		_w20232_
	);
	LUT2 #(
		.INIT('h1)
	) name9721 (
		\m_wb_adr_o[23]_pad ,
		_w20224_,
		_w20233_
	);
	LUT2 #(
		.INIT('h8)
	) name9722 (
		\m_wb_adr_o[23]_pad ,
		_w20224_,
		_w20234_
	);
	LUT2 #(
		.INIT('h1)
	) name9723 (
		_w14591_,
		_w20233_,
		_w20235_
	);
	LUT2 #(
		.INIT('h4)
	) name9724 (
		_w20234_,
		_w20235_,
		_w20236_
	);
	LUT2 #(
		.INIT('h8)
	) name9725 (
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w12634_,
		_w20237_
	);
	LUT2 #(
		.INIT('h8)
	) name9726 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		_w12577_,
		_w20238_
	);
	LUT2 #(
		.INIT('h1)
	) name9727 (
		_w20232_,
		_w20237_,
		_w20239_
	);
	LUT2 #(
		.INIT('h4)
	) name9728 (
		_w20238_,
		_w20239_,
		_w20240_
	);
	LUT2 #(
		.INIT('h4)
	) name9729 (
		_w20236_,
		_w20240_,
		_w20241_
	);
	LUT2 #(
		.INIT('h8)
	) name9730 (
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w12577_,
		_w20242_
	);
	LUT2 #(
		.INIT('h4)
	) name9731 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w12608_,
		_w20243_
	);
	LUT2 #(
		.INIT('h2)
	) name9732 (
		_w12621_,
		_w20243_,
		_w20244_
	);
	LUT2 #(
		.INIT('h1)
	) name9733 (
		_w12623_,
		_w20244_,
		_w20245_
	);
	LUT2 #(
		.INIT('h1)
	) name9734 (
		\m_wb_adr_o[24]_pad ,
		_w20234_,
		_w20246_
	);
	LUT2 #(
		.INIT('h1)
	) name9735 (
		_w15125_,
		_w20245_,
		_w20247_
	);
	LUT2 #(
		.INIT('h4)
	) name9736 (
		_w20246_,
		_w20247_,
		_w20248_
	);
	LUT2 #(
		.INIT('h8)
	) name9737 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w12634_,
		_w20249_
	);
	LUT2 #(
		.INIT('h8)
	) name9738 (
		\m_wb_adr_o[24]_pad ,
		_w12636_,
		_w20250_
	);
	LUT2 #(
		.INIT('h1)
	) name9739 (
		_w20242_,
		_w20249_,
		_w20251_
	);
	LUT2 #(
		.INIT('h4)
	) name9740 (
		_w20250_,
		_w20251_,
		_w20252_
	);
	LUT2 #(
		.INIT('h4)
	) name9741 (
		_w20248_,
		_w20252_,
		_w20253_
	);
	LUT2 #(
		.INIT('h4)
	) name9742 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w12575_,
		_w20254_
	);
	LUT2 #(
		.INIT('h1)
	) name9743 (
		\m_wb_adr_o[25]_pad ,
		_w15125_,
		_w20255_
	);
	LUT2 #(
		.INIT('h1)
	) name9744 (
		_w15126_,
		_w20255_,
		_w20256_
	);
	LUT2 #(
		.INIT('h1)
	) name9745 (
		_w12575_,
		_w20256_,
		_w20257_
	);
	LUT2 #(
		.INIT('h2)
	) name9746 (
		_w12561_,
		_w20254_,
		_w20258_
	);
	LUT2 #(
		.INIT('h4)
	) name9747 (
		_w20257_,
		_w20258_,
		_w20259_
	);
	LUT2 #(
		.INIT('h8)
	) name9748 (
		\m_wb_adr_o[25]_pad ,
		_w12636_,
		_w20260_
	);
	LUT2 #(
		.INIT('h8)
	) name9749 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		_w12631_,
		_w20261_
	);
	LUT2 #(
		.INIT('h8)
	) name9750 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w12572_,
		_w20262_
	);
	LUT2 #(
		.INIT('h4)
	) name9751 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		_w12608_,
		_w20263_
	);
	LUT2 #(
		.INIT('h1)
	) name9752 (
		_w12608_,
		_w20256_,
		_w20264_
	);
	LUT2 #(
		.INIT('h2)
	) name9753 (
		_w12621_,
		_w20263_,
		_w20265_
	);
	LUT2 #(
		.INIT('h4)
	) name9754 (
		_w20264_,
		_w20265_,
		_w20266_
	);
	LUT2 #(
		.INIT('h1)
	) name9755 (
		_w20261_,
		_w20262_,
		_w20267_
	);
	LUT2 #(
		.INIT('h4)
	) name9756 (
		_w20260_,
		_w20267_,
		_w20268_
	);
	LUT2 #(
		.INIT('h4)
	) name9757 (
		_w20259_,
		_w20268_,
		_w20269_
	);
	LUT2 #(
		.INIT('h4)
	) name9758 (
		_w20266_,
		_w20269_,
		_w20270_
	);
	LUT2 #(
		.INIT('h8)
	) name9759 (
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w12577_,
		_w20271_
	);
	LUT2 #(
		.INIT('h4)
	) name9760 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w12608_,
		_w20272_
	);
	LUT2 #(
		.INIT('h2)
	) name9761 (
		_w12621_,
		_w20272_,
		_w20273_
	);
	LUT2 #(
		.INIT('h1)
	) name9762 (
		_w12623_,
		_w20273_,
		_w20274_
	);
	LUT2 #(
		.INIT('h1)
	) name9763 (
		\m_wb_adr_o[28]_pad ,
		_w18019_,
		_w20275_
	);
	LUT2 #(
		.INIT('h1)
	) name9764 (
		_w12604_,
		_w20274_,
		_w20276_
	);
	LUT2 #(
		.INIT('h4)
	) name9765 (
		_w20275_,
		_w20276_,
		_w20277_
	);
	LUT2 #(
		.INIT('h8)
	) name9766 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w12634_,
		_w20278_
	);
	LUT2 #(
		.INIT('h8)
	) name9767 (
		\m_wb_adr_o[28]_pad ,
		_w12636_,
		_w20279_
	);
	LUT2 #(
		.INIT('h1)
	) name9768 (
		_w20271_,
		_w20278_,
		_w20280_
	);
	LUT2 #(
		.INIT('h4)
	) name9769 (
		_w20279_,
		_w20280_,
		_w20281_
	);
	LUT2 #(
		.INIT('h4)
	) name9770 (
		_w20277_,
		_w20281_,
		_w20282_
	);
	LUT2 #(
		.INIT('h8)
	) name9771 (
		\m_wb_adr_o[29]_pad ,
		_w12636_,
		_w20283_
	);
	LUT2 #(
		.INIT('h1)
	) name9772 (
		\m_wb_adr_o[29]_pad ,
		_w12604_,
		_w20284_
	);
	LUT2 #(
		.INIT('h4)
	) name9773 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w12608_,
		_w20285_
	);
	LUT2 #(
		.INIT('h2)
	) name9774 (
		_w12621_,
		_w20285_,
		_w20286_
	);
	LUT2 #(
		.INIT('h1)
	) name9775 (
		_w12623_,
		_w20286_,
		_w20287_
	);
	LUT2 #(
		.INIT('h1)
	) name9776 (
		_w12605_,
		_w20287_,
		_w20288_
	);
	LUT2 #(
		.INIT('h4)
	) name9777 (
		_w20284_,
		_w20288_,
		_w20289_
	);
	LUT2 #(
		.INIT('h8)
	) name9778 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w12634_,
		_w20290_
	);
	LUT2 #(
		.INIT('h8)
	) name9779 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		_w12577_,
		_w20291_
	);
	LUT2 #(
		.INIT('h1)
	) name9780 (
		_w20283_,
		_w20290_,
		_w20292_
	);
	LUT2 #(
		.INIT('h4)
	) name9781 (
		_w20291_,
		_w20292_,
		_w20293_
	);
	LUT2 #(
		.INIT('h4)
	) name9782 (
		_w20289_,
		_w20293_,
		_w20294_
	);
	LUT2 #(
		.INIT('h8)
	) name9783 (
		\m_wb_adr_o[5]_pad ,
		_w12636_,
		_w20295_
	);
	LUT2 #(
		.INIT('h8)
	) name9784 (
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w12577_,
		_w20296_
	);
	LUT2 #(
		.INIT('h8)
	) name9785 (
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w12634_,
		_w20297_
	);
	LUT2 #(
		.INIT('h1)
	) name9786 (
		\m_wb_adr_o[5]_pad ,
		_w12580_,
		_w20298_
	);
	LUT2 #(
		.INIT('h1)
	) name9787 (
		_w12581_,
		_w20298_,
		_w20299_
	);
	LUT2 #(
		.INIT('h4)
	) name9788 (
		_w14591_,
		_w20299_,
		_w20300_
	);
	LUT2 #(
		.INIT('h1)
	) name9789 (
		_w20295_,
		_w20297_,
		_w20301_
	);
	LUT2 #(
		.INIT('h1)
	) name9790 (
		_w20296_,
		_w20300_,
		_w20302_
	);
	LUT2 #(
		.INIT('h8)
	) name9791 (
		_w20301_,
		_w20302_,
		_w20303_
	);
	LUT2 #(
		.INIT('h8)
	) name9792 (
		\m_wb_adr_o[6]_pad ,
		_w12636_,
		_w20304_
	);
	LUT2 #(
		.INIT('h8)
	) name9793 (
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w12577_,
		_w20305_
	);
	LUT2 #(
		.INIT('h8)
	) name9794 (
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w12634_,
		_w20306_
	);
	LUT2 #(
		.INIT('h1)
	) name9795 (
		\m_wb_adr_o[6]_pad ,
		_w12581_,
		_w20307_
	);
	LUT2 #(
		.INIT('h1)
	) name9796 (
		_w12582_,
		_w20307_,
		_w20308_
	);
	LUT2 #(
		.INIT('h4)
	) name9797 (
		_w14591_,
		_w20308_,
		_w20309_
	);
	LUT2 #(
		.INIT('h1)
	) name9798 (
		_w20304_,
		_w20306_,
		_w20310_
	);
	LUT2 #(
		.INIT('h1)
	) name9799 (
		_w20305_,
		_w20309_,
		_w20311_
	);
	LUT2 #(
		.INIT('h8)
	) name9800 (
		_w20310_,
		_w20311_,
		_w20312_
	);
	LUT2 #(
		.INIT('h8)
	) name9801 (
		\m_wb_adr_o[7]_pad ,
		_w12636_,
		_w20313_
	);
	LUT2 #(
		.INIT('h8)
	) name9802 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		_w12577_,
		_w20314_
	);
	LUT2 #(
		.INIT('h8)
	) name9803 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		_w12634_,
		_w20315_
	);
	LUT2 #(
		.INIT('h1)
	) name9804 (
		\m_wb_adr_o[7]_pad ,
		_w12582_,
		_w20316_
	);
	LUT2 #(
		.INIT('h1)
	) name9805 (
		_w12583_,
		_w20316_,
		_w20317_
	);
	LUT2 #(
		.INIT('h4)
	) name9806 (
		_w14591_,
		_w20317_,
		_w20318_
	);
	LUT2 #(
		.INIT('h1)
	) name9807 (
		_w20313_,
		_w20315_,
		_w20319_
	);
	LUT2 #(
		.INIT('h1)
	) name9808 (
		_w20314_,
		_w20318_,
		_w20320_
	);
	LUT2 #(
		.INIT('h8)
	) name9809 (
		_w20319_,
		_w20320_,
		_w20321_
	);
	LUT2 #(
		.INIT('h8)
	) name9810 (
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w12577_,
		_w20322_
	);
	LUT2 #(
		.INIT('h8)
	) name9811 (
		\m_wb_adr_o[9]_pad ,
		_w12636_,
		_w20323_
	);
	LUT2 #(
		.INIT('h8)
	) name9812 (
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w12634_,
		_w20324_
	);
	LUT2 #(
		.INIT('h1)
	) name9813 (
		\m_wb_adr_o[9]_pad ,
		_w12584_,
		_w20325_
	);
	LUT2 #(
		.INIT('h1)
	) name9814 (
		_w12585_,
		_w20325_,
		_w20326_
	);
	LUT2 #(
		.INIT('h4)
	) name9815 (
		_w14591_,
		_w20326_,
		_w20327_
	);
	LUT2 #(
		.INIT('h1)
	) name9816 (
		_w20322_,
		_w20324_,
		_w20328_
	);
	LUT2 #(
		.INIT('h1)
	) name9817 (
		_w20323_,
		_w20327_,
		_w20329_
	);
	LUT2 #(
		.INIT('h8)
	) name9818 (
		_w20328_,
		_w20329_,
		_w20330_
	);
	LUT2 #(
		.INIT('h8)
	) name9819 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		_w12577_,
		_w20331_
	);
	LUT2 #(
		.INIT('h8)
	) name9820 (
		\m_wb_adr_o[10]_pad ,
		_w12636_,
		_w20332_
	);
	LUT2 #(
		.INIT('h8)
	) name9821 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		_w12634_,
		_w20333_
	);
	LUT2 #(
		.INIT('h1)
	) name9822 (
		\m_wb_adr_o[10]_pad ,
		_w12585_,
		_w20334_
	);
	LUT2 #(
		.INIT('h1)
	) name9823 (
		_w12586_,
		_w20334_,
		_w20335_
	);
	LUT2 #(
		.INIT('h4)
	) name9824 (
		_w14591_,
		_w20335_,
		_w20336_
	);
	LUT2 #(
		.INIT('h1)
	) name9825 (
		_w20331_,
		_w20333_,
		_w20337_
	);
	LUT2 #(
		.INIT('h1)
	) name9826 (
		_w20332_,
		_w20336_,
		_w20338_
	);
	LUT2 #(
		.INIT('h8)
	) name9827 (
		_w20337_,
		_w20338_,
		_w20339_
	);
	LUT2 #(
		.INIT('h2)
	) name9828 (
		\wishbone_LatchedTxLength_reg[0]/NET0131 ,
		_w12656_,
		_w20340_
	);
	LUT2 #(
		.INIT('h1)
	) name9829 (
		_w19089_,
		_w20340_,
		_w20341_
	);
	LUT2 #(
		.INIT('h2)
	) name9830 (
		\wishbone_LatchedTxLength_reg[10]/NET0131 ,
		_w12656_,
		_w20342_
	);
	LUT2 #(
		.INIT('h1)
	) name9831 (
		_w17288_,
		_w20342_,
		_w20343_
	);
	LUT2 #(
		.INIT('h2)
	) name9832 (
		\wishbone_LatchedTxLength_reg[11]/NET0131 ,
		_w12656_,
		_w20344_
	);
	LUT2 #(
		.INIT('h8)
	) name9833 (
		\wishbone_bd_ram_mem3_reg[30][27]/P0001 ,
		_w13104_,
		_w20345_
	);
	LUT2 #(
		.INIT('h8)
	) name9834 (
		\wishbone_bd_ram_mem3_reg[26][27]/P0001 ,
		_w12699_,
		_w20346_
	);
	LUT2 #(
		.INIT('h8)
	) name9835 (
		\wishbone_bd_ram_mem3_reg[24][27]/P0001 ,
		_w13084_,
		_w20347_
	);
	LUT2 #(
		.INIT('h8)
	) name9836 (
		\wishbone_bd_ram_mem3_reg[104][27]/P0001 ,
		_w13148_,
		_w20348_
	);
	LUT2 #(
		.INIT('h8)
	) name9837 (
		\wishbone_bd_ram_mem3_reg[118][27]/P0001 ,
		_w12830_,
		_w20349_
	);
	LUT2 #(
		.INIT('h8)
	) name9838 (
		\wishbone_bd_ram_mem3_reg[203][27]/P0001 ,
		_w13158_,
		_w20350_
	);
	LUT2 #(
		.INIT('h8)
	) name9839 (
		\wishbone_bd_ram_mem3_reg[131][27]/P0001 ,
		_w12852_,
		_w20351_
	);
	LUT2 #(
		.INIT('h8)
	) name9840 (
		\wishbone_bd_ram_mem3_reg[70][27]/P0001 ,
		_w12840_,
		_w20352_
	);
	LUT2 #(
		.INIT('h8)
	) name9841 (
		\wishbone_bd_ram_mem3_reg[103][27]/P0001 ,
		_w12846_,
		_w20353_
	);
	LUT2 #(
		.INIT('h8)
	) name9842 (
		\wishbone_bd_ram_mem3_reg[216][27]/P0001 ,
		_w13028_,
		_w20354_
	);
	LUT2 #(
		.INIT('h8)
	) name9843 (
		\wishbone_bd_ram_mem3_reg[212][27]/P0001 ,
		_w12796_,
		_w20355_
	);
	LUT2 #(
		.INIT('h8)
	) name9844 (
		\wishbone_bd_ram_mem3_reg[155][27]/P0001 ,
		_w13122_,
		_w20356_
	);
	LUT2 #(
		.INIT('h8)
	) name9845 (
		\wishbone_bd_ram_mem3_reg[4][27]/P0001 ,
		_w12666_,
		_w20357_
	);
	LUT2 #(
		.INIT('h8)
	) name9846 (
		\wishbone_bd_ram_mem3_reg[94][27]/P0001 ,
		_w13186_,
		_w20358_
	);
	LUT2 #(
		.INIT('h8)
	) name9847 (
		\wishbone_bd_ram_mem3_reg[77][27]/P0001 ,
		_w12982_,
		_w20359_
	);
	LUT2 #(
		.INIT('h8)
	) name9848 (
		\wishbone_bd_ram_mem3_reg[32][27]/P0001 ,
		_w13120_,
		_w20360_
	);
	LUT2 #(
		.INIT('h8)
	) name9849 (
		\wishbone_bd_ram_mem3_reg[247][27]/P0001 ,
		_w12818_,
		_w20361_
	);
	LUT2 #(
		.INIT('h8)
	) name9850 (
		\wishbone_bd_ram_mem3_reg[232][27]/P0001 ,
		_w12758_,
		_w20362_
	);
	LUT2 #(
		.INIT('h8)
	) name9851 (
		\wishbone_bd_ram_mem3_reg[34][27]/P0001 ,
		_w12930_,
		_w20363_
	);
	LUT2 #(
		.INIT('h8)
	) name9852 (
		\wishbone_bd_ram_mem3_reg[8][27]/P0001 ,
		_w12920_,
		_w20364_
	);
	LUT2 #(
		.INIT('h8)
	) name9853 (
		\wishbone_bd_ram_mem3_reg[160][27]/P0001 ,
		_w12872_,
		_w20365_
	);
	LUT2 #(
		.INIT('h8)
	) name9854 (
		\wishbone_bd_ram_mem3_reg[198][27]/P0001 ,
		_w12832_,
		_w20366_
	);
	LUT2 #(
		.INIT('h8)
	) name9855 (
		\wishbone_bd_ram_mem3_reg[183][27]/P0001 ,
		_w12787_,
		_w20367_
	);
	LUT2 #(
		.INIT('h8)
	) name9856 (
		\wishbone_bd_ram_mem3_reg[121][27]/P0001 ,
		_w13078_,
		_w20368_
	);
	LUT2 #(
		.INIT('h8)
	) name9857 (
		\wishbone_bd_ram_mem3_reg[176][27]/P0001 ,
		_w12868_,
		_w20369_
	);
	LUT2 #(
		.INIT('h8)
	) name9858 (
		\wishbone_bd_ram_mem3_reg[148][27]/P0001 ,
		_w13000_,
		_w20370_
	);
	LUT2 #(
		.INIT('h8)
	) name9859 (
		\wishbone_bd_ram_mem3_reg[96][27]/P0001 ,
		_w12912_,
		_w20371_
	);
	LUT2 #(
		.INIT('h8)
	) name9860 (
		\wishbone_bd_ram_mem3_reg[184][27]/P0001 ,
		_w13062_,
		_w20372_
	);
	LUT2 #(
		.INIT('h8)
	) name9861 (
		\wishbone_bd_ram_mem3_reg[111][27]/P0001 ,
		_w12744_,
		_w20373_
	);
	LUT2 #(
		.INIT('h8)
	) name9862 (
		\wishbone_bd_ram_mem3_reg[117][27]/P0001 ,
		_w12715_,
		_w20374_
	);
	LUT2 #(
		.INIT('h8)
	) name9863 (
		\wishbone_bd_ram_mem3_reg[193][27]/P0001 ,
		_w13056_,
		_w20375_
	);
	LUT2 #(
		.INIT('h8)
	) name9864 (
		\wishbone_bd_ram_mem3_reg[220][27]/P0001 ,
		_w13066_,
		_w20376_
	);
	LUT2 #(
		.INIT('h8)
	) name9865 (
		\wishbone_bd_ram_mem3_reg[134][27]/P0001 ,
		_w12763_,
		_w20377_
	);
	LUT2 #(
		.INIT('h8)
	) name9866 (
		\wishbone_bd_ram_mem3_reg[187][27]/P0001 ,
		_w13196_,
		_w20378_
	);
	LUT2 #(
		.INIT('h8)
	) name9867 (
		\wishbone_bd_ram_mem3_reg[7][27]/P0001 ,
		_w12728_,
		_w20379_
	);
	LUT2 #(
		.INIT('h8)
	) name9868 (
		\wishbone_bd_ram_mem3_reg[63][27]/P0001 ,
		_w12850_,
		_w20380_
	);
	LUT2 #(
		.INIT('h8)
	) name9869 (
		\wishbone_bd_ram_mem3_reg[49][27]/P0001 ,
		_w12994_,
		_w20381_
	);
	LUT2 #(
		.INIT('h8)
	) name9870 (
		\wishbone_bd_ram_mem3_reg[53][27]/P0001 ,
		_w13020_,
		_w20382_
	);
	LUT2 #(
		.INIT('h8)
	) name9871 (
		\wishbone_bd_ram_mem3_reg[222][27]/P0001 ,
		_w13094_,
		_w20383_
	);
	LUT2 #(
		.INIT('h8)
	) name9872 (
		\wishbone_bd_ram_mem3_reg[31][27]/P0001 ,
		_w13198_,
		_w20384_
	);
	LUT2 #(
		.INIT('h8)
	) name9873 (
		\wishbone_bd_ram_mem3_reg[179][27]/P0001 ,
		_w13050_,
		_w20385_
	);
	LUT2 #(
		.INIT('h8)
	) name9874 (
		\wishbone_bd_ram_mem3_reg[190][27]/P0001 ,
		_w12858_,
		_w20386_
	);
	LUT2 #(
		.INIT('h8)
	) name9875 (
		\wishbone_bd_ram_mem3_reg[130][27]/P0001 ,
		_w12914_,
		_w20387_
	);
	LUT2 #(
		.INIT('h8)
	) name9876 (
		\wishbone_bd_ram_mem3_reg[39][27]/P0001 ,
		_w13018_,
		_w20388_
	);
	LUT2 #(
		.INIT('h8)
	) name9877 (
		\wishbone_bd_ram_mem3_reg[127][27]/P0001 ,
		_w13164_,
		_w20389_
	);
	LUT2 #(
		.INIT('h8)
	) name9878 (
		\wishbone_bd_ram_mem3_reg[116][27]/P0001 ,
		_w12998_,
		_w20390_
	);
	LUT2 #(
		.INIT('h8)
	) name9879 (
		\wishbone_bd_ram_mem3_reg[159][27]/P0001 ,
		_w12774_,
		_w20391_
	);
	LUT2 #(
		.INIT('h8)
	) name9880 (
		\wishbone_bd_ram_mem3_reg[233][27]/P0001 ,
		_w12836_,
		_w20392_
	);
	LUT2 #(
		.INIT('h8)
	) name9881 (
		\wishbone_bd_ram_mem3_reg[204][27]/P0001 ,
		_w13162_,
		_w20393_
	);
	LUT2 #(
		.INIT('h8)
	) name9882 (
		\wishbone_bd_ram_mem3_reg[213][27]/P0001 ,
		_w13002_,
		_w20394_
	);
	LUT2 #(
		.INIT('h8)
	) name9883 (
		\wishbone_bd_ram_mem3_reg[5][27]/P0001 ,
		_w12878_,
		_w20395_
	);
	LUT2 #(
		.INIT('h8)
	) name9884 (
		\wishbone_bd_ram_mem3_reg[61][27]/P0001 ,
		_w12725_,
		_w20396_
	);
	LUT2 #(
		.INIT('h8)
	) name9885 (
		\wishbone_bd_ram_mem3_reg[6][27]/P0001 ,
		_w12968_,
		_w20397_
	);
	LUT2 #(
		.INIT('h8)
	) name9886 (
		\wishbone_bd_ram_mem3_reg[110][27]/P0001 ,
		_w13046_,
		_w20398_
	);
	LUT2 #(
		.INIT('h8)
	) name9887 (
		\wishbone_bd_ram_mem3_reg[143][27]/P0001 ,
		_w12922_,
		_w20399_
	);
	LUT2 #(
		.INIT('h8)
	) name9888 (
		\wishbone_bd_ram_mem3_reg[173][27]/P0001 ,
		_w12854_,
		_w20400_
	);
	LUT2 #(
		.INIT('h8)
	) name9889 (
		\wishbone_bd_ram_mem3_reg[189][27]/P0001 ,
		_w13042_,
		_w20401_
	);
	LUT2 #(
		.INIT('h8)
	) name9890 (
		\wishbone_bd_ram_mem3_reg[249][27]/P0001 ,
		_w12900_,
		_w20402_
	);
	LUT2 #(
		.INIT('h8)
	) name9891 (
		\wishbone_bd_ram_mem3_reg[138][27]/P0001 ,
		_w12958_,
		_w20403_
	);
	LUT2 #(
		.INIT('h8)
	) name9892 (
		\wishbone_bd_ram_mem3_reg[99][27]/P0001 ,
		_w13038_,
		_w20404_
	);
	LUT2 #(
		.INIT('h8)
	) name9893 (
		\wishbone_bd_ram_mem3_reg[239][27]/P0001 ,
		_w12862_,
		_w20405_
	);
	LUT2 #(
		.INIT('h8)
	) name9894 (
		\wishbone_bd_ram_mem3_reg[164][27]/P0001 ,
		_w12876_,
		_w20406_
	);
	LUT2 #(
		.INIT('h8)
	) name9895 (
		\wishbone_bd_ram_mem3_reg[154][27]/P0001 ,
		_w12962_,
		_w20407_
	);
	LUT2 #(
		.INIT('h8)
	) name9896 (
		\wishbone_bd_ram_mem3_reg[244][27]/P0001 ,
		_w12747_,
		_w20408_
	);
	LUT2 #(
		.INIT('h8)
	) name9897 (
		\wishbone_bd_ram_mem3_reg[225][27]/P0001 ,
		_w13092_,
		_w20409_
	);
	LUT2 #(
		.INIT('h8)
	) name9898 (
		\wishbone_bd_ram_mem3_reg[242][27]/P0001 ,
		_w12932_,
		_w20410_
	);
	LUT2 #(
		.INIT('h8)
	) name9899 (
		\wishbone_bd_ram_mem3_reg[74][27]/P0001 ,
		_w12812_,
		_w20411_
	);
	LUT2 #(
		.INIT('h8)
	) name9900 (
		\wishbone_bd_ram_mem3_reg[37][27]/P0001 ,
		_w13102_,
		_w20412_
	);
	LUT2 #(
		.INIT('h8)
	) name9901 (
		\wishbone_bd_ram_mem3_reg[120][27]/P0001 ,
		_w12707_,
		_w20413_
	);
	LUT2 #(
		.INIT('h8)
	) name9902 (
		\wishbone_bd_ram_mem3_reg[177][27]/P0001 ,
		_w12996_,
		_w20414_
	);
	LUT2 #(
		.INIT('h8)
	) name9903 (
		\wishbone_bd_ram_mem3_reg[68][27]/P0001 ,
		_w12946_,
		_w20415_
	);
	LUT2 #(
		.INIT('h8)
	) name9904 (
		\wishbone_bd_ram_mem3_reg[136][27]/P0001 ,
		_w13064_,
		_w20416_
	);
	LUT2 #(
		.INIT('h8)
	) name9905 (
		\wishbone_bd_ram_mem3_reg[16][27]/P0001 ,
		_w13140_,
		_w20417_
	);
	LUT2 #(
		.INIT('h8)
	) name9906 (
		\wishbone_bd_ram_mem3_reg[175][27]/P0001 ,
		_w13126_,
		_w20418_
	);
	LUT2 #(
		.INIT('h8)
	) name9907 (
		\wishbone_bd_ram_mem3_reg[107][27]/P0001 ,
		_w12749_,
		_w20419_
	);
	LUT2 #(
		.INIT('h8)
	) name9908 (
		\wishbone_bd_ram_mem3_reg[181][27]/P0001 ,
		_w12828_,
		_w20420_
	);
	LUT2 #(
		.INIT('h8)
	) name9909 (
		\wishbone_bd_ram_mem3_reg[89][27]/P0001 ,
		_w12964_,
		_w20421_
	);
	LUT2 #(
		.INIT('h8)
	) name9910 (
		\wishbone_bd_ram_mem3_reg[252][27]/P0001 ,
		_w13080_,
		_w20422_
	);
	LUT2 #(
		.INIT('h8)
	) name9911 (
		\wishbone_bd_ram_mem3_reg[227][27]/P0001 ,
		_w12936_,
		_w20423_
	);
	LUT2 #(
		.INIT('h8)
	) name9912 (
		\wishbone_bd_ram_mem3_reg[13][27]/P0001 ,
		_w13178_,
		_w20424_
	);
	LUT2 #(
		.INIT('h8)
	) name9913 (
		\wishbone_bd_ram_mem3_reg[124][27]/P0001 ,
		_w13058_,
		_w20425_
	);
	LUT2 #(
		.INIT('h8)
	) name9914 (
		\wishbone_bd_ram_mem3_reg[169][27]/P0001 ,
		_w12722_,
		_w20426_
	);
	LUT2 #(
		.INIT('h8)
	) name9915 (
		\wishbone_bd_ram_mem3_reg[128][27]/P0001 ,
		_w12793_,
		_w20427_
	);
	LUT2 #(
		.INIT('h8)
	) name9916 (
		\wishbone_bd_ram_mem3_reg[200][27]/P0001 ,
		_w12988_,
		_w20428_
	);
	LUT2 #(
		.INIT('h8)
	) name9917 (
		\wishbone_bd_ram_mem3_reg[80][27]/P0001 ,
		_w12689_,
		_w20429_
	);
	LUT2 #(
		.INIT('h8)
	) name9918 (
		\wishbone_bd_ram_mem3_reg[3][27]/P0001 ,
		_w12866_,
		_w20430_
	);
	LUT2 #(
		.INIT('h8)
	) name9919 (
		\wishbone_bd_ram_mem3_reg[52][27]/P0001 ,
		_w13082_,
		_w20431_
	);
	LUT2 #(
		.INIT('h8)
	) name9920 (
		\wishbone_bd_ram_mem3_reg[73][27]/P0001 ,
		_w12918_,
		_w20432_
	);
	LUT2 #(
		.INIT('h8)
	) name9921 (
		\wishbone_bd_ram_mem3_reg[55][27]/P0001 ,
		_w12785_,
		_w20433_
	);
	LUT2 #(
		.INIT('h8)
	) name9922 (
		\wishbone_bd_ram_mem3_reg[219][27]/P0001 ,
		_w12806_,
		_w20434_
	);
	LUT2 #(
		.INIT('h8)
	) name9923 (
		\wishbone_bd_ram_mem3_reg[147][27]/P0001 ,
		_w13146_,
		_w20435_
	);
	LUT2 #(
		.INIT('h8)
	) name9924 (
		\wishbone_bd_ram_mem3_reg[180][27]/P0001 ,
		_w12791_,
		_w20436_
	);
	LUT2 #(
		.INIT('h8)
	) name9925 (
		\wishbone_bd_ram_mem3_reg[214][27]/P0001 ,
		_w12984_,
		_w20437_
	);
	LUT2 #(
		.INIT('h8)
	) name9926 (
		\wishbone_bd_ram_mem3_reg[113][27]/P0001 ,
		_w13026_,
		_w20438_
	);
	LUT2 #(
		.INIT('h8)
	) name9927 (
		\wishbone_bd_ram_mem3_reg[119][27]/P0001 ,
		_w13048_,
		_w20439_
	);
	LUT2 #(
		.INIT('h8)
	) name9928 (
		\wishbone_bd_ram_mem3_reg[132][27]/P0001 ,
		_w12992_,
		_w20440_
	);
	LUT2 #(
		.INIT('h8)
	) name9929 (
		\wishbone_bd_ram_mem3_reg[248][27]/P0001 ,
		_w12789_,
		_w20441_
	);
	LUT2 #(
		.INIT('h8)
	) name9930 (
		\wishbone_bd_ram_mem3_reg[126][27]/P0001 ,
		_w13218_,
		_w20442_
	);
	LUT2 #(
		.INIT('h8)
	) name9931 (
		\wishbone_bd_ram_mem3_reg[62][27]/P0001 ,
		_w12673_,
		_w20443_
	);
	LUT2 #(
		.INIT('h8)
	) name9932 (
		\wishbone_bd_ram_mem3_reg[58][27]/P0001 ,
		_w13070_,
		_w20444_
	);
	LUT2 #(
		.INIT('h8)
	) name9933 (
		\wishbone_bd_ram_mem3_reg[208][27]/P0001 ,
		_w13032_,
		_w20445_
	);
	LUT2 #(
		.INIT('h8)
	) name9934 (
		\wishbone_bd_ram_mem3_reg[192][27]/P0001 ,
		_w12938_,
		_w20446_
	);
	LUT2 #(
		.INIT('h8)
	) name9935 (
		\wishbone_bd_ram_mem3_reg[171][27]/P0001 ,
		_w12910_,
		_w20447_
	);
	LUT2 #(
		.INIT('h8)
	) name9936 (
		\wishbone_bd_ram_mem3_reg[98][27]/P0001 ,
		_w12816_,
		_w20448_
	);
	LUT2 #(
		.INIT('h8)
	) name9937 (
		\wishbone_bd_ram_mem3_reg[75][27]/P0001 ,
		_w12826_,
		_w20449_
	);
	LUT2 #(
		.INIT('h8)
	) name9938 (
		\wishbone_bd_ram_mem3_reg[25][27]/P0001 ,
		_w13108_,
		_w20450_
	);
	LUT2 #(
		.INIT('h8)
	) name9939 (
		\wishbone_bd_ram_mem3_reg[43][27]/P0001 ,
		_w13200_,
		_w20451_
	);
	LUT2 #(
		.INIT('h8)
	) name9940 (
		\wishbone_bd_ram_mem3_reg[153][27]/P0001 ,
		_w12890_,
		_w20452_
	);
	LUT2 #(
		.INIT('h8)
	) name9941 (
		\wishbone_bd_ram_mem3_reg[133][27]/P0001 ,
		_w12761_,
		_w20453_
	);
	LUT2 #(
		.INIT('h8)
	) name9942 (
		\wishbone_bd_ram_mem3_reg[60][27]/P0001 ,
		_w13204_,
		_w20454_
	);
	LUT2 #(
		.INIT('h8)
	) name9943 (
		\wishbone_bd_ram_mem3_reg[123][27]/P0001 ,
		_w13114_,
		_w20455_
	);
	LUT2 #(
		.INIT('h8)
	) name9944 (
		\wishbone_bd_ram_mem3_reg[84][27]/P0001 ,
		_w12934_,
		_w20456_
	);
	LUT2 #(
		.INIT('h8)
	) name9945 (
		\wishbone_bd_ram_mem3_reg[205][27]/P0001 ,
		_w13068_,
		_w20457_
	);
	LUT2 #(
		.INIT('h8)
	) name9946 (
		\wishbone_bd_ram_mem3_reg[78][27]/P0001 ,
		_w12874_,
		_w20458_
	);
	LUT2 #(
		.INIT('h8)
	) name9947 (
		\wishbone_bd_ram_mem3_reg[221][27]/P0001 ,
		_w12802_,
		_w20459_
	);
	LUT2 #(
		.INIT('h8)
	) name9948 (
		\wishbone_bd_ram_mem3_reg[88][27]/P0001 ,
		_w12860_,
		_w20460_
	);
	LUT2 #(
		.INIT('h8)
	) name9949 (
		\wishbone_bd_ram_mem3_reg[243][27]/P0001 ,
		_w12804_,
		_w20461_
	);
	LUT2 #(
		.INIT('h8)
	) name9950 (
		\wishbone_bd_ram_mem3_reg[122][27]/P0001 ,
		_w13130_,
		_w20462_
	);
	LUT2 #(
		.INIT('h8)
	) name9951 (
		\wishbone_bd_ram_mem3_reg[91][27]/P0001 ,
		_w13074_,
		_w20463_
	);
	LUT2 #(
		.INIT('h8)
	) name9952 (
		\wishbone_bd_ram_mem3_reg[65][27]/P0001 ,
		_w13176_,
		_w20464_
	);
	LUT2 #(
		.INIT('h8)
	) name9953 (
		\wishbone_bd_ram_mem3_reg[162][27]/P0001 ,
		_w13098_,
		_w20465_
	);
	LUT2 #(
		.INIT('h8)
	) name9954 (
		\wishbone_bd_ram_mem3_reg[238][27]/P0001 ,
		_w13160_,
		_w20466_
	);
	LUT2 #(
		.INIT('h8)
	) name9955 (
		\wishbone_bd_ram_mem3_reg[47][27]/P0001 ,
		_w12904_,
		_w20467_
	);
	LUT2 #(
		.INIT('h8)
	) name9956 (
		\wishbone_bd_ram_mem3_reg[201][27]/P0001 ,
		_w12822_,
		_w20468_
	);
	LUT2 #(
		.INIT('h8)
	) name9957 (
		\wishbone_bd_ram_mem3_reg[182][27]/P0001 ,
		_w12820_,
		_w20469_
	);
	LUT2 #(
		.INIT('h8)
	) name9958 (
		\wishbone_bd_ram_mem3_reg[51][27]/P0001 ,
		_w13024_,
		_w20470_
	);
	LUT2 #(
		.INIT('h8)
	) name9959 (
		\wishbone_bd_ram_mem3_reg[101][27]/P0001 ,
		_w13192_,
		_w20471_
	);
	LUT2 #(
		.INIT('h8)
	) name9960 (
		\wishbone_bd_ram_mem3_reg[210][27]/P0001 ,
		_w12924_,
		_w20472_
	);
	LUT2 #(
		.INIT('h8)
	) name9961 (
		\wishbone_bd_ram_mem3_reg[144][27]/P0001 ,
		_w12756_,
		_w20473_
	);
	LUT2 #(
		.INIT('h8)
	) name9962 (
		\wishbone_bd_ram_mem3_reg[142][27]/P0001 ,
		_w12928_,
		_w20474_
	);
	LUT2 #(
		.INIT('h8)
	) name9963 (
		\wishbone_bd_ram_mem3_reg[83][27]/P0001 ,
		_w12916_,
		_w20475_
	);
	LUT2 #(
		.INIT('h8)
	) name9964 (
		\wishbone_bd_ram_mem3_reg[76][27]/P0001 ,
		_w13184_,
		_w20476_
	);
	LUT2 #(
		.INIT('h8)
	) name9965 (
		\wishbone_bd_ram_mem3_reg[102][27]/P0001 ,
		_w12685_,
		_w20477_
	);
	LUT2 #(
		.INIT('h8)
	) name9966 (
		\wishbone_bd_ram_mem3_reg[35][27]/P0001 ,
		_w12703_,
		_w20478_
	);
	LUT2 #(
		.INIT('h8)
	) name9967 (
		\wishbone_bd_ram_mem3_reg[29][27]/P0001 ,
		_w12952_,
		_w20479_
	);
	LUT2 #(
		.INIT('h8)
	) name9968 (
		\wishbone_bd_ram_mem3_reg[151][27]/P0001 ,
		_w13142_,
		_w20480_
	);
	LUT2 #(
		.INIT('h8)
	) name9969 (
		\wishbone_bd_ram_mem3_reg[12][27]/P0001 ,
		_w13118_,
		_w20481_
	);
	LUT2 #(
		.INIT('h8)
	) name9970 (
		\wishbone_bd_ram_mem3_reg[86][27]/P0001 ,
		_w12735_,
		_w20482_
	);
	LUT2 #(
		.INIT('h8)
	) name9971 (
		\wishbone_bd_ram_mem3_reg[215][27]/P0001 ,
		_w12974_,
		_w20483_
	);
	LUT2 #(
		.INIT('h8)
	) name9972 (
		\wishbone_bd_ram_mem3_reg[129][27]/P0001 ,
		_w12776_,
		_w20484_
	);
	LUT2 #(
		.INIT('h8)
	) name9973 (
		\wishbone_bd_ram_mem3_reg[209][27]/P0001 ,
		_w13152_,
		_w20485_
	);
	LUT2 #(
		.INIT('h8)
	) name9974 (
		\wishbone_bd_ram_mem3_reg[158][27]/P0001 ,
		_w12898_,
		_w20486_
	);
	LUT2 #(
		.INIT('h8)
	) name9975 (
		\wishbone_bd_ram_mem3_reg[112][27]/P0001 ,
		_w12733_,
		_w20487_
	);
	LUT2 #(
		.INIT('h8)
	) name9976 (
		\wishbone_bd_ram_mem3_reg[85][27]/P0001 ,
		_w13216_,
		_w20488_
	);
	LUT2 #(
		.INIT('h8)
	) name9977 (
		\wishbone_bd_ram_mem3_reg[125][27]/P0001 ,
		_w12956_,
		_w20489_
	);
	LUT2 #(
		.INIT('h8)
	) name9978 (
		\wishbone_bd_ram_mem3_reg[54][27]/P0001 ,
		_w12770_,
		_w20490_
	);
	LUT2 #(
		.INIT('h8)
	) name9979 (
		\wishbone_bd_ram_mem3_reg[141][27]/P0001 ,
		_w13004_,
		_w20491_
	);
	LUT2 #(
		.INIT('h8)
	) name9980 (
		\wishbone_bd_ram_mem3_reg[178][27]/P0001 ,
		_w12886_,
		_w20492_
	);
	LUT2 #(
		.INIT('h8)
	) name9981 (
		\wishbone_bd_ram_mem3_reg[20][27]/P0001 ,
		_w13174_,
		_w20493_
	);
	LUT2 #(
		.INIT('h8)
	) name9982 (
		\wishbone_bd_ram_mem3_reg[172][27]/P0001 ,
		_w12944_,
		_w20494_
	);
	LUT2 #(
		.INIT('h8)
	) name9983 (
		\wishbone_bd_ram_mem3_reg[218][27]/P0001 ,
		_w13206_,
		_w20495_
	);
	LUT2 #(
		.INIT('h8)
	) name9984 (
		\wishbone_bd_ram_mem3_reg[93][27]/P0001 ,
		_w13016_,
		_w20496_
	);
	LUT2 #(
		.INIT('h8)
	) name9985 (
		\wishbone_bd_ram_mem3_reg[11][27]/P0001 ,
		_w13194_,
		_w20497_
	);
	LUT2 #(
		.INIT('h8)
	) name9986 (
		\wishbone_bd_ram_mem3_reg[79][27]/P0001 ,
		_w13212_,
		_w20498_
	);
	LUT2 #(
		.INIT('h8)
	) name9987 (
		\wishbone_bd_ram_mem3_reg[137][27]/P0001 ,
		_w13168_,
		_w20499_
	);
	LUT2 #(
		.INIT('h8)
	) name9988 (
		\wishbone_bd_ram_mem3_reg[135][27]/P0001 ,
		_w13124_,
		_w20500_
	);
	LUT2 #(
		.INIT('h8)
	) name9989 (
		\wishbone_bd_ram_mem3_reg[168][27]/P0001 ,
		_w13208_,
		_w20501_
	);
	LUT2 #(
		.INIT('h8)
	) name9990 (
		\wishbone_bd_ram_mem3_reg[254][27]/P0001 ,
		_w12892_,
		_w20502_
	);
	LUT2 #(
		.INIT('h8)
	) name9991 (
		\wishbone_bd_ram_mem3_reg[46][27]/P0001 ,
		_w12884_,
		_w20503_
	);
	LUT2 #(
		.INIT('h8)
	) name9992 (
		\wishbone_bd_ram_mem3_reg[223][27]/P0001 ,
		_w12838_,
		_w20504_
	);
	LUT2 #(
		.INIT('h8)
	) name9993 (
		\wishbone_bd_ram_mem3_reg[251][27]/P0001 ,
		_w13054_,
		_w20505_
	);
	LUT2 #(
		.INIT('h8)
	) name9994 (
		\wishbone_bd_ram_mem3_reg[235][27]/P0001 ,
		_w12696_,
		_w20506_
	);
	LUT2 #(
		.INIT('h8)
	) name9995 (
		\wishbone_bd_ram_mem3_reg[152][27]/P0001 ,
		_w12966_,
		_w20507_
	);
	LUT2 #(
		.INIT('h8)
	) name9996 (
		\wishbone_bd_ram_mem3_reg[224][27]/P0001 ,
		_w12902_,
		_w20508_
	);
	LUT2 #(
		.INIT('h8)
	) name9997 (
		\wishbone_bd_ram_mem3_reg[156][27]/P0001 ,
		_w13190_,
		_w20509_
	);
	LUT2 #(
		.INIT('h8)
	) name9998 (
		\wishbone_bd_ram_mem3_reg[92][27]/P0001 ,
		_w13010_,
		_w20510_
	);
	LUT2 #(
		.INIT('h8)
	) name9999 (
		\wishbone_bd_ram_mem3_reg[90][27]/P0001 ,
		_w12978_,
		_w20511_
	);
	LUT2 #(
		.INIT('h8)
	) name10000 (
		\wishbone_bd_ram_mem3_reg[231][27]/P0001 ,
		_w12856_,
		_w20512_
	);
	LUT2 #(
		.INIT('h8)
	) name10001 (
		\wishbone_bd_ram_mem3_reg[82][27]/P0001 ,
		_w12942_,
		_w20513_
	);
	LUT2 #(
		.INIT('h8)
	) name10002 (
		\wishbone_bd_ram_mem3_reg[195][27]/P0001 ,
		_w13144_,
		_w20514_
	);
	LUT2 #(
		.INIT('h8)
	) name10003 (
		\wishbone_bd_ram_mem3_reg[50][27]/P0001 ,
		_w13150_,
		_w20515_
	);
	LUT2 #(
		.INIT('h8)
	) name10004 (
		\wishbone_bd_ram_mem3_reg[185][27]/P0001 ,
		_w12940_,
		_w20516_
	);
	LUT2 #(
		.INIT('h8)
	) name10005 (
		\wishbone_bd_ram_mem3_reg[19][27]/P0001 ,
		_w13012_,
		_w20517_
	);
	LUT2 #(
		.INIT('h8)
	) name10006 (
		\wishbone_bd_ram_mem3_reg[229][27]/P0001 ,
		_w12711_,
		_w20518_
	);
	LUT2 #(
		.INIT('h8)
	) name10007 (
		\wishbone_bd_ram_mem3_reg[196][27]/P0001 ,
		_w13090_,
		_w20519_
	);
	LUT2 #(
		.INIT('h8)
	) name10008 (
		\wishbone_bd_ram_mem3_reg[105][27]/P0001 ,
		_w12751_,
		_w20520_
	);
	LUT2 #(
		.INIT('h8)
	) name10009 (
		\wishbone_bd_ram_mem3_reg[145][27]/P0001 ,
		_w13106_,
		_w20521_
	);
	LUT2 #(
		.INIT('h8)
	) name10010 (
		\wishbone_bd_ram_mem3_reg[186][27]/P0001 ,
		_w12783_,
		_w20522_
	);
	LUT2 #(
		.INIT('h8)
	) name10011 (
		\wishbone_bd_ram_mem3_reg[150][27]/P0001 ,
		_w13136_,
		_w20523_
	);
	LUT2 #(
		.INIT('h8)
	) name10012 (
		\wishbone_bd_ram_mem3_reg[211][27]/P0001 ,
		_w13166_,
		_w20524_
	);
	LUT2 #(
		.INIT('h8)
	) name10013 (
		\wishbone_bd_ram_mem3_reg[197][27]/P0001 ,
		_w12834_,
		_w20525_
	);
	LUT2 #(
		.INIT('h8)
	) name10014 (
		\wishbone_bd_ram_mem3_reg[67][27]/P0001 ,
		_w13134_,
		_w20526_
	);
	LUT2 #(
		.INIT('h8)
	) name10015 (
		\wishbone_bd_ram_mem3_reg[114][27]/P0001 ,
		_w13202_,
		_w20527_
	);
	LUT2 #(
		.INIT('h8)
	) name10016 (
		\wishbone_bd_ram_mem3_reg[188][27]/P0001 ,
		_w12948_,
		_w20528_
	);
	LUT2 #(
		.INIT('h8)
	) name10017 (
		\wishbone_bd_ram_mem3_reg[226][27]/P0001 ,
		_w13138_,
		_w20529_
	);
	LUT2 #(
		.INIT('h8)
	) name10018 (
		\wishbone_bd_ram_mem3_reg[108][27]/P0001 ,
		_w13156_,
		_w20530_
	);
	LUT2 #(
		.INIT('h8)
	) name10019 (
		\wishbone_bd_ram_mem3_reg[246][27]/P0001 ,
		_w13076_,
		_w20531_
	);
	LUT2 #(
		.INIT('h8)
	) name10020 (
		\wishbone_bd_ram_mem3_reg[0][27]/P0001 ,
		_w12717_,
		_w20532_
	);
	LUT2 #(
		.INIT('h8)
	) name10021 (
		\wishbone_bd_ram_mem3_reg[42][27]/P0001 ,
		_w12842_,
		_w20533_
	);
	LUT2 #(
		.INIT('h8)
	) name10022 (
		\wishbone_bd_ram_mem3_reg[48][27]/P0001 ,
		_w12970_,
		_w20534_
	);
	LUT2 #(
		.INIT('h8)
	) name10023 (
		\wishbone_bd_ram_mem3_reg[44][27]/P0001 ,
		_w12896_,
		_w20535_
	);
	LUT2 #(
		.INIT('h8)
	) name10024 (
		\wishbone_bd_ram_mem3_reg[237][27]/P0001 ,
		_w12990_,
		_w20536_
	);
	LUT2 #(
		.INIT('h8)
	) name10025 (
		\wishbone_bd_ram_mem3_reg[240][27]/P0001 ,
		_w12864_,
		_w20537_
	);
	LUT2 #(
		.INIT('h8)
	) name10026 (
		\wishbone_bd_ram_mem3_reg[97][27]/P0001 ,
		_w13096_,
		_w20538_
	);
	LUT2 #(
		.INIT('h8)
	) name10027 (
		\wishbone_bd_ram_mem3_reg[139][27]/P0001 ,
		_w12814_,
		_w20539_
	);
	LUT2 #(
		.INIT('h8)
	) name10028 (
		\wishbone_bd_ram_mem3_reg[234][27]/P0001 ,
		_w13214_,
		_w20540_
	);
	LUT2 #(
		.INIT('h8)
	) name10029 (
		\wishbone_bd_ram_mem3_reg[206][27]/P0001 ,
		_w12954_,
		_w20541_
	);
	LUT2 #(
		.INIT('h8)
	) name10030 (
		\wishbone_bd_ram_mem3_reg[9][27]/P0001 ,
		_w12808_,
		_w20542_
	);
	LUT2 #(
		.INIT('h8)
	) name10031 (
		\wishbone_bd_ram_mem3_reg[27][27]/P0001 ,
		_w12880_,
		_w20543_
	);
	LUT2 #(
		.INIT('h8)
	) name10032 (
		\wishbone_bd_ram_mem3_reg[95][27]/P0001 ,
		_w12844_,
		_w20544_
	);
	LUT2 #(
		.INIT('h8)
	) name10033 (
		\wishbone_bd_ram_mem3_reg[163][27]/P0001 ,
		_w12882_,
		_w20545_
	);
	LUT2 #(
		.INIT('h8)
	) name10034 (
		\wishbone_bd_ram_mem3_reg[41][27]/P0001 ,
		_w13052_,
		_w20546_
	);
	LUT2 #(
		.INIT('h8)
	) name10035 (
		\wishbone_bd_ram_mem3_reg[36][27]/P0001 ,
		_w12800_,
		_w20547_
	);
	LUT2 #(
		.INIT('h8)
	) name10036 (
		\wishbone_bd_ram_mem3_reg[71][27]/P0001 ,
		_w12798_,
		_w20548_
	);
	LUT2 #(
		.INIT('h8)
	) name10037 (
		\wishbone_bd_ram_mem3_reg[38][27]/P0001 ,
		_w13182_,
		_w20549_
	);
	LUT2 #(
		.INIT('h8)
	) name10038 (
		\wishbone_bd_ram_mem3_reg[2][27]/P0001 ,
		_w13088_,
		_w20550_
	);
	LUT2 #(
		.INIT('h8)
	) name10039 (
		\wishbone_bd_ram_mem3_reg[115][27]/P0001 ,
		_w13112_,
		_w20551_
	);
	LUT2 #(
		.INIT('h8)
	) name10040 (
		\wishbone_bd_ram_mem3_reg[23][27]/P0001 ,
		_w13008_,
		_w20552_
	);
	LUT2 #(
		.INIT('h8)
	) name10041 (
		\wishbone_bd_ram_mem3_reg[149][27]/P0001 ,
		_w12741_,
		_w20553_
	);
	LUT2 #(
		.INIT('h8)
	) name10042 (
		\wishbone_bd_ram_mem3_reg[21][27]/P0001 ,
		_w12906_,
		_w20554_
	);
	LUT2 #(
		.INIT('h8)
	) name10043 (
		\wishbone_bd_ram_mem3_reg[207][27]/P0001 ,
		_w13180_,
		_w20555_
	);
	LUT2 #(
		.INIT('h8)
	) name10044 (
		\wishbone_bd_ram_mem3_reg[165][27]/P0001 ,
		_w13044_,
		_w20556_
	);
	LUT2 #(
		.INIT('h8)
	) name10045 (
		\wishbone_bd_ram_mem3_reg[18][27]/P0001 ,
		_w12679_,
		_w20557_
	);
	LUT2 #(
		.INIT('h8)
	) name10046 (
		\wishbone_bd_ram_mem3_reg[1][27]/P0001 ,
		_w13014_,
		_w20558_
	);
	LUT2 #(
		.INIT('h8)
	) name10047 (
		\wishbone_bd_ram_mem3_reg[167][27]/P0001 ,
		_w12986_,
		_w20559_
	);
	LUT2 #(
		.INIT('h8)
	) name10048 (
		\wishbone_bd_ram_mem3_reg[250][27]/P0001 ,
		_w13128_,
		_w20560_
	);
	LUT2 #(
		.INIT('h8)
	) name10049 (
		\wishbone_bd_ram_mem3_reg[157][27]/P0001 ,
		_w12926_,
		_w20561_
	);
	LUT2 #(
		.INIT('h8)
	) name10050 (
		\wishbone_bd_ram_mem3_reg[166][27]/P0001 ,
		_w13040_,
		_w20562_
	);
	LUT2 #(
		.INIT('h8)
	) name10051 (
		\wishbone_bd_ram_mem3_reg[228][27]/P0001 ,
		_w12765_,
		_w20563_
	);
	LUT2 #(
		.INIT('h8)
	) name10052 (
		\wishbone_bd_ram_mem3_reg[28][27]/P0001 ,
		_w13170_,
		_w20564_
	);
	LUT2 #(
		.INIT('h8)
	) name10053 (
		\wishbone_bd_ram_mem3_reg[174][27]/P0001 ,
		_w12972_,
		_w20565_
	);
	LUT2 #(
		.INIT('h8)
	) name10054 (
		\wishbone_bd_ram_mem3_reg[40][27]/P0001 ,
		_w13132_,
		_w20566_
	);
	LUT2 #(
		.INIT('h8)
	) name10055 (
		\wishbone_bd_ram_mem3_reg[236][27]/P0001 ,
		_w12731_,
		_w20567_
	);
	LUT2 #(
		.INIT('h8)
	) name10056 (
		\wishbone_bd_ram_mem3_reg[81][27]/P0001 ,
		_w12950_,
		_w20568_
	);
	LUT2 #(
		.INIT('h8)
	) name10057 (
		\wishbone_bd_ram_mem3_reg[230][27]/P0001 ,
		_w13036_,
		_w20569_
	);
	LUT2 #(
		.INIT('h8)
	) name10058 (
		\wishbone_bd_ram_mem3_reg[170][27]/P0001 ,
		_w13030_,
		_w20570_
	);
	LUT2 #(
		.INIT('h8)
	) name10059 (
		\wishbone_bd_ram_mem3_reg[217][27]/P0001 ,
		_w13188_,
		_w20571_
	);
	LUT2 #(
		.INIT('h8)
	) name10060 (
		\wishbone_bd_ram_mem3_reg[191][27]/P0001 ,
		_w13034_,
		_w20572_
	);
	LUT2 #(
		.INIT('h8)
	) name10061 (
		\wishbone_bd_ram_mem3_reg[106][27]/P0001 ,
		_w12713_,
		_w20573_
	);
	LUT2 #(
		.INIT('h8)
	) name10062 (
		\wishbone_bd_ram_mem3_reg[255][27]/P0001 ,
		_w13072_,
		_w20574_
	);
	LUT2 #(
		.INIT('h8)
	) name10063 (
		\wishbone_bd_ram_mem3_reg[87][27]/P0001 ,
		_w13154_,
		_w20575_
	);
	LUT2 #(
		.INIT('h8)
	) name10064 (
		\wishbone_bd_ram_mem3_reg[15][27]/P0001 ,
		_w13210_,
		_w20576_
	);
	LUT2 #(
		.INIT('h8)
	) name10065 (
		\wishbone_bd_ram_mem3_reg[22][27]/P0001 ,
		_w13110_,
		_w20577_
	);
	LUT2 #(
		.INIT('h8)
	) name10066 (
		\wishbone_bd_ram_mem3_reg[64][27]/P0001 ,
		_w12976_,
		_w20578_
	);
	LUT2 #(
		.INIT('h8)
	) name10067 (
		\wishbone_bd_ram_mem3_reg[17][27]/P0001 ,
		_w12848_,
		_w20579_
	);
	LUT2 #(
		.INIT('h8)
	) name10068 (
		\wishbone_bd_ram_mem3_reg[33][27]/P0001 ,
		_w12980_,
		_w20580_
	);
	LUT2 #(
		.INIT('h8)
	) name10069 (
		\wishbone_bd_ram_mem3_reg[194][27]/P0001 ,
		_w12772_,
		_w20581_
	);
	LUT2 #(
		.INIT('h8)
	) name10070 (
		\wishbone_bd_ram_mem3_reg[161][27]/P0001 ,
		_w12754_,
		_w20582_
	);
	LUT2 #(
		.INIT('h8)
	) name10071 (
		\wishbone_bd_ram_mem3_reg[14][27]/P0001 ,
		_w13086_,
		_w20583_
	);
	LUT2 #(
		.INIT('h8)
	) name10072 (
		\wishbone_bd_ram_mem3_reg[202][27]/P0001 ,
		_w12870_,
		_w20584_
	);
	LUT2 #(
		.INIT('h8)
	) name10073 (
		\wishbone_bd_ram_mem3_reg[245][27]/P0001 ,
		_w13022_,
		_w20585_
	);
	LUT2 #(
		.INIT('h8)
	) name10074 (
		\wishbone_bd_ram_mem3_reg[146][27]/P0001 ,
		_w13060_,
		_w20586_
	);
	LUT2 #(
		.INIT('h8)
	) name10075 (
		\wishbone_bd_ram_mem3_reg[45][27]/P0001 ,
		_w12908_,
		_w20587_
	);
	LUT2 #(
		.INIT('h8)
	) name10076 (
		\wishbone_bd_ram_mem3_reg[66][27]/P0001 ,
		_w12824_,
		_w20588_
	);
	LUT2 #(
		.INIT('h8)
	) name10077 (
		\wishbone_bd_ram_mem3_reg[253][27]/P0001 ,
		_w13100_,
		_w20589_
	);
	LUT2 #(
		.INIT('h8)
	) name10078 (
		\wishbone_bd_ram_mem3_reg[109][27]/P0001 ,
		_w12888_,
		_w20590_
	);
	LUT2 #(
		.INIT('h8)
	) name10079 (
		\wishbone_bd_ram_mem3_reg[69][27]/P0001 ,
		_w12738_,
		_w20591_
	);
	LUT2 #(
		.INIT('h8)
	) name10080 (
		\wishbone_bd_ram_mem3_reg[199][27]/P0001 ,
		_w12768_,
		_w20592_
	);
	LUT2 #(
		.INIT('h8)
	) name10081 (
		\wishbone_bd_ram_mem3_reg[57][27]/P0001 ,
		_w13116_,
		_w20593_
	);
	LUT2 #(
		.INIT('h8)
	) name10082 (
		\wishbone_bd_ram_mem3_reg[100][27]/P0001 ,
		_w12960_,
		_w20594_
	);
	LUT2 #(
		.INIT('h8)
	) name10083 (
		\wishbone_bd_ram_mem3_reg[59][27]/P0001 ,
		_w12780_,
		_w20595_
	);
	LUT2 #(
		.INIT('h8)
	) name10084 (
		\wishbone_bd_ram_mem3_reg[10][27]/P0001 ,
		_w13172_,
		_w20596_
	);
	LUT2 #(
		.INIT('h8)
	) name10085 (
		\wishbone_bd_ram_mem3_reg[72][27]/P0001 ,
		_w12810_,
		_w20597_
	);
	LUT2 #(
		.INIT('h8)
	) name10086 (
		\wishbone_bd_ram_mem3_reg[241][27]/P0001 ,
		_w13006_,
		_w20598_
	);
	LUT2 #(
		.INIT('h8)
	) name10087 (
		\wishbone_bd_ram_mem3_reg[56][27]/P0001 ,
		_w12778_,
		_w20599_
	);
	LUT2 #(
		.INIT('h8)
	) name10088 (
		\wishbone_bd_ram_mem3_reg[140][27]/P0001 ,
		_w12894_,
		_w20600_
	);
	LUT2 #(
		.INIT('h1)
	) name10089 (
		_w20345_,
		_w20346_,
		_w20601_
	);
	LUT2 #(
		.INIT('h1)
	) name10090 (
		_w20347_,
		_w20348_,
		_w20602_
	);
	LUT2 #(
		.INIT('h1)
	) name10091 (
		_w20349_,
		_w20350_,
		_w20603_
	);
	LUT2 #(
		.INIT('h1)
	) name10092 (
		_w20351_,
		_w20352_,
		_w20604_
	);
	LUT2 #(
		.INIT('h1)
	) name10093 (
		_w20353_,
		_w20354_,
		_w20605_
	);
	LUT2 #(
		.INIT('h1)
	) name10094 (
		_w20355_,
		_w20356_,
		_w20606_
	);
	LUT2 #(
		.INIT('h1)
	) name10095 (
		_w20357_,
		_w20358_,
		_w20607_
	);
	LUT2 #(
		.INIT('h1)
	) name10096 (
		_w20359_,
		_w20360_,
		_w20608_
	);
	LUT2 #(
		.INIT('h1)
	) name10097 (
		_w20361_,
		_w20362_,
		_w20609_
	);
	LUT2 #(
		.INIT('h1)
	) name10098 (
		_w20363_,
		_w20364_,
		_w20610_
	);
	LUT2 #(
		.INIT('h1)
	) name10099 (
		_w20365_,
		_w20366_,
		_w20611_
	);
	LUT2 #(
		.INIT('h1)
	) name10100 (
		_w20367_,
		_w20368_,
		_w20612_
	);
	LUT2 #(
		.INIT('h1)
	) name10101 (
		_w20369_,
		_w20370_,
		_w20613_
	);
	LUT2 #(
		.INIT('h1)
	) name10102 (
		_w20371_,
		_w20372_,
		_w20614_
	);
	LUT2 #(
		.INIT('h1)
	) name10103 (
		_w20373_,
		_w20374_,
		_w20615_
	);
	LUT2 #(
		.INIT('h1)
	) name10104 (
		_w20375_,
		_w20376_,
		_w20616_
	);
	LUT2 #(
		.INIT('h1)
	) name10105 (
		_w20377_,
		_w20378_,
		_w20617_
	);
	LUT2 #(
		.INIT('h1)
	) name10106 (
		_w20379_,
		_w20380_,
		_w20618_
	);
	LUT2 #(
		.INIT('h1)
	) name10107 (
		_w20381_,
		_w20382_,
		_w20619_
	);
	LUT2 #(
		.INIT('h1)
	) name10108 (
		_w20383_,
		_w20384_,
		_w20620_
	);
	LUT2 #(
		.INIT('h1)
	) name10109 (
		_w20385_,
		_w20386_,
		_w20621_
	);
	LUT2 #(
		.INIT('h1)
	) name10110 (
		_w20387_,
		_w20388_,
		_w20622_
	);
	LUT2 #(
		.INIT('h1)
	) name10111 (
		_w20389_,
		_w20390_,
		_w20623_
	);
	LUT2 #(
		.INIT('h1)
	) name10112 (
		_w20391_,
		_w20392_,
		_w20624_
	);
	LUT2 #(
		.INIT('h1)
	) name10113 (
		_w20393_,
		_w20394_,
		_w20625_
	);
	LUT2 #(
		.INIT('h1)
	) name10114 (
		_w20395_,
		_w20396_,
		_w20626_
	);
	LUT2 #(
		.INIT('h1)
	) name10115 (
		_w20397_,
		_w20398_,
		_w20627_
	);
	LUT2 #(
		.INIT('h1)
	) name10116 (
		_w20399_,
		_w20400_,
		_w20628_
	);
	LUT2 #(
		.INIT('h1)
	) name10117 (
		_w20401_,
		_w20402_,
		_w20629_
	);
	LUT2 #(
		.INIT('h1)
	) name10118 (
		_w20403_,
		_w20404_,
		_w20630_
	);
	LUT2 #(
		.INIT('h1)
	) name10119 (
		_w20405_,
		_w20406_,
		_w20631_
	);
	LUT2 #(
		.INIT('h1)
	) name10120 (
		_w20407_,
		_w20408_,
		_w20632_
	);
	LUT2 #(
		.INIT('h1)
	) name10121 (
		_w20409_,
		_w20410_,
		_w20633_
	);
	LUT2 #(
		.INIT('h1)
	) name10122 (
		_w20411_,
		_w20412_,
		_w20634_
	);
	LUT2 #(
		.INIT('h1)
	) name10123 (
		_w20413_,
		_w20414_,
		_w20635_
	);
	LUT2 #(
		.INIT('h1)
	) name10124 (
		_w20415_,
		_w20416_,
		_w20636_
	);
	LUT2 #(
		.INIT('h1)
	) name10125 (
		_w20417_,
		_w20418_,
		_w20637_
	);
	LUT2 #(
		.INIT('h1)
	) name10126 (
		_w20419_,
		_w20420_,
		_w20638_
	);
	LUT2 #(
		.INIT('h1)
	) name10127 (
		_w20421_,
		_w20422_,
		_w20639_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w20423_,
		_w20424_,
		_w20640_
	);
	LUT2 #(
		.INIT('h1)
	) name10129 (
		_w20425_,
		_w20426_,
		_w20641_
	);
	LUT2 #(
		.INIT('h1)
	) name10130 (
		_w20427_,
		_w20428_,
		_w20642_
	);
	LUT2 #(
		.INIT('h1)
	) name10131 (
		_w20429_,
		_w20430_,
		_w20643_
	);
	LUT2 #(
		.INIT('h1)
	) name10132 (
		_w20431_,
		_w20432_,
		_w20644_
	);
	LUT2 #(
		.INIT('h1)
	) name10133 (
		_w20433_,
		_w20434_,
		_w20645_
	);
	LUT2 #(
		.INIT('h1)
	) name10134 (
		_w20435_,
		_w20436_,
		_w20646_
	);
	LUT2 #(
		.INIT('h1)
	) name10135 (
		_w20437_,
		_w20438_,
		_w20647_
	);
	LUT2 #(
		.INIT('h1)
	) name10136 (
		_w20439_,
		_w20440_,
		_w20648_
	);
	LUT2 #(
		.INIT('h1)
	) name10137 (
		_w20441_,
		_w20442_,
		_w20649_
	);
	LUT2 #(
		.INIT('h1)
	) name10138 (
		_w20443_,
		_w20444_,
		_w20650_
	);
	LUT2 #(
		.INIT('h1)
	) name10139 (
		_w20445_,
		_w20446_,
		_w20651_
	);
	LUT2 #(
		.INIT('h1)
	) name10140 (
		_w20447_,
		_w20448_,
		_w20652_
	);
	LUT2 #(
		.INIT('h1)
	) name10141 (
		_w20449_,
		_w20450_,
		_w20653_
	);
	LUT2 #(
		.INIT('h1)
	) name10142 (
		_w20451_,
		_w20452_,
		_w20654_
	);
	LUT2 #(
		.INIT('h1)
	) name10143 (
		_w20453_,
		_w20454_,
		_w20655_
	);
	LUT2 #(
		.INIT('h1)
	) name10144 (
		_w20455_,
		_w20456_,
		_w20656_
	);
	LUT2 #(
		.INIT('h1)
	) name10145 (
		_w20457_,
		_w20458_,
		_w20657_
	);
	LUT2 #(
		.INIT('h1)
	) name10146 (
		_w20459_,
		_w20460_,
		_w20658_
	);
	LUT2 #(
		.INIT('h1)
	) name10147 (
		_w20461_,
		_w20462_,
		_w20659_
	);
	LUT2 #(
		.INIT('h1)
	) name10148 (
		_w20463_,
		_w20464_,
		_w20660_
	);
	LUT2 #(
		.INIT('h1)
	) name10149 (
		_w20465_,
		_w20466_,
		_w20661_
	);
	LUT2 #(
		.INIT('h1)
	) name10150 (
		_w20467_,
		_w20468_,
		_w20662_
	);
	LUT2 #(
		.INIT('h1)
	) name10151 (
		_w20469_,
		_w20470_,
		_w20663_
	);
	LUT2 #(
		.INIT('h1)
	) name10152 (
		_w20471_,
		_w20472_,
		_w20664_
	);
	LUT2 #(
		.INIT('h1)
	) name10153 (
		_w20473_,
		_w20474_,
		_w20665_
	);
	LUT2 #(
		.INIT('h1)
	) name10154 (
		_w20475_,
		_w20476_,
		_w20666_
	);
	LUT2 #(
		.INIT('h1)
	) name10155 (
		_w20477_,
		_w20478_,
		_w20667_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w20479_,
		_w20480_,
		_w20668_
	);
	LUT2 #(
		.INIT('h1)
	) name10157 (
		_w20481_,
		_w20482_,
		_w20669_
	);
	LUT2 #(
		.INIT('h1)
	) name10158 (
		_w20483_,
		_w20484_,
		_w20670_
	);
	LUT2 #(
		.INIT('h1)
	) name10159 (
		_w20485_,
		_w20486_,
		_w20671_
	);
	LUT2 #(
		.INIT('h1)
	) name10160 (
		_w20487_,
		_w20488_,
		_w20672_
	);
	LUT2 #(
		.INIT('h1)
	) name10161 (
		_w20489_,
		_w20490_,
		_w20673_
	);
	LUT2 #(
		.INIT('h1)
	) name10162 (
		_w20491_,
		_w20492_,
		_w20674_
	);
	LUT2 #(
		.INIT('h1)
	) name10163 (
		_w20493_,
		_w20494_,
		_w20675_
	);
	LUT2 #(
		.INIT('h1)
	) name10164 (
		_w20495_,
		_w20496_,
		_w20676_
	);
	LUT2 #(
		.INIT('h1)
	) name10165 (
		_w20497_,
		_w20498_,
		_w20677_
	);
	LUT2 #(
		.INIT('h1)
	) name10166 (
		_w20499_,
		_w20500_,
		_w20678_
	);
	LUT2 #(
		.INIT('h1)
	) name10167 (
		_w20501_,
		_w20502_,
		_w20679_
	);
	LUT2 #(
		.INIT('h1)
	) name10168 (
		_w20503_,
		_w20504_,
		_w20680_
	);
	LUT2 #(
		.INIT('h1)
	) name10169 (
		_w20505_,
		_w20506_,
		_w20681_
	);
	LUT2 #(
		.INIT('h1)
	) name10170 (
		_w20507_,
		_w20508_,
		_w20682_
	);
	LUT2 #(
		.INIT('h1)
	) name10171 (
		_w20509_,
		_w20510_,
		_w20683_
	);
	LUT2 #(
		.INIT('h1)
	) name10172 (
		_w20511_,
		_w20512_,
		_w20684_
	);
	LUT2 #(
		.INIT('h1)
	) name10173 (
		_w20513_,
		_w20514_,
		_w20685_
	);
	LUT2 #(
		.INIT('h1)
	) name10174 (
		_w20515_,
		_w20516_,
		_w20686_
	);
	LUT2 #(
		.INIT('h1)
	) name10175 (
		_w20517_,
		_w20518_,
		_w20687_
	);
	LUT2 #(
		.INIT('h1)
	) name10176 (
		_w20519_,
		_w20520_,
		_w20688_
	);
	LUT2 #(
		.INIT('h1)
	) name10177 (
		_w20521_,
		_w20522_,
		_w20689_
	);
	LUT2 #(
		.INIT('h1)
	) name10178 (
		_w20523_,
		_w20524_,
		_w20690_
	);
	LUT2 #(
		.INIT('h1)
	) name10179 (
		_w20525_,
		_w20526_,
		_w20691_
	);
	LUT2 #(
		.INIT('h1)
	) name10180 (
		_w20527_,
		_w20528_,
		_w20692_
	);
	LUT2 #(
		.INIT('h1)
	) name10181 (
		_w20529_,
		_w20530_,
		_w20693_
	);
	LUT2 #(
		.INIT('h1)
	) name10182 (
		_w20531_,
		_w20532_,
		_w20694_
	);
	LUT2 #(
		.INIT('h1)
	) name10183 (
		_w20533_,
		_w20534_,
		_w20695_
	);
	LUT2 #(
		.INIT('h1)
	) name10184 (
		_w20535_,
		_w20536_,
		_w20696_
	);
	LUT2 #(
		.INIT('h1)
	) name10185 (
		_w20537_,
		_w20538_,
		_w20697_
	);
	LUT2 #(
		.INIT('h1)
	) name10186 (
		_w20539_,
		_w20540_,
		_w20698_
	);
	LUT2 #(
		.INIT('h1)
	) name10187 (
		_w20541_,
		_w20542_,
		_w20699_
	);
	LUT2 #(
		.INIT('h1)
	) name10188 (
		_w20543_,
		_w20544_,
		_w20700_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		_w20545_,
		_w20546_,
		_w20701_
	);
	LUT2 #(
		.INIT('h1)
	) name10190 (
		_w20547_,
		_w20548_,
		_w20702_
	);
	LUT2 #(
		.INIT('h1)
	) name10191 (
		_w20549_,
		_w20550_,
		_w20703_
	);
	LUT2 #(
		.INIT('h1)
	) name10192 (
		_w20551_,
		_w20552_,
		_w20704_
	);
	LUT2 #(
		.INIT('h1)
	) name10193 (
		_w20553_,
		_w20554_,
		_w20705_
	);
	LUT2 #(
		.INIT('h1)
	) name10194 (
		_w20555_,
		_w20556_,
		_w20706_
	);
	LUT2 #(
		.INIT('h1)
	) name10195 (
		_w20557_,
		_w20558_,
		_w20707_
	);
	LUT2 #(
		.INIT('h1)
	) name10196 (
		_w20559_,
		_w20560_,
		_w20708_
	);
	LUT2 #(
		.INIT('h1)
	) name10197 (
		_w20561_,
		_w20562_,
		_w20709_
	);
	LUT2 #(
		.INIT('h1)
	) name10198 (
		_w20563_,
		_w20564_,
		_w20710_
	);
	LUT2 #(
		.INIT('h1)
	) name10199 (
		_w20565_,
		_w20566_,
		_w20711_
	);
	LUT2 #(
		.INIT('h1)
	) name10200 (
		_w20567_,
		_w20568_,
		_w20712_
	);
	LUT2 #(
		.INIT('h1)
	) name10201 (
		_w20569_,
		_w20570_,
		_w20713_
	);
	LUT2 #(
		.INIT('h1)
	) name10202 (
		_w20571_,
		_w20572_,
		_w20714_
	);
	LUT2 #(
		.INIT('h1)
	) name10203 (
		_w20573_,
		_w20574_,
		_w20715_
	);
	LUT2 #(
		.INIT('h1)
	) name10204 (
		_w20575_,
		_w20576_,
		_w20716_
	);
	LUT2 #(
		.INIT('h1)
	) name10205 (
		_w20577_,
		_w20578_,
		_w20717_
	);
	LUT2 #(
		.INIT('h1)
	) name10206 (
		_w20579_,
		_w20580_,
		_w20718_
	);
	LUT2 #(
		.INIT('h1)
	) name10207 (
		_w20581_,
		_w20582_,
		_w20719_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w20583_,
		_w20584_,
		_w20720_
	);
	LUT2 #(
		.INIT('h1)
	) name10209 (
		_w20585_,
		_w20586_,
		_w20721_
	);
	LUT2 #(
		.INIT('h1)
	) name10210 (
		_w20587_,
		_w20588_,
		_w20722_
	);
	LUT2 #(
		.INIT('h1)
	) name10211 (
		_w20589_,
		_w20590_,
		_w20723_
	);
	LUT2 #(
		.INIT('h1)
	) name10212 (
		_w20591_,
		_w20592_,
		_w20724_
	);
	LUT2 #(
		.INIT('h1)
	) name10213 (
		_w20593_,
		_w20594_,
		_w20725_
	);
	LUT2 #(
		.INIT('h1)
	) name10214 (
		_w20595_,
		_w20596_,
		_w20726_
	);
	LUT2 #(
		.INIT('h1)
	) name10215 (
		_w20597_,
		_w20598_,
		_w20727_
	);
	LUT2 #(
		.INIT('h1)
	) name10216 (
		_w20599_,
		_w20600_,
		_w20728_
	);
	LUT2 #(
		.INIT('h8)
	) name10217 (
		_w20727_,
		_w20728_,
		_w20729_
	);
	LUT2 #(
		.INIT('h8)
	) name10218 (
		_w20725_,
		_w20726_,
		_w20730_
	);
	LUT2 #(
		.INIT('h8)
	) name10219 (
		_w20723_,
		_w20724_,
		_w20731_
	);
	LUT2 #(
		.INIT('h8)
	) name10220 (
		_w20721_,
		_w20722_,
		_w20732_
	);
	LUT2 #(
		.INIT('h8)
	) name10221 (
		_w20719_,
		_w20720_,
		_w20733_
	);
	LUT2 #(
		.INIT('h8)
	) name10222 (
		_w20717_,
		_w20718_,
		_w20734_
	);
	LUT2 #(
		.INIT('h8)
	) name10223 (
		_w20715_,
		_w20716_,
		_w20735_
	);
	LUT2 #(
		.INIT('h8)
	) name10224 (
		_w20713_,
		_w20714_,
		_w20736_
	);
	LUT2 #(
		.INIT('h8)
	) name10225 (
		_w20711_,
		_w20712_,
		_w20737_
	);
	LUT2 #(
		.INIT('h8)
	) name10226 (
		_w20709_,
		_w20710_,
		_w20738_
	);
	LUT2 #(
		.INIT('h8)
	) name10227 (
		_w20707_,
		_w20708_,
		_w20739_
	);
	LUT2 #(
		.INIT('h8)
	) name10228 (
		_w20705_,
		_w20706_,
		_w20740_
	);
	LUT2 #(
		.INIT('h8)
	) name10229 (
		_w20703_,
		_w20704_,
		_w20741_
	);
	LUT2 #(
		.INIT('h8)
	) name10230 (
		_w20701_,
		_w20702_,
		_w20742_
	);
	LUT2 #(
		.INIT('h8)
	) name10231 (
		_w20699_,
		_w20700_,
		_w20743_
	);
	LUT2 #(
		.INIT('h8)
	) name10232 (
		_w20697_,
		_w20698_,
		_w20744_
	);
	LUT2 #(
		.INIT('h8)
	) name10233 (
		_w20695_,
		_w20696_,
		_w20745_
	);
	LUT2 #(
		.INIT('h8)
	) name10234 (
		_w20693_,
		_w20694_,
		_w20746_
	);
	LUT2 #(
		.INIT('h8)
	) name10235 (
		_w20691_,
		_w20692_,
		_w20747_
	);
	LUT2 #(
		.INIT('h8)
	) name10236 (
		_w20689_,
		_w20690_,
		_w20748_
	);
	LUT2 #(
		.INIT('h8)
	) name10237 (
		_w20687_,
		_w20688_,
		_w20749_
	);
	LUT2 #(
		.INIT('h8)
	) name10238 (
		_w20685_,
		_w20686_,
		_w20750_
	);
	LUT2 #(
		.INIT('h8)
	) name10239 (
		_w20683_,
		_w20684_,
		_w20751_
	);
	LUT2 #(
		.INIT('h8)
	) name10240 (
		_w20681_,
		_w20682_,
		_w20752_
	);
	LUT2 #(
		.INIT('h8)
	) name10241 (
		_w20679_,
		_w20680_,
		_w20753_
	);
	LUT2 #(
		.INIT('h8)
	) name10242 (
		_w20677_,
		_w20678_,
		_w20754_
	);
	LUT2 #(
		.INIT('h8)
	) name10243 (
		_w20675_,
		_w20676_,
		_w20755_
	);
	LUT2 #(
		.INIT('h8)
	) name10244 (
		_w20673_,
		_w20674_,
		_w20756_
	);
	LUT2 #(
		.INIT('h8)
	) name10245 (
		_w20671_,
		_w20672_,
		_w20757_
	);
	LUT2 #(
		.INIT('h8)
	) name10246 (
		_w20669_,
		_w20670_,
		_w20758_
	);
	LUT2 #(
		.INIT('h8)
	) name10247 (
		_w20667_,
		_w20668_,
		_w20759_
	);
	LUT2 #(
		.INIT('h8)
	) name10248 (
		_w20665_,
		_w20666_,
		_w20760_
	);
	LUT2 #(
		.INIT('h8)
	) name10249 (
		_w20663_,
		_w20664_,
		_w20761_
	);
	LUT2 #(
		.INIT('h8)
	) name10250 (
		_w20661_,
		_w20662_,
		_w20762_
	);
	LUT2 #(
		.INIT('h8)
	) name10251 (
		_w20659_,
		_w20660_,
		_w20763_
	);
	LUT2 #(
		.INIT('h8)
	) name10252 (
		_w20657_,
		_w20658_,
		_w20764_
	);
	LUT2 #(
		.INIT('h8)
	) name10253 (
		_w20655_,
		_w20656_,
		_w20765_
	);
	LUT2 #(
		.INIT('h8)
	) name10254 (
		_w20653_,
		_w20654_,
		_w20766_
	);
	LUT2 #(
		.INIT('h8)
	) name10255 (
		_w20651_,
		_w20652_,
		_w20767_
	);
	LUT2 #(
		.INIT('h8)
	) name10256 (
		_w20649_,
		_w20650_,
		_w20768_
	);
	LUT2 #(
		.INIT('h8)
	) name10257 (
		_w20647_,
		_w20648_,
		_w20769_
	);
	LUT2 #(
		.INIT('h8)
	) name10258 (
		_w20645_,
		_w20646_,
		_w20770_
	);
	LUT2 #(
		.INIT('h8)
	) name10259 (
		_w20643_,
		_w20644_,
		_w20771_
	);
	LUT2 #(
		.INIT('h8)
	) name10260 (
		_w20641_,
		_w20642_,
		_w20772_
	);
	LUT2 #(
		.INIT('h8)
	) name10261 (
		_w20639_,
		_w20640_,
		_w20773_
	);
	LUT2 #(
		.INIT('h8)
	) name10262 (
		_w20637_,
		_w20638_,
		_w20774_
	);
	LUT2 #(
		.INIT('h8)
	) name10263 (
		_w20635_,
		_w20636_,
		_w20775_
	);
	LUT2 #(
		.INIT('h8)
	) name10264 (
		_w20633_,
		_w20634_,
		_w20776_
	);
	LUT2 #(
		.INIT('h8)
	) name10265 (
		_w20631_,
		_w20632_,
		_w20777_
	);
	LUT2 #(
		.INIT('h8)
	) name10266 (
		_w20629_,
		_w20630_,
		_w20778_
	);
	LUT2 #(
		.INIT('h8)
	) name10267 (
		_w20627_,
		_w20628_,
		_w20779_
	);
	LUT2 #(
		.INIT('h8)
	) name10268 (
		_w20625_,
		_w20626_,
		_w20780_
	);
	LUT2 #(
		.INIT('h8)
	) name10269 (
		_w20623_,
		_w20624_,
		_w20781_
	);
	LUT2 #(
		.INIT('h8)
	) name10270 (
		_w20621_,
		_w20622_,
		_w20782_
	);
	LUT2 #(
		.INIT('h8)
	) name10271 (
		_w20619_,
		_w20620_,
		_w20783_
	);
	LUT2 #(
		.INIT('h8)
	) name10272 (
		_w20617_,
		_w20618_,
		_w20784_
	);
	LUT2 #(
		.INIT('h8)
	) name10273 (
		_w20615_,
		_w20616_,
		_w20785_
	);
	LUT2 #(
		.INIT('h8)
	) name10274 (
		_w20613_,
		_w20614_,
		_w20786_
	);
	LUT2 #(
		.INIT('h8)
	) name10275 (
		_w20611_,
		_w20612_,
		_w20787_
	);
	LUT2 #(
		.INIT('h8)
	) name10276 (
		_w20609_,
		_w20610_,
		_w20788_
	);
	LUT2 #(
		.INIT('h8)
	) name10277 (
		_w20607_,
		_w20608_,
		_w20789_
	);
	LUT2 #(
		.INIT('h8)
	) name10278 (
		_w20605_,
		_w20606_,
		_w20790_
	);
	LUT2 #(
		.INIT('h8)
	) name10279 (
		_w20603_,
		_w20604_,
		_w20791_
	);
	LUT2 #(
		.INIT('h8)
	) name10280 (
		_w20601_,
		_w20602_,
		_w20792_
	);
	LUT2 #(
		.INIT('h8)
	) name10281 (
		_w20791_,
		_w20792_,
		_w20793_
	);
	LUT2 #(
		.INIT('h8)
	) name10282 (
		_w20789_,
		_w20790_,
		_w20794_
	);
	LUT2 #(
		.INIT('h8)
	) name10283 (
		_w20787_,
		_w20788_,
		_w20795_
	);
	LUT2 #(
		.INIT('h8)
	) name10284 (
		_w20785_,
		_w20786_,
		_w20796_
	);
	LUT2 #(
		.INIT('h8)
	) name10285 (
		_w20783_,
		_w20784_,
		_w20797_
	);
	LUT2 #(
		.INIT('h8)
	) name10286 (
		_w20781_,
		_w20782_,
		_w20798_
	);
	LUT2 #(
		.INIT('h8)
	) name10287 (
		_w20779_,
		_w20780_,
		_w20799_
	);
	LUT2 #(
		.INIT('h8)
	) name10288 (
		_w20777_,
		_w20778_,
		_w20800_
	);
	LUT2 #(
		.INIT('h8)
	) name10289 (
		_w20775_,
		_w20776_,
		_w20801_
	);
	LUT2 #(
		.INIT('h8)
	) name10290 (
		_w20773_,
		_w20774_,
		_w20802_
	);
	LUT2 #(
		.INIT('h8)
	) name10291 (
		_w20771_,
		_w20772_,
		_w20803_
	);
	LUT2 #(
		.INIT('h8)
	) name10292 (
		_w20769_,
		_w20770_,
		_w20804_
	);
	LUT2 #(
		.INIT('h8)
	) name10293 (
		_w20767_,
		_w20768_,
		_w20805_
	);
	LUT2 #(
		.INIT('h8)
	) name10294 (
		_w20765_,
		_w20766_,
		_w20806_
	);
	LUT2 #(
		.INIT('h8)
	) name10295 (
		_w20763_,
		_w20764_,
		_w20807_
	);
	LUT2 #(
		.INIT('h8)
	) name10296 (
		_w20761_,
		_w20762_,
		_w20808_
	);
	LUT2 #(
		.INIT('h8)
	) name10297 (
		_w20759_,
		_w20760_,
		_w20809_
	);
	LUT2 #(
		.INIT('h8)
	) name10298 (
		_w20757_,
		_w20758_,
		_w20810_
	);
	LUT2 #(
		.INIT('h8)
	) name10299 (
		_w20755_,
		_w20756_,
		_w20811_
	);
	LUT2 #(
		.INIT('h8)
	) name10300 (
		_w20753_,
		_w20754_,
		_w20812_
	);
	LUT2 #(
		.INIT('h8)
	) name10301 (
		_w20751_,
		_w20752_,
		_w20813_
	);
	LUT2 #(
		.INIT('h8)
	) name10302 (
		_w20749_,
		_w20750_,
		_w20814_
	);
	LUT2 #(
		.INIT('h8)
	) name10303 (
		_w20747_,
		_w20748_,
		_w20815_
	);
	LUT2 #(
		.INIT('h8)
	) name10304 (
		_w20745_,
		_w20746_,
		_w20816_
	);
	LUT2 #(
		.INIT('h8)
	) name10305 (
		_w20743_,
		_w20744_,
		_w20817_
	);
	LUT2 #(
		.INIT('h8)
	) name10306 (
		_w20741_,
		_w20742_,
		_w20818_
	);
	LUT2 #(
		.INIT('h8)
	) name10307 (
		_w20739_,
		_w20740_,
		_w20819_
	);
	LUT2 #(
		.INIT('h8)
	) name10308 (
		_w20737_,
		_w20738_,
		_w20820_
	);
	LUT2 #(
		.INIT('h8)
	) name10309 (
		_w20735_,
		_w20736_,
		_w20821_
	);
	LUT2 #(
		.INIT('h8)
	) name10310 (
		_w20733_,
		_w20734_,
		_w20822_
	);
	LUT2 #(
		.INIT('h8)
	) name10311 (
		_w20731_,
		_w20732_,
		_w20823_
	);
	LUT2 #(
		.INIT('h8)
	) name10312 (
		_w20729_,
		_w20730_,
		_w20824_
	);
	LUT2 #(
		.INIT('h8)
	) name10313 (
		_w20823_,
		_w20824_,
		_w20825_
	);
	LUT2 #(
		.INIT('h8)
	) name10314 (
		_w20821_,
		_w20822_,
		_w20826_
	);
	LUT2 #(
		.INIT('h8)
	) name10315 (
		_w20819_,
		_w20820_,
		_w20827_
	);
	LUT2 #(
		.INIT('h8)
	) name10316 (
		_w20817_,
		_w20818_,
		_w20828_
	);
	LUT2 #(
		.INIT('h8)
	) name10317 (
		_w20815_,
		_w20816_,
		_w20829_
	);
	LUT2 #(
		.INIT('h8)
	) name10318 (
		_w20813_,
		_w20814_,
		_w20830_
	);
	LUT2 #(
		.INIT('h8)
	) name10319 (
		_w20811_,
		_w20812_,
		_w20831_
	);
	LUT2 #(
		.INIT('h8)
	) name10320 (
		_w20809_,
		_w20810_,
		_w20832_
	);
	LUT2 #(
		.INIT('h8)
	) name10321 (
		_w20807_,
		_w20808_,
		_w20833_
	);
	LUT2 #(
		.INIT('h8)
	) name10322 (
		_w20805_,
		_w20806_,
		_w20834_
	);
	LUT2 #(
		.INIT('h8)
	) name10323 (
		_w20803_,
		_w20804_,
		_w20835_
	);
	LUT2 #(
		.INIT('h8)
	) name10324 (
		_w20801_,
		_w20802_,
		_w20836_
	);
	LUT2 #(
		.INIT('h8)
	) name10325 (
		_w20799_,
		_w20800_,
		_w20837_
	);
	LUT2 #(
		.INIT('h8)
	) name10326 (
		_w20797_,
		_w20798_,
		_w20838_
	);
	LUT2 #(
		.INIT('h8)
	) name10327 (
		_w20795_,
		_w20796_,
		_w20839_
	);
	LUT2 #(
		.INIT('h8)
	) name10328 (
		_w20793_,
		_w20794_,
		_w20840_
	);
	LUT2 #(
		.INIT('h8)
	) name10329 (
		_w20839_,
		_w20840_,
		_w20841_
	);
	LUT2 #(
		.INIT('h8)
	) name10330 (
		_w20837_,
		_w20838_,
		_w20842_
	);
	LUT2 #(
		.INIT('h8)
	) name10331 (
		_w20835_,
		_w20836_,
		_w20843_
	);
	LUT2 #(
		.INIT('h8)
	) name10332 (
		_w20833_,
		_w20834_,
		_w20844_
	);
	LUT2 #(
		.INIT('h8)
	) name10333 (
		_w20831_,
		_w20832_,
		_w20845_
	);
	LUT2 #(
		.INIT('h8)
	) name10334 (
		_w20829_,
		_w20830_,
		_w20846_
	);
	LUT2 #(
		.INIT('h8)
	) name10335 (
		_w20827_,
		_w20828_,
		_w20847_
	);
	LUT2 #(
		.INIT('h8)
	) name10336 (
		_w20825_,
		_w20826_,
		_w20848_
	);
	LUT2 #(
		.INIT('h8)
	) name10337 (
		_w20847_,
		_w20848_,
		_w20849_
	);
	LUT2 #(
		.INIT('h8)
	) name10338 (
		_w20845_,
		_w20846_,
		_w20850_
	);
	LUT2 #(
		.INIT('h8)
	) name10339 (
		_w20843_,
		_w20844_,
		_w20851_
	);
	LUT2 #(
		.INIT('h8)
	) name10340 (
		_w20841_,
		_w20842_,
		_w20852_
	);
	LUT2 #(
		.INIT('h8)
	) name10341 (
		_w20851_,
		_w20852_,
		_w20853_
	);
	LUT2 #(
		.INIT('h8)
	) name10342 (
		_w20849_,
		_w20850_,
		_w20854_
	);
	LUT2 #(
		.INIT('h8)
	) name10343 (
		_w20853_,
		_w20854_,
		_w20855_
	);
	LUT2 #(
		.INIT('h1)
	) name10344 (
		wb_rst_i_pad,
		_w20855_,
		_w20856_
	);
	LUT2 #(
		.INIT('h8)
	) name10345 (
		_w12656_,
		_w20856_,
		_w20857_
	);
	LUT2 #(
		.INIT('h1)
	) name10346 (
		_w20344_,
		_w20857_,
		_w20858_
	);
	LUT2 #(
		.INIT('h2)
	) name10347 (
		\wishbone_LatchedTxLength_reg[12]/NET0131 ,
		_w12656_,
		_w20859_
	);
	LUT2 #(
		.INIT('h1)
	) name10348 (
		_w13476_,
		_w20859_,
		_w20860_
	);
	LUT2 #(
		.INIT('h2)
	) name10349 (
		\wishbone_LatchedTxLength_reg[13]/NET0131 ,
		_w12656_,
		_w20861_
	);
	LUT2 #(
		.INIT('h1)
	) name10350 (
		_w14020_,
		_w20861_,
		_w20862_
	);
	LUT2 #(
		.INIT('h2)
	) name10351 (
		\wishbone_LatchedTxLength_reg[14]/NET0131 ,
		_w12656_,
		_w20863_
	);
	LUT2 #(
		.INIT('h1)
	) name10352 (
		_w14537_,
		_w20863_,
		_w20864_
	);
	LUT2 #(
		.INIT('h1)
	) name10353 (
		\wishbone_LatchedTxLength_reg[15]/NET0131 ,
		_w12656_,
		_w20865_
	);
	LUT2 #(
		.INIT('h1)
	) name10354 (
		_w19605_,
		_w20865_,
		_w20866_
	);
	LUT2 #(
		.INIT('h2)
	) name10355 (
		\wishbone_LatchedTxLength_reg[1]/NET0131 ,
		_w12656_,
		_w20867_
	);
	LUT2 #(
		.INIT('h1)
	) name10356 (
		_w20127_,
		_w20867_,
		_w20868_
	);
	LUT2 #(
		.INIT('h2)
	) name10357 (
		\wishbone_LatchedTxLength_reg[2]/NET0131 ,
		_w12656_,
		_w20869_
	);
	LUT2 #(
		.INIT('h1)
	) name10358 (
		_w18565_,
		_w20869_,
		_w20870_
	);
	LUT2 #(
		.INIT('h2)
	) name10359 (
		\wishbone_LatchedTxLength_reg[3]/NET0131 ,
		_w12656_,
		_w20871_
	);
	LUT2 #(
		.INIT('h8)
	) name10360 (
		\wishbone_bd_ram_mem2_reg[96][19]/P0001 ,
		_w12912_,
		_w20872_
	);
	LUT2 #(
		.INIT('h8)
	) name10361 (
		\wishbone_bd_ram_mem2_reg[121][19]/P0001 ,
		_w13078_,
		_w20873_
	);
	LUT2 #(
		.INIT('h8)
	) name10362 (
		\wishbone_bd_ram_mem2_reg[191][19]/P0001 ,
		_w13034_,
		_w20874_
	);
	LUT2 #(
		.INIT('h8)
	) name10363 (
		\wishbone_bd_ram_mem2_reg[98][19]/P0001 ,
		_w12816_,
		_w20875_
	);
	LUT2 #(
		.INIT('h8)
	) name10364 (
		\wishbone_bd_ram_mem2_reg[89][19]/P0001 ,
		_w12964_,
		_w20876_
	);
	LUT2 #(
		.INIT('h8)
	) name10365 (
		\wishbone_bd_ram_mem2_reg[72][19]/P0001 ,
		_w12810_,
		_w20877_
	);
	LUT2 #(
		.INIT('h8)
	) name10366 (
		\wishbone_bd_ram_mem2_reg[180][19]/P0001 ,
		_w12791_,
		_w20878_
	);
	LUT2 #(
		.INIT('h8)
	) name10367 (
		\wishbone_bd_ram_mem2_reg[248][19]/P0001 ,
		_w12789_,
		_w20879_
	);
	LUT2 #(
		.INIT('h8)
	) name10368 (
		\wishbone_bd_ram_mem2_reg[161][19]/P0001 ,
		_w12754_,
		_w20880_
	);
	LUT2 #(
		.INIT('h8)
	) name10369 (
		\wishbone_bd_ram_mem2_reg[31][19]/P0001 ,
		_w13198_,
		_w20881_
	);
	LUT2 #(
		.INIT('h8)
	) name10370 (
		\wishbone_bd_ram_mem2_reg[27][19]/P0001 ,
		_w12880_,
		_w20882_
	);
	LUT2 #(
		.INIT('h8)
	) name10371 (
		\wishbone_bd_ram_mem2_reg[210][19]/P0001 ,
		_w12924_,
		_w20883_
	);
	LUT2 #(
		.INIT('h8)
	) name10372 (
		\wishbone_bd_ram_mem2_reg[107][19]/P0001 ,
		_w12749_,
		_w20884_
	);
	LUT2 #(
		.INIT('h8)
	) name10373 (
		\wishbone_bd_ram_mem2_reg[54][19]/P0001 ,
		_w12770_,
		_w20885_
	);
	LUT2 #(
		.INIT('h8)
	) name10374 (
		\wishbone_bd_ram_mem2_reg[64][19]/P0001 ,
		_w12976_,
		_w20886_
	);
	LUT2 #(
		.INIT('h8)
	) name10375 (
		\wishbone_bd_ram_mem2_reg[158][19]/P0001 ,
		_w12898_,
		_w20887_
	);
	LUT2 #(
		.INIT('h8)
	) name10376 (
		\wishbone_bd_ram_mem2_reg[69][19]/P0001 ,
		_w12738_,
		_w20888_
	);
	LUT2 #(
		.INIT('h8)
	) name10377 (
		\wishbone_bd_ram_mem2_reg[87][19]/P0001 ,
		_w13154_,
		_w20889_
	);
	LUT2 #(
		.INIT('h8)
	) name10378 (
		\wishbone_bd_ram_mem2_reg[85][19]/P0001 ,
		_w13216_,
		_w20890_
	);
	LUT2 #(
		.INIT('h8)
	) name10379 (
		\wishbone_bd_ram_mem2_reg[235][19]/P0001 ,
		_w12696_,
		_w20891_
	);
	LUT2 #(
		.INIT('h8)
	) name10380 (
		\wishbone_bd_ram_mem2_reg[151][19]/P0001 ,
		_w13142_,
		_w20892_
	);
	LUT2 #(
		.INIT('h8)
	) name10381 (
		\wishbone_bd_ram_mem2_reg[92][19]/P0001 ,
		_w13010_,
		_w20893_
	);
	LUT2 #(
		.INIT('h8)
	) name10382 (
		\wishbone_bd_ram_mem2_reg[144][19]/P0001 ,
		_w12756_,
		_w20894_
	);
	LUT2 #(
		.INIT('h8)
	) name10383 (
		\wishbone_bd_ram_mem2_reg[5][19]/P0001 ,
		_w12878_,
		_w20895_
	);
	LUT2 #(
		.INIT('h8)
	) name10384 (
		\wishbone_bd_ram_mem2_reg[150][19]/P0001 ,
		_w13136_,
		_w20896_
	);
	LUT2 #(
		.INIT('h8)
	) name10385 (
		\wishbone_bd_ram_mem2_reg[143][19]/P0001 ,
		_w12922_,
		_w20897_
	);
	LUT2 #(
		.INIT('h8)
	) name10386 (
		\wishbone_bd_ram_mem2_reg[3][19]/P0001 ,
		_w12866_,
		_w20898_
	);
	LUT2 #(
		.INIT('h8)
	) name10387 (
		\wishbone_bd_ram_mem2_reg[227][19]/P0001 ,
		_w12936_,
		_w20899_
	);
	LUT2 #(
		.INIT('h8)
	) name10388 (
		\wishbone_bd_ram_mem2_reg[207][19]/P0001 ,
		_w13180_,
		_w20900_
	);
	LUT2 #(
		.INIT('h8)
	) name10389 (
		\wishbone_bd_ram_mem2_reg[132][19]/P0001 ,
		_w12992_,
		_w20901_
	);
	LUT2 #(
		.INIT('h8)
	) name10390 (
		\wishbone_bd_ram_mem2_reg[159][19]/P0001 ,
		_w12774_,
		_w20902_
	);
	LUT2 #(
		.INIT('h8)
	) name10391 (
		\wishbone_bd_ram_mem2_reg[16][19]/P0001 ,
		_w13140_,
		_w20903_
	);
	LUT2 #(
		.INIT('h8)
	) name10392 (
		\wishbone_bd_ram_mem2_reg[124][19]/P0001 ,
		_w13058_,
		_w20904_
	);
	LUT2 #(
		.INIT('h8)
	) name10393 (
		\wishbone_bd_ram_mem2_reg[28][19]/P0001 ,
		_w13170_,
		_w20905_
	);
	LUT2 #(
		.INIT('h8)
	) name10394 (
		\wishbone_bd_ram_mem2_reg[228][19]/P0001 ,
		_w12765_,
		_w20906_
	);
	LUT2 #(
		.INIT('h8)
	) name10395 (
		\wishbone_bd_ram_mem2_reg[100][19]/P0001 ,
		_w12960_,
		_w20907_
	);
	LUT2 #(
		.INIT('h8)
	) name10396 (
		\wishbone_bd_ram_mem2_reg[39][19]/P0001 ,
		_w13018_,
		_w20908_
	);
	LUT2 #(
		.INIT('h8)
	) name10397 (
		\wishbone_bd_ram_mem2_reg[63][19]/P0001 ,
		_w12850_,
		_w20909_
	);
	LUT2 #(
		.INIT('h8)
	) name10398 (
		\wishbone_bd_ram_mem2_reg[129][19]/P0001 ,
		_w12776_,
		_w20910_
	);
	LUT2 #(
		.INIT('h8)
	) name10399 (
		\wishbone_bd_ram_mem2_reg[201][19]/P0001 ,
		_w12822_,
		_w20911_
	);
	LUT2 #(
		.INIT('h8)
	) name10400 (
		\wishbone_bd_ram_mem2_reg[20][19]/P0001 ,
		_w13174_,
		_w20912_
	);
	LUT2 #(
		.INIT('h8)
	) name10401 (
		\wishbone_bd_ram_mem2_reg[163][19]/P0001 ,
		_w12882_,
		_w20913_
	);
	LUT2 #(
		.INIT('h8)
	) name10402 (
		\wishbone_bd_ram_mem2_reg[242][19]/P0001 ,
		_w12932_,
		_w20914_
	);
	LUT2 #(
		.INIT('h8)
	) name10403 (
		\wishbone_bd_ram_mem2_reg[60][19]/P0001 ,
		_w13204_,
		_w20915_
	);
	LUT2 #(
		.INIT('h8)
	) name10404 (
		\wishbone_bd_ram_mem2_reg[80][19]/P0001 ,
		_w12689_,
		_w20916_
	);
	LUT2 #(
		.INIT('h8)
	) name10405 (
		\wishbone_bd_ram_mem2_reg[169][19]/P0001 ,
		_w12722_,
		_w20917_
	);
	LUT2 #(
		.INIT('h8)
	) name10406 (
		\wishbone_bd_ram_mem2_reg[229][19]/P0001 ,
		_w12711_,
		_w20918_
	);
	LUT2 #(
		.INIT('h8)
	) name10407 (
		\wishbone_bd_ram_mem2_reg[25][19]/P0001 ,
		_w13108_,
		_w20919_
	);
	LUT2 #(
		.INIT('h8)
	) name10408 (
		\wishbone_bd_ram_mem2_reg[30][19]/P0001 ,
		_w13104_,
		_w20920_
	);
	LUT2 #(
		.INIT('h8)
	) name10409 (
		\wishbone_bd_ram_mem2_reg[36][19]/P0001 ,
		_w12800_,
		_w20921_
	);
	LUT2 #(
		.INIT('h8)
	) name10410 (
		\wishbone_bd_ram_mem2_reg[130][19]/P0001 ,
		_w12914_,
		_w20922_
	);
	LUT2 #(
		.INIT('h8)
	) name10411 (
		\wishbone_bd_ram_mem2_reg[236][19]/P0001 ,
		_w12731_,
		_w20923_
	);
	LUT2 #(
		.INIT('h8)
	) name10412 (
		\wishbone_bd_ram_mem2_reg[176][19]/P0001 ,
		_w12868_,
		_w20924_
	);
	LUT2 #(
		.INIT('h8)
	) name10413 (
		\wishbone_bd_ram_mem2_reg[208][19]/P0001 ,
		_w13032_,
		_w20925_
	);
	LUT2 #(
		.INIT('h8)
	) name10414 (
		\wishbone_bd_ram_mem2_reg[77][19]/P0001 ,
		_w12982_,
		_w20926_
	);
	LUT2 #(
		.INIT('h8)
	) name10415 (
		\wishbone_bd_ram_mem2_reg[182][19]/P0001 ,
		_w12820_,
		_w20927_
	);
	LUT2 #(
		.INIT('h8)
	) name10416 (
		\wishbone_bd_ram_mem2_reg[49][19]/P0001 ,
		_w12994_,
		_w20928_
	);
	LUT2 #(
		.INIT('h8)
	) name10417 (
		\wishbone_bd_ram_mem2_reg[7][19]/P0001 ,
		_w12728_,
		_w20929_
	);
	LUT2 #(
		.INIT('h8)
	) name10418 (
		\wishbone_bd_ram_mem2_reg[219][19]/P0001 ,
		_w12806_,
		_w20930_
	);
	LUT2 #(
		.INIT('h8)
	) name10419 (
		\wishbone_bd_ram_mem2_reg[245][19]/P0001 ,
		_w13022_,
		_w20931_
	);
	LUT2 #(
		.INIT('h8)
	) name10420 (
		\wishbone_bd_ram_mem2_reg[14][19]/P0001 ,
		_w13086_,
		_w20932_
	);
	LUT2 #(
		.INIT('h8)
	) name10421 (
		\wishbone_bd_ram_mem2_reg[38][19]/P0001 ,
		_w13182_,
		_w20933_
	);
	LUT2 #(
		.INIT('h8)
	) name10422 (
		\wishbone_bd_ram_mem2_reg[138][19]/P0001 ,
		_w12958_,
		_w20934_
	);
	LUT2 #(
		.INIT('h8)
	) name10423 (
		\wishbone_bd_ram_mem2_reg[13][19]/P0001 ,
		_w13178_,
		_w20935_
	);
	LUT2 #(
		.INIT('h8)
	) name10424 (
		\wishbone_bd_ram_mem2_reg[11][19]/P0001 ,
		_w13194_,
		_w20936_
	);
	LUT2 #(
		.INIT('h8)
	) name10425 (
		\wishbone_bd_ram_mem2_reg[18][19]/P0001 ,
		_w12679_,
		_w20937_
	);
	LUT2 #(
		.INIT('h8)
	) name10426 (
		\wishbone_bd_ram_mem2_reg[237][19]/P0001 ,
		_w12990_,
		_w20938_
	);
	LUT2 #(
		.INIT('h8)
	) name10427 (
		\wishbone_bd_ram_mem2_reg[135][19]/P0001 ,
		_w13124_,
		_w20939_
	);
	LUT2 #(
		.INIT('h8)
	) name10428 (
		\wishbone_bd_ram_mem2_reg[164][19]/P0001 ,
		_w12876_,
		_w20940_
	);
	LUT2 #(
		.INIT('h8)
	) name10429 (
		\wishbone_bd_ram_mem2_reg[56][19]/P0001 ,
		_w12778_,
		_w20941_
	);
	LUT2 #(
		.INIT('h8)
	) name10430 (
		\wishbone_bd_ram_mem2_reg[108][19]/P0001 ,
		_w13156_,
		_w20942_
	);
	LUT2 #(
		.INIT('h8)
	) name10431 (
		\wishbone_bd_ram_mem2_reg[217][19]/P0001 ,
		_w13188_,
		_w20943_
	);
	LUT2 #(
		.INIT('h8)
	) name10432 (
		\wishbone_bd_ram_mem2_reg[104][19]/P0001 ,
		_w13148_,
		_w20944_
	);
	LUT2 #(
		.INIT('h8)
	) name10433 (
		\wishbone_bd_ram_mem2_reg[156][19]/P0001 ,
		_w13190_,
		_w20945_
	);
	LUT2 #(
		.INIT('h8)
	) name10434 (
		\wishbone_bd_ram_mem2_reg[61][19]/P0001 ,
		_w12725_,
		_w20946_
	);
	LUT2 #(
		.INIT('h8)
	) name10435 (
		\wishbone_bd_ram_mem2_reg[109][19]/P0001 ,
		_w12888_,
		_w20947_
	);
	LUT2 #(
		.INIT('h8)
	) name10436 (
		\wishbone_bd_ram_mem2_reg[37][19]/P0001 ,
		_w13102_,
		_w20948_
	);
	LUT2 #(
		.INIT('h8)
	) name10437 (
		\wishbone_bd_ram_mem2_reg[55][19]/P0001 ,
		_w12785_,
		_w20949_
	);
	LUT2 #(
		.INIT('h8)
	) name10438 (
		\wishbone_bd_ram_mem2_reg[70][19]/P0001 ,
		_w12840_,
		_w20950_
	);
	LUT2 #(
		.INIT('h8)
	) name10439 (
		\wishbone_bd_ram_mem2_reg[170][19]/P0001 ,
		_w13030_,
		_w20951_
	);
	LUT2 #(
		.INIT('h8)
	) name10440 (
		\wishbone_bd_ram_mem2_reg[73][19]/P0001 ,
		_w12918_,
		_w20952_
	);
	LUT2 #(
		.INIT('h8)
	) name10441 (
		\wishbone_bd_ram_mem2_reg[187][19]/P0001 ,
		_w13196_,
		_w20953_
	);
	LUT2 #(
		.INIT('h8)
	) name10442 (
		\wishbone_bd_ram_mem2_reg[26][19]/P0001 ,
		_w12699_,
		_w20954_
	);
	LUT2 #(
		.INIT('h8)
	) name10443 (
		\wishbone_bd_ram_mem2_reg[67][19]/P0001 ,
		_w13134_,
		_w20955_
	);
	LUT2 #(
		.INIT('h8)
	) name10444 (
		\wishbone_bd_ram_mem2_reg[103][19]/P0001 ,
		_w12846_,
		_w20956_
	);
	LUT2 #(
		.INIT('h8)
	) name10445 (
		\wishbone_bd_ram_mem2_reg[223][19]/P0001 ,
		_w12838_,
		_w20957_
	);
	LUT2 #(
		.INIT('h8)
	) name10446 (
		\wishbone_bd_ram_mem2_reg[203][19]/P0001 ,
		_w13158_,
		_w20958_
	);
	LUT2 #(
		.INIT('h8)
	) name10447 (
		\wishbone_bd_ram_mem2_reg[181][19]/P0001 ,
		_w12828_,
		_w20959_
	);
	LUT2 #(
		.INIT('h8)
	) name10448 (
		\wishbone_bd_ram_mem2_reg[249][19]/P0001 ,
		_w12900_,
		_w20960_
	);
	LUT2 #(
		.INIT('h8)
	) name10449 (
		\wishbone_bd_ram_mem2_reg[32][19]/P0001 ,
		_w13120_,
		_w20961_
	);
	LUT2 #(
		.INIT('h8)
	) name10450 (
		\wishbone_bd_ram_mem2_reg[136][19]/P0001 ,
		_w13064_,
		_w20962_
	);
	LUT2 #(
		.INIT('h8)
	) name10451 (
		\wishbone_bd_ram_mem2_reg[118][19]/P0001 ,
		_w12830_,
		_w20963_
	);
	LUT2 #(
		.INIT('h8)
	) name10452 (
		\wishbone_bd_ram_mem2_reg[193][19]/P0001 ,
		_w13056_,
		_w20964_
	);
	LUT2 #(
		.INIT('h8)
	) name10453 (
		\wishbone_bd_ram_mem2_reg[42][19]/P0001 ,
		_w12842_,
		_w20965_
	);
	LUT2 #(
		.INIT('h8)
	) name10454 (
		\wishbone_bd_ram_mem2_reg[106][19]/P0001 ,
		_w12713_,
		_w20966_
	);
	LUT2 #(
		.INIT('h8)
	) name10455 (
		\wishbone_bd_ram_mem2_reg[15][19]/P0001 ,
		_w13210_,
		_w20967_
	);
	LUT2 #(
		.INIT('h8)
	) name10456 (
		\wishbone_bd_ram_mem2_reg[134][19]/P0001 ,
		_w12763_,
		_w20968_
	);
	LUT2 #(
		.INIT('h8)
	) name10457 (
		\wishbone_bd_ram_mem2_reg[62][19]/P0001 ,
		_w12673_,
		_w20969_
	);
	LUT2 #(
		.INIT('h8)
	) name10458 (
		\wishbone_bd_ram_mem2_reg[102][19]/P0001 ,
		_w12685_,
		_w20970_
	);
	LUT2 #(
		.INIT('h8)
	) name10459 (
		\wishbone_bd_ram_mem2_reg[126][19]/P0001 ,
		_w13218_,
		_w20971_
	);
	LUT2 #(
		.INIT('h8)
	) name10460 (
		\wishbone_bd_ram_mem2_reg[172][19]/P0001 ,
		_w12944_,
		_w20972_
	);
	LUT2 #(
		.INIT('h8)
	) name10461 (
		\wishbone_bd_ram_mem2_reg[212][19]/P0001 ,
		_w12796_,
		_w20973_
	);
	LUT2 #(
		.INIT('h8)
	) name10462 (
		\wishbone_bd_ram_mem2_reg[157][19]/P0001 ,
		_w12926_,
		_w20974_
	);
	LUT2 #(
		.INIT('h8)
	) name10463 (
		\wishbone_bd_ram_mem2_reg[183][19]/P0001 ,
		_w12787_,
		_w20975_
	);
	LUT2 #(
		.INIT('h8)
	) name10464 (
		\wishbone_bd_ram_mem2_reg[206][19]/P0001 ,
		_w12954_,
		_w20976_
	);
	LUT2 #(
		.INIT('h8)
	) name10465 (
		\wishbone_bd_ram_mem2_reg[215][19]/P0001 ,
		_w12974_,
		_w20977_
	);
	LUT2 #(
		.INIT('h8)
	) name10466 (
		\wishbone_bd_ram_mem2_reg[114][19]/P0001 ,
		_w13202_,
		_w20978_
	);
	LUT2 #(
		.INIT('h8)
	) name10467 (
		\wishbone_bd_ram_mem2_reg[119][19]/P0001 ,
		_w13048_,
		_w20979_
	);
	LUT2 #(
		.INIT('h8)
	) name10468 (
		\wishbone_bd_ram_mem2_reg[252][19]/P0001 ,
		_w13080_,
		_w20980_
	);
	LUT2 #(
		.INIT('h8)
	) name10469 (
		\wishbone_bd_ram_mem2_reg[21][19]/P0001 ,
		_w12906_,
		_w20981_
	);
	LUT2 #(
		.INIT('h8)
	) name10470 (
		\wishbone_bd_ram_mem2_reg[225][19]/P0001 ,
		_w13092_,
		_w20982_
	);
	LUT2 #(
		.INIT('h8)
	) name10471 (
		\wishbone_bd_ram_mem2_reg[205][19]/P0001 ,
		_w13068_,
		_w20983_
	);
	LUT2 #(
		.INIT('h8)
	) name10472 (
		\wishbone_bd_ram_mem2_reg[160][19]/P0001 ,
		_w12872_,
		_w20984_
	);
	LUT2 #(
		.INIT('h8)
	) name10473 (
		\wishbone_bd_ram_mem2_reg[148][19]/P0001 ,
		_w13000_,
		_w20985_
	);
	LUT2 #(
		.INIT('h8)
	) name10474 (
		\wishbone_bd_ram_mem2_reg[23][19]/P0001 ,
		_w13008_,
		_w20986_
	);
	LUT2 #(
		.INIT('h8)
	) name10475 (
		\wishbone_bd_ram_mem2_reg[131][19]/P0001 ,
		_w12852_,
		_w20987_
	);
	LUT2 #(
		.INIT('h8)
	) name10476 (
		\wishbone_bd_ram_mem2_reg[79][19]/P0001 ,
		_w13212_,
		_w20988_
	);
	LUT2 #(
		.INIT('h8)
	) name10477 (
		\wishbone_bd_ram_mem2_reg[91][19]/P0001 ,
		_w13074_,
		_w20989_
	);
	LUT2 #(
		.INIT('h8)
	) name10478 (
		\wishbone_bd_ram_mem2_reg[147][19]/P0001 ,
		_w13146_,
		_w20990_
	);
	LUT2 #(
		.INIT('h8)
	) name10479 (
		\wishbone_bd_ram_mem2_reg[113][19]/P0001 ,
		_w13026_,
		_w20991_
	);
	LUT2 #(
		.INIT('h8)
	) name10480 (
		\wishbone_bd_ram_mem2_reg[10][19]/P0001 ,
		_w13172_,
		_w20992_
	);
	LUT2 #(
		.INIT('h8)
	) name10481 (
		\wishbone_bd_ram_mem2_reg[74][19]/P0001 ,
		_w12812_,
		_w20993_
	);
	LUT2 #(
		.INIT('h8)
	) name10482 (
		\wishbone_bd_ram_mem2_reg[230][19]/P0001 ,
		_w13036_,
		_w20994_
	);
	LUT2 #(
		.INIT('h8)
	) name10483 (
		\wishbone_bd_ram_mem2_reg[6][19]/P0001 ,
		_w12968_,
		_w20995_
	);
	LUT2 #(
		.INIT('h8)
	) name10484 (
		\wishbone_bd_ram_mem2_reg[52][19]/P0001 ,
		_w13082_,
		_w20996_
	);
	LUT2 #(
		.INIT('h8)
	) name10485 (
		\wishbone_bd_ram_mem2_reg[190][19]/P0001 ,
		_w12858_,
		_w20997_
	);
	LUT2 #(
		.INIT('h8)
	) name10486 (
		\wishbone_bd_ram_mem2_reg[222][19]/P0001 ,
		_w13094_,
		_w20998_
	);
	LUT2 #(
		.INIT('h8)
	) name10487 (
		\wishbone_bd_ram_mem2_reg[122][19]/P0001 ,
		_w13130_,
		_w20999_
	);
	LUT2 #(
		.INIT('h8)
	) name10488 (
		\wishbone_bd_ram_mem2_reg[86][19]/P0001 ,
		_w12735_,
		_w21000_
	);
	LUT2 #(
		.INIT('h8)
	) name10489 (
		\wishbone_bd_ram_mem2_reg[137][19]/P0001 ,
		_w13168_,
		_w21001_
	);
	LUT2 #(
		.INIT('h8)
	) name10490 (
		\wishbone_bd_ram_mem2_reg[66][19]/P0001 ,
		_w12824_,
		_w21002_
	);
	LUT2 #(
		.INIT('h8)
	) name10491 (
		\wishbone_bd_ram_mem2_reg[221][19]/P0001 ,
		_w12802_,
		_w21003_
	);
	LUT2 #(
		.INIT('h8)
	) name10492 (
		\wishbone_bd_ram_mem2_reg[65][19]/P0001 ,
		_w13176_,
		_w21004_
	);
	LUT2 #(
		.INIT('h8)
	) name10493 (
		\wishbone_bd_ram_mem2_reg[234][19]/P0001 ,
		_w13214_,
		_w21005_
	);
	LUT2 #(
		.INIT('h8)
	) name10494 (
		\wishbone_bd_ram_mem2_reg[166][19]/P0001 ,
		_w13040_,
		_w21006_
	);
	LUT2 #(
		.INIT('h8)
	) name10495 (
		\wishbone_bd_ram_mem2_reg[78][19]/P0001 ,
		_w12874_,
		_w21007_
	);
	LUT2 #(
		.INIT('h8)
	) name10496 (
		\wishbone_bd_ram_mem2_reg[127][19]/P0001 ,
		_w13164_,
		_w21008_
	);
	LUT2 #(
		.INIT('h8)
	) name10497 (
		\wishbone_bd_ram_mem2_reg[244][19]/P0001 ,
		_w12747_,
		_w21009_
	);
	LUT2 #(
		.INIT('h8)
	) name10498 (
		\wishbone_bd_ram_mem2_reg[184][19]/P0001 ,
		_w13062_,
		_w21010_
	);
	LUT2 #(
		.INIT('h8)
	) name10499 (
		\wishbone_bd_ram_mem2_reg[117][19]/P0001 ,
		_w12715_,
		_w21011_
	);
	LUT2 #(
		.INIT('h8)
	) name10500 (
		\wishbone_bd_ram_mem2_reg[95][19]/P0001 ,
		_w12844_,
		_w21012_
	);
	LUT2 #(
		.INIT('h8)
	) name10501 (
		\wishbone_bd_ram_mem2_reg[99][19]/P0001 ,
		_w13038_,
		_w21013_
	);
	LUT2 #(
		.INIT('h8)
	) name10502 (
		\wishbone_bd_ram_mem2_reg[142][19]/P0001 ,
		_w12928_,
		_w21014_
	);
	LUT2 #(
		.INIT('h8)
	) name10503 (
		\wishbone_bd_ram_mem2_reg[153][19]/P0001 ,
		_w12890_,
		_w21015_
	);
	LUT2 #(
		.INIT('h8)
	) name10504 (
		\wishbone_bd_ram_mem2_reg[57][19]/P0001 ,
		_w13116_,
		_w21016_
	);
	LUT2 #(
		.INIT('h8)
	) name10505 (
		\wishbone_bd_ram_mem2_reg[232][19]/P0001 ,
		_w12758_,
		_w21017_
	);
	LUT2 #(
		.INIT('h8)
	) name10506 (
		\wishbone_bd_ram_mem2_reg[34][19]/P0001 ,
		_w12930_,
		_w21018_
	);
	LUT2 #(
		.INIT('h8)
	) name10507 (
		\wishbone_bd_ram_mem2_reg[82][19]/P0001 ,
		_w12942_,
		_w21019_
	);
	LUT2 #(
		.INIT('h8)
	) name10508 (
		\wishbone_bd_ram_mem2_reg[255][19]/P0001 ,
		_w13072_,
		_w21020_
	);
	LUT2 #(
		.INIT('h8)
	) name10509 (
		\wishbone_bd_ram_mem2_reg[155][19]/P0001 ,
		_w13122_,
		_w21021_
	);
	LUT2 #(
		.INIT('h8)
	) name10510 (
		\wishbone_bd_ram_mem2_reg[139][19]/P0001 ,
		_w12814_,
		_w21022_
	);
	LUT2 #(
		.INIT('h8)
	) name10511 (
		\wishbone_bd_ram_mem2_reg[250][19]/P0001 ,
		_w13128_,
		_w21023_
	);
	LUT2 #(
		.INIT('h8)
	) name10512 (
		\wishbone_bd_ram_mem2_reg[194][19]/P0001 ,
		_w12772_,
		_w21024_
	);
	LUT2 #(
		.INIT('h8)
	) name10513 (
		\wishbone_bd_ram_mem2_reg[44][19]/P0001 ,
		_w12896_,
		_w21025_
	);
	LUT2 #(
		.INIT('h8)
	) name10514 (
		\wishbone_bd_ram_mem2_reg[168][19]/P0001 ,
		_w13208_,
		_w21026_
	);
	LUT2 #(
		.INIT('h8)
	) name10515 (
		\wishbone_bd_ram_mem2_reg[209][19]/P0001 ,
		_w13152_,
		_w21027_
	);
	LUT2 #(
		.INIT('h8)
	) name10516 (
		\wishbone_bd_ram_mem2_reg[154][19]/P0001 ,
		_w12962_,
		_w21028_
	);
	LUT2 #(
		.INIT('h8)
	) name10517 (
		\wishbone_bd_ram_mem2_reg[76][19]/P0001 ,
		_w13184_,
		_w21029_
	);
	LUT2 #(
		.INIT('h8)
	) name10518 (
		\wishbone_bd_ram_mem2_reg[238][19]/P0001 ,
		_w13160_,
		_w21030_
	);
	LUT2 #(
		.INIT('h8)
	) name10519 (
		\wishbone_bd_ram_mem2_reg[8][19]/P0001 ,
		_w12920_,
		_w21031_
	);
	LUT2 #(
		.INIT('h8)
	) name10520 (
		\wishbone_bd_ram_mem2_reg[41][19]/P0001 ,
		_w13052_,
		_w21032_
	);
	LUT2 #(
		.INIT('h8)
	) name10521 (
		\wishbone_bd_ram_mem2_reg[33][19]/P0001 ,
		_w12980_,
		_w21033_
	);
	LUT2 #(
		.INIT('h8)
	) name10522 (
		\wishbone_bd_ram_mem2_reg[198][19]/P0001 ,
		_w12832_,
		_w21034_
	);
	LUT2 #(
		.INIT('h8)
	) name10523 (
		\wishbone_bd_ram_mem2_reg[0][19]/P0001 ,
		_w12717_,
		_w21035_
	);
	LUT2 #(
		.INIT('h8)
	) name10524 (
		\wishbone_bd_ram_mem2_reg[199][19]/P0001 ,
		_w12768_,
		_w21036_
	);
	LUT2 #(
		.INIT('h8)
	) name10525 (
		\wishbone_bd_ram_mem2_reg[71][19]/P0001 ,
		_w12798_,
		_w21037_
	);
	LUT2 #(
		.INIT('h8)
	) name10526 (
		\wishbone_bd_ram_mem2_reg[47][19]/P0001 ,
		_w12904_,
		_w21038_
	);
	LUT2 #(
		.INIT('h8)
	) name10527 (
		\wishbone_bd_ram_mem2_reg[29][19]/P0001 ,
		_w12952_,
		_w21039_
	);
	LUT2 #(
		.INIT('h8)
	) name10528 (
		\wishbone_bd_ram_mem2_reg[110][19]/P0001 ,
		_w13046_,
		_w21040_
	);
	LUT2 #(
		.INIT('h8)
	) name10529 (
		\wishbone_bd_ram_mem2_reg[59][19]/P0001 ,
		_w12780_,
		_w21041_
	);
	LUT2 #(
		.INIT('h8)
	) name10530 (
		\wishbone_bd_ram_mem2_reg[140][19]/P0001 ,
		_w12894_,
		_w21042_
	);
	LUT2 #(
		.INIT('h8)
	) name10531 (
		\wishbone_bd_ram_mem2_reg[9][19]/P0001 ,
		_w12808_,
		_w21043_
	);
	LUT2 #(
		.INIT('h8)
	) name10532 (
		\wishbone_bd_ram_mem2_reg[178][19]/P0001 ,
		_w12886_,
		_w21044_
	);
	LUT2 #(
		.INIT('h8)
	) name10533 (
		\wishbone_bd_ram_mem2_reg[75][19]/P0001 ,
		_w12826_,
		_w21045_
	);
	LUT2 #(
		.INIT('h8)
	) name10534 (
		\wishbone_bd_ram_mem2_reg[53][19]/P0001 ,
		_w13020_,
		_w21046_
	);
	LUT2 #(
		.INIT('h8)
	) name10535 (
		\wishbone_bd_ram_mem2_reg[111][19]/P0001 ,
		_w12744_,
		_w21047_
	);
	LUT2 #(
		.INIT('h8)
	) name10536 (
		\wishbone_bd_ram_mem2_reg[128][19]/P0001 ,
		_w12793_,
		_w21048_
	);
	LUT2 #(
		.INIT('h8)
	) name10537 (
		\wishbone_bd_ram_mem2_reg[254][19]/P0001 ,
		_w12892_,
		_w21049_
	);
	LUT2 #(
		.INIT('h8)
	) name10538 (
		\wishbone_bd_ram_mem2_reg[196][19]/P0001 ,
		_w13090_,
		_w21050_
	);
	LUT2 #(
		.INIT('h8)
	) name10539 (
		\wishbone_bd_ram_mem2_reg[17][19]/P0001 ,
		_w12848_,
		_w21051_
	);
	LUT2 #(
		.INIT('h8)
	) name10540 (
		\wishbone_bd_ram_mem2_reg[43][19]/P0001 ,
		_w13200_,
		_w21052_
	);
	LUT2 #(
		.INIT('h8)
	) name10541 (
		\wishbone_bd_ram_mem2_reg[231][19]/P0001 ,
		_w12856_,
		_w21053_
	);
	LUT2 #(
		.INIT('h8)
	) name10542 (
		\wishbone_bd_ram_mem2_reg[40][19]/P0001 ,
		_w13132_,
		_w21054_
	);
	LUT2 #(
		.INIT('h8)
	) name10543 (
		\wishbone_bd_ram_mem2_reg[93][19]/P0001 ,
		_w13016_,
		_w21055_
	);
	LUT2 #(
		.INIT('h8)
	) name10544 (
		\wishbone_bd_ram_mem2_reg[48][19]/P0001 ,
		_w12970_,
		_w21056_
	);
	LUT2 #(
		.INIT('h8)
	) name10545 (
		\wishbone_bd_ram_mem2_reg[141][19]/P0001 ,
		_w13004_,
		_w21057_
	);
	LUT2 #(
		.INIT('h8)
	) name10546 (
		\wishbone_bd_ram_mem2_reg[167][19]/P0001 ,
		_w12986_,
		_w21058_
	);
	LUT2 #(
		.INIT('h8)
	) name10547 (
		\wishbone_bd_ram_mem2_reg[125][19]/P0001 ,
		_w12956_,
		_w21059_
	);
	LUT2 #(
		.INIT('h8)
	) name10548 (
		\wishbone_bd_ram_mem2_reg[173][19]/P0001 ,
		_w12854_,
		_w21060_
	);
	LUT2 #(
		.INIT('h8)
	) name10549 (
		\wishbone_bd_ram_mem2_reg[240][19]/P0001 ,
		_w12864_,
		_w21061_
	);
	LUT2 #(
		.INIT('h8)
	) name10550 (
		\wishbone_bd_ram_mem2_reg[211][19]/P0001 ,
		_w13166_,
		_w21062_
	);
	LUT2 #(
		.INIT('h8)
	) name10551 (
		\wishbone_bd_ram_mem2_reg[116][19]/P0001 ,
		_w12998_,
		_w21063_
	);
	LUT2 #(
		.INIT('h8)
	) name10552 (
		\wishbone_bd_ram_mem2_reg[46][19]/P0001 ,
		_w12884_,
		_w21064_
	);
	LUT2 #(
		.INIT('h8)
	) name10553 (
		\wishbone_bd_ram_mem2_reg[19][19]/P0001 ,
		_w13012_,
		_w21065_
	);
	LUT2 #(
		.INIT('h8)
	) name10554 (
		\wishbone_bd_ram_mem2_reg[165][19]/P0001 ,
		_w13044_,
		_w21066_
	);
	LUT2 #(
		.INIT('h8)
	) name10555 (
		\wishbone_bd_ram_mem2_reg[218][19]/P0001 ,
		_w13206_,
		_w21067_
	);
	LUT2 #(
		.INIT('h8)
	) name10556 (
		\wishbone_bd_ram_mem2_reg[115][19]/P0001 ,
		_w13112_,
		_w21068_
	);
	LUT2 #(
		.INIT('h8)
	) name10557 (
		\wishbone_bd_ram_mem2_reg[192][19]/P0001 ,
		_w12938_,
		_w21069_
	);
	LUT2 #(
		.INIT('h8)
	) name10558 (
		\wishbone_bd_ram_mem2_reg[197][19]/P0001 ,
		_w12834_,
		_w21070_
	);
	LUT2 #(
		.INIT('h8)
	) name10559 (
		\wishbone_bd_ram_mem2_reg[12][19]/P0001 ,
		_w13118_,
		_w21071_
	);
	LUT2 #(
		.INIT('h8)
	) name10560 (
		\wishbone_bd_ram_mem2_reg[112][19]/P0001 ,
		_w12733_,
		_w21072_
	);
	LUT2 #(
		.INIT('h8)
	) name10561 (
		\wishbone_bd_ram_mem2_reg[253][19]/P0001 ,
		_w13100_,
		_w21073_
	);
	LUT2 #(
		.INIT('h8)
	) name10562 (
		\wishbone_bd_ram_mem2_reg[226][19]/P0001 ,
		_w13138_,
		_w21074_
	);
	LUT2 #(
		.INIT('h8)
	) name10563 (
		\wishbone_bd_ram_mem2_reg[195][19]/P0001 ,
		_w13144_,
		_w21075_
	);
	LUT2 #(
		.INIT('h8)
	) name10564 (
		\wishbone_bd_ram_mem2_reg[146][19]/P0001 ,
		_w13060_,
		_w21076_
	);
	LUT2 #(
		.INIT('h8)
	) name10565 (
		\wishbone_bd_ram_mem2_reg[179][19]/P0001 ,
		_w13050_,
		_w21077_
	);
	LUT2 #(
		.INIT('h8)
	) name10566 (
		\wishbone_bd_ram_mem2_reg[162][19]/P0001 ,
		_w13098_,
		_w21078_
	);
	LUT2 #(
		.INIT('h8)
	) name10567 (
		\wishbone_bd_ram_mem2_reg[105][19]/P0001 ,
		_w12751_,
		_w21079_
	);
	LUT2 #(
		.INIT('h8)
	) name10568 (
		\wishbone_bd_ram_mem2_reg[189][19]/P0001 ,
		_w13042_,
		_w21080_
	);
	LUT2 #(
		.INIT('h8)
	) name10569 (
		\wishbone_bd_ram_mem2_reg[171][19]/P0001 ,
		_w12910_,
		_w21081_
	);
	LUT2 #(
		.INIT('h8)
	) name10570 (
		\wishbone_bd_ram_mem2_reg[188][19]/P0001 ,
		_w12948_,
		_w21082_
	);
	LUT2 #(
		.INIT('h8)
	) name10571 (
		\wishbone_bd_ram_mem2_reg[45][19]/P0001 ,
		_w12908_,
		_w21083_
	);
	LUT2 #(
		.INIT('h8)
	) name10572 (
		\wishbone_bd_ram_mem2_reg[224][19]/P0001 ,
		_w12902_,
		_w21084_
	);
	LUT2 #(
		.INIT('h8)
	) name10573 (
		\wishbone_bd_ram_mem2_reg[174][19]/P0001 ,
		_w12972_,
		_w21085_
	);
	LUT2 #(
		.INIT('h8)
	) name10574 (
		\wishbone_bd_ram_mem2_reg[202][19]/P0001 ,
		_w12870_,
		_w21086_
	);
	LUT2 #(
		.INIT('h8)
	) name10575 (
		\wishbone_bd_ram_mem2_reg[22][19]/P0001 ,
		_w13110_,
		_w21087_
	);
	LUT2 #(
		.INIT('h8)
	) name10576 (
		\wishbone_bd_ram_mem2_reg[120][19]/P0001 ,
		_w12707_,
		_w21088_
	);
	LUT2 #(
		.INIT('h8)
	) name10577 (
		\wishbone_bd_ram_mem2_reg[185][19]/P0001 ,
		_w12940_,
		_w21089_
	);
	LUT2 #(
		.INIT('h8)
	) name10578 (
		\wishbone_bd_ram_mem2_reg[101][19]/P0001 ,
		_w13192_,
		_w21090_
	);
	LUT2 #(
		.INIT('h8)
	) name10579 (
		\wishbone_bd_ram_mem2_reg[241][19]/P0001 ,
		_w13006_,
		_w21091_
	);
	LUT2 #(
		.INIT('h8)
	) name10580 (
		\wishbone_bd_ram_mem2_reg[149][19]/P0001 ,
		_w12741_,
		_w21092_
	);
	LUT2 #(
		.INIT('h8)
	) name10581 (
		\wishbone_bd_ram_mem2_reg[200][19]/P0001 ,
		_w12988_,
		_w21093_
	);
	LUT2 #(
		.INIT('h8)
	) name10582 (
		\wishbone_bd_ram_mem2_reg[50][19]/P0001 ,
		_w13150_,
		_w21094_
	);
	LUT2 #(
		.INIT('h8)
	) name10583 (
		\wishbone_bd_ram_mem2_reg[152][19]/P0001 ,
		_w12966_,
		_w21095_
	);
	LUT2 #(
		.INIT('h8)
	) name10584 (
		\wishbone_bd_ram_mem2_reg[84][19]/P0001 ,
		_w12934_,
		_w21096_
	);
	LUT2 #(
		.INIT('h8)
	) name10585 (
		\wishbone_bd_ram_mem2_reg[24][19]/P0001 ,
		_w13084_,
		_w21097_
	);
	LUT2 #(
		.INIT('h8)
	) name10586 (
		\wishbone_bd_ram_mem2_reg[97][19]/P0001 ,
		_w13096_,
		_w21098_
	);
	LUT2 #(
		.INIT('h8)
	) name10587 (
		\wishbone_bd_ram_mem2_reg[1][19]/P0001 ,
		_w13014_,
		_w21099_
	);
	LUT2 #(
		.INIT('h8)
	) name10588 (
		\wishbone_bd_ram_mem2_reg[4][19]/P0001 ,
		_w12666_,
		_w21100_
	);
	LUT2 #(
		.INIT('h8)
	) name10589 (
		\wishbone_bd_ram_mem2_reg[2][19]/P0001 ,
		_w13088_,
		_w21101_
	);
	LUT2 #(
		.INIT('h8)
	) name10590 (
		\wishbone_bd_ram_mem2_reg[246][19]/P0001 ,
		_w13076_,
		_w21102_
	);
	LUT2 #(
		.INIT('h8)
	) name10591 (
		\wishbone_bd_ram_mem2_reg[133][19]/P0001 ,
		_w12761_,
		_w21103_
	);
	LUT2 #(
		.INIT('h8)
	) name10592 (
		\wishbone_bd_ram_mem2_reg[216][19]/P0001 ,
		_w13028_,
		_w21104_
	);
	LUT2 #(
		.INIT('h8)
	) name10593 (
		\wishbone_bd_ram_mem2_reg[177][19]/P0001 ,
		_w12996_,
		_w21105_
	);
	LUT2 #(
		.INIT('h8)
	) name10594 (
		\wishbone_bd_ram_mem2_reg[175][19]/P0001 ,
		_w13126_,
		_w21106_
	);
	LUT2 #(
		.INIT('h8)
	) name10595 (
		\wishbone_bd_ram_mem2_reg[243][19]/P0001 ,
		_w12804_,
		_w21107_
	);
	LUT2 #(
		.INIT('h8)
	) name10596 (
		\wishbone_bd_ram_mem2_reg[123][19]/P0001 ,
		_w13114_,
		_w21108_
	);
	LUT2 #(
		.INIT('h8)
	) name10597 (
		\wishbone_bd_ram_mem2_reg[88][19]/P0001 ,
		_w12860_,
		_w21109_
	);
	LUT2 #(
		.INIT('h8)
	) name10598 (
		\wishbone_bd_ram_mem2_reg[251][19]/P0001 ,
		_w13054_,
		_w21110_
	);
	LUT2 #(
		.INIT('h8)
	) name10599 (
		\wishbone_bd_ram_mem2_reg[81][19]/P0001 ,
		_w12950_,
		_w21111_
	);
	LUT2 #(
		.INIT('h8)
	) name10600 (
		\wishbone_bd_ram_mem2_reg[51][19]/P0001 ,
		_w13024_,
		_w21112_
	);
	LUT2 #(
		.INIT('h8)
	) name10601 (
		\wishbone_bd_ram_mem2_reg[247][19]/P0001 ,
		_w12818_,
		_w21113_
	);
	LUT2 #(
		.INIT('h8)
	) name10602 (
		\wishbone_bd_ram_mem2_reg[186][19]/P0001 ,
		_w12783_,
		_w21114_
	);
	LUT2 #(
		.INIT('h8)
	) name10603 (
		\wishbone_bd_ram_mem2_reg[233][19]/P0001 ,
		_w12836_,
		_w21115_
	);
	LUT2 #(
		.INIT('h8)
	) name10604 (
		\wishbone_bd_ram_mem2_reg[83][19]/P0001 ,
		_w12916_,
		_w21116_
	);
	LUT2 #(
		.INIT('h8)
	) name10605 (
		\wishbone_bd_ram_mem2_reg[214][19]/P0001 ,
		_w12984_,
		_w21117_
	);
	LUT2 #(
		.INIT('h8)
	) name10606 (
		\wishbone_bd_ram_mem2_reg[220][19]/P0001 ,
		_w13066_,
		_w21118_
	);
	LUT2 #(
		.INIT('h8)
	) name10607 (
		\wishbone_bd_ram_mem2_reg[58][19]/P0001 ,
		_w13070_,
		_w21119_
	);
	LUT2 #(
		.INIT('h8)
	) name10608 (
		\wishbone_bd_ram_mem2_reg[145][19]/P0001 ,
		_w13106_,
		_w21120_
	);
	LUT2 #(
		.INIT('h8)
	) name10609 (
		\wishbone_bd_ram_mem2_reg[35][19]/P0001 ,
		_w12703_,
		_w21121_
	);
	LUT2 #(
		.INIT('h8)
	) name10610 (
		\wishbone_bd_ram_mem2_reg[94][19]/P0001 ,
		_w13186_,
		_w21122_
	);
	LUT2 #(
		.INIT('h8)
	) name10611 (
		\wishbone_bd_ram_mem2_reg[239][19]/P0001 ,
		_w12862_,
		_w21123_
	);
	LUT2 #(
		.INIT('h8)
	) name10612 (
		\wishbone_bd_ram_mem2_reg[204][19]/P0001 ,
		_w13162_,
		_w21124_
	);
	LUT2 #(
		.INIT('h8)
	) name10613 (
		\wishbone_bd_ram_mem2_reg[213][19]/P0001 ,
		_w13002_,
		_w21125_
	);
	LUT2 #(
		.INIT('h8)
	) name10614 (
		\wishbone_bd_ram_mem2_reg[90][19]/P0001 ,
		_w12978_,
		_w21126_
	);
	LUT2 #(
		.INIT('h8)
	) name10615 (
		\wishbone_bd_ram_mem2_reg[68][19]/P0001 ,
		_w12946_,
		_w21127_
	);
	LUT2 #(
		.INIT('h1)
	) name10616 (
		_w20872_,
		_w20873_,
		_w21128_
	);
	LUT2 #(
		.INIT('h1)
	) name10617 (
		_w20874_,
		_w20875_,
		_w21129_
	);
	LUT2 #(
		.INIT('h1)
	) name10618 (
		_w20876_,
		_w20877_,
		_w21130_
	);
	LUT2 #(
		.INIT('h1)
	) name10619 (
		_w20878_,
		_w20879_,
		_w21131_
	);
	LUT2 #(
		.INIT('h1)
	) name10620 (
		_w20880_,
		_w20881_,
		_w21132_
	);
	LUT2 #(
		.INIT('h1)
	) name10621 (
		_w20882_,
		_w20883_,
		_w21133_
	);
	LUT2 #(
		.INIT('h1)
	) name10622 (
		_w20884_,
		_w20885_,
		_w21134_
	);
	LUT2 #(
		.INIT('h1)
	) name10623 (
		_w20886_,
		_w20887_,
		_w21135_
	);
	LUT2 #(
		.INIT('h1)
	) name10624 (
		_w20888_,
		_w20889_,
		_w21136_
	);
	LUT2 #(
		.INIT('h1)
	) name10625 (
		_w20890_,
		_w20891_,
		_w21137_
	);
	LUT2 #(
		.INIT('h1)
	) name10626 (
		_w20892_,
		_w20893_,
		_w21138_
	);
	LUT2 #(
		.INIT('h1)
	) name10627 (
		_w20894_,
		_w20895_,
		_w21139_
	);
	LUT2 #(
		.INIT('h1)
	) name10628 (
		_w20896_,
		_w20897_,
		_w21140_
	);
	LUT2 #(
		.INIT('h1)
	) name10629 (
		_w20898_,
		_w20899_,
		_w21141_
	);
	LUT2 #(
		.INIT('h1)
	) name10630 (
		_w20900_,
		_w20901_,
		_w21142_
	);
	LUT2 #(
		.INIT('h1)
	) name10631 (
		_w20902_,
		_w20903_,
		_w21143_
	);
	LUT2 #(
		.INIT('h1)
	) name10632 (
		_w20904_,
		_w20905_,
		_w21144_
	);
	LUT2 #(
		.INIT('h1)
	) name10633 (
		_w20906_,
		_w20907_,
		_w21145_
	);
	LUT2 #(
		.INIT('h1)
	) name10634 (
		_w20908_,
		_w20909_,
		_w21146_
	);
	LUT2 #(
		.INIT('h1)
	) name10635 (
		_w20910_,
		_w20911_,
		_w21147_
	);
	LUT2 #(
		.INIT('h1)
	) name10636 (
		_w20912_,
		_w20913_,
		_w21148_
	);
	LUT2 #(
		.INIT('h1)
	) name10637 (
		_w20914_,
		_w20915_,
		_w21149_
	);
	LUT2 #(
		.INIT('h1)
	) name10638 (
		_w20916_,
		_w20917_,
		_w21150_
	);
	LUT2 #(
		.INIT('h1)
	) name10639 (
		_w20918_,
		_w20919_,
		_w21151_
	);
	LUT2 #(
		.INIT('h1)
	) name10640 (
		_w20920_,
		_w20921_,
		_w21152_
	);
	LUT2 #(
		.INIT('h1)
	) name10641 (
		_w20922_,
		_w20923_,
		_w21153_
	);
	LUT2 #(
		.INIT('h1)
	) name10642 (
		_w20924_,
		_w20925_,
		_w21154_
	);
	LUT2 #(
		.INIT('h1)
	) name10643 (
		_w20926_,
		_w20927_,
		_w21155_
	);
	LUT2 #(
		.INIT('h1)
	) name10644 (
		_w20928_,
		_w20929_,
		_w21156_
	);
	LUT2 #(
		.INIT('h1)
	) name10645 (
		_w20930_,
		_w20931_,
		_w21157_
	);
	LUT2 #(
		.INIT('h1)
	) name10646 (
		_w20932_,
		_w20933_,
		_w21158_
	);
	LUT2 #(
		.INIT('h1)
	) name10647 (
		_w20934_,
		_w20935_,
		_w21159_
	);
	LUT2 #(
		.INIT('h1)
	) name10648 (
		_w20936_,
		_w20937_,
		_w21160_
	);
	LUT2 #(
		.INIT('h1)
	) name10649 (
		_w20938_,
		_w20939_,
		_w21161_
	);
	LUT2 #(
		.INIT('h1)
	) name10650 (
		_w20940_,
		_w20941_,
		_w21162_
	);
	LUT2 #(
		.INIT('h1)
	) name10651 (
		_w20942_,
		_w20943_,
		_w21163_
	);
	LUT2 #(
		.INIT('h1)
	) name10652 (
		_w20944_,
		_w20945_,
		_w21164_
	);
	LUT2 #(
		.INIT('h1)
	) name10653 (
		_w20946_,
		_w20947_,
		_w21165_
	);
	LUT2 #(
		.INIT('h1)
	) name10654 (
		_w20948_,
		_w20949_,
		_w21166_
	);
	LUT2 #(
		.INIT('h1)
	) name10655 (
		_w20950_,
		_w20951_,
		_w21167_
	);
	LUT2 #(
		.INIT('h1)
	) name10656 (
		_w20952_,
		_w20953_,
		_w21168_
	);
	LUT2 #(
		.INIT('h1)
	) name10657 (
		_w20954_,
		_w20955_,
		_w21169_
	);
	LUT2 #(
		.INIT('h1)
	) name10658 (
		_w20956_,
		_w20957_,
		_w21170_
	);
	LUT2 #(
		.INIT('h1)
	) name10659 (
		_w20958_,
		_w20959_,
		_w21171_
	);
	LUT2 #(
		.INIT('h1)
	) name10660 (
		_w20960_,
		_w20961_,
		_w21172_
	);
	LUT2 #(
		.INIT('h1)
	) name10661 (
		_w20962_,
		_w20963_,
		_w21173_
	);
	LUT2 #(
		.INIT('h1)
	) name10662 (
		_w20964_,
		_w20965_,
		_w21174_
	);
	LUT2 #(
		.INIT('h1)
	) name10663 (
		_w20966_,
		_w20967_,
		_w21175_
	);
	LUT2 #(
		.INIT('h1)
	) name10664 (
		_w20968_,
		_w20969_,
		_w21176_
	);
	LUT2 #(
		.INIT('h1)
	) name10665 (
		_w20970_,
		_w20971_,
		_w21177_
	);
	LUT2 #(
		.INIT('h1)
	) name10666 (
		_w20972_,
		_w20973_,
		_w21178_
	);
	LUT2 #(
		.INIT('h1)
	) name10667 (
		_w20974_,
		_w20975_,
		_w21179_
	);
	LUT2 #(
		.INIT('h1)
	) name10668 (
		_w20976_,
		_w20977_,
		_w21180_
	);
	LUT2 #(
		.INIT('h1)
	) name10669 (
		_w20978_,
		_w20979_,
		_w21181_
	);
	LUT2 #(
		.INIT('h1)
	) name10670 (
		_w20980_,
		_w20981_,
		_w21182_
	);
	LUT2 #(
		.INIT('h1)
	) name10671 (
		_w20982_,
		_w20983_,
		_w21183_
	);
	LUT2 #(
		.INIT('h1)
	) name10672 (
		_w20984_,
		_w20985_,
		_w21184_
	);
	LUT2 #(
		.INIT('h1)
	) name10673 (
		_w20986_,
		_w20987_,
		_w21185_
	);
	LUT2 #(
		.INIT('h1)
	) name10674 (
		_w20988_,
		_w20989_,
		_w21186_
	);
	LUT2 #(
		.INIT('h1)
	) name10675 (
		_w20990_,
		_w20991_,
		_w21187_
	);
	LUT2 #(
		.INIT('h1)
	) name10676 (
		_w20992_,
		_w20993_,
		_w21188_
	);
	LUT2 #(
		.INIT('h1)
	) name10677 (
		_w20994_,
		_w20995_,
		_w21189_
	);
	LUT2 #(
		.INIT('h1)
	) name10678 (
		_w20996_,
		_w20997_,
		_w21190_
	);
	LUT2 #(
		.INIT('h1)
	) name10679 (
		_w20998_,
		_w20999_,
		_w21191_
	);
	LUT2 #(
		.INIT('h1)
	) name10680 (
		_w21000_,
		_w21001_,
		_w21192_
	);
	LUT2 #(
		.INIT('h1)
	) name10681 (
		_w21002_,
		_w21003_,
		_w21193_
	);
	LUT2 #(
		.INIT('h1)
	) name10682 (
		_w21004_,
		_w21005_,
		_w21194_
	);
	LUT2 #(
		.INIT('h1)
	) name10683 (
		_w21006_,
		_w21007_,
		_w21195_
	);
	LUT2 #(
		.INIT('h1)
	) name10684 (
		_w21008_,
		_w21009_,
		_w21196_
	);
	LUT2 #(
		.INIT('h1)
	) name10685 (
		_w21010_,
		_w21011_,
		_w21197_
	);
	LUT2 #(
		.INIT('h1)
	) name10686 (
		_w21012_,
		_w21013_,
		_w21198_
	);
	LUT2 #(
		.INIT('h1)
	) name10687 (
		_w21014_,
		_w21015_,
		_w21199_
	);
	LUT2 #(
		.INIT('h1)
	) name10688 (
		_w21016_,
		_w21017_,
		_w21200_
	);
	LUT2 #(
		.INIT('h1)
	) name10689 (
		_w21018_,
		_w21019_,
		_w21201_
	);
	LUT2 #(
		.INIT('h1)
	) name10690 (
		_w21020_,
		_w21021_,
		_w21202_
	);
	LUT2 #(
		.INIT('h1)
	) name10691 (
		_w21022_,
		_w21023_,
		_w21203_
	);
	LUT2 #(
		.INIT('h1)
	) name10692 (
		_w21024_,
		_w21025_,
		_w21204_
	);
	LUT2 #(
		.INIT('h1)
	) name10693 (
		_w21026_,
		_w21027_,
		_w21205_
	);
	LUT2 #(
		.INIT('h1)
	) name10694 (
		_w21028_,
		_w21029_,
		_w21206_
	);
	LUT2 #(
		.INIT('h1)
	) name10695 (
		_w21030_,
		_w21031_,
		_w21207_
	);
	LUT2 #(
		.INIT('h1)
	) name10696 (
		_w21032_,
		_w21033_,
		_w21208_
	);
	LUT2 #(
		.INIT('h1)
	) name10697 (
		_w21034_,
		_w21035_,
		_w21209_
	);
	LUT2 #(
		.INIT('h1)
	) name10698 (
		_w21036_,
		_w21037_,
		_w21210_
	);
	LUT2 #(
		.INIT('h1)
	) name10699 (
		_w21038_,
		_w21039_,
		_w21211_
	);
	LUT2 #(
		.INIT('h1)
	) name10700 (
		_w21040_,
		_w21041_,
		_w21212_
	);
	LUT2 #(
		.INIT('h1)
	) name10701 (
		_w21042_,
		_w21043_,
		_w21213_
	);
	LUT2 #(
		.INIT('h1)
	) name10702 (
		_w21044_,
		_w21045_,
		_w21214_
	);
	LUT2 #(
		.INIT('h1)
	) name10703 (
		_w21046_,
		_w21047_,
		_w21215_
	);
	LUT2 #(
		.INIT('h1)
	) name10704 (
		_w21048_,
		_w21049_,
		_w21216_
	);
	LUT2 #(
		.INIT('h1)
	) name10705 (
		_w21050_,
		_w21051_,
		_w21217_
	);
	LUT2 #(
		.INIT('h1)
	) name10706 (
		_w21052_,
		_w21053_,
		_w21218_
	);
	LUT2 #(
		.INIT('h1)
	) name10707 (
		_w21054_,
		_w21055_,
		_w21219_
	);
	LUT2 #(
		.INIT('h1)
	) name10708 (
		_w21056_,
		_w21057_,
		_w21220_
	);
	LUT2 #(
		.INIT('h1)
	) name10709 (
		_w21058_,
		_w21059_,
		_w21221_
	);
	LUT2 #(
		.INIT('h1)
	) name10710 (
		_w21060_,
		_w21061_,
		_w21222_
	);
	LUT2 #(
		.INIT('h1)
	) name10711 (
		_w21062_,
		_w21063_,
		_w21223_
	);
	LUT2 #(
		.INIT('h1)
	) name10712 (
		_w21064_,
		_w21065_,
		_w21224_
	);
	LUT2 #(
		.INIT('h1)
	) name10713 (
		_w21066_,
		_w21067_,
		_w21225_
	);
	LUT2 #(
		.INIT('h1)
	) name10714 (
		_w21068_,
		_w21069_,
		_w21226_
	);
	LUT2 #(
		.INIT('h1)
	) name10715 (
		_w21070_,
		_w21071_,
		_w21227_
	);
	LUT2 #(
		.INIT('h1)
	) name10716 (
		_w21072_,
		_w21073_,
		_w21228_
	);
	LUT2 #(
		.INIT('h1)
	) name10717 (
		_w21074_,
		_w21075_,
		_w21229_
	);
	LUT2 #(
		.INIT('h1)
	) name10718 (
		_w21076_,
		_w21077_,
		_w21230_
	);
	LUT2 #(
		.INIT('h1)
	) name10719 (
		_w21078_,
		_w21079_,
		_w21231_
	);
	LUT2 #(
		.INIT('h1)
	) name10720 (
		_w21080_,
		_w21081_,
		_w21232_
	);
	LUT2 #(
		.INIT('h1)
	) name10721 (
		_w21082_,
		_w21083_,
		_w21233_
	);
	LUT2 #(
		.INIT('h1)
	) name10722 (
		_w21084_,
		_w21085_,
		_w21234_
	);
	LUT2 #(
		.INIT('h1)
	) name10723 (
		_w21086_,
		_w21087_,
		_w21235_
	);
	LUT2 #(
		.INIT('h1)
	) name10724 (
		_w21088_,
		_w21089_,
		_w21236_
	);
	LUT2 #(
		.INIT('h1)
	) name10725 (
		_w21090_,
		_w21091_,
		_w21237_
	);
	LUT2 #(
		.INIT('h1)
	) name10726 (
		_w21092_,
		_w21093_,
		_w21238_
	);
	LUT2 #(
		.INIT('h1)
	) name10727 (
		_w21094_,
		_w21095_,
		_w21239_
	);
	LUT2 #(
		.INIT('h1)
	) name10728 (
		_w21096_,
		_w21097_,
		_w21240_
	);
	LUT2 #(
		.INIT('h1)
	) name10729 (
		_w21098_,
		_w21099_,
		_w21241_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		_w21100_,
		_w21101_,
		_w21242_
	);
	LUT2 #(
		.INIT('h1)
	) name10731 (
		_w21102_,
		_w21103_,
		_w21243_
	);
	LUT2 #(
		.INIT('h1)
	) name10732 (
		_w21104_,
		_w21105_,
		_w21244_
	);
	LUT2 #(
		.INIT('h1)
	) name10733 (
		_w21106_,
		_w21107_,
		_w21245_
	);
	LUT2 #(
		.INIT('h1)
	) name10734 (
		_w21108_,
		_w21109_,
		_w21246_
	);
	LUT2 #(
		.INIT('h1)
	) name10735 (
		_w21110_,
		_w21111_,
		_w21247_
	);
	LUT2 #(
		.INIT('h1)
	) name10736 (
		_w21112_,
		_w21113_,
		_w21248_
	);
	LUT2 #(
		.INIT('h1)
	) name10737 (
		_w21114_,
		_w21115_,
		_w21249_
	);
	LUT2 #(
		.INIT('h1)
	) name10738 (
		_w21116_,
		_w21117_,
		_w21250_
	);
	LUT2 #(
		.INIT('h1)
	) name10739 (
		_w21118_,
		_w21119_,
		_w21251_
	);
	LUT2 #(
		.INIT('h1)
	) name10740 (
		_w21120_,
		_w21121_,
		_w21252_
	);
	LUT2 #(
		.INIT('h1)
	) name10741 (
		_w21122_,
		_w21123_,
		_w21253_
	);
	LUT2 #(
		.INIT('h1)
	) name10742 (
		_w21124_,
		_w21125_,
		_w21254_
	);
	LUT2 #(
		.INIT('h1)
	) name10743 (
		_w21126_,
		_w21127_,
		_w21255_
	);
	LUT2 #(
		.INIT('h8)
	) name10744 (
		_w21254_,
		_w21255_,
		_w21256_
	);
	LUT2 #(
		.INIT('h8)
	) name10745 (
		_w21252_,
		_w21253_,
		_w21257_
	);
	LUT2 #(
		.INIT('h8)
	) name10746 (
		_w21250_,
		_w21251_,
		_w21258_
	);
	LUT2 #(
		.INIT('h8)
	) name10747 (
		_w21248_,
		_w21249_,
		_w21259_
	);
	LUT2 #(
		.INIT('h8)
	) name10748 (
		_w21246_,
		_w21247_,
		_w21260_
	);
	LUT2 #(
		.INIT('h8)
	) name10749 (
		_w21244_,
		_w21245_,
		_w21261_
	);
	LUT2 #(
		.INIT('h8)
	) name10750 (
		_w21242_,
		_w21243_,
		_w21262_
	);
	LUT2 #(
		.INIT('h8)
	) name10751 (
		_w21240_,
		_w21241_,
		_w21263_
	);
	LUT2 #(
		.INIT('h8)
	) name10752 (
		_w21238_,
		_w21239_,
		_w21264_
	);
	LUT2 #(
		.INIT('h8)
	) name10753 (
		_w21236_,
		_w21237_,
		_w21265_
	);
	LUT2 #(
		.INIT('h8)
	) name10754 (
		_w21234_,
		_w21235_,
		_w21266_
	);
	LUT2 #(
		.INIT('h8)
	) name10755 (
		_w21232_,
		_w21233_,
		_w21267_
	);
	LUT2 #(
		.INIT('h8)
	) name10756 (
		_w21230_,
		_w21231_,
		_w21268_
	);
	LUT2 #(
		.INIT('h8)
	) name10757 (
		_w21228_,
		_w21229_,
		_w21269_
	);
	LUT2 #(
		.INIT('h8)
	) name10758 (
		_w21226_,
		_w21227_,
		_w21270_
	);
	LUT2 #(
		.INIT('h8)
	) name10759 (
		_w21224_,
		_w21225_,
		_w21271_
	);
	LUT2 #(
		.INIT('h8)
	) name10760 (
		_w21222_,
		_w21223_,
		_w21272_
	);
	LUT2 #(
		.INIT('h8)
	) name10761 (
		_w21220_,
		_w21221_,
		_w21273_
	);
	LUT2 #(
		.INIT('h8)
	) name10762 (
		_w21218_,
		_w21219_,
		_w21274_
	);
	LUT2 #(
		.INIT('h8)
	) name10763 (
		_w21216_,
		_w21217_,
		_w21275_
	);
	LUT2 #(
		.INIT('h8)
	) name10764 (
		_w21214_,
		_w21215_,
		_w21276_
	);
	LUT2 #(
		.INIT('h8)
	) name10765 (
		_w21212_,
		_w21213_,
		_w21277_
	);
	LUT2 #(
		.INIT('h8)
	) name10766 (
		_w21210_,
		_w21211_,
		_w21278_
	);
	LUT2 #(
		.INIT('h8)
	) name10767 (
		_w21208_,
		_w21209_,
		_w21279_
	);
	LUT2 #(
		.INIT('h8)
	) name10768 (
		_w21206_,
		_w21207_,
		_w21280_
	);
	LUT2 #(
		.INIT('h8)
	) name10769 (
		_w21204_,
		_w21205_,
		_w21281_
	);
	LUT2 #(
		.INIT('h8)
	) name10770 (
		_w21202_,
		_w21203_,
		_w21282_
	);
	LUT2 #(
		.INIT('h8)
	) name10771 (
		_w21200_,
		_w21201_,
		_w21283_
	);
	LUT2 #(
		.INIT('h8)
	) name10772 (
		_w21198_,
		_w21199_,
		_w21284_
	);
	LUT2 #(
		.INIT('h8)
	) name10773 (
		_w21196_,
		_w21197_,
		_w21285_
	);
	LUT2 #(
		.INIT('h8)
	) name10774 (
		_w21194_,
		_w21195_,
		_w21286_
	);
	LUT2 #(
		.INIT('h8)
	) name10775 (
		_w21192_,
		_w21193_,
		_w21287_
	);
	LUT2 #(
		.INIT('h8)
	) name10776 (
		_w21190_,
		_w21191_,
		_w21288_
	);
	LUT2 #(
		.INIT('h8)
	) name10777 (
		_w21188_,
		_w21189_,
		_w21289_
	);
	LUT2 #(
		.INIT('h8)
	) name10778 (
		_w21186_,
		_w21187_,
		_w21290_
	);
	LUT2 #(
		.INIT('h8)
	) name10779 (
		_w21184_,
		_w21185_,
		_w21291_
	);
	LUT2 #(
		.INIT('h8)
	) name10780 (
		_w21182_,
		_w21183_,
		_w21292_
	);
	LUT2 #(
		.INIT('h8)
	) name10781 (
		_w21180_,
		_w21181_,
		_w21293_
	);
	LUT2 #(
		.INIT('h8)
	) name10782 (
		_w21178_,
		_w21179_,
		_w21294_
	);
	LUT2 #(
		.INIT('h8)
	) name10783 (
		_w21176_,
		_w21177_,
		_w21295_
	);
	LUT2 #(
		.INIT('h8)
	) name10784 (
		_w21174_,
		_w21175_,
		_w21296_
	);
	LUT2 #(
		.INIT('h8)
	) name10785 (
		_w21172_,
		_w21173_,
		_w21297_
	);
	LUT2 #(
		.INIT('h8)
	) name10786 (
		_w21170_,
		_w21171_,
		_w21298_
	);
	LUT2 #(
		.INIT('h8)
	) name10787 (
		_w21168_,
		_w21169_,
		_w21299_
	);
	LUT2 #(
		.INIT('h8)
	) name10788 (
		_w21166_,
		_w21167_,
		_w21300_
	);
	LUT2 #(
		.INIT('h8)
	) name10789 (
		_w21164_,
		_w21165_,
		_w21301_
	);
	LUT2 #(
		.INIT('h8)
	) name10790 (
		_w21162_,
		_w21163_,
		_w21302_
	);
	LUT2 #(
		.INIT('h8)
	) name10791 (
		_w21160_,
		_w21161_,
		_w21303_
	);
	LUT2 #(
		.INIT('h8)
	) name10792 (
		_w21158_,
		_w21159_,
		_w21304_
	);
	LUT2 #(
		.INIT('h8)
	) name10793 (
		_w21156_,
		_w21157_,
		_w21305_
	);
	LUT2 #(
		.INIT('h8)
	) name10794 (
		_w21154_,
		_w21155_,
		_w21306_
	);
	LUT2 #(
		.INIT('h8)
	) name10795 (
		_w21152_,
		_w21153_,
		_w21307_
	);
	LUT2 #(
		.INIT('h8)
	) name10796 (
		_w21150_,
		_w21151_,
		_w21308_
	);
	LUT2 #(
		.INIT('h8)
	) name10797 (
		_w21148_,
		_w21149_,
		_w21309_
	);
	LUT2 #(
		.INIT('h8)
	) name10798 (
		_w21146_,
		_w21147_,
		_w21310_
	);
	LUT2 #(
		.INIT('h8)
	) name10799 (
		_w21144_,
		_w21145_,
		_w21311_
	);
	LUT2 #(
		.INIT('h8)
	) name10800 (
		_w21142_,
		_w21143_,
		_w21312_
	);
	LUT2 #(
		.INIT('h8)
	) name10801 (
		_w21140_,
		_w21141_,
		_w21313_
	);
	LUT2 #(
		.INIT('h8)
	) name10802 (
		_w21138_,
		_w21139_,
		_w21314_
	);
	LUT2 #(
		.INIT('h8)
	) name10803 (
		_w21136_,
		_w21137_,
		_w21315_
	);
	LUT2 #(
		.INIT('h8)
	) name10804 (
		_w21134_,
		_w21135_,
		_w21316_
	);
	LUT2 #(
		.INIT('h8)
	) name10805 (
		_w21132_,
		_w21133_,
		_w21317_
	);
	LUT2 #(
		.INIT('h8)
	) name10806 (
		_w21130_,
		_w21131_,
		_w21318_
	);
	LUT2 #(
		.INIT('h8)
	) name10807 (
		_w21128_,
		_w21129_,
		_w21319_
	);
	LUT2 #(
		.INIT('h8)
	) name10808 (
		_w21318_,
		_w21319_,
		_w21320_
	);
	LUT2 #(
		.INIT('h8)
	) name10809 (
		_w21316_,
		_w21317_,
		_w21321_
	);
	LUT2 #(
		.INIT('h8)
	) name10810 (
		_w21314_,
		_w21315_,
		_w21322_
	);
	LUT2 #(
		.INIT('h8)
	) name10811 (
		_w21312_,
		_w21313_,
		_w21323_
	);
	LUT2 #(
		.INIT('h8)
	) name10812 (
		_w21310_,
		_w21311_,
		_w21324_
	);
	LUT2 #(
		.INIT('h8)
	) name10813 (
		_w21308_,
		_w21309_,
		_w21325_
	);
	LUT2 #(
		.INIT('h8)
	) name10814 (
		_w21306_,
		_w21307_,
		_w21326_
	);
	LUT2 #(
		.INIT('h8)
	) name10815 (
		_w21304_,
		_w21305_,
		_w21327_
	);
	LUT2 #(
		.INIT('h8)
	) name10816 (
		_w21302_,
		_w21303_,
		_w21328_
	);
	LUT2 #(
		.INIT('h8)
	) name10817 (
		_w21300_,
		_w21301_,
		_w21329_
	);
	LUT2 #(
		.INIT('h8)
	) name10818 (
		_w21298_,
		_w21299_,
		_w21330_
	);
	LUT2 #(
		.INIT('h8)
	) name10819 (
		_w21296_,
		_w21297_,
		_w21331_
	);
	LUT2 #(
		.INIT('h8)
	) name10820 (
		_w21294_,
		_w21295_,
		_w21332_
	);
	LUT2 #(
		.INIT('h8)
	) name10821 (
		_w21292_,
		_w21293_,
		_w21333_
	);
	LUT2 #(
		.INIT('h8)
	) name10822 (
		_w21290_,
		_w21291_,
		_w21334_
	);
	LUT2 #(
		.INIT('h8)
	) name10823 (
		_w21288_,
		_w21289_,
		_w21335_
	);
	LUT2 #(
		.INIT('h8)
	) name10824 (
		_w21286_,
		_w21287_,
		_w21336_
	);
	LUT2 #(
		.INIT('h8)
	) name10825 (
		_w21284_,
		_w21285_,
		_w21337_
	);
	LUT2 #(
		.INIT('h8)
	) name10826 (
		_w21282_,
		_w21283_,
		_w21338_
	);
	LUT2 #(
		.INIT('h8)
	) name10827 (
		_w21280_,
		_w21281_,
		_w21339_
	);
	LUT2 #(
		.INIT('h8)
	) name10828 (
		_w21278_,
		_w21279_,
		_w21340_
	);
	LUT2 #(
		.INIT('h8)
	) name10829 (
		_w21276_,
		_w21277_,
		_w21341_
	);
	LUT2 #(
		.INIT('h8)
	) name10830 (
		_w21274_,
		_w21275_,
		_w21342_
	);
	LUT2 #(
		.INIT('h8)
	) name10831 (
		_w21272_,
		_w21273_,
		_w21343_
	);
	LUT2 #(
		.INIT('h8)
	) name10832 (
		_w21270_,
		_w21271_,
		_w21344_
	);
	LUT2 #(
		.INIT('h8)
	) name10833 (
		_w21268_,
		_w21269_,
		_w21345_
	);
	LUT2 #(
		.INIT('h8)
	) name10834 (
		_w21266_,
		_w21267_,
		_w21346_
	);
	LUT2 #(
		.INIT('h8)
	) name10835 (
		_w21264_,
		_w21265_,
		_w21347_
	);
	LUT2 #(
		.INIT('h8)
	) name10836 (
		_w21262_,
		_w21263_,
		_w21348_
	);
	LUT2 #(
		.INIT('h8)
	) name10837 (
		_w21260_,
		_w21261_,
		_w21349_
	);
	LUT2 #(
		.INIT('h8)
	) name10838 (
		_w21258_,
		_w21259_,
		_w21350_
	);
	LUT2 #(
		.INIT('h8)
	) name10839 (
		_w21256_,
		_w21257_,
		_w21351_
	);
	LUT2 #(
		.INIT('h8)
	) name10840 (
		_w21350_,
		_w21351_,
		_w21352_
	);
	LUT2 #(
		.INIT('h8)
	) name10841 (
		_w21348_,
		_w21349_,
		_w21353_
	);
	LUT2 #(
		.INIT('h8)
	) name10842 (
		_w21346_,
		_w21347_,
		_w21354_
	);
	LUT2 #(
		.INIT('h8)
	) name10843 (
		_w21344_,
		_w21345_,
		_w21355_
	);
	LUT2 #(
		.INIT('h8)
	) name10844 (
		_w21342_,
		_w21343_,
		_w21356_
	);
	LUT2 #(
		.INIT('h8)
	) name10845 (
		_w21340_,
		_w21341_,
		_w21357_
	);
	LUT2 #(
		.INIT('h8)
	) name10846 (
		_w21338_,
		_w21339_,
		_w21358_
	);
	LUT2 #(
		.INIT('h8)
	) name10847 (
		_w21336_,
		_w21337_,
		_w21359_
	);
	LUT2 #(
		.INIT('h8)
	) name10848 (
		_w21334_,
		_w21335_,
		_w21360_
	);
	LUT2 #(
		.INIT('h8)
	) name10849 (
		_w21332_,
		_w21333_,
		_w21361_
	);
	LUT2 #(
		.INIT('h8)
	) name10850 (
		_w21330_,
		_w21331_,
		_w21362_
	);
	LUT2 #(
		.INIT('h8)
	) name10851 (
		_w21328_,
		_w21329_,
		_w21363_
	);
	LUT2 #(
		.INIT('h8)
	) name10852 (
		_w21326_,
		_w21327_,
		_w21364_
	);
	LUT2 #(
		.INIT('h8)
	) name10853 (
		_w21324_,
		_w21325_,
		_w21365_
	);
	LUT2 #(
		.INIT('h8)
	) name10854 (
		_w21322_,
		_w21323_,
		_w21366_
	);
	LUT2 #(
		.INIT('h8)
	) name10855 (
		_w21320_,
		_w21321_,
		_w21367_
	);
	LUT2 #(
		.INIT('h8)
	) name10856 (
		_w21366_,
		_w21367_,
		_w21368_
	);
	LUT2 #(
		.INIT('h8)
	) name10857 (
		_w21364_,
		_w21365_,
		_w21369_
	);
	LUT2 #(
		.INIT('h8)
	) name10858 (
		_w21362_,
		_w21363_,
		_w21370_
	);
	LUT2 #(
		.INIT('h8)
	) name10859 (
		_w21360_,
		_w21361_,
		_w21371_
	);
	LUT2 #(
		.INIT('h8)
	) name10860 (
		_w21358_,
		_w21359_,
		_w21372_
	);
	LUT2 #(
		.INIT('h8)
	) name10861 (
		_w21356_,
		_w21357_,
		_w21373_
	);
	LUT2 #(
		.INIT('h8)
	) name10862 (
		_w21354_,
		_w21355_,
		_w21374_
	);
	LUT2 #(
		.INIT('h8)
	) name10863 (
		_w21352_,
		_w21353_,
		_w21375_
	);
	LUT2 #(
		.INIT('h8)
	) name10864 (
		_w21374_,
		_w21375_,
		_w21376_
	);
	LUT2 #(
		.INIT('h8)
	) name10865 (
		_w21372_,
		_w21373_,
		_w21377_
	);
	LUT2 #(
		.INIT('h8)
	) name10866 (
		_w21370_,
		_w21371_,
		_w21378_
	);
	LUT2 #(
		.INIT('h8)
	) name10867 (
		_w21368_,
		_w21369_,
		_w21379_
	);
	LUT2 #(
		.INIT('h8)
	) name10868 (
		_w21378_,
		_w21379_,
		_w21380_
	);
	LUT2 #(
		.INIT('h8)
	) name10869 (
		_w21376_,
		_w21377_,
		_w21381_
	);
	LUT2 #(
		.INIT('h8)
	) name10870 (
		_w21380_,
		_w21381_,
		_w21382_
	);
	LUT2 #(
		.INIT('h1)
	) name10871 (
		wb_rst_i_pad,
		_w21382_,
		_w21383_
	);
	LUT2 #(
		.INIT('h8)
	) name10872 (
		_w12656_,
		_w21383_,
		_w21384_
	);
	LUT2 #(
		.INIT('h1)
	) name10873 (
		_w20871_,
		_w21384_,
		_w21385_
	);
	LUT2 #(
		.INIT('h2)
	) name10874 (
		\wishbone_LatchedTxLength_reg[4]/NET0131 ,
		_w12656_,
		_w21386_
	);
	LUT2 #(
		.INIT('h1)
	) name10875 (
		_w16744_,
		_w21386_,
		_w21387_
	);
	LUT2 #(
		.INIT('h2)
	) name10876 (
		\wishbone_LatchedTxLength_reg[5]/NET0131 ,
		_w12656_,
		_w21388_
	);
	LUT2 #(
		.INIT('h8)
	) name10877 (
		\wishbone_bd_ram_mem2_reg[44][21]/P0001 ,
		_w12896_,
		_w21389_
	);
	LUT2 #(
		.INIT('h8)
	) name10878 (
		\wishbone_bd_ram_mem2_reg[30][21]/P0001 ,
		_w13104_,
		_w21390_
	);
	LUT2 #(
		.INIT('h8)
	) name10879 (
		\wishbone_bd_ram_mem2_reg[171][21]/P0001 ,
		_w12910_,
		_w21391_
	);
	LUT2 #(
		.INIT('h8)
	) name10880 (
		\wishbone_bd_ram_mem2_reg[17][21]/P0001 ,
		_w12848_,
		_w21392_
	);
	LUT2 #(
		.INIT('h8)
	) name10881 (
		\wishbone_bd_ram_mem2_reg[128][21]/P0001 ,
		_w12793_,
		_w21393_
	);
	LUT2 #(
		.INIT('h8)
	) name10882 (
		\wishbone_bd_ram_mem2_reg[255][21]/P0001 ,
		_w13072_,
		_w21394_
	);
	LUT2 #(
		.INIT('h8)
	) name10883 (
		\wishbone_bd_ram_mem2_reg[90][21]/P0001 ,
		_w12978_,
		_w21395_
	);
	LUT2 #(
		.INIT('h8)
	) name10884 (
		\wishbone_bd_ram_mem2_reg[178][21]/P0001 ,
		_w12886_,
		_w21396_
	);
	LUT2 #(
		.INIT('h8)
	) name10885 (
		\wishbone_bd_ram_mem2_reg[60][21]/P0001 ,
		_w13204_,
		_w21397_
	);
	LUT2 #(
		.INIT('h8)
	) name10886 (
		\wishbone_bd_ram_mem2_reg[238][21]/P0001 ,
		_w13160_,
		_w21398_
	);
	LUT2 #(
		.INIT('h8)
	) name10887 (
		\wishbone_bd_ram_mem2_reg[173][21]/P0001 ,
		_w12854_,
		_w21399_
	);
	LUT2 #(
		.INIT('h8)
	) name10888 (
		\wishbone_bd_ram_mem2_reg[94][21]/P0001 ,
		_w13186_,
		_w21400_
	);
	LUT2 #(
		.INIT('h8)
	) name10889 (
		\wishbone_bd_ram_mem2_reg[212][21]/P0001 ,
		_w12796_,
		_w21401_
	);
	LUT2 #(
		.INIT('h8)
	) name10890 (
		\wishbone_bd_ram_mem2_reg[165][21]/P0001 ,
		_w13044_,
		_w21402_
	);
	LUT2 #(
		.INIT('h8)
	) name10891 (
		\wishbone_bd_ram_mem2_reg[102][21]/P0001 ,
		_w12685_,
		_w21403_
	);
	LUT2 #(
		.INIT('h8)
	) name10892 (
		\wishbone_bd_ram_mem2_reg[213][21]/P0001 ,
		_w13002_,
		_w21404_
	);
	LUT2 #(
		.INIT('h8)
	) name10893 (
		\wishbone_bd_ram_mem2_reg[242][21]/P0001 ,
		_w12932_,
		_w21405_
	);
	LUT2 #(
		.INIT('h8)
	) name10894 (
		\wishbone_bd_ram_mem2_reg[111][21]/P0001 ,
		_w12744_,
		_w21406_
	);
	LUT2 #(
		.INIT('h8)
	) name10895 (
		\wishbone_bd_ram_mem2_reg[2][21]/P0001 ,
		_w13088_,
		_w21407_
	);
	LUT2 #(
		.INIT('h8)
	) name10896 (
		\wishbone_bd_ram_mem2_reg[179][21]/P0001 ,
		_w13050_,
		_w21408_
	);
	LUT2 #(
		.INIT('h8)
	) name10897 (
		\wishbone_bd_ram_mem2_reg[148][21]/P0001 ,
		_w13000_,
		_w21409_
	);
	LUT2 #(
		.INIT('h8)
	) name10898 (
		\wishbone_bd_ram_mem2_reg[193][21]/P0001 ,
		_w13056_,
		_w21410_
	);
	LUT2 #(
		.INIT('h8)
	) name10899 (
		\wishbone_bd_ram_mem2_reg[220][21]/P0001 ,
		_w13066_,
		_w21411_
	);
	LUT2 #(
		.INIT('h8)
	) name10900 (
		\wishbone_bd_ram_mem2_reg[230][21]/P0001 ,
		_w13036_,
		_w21412_
	);
	LUT2 #(
		.INIT('h8)
	) name10901 (
		\wishbone_bd_ram_mem2_reg[87][21]/P0001 ,
		_w13154_,
		_w21413_
	);
	LUT2 #(
		.INIT('h8)
	) name10902 (
		\wishbone_bd_ram_mem2_reg[141][21]/P0001 ,
		_w13004_,
		_w21414_
	);
	LUT2 #(
		.INIT('h8)
	) name10903 (
		\wishbone_bd_ram_mem2_reg[8][21]/P0001 ,
		_w12920_,
		_w21415_
	);
	LUT2 #(
		.INIT('h8)
	) name10904 (
		\wishbone_bd_ram_mem2_reg[186][21]/P0001 ,
		_w12783_,
		_w21416_
	);
	LUT2 #(
		.INIT('h8)
	) name10905 (
		\wishbone_bd_ram_mem2_reg[168][21]/P0001 ,
		_w13208_,
		_w21417_
	);
	LUT2 #(
		.INIT('h8)
	) name10906 (
		\wishbone_bd_ram_mem2_reg[115][21]/P0001 ,
		_w13112_,
		_w21418_
	);
	LUT2 #(
		.INIT('h8)
	) name10907 (
		\wishbone_bd_ram_mem2_reg[82][21]/P0001 ,
		_w12942_,
		_w21419_
	);
	LUT2 #(
		.INIT('h8)
	) name10908 (
		\wishbone_bd_ram_mem2_reg[177][21]/P0001 ,
		_w12996_,
		_w21420_
	);
	LUT2 #(
		.INIT('h8)
	) name10909 (
		\wishbone_bd_ram_mem2_reg[51][21]/P0001 ,
		_w13024_,
		_w21421_
	);
	LUT2 #(
		.INIT('h8)
	) name10910 (
		\wishbone_bd_ram_mem2_reg[93][21]/P0001 ,
		_w13016_,
		_w21422_
	);
	LUT2 #(
		.INIT('h8)
	) name10911 (
		\wishbone_bd_ram_mem2_reg[226][21]/P0001 ,
		_w13138_,
		_w21423_
	);
	LUT2 #(
		.INIT('h8)
	) name10912 (
		\wishbone_bd_ram_mem2_reg[176][21]/P0001 ,
		_w12868_,
		_w21424_
	);
	LUT2 #(
		.INIT('h8)
	) name10913 (
		\wishbone_bd_ram_mem2_reg[203][21]/P0001 ,
		_w13158_,
		_w21425_
	);
	LUT2 #(
		.INIT('h8)
	) name10914 (
		\wishbone_bd_ram_mem2_reg[229][21]/P0001 ,
		_w12711_,
		_w21426_
	);
	LUT2 #(
		.INIT('h8)
	) name10915 (
		\wishbone_bd_ram_mem2_reg[116][21]/P0001 ,
		_w12998_,
		_w21427_
	);
	LUT2 #(
		.INIT('h8)
	) name10916 (
		\wishbone_bd_ram_mem2_reg[234][21]/P0001 ,
		_w13214_,
		_w21428_
	);
	LUT2 #(
		.INIT('h8)
	) name10917 (
		\wishbone_bd_ram_mem2_reg[243][21]/P0001 ,
		_w12804_,
		_w21429_
	);
	LUT2 #(
		.INIT('h8)
	) name10918 (
		\wishbone_bd_ram_mem2_reg[248][21]/P0001 ,
		_w12789_,
		_w21430_
	);
	LUT2 #(
		.INIT('h8)
	) name10919 (
		\wishbone_bd_ram_mem2_reg[189][21]/P0001 ,
		_w13042_,
		_w21431_
	);
	LUT2 #(
		.INIT('h8)
	) name10920 (
		\wishbone_bd_ram_mem2_reg[174][21]/P0001 ,
		_w12972_,
		_w21432_
	);
	LUT2 #(
		.INIT('h8)
	) name10921 (
		\wishbone_bd_ram_mem2_reg[121][21]/P0001 ,
		_w13078_,
		_w21433_
	);
	LUT2 #(
		.INIT('h8)
	) name10922 (
		\wishbone_bd_ram_mem2_reg[10][21]/P0001 ,
		_w13172_,
		_w21434_
	);
	LUT2 #(
		.INIT('h8)
	) name10923 (
		\wishbone_bd_ram_mem2_reg[147][21]/P0001 ,
		_w13146_,
		_w21435_
	);
	LUT2 #(
		.INIT('h8)
	) name10924 (
		\wishbone_bd_ram_mem2_reg[206][21]/P0001 ,
		_w12954_,
		_w21436_
	);
	LUT2 #(
		.INIT('h8)
	) name10925 (
		\wishbone_bd_ram_mem2_reg[191][21]/P0001 ,
		_w13034_,
		_w21437_
	);
	LUT2 #(
		.INIT('h8)
	) name10926 (
		\wishbone_bd_ram_mem2_reg[214][21]/P0001 ,
		_w12984_,
		_w21438_
	);
	LUT2 #(
		.INIT('h8)
	) name10927 (
		\wishbone_bd_ram_mem2_reg[120][21]/P0001 ,
		_w12707_,
		_w21439_
	);
	LUT2 #(
		.INIT('h8)
	) name10928 (
		\wishbone_bd_ram_mem2_reg[5][21]/P0001 ,
		_w12878_,
		_w21440_
	);
	LUT2 #(
		.INIT('h8)
	) name10929 (
		\wishbone_bd_ram_mem2_reg[117][21]/P0001 ,
		_w12715_,
		_w21441_
	);
	LUT2 #(
		.INIT('h8)
	) name10930 (
		\wishbone_bd_ram_mem2_reg[100][21]/P0001 ,
		_w12960_,
		_w21442_
	);
	LUT2 #(
		.INIT('h8)
	) name10931 (
		\wishbone_bd_ram_mem2_reg[182][21]/P0001 ,
		_w12820_,
		_w21443_
	);
	LUT2 #(
		.INIT('h8)
	) name10932 (
		\wishbone_bd_ram_mem2_reg[247][21]/P0001 ,
		_w12818_,
		_w21444_
	);
	LUT2 #(
		.INIT('h8)
	) name10933 (
		\wishbone_bd_ram_mem2_reg[108][21]/P0001 ,
		_w13156_,
		_w21445_
	);
	LUT2 #(
		.INIT('h8)
	) name10934 (
		\wishbone_bd_ram_mem2_reg[190][21]/P0001 ,
		_w12858_,
		_w21446_
	);
	LUT2 #(
		.INIT('h8)
	) name10935 (
		\wishbone_bd_ram_mem2_reg[45][21]/P0001 ,
		_w12908_,
		_w21447_
	);
	LUT2 #(
		.INIT('h8)
	) name10936 (
		\wishbone_bd_ram_mem2_reg[15][21]/P0001 ,
		_w13210_,
		_w21448_
	);
	LUT2 #(
		.INIT('h8)
	) name10937 (
		\wishbone_bd_ram_mem2_reg[237][21]/P0001 ,
		_w12990_,
		_w21449_
	);
	LUT2 #(
		.INIT('h8)
	) name10938 (
		\wishbone_bd_ram_mem2_reg[21][21]/P0001 ,
		_w12906_,
		_w21450_
	);
	LUT2 #(
		.INIT('h8)
	) name10939 (
		\wishbone_bd_ram_mem2_reg[134][21]/P0001 ,
		_w12763_,
		_w21451_
	);
	LUT2 #(
		.INIT('h8)
	) name10940 (
		\wishbone_bd_ram_mem2_reg[211][21]/P0001 ,
		_w13166_,
		_w21452_
	);
	LUT2 #(
		.INIT('h8)
	) name10941 (
		\wishbone_bd_ram_mem2_reg[23][21]/P0001 ,
		_w13008_,
		_w21453_
	);
	LUT2 #(
		.INIT('h8)
	) name10942 (
		\wishbone_bd_ram_mem2_reg[143][21]/P0001 ,
		_w12922_,
		_w21454_
	);
	LUT2 #(
		.INIT('h8)
	) name10943 (
		\wishbone_bd_ram_mem2_reg[48][21]/P0001 ,
		_w12970_,
		_w21455_
	);
	LUT2 #(
		.INIT('h8)
	) name10944 (
		\wishbone_bd_ram_mem2_reg[9][21]/P0001 ,
		_w12808_,
		_w21456_
	);
	LUT2 #(
		.INIT('h8)
	) name10945 (
		\wishbone_bd_ram_mem2_reg[64][21]/P0001 ,
		_w12976_,
		_w21457_
	);
	LUT2 #(
		.INIT('h8)
	) name10946 (
		\wishbone_bd_ram_mem2_reg[157][21]/P0001 ,
		_w12926_,
		_w21458_
	);
	LUT2 #(
		.INIT('h8)
	) name10947 (
		\wishbone_bd_ram_mem2_reg[144][21]/P0001 ,
		_w12756_,
		_w21459_
	);
	LUT2 #(
		.INIT('h8)
	) name10948 (
		\wishbone_bd_ram_mem2_reg[155][21]/P0001 ,
		_w13122_,
		_w21460_
	);
	LUT2 #(
		.INIT('h8)
	) name10949 (
		\wishbone_bd_ram_mem2_reg[24][21]/P0001 ,
		_w13084_,
		_w21461_
	);
	LUT2 #(
		.INIT('h8)
	) name10950 (
		\wishbone_bd_ram_mem2_reg[209][21]/P0001 ,
		_w13152_,
		_w21462_
	);
	LUT2 #(
		.INIT('h8)
	) name10951 (
		\wishbone_bd_ram_mem2_reg[149][21]/P0001 ,
		_w12741_,
		_w21463_
	);
	LUT2 #(
		.INIT('h8)
	) name10952 (
		\wishbone_bd_ram_mem2_reg[207][21]/P0001 ,
		_w13180_,
		_w21464_
	);
	LUT2 #(
		.INIT('h8)
	) name10953 (
		\wishbone_bd_ram_mem2_reg[58][21]/P0001 ,
		_w13070_,
		_w21465_
	);
	LUT2 #(
		.INIT('h8)
	) name10954 (
		\wishbone_bd_ram_mem2_reg[198][21]/P0001 ,
		_w12832_,
		_w21466_
	);
	LUT2 #(
		.INIT('h8)
	) name10955 (
		\wishbone_bd_ram_mem2_reg[246][21]/P0001 ,
		_w13076_,
		_w21467_
	);
	LUT2 #(
		.INIT('h8)
	) name10956 (
		\wishbone_bd_ram_mem2_reg[95][21]/P0001 ,
		_w12844_,
		_w21468_
	);
	LUT2 #(
		.INIT('h8)
	) name10957 (
		\wishbone_bd_ram_mem2_reg[101][21]/P0001 ,
		_w13192_,
		_w21469_
	);
	LUT2 #(
		.INIT('h8)
	) name10958 (
		\wishbone_bd_ram_mem2_reg[99][21]/P0001 ,
		_w13038_,
		_w21470_
	);
	LUT2 #(
		.INIT('h8)
	) name10959 (
		\wishbone_bd_ram_mem2_reg[119][21]/P0001 ,
		_w13048_,
		_w21471_
	);
	LUT2 #(
		.INIT('h8)
	) name10960 (
		\wishbone_bd_ram_mem2_reg[145][21]/P0001 ,
		_w13106_,
		_w21472_
	);
	LUT2 #(
		.INIT('h8)
	) name10961 (
		\wishbone_bd_ram_mem2_reg[68][21]/P0001 ,
		_w12946_,
		_w21473_
	);
	LUT2 #(
		.INIT('h8)
	) name10962 (
		\wishbone_bd_ram_mem2_reg[175][21]/P0001 ,
		_w13126_,
		_w21474_
	);
	LUT2 #(
		.INIT('h8)
	) name10963 (
		\wishbone_bd_ram_mem2_reg[37][21]/P0001 ,
		_w13102_,
		_w21475_
	);
	LUT2 #(
		.INIT('h8)
	) name10964 (
		\wishbone_bd_ram_mem2_reg[169][21]/P0001 ,
		_w12722_,
		_w21476_
	);
	LUT2 #(
		.INIT('h8)
	) name10965 (
		\wishbone_bd_ram_mem2_reg[109][21]/P0001 ,
		_w12888_,
		_w21477_
	);
	LUT2 #(
		.INIT('h8)
	) name10966 (
		\wishbone_bd_ram_mem2_reg[122][21]/P0001 ,
		_w13130_,
		_w21478_
	);
	LUT2 #(
		.INIT('h8)
	) name10967 (
		\wishbone_bd_ram_mem2_reg[28][21]/P0001 ,
		_w13170_,
		_w21479_
	);
	LUT2 #(
		.INIT('h8)
	) name10968 (
		\wishbone_bd_ram_mem2_reg[156][21]/P0001 ,
		_w13190_,
		_w21480_
	);
	LUT2 #(
		.INIT('h8)
	) name10969 (
		\wishbone_bd_ram_mem2_reg[254][21]/P0001 ,
		_w12892_,
		_w21481_
	);
	LUT2 #(
		.INIT('h8)
	) name10970 (
		\wishbone_bd_ram_mem2_reg[183][21]/P0001 ,
		_w12787_,
		_w21482_
	);
	LUT2 #(
		.INIT('h8)
	) name10971 (
		\wishbone_bd_ram_mem2_reg[38][21]/P0001 ,
		_w13182_,
		_w21483_
	);
	LUT2 #(
		.INIT('h8)
	) name10972 (
		\wishbone_bd_ram_mem2_reg[232][21]/P0001 ,
		_w12758_,
		_w21484_
	);
	LUT2 #(
		.INIT('h8)
	) name10973 (
		\wishbone_bd_ram_mem2_reg[81][21]/P0001 ,
		_w12950_,
		_w21485_
	);
	LUT2 #(
		.INIT('h8)
	) name10974 (
		\wishbone_bd_ram_mem2_reg[78][21]/P0001 ,
		_w12874_,
		_w21486_
	);
	LUT2 #(
		.INIT('h8)
	) name10975 (
		\wishbone_bd_ram_mem2_reg[50][21]/P0001 ,
		_w13150_,
		_w21487_
	);
	LUT2 #(
		.INIT('h8)
	) name10976 (
		\wishbone_bd_ram_mem2_reg[127][21]/P0001 ,
		_w13164_,
		_w21488_
	);
	LUT2 #(
		.INIT('h8)
	) name10977 (
		\wishbone_bd_ram_mem2_reg[63][21]/P0001 ,
		_w12850_,
		_w21489_
	);
	LUT2 #(
		.INIT('h8)
	) name10978 (
		\wishbone_bd_ram_mem2_reg[125][21]/P0001 ,
		_w12956_,
		_w21490_
	);
	LUT2 #(
		.INIT('h8)
	) name10979 (
		\wishbone_bd_ram_mem2_reg[104][21]/P0001 ,
		_w13148_,
		_w21491_
	);
	LUT2 #(
		.INIT('h8)
	) name10980 (
		\wishbone_bd_ram_mem2_reg[85][21]/P0001 ,
		_w13216_,
		_w21492_
	);
	LUT2 #(
		.INIT('h8)
	) name10981 (
		\wishbone_bd_ram_mem2_reg[162][21]/P0001 ,
		_w13098_,
		_w21493_
	);
	LUT2 #(
		.INIT('h8)
	) name10982 (
		\wishbone_bd_ram_mem2_reg[7][21]/P0001 ,
		_w12728_,
		_w21494_
	);
	LUT2 #(
		.INIT('h8)
	) name10983 (
		\wishbone_bd_ram_mem2_reg[151][21]/P0001 ,
		_w13142_,
		_w21495_
	);
	LUT2 #(
		.INIT('h8)
	) name10984 (
		\wishbone_bd_ram_mem2_reg[62][21]/P0001 ,
		_w12673_,
		_w21496_
	);
	LUT2 #(
		.INIT('h8)
	) name10985 (
		\wishbone_bd_ram_mem2_reg[196][21]/P0001 ,
		_w13090_,
		_w21497_
	);
	LUT2 #(
		.INIT('h8)
	) name10986 (
		\wishbone_bd_ram_mem2_reg[27][21]/P0001 ,
		_w12880_,
		_w21498_
	);
	LUT2 #(
		.INIT('h8)
	) name10987 (
		\wishbone_bd_ram_mem2_reg[22][21]/P0001 ,
		_w13110_,
		_w21499_
	);
	LUT2 #(
		.INIT('h8)
	) name10988 (
		\wishbone_bd_ram_mem2_reg[1][21]/P0001 ,
		_w13014_,
		_w21500_
	);
	LUT2 #(
		.INIT('h8)
	) name10989 (
		\wishbone_bd_ram_mem2_reg[65][21]/P0001 ,
		_w13176_,
		_w21501_
	);
	LUT2 #(
		.INIT('h8)
	) name10990 (
		\wishbone_bd_ram_mem2_reg[77][21]/P0001 ,
		_w12982_,
		_w21502_
	);
	LUT2 #(
		.INIT('h8)
	) name10991 (
		\wishbone_bd_ram_mem2_reg[195][21]/P0001 ,
		_w13144_,
		_w21503_
	);
	LUT2 #(
		.INIT('h8)
	) name10992 (
		\wishbone_bd_ram_mem2_reg[192][21]/P0001 ,
		_w12938_,
		_w21504_
	);
	LUT2 #(
		.INIT('h8)
	) name10993 (
		\wishbone_bd_ram_mem2_reg[114][21]/P0001 ,
		_w13202_,
		_w21505_
	);
	LUT2 #(
		.INIT('h8)
	) name10994 (
		\wishbone_bd_ram_mem2_reg[129][21]/P0001 ,
		_w12776_,
		_w21506_
	);
	LUT2 #(
		.INIT('h8)
	) name10995 (
		\wishbone_bd_ram_mem2_reg[70][21]/P0001 ,
		_w12840_,
		_w21507_
	);
	LUT2 #(
		.INIT('h8)
	) name10996 (
		\wishbone_bd_ram_mem2_reg[166][21]/P0001 ,
		_w13040_,
		_w21508_
	);
	LUT2 #(
		.INIT('h8)
	) name10997 (
		\wishbone_bd_ram_mem2_reg[14][21]/P0001 ,
		_w13086_,
		_w21509_
	);
	LUT2 #(
		.INIT('h8)
	) name10998 (
		\wishbone_bd_ram_mem2_reg[222][21]/P0001 ,
		_w13094_,
		_w21510_
	);
	LUT2 #(
		.INIT('h8)
	) name10999 (
		\wishbone_bd_ram_mem2_reg[40][21]/P0001 ,
		_w13132_,
		_w21511_
	);
	LUT2 #(
		.INIT('h8)
	) name11000 (
		\wishbone_bd_ram_mem2_reg[181][21]/P0001 ,
		_w12828_,
		_w21512_
	);
	LUT2 #(
		.INIT('h8)
	) name11001 (
		\wishbone_bd_ram_mem2_reg[80][21]/P0001 ,
		_w12689_,
		_w21513_
	);
	LUT2 #(
		.INIT('h8)
	) name11002 (
		\wishbone_bd_ram_mem2_reg[210][21]/P0001 ,
		_w12924_,
		_w21514_
	);
	LUT2 #(
		.INIT('h8)
	) name11003 (
		\wishbone_bd_ram_mem2_reg[208][21]/P0001 ,
		_w13032_,
		_w21515_
	);
	LUT2 #(
		.INIT('h8)
	) name11004 (
		\wishbone_bd_ram_mem2_reg[184][21]/P0001 ,
		_w13062_,
		_w21516_
	);
	LUT2 #(
		.INIT('h8)
	) name11005 (
		\wishbone_bd_ram_mem2_reg[224][21]/P0001 ,
		_w12902_,
		_w21517_
	);
	LUT2 #(
		.INIT('h8)
	) name11006 (
		\wishbone_bd_ram_mem2_reg[54][21]/P0001 ,
		_w12770_,
		_w21518_
	);
	LUT2 #(
		.INIT('h8)
	) name11007 (
		\wishbone_bd_ram_mem2_reg[137][21]/P0001 ,
		_w13168_,
		_w21519_
	);
	LUT2 #(
		.INIT('h8)
	) name11008 (
		\wishbone_bd_ram_mem2_reg[172][21]/P0001 ,
		_w12944_,
		_w21520_
	);
	LUT2 #(
		.INIT('h8)
	) name11009 (
		\wishbone_bd_ram_mem2_reg[57][21]/P0001 ,
		_w13116_,
		_w21521_
	);
	LUT2 #(
		.INIT('h8)
	) name11010 (
		\wishbone_bd_ram_mem2_reg[123][21]/P0001 ,
		_w13114_,
		_w21522_
	);
	LUT2 #(
		.INIT('h8)
	) name11011 (
		\wishbone_bd_ram_mem2_reg[3][21]/P0001 ,
		_w12866_,
		_w21523_
	);
	LUT2 #(
		.INIT('h8)
	) name11012 (
		\wishbone_bd_ram_mem2_reg[130][21]/P0001 ,
		_w12914_,
		_w21524_
	);
	LUT2 #(
		.INIT('h8)
	) name11013 (
		\wishbone_bd_ram_mem2_reg[244][21]/P0001 ,
		_w12747_,
		_w21525_
	);
	LUT2 #(
		.INIT('h8)
	) name11014 (
		\wishbone_bd_ram_mem2_reg[49][21]/P0001 ,
		_w12994_,
		_w21526_
	);
	LUT2 #(
		.INIT('h8)
	) name11015 (
		\wishbone_bd_ram_mem2_reg[217][21]/P0001 ,
		_w13188_,
		_w21527_
	);
	LUT2 #(
		.INIT('h8)
	) name11016 (
		\wishbone_bd_ram_mem2_reg[138][21]/P0001 ,
		_w12958_,
		_w21528_
	);
	LUT2 #(
		.INIT('h8)
	) name11017 (
		\wishbone_bd_ram_mem2_reg[56][21]/P0001 ,
		_w12778_,
		_w21529_
	);
	LUT2 #(
		.INIT('h8)
	) name11018 (
		\wishbone_bd_ram_mem2_reg[150][21]/P0001 ,
		_w13136_,
		_w21530_
	);
	LUT2 #(
		.INIT('h8)
	) name11019 (
		\wishbone_bd_ram_mem2_reg[74][21]/P0001 ,
		_w12812_,
		_w21531_
	);
	LUT2 #(
		.INIT('h8)
	) name11020 (
		\wishbone_bd_ram_mem2_reg[79][21]/P0001 ,
		_w13212_,
		_w21532_
	);
	LUT2 #(
		.INIT('h8)
	) name11021 (
		\wishbone_bd_ram_mem2_reg[135][21]/P0001 ,
		_w13124_,
		_w21533_
	);
	LUT2 #(
		.INIT('h8)
	) name11022 (
		\wishbone_bd_ram_mem2_reg[46][21]/P0001 ,
		_w12884_,
		_w21534_
	);
	LUT2 #(
		.INIT('h8)
	) name11023 (
		\wishbone_bd_ram_mem2_reg[47][21]/P0001 ,
		_w12904_,
		_w21535_
	);
	LUT2 #(
		.INIT('h8)
	) name11024 (
		\wishbone_bd_ram_mem2_reg[132][21]/P0001 ,
		_w12992_,
		_w21536_
	);
	LUT2 #(
		.INIT('h8)
	) name11025 (
		\wishbone_bd_ram_mem2_reg[13][21]/P0001 ,
		_w13178_,
		_w21537_
	);
	LUT2 #(
		.INIT('h8)
	) name11026 (
		\wishbone_bd_ram_mem2_reg[241][21]/P0001 ,
		_w13006_,
		_w21538_
	);
	LUT2 #(
		.INIT('h8)
	) name11027 (
		\wishbone_bd_ram_mem2_reg[167][21]/P0001 ,
		_w12986_,
		_w21539_
	);
	LUT2 #(
		.INIT('h8)
	) name11028 (
		\wishbone_bd_ram_mem2_reg[53][21]/P0001 ,
		_w13020_,
		_w21540_
	);
	LUT2 #(
		.INIT('h8)
	) name11029 (
		\wishbone_bd_ram_mem2_reg[227][21]/P0001 ,
		_w12936_,
		_w21541_
	);
	LUT2 #(
		.INIT('h8)
	) name11030 (
		\wishbone_bd_ram_mem2_reg[34][21]/P0001 ,
		_w12930_,
		_w21542_
	);
	LUT2 #(
		.INIT('h8)
	) name11031 (
		\wishbone_bd_ram_mem2_reg[11][21]/P0001 ,
		_w13194_,
		_w21543_
	);
	LUT2 #(
		.INIT('h8)
	) name11032 (
		\wishbone_bd_ram_mem2_reg[131][21]/P0001 ,
		_w12852_,
		_w21544_
	);
	LUT2 #(
		.INIT('h8)
	) name11033 (
		\wishbone_bd_ram_mem2_reg[83][21]/P0001 ,
		_w12916_,
		_w21545_
	);
	LUT2 #(
		.INIT('h8)
	) name11034 (
		\wishbone_bd_ram_mem2_reg[252][21]/P0001 ,
		_w13080_,
		_w21546_
	);
	LUT2 #(
		.INIT('h8)
	) name11035 (
		\wishbone_bd_ram_mem2_reg[154][21]/P0001 ,
		_w12962_,
		_w21547_
	);
	LUT2 #(
		.INIT('h8)
	) name11036 (
		\wishbone_bd_ram_mem2_reg[231][21]/P0001 ,
		_w12856_,
		_w21548_
	);
	LUT2 #(
		.INIT('h8)
	) name11037 (
		\wishbone_bd_ram_mem2_reg[216][21]/P0001 ,
		_w13028_,
		_w21549_
	);
	LUT2 #(
		.INIT('h8)
	) name11038 (
		\wishbone_bd_ram_mem2_reg[170][21]/P0001 ,
		_w13030_,
		_w21550_
	);
	LUT2 #(
		.INIT('h8)
	) name11039 (
		\wishbone_bd_ram_mem2_reg[142][21]/P0001 ,
		_w12928_,
		_w21551_
	);
	LUT2 #(
		.INIT('h8)
	) name11040 (
		\wishbone_bd_ram_mem2_reg[140][21]/P0001 ,
		_w12894_,
		_w21552_
	);
	LUT2 #(
		.INIT('h8)
	) name11041 (
		\wishbone_bd_ram_mem2_reg[146][21]/P0001 ,
		_w13060_,
		_w21553_
	);
	LUT2 #(
		.INIT('h8)
	) name11042 (
		\wishbone_bd_ram_mem2_reg[124][21]/P0001 ,
		_w13058_,
		_w21554_
	);
	LUT2 #(
		.INIT('h8)
	) name11043 (
		\wishbone_bd_ram_mem2_reg[164][21]/P0001 ,
		_w12876_,
		_w21555_
	);
	LUT2 #(
		.INIT('h8)
	) name11044 (
		\wishbone_bd_ram_mem2_reg[52][21]/P0001 ,
		_w13082_,
		_w21556_
	);
	LUT2 #(
		.INIT('h8)
	) name11045 (
		\wishbone_bd_ram_mem2_reg[163][21]/P0001 ,
		_w12882_,
		_w21557_
	);
	LUT2 #(
		.INIT('h8)
	) name11046 (
		\wishbone_bd_ram_mem2_reg[218][21]/P0001 ,
		_w13206_,
		_w21558_
	);
	LUT2 #(
		.INIT('h8)
	) name11047 (
		\wishbone_bd_ram_mem2_reg[180][21]/P0001 ,
		_w12791_,
		_w21559_
	);
	LUT2 #(
		.INIT('h8)
	) name11048 (
		\wishbone_bd_ram_mem2_reg[86][21]/P0001 ,
		_w12735_,
		_w21560_
	);
	LUT2 #(
		.INIT('h8)
	) name11049 (
		\wishbone_bd_ram_mem2_reg[250][21]/P0001 ,
		_w13128_,
		_w21561_
	);
	LUT2 #(
		.INIT('h8)
	) name11050 (
		\wishbone_bd_ram_mem2_reg[225][21]/P0001 ,
		_w13092_,
		_w21562_
	);
	LUT2 #(
		.INIT('h8)
	) name11051 (
		\wishbone_bd_ram_mem2_reg[112][21]/P0001 ,
		_w12733_,
		_w21563_
	);
	LUT2 #(
		.INIT('h8)
	) name11052 (
		\wishbone_bd_ram_mem2_reg[25][21]/P0001 ,
		_w13108_,
		_w21564_
	);
	LUT2 #(
		.INIT('h8)
	) name11053 (
		\wishbone_bd_ram_mem2_reg[29][21]/P0001 ,
		_w12952_,
		_w21565_
	);
	LUT2 #(
		.INIT('h8)
	) name11054 (
		\wishbone_bd_ram_mem2_reg[110][21]/P0001 ,
		_w13046_,
		_w21566_
	);
	LUT2 #(
		.INIT('h8)
	) name11055 (
		\wishbone_bd_ram_mem2_reg[19][21]/P0001 ,
		_w13012_,
		_w21567_
	);
	LUT2 #(
		.INIT('h8)
	) name11056 (
		\wishbone_bd_ram_mem2_reg[204][21]/P0001 ,
		_w13162_,
		_w21568_
	);
	LUT2 #(
		.INIT('h8)
	) name11057 (
		\wishbone_bd_ram_mem2_reg[185][21]/P0001 ,
		_w12940_,
		_w21569_
	);
	LUT2 #(
		.INIT('h8)
	) name11058 (
		\wishbone_bd_ram_mem2_reg[43][21]/P0001 ,
		_w13200_,
		_w21570_
	);
	LUT2 #(
		.INIT('h8)
	) name11059 (
		\wishbone_bd_ram_mem2_reg[69][21]/P0001 ,
		_w12738_,
		_w21571_
	);
	LUT2 #(
		.INIT('h8)
	) name11060 (
		\wishbone_bd_ram_mem2_reg[249][21]/P0001 ,
		_w12900_,
		_w21572_
	);
	LUT2 #(
		.INIT('h8)
	) name11061 (
		\wishbone_bd_ram_mem2_reg[187][21]/P0001 ,
		_w13196_,
		_w21573_
	);
	LUT2 #(
		.INIT('h8)
	) name11062 (
		\wishbone_bd_ram_mem2_reg[67][21]/P0001 ,
		_w13134_,
		_w21574_
	);
	LUT2 #(
		.INIT('h8)
	) name11063 (
		\wishbone_bd_ram_mem2_reg[73][21]/P0001 ,
		_w12918_,
		_w21575_
	);
	LUT2 #(
		.INIT('h8)
	) name11064 (
		\wishbone_bd_ram_mem2_reg[197][21]/P0001 ,
		_w12834_,
		_w21576_
	);
	LUT2 #(
		.INIT('h8)
	) name11065 (
		\wishbone_bd_ram_mem2_reg[4][21]/P0001 ,
		_w12666_,
		_w21577_
	);
	LUT2 #(
		.INIT('h8)
	) name11066 (
		\wishbone_bd_ram_mem2_reg[202][21]/P0001 ,
		_w12870_,
		_w21578_
	);
	LUT2 #(
		.INIT('h8)
	) name11067 (
		\wishbone_bd_ram_mem2_reg[235][21]/P0001 ,
		_w12696_,
		_w21579_
	);
	LUT2 #(
		.INIT('h8)
	) name11068 (
		\wishbone_bd_ram_mem2_reg[159][21]/P0001 ,
		_w12774_,
		_w21580_
	);
	LUT2 #(
		.INIT('h8)
	) name11069 (
		\wishbone_bd_ram_mem2_reg[76][21]/P0001 ,
		_w13184_,
		_w21581_
	);
	LUT2 #(
		.INIT('h8)
	) name11070 (
		\wishbone_bd_ram_mem2_reg[75][21]/P0001 ,
		_w12826_,
		_w21582_
	);
	LUT2 #(
		.INIT('h8)
	) name11071 (
		\wishbone_bd_ram_mem2_reg[71][21]/P0001 ,
		_w12798_,
		_w21583_
	);
	LUT2 #(
		.INIT('h8)
	) name11072 (
		\wishbone_bd_ram_mem2_reg[105][21]/P0001 ,
		_w12751_,
		_w21584_
	);
	LUT2 #(
		.INIT('h8)
	) name11073 (
		\wishbone_bd_ram_mem2_reg[201][21]/P0001 ,
		_w12822_,
		_w21585_
	);
	LUT2 #(
		.INIT('h8)
	) name11074 (
		\wishbone_bd_ram_mem2_reg[33][21]/P0001 ,
		_w12980_,
		_w21586_
	);
	LUT2 #(
		.INIT('h8)
	) name11075 (
		\wishbone_bd_ram_mem2_reg[223][21]/P0001 ,
		_w12838_,
		_w21587_
	);
	LUT2 #(
		.INIT('h8)
	) name11076 (
		\wishbone_bd_ram_mem2_reg[72][21]/P0001 ,
		_w12810_,
		_w21588_
	);
	LUT2 #(
		.INIT('h8)
	) name11077 (
		\wishbone_bd_ram_mem2_reg[188][21]/P0001 ,
		_w12948_,
		_w21589_
	);
	LUT2 #(
		.INIT('h8)
	) name11078 (
		\wishbone_bd_ram_mem2_reg[158][21]/P0001 ,
		_w12898_,
		_w21590_
	);
	LUT2 #(
		.INIT('h8)
	) name11079 (
		\wishbone_bd_ram_mem2_reg[239][21]/P0001 ,
		_w12862_,
		_w21591_
	);
	LUT2 #(
		.INIT('h8)
	) name11080 (
		\wishbone_bd_ram_mem2_reg[91][21]/P0001 ,
		_w13074_,
		_w21592_
	);
	LUT2 #(
		.INIT('h8)
	) name11081 (
		\wishbone_bd_ram_mem2_reg[236][21]/P0001 ,
		_w12731_,
		_w21593_
	);
	LUT2 #(
		.INIT('h8)
	) name11082 (
		\wishbone_bd_ram_mem2_reg[199][21]/P0001 ,
		_w12768_,
		_w21594_
	);
	LUT2 #(
		.INIT('h8)
	) name11083 (
		\wishbone_bd_ram_mem2_reg[66][21]/P0001 ,
		_w12824_,
		_w21595_
	);
	LUT2 #(
		.INIT('h8)
	) name11084 (
		\wishbone_bd_ram_mem2_reg[31][21]/P0001 ,
		_w13198_,
		_w21596_
	);
	LUT2 #(
		.INIT('h8)
	) name11085 (
		\wishbone_bd_ram_mem2_reg[12][21]/P0001 ,
		_w13118_,
		_w21597_
	);
	LUT2 #(
		.INIT('h8)
	) name11086 (
		\wishbone_bd_ram_mem2_reg[20][21]/P0001 ,
		_w13174_,
		_w21598_
	);
	LUT2 #(
		.INIT('h8)
	) name11087 (
		\wishbone_bd_ram_mem2_reg[221][21]/P0001 ,
		_w12802_,
		_w21599_
	);
	LUT2 #(
		.INIT('h8)
	) name11088 (
		\wishbone_bd_ram_mem2_reg[35][21]/P0001 ,
		_w12703_,
		_w21600_
	);
	LUT2 #(
		.INIT('h8)
	) name11089 (
		\wishbone_bd_ram_mem2_reg[42][21]/P0001 ,
		_w12842_,
		_w21601_
	);
	LUT2 #(
		.INIT('h8)
	) name11090 (
		\wishbone_bd_ram_mem2_reg[26][21]/P0001 ,
		_w12699_,
		_w21602_
	);
	LUT2 #(
		.INIT('h8)
	) name11091 (
		\wishbone_bd_ram_mem2_reg[152][21]/P0001 ,
		_w12966_,
		_w21603_
	);
	LUT2 #(
		.INIT('h8)
	) name11092 (
		\wishbone_bd_ram_mem2_reg[233][21]/P0001 ,
		_w12836_,
		_w21604_
	);
	LUT2 #(
		.INIT('h8)
	) name11093 (
		\wishbone_bd_ram_mem2_reg[160][21]/P0001 ,
		_w12872_,
		_w21605_
	);
	LUT2 #(
		.INIT('h8)
	) name11094 (
		\wishbone_bd_ram_mem2_reg[61][21]/P0001 ,
		_w12725_,
		_w21606_
	);
	LUT2 #(
		.INIT('h8)
	) name11095 (
		\wishbone_bd_ram_mem2_reg[136][21]/P0001 ,
		_w13064_,
		_w21607_
	);
	LUT2 #(
		.INIT('h8)
	) name11096 (
		\wishbone_bd_ram_mem2_reg[41][21]/P0001 ,
		_w13052_,
		_w21608_
	);
	LUT2 #(
		.INIT('h8)
	) name11097 (
		\wishbone_bd_ram_mem2_reg[84][21]/P0001 ,
		_w12934_,
		_w21609_
	);
	LUT2 #(
		.INIT('h8)
	) name11098 (
		\wishbone_bd_ram_mem2_reg[153][21]/P0001 ,
		_w12890_,
		_w21610_
	);
	LUT2 #(
		.INIT('h8)
	) name11099 (
		\wishbone_bd_ram_mem2_reg[106][21]/P0001 ,
		_w12713_,
		_w21611_
	);
	LUT2 #(
		.INIT('h8)
	) name11100 (
		\wishbone_bd_ram_mem2_reg[92][21]/P0001 ,
		_w13010_,
		_w21612_
	);
	LUT2 #(
		.INIT('h8)
	) name11101 (
		\wishbone_bd_ram_mem2_reg[98][21]/P0001 ,
		_w12816_,
		_w21613_
	);
	LUT2 #(
		.INIT('h8)
	) name11102 (
		\wishbone_bd_ram_mem2_reg[200][21]/P0001 ,
		_w12988_,
		_w21614_
	);
	LUT2 #(
		.INIT('h8)
	) name11103 (
		\wishbone_bd_ram_mem2_reg[59][21]/P0001 ,
		_w12780_,
		_w21615_
	);
	LUT2 #(
		.INIT('h8)
	) name11104 (
		\wishbone_bd_ram_mem2_reg[113][21]/P0001 ,
		_w13026_,
		_w21616_
	);
	LUT2 #(
		.INIT('h8)
	) name11105 (
		\wishbone_bd_ram_mem2_reg[118][21]/P0001 ,
		_w12830_,
		_w21617_
	);
	LUT2 #(
		.INIT('h8)
	) name11106 (
		\wishbone_bd_ram_mem2_reg[16][21]/P0001 ,
		_w13140_,
		_w21618_
	);
	LUT2 #(
		.INIT('h8)
	) name11107 (
		\wishbone_bd_ram_mem2_reg[6][21]/P0001 ,
		_w12968_,
		_w21619_
	);
	LUT2 #(
		.INIT('h8)
	) name11108 (
		\wishbone_bd_ram_mem2_reg[139][21]/P0001 ,
		_w12814_,
		_w21620_
	);
	LUT2 #(
		.INIT('h8)
	) name11109 (
		\wishbone_bd_ram_mem2_reg[97][21]/P0001 ,
		_w13096_,
		_w21621_
	);
	LUT2 #(
		.INIT('h8)
	) name11110 (
		\wishbone_bd_ram_mem2_reg[89][21]/P0001 ,
		_w12964_,
		_w21622_
	);
	LUT2 #(
		.INIT('h8)
	) name11111 (
		\wishbone_bd_ram_mem2_reg[0][21]/P0001 ,
		_w12717_,
		_w21623_
	);
	LUT2 #(
		.INIT('h8)
	) name11112 (
		\wishbone_bd_ram_mem2_reg[107][21]/P0001 ,
		_w12749_,
		_w21624_
	);
	LUT2 #(
		.INIT('h8)
	) name11113 (
		\wishbone_bd_ram_mem2_reg[253][21]/P0001 ,
		_w13100_,
		_w21625_
	);
	LUT2 #(
		.INIT('h8)
	) name11114 (
		\wishbone_bd_ram_mem2_reg[39][21]/P0001 ,
		_w13018_,
		_w21626_
	);
	LUT2 #(
		.INIT('h8)
	) name11115 (
		\wishbone_bd_ram_mem2_reg[194][21]/P0001 ,
		_w12772_,
		_w21627_
	);
	LUT2 #(
		.INIT('h8)
	) name11116 (
		\wishbone_bd_ram_mem2_reg[133][21]/P0001 ,
		_w12761_,
		_w21628_
	);
	LUT2 #(
		.INIT('h8)
	) name11117 (
		\wishbone_bd_ram_mem2_reg[219][21]/P0001 ,
		_w12806_,
		_w21629_
	);
	LUT2 #(
		.INIT('h8)
	) name11118 (
		\wishbone_bd_ram_mem2_reg[103][21]/P0001 ,
		_w12846_,
		_w21630_
	);
	LUT2 #(
		.INIT('h8)
	) name11119 (
		\wishbone_bd_ram_mem2_reg[245][21]/P0001 ,
		_w13022_,
		_w21631_
	);
	LUT2 #(
		.INIT('h8)
	) name11120 (
		\wishbone_bd_ram_mem2_reg[251][21]/P0001 ,
		_w13054_,
		_w21632_
	);
	LUT2 #(
		.INIT('h8)
	) name11121 (
		\wishbone_bd_ram_mem2_reg[240][21]/P0001 ,
		_w12864_,
		_w21633_
	);
	LUT2 #(
		.INIT('h8)
	) name11122 (
		\wishbone_bd_ram_mem2_reg[32][21]/P0001 ,
		_w13120_,
		_w21634_
	);
	LUT2 #(
		.INIT('h8)
	) name11123 (
		\wishbone_bd_ram_mem2_reg[88][21]/P0001 ,
		_w12860_,
		_w21635_
	);
	LUT2 #(
		.INIT('h8)
	) name11124 (
		\wishbone_bd_ram_mem2_reg[205][21]/P0001 ,
		_w13068_,
		_w21636_
	);
	LUT2 #(
		.INIT('h8)
	) name11125 (
		\wishbone_bd_ram_mem2_reg[161][21]/P0001 ,
		_w12754_,
		_w21637_
	);
	LUT2 #(
		.INIT('h8)
	) name11126 (
		\wishbone_bd_ram_mem2_reg[36][21]/P0001 ,
		_w12800_,
		_w21638_
	);
	LUT2 #(
		.INIT('h8)
	) name11127 (
		\wishbone_bd_ram_mem2_reg[55][21]/P0001 ,
		_w12785_,
		_w21639_
	);
	LUT2 #(
		.INIT('h8)
	) name11128 (
		\wishbone_bd_ram_mem2_reg[215][21]/P0001 ,
		_w12974_,
		_w21640_
	);
	LUT2 #(
		.INIT('h8)
	) name11129 (
		\wishbone_bd_ram_mem2_reg[96][21]/P0001 ,
		_w12912_,
		_w21641_
	);
	LUT2 #(
		.INIT('h8)
	) name11130 (
		\wishbone_bd_ram_mem2_reg[228][21]/P0001 ,
		_w12765_,
		_w21642_
	);
	LUT2 #(
		.INIT('h8)
	) name11131 (
		\wishbone_bd_ram_mem2_reg[18][21]/P0001 ,
		_w12679_,
		_w21643_
	);
	LUT2 #(
		.INIT('h8)
	) name11132 (
		\wishbone_bd_ram_mem2_reg[126][21]/P0001 ,
		_w13218_,
		_w21644_
	);
	LUT2 #(
		.INIT('h1)
	) name11133 (
		_w21389_,
		_w21390_,
		_w21645_
	);
	LUT2 #(
		.INIT('h1)
	) name11134 (
		_w21391_,
		_w21392_,
		_w21646_
	);
	LUT2 #(
		.INIT('h1)
	) name11135 (
		_w21393_,
		_w21394_,
		_w21647_
	);
	LUT2 #(
		.INIT('h1)
	) name11136 (
		_w21395_,
		_w21396_,
		_w21648_
	);
	LUT2 #(
		.INIT('h1)
	) name11137 (
		_w21397_,
		_w21398_,
		_w21649_
	);
	LUT2 #(
		.INIT('h1)
	) name11138 (
		_w21399_,
		_w21400_,
		_w21650_
	);
	LUT2 #(
		.INIT('h1)
	) name11139 (
		_w21401_,
		_w21402_,
		_w21651_
	);
	LUT2 #(
		.INIT('h1)
	) name11140 (
		_w21403_,
		_w21404_,
		_w21652_
	);
	LUT2 #(
		.INIT('h1)
	) name11141 (
		_w21405_,
		_w21406_,
		_w21653_
	);
	LUT2 #(
		.INIT('h1)
	) name11142 (
		_w21407_,
		_w21408_,
		_w21654_
	);
	LUT2 #(
		.INIT('h1)
	) name11143 (
		_w21409_,
		_w21410_,
		_w21655_
	);
	LUT2 #(
		.INIT('h1)
	) name11144 (
		_w21411_,
		_w21412_,
		_w21656_
	);
	LUT2 #(
		.INIT('h1)
	) name11145 (
		_w21413_,
		_w21414_,
		_w21657_
	);
	LUT2 #(
		.INIT('h1)
	) name11146 (
		_w21415_,
		_w21416_,
		_w21658_
	);
	LUT2 #(
		.INIT('h1)
	) name11147 (
		_w21417_,
		_w21418_,
		_w21659_
	);
	LUT2 #(
		.INIT('h1)
	) name11148 (
		_w21419_,
		_w21420_,
		_w21660_
	);
	LUT2 #(
		.INIT('h1)
	) name11149 (
		_w21421_,
		_w21422_,
		_w21661_
	);
	LUT2 #(
		.INIT('h1)
	) name11150 (
		_w21423_,
		_w21424_,
		_w21662_
	);
	LUT2 #(
		.INIT('h1)
	) name11151 (
		_w21425_,
		_w21426_,
		_w21663_
	);
	LUT2 #(
		.INIT('h1)
	) name11152 (
		_w21427_,
		_w21428_,
		_w21664_
	);
	LUT2 #(
		.INIT('h1)
	) name11153 (
		_w21429_,
		_w21430_,
		_w21665_
	);
	LUT2 #(
		.INIT('h1)
	) name11154 (
		_w21431_,
		_w21432_,
		_w21666_
	);
	LUT2 #(
		.INIT('h1)
	) name11155 (
		_w21433_,
		_w21434_,
		_w21667_
	);
	LUT2 #(
		.INIT('h1)
	) name11156 (
		_w21435_,
		_w21436_,
		_w21668_
	);
	LUT2 #(
		.INIT('h1)
	) name11157 (
		_w21437_,
		_w21438_,
		_w21669_
	);
	LUT2 #(
		.INIT('h1)
	) name11158 (
		_w21439_,
		_w21440_,
		_w21670_
	);
	LUT2 #(
		.INIT('h1)
	) name11159 (
		_w21441_,
		_w21442_,
		_w21671_
	);
	LUT2 #(
		.INIT('h1)
	) name11160 (
		_w21443_,
		_w21444_,
		_w21672_
	);
	LUT2 #(
		.INIT('h1)
	) name11161 (
		_w21445_,
		_w21446_,
		_w21673_
	);
	LUT2 #(
		.INIT('h1)
	) name11162 (
		_w21447_,
		_w21448_,
		_w21674_
	);
	LUT2 #(
		.INIT('h1)
	) name11163 (
		_w21449_,
		_w21450_,
		_w21675_
	);
	LUT2 #(
		.INIT('h1)
	) name11164 (
		_w21451_,
		_w21452_,
		_w21676_
	);
	LUT2 #(
		.INIT('h1)
	) name11165 (
		_w21453_,
		_w21454_,
		_w21677_
	);
	LUT2 #(
		.INIT('h1)
	) name11166 (
		_w21455_,
		_w21456_,
		_w21678_
	);
	LUT2 #(
		.INIT('h1)
	) name11167 (
		_w21457_,
		_w21458_,
		_w21679_
	);
	LUT2 #(
		.INIT('h1)
	) name11168 (
		_w21459_,
		_w21460_,
		_w21680_
	);
	LUT2 #(
		.INIT('h1)
	) name11169 (
		_w21461_,
		_w21462_,
		_w21681_
	);
	LUT2 #(
		.INIT('h1)
	) name11170 (
		_w21463_,
		_w21464_,
		_w21682_
	);
	LUT2 #(
		.INIT('h1)
	) name11171 (
		_w21465_,
		_w21466_,
		_w21683_
	);
	LUT2 #(
		.INIT('h1)
	) name11172 (
		_w21467_,
		_w21468_,
		_w21684_
	);
	LUT2 #(
		.INIT('h1)
	) name11173 (
		_w21469_,
		_w21470_,
		_w21685_
	);
	LUT2 #(
		.INIT('h1)
	) name11174 (
		_w21471_,
		_w21472_,
		_w21686_
	);
	LUT2 #(
		.INIT('h1)
	) name11175 (
		_w21473_,
		_w21474_,
		_w21687_
	);
	LUT2 #(
		.INIT('h1)
	) name11176 (
		_w21475_,
		_w21476_,
		_w21688_
	);
	LUT2 #(
		.INIT('h1)
	) name11177 (
		_w21477_,
		_w21478_,
		_w21689_
	);
	LUT2 #(
		.INIT('h1)
	) name11178 (
		_w21479_,
		_w21480_,
		_w21690_
	);
	LUT2 #(
		.INIT('h1)
	) name11179 (
		_w21481_,
		_w21482_,
		_w21691_
	);
	LUT2 #(
		.INIT('h1)
	) name11180 (
		_w21483_,
		_w21484_,
		_w21692_
	);
	LUT2 #(
		.INIT('h1)
	) name11181 (
		_w21485_,
		_w21486_,
		_w21693_
	);
	LUT2 #(
		.INIT('h1)
	) name11182 (
		_w21487_,
		_w21488_,
		_w21694_
	);
	LUT2 #(
		.INIT('h1)
	) name11183 (
		_w21489_,
		_w21490_,
		_w21695_
	);
	LUT2 #(
		.INIT('h1)
	) name11184 (
		_w21491_,
		_w21492_,
		_w21696_
	);
	LUT2 #(
		.INIT('h1)
	) name11185 (
		_w21493_,
		_w21494_,
		_w21697_
	);
	LUT2 #(
		.INIT('h1)
	) name11186 (
		_w21495_,
		_w21496_,
		_w21698_
	);
	LUT2 #(
		.INIT('h1)
	) name11187 (
		_w21497_,
		_w21498_,
		_w21699_
	);
	LUT2 #(
		.INIT('h1)
	) name11188 (
		_w21499_,
		_w21500_,
		_w21700_
	);
	LUT2 #(
		.INIT('h1)
	) name11189 (
		_w21501_,
		_w21502_,
		_w21701_
	);
	LUT2 #(
		.INIT('h1)
	) name11190 (
		_w21503_,
		_w21504_,
		_w21702_
	);
	LUT2 #(
		.INIT('h1)
	) name11191 (
		_w21505_,
		_w21506_,
		_w21703_
	);
	LUT2 #(
		.INIT('h1)
	) name11192 (
		_w21507_,
		_w21508_,
		_w21704_
	);
	LUT2 #(
		.INIT('h1)
	) name11193 (
		_w21509_,
		_w21510_,
		_w21705_
	);
	LUT2 #(
		.INIT('h1)
	) name11194 (
		_w21511_,
		_w21512_,
		_w21706_
	);
	LUT2 #(
		.INIT('h1)
	) name11195 (
		_w21513_,
		_w21514_,
		_w21707_
	);
	LUT2 #(
		.INIT('h1)
	) name11196 (
		_w21515_,
		_w21516_,
		_w21708_
	);
	LUT2 #(
		.INIT('h1)
	) name11197 (
		_w21517_,
		_w21518_,
		_w21709_
	);
	LUT2 #(
		.INIT('h1)
	) name11198 (
		_w21519_,
		_w21520_,
		_w21710_
	);
	LUT2 #(
		.INIT('h1)
	) name11199 (
		_w21521_,
		_w21522_,
		_w21711_
	);
	LUT2 #(
		.INIT('h1)
	) name11200 (
		_w21523_,
		_w21524_,
		_w21712_
	);
	LUT2 #(
		.INIT('h1)
	) name11201 (
		_w21525_,
		_w21526_,
		_w21713_
	);
	LUT2 #(
		.INIT('h1)
	) name11202 (
		_w21527_,
		_w21528_,
		_w21714_
	);
	LUT2 #(
		.INIT('h1)
	) name11203 (
		_w21529_,
		_w21530_,
		_w21715_
	);
	LUT2 #(
		.INIT('h1)
	) name11204 (
		_w21531_,
		_w21532_,
		_w21716_
	);
	LUT2 #(
		.INIT('h1)
	) name11205 (
		_w21533_,
		_w21534_,
		_w21717_
	);
	LUT2 #(
		.INIT('h1)
	) name11206 (
		_w21535_,
		_w21536_,
		_w21718_
	);
	LUT2 #(
		.INIT('h1)
	) name11207 (
		_w21537_,
		_w21538_,
		_w21719_
	);
	LUT2 #(
		.INIT('h1)
	) name11208 (
		_w21539_,
		_w21540_,
		_w21720_
	);
	LUT2 #(
		.INIT('h1)
	) name11209 (
		_w21541_,
		_w21542_,
		_w21721_
	);
	LUT2 #(
		.INIT('h1)
	) name11210 (
		_w21543_,
		_w21544_,
		_w21722_
	);
	LUT2 #(
		.INIT('h1)
	) name11211 (
		_w21545_,
		_w21546_,
		_w21723_
	);
	LUT2 #(
		.INIT('h1)
	) name11212 (
		_w21547_,
		_w21548_,
		_w21724_
	);
	LUT2 #(
		.INIT('h1)
	) name11213 (
		_w21549_,
		_w21550_,
		_w21725_
	);
	LUT2 #(
		.INIT('h1)
	) name11214 (
		_w21551_,
		_w21552_,
		_w21726_
	);
	LUT2 #(
		.INIT('h1)
	) name11215 (
		_w21553_,
		_w21554_,
		_w21727_
	);
	LUT2 #(
		.INIT('h1)
	) name11216 (
		_w21555_,
		_w21556_,
		_w21728_
	);
	LUT2 #(
		.INIT('h1)
	) name11217 (
		_w21557_,
		_w21558_,
		_w21729_
	);
	LUT2 #(
		.INIT('h1)
	) name11218 (
		_w21559_,
		_w21560_,
		_w21730_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		_w21561_,
		_w21562_,
		_w21731_
	);
	LUT2 #(
		.INIT('h1)
	) name11220 (
		_w21563_,
		_w21564_,
		_w21732_
	);
	LUT2 #(
		.INIT('h1)
	) name11221 (
		_w21565_,
		_w21566_,
		_w21733_
	);
	LUT2 #(
		.INIT('h1)
	) name11222 (
		_w21567_,
		_w21568_,
		_w21734_
	);
	LUT2 #(
		.INIT('h1)
	) name11223 (
		_w21569_,
		_w21570_,
		_w21735_
	);
	LUT2 #(
		.INIT('h1)
	) name11224 (
		_w21571_,
		_w21572_,
		_w21736_
	);
	LUT2 #(
		.INIT('h1)
	) name11225 (
		_w21573_,
		_w21574_,
		_w21737_
	);
	LUT2 #(
		.INIT('h1)
	) name11226 (
		_w21575_,
		_w21576_,
		_w21738_
	);
	LUT2 #(
		.INIT('h1)
	) name11227 (
		_w21577_,
		_w21578_,
		_w21739_
	);
	LUT2 #(
		.INIT('h1)
	) name11228 (
		_w21579_,
		_w21580_,
		_w21740_
	);
	LUT2 #(
		.INIT('h1)
	) name11229 (
		_w21581_,
		_w21582_,
		_w21741_
	);
	LUT2 #(
		.INIT('h1)
	) name11230 (
		_w21583_,
		_w21584_,
		_w21742_
	);
	LUT2 #(
		.INIT('h1)
	) name11231 (
		_w21585_,
		_w21586_,
		_w21743_
	);
	LUT2 #(
		.INIT('h1)
	) name11232 (
		_w21587_,
		_w21588_,
		_w21744_
	);
	LUT2 #(
		.INIT('h1)
	) name11233 (
		_w21589_,
		_w21590_,
		_w21745_
	);
	LUT2 #(
		.INIT('h1)
	) name11234 (
		_w21591_,
		_w21592_,
		_w21746_
	);
	LUT2 #(
		.INIT('h1)
	) name11235 (
		_w21593_,
		_w21594_,
		_w21747_
	);
	LUT2 #(
		.INIT('h1)
	) name11236 (
		_w21595_,
		_w21596_,
		_w21748_
	);
	LUT2 #(
		.INIT('h1)
	) name11237 (
		_w21597_,
		_w21598_,
		_w21749_
	);
	LUT2 #(
		.INIT('h1)
	) name11238 (
		_w21599_,
		_w21600_,
		_w21750_
	);
	LUT2 #(
		.INIT('h1)
	) name11239 (
		_w21601_,
		_w21602_,
		_w21751_
	);
	LUT2 #(
		.INIT('h1)
	) name11240 (
		_w21603_,
		_w21604_,
		_w21752_
	);
	LUT2 #(
		.INIT('h1)
	) name11241 (
		_w21605_,
		_w21606_,
		_w21753_
	);
	LUT2 #(
		.INIT('h1)
	) name11242 (
		_w21607_,
		_w21608_,
		_w21754_
	);
	LUT2 #(
		.INIT('h1)
	) name11243 (
		_w21609_,
		_w21610_,
		_w21755_
	);
	LUT2 #(
		.INIT('h1)
	) name11244 (
		_w21611_,
		_w21612_,
		_w21756_
	);
	LUT2 #(
		.INIT('h1)
	) name11245 (
		_w21613_,
		_w21614_,
		_w21757_
	);
	LUT2 #(
		.INIT('h1)
	) name11246 (
		_w21615_,
		_w21616_,
		_w21758_
	);
	LUT2 #(
		.INIT('h1)
	) name11247 (
		_w21617_,
		_w21618_,
		_w21759_
	);
	LUT2 #(
		.INIT('h1)
	) name11248 (
		_w21619_,
		_w21620_,
		_w21760_
	);
	LUT2 #(
		.INIT('h1)
	) name11249 (
		_w21621_,
		_w21622_,
		_w21761_
	);
	LUT2 #(
		.INIT('h1)
	) name11250 (
		_w21623_,
		_w21624_,
		_w21762_
	);
	LUT2 #(
		.INIT('h1)
	) name11251 (
		_w21625_,
		_w21626_,
		_w21763_
	);
	LUT2 #(
		.INIT('h1)
	) name11252 (
		_w21627_,
		_w21628_,
		_w21764_
	);
	LUT2 #(
		.INIT('h1)
	) name11253 (
		_w21629_,
		_w21630_,
		_w21765_
	);
	LUT2 #(
		.INIT('h1)
	) name11254 (
		_w21631_,
		_w21632_,
		_w21766_
	);
	LUT2 #(
		.INIT('h1)
	) name11255 (
		_w21633_,
		_w21634_,
		_w21767_
	);
	LUT2 #(
		.INIT('h1)
	) name11256 (
		_w21635_,
		_w21636_,
		_w21768_
	);
	LUT2 #(
		.INIT('h1)
	) name11257 (
		_w21637_,
		_w21638_,
		_w21769_
	);
	LUT2 #(
		.INIT('h1)
	) name11258 (
		_w21639_,
		_w21640_,
		_w21770_
	);
	LUT2 #(
		.INIT('h1)
	) name11259 (
		_w21641_,
		_w21642_,
		_w21771_
	);
	LUT2 #(
		.INIT('h1)
	) name11260 (
		_w21643_,
		_w21644_,
		_w21772_
	);
	LUT2 #(
		.INIT('h8)
	) name11261 (
		_w21771_,
		_w21772_,
		_w21773_
	);
	LUT2 #(
		.INIT('h8)
	) name11262 (
		_w21769_,
		_w21770_,
		_w21774_
	);
	LUT2 #(
		.INIT('h8)
	) name11263 (
		_w21767_,
		_w21768_,
		_w21775_
	);
	LUT2 #(
		.INIT('h8)
	) name11264 (
		_w21765_,
		_w21766_,
		_w21776_
	);
	LUT2 #(
		.INIT('h8)
	) name11265 (
		_w21763_,
		_w21764_,
		_w21777_
	);
	LUT2 #(
		.INIT('h8)
	) name11266 (
		_w21761_,
		_w21762_,
		_w21778_
	);
	LUT2 #(
		.INIT('h8)
	) name11267 (
		_w21759_,
		_w21760_,
		_w21779_
	);
	LUT2 #(
		.INIT('h8)
	) name11268 (
		_w21757_,
		_w21758_,
		_w21780_
	);
	LUT2 #(
		.INIT('h8)
	) name11269 (
		_w21755_,
		_w21756_,
		_w21781_
	);
	LUT2 #(
		.INIT('h8)
	) name11270 (
		_w21753_,
		_w21754_,
		_w21782_
	);
	LUT2 #(
		.INIT('h8)
	) name11271 (
		_w21751_,
		_w21752_,
		_w21783_
	);
	LUT2 #(
		.INIT('h8)
	) name11272 (
		_w21749_,
		_w21750_,
		_w21784_
	);
	LUT2 #(
		.INIT('h8)
	) name11273 (
		_w21747_,
		_w21748_,
		_w21785_
	);
	LUT2 #(
		.INIT('h8)
	) name11274 (
		_w21745_,
		_w21746_,
		_w21786_
	);
	LUT2 #(
		.INIT('h8)
	) name11275 (
		_w21743_,
		_w21744_,
		_w21787_
	);
	LUT2 #(
		.INIT('h8)
	) name11276 (
		_w21741_,
		_w21742_,
		_w21788_
	);
	LUT2 #(
		.INIT('h8)
	) name11277 (
		_w21739_,
		_w21740_,
		_w21789_
	);
	LUT2 #(
		.INIT('h8)
	) name11278 (
		_w21737_,
		_w21738_,
		_w21790_
	);
	LUT2 #(
		.INIT('h8)
	) name11279 (
		_w21735_,
		_w21736_,
		_w21791_
	);
	LUT2 #(
		.INIT('h8)
	) name11280 (
		_w21733_,
		_w21734_,
		_w21792_
	);
	LUT2 #(
		.INIT('h8)
	) name11281 (
		_w21731_,
		_w21732_,
		_w21793_
	);
	LUT2 #(
		.INIT('h8)
	) name11282 (
		_w21729_,
		_w21730_,
		_w21794_
	);
	LUT2 #(
		.INIT('h8)
	) name11283 (
		_w21727_,
		_w21728_,
		_w21795_
	);
	LUT2 #(
		.INIT('h8)
	) name11284 (
		_w21725_,
		_w21726_,
		_w21796_
	);
	LUT2 #(
		.INIT('h8)
	) name11285 (
		_w21723_,
		_w21724_,
		_w21797_
	);
	LUT2 #(
		.INIT('h8)
	) name11286 (
		_w21721_,
		_w21722_,
		_w21798_
	);
	LUT2 #(
		.INIT('h8)
	) name11287 (
		_w21719_,
		_w21720_,
		_w21799_
	);
	LUT2 #(
		.INIT('h8)
	) name11288 (
		_w21717_,
		_w21718_,
		_w21800_
	);
	LUT2 #(
		.INIT('h8)
	) name11289 (
		_w21715_,
		_w21716_,
		_w21801_
	);
	LUT2 #(
		.INIT('h8)
	) name11290 (
		_w21713_,
		_w21714_,
		_w21802_
	);
	LUT2 #(
		.INIT('h8)
	) name11291 (
		_w21711_,
		_w21712_,
		_w21803_
	);
	LUT2 #(
		.INIT('h8)
	) name11292 (
		_w21709_,
		_w21710_,
		_w21804_
	);
	LUT2 #(
		.INIT('h8)
	) name11293 (
		_w21707_,
		_w21708_,
		_w21805_
	);
	LUT2 #(
		.INIT('h8)
	) name11294 (
		_w21705_,
		_w21706_,
		_w21806_
	);
	LUT2 #(
		.INIT('h8)
	) name11295 (
		_w21703_,
		_w21704_,
		_w21807_
	);
	LUT2 #(
		.INIT('h8)
	) name11296 (
		_w21701_,
		_w21702_,
		_w21808_
	);
	LUT2 #(
		.INIT('h8)
	) name11297 (
		_w21699_,
		_w21700_,
		_w21809_
	);
	LUT2 #(
		.INIT('h8)
	) name11298 (
		_w21697_,
		_w21698_,
		_w21810_
	);
	LUT2 #(
		.INIT('h8)
	) name11299 (
		_w21695_,
		_w21696_,
		_w21811_
	);
	LUT2 #(
		.INIT('h8)
	) name11300 (
		_w21693_,
		_w21694_,
		_w21812_
	);
	LUT2 #(
		.INIT('h8)
	) name11301 (
		_w21691_,
		_w21692_,
		_w21813_
	);
	LUT2 #(
		.INIT('h8)
	) name11302 (
		_w21689_,
		_w21690_,
		_w21814_
	);
	LUT2 #(
		.INIT('h8)
	) name11303 (
		_w21687_,
		_w21688_,
		_w21815_
	);
	LUT2 #(
		.INIT('h8)
	) name11304 (
		_w21685_,
		_w21686_,
		_w21816_
	);
	LUT2 #(
		.INIT('h8)
	) name11305 (
		_w21683_,
		_w21684_,
		_w21817_
	);
	LUT2 #(
		.INIT('h8)
	) name11306 (
		_w21681_,
		_w21682_,
		_w21818_
	);
	LUT2 #(
		.INIT('h8)
	) name11307 (
		_w21679_,
		_w21680_,
		_w21819_
	);
	LUT2 #(
		.INIT('h8)
	) name11308 (
		_w21677_,
		_w21678_,
		_w21820_
	);
	LUT2 #(
		.INIT('h8)
	) name11309 (
		_w21675_,
		_w21676_,
		_w21821_
	);
	LUT2 #(
		.INIT('h8)
	) name11310 (
		_w21673_,
		_w21674_,
		_w21822_
	);
	LUT2 #(
		.INIT('h8)
	) name11311 (
		_w21671_,
		_w21672_,
		_w21823_
	);
	LUT2 #(
		.INIT('h8)
	) name11312 (
		_w21669_,
		_w21670_,
		_w21824_
	);
	LUT2 #(
		.INIT('h8)
	) name11313 (
		_w21667_,
		_w21668_,
		_w21825_
	);
	LUT2 #(
		.INIT('h8)
	) name11314 (
		_w21665_,
		_w21666_,
		_w21826_
	);
	LUT2 #(
		.INIT('h8)
	) name11315 (
		_w21663_,
		_w21664_,
		_w21827_
	);
	LUT2 #(
		.INIT('h8)
	) name11316 (
		_w21661_,
		_w21662_,
		_w21828_
	);
	LUT2 #(
		.INIT('h8)
	) name11317 (
		_w21659_,
		_w21660_,
		_w21829_
	);
	LUT2 #(
		.INIT('h8)
	) name11318 (
		_w21657_,
		_w21658_,
		_w21830_
	);
	LUT2 #(
		.INIT('h8)
	) name11319 (
		_w21655_,
		_w21656_,
		_w21831_
	);
	LUT2 #(
		.INIT('h8)
	) name11320 (
		_w21653_,
		_w21654_,
		_w21832_
	);
	LUT2 #(
		.INIT('h8)
	) name11321 (
		_w21651_,
		_w21652_,
		_w21833_
	);
	LUT2 #(
		.INIT('h8)
	) name11322 (
		_w21649_,
		_w21650_,
		_w21834_
	);
	LUT2 #(
		.INIT('h8)
	) name11323 (
		_w21647_,
		_w21648_,
		_w21835_
	);
	LUT2 #(
		.INIT('h8)
	) name11324 (
		_w21645_,
		_w21646_,
		_w21836_
	);
	LUT2 #(
		.INIT('h8)
	) name11325 (
		_w21835_,
		_w21836_,
		_w21837_
	);
	LUT2 #(
		.INIT('h8)
	) name11326 (
		_w21833_,
		_w21834_,
		_w21838_
	);
	LUT2 #(
		.INIT('h8)
	) name11327 (
		_w21831_,
		_w21832_,
		_w21839_
	);
	LUT2 #(
		.INIT('h8)
	) name11328 (
		_w21829_,
		_w21830_,
		_w21840_
	);
	LUT2 #(
		.INIT('h8)
	) name11329 (
		_w21827_,
		_w21828_,
		_w21841_
	);
	LUT2 #(
		.INIT('h8)
	) name11330 (
		_w21825_,
		_w21826_,
		_w21842_
	);
	LUT2 #(
		.INIT('h8)
	) name11331 (
		_w21823_,
		_w21824_,
		_w21843_
	);
	LUT2 #(
		.INIT('h8)
	) name11332 (
		_w21821_,
		_w21822_,
		_w21844_
	);
	LUT2 #(
		.INIT('h8)
	) name11333 (
		_w21819_,
		_w21820_,
		_w21845_
	);
	LUT2 #(
		.INIT('h8)
	) name11334 (
		_w21817_,
		_w21818_,
		_w21846_
	);
	LUT2 #(
		.INIT('h8)
	) name11335 (
		_w21815_,
		_w21816_,
		_w21847_
	);
	LUT2 #(
		.INIT('h8)
	) name11336 (
		_w21813_,
		_w21814_,
		_w21848_
	);
	LUT2 #(
		.INIT('h8)
	) name11337 (
		_w21811_,
		_w21812_,
		_w21849_
	);
	LUT2 #(
		.INIT('h8)
	) name11338 (
		_w21809_,
		_w21810_,
		_w21850_
	);
	LUT2 #(
		.INIT('h8)
	) name11339 (
		_w21807_,
		_w21808_,
		_w21851_
	);
	LUT2 #(
		.INIT('h8)
	) name11340 (
		_w21805_,
		_w21806_,
		_w21852_
	);
	LUT2 #(
		.INIT('h8)
	) name11341 (
		_w21803_,
		_w21804_,
		_w21853_
	);
	LUT2 #(
		.INIT('h8)
	) name11342 (
		_w21801_,
		_w21802_,
		_w21854_
	);
	LUT2 #(
		.INIT('h8)
	) name11343 (
		_w21799_,
		_w21800_,
		_w21855_
	);
	LUT2 #(
		.INIT('h8)
	) name11344 (
		_w21797_,
		_w21798_,
		_w21856_
	);
	LUT2 #(
		.INIT('h8)
	) name11345 (
		_w21795_,
		_w21796_,
		_w21857_
	);
	LUT2 #(
		.INIT('h8)
	) name11346 (
		_w21793_,
		_w21794_,
		_w21858_
	);
	LUT2 #(
		.INIT('h8)
	) name11347 (
		_w21791_,
		_w21792_,
		_w21859_
	);
	LUT2 #(
		.INIT('h8)
	) name11348 (
		_w21789_,
		_w21790_,
		_w21860_
	);
	LUT2 #(
		.INIT('h8)
	) name11349 (
		_w21787_,
		_w21788_,
		_w21861_
	);
	LUT2 #(
		.INIT('h8)
	) name11350 (
		_w21785_,
		_w21786_,
		_w21862_
	);
	LUT2 #(
		.INIT('h8)
	) name11351 (
		_w21783_,
		_w21784_,
		_w21863_
	);
	LUT2 #(
		.INIT('h8)
	) name11352 (
		_w21781_,
		_w21782_,
		_w21864_
	);
	LUT2 #(
		.INIT('h8)
	) name11353 (
		_w21779_,
		_w21780_,
		_w21865_
	);
	LUT2 #(
		.INIT('h8)
	) name11354 (
		_w21777_,
		_w21778_,
		_w21866_
	);
	LUT2 #(
		.INIT('h8)
	) name11355 (
		_w21775_,
		_w21776_,
		_w21867_
	);
	LUT2 #(
		.INIT('h8)
	) name11356 (
		_w21773_,
		_w21774_,
		_w21868_
	);
	LUT2 #(
		.INIT('h8)
	) name11357 (
		_w21867_,
		_w21868_,
		_w21869_
	);
	LUT2 #(
		.INIT('h8)
	) name11358 (
		_w21865_,
		_w21866_,
		_w21870_
	);
	LUT2 #(
		.INIT('h8)
	) name11359 (
		_w21863_,
		_w21864_,
		_w21871_
	);
	LUT2 #(
		.INIT('h8)
	) name11360 (
		_w21861_,
		_w21862_,
		_w21872_
	);
	LUT2 #(
		.INIT('h8)
	) name11361 (
		_w21859_,
		_w21860_,
		_w21873_
	);
	LUT2 #(
		.INIT('h8)
	) name11362 (
		_w21857_,
		_w21858_,
		_w21874_
	);
	LUT2 #(
		.INIT('h8)
	) name11363 (
		_w21855_,
		_w21856_,
		_w21875_
	);
	LUT2 #(
		.INIT('h8)
	) name11364 (
		_w21853_,
		_w21854_,
		_w21876_
	);
	LUT2 #(
		.INIT('h8)
	) name11365 (
		_w21851_,
		_w21852_,
		_w21877_
	);
	LUT2 #(
		.INIT('h8)
	) name11366 (
		_w21849_,
		_w21850_,
		_w21878_
	);
	LUT2 #(
		.INIT('h8)
	) name11367 (
		_w21847_,
		_w21848_,
		_w21879_
	);
	LUT2 #(
		.INIT('h8)
	) name11368 (
		_w21845_,
		_w21846_,
		_w21880_
	);
	LUT2 #(
		.INIT('h8)
	) name11369 (
		_w21843_,
		_w21844_,
		_w21881_
	);
	LUT2 #(
		.INIT('h8)
	) name11370 (
		_w21841_,
		_w21842_,
		_w21882_
	);
	LUT2 #(
		.INIT('h8)
	) name11371 (
		_w21839_,
		_w21840_,
		_w21883_
	);
	LUT2 #(
		.INIT('h8)
	) name11372 (
		_w21837_,
		_w21838_,
		_w21884_
	);
	LUT2 #(
		.INIT('h8)
	) name11373 (
		_w21883_,
		_w21884_,
		_w21885_
	);
	LUT2 #(
		.INIT('h8)
	) name11374 (
		_w21881_,
		_w21882_,
		_w21886_
	);
	LUT2 #(
		.INIT('h8)
	) name11375 (
		_w21879_,
		_w21880_,
		_w21887_
	);
	LUT2 #(
		.INIT('h8)
	) name11376 (
		_w21877_,
		_w21878_,
		_w21888_
	);
	LUT2 #(
		.INIT('h8)
	) name11377 (
		_w21875_,
		_w21876_,
		_w21889_
	);
	LUT2 #(
		.INIT('h8)
	) name11378 (
		_w21873_,
		_w21874_,
		_w21890_
	);
	LUT2 #(
		.INIT('h8)
	) name11379 (
		_w21871_,
		_w21872_,
		_w21891_
	);
	LUT2 #(
		.INIT('h8)
	) name11380 (
		_w21869_,
		_w21870_,
		_w21892_
	);
	LUT2 #(
		.INIT('h8)
	) name11381 (
		_w21891_,
		_w21892_,
		_w21893_
	);
	LUT2 #(
		.INIT('h8)
	) name11382 (
		_w21889_,
		_w21890_,
		_w21894_
	);
	LUT2 #(
		.INIT('h8)
	) name11383 (
		_w21887_,
		_w21888_,
		_w21895_
	);
	LUT2 #(
		.INIT('h8)
	) name11384 (
		_w21885_,
		_w21886_,
		_w21896_
	);
	LUT2 #(
		.INIT('h8)
	) name11385 (
		_w21895_,
		_w21896_,
		_w21897_
	);
	LUT2 #(
		.INIT('h8)
	) name11386 (
		_w21893_,
		_w21894_,
		_w21898_
	);
	LUT2 #(
		.INIT('h8)
	) name11387 (
		_w21897_,
		_w21898_,
		_w21899_
	);
	LUT2 #(
		.INIT('h1)
	) name11388 (
		wb_rst_i_pad,
		_w21899_,
		_w21900_
	);
	LUT2 #(
		.INIT('h8)
	) name11389 (
		_w12656_,
		_w21900_,
		_w21901_
	);
	LUT2 #(
		.INIT('h1)
	) name11390 (
		_w21388_,
		_w21901_,
		_w21902_
	);
	LUT2 #(
		.INIT('h2)
	) name11391 (
		\wishbone_LatchedTxLength_reg[7]/NET0131 ,
		_w12656_,
		_w21903_
	);
	LUT2 #(
		.INIT('h8)
	) name11392 (
		\wishbone_bd_ram_mem2_reg[43][23]/P0001 ,
		_w13200_,
		_w21904_
	);
	LUT2 #(
		.INIT('h8)
	) name11393 (
		\wishbone_bd_ram_mem2_reg[18][23]/P0001 ,
		_w12679_,
		_w21905_
	);
	LUT2 #(
		.INIT('h8)
	) name11394 (
		\wishbone_bd_ram_mem2_reg[236][23]/P0001 ,
		_w12731_,
		_w21906_
	);
	LUT2 #(
		.INIT('h8)
	) name11395 (
		\wishbone_bd_ram_mem2_reg[102][23]/P0001 ,
		_w12685_,
		_w21907_
	);
	LUT2 #(
		.INIT('h8)
	) name11396 (
		\wishbone_bd_ram_mem2_reg[189][23]/P0001 ,
		_w13042_,
		_w21908_
	);
	LUT2 #(
		.INIT('h8)
	) name11397 (
		\wishbone_bd_ram_mem2_reg[197][23]/P0001 ,
		_w12834_,
		_w21909_
	);
	LUT2 #(
		.INIT('h8)
	) name11398 (
		\wishbone_bd_ram_mem2_reg[72][23]/P0001 ,
		_w12810_,
		_w21910_
	);
	LUT2 #(
		.INIT('h8)
	) name11399 (
		\wishbone_bd_ram_mem2_reg[6][23]/P0001 ,
		_w12968_,
		_w21911_
	);
	LUT2 #(
		.INIT('h8)
	) name11400 (
		\wishbone_bd_ram_mem2_reg[141][23]/P0001 ,
		_w13004_,
		_w21912_
	);
	LUT2 #(
		.INIT('h8)
	) name11401 (
		\wishbone_bd_ram_mem2_reg[238][23]/P0001 ,
		_w13160_,
		_w21913_
	);
	LUT2 #(
		.INIT('h8)
	) name11402 (
		\wishbone_bd_ram_mem2_reg[114][23]/P0001 ,
		_w13202_,
		_w21914_
	);
	LUT2 #(
		.INIT('h8)
	) name11403 (
		\wishbone_bd_ram_mem2_reg[75][23]/P0001 ,
		_w12826_,
		_w21915_
	);
	LUT2 #(
		.INIT('h8)
	) name11404 (
		\wishbone_bd_ram_mem2_reg[235][23]/P0001 ,
		_w12696_,
		_w21916_
	);
	LUT2 #(
		.INIT('h8)
	) name11405 (
		\wishbone_bd_ram_mem2_reg[112][23]/P0001 ,
		_w12733_,
		_w21917_
	);
	LUT2 #(
		.INIT('h8)
	) name11406 (
		\wishbone_bd_ram_mem2_reg[34][23]/P0001 ,
		_w12930_,
		_w21918_
	);
	LUT2 #(
		.INIT('h8)
	) name11407 (
		\wishbone_bd_ram_mem2_reg[251][23]/P0001 ,
		_w13054_,
		_w21919_
	);
	LUT2 #(
		.INIT('h8)
	) name11408 (
		\wishbone_bd_ram_mem2_reg[243][23]/P0001 ,
		_w12804_,
		_w21920_
	);
	LUT2 #(
		.INIT('h8)
	) name11409 (
		\wishbone_bd_ram_mem2_reg[70][23]/P0001 ,
		_w12840_,
		_w21921_
	);
	LUT2 #(
		.INIT('h8)
	) name11410 (
		\wishbone_bd_ram_mem2_reg[161][23]/P0001 ,
		_w12754_,
		_w21922_
	);
	LUT2 #(
		.INIT('h8)
	) name11411 (
		\wishbone_bd_ram_mem2_reg[29][23]/P0001 ,
		_w12952_,
		_w21923_
	);
	LUT2 #(
		.INIT('h8)
	) name11412 (
		\wishbone_bd_ram_mem2_reg[157][23]/P0001 ,
		_w12926_,
		_w21924_
	);
	LUT2 #(
		.INIT('h8)
	) name11413 (
		\wishbone_bd_ram_mem2_reg[105][23]/P0001 ,
		_w12751_,
		_w21925_
	);
	LUT2 #(
		.INIT('h8)
	) name11414 (
		\wishbone_bd_ram_mem2_reg[220][23]/P0001 ,
		_w13066_,
		_w21926_
	);
	LUT2 #(
		.INIT('h8)
	) name11415 (
		\wishbone_bd_ram_mem2_reg[125][23]/P0001 ,
		_w12956_,
		_w21927_
	);
	LUT2 #(
		.INIT('h8)
	) name11416 (
		\wishbone_bd_ram_mem2_reg[111][23]/P0001 ,
		_w12744_,
		_w21928_
	);
	LUT2 #(
		.INIT('h8)
	) name11417 (
		\wishbone_bd_ram_mem2_reg[160][23]/P0001 ,
		_w12872_,
		_w21929_
	);
	LUT2 #(
		.INIT('h8)
	) name11418 (
		\wishbone_bd_ram_mem2_reg[192][23]/P0001 ,
		_w12938_,
		_w21930_
	);
	LUT2 #(
		.INIT('h8)
	) name11419 (
		\wishbone_bd_ram_mem2_reg[159][23]/P0001 ,
		_w12774_,
		_w21931_
	);
	LUT2 #(
		.INIT('h8)
	) name11420 (
		\wishbone_bd_ram_mem2_reg[82][23]/P0001 ,
		_w12942_,
		_w21932_
	);
	LUT2 #(
		.INIT('h8)
	) name11421 (
		\wishbone_bd_ram_mem2_reg[55][23]/P0001 ,
		_w12785_,
		_w21933_
	);
	LUT2 #(
		.INIT('h8)
	) name11422 (
		\wishbone_bd_ram_mem2_reg[81][23]/P0001 ,
		_w12950_,
		_w21934_
	);
	LUT2 #(
		.INIT('h8)
	) name11423 (
		\wishbone_bd_ram_mem2_reg[223][23]/P0001 ,
		_w12838_,
		_w21935_
	);
	LUT2 #(
		.INIT('h8)
	) name11424 (
		\wishbone_bd_ram_mem2_reg[54][23]/P0001 ,
		_w12770_,
		_w21936_
	);
	LUT2 #(
		.INIT('h8)
	) name11425 (
		\wishbone_bd_ram_mem2_reg[234][23]/P0001 ,
		_w13214_,
		_w21937_
	);
	LUT2 #(
		.INIT('h8)
	) name11426 (
		\wishbone_bd_ram_mem2_reg[222][23]/P0001 ,
		_w13094_,
		_w21938_
	);
	LUT2 #(
		.INIT('h8)
	) name11427 (
		\wishbone_bd_ram_mem2_reg[73][23]/P0001 ,
		_w12918_,
		_w21939_
	);
	LUT2 #(
		.INIT('h8)
	) name11428 (
		\wishbone_bd_ram_mem2_reg[56][23]/P0001 ,
		_w12778_,
		_w21940_
	);
	LUT2 #(
		.INIT('h8)
	) name11429 (
		\wishbone_bd_ram_mem2_reg[59][23]/P0001 ,
		_w12780_,
		_w21941_
	);
	LUT2 #(
		.INIT('h8)
	) name11430 (
		\wishbone_bd_ram_mem2_reg[129][23]/P0001 ,
		_w12776_,
		_w21942_
	);
	LUT2 #(
		.INIT('h8)
	) name11431 (
		\wishbone_bd_ram_mem2_reg[245][23]/P0001 ,
		_w13022_,
		_w21943_
	);
	LUT2 #(
		.INIT('h8)
	) name11432 (
		\wishbone_bd_ram_mem2_reg[242][23]/P0001 ,
		_w12932_,
		_w21944_
	);
	LUT2 #(
		.INIT('h8)
	) name11433 (
		\wishbone_bd_ram_mem2_reg[214][23]/P0001 ,
		_w12984_,
		_w21945_
	);
	LUT2 #(
		.INIT('h8)
	) name11434 (
		\wishbone_bd_ram_mem2_reg[20][23]/P0001 ,
		_w13174_,
		_w21946_
	);
	LUT2 #(
		.INIT('h8)
	) name11435 (
		\wishbone_bd_ram_mem2_reg[65][23]/P0001 ,
		_w13176_,
		_w21947_
	);
	LUT2 #(
		.INIT('h8)
	) name11436 (
		\wishbone_bd_ram_mem2_reg[140][23]/P0001 ,
		_w12894_,
		_w21948_
	);
	LUT2 #(
		.INIT('h8)
	) name11437 (
		\wishbone_bd_ram_mem2_reg[87][23]/P0001 ,
		_w13154_,
		_w21949_
	);
	LUT2 #(
		.INIT('h8)
	) name11438 (
		\wishbone_bd_ram_mem2_reg[51][23]/P0001 ,
		_w13024_,
		_w21950_
	);
	LUT2 #(
		.INIT('h8)
	) name11439 (
		\wishbone_bd_ram_mem2_reg[250][23]/P0001 ,
		_w13128_,
		_w21951_
	);
	LUT2 #(
		.INIT('h8)
	) name11440 (
		\wishbone_bd_ram_mem2_reg[211][23]/P0001 ,
		_w13166_,
		_w21952_
	);
	LUT2 #(
		.INIT('h8)
	) name11441 (
		\wishbone_bd_ram_mem2_reg[240][23]/P0001 ,
		_w12864_,
		_w21953_
	);
	LUT2 #(
		.INIT('h8)
	) name11442 (
		\wishbone_bd_ram_mem2_reg[255][23]/P0001 ,
		_w13072_,
		_w21954_
	);
	LUT2 #(
		.INIT('h8)
	) name11443 (
		\wishbone_bd_ram_mem2_reg[135][23]/P0001 ,
		_w13124_,
		_w21955_
	);
	LUT2 #(
		.INIT('h8)
	) name11444 (
		\wishbone_bd_ram_mem2_reg[109][23]/P0001 ,
		_w12888_,
		_w21956_
	);
	LUT2 #(
		.INIT('h8)
	) name11445 (
		\wishbone_bd_ram_mem2_reg[142][23]/P0001 ,
		_w12928_,
		_w21957_
	);
	LUT2 #(
		.INIT('h8)
	) name11446 (
		\wishbone_bd_ram_mem2_reg[104][23]/P0001 ,
		_w13148_,
		_w21958_
	);
	LUT2 #(
		.INIT('h8)
	) name11447 (
		\wishbone_bd_ram_mem2_reg[151][23]/P0001 ,
		_w13142_,
		_w21959_
	);
	LUT2 #(
		.INIT('h8)
	) name11448 (
		\wishbone_bd_ram_mem2_reg[164][23]/P0001 ,
		_w12876_,
		_w21960_
	);
	LUT2 #(
		.INIT('h8)
	) name11449 (
		\wishbone_bd_ram_mem2_reg[133][23]/P0001 ,
		_w12761_,
		_w21961_
	);
	LUT2 #(
		.INIT('h8)
	) name11450 (
		\wishbone_bd_ram_mem2_reg[163][23]/P0001 ,
		_w12882_,
		_w21962_
	);
	LUT2 #(
		.INIT('h8)
	) name11451 (
		\wishbone_bd_ram_mem2_reg[136][23]/P0001 ,
		_w13064_,
		_w21963_
	);
	LUT2 #(
		.INIT('h8)
	) name11452 (
		\wishbone_bd_ram_mem2_reg[181][23]/P0001 ,
		_w12828_,
		_w21964_
	);
	LUT2 #(
		.INIT('h8)
	) name11453 (
		\wishbone_bd_ram_mem2_reg[144][23]/P0001 ,
		_w12756_,
		_w21965_
	);
	LUT2 #(
		.INIT('h8)
	) name11454 (
		\wishbone_bd_ram_mem2_reg[134][23]/P0001 ,
		_w12763_,
		_w21966_
	);
	LUT2 #(
		.INIT('h8)
	) name11455 (
		\wishbone_bd_ram_mem2_reg[107][23]/P0001 ,
		_w12749_,
		_w21967_
	);
	LUT2 #(
		.INIT('h8)
	) name11456 (
		\wishbone_bd_ram_mem2_reg[249][23]/P0001 ,
		_w12900_,
		_w21968_
	);
	LUT2 #(
		.INIT('h8)
	) name11457 (
		\wishbone_bd_ram_mem2_reg[179][23]/P0001 ,
		_w13050_,
		_w21969_
	);
	LUT2 #(
		.INIT('h8)
	) name11458 (
		\wishbone_bd_ram_mem2_reg[66][23]/P0001 ,
		_w12824_,
		_w21970_
	);
	LUT2 #(
		.INIT('h8)
	) name11459 (
		\wishbone_bd_ram_mem2_reg[180][23]/P0001 ,
		_w12791_,
		_w21971_
	);
	LUT2 #(
		.INIT('h8)
	) name11460 (
		\wishbone_bd_ram_mem2_reg[88][23]/P0001 ,
		_w12860_,
		_w21972_
	);
	LUT2 #(
		.INIT('h8)
	) name11461 (
		\wishbone_bd_ram_mem2_reg[103][23]/P0001 ,
		_w12846_,
		_w21973_
	);
	LUT2 #(
		.INIT('h8)
	) name11462 (
		\wishbone_bd_ram_mem2_reg[61][23]/P0001 ,
		_w12725_,
		_w21974_
	);
	LUT2 #(
		.INIT('h8)
	) name11463 (
		\wishbone_bd_ram_mem2_reg[53][23]/P0001 ,
		_w13020_,
		_w21975_
	);
	LUT2 #(
		.INIT('h8)
	) name11464 (
		\wishbone_bd_ram_mem2_reg[166][23]/P0001 ,
		_w13040_,
		_w21976_
	);
	LUT2 #(
		.INIT('h8)
	) name11465 (
		\wishbone_bd_ram_mem2_reg[126][23]/P0001 ,
		_w13218_,
		_w21977_
	);
	LUT2 #(
		.INIT('h8)
	) name11466 (
		\wishbone_bd_ram_mem2_reg[153][23]/P0001 ,
		_w12890_,
		_w21978_
	);
	LUT2 #(
		.INIT('h8)
	) name11467 (
		\wishbone_bd_ram_mem2_reg[201][23]/P0001 ,
		_w12822_,
		_w21979_
	);
	LUT2 #(
		.INIT('h8)
	) name11468 (
		\wishbone_bd_ram_mem2_reg[3][23]/P0001 ,
		_w12866_,
		_w21980_
	);
	LUT2 #(
		.INIT('h8)
	) name11469 (
		\wishbone_bd_ram_mem2_reg[194][23]/P0001 ,
		_w12772_,
		_w21981_
	);
	LUT2 #(
		.INIT('h8)
	) name11470 (
		\wishbone_bd_ram_mem2_reg[219][23]/P0001 ,
		_w12806_,
		_w21982_
	);
	LUT2 #(
		.INIT('h8)
	) name11471 (
		\wishbone_bd_ram_mem2_reg[79][23]/P0001 ,
		_w13212_,
		_w21983_
	);
	LUT2 #(
		.INIT('h8)
	) name11472 (
		\wishbone_bd_ram_mem2_reg[139][23]/P0001 ,
		_w12814_,
		_w21984_
	);
	LUT2 #(
		.INIT('h8)
	) name11473 (
		\wishbone_bd_ram_mem2_reg[35][23]/P0001 ,
		_w12703_,
		_w21985_
	);
	LUT2 #(
		.INIT('h8)
	) name11474 (
		\wishbone_bd_ram_mem2_reg[5][23]/P0001 ,
		_w12878_,
		_w21986_
	);
	LUT2 #(
		.INIT('h8)
	) name11475 (
		\wishbone_bd_ram_mem2_reg[199][23]/P0001 ,
		_w12768_,
		_w21987_
	);
	LUT2 #(
		.INIT('h8)
	) name11476 (
		\wishbone_bd_ram_mem2_reg[38][23]/P0001 ,
		_w13182_,
		_w21988_
	);
	LUT2 #(
		.INIT('h8)
	) name11477 (
		\wishbone_bd_ram_mem2_reg[85][23]/P0001 ,
		_w13216_,
		_w21989_
	);
	LUT2 #(
		.INIT('h8)
	) name11478 (
		\wishbone_bd_ram_mem2_reg[50][23]/P0001 ,
		_w13150_,
		_w21990_
	);
	LUT2 #(
		.INIT('h8)
	) name11479 (
		\wishbone_bd_ram_mem2_reg[31][23]/P0001 ,
		_w13198_,
		_w21991_
	);
	LUT2 #(
		.INIT('h8)
	) name11480 (
		\wishbone_bd_ram_mem2_reg[11][23]/P0001 ,
		_w13194_,
		_w21992_
	);
	LUT2 #(
		.INIT('h8)
	) name11481 (
		\wishbone_bd_ram_mem2_reg[178][23]/P0001 ,
		_w12886_,
		_w21993_
	);
	LUT2 #(
		.INIT('h8)
	) name11482 (
		\wishbone_bd_ram_mem2_reg[210][23]/P0001 ,
		_w12924_,
		_w21994_
	);
	LUT2 #(
		.INIT('h8)
	) name11483 (
		\wishbone_bd_ram_mem2_reg[231][23]/P0001 ,
		_w12856_,
		_w21995_
	);
	LUT2 #(
		.INIT('h8)
	) name11484 (
		\wishbone_bd_ram_mem2_reg[202][23]/P0001 ,
		_w12870_,
		_w21996_
	);
	LUT2 #(
		.INIT('h8)
	) name11485 (
		\wishbone_bd_ram_mem2_reg[191][23]/P0001 ,
		_w13034_,
		_w21997_
	);
	LUT2 #(
		.INIT('h8)
	) name11486 (
		\wishbone_bd_ram_mem2_reg[68][23]/P0001 ,
		_w12946_,
		_w21998_
	);
	LUT2 #(
		.INIT('h8)
	) name11487 (
		\wishbone_bd_ram_mem2_reg[228][23]/P0001 ,
		_w12765_,
		_w21999_
	);
	LUT2 #(
		.INIT('h8)
	) name11488 (
		\wishbone_bd_ram_mem2_reg[213][23]/P0001 ,
		_w13002_,
		_w22000_
	);
	LUT2 #(
		.INIT('h8)
	) name11489 (
		\wishbone_bd_ram_mem2_reg[212][23]/P0001 ,
		_w12796_,
		_w22001_
	);
	LUT2 #(
		.INIT('h8)
	) name11490 (
		\wishbone_bd_ram_mem2_reg[47][23]/P0001 ,
		_w12904_,
		_w22002_
	);
	LUT2 #(
		.INIT('h8)
	) name11491 (
		\wishbone_bd_ram_mem2_reg[1][23]/P0001 ,
		_w13014_,
		_w22003_
	);
	LUT2 #(
		.INIT('h8)
	) name11492 (
		\wishbone_bd_ram_mem2_reg[92][23]/P0001 ,
		_w13010_,
		_w22004_
	);
	LUT2 #(
		.INIT('h8)
	) name11493 (
		\wishbone_bd_ram_mem2_reg[230][23]/P0001 ,
		_w13036_,
		_w22005_
	);
	LUT2 #(
		.INIT('h8)
	) name11494 (
		\wishbone_bd_ram_mem2_reg[182][23]/P0001 ,
		_w12820_,
		_w22006_
	);
	LUT2 #(
		.INIT('h8)
	) name11495 (
		\wishbone_bd_ram_mem2_reg[80][23]/P0001 ,
		_w12689_,
		_w22007_
	);
	LUT2 #(
		.INIT('h8)
	) name11496 (
		\wishbone_bd_ram_mem2_reg[97][23]/P0001 ,
		_w13096_,
		_w22008_
	);
	LUT2 #(
		.INIT('h8)
	) name11497 (
		\wishbone_bd_ram_mem2_reg[138][23]/P0001 ,
		_w12958_,
		_w22009_
	);
	LUT2 #(
		.INIT('h8)
	) name11498 (
		\wishbone_bd_ram_mem2_reg[8][23]/P0001 ,
		_w12920_,
		_w22010_
	);
	LUT2 #(
		.INIT('h8)
	) name11499 (
		\wishbone_bd_ram_mem2_reg[62][23]/P0001 ,
		_w12673_,
		_w22011_
	);
	LUT2 #(
		.INIT('h8)
	) name11500 (
		\wishbone_bd_ram_mem2_reg[123][23]/P0001 ,
		_w13114_,
		_w22012_
	);
	LUT2 #(
		.INIT('h8)
	) name11501 (
		\wishbone_bd_ram_mem2_reg[149][23]/P0001 ,
		_w12741_,
		_w22013_
	);
	LUT2 #(
		.INIT('h8)
	) name11502 (
		\wishbone_bd_ram_mem2_reg[7][23]/P0001 ,
		_w12728_,
		_w22014_
	);
	LUT2 #(
		.INIT('h8)
	) name11503 (
		\wishbone_bd_ram_mem2_reg[203][23]/P0001 ,
		_w13158_,
		_w22015_
	);
	LUT2 #(
		.INIT('h8)
	) name11504 (
		\wishbone_bd_ram_mem2_reg[175][23]/P0001 ,
		_w13126_,
		_w22016_
	);
	LUT2 #(
		.INIT('h8)
	) name11505 (
		\wishbone_bd_ram_mem2_reg[64][23]/P0001 ,
		_w12976_,
		_w22017_
	);
	LUT2 #(
		.INIT('h8)
	) name11506 (
		\wishbone_bd_ram_mem2_reg[239][23]/P0001 ,
		_w12862_,
		_w22018_
	);
	LUT2 #(
		.INIT('h8)
	) name11507 (
		\wishbone_bd_ram_mem2_reg[118][23]/P0001 ,
		_w12830_,
		_w22019_
	);
	LUT2 #(
		.INIT('h8)
	) name11508 (
		\wishbone_bd_ram_mem2_reg[209][23]/P0001 ,
		_w13152_,
		_w22020_
	);
	LUT2 #(
		.INIT('h8)
	) name11509 (
		\wishbone_bd_ram_mem2_reg[196][23]/P0001 ,
		_w13090_,
		_w22021_
	);
	LUT2 #(
		.INIT('h8)
	) name11510 (
		\wishbone_bd_ram_mem2_reg[10][23]/P0001 ,
		_w13172_,
		_w22022_
	);
	LUT2 #(
		.INIT('h8)
	) name11511 (
		\wishbone_bd_ram_mem2_reg[24][23]/P0001 ,
		_w13084_,
		_w22023_
	);
	LUT2 #(
		.INIT('h8)
	) name11512 (
		\wishbone_bd_ram_mem2_reg[241][23]/P0001 ,
		_w13006_,
		_w22024_
	);
	LUT2 #(
		.INIT('h8)
	) name11513 (
		\wishbone_bd_ram_mem2_reg[227][23]/P0001 ,
		_w12936_,
		_w22025_
	);
	LUT2 #(
		.INIT('h8)
	) name11514 (
		\wishbone_bd_ram_mem2_reg[9][23]/P0001 ,
		_w12808_,
		_w22026_
	);
	LUT2 #(
		.INIT('h8)
	) name11515 (
		\wishbone_bd_ram_mem2_reg[206][23]/P0001 ,
		_w12954_,
		_w22027_
	);
	LUT2 #(
		.INIT('h8)
	) name11516 (
		\wishbone_bd_ram_mem2_reg[78][23]/P0001 ,
		_w12874_,
		_w22028_
	);
	LUT2 #(
		.INIT('h8)
	) name11517 (
		\wishbone_bd_ram_mem2_reg[207][23]/P0001 ,
		_w13180_,
		_w22029_
	);
	LUT2 #(
		.INIT('h8)
	) name11518 (
		\wishbone_bd_ram_mem2_reg[117][23]/P0001 ,
		_w12715_,
		_w22030_
	);
	LUT2 #(
		.INIT('h8)
	) name11519 (
		\wishbone_bd_ram_mem2_reg[237][23]/P0001 ,
		_w12990_,
		_w22031_
	);
	LUT2 #(
		.INIT('h8)
	) name11520 (
		\wishbone_bd_ram_mem2_reg[143][23]/P0001 ,
		_w12922_,
		_w22032_
	);
	LUT2 #(
		.INIT('h8)
	) name11521 (
		\wishbone_bd_ram_mem2_reg[152][23]/P0001 ,
		_w12966_,
		_w22033_
	);
	LUT2 #(
		.INIT('h8)
	) name11522 (
		\wishbone_bd_ram_mem2_reg[25][23]/P0001 ,
		_w13108_,
		_w22034_
	);
	LUT2 #(
		.INIT('h8)
	) name11523 (
		\wishbone_bd_ram_mem2_reg[32][23]/P0001 ,
		_w13120_,
		_w22035_
	);
	LUT2 #(
		.INIT('h8)
	) name11524 (
		\wishbone_bd_ram_mem2_reg[120][23]/P0001 ,
		_w12707_,
		_w22036_
	);
	LUT2 #(
		.INIT('h8)
	) name11525 (
		\wishbone_bd_ram_mem2_reg[115][23]/P0001 ,
		_w13112_,
		_w22037_
	);
	LUT2 #(
		.INIT('h8)
	) name11526 (
		\wishbone_bd_ram_mem2_reg[84][23]/P0001 ,
		_w12934_,
		_w22038_
	);
	LUT2 #(
		.INIT('h8)
	) name11527 (
		\wishbone_bd_ram_mem2_reg[16][23]/P0001 ,
		_w13140_,
		_w22039_
	);
	LUT2 #(
		.INIT('h8)
	) name11528 (
		\wishbone_bd_ram_mem2_reg[33][23]/P0001 ,
		_w12980_,
		_w22040_
	);
	LUT2 #(
		.INIT('h8)
	) name11529 (
		\wishbone_bd_ram_mem2_reg[131][23]/P0001 ,
		_w12852_,
		_w22041_
	);
	LUT2 #(
		.INIT('h8)
	) name11530 (
		\wishbone_bd_ram_mem2_reg[248][23]/P0001 ,
		_w12789_,
		_w22042_
	);
	LUT2 #(
		.INIT('h8)
	) name11531 (
		\wishbone_bd_ram_mem2_reg[15][23]/P0001 ,
		_w13210_,
		_w22043_
	);
	LUT2 #(
		.INIT('h8)
	) name11532 (
		\wishbone_bd_ram_mem2_reg[247][23]/P0001 ,
		_w12818_,
		_w22044_
	);
	LUT2 #(
		.INIT('h8)
	) name11533 (
		\wishbone_bd_ram_mem2_reg[154][23]/P0001 ,
		_w12962_,
		_w22045_
	);
	LUT2 #(
		.INIT('h8)
	) name11534 (
		\wishbone_bd_ram_mem2_reg[93][23]/P0001 ,
		_w13016_,
		_w22046_
	);
	LUT2 #(
		.INIT('h8)
	) name11535 (
		\wishbone_bd_ram_mem2_reg[39][23]/P0001 ,
		_w13018_,
		_w22047_
	);
	LUT2 #(
		.INIT('h8)
	) name11536 (
		\wishbone_bd_ram_mem2_reg[57][23]/P0001 ,
		_w13116_,
		_w22048_
	);
	LUT2 #(
		.INIT('h8)
	) name11537 (
		\wishbone_bd_ram_mem2_reg[28][23]/P0001 ,
		_w13170_,
		_w22049_
	);
	LUT2 #(
		.INIT('h8)
	) name11538 (
		\wishbone_bd_ram_mem2_reg[148][23]/P0001 ,
		_w13000_,
		_w22050_
	);
	LUT2 #(
		.INIT('h8)
	) name11539 (
		\wishbone_bd_ram_mem2_reg[190][23]/P0001 ,
		_w12858_,
		_w22051_
	);
	LUT2 #(
		.INIT('h8)
	) name11540 (
		\wishbone_bd_ram_mem2_reg[0][23]/P0001 ,
		_w12717_,
		_w22052_
	);
	LUT2 #(
		.INIT('h8)
	) name11541 (
		\wishbone_bd_ram_mem2_reg[122][23]/P0001 ,
		_w13130_,
		_w22053_
	);
	LUT2 #(
		.INIT('h8)
	) name11542 (
		\wishbone_bd_ram_mem2_reg[46][23]/P0001 ,
		_w12884_,
		_w22054_
	);
	LUT2 #(
		.INIT('h8)
	) name11543 (
		\wishbone_bd_ram_mem2_reg[155][23]/P0001 ,
		_w13122_,
		_w22055_
	);
	LUT2 #(
		.INIT('h8)
	) name11544 (
		\wishbone_bd_ram_mem2_reg[132][23]/P0001 ,
		_w12992_,
		_w22056_
	);
	LUT2 #(
		.INIT('h8)
	) name11545 (
		\wishbone_bd_ram_mem2_reg[17][23]/P0001 ,
		_w12848_,
		_w22057_
	);
	LUT2 #(
		.INIT('h8)
	) name11546 (
		\wishbone_bd_ram_mem2_reg[208][23]/P0001 ,
		_w13032_,
		_w22058_
	);
	LUT2 #(
		.INIT('h8)
	) name11547 (
		\wishbone_bd_ram_mem2_reg[49][23]/P0001 ,
		_w12994_,
		_w22059_
	);
	LUT2 #(
		.INIT('h8)
	) name11548 (
		\wishbone_bd_ram_mem2_reg[63][23]/P0001 ,
		_w12850_,
		_w22060_
	);
	LUT2 #(
		.INIT('h8)
	) name11549 (
		\wishbone_bd_ram_mem2_reg[253][23]/P0001 ,
		_w13100_,
		_w22061_
	);
	LUT2 #(
		.INIT('h8)
	) name11550 (
		\wishbone_bd_ram_mem2_reg[36][23]/P0001 ,
		_w12800_,
		_w22062_
	);
	LUT2 #(
		.INIT('h8)
	) name11551 (
		\wishbone_bd_ram_mem2_reg[113][23]/P0001 ,
		_w13026_,
		_w22063_
	);
	LUT2 #(
		.INIT('h8)
	) name11552 (
		\wishbone_bd_ram_mem2_reg[187][23]/P0001 ,
		_w13196_,
		_w22064_
	);
	LUT2 #(
		.INIT('h8)
	) name11553 (
		\wishbone_bd_ram_mem2_reg[185][23]/P0001 ,
		_w12940_,
		_w22065_
	);
	LUT2 #(
		.INIT('h8)
	) name11554 (
		\wishbone_bd_ram_mem2_reg[167][23]/P0001 ,
		_w12986_,
		_w22066_
	);
	LUT2 #(
		.INIT('h8)
	) name11555 (
		\wishbone_bd_ram_mem2_reg[130][23]/P0001 ,
		_w12914_,
		_w22067_
	);
	LUT2 #(
		.INIT('h8)
	) name11556 (
		\wishbone_bd_ram_mem2_reg[52][23]/P0001 ,
		_w13082_,
		_w22068_
	);
	LUT2 #(
		.INIT('h8)
	) name11557 (
		\wishbone_bd_ram_mem2_reg[137][23]/P0001 ,
		_w13168_,
		_w22069_
	);
	LUT2 #(
		.INIT('h8)
	) name11558 (
		\wishbone_bd_ram_mem2_reg[108][23]/P0001 ,
		_w13156_,
		_w22070_
	);
	LUT2 #(
		.INIT('h8)
	) name11559 (
		\wishbone_bd_ram_mem2_reg[60][23]/P0001 ,
		_w13204_,
		_w22071_
	);
	LUT2 #(
		.INIT('h8)
	) name11560 (
		\wishbone_bd_ram_mem2_reg[45][23]/P0001 ,
		_w12908_,
		_w22072_
	);
	LUT2 #(
		.INIT('h8)
	) name11561 (
		\wishbone_bd_ram_mem2_reg[110][23]/P0001 ,
		_w13046_,
		_w22073_
	);
	LUT2 #(
		.INIT('h8)
	) name11562 (
		\wishbone_bd_ram_mem2_reg[183][23]/P0001 ,
		_w12787_,
		_w22074_
	);
	LUT2 #(
		.INIT('h8)
	) name11563 (
		\wishbone_bd_ram_mem2_reg[171][23]/P0001 ,
		_w12910_,
		_w22075_
	);
	LUT2 #(
		.INIT('h8)
	) name11564 (
		\wishbone_bd_ram_mem2_reg[41][23]/P0001 ,
		_w13052_,
		_w22076_
	);
	LUT2 #(
		.INIT('h8)
	) name11565 (
		\wishbone_bd_ram_mem2_reg[226][23]/P0001 ,
		_w13138_,
		_w22077_
	);
	LUT2 #(
		.INIT('h8)
	) name11566 (
		\wishbone_bd_ram_mem2_reg[165][23]/P0001 ,
		_w13044_,
		_w22078_
	);
	LUT2 #(
		.INIT('h8)
	) name11567 (
		\wishbone_bd_ram_mem2_reg[124][23]/P0001 ,
		_w13058_,
		_w22079_
	);
	LUT2 #(
		.INIT('h8)
	) name11568 (
		\wishbone_bd_ram_mem2_reg[128][23]/P0001 ,
		_w12793_,
		_w22080_
	);
	LUT2 #(
		.INIT('h8)
	) name11569 (
		\wishbone_bd_ram_mem2_reg[184][23]/P0001 ,
		_w13062_,
		_w22081_
	);
	LUT2 #(
		.INIT('h8)
	) name11570 (
		\wishbone_bd_ram_mem2_reg[19][23]/P0001 ,
		_w13012_,
		_w22082_
	);
	LUT2 #(
		.INIT('h8)
	) name11571 (
		\wishbone_bd_ram_mem2_reg[244][23]/P0001 ,
		_w12747_,
		_w22083_
	);
	LUT2 #(
		.INIT('h8)
	) name11572 (
		\wishbone_bd_ram_mem2_reg[170][23]/P0001 ,
		_w13030_,
		_w22084_
	);
	LUT2 #(
		.INIT('h8)
	) name11573 (
		\wishbone_bd_ram_mem2_reg[44][23]/P0001 ,
		_w12896_,
		_w22085_
	);
	LUT2 #(
		.INIT('h8)
	) name11574 (
		\wishbone_bd_ram_mem2_reg[90][23]/P0001 ,
		_w12978_,
		_w22086_
	);
	LUT2 #(
		.INIT('h8)
	) name11575 (
		\wishbone_bd_ram_mem2_reg[198][23]/P0001 ,
		_w12832_,
		_w22087_
	);
	LUT2 #(
		.INIT('h8)
	) name11576 (
		\wishbone_bd_ram_mem2_reg[216][23]/P0001 ,
		_w13028_,
		_w22088_
	);
	LUT2 #(
		.INIT('h8)
	) name11577 (
		\wishbone_bd_ram_mem2_reg[86][23]/P0001 ,
		_w12735_,
		_w22089_
	);
	LUT2 #(
		.INIT('h8)
	) name11578 (
		\wishbone_bd_ram_mem2_reg[215][23]/P0001 ,
		_w12974_,
		_w22090_
	);
	LUT2 #(
		.INIT('h8)
	) name11579 (
		\wishbone_bd_ram_mem2_reg[145][23]/P0001 ,
		_w13106_,
		_w22091_
	);
	LUT2 #(
		.INIT('h8)
	) name11580 (
		\wishbone_bd_ram_mem2_reg[96][23]/P0001 ,
		_w12912_,
		_w22092_
	);
	LUT2 #(
		.INIT('h8)
	) name11581 (
		\wishbone_bd_ram_mem2_reg[14][23]/P0001 ,
		_w13086_,
		_w22093_
	);
	LUT2 #(
		.INIT('h8)
	) name11582 (
		\wishbone_bd_ram_mem2_reg[89][23]/P0001 ,
		_w12964_,
		_w22094_
	);
	LUT2 #(
		.INIT('h8)
	) name11583 (
		\wishbone_bd_ram_mem2_reg[100][23]/P0001 ,
		_w12960_,
		_w22095_
	);
	LUT2 #(
		.INIT('h8)
	) name11584 (
		\wishbone_bd_ram_mem2_reg[94][23]/P0001 ,
		_w13186_,
		_w22096_
	);
	LUT2 #(
		.INIT('h8)
	) name11585 (
		\wishbone_bd_ram_mem2_reg[176][23]/P0001 ,
		_w12868_,
		_w22097_
	);
	LUT2 #(
		.INIT('h8)
	) name11586 (
		\wishbone_bd_ram_mem2_reg[172][23]/P0001 ,
		_w12944_,
		_w22098_
	);
	LUT2 #(
		.INIT('h8)
	) name11587 (
		\wishbone_bd_ram_mem2_reg[193][23]/P0001 ,
		_w13056_,
		_w22099_
	);
	LUT2 #(
		.INIT('h8)
	) name11588 (
		\wishbone_bd_ram_mem2_reg[233][23]/P0001 ,
		_w12836_,
		_w22100_
	);
	LUT2 #(
		.INIT('h8)
	) name11589 (
		\wishbone_bd_ram_mem2_reg[37][23]/P0001 ,
		_w13102_,
		_w22101_
	);
	LUT2 #(
		.INIT('h8)
	) name11590 (
		\wishbone_bd_ram_mem2_reg[177][23]/P0001 ,
		_w12996_,
		_w22102_
	);
	LUT2 #(
		.INIT('h8)
	) name11591 (
		\wishbone_bd_ram_mem2_reg[174][23]/P0001 ,
		_w12972_,
		_w22103_
	);
	LUT2 #(
		.INIT('h8)
	) name11592 (
		\wishbone_bd_ram_mem2_reg[99][23]/P0001 ,
		_w13038_,
		_w22104_
	);
	LUT2 #(
		.INIT('h8)
	) name11593 (
		\wishbone_bd_ram_mem2_reg[186][23]/P0001 ,
		_w12783_,
		_w22105_
	);
	LUT2 #(
		.INIT('h8)
	) name11594 (
		\wishbone_bd_ram_mem2_reg[195][23]/P0001 ,
		_w13144_,
		_w22106_
	);
	LUT2 #(
		.INIT('h8)
	) name11595 (
		\wishbone_bd_ram_mem2_reg[76][23]/P0001 ,
		_w13184_,
		_w22107_
	);
	LUT2 #(
		.INIT('h8)
	) name11596 (
		\wishbone_bd_ram_mem2_reg[67][23]/P0001 ,
		_w13134_,
		_w22108_
	);
	LUT2 #(
		.INIT('h8)
	) name11597 (
		\wishbone_bd_ram_mem2_reg[121][23]/P0001 ,
		_w13078_,
		_w22109_
	);
	LUT2 #(
		.INIT('h8)
	) name11598 (
		\wishbone_bd_ram_mem2_reg[48][23]/P0001 ,
		_w12970_,
		_w22110_
	);
	LUT2 #(
		.INIT('h8)
	) name11599 (
		\wishbone_bd_ram_mem2_reg[169][23]/P0001 ,
		_w12722_,
		_w22111_
	);
	LUT2 #(
		.INIT('h8)
	) name11600 (
		\wishbone_bd_ram_mem2_reg[12][23]/P0001 ,
		_w13118_,
		_w22112_
	);
	LUT2 #(
		.INIT('h8)
	) name11601 (
		\wishbone_bd_ram_mem2_reg[30][23]/P0001 ,
		_w13104_,
		_w22113_
	);
	LUT2 #(
		.INIT('h8)
	) name11602 (
		\wishbone_bd_ram_mem2_reg[221][23]/P0001 ,
		_w12802_,
		_w22114_
	);
	LUT2 #(
		.INIT('h8)
	) name11603 (
		\wishbone_bd_ram_mem2_reg[188][23]/P0001 ,
		_w12948_,
		_w22115_
	);
	LUT2 #(
		.INIT('h8)
	) name11604 (
		\wishbone_bd_ram_mem2_reg[2][23]/P0001 ,
		_w13088_,
		_w22116_
	);
	LUT2 #(
		.INIT('h8)
	) name11605 (
		\wishbone_bd_ram_mem2_reg[42][23]/P0001 ,
		_w12842_,
		_w22117_
	);
	LUT2 #(
		.INIT('h8)
	) name11606 (
		\wishbone_bd_ram_mem2_reg[218][23]/P0001 ,
		_w13206_,
		_w22118_
	);
	LUT2 #(
		.INIT('h8)
	) name11607 (
		\wishbone_bd_ram_mem2_reg[158][23]/P0001 ,
		_w12898_,
		_w22119_
	);
	LUT2 #(
		.INIT('h8)
	) name11608 (
		\wishbone_bd_ram_mem2_reg[40][23]/P0001 ,
		_w13132_,
		_w22120_
	);
	LUT2 #(
		.INIT('h8)
	) name11609 (
		\wishbone_bd_ram_mem2_reg[21][23]/P0001 ,
		_w12906_,
		_w22121_
	);
	LUT2 #(
		.INIT('h8)
	) name11610 (
		\wishbone_bd_ram_mem2_reg[101][23]/P0001 ,
		_w13192_,
		_w22122_
	);
	LUT2 #(
		.INIT('h8)
	) name11611 (
		\wishbone_bd_ram_mem2_reg[147][23]/P0001 ,
		_w13146_,
		_w22123_
	);
	LUT2 #(
		.INIT('h8)
	) name11612 (
		\wishbone_bd_ram_mem2_reg[98][23]/P0001 ,
		_w12816_,
		_w22124_
	);
	LUT2 #(
		.INIT('h8)
	) name11613 (
		\wishbone_bd_ram_mem2_reg[27][23]/P0001 ,
		_w12880_,
		_w22125_
	);
	LUT2 #(
		.INIT('h8)
	) name11614 (
		\wishbone_bd_ram_mem2_reg[205][23]/P0001 ,
		_w13068_,
		_w22126_
	);
	LUT2 #(
		.INIT('h8)
	) name11615 (
		\wishbone_bd_ram_mem2_reg[71][23]/P0001 ,
		_w12798_,
		_w22127_
	);
	LUT2 #(
		.INIT('h8)
	) name11616 (
		\wishbone_bd_ram_mem2_reg[58][23]/P0001 ,
		_w13070_,
		_w22128_
	);
	LUT2 #(
		.INIT('h8)
	) name11617 (
		\wishbone_bd_ram_mem2_reg[200][23]/P0001 ,
		_w12988_,
		_w22129_
	);
	LUT2 #(
		.INIT('h8)
	) name11618 (
		\wishbone_bd_ram_mem2_reg[254][23]/P0001 ,
		_w12892_,
		_w22130_
	);
	LUT2 #(
		.INIT('h8)
	) name11619 (
		\wishbone_bd_ram_mem2_reg[204][23]/P0001 ,
		_w13162_,
		_w22131_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		\wishbone_bd_ram_mem2_reg[127][23]/P0001 ,
		_w13164_,
		_w22132_
	);
	LUT2 #(
		.INIT('h8)
	) name11621 (
		\wishbone_bd_ram_mem2_reg[224][23]/P0001 ,
		_w12902_,
		_w22133_
	);
	LUT2 #(
		.INIT('h8)
	) name11622 (
		\wishbone_bd_ram_mem2_reg[229][23]/P0001 ,
		_w12711_,
		_w22134_
	);
	LUT2 #(
		.INIT('h8)
	) name11623 (
		\wishbone_bd_ram_mem2_reg[225][23]/P0001 ,
		_w13092_,
		_w22135_
	);
	LUT2 #(
		.INIT('h8)
	) name11624 (
		\wishbone_bd_ram_mem2_reg[83][23]/P0001 ,
		_w12916_,
		_w22136_
	);
	LUT2 #(
		.INIT('h8)
	) name11625 (
		\wishbone_bd_ram_mem2_reg[69][23]/P0001 ,
		_w12738_,
		_w22137_
	);
	LUT2 #(
		.INIT('h8)
	) name11626 (
		\wishbone_bd_ram_mem2_reg[119][23]/P0001 ,
		_w13048_,
		_w22138_
	);
	LUT2 #(
		.INIT('h8)
	) name11627 (
		\wishbone_bd_ram_mem2_reg[146][23]/P0001 ,
		_w13060_,
		_w22139_
	);
	LUT2 #(
		.INIT('h8)
	) name11628 (
		\wishbone_bd_ram_mem2_reg[252][23]/P0001 ,
		_w13080_,
		_w22140_
	);
	LUT2 #(
		.INIT('h8)
	) name11629 (
		\wishbone_bd_ram_mem2_reg[77][23]/P0001 ,
		_w12982_,
		_w22141_
	);
	LUT2 #(
		.INIT('h8)
	) name11630 (
		\wishbone_bd_ram_mem2_reg[116][23]/P0001 ,
		_w12998_,
		_w22142_
	);
	LUT2 #(
		.INIT('h8)
	) name11631 (
		\wishbone_bd_ram_mem2_reg[23][23]/P0001 ,
		_w13008_,
		_w22143_
	);
	LUT2 #(
		.INIT('h8)
	) name11632 (
		\wishbone_bd_ram_mem2_reg[246][23]/P0001 ,
		_w13076_,
		_w22144_
	);
	LUT2 #(
		.INIT('h8)
	) name11633 (
		\wishbone_bd_ram_mem2_reg[156][23]/P0001 ,
		_w13190_,
		_w22145_
	);
	LUT2 #(
		.INIT('h8)
	) name11634 (
		\wishbone_bd_ram_mem2_reg[74][23]/P0001 ,
		_w12812_,
		_w22146_
	);
	LUT2 #(
		.INIT('h8)
	) name11635 (
		\wishbone_bd_ram_mem2_reg[91][23]/P0001 ,
		_w13074_,
		_w22147_
	);
	LUT2 #(
		.INIT('h8)
	) name11636 (
		\wishbone_bd_ram_mem2_reg[217][23]/P0001 ,
		_w13188_,
		_w22148_
	);
	LUT2 #(
		.INIT('h8)
	) name11637 (
		\wishbone_bd_ram_mem2_reg[162][23]/P0001 ,
		_w13098_,
		_w22149_
	);
	LUT2 #(
		.INIT('h8)
	) name11638 (
		\wishbone_bd_ram_mem2_reg[4][23]/P0001 ,
		_w12666_,
		_w22150_
	);
	LUT2 #(
		.INIT('h8)
	) name11639 (
		\wishbone_bd_ram_mem2_reg[106][23]/P0001 ,
		_w12713_,
		_w22151_
	);
	LUT2 #(
		.INIT('h8)
	) name11640 (
		\wishbone_bd_ram_mem2_reg[26][23]/P0001 ,
		_w12699_,
		_w22152_
	);
	LUT2 #(
		.INIT('h8)
	) name11641 (
		\wishbone_bd_ram_mem2_reg[150][23]/P0001 ,
		_w13136_,
		_w22153_
	);
	LUT2 #(
		.INIT('h8)
	) name11642 (
		\wishbone_bd_ram_mem2_reg[22][23]/P0001 ,
		_w13110_,
		_w22154_
	);
	LUT2 #(
		.INIT('h8)
	) name11643 (
		\wishbone_bd_ram_mem2_reg[168][23]/P0001 ,
		_w13208_,
		_w22155_
	);
	LUT2 #(
		.INIT('h8)
	) name11644 (
		\wishbone_bd_ram_mem2_reg[95][23]/P0001 ,
		_w12844_,
		_w22156_
	);
	LUT2 #(
		.INIT('h8)
	) name11645 (
		\wishbone_bd_ram_mem2_reg[232][23]/P0001 ,
		_w12758_,
		_w22157_
	);
	LUT2 #(
		.INIT('h8)
	) name11646 (
		\wishbone_bd_ram_mem2_reg[13][23]/P0001 ,
		_w13178_,
		_w22158_
	);
	LUT2 #(
		.INIT('h8)
	) name11647 (
		\wishbone_bd_ram_mem2_reg[173][23]/P0001 ,
		_w12854_,
		_w22159_
	);
	LUT2 #(
		.INIT('h1)
	) name11648 (
		_w21904_,
		_w21905_,
		_w22160_
	);
	LUT2 #(
		.INIT('h1)
	) name11649 (
		_w21906_,
		_w21907_,
		_w22161_
	);
	LUT2 #(
		.INIT('h1)
	) name11650 (
		_w21908_,
		_w21909_,
		_w22162_
	);
	LUT2 #(
		.INIT('h1)
	) name11651 (
		_w21910_,
		_w21911_,
		_w22163_
	);
	LUT2 #(
		.INIT('h1)
	) name11652 (
		_w21912_,
		_w21913_,
		_w22164_
	);
	LUT2 #(
		.INIT('h1)
	) name11653 (
		_w21914_,
		_w21915_,
		_w22165_
	);
	LUT2 #(
		.INIT('h1)
	) name11654 (
		_w21916_,
		_w21917_,
		_w22166_
	);
	LUT2 #(
		.INIT('h1)
	) name11655 (
		_w21918_,
		_w21919_,
		_w22167_
	);
	LUT2 #(
		.INIT('h1)
	) name11656 (
		_w21920_,
		_w21921_,
		_w22168_
	);
	LUT2 #(
		.INIT('h1)
	) name11657 (
		_w21922_,
		_w21923_,
		_w22169_
	);
	LUT2 #(
		.INIT('h1)
	) name11658 (
		_w21924_,
		_w21925_,
		_w22170_
	);
	LUT2 #(
		.INIT('h1)
	) name11659 (
		_w21926_,
		_w21927_,
		_w22171_
	);
	LUT2 #(
		.INIT('h1)
	) name11660 (
		_w21928_,
		_w21929_,
		_w22172_
	);
	LUT2 #(
		.INIT('h1)
	) name11661 (
		_w21930_,
		_w21931_,
		_w22173_
	);
	LUT2 #(
		.INIT('h1)
	) name11662 (
		_w21932_,
		_w21933_,
		_w22174_
	);
	LUT2 #(
		.INIT('h1)
	) name11663 (
		_w21934_,
		_w21935_,
		_w22175_
	);
	LUT2 #(
		.INIT('h1)
	) name11664 (
		_w21936_,
		_w21937_,
		_w22176_
	);
	LUT2 #(
		.INIT('h1)
	) name11665 (
		_w21938_,
		_w21939_,
		_w22177_
	);
	LUT2 #(
		.INIT('h1)
	) name11666 (
		_w21940_,
		_w21941_,
		_w22178_
	);
	LUT2 #(
		.INIT('h1)
	) name11667 (
		_w21942_,
		_w21943_,
		_w22179_
	);
	LUT2 #(
		.INIT('h1)
	) name11668 (
		_w21944_,
		_w21945_,
		_w22180_
	);
	LUT2 #(
		.INIT('h1)
	) name11669 (
		_w21946_,
		_w21947_,
		_w22181_
	);
	LUT2 #(
		.INIT('h1)
	) name11670 (
		_w21948_,
		_w21949_,
		_w22182_
	);
	LUT2 #(
		.INIT('h1)
	) name11671 (
		_w21950_,
		_w21951_,
		_w22183_
	);
	LUT2 #(
		.INIT('h1)
	) name11672 (
		_w21952_,
		_w21953_,
		_w22184_
	);
	LUT2 #(
		.INIT('h1)
	) name11673 (
		_w21954_,
		_w21955_,
		_w22185_
	);
	LUT2 #(
		.INIT('h1)
	) name11674 (
		_w21956_,
		_w21957_,
		_w22186_
	);
	LUT2 #(
		.INIT('h1)
	) name11675 (
		_w21958_,
		_w21959_,
		_w22187_
	);
	LUT2 #(
		.INIT('h1)
	) name11676 (
		_w21960_,
		_w21961_,
		_w22188_
	);
	LUT2 #(
		.INIT('h1)
	) name11677 (
		_w21962_,
		_w21963_,
		_w22189_
	);
	LUT2 #(
		.INIT('h1)
	) name11678 (
		_w21964_,
		_w21965_,
		_w22190_
	);
	LUT2 #(
		.INIT('h1)
	) name11679 (
		_w21966_,
		_w21967_,
		_w22191_
	);
	LUT2 #(
		.INIT('h1)
	) name11680 (
		_w21968_,
		_w21969_,
		_w22192_
	);
	LUT2 #(
		.INIT('h1)
	) name11681 (
		_w21970_,
		_w21971_,
		_w22193_
	);
	LUT2 #(
		.INIT('h1)
	) name11682 (
		_w21972_,
		_w21973_,
		_w22194_
	);
	LUT2 #(
		.INIT('h1)
	) name11683 (
		_w21974_,
		_w21975_,
		_w22195_
	);
	LUT2 #(
		.INIT('h1)
	) name11684 (
		_w21976_,
		_w21977_,
		_w22196_
	);
	LUT2 #(
		.INIT('h1)
	) name11685 (
		_w21978_,
		_w21979_,
		_w22197_
	);
	LUT2 #(
		.INIT('h1)
	) name11686 (
		_w21980_,
		_w21981_,
		_w22198_
	);
	LUT2 #(
		.INIT('h1)
	) name11687 (
		_w21982_,
		_w21983_,
		_w22199_
	);
	LUT2 #(
		.INIT('h1)
	) name11688 (
		_w21984_,
		_w21985_,
		_w22200_
	);
	LUT2 #(
		.INIT('h1)
	) name11689 (
		_w21986_,
		_w21987_,
		_w22201_
	);
	LUT2 #(
		.INIT('h1)
	) name11690 (
		_w21988_,
		_w21989_,
		_w22202_
	);
	LUT2 #(
		.INIT('h1)
	) name11691 (
		_w21990_,
		_w21991_,
		_w22203_
	);
	LUT2 #(
		.INIT('h1)
	) name11692 (
		_w21992_,
		_w21993_,
		_w22204_
	);
	LUT2 #(
		.INIT('h1)
	) name11693 (
		_w21994_,
		_w21995_,
		_w22205_
	);
	LUT2 #(
		.INIT('h1)
	) name11694 (
		_w21996_,
		_w21997_,
		_w22206_
	);
	LUT2 #(
		.INIT('h1)
	) name11695 (
		_w21998_,
		_w21999_,
		_w22207_
	);
	LUT2 #(
		.INIT('h1)
	) name11696 (
		_w22000_,
		_w22001_,
		_w22208_
	);
	LUT2 #(
		.INIT('h1)
	) name11697 (
		_w22002_,
		_w22003_,
		_w22209_
	);
	LUT2 #(
		.INIT('h1)
	) name11698 (
		_w22004_,
		_w22005_,
		_w22210_
	);
	LUT2 #(
		.INIT('h1)
	) name11699 (
		_w22006_,
		_w22007_,
		_w22211_
	);
	LUT2 #(
		.INIT('h1)
	) name11700 (
		_w22008_,
		_w22009_,
		_w22212_
	);
	LUT2 #(
		.INIT('h1)
	) name11701 (
		_w22010_,
		_w22011_,
		_w22213_
	);
	LUT2 #(
		.INIT('h1)
	) name11702 (
		_w22012_,
		_w22013_,
		_w22214_
	);
	LUT2 #(
		.INIT('h1)
	) name11703 (
		_w22014_,
		_w22015_,
		_w22215_
	);
	LUT2 #(
		.INIT('h1)
	) name11704 (
		_w22016_,
		_w22017_,
		_w22216_
	);
	LUT2 #(
		.INIT('h1)
	) name11705 (
		_w22018_,
		_w22019_,
		_w22217_
	);
	LUT2 #(
		.INIT('h1)
	) name11706 (
		_w22020_,
		_w22021_,
		_w22218_
	);
	LUT2 #(
		.INIT('h1)
	) name11707 (
		_w22022_,
		_w22023_,
		_w22219_
	);
	LUT2 #(
		.INIT('h1)
	) name11708 (
		_w22024_,
		_w22025_,
		_w22220_
	);
	LUT2 #(
		.INIT('h1)
	) name11709 (
		_w22026_,
		_w22027_,
		_w22221_
	);
	LUT2 #(
		.INIT('h1)
	) name11710 (
		_w22028_,
		_w22029_,
		_w22222_
	);
	LUT2 #(
		.INIT('h1)
	) name11711 (
		_w22030_,
		_w22031_,
		_w22223_
	);
	LUT2 #(
		.INIT('h1)
	) name11712 (
		_w22032_,
		_w22033_,
		_w22224_
	);
	LUT2 #(
		.INIT('h1)
	) name11713 (
		_w22034_,
		_w22035_,
		_w22225_
	);
	LUT2 #(
		.INIT('h1)
	) name11714 (
		_w22036_,
		_w22037_,
		_w22226_
	);
	LUT2 #(
		.INIT('h1)
	) name11715 (
		_w22038_,
		_w22039_,
		_w22227_
	);
	LUT2 #(
		.INIT('h1)
	) name11716 (
		_w22040_,
		_w22041_,
		_w22228_
	);
	LUT2 #(
		.INIT('h1)
	) name11717 (
		_w22042_,
		_w22043_,
		_w22229_
	);
	LUT2 #(
		.INIT('h1)
	) name11718 (
		_w22044_,
		_w22045_,
		_w22230_
	);
	LUT2 #(
		.INIT('h1)
	) name11719 (
		_w22046_,
		_w22047_,
		_w22231_
	);
	LUT2 #(
		.INIT('h1)
	) name11720 (
		_w22048_,
		_w22049_,
		_w22232_
	);
	LUT2 #(
		.INIT('h1)
	) name11721 (
		_w22050_,
		_w22051_,
		_w22233_
	);
	LUT2 #(
		.INIT('h1)
	) name11722 (
		_w22052_,
		_w22053_,
		_w22234_
	);
	LUT2 #(
		.INIT('h1)
	) name11723 (
		_w22054_,
		_w22055_,
		_w22235_
	);
	LUT2 #(
		.INIT('h1)
	) name11724 (
		_w22056_,
		_w22057_,
		_w22236_
	);
	LUT2 #(
		.INIT('h1)
	) name11725 (
		_w22058_,
		_w22059_,
		_w22237_
	);
	LUT2 #(
		.INIT('h1)
	) name11726 (
		_w22060_,
		_w22061_,
		_w22238_
	);
	LUT2 #(
		.INIT('h1)
	) name11727 (
		_w22062_,
		_w22063_,
		_w22239_
	);
	LUT2 #(
		.INIT('h1)
	) name11728 (
		_w22064_,
		_w22065_,
		_w22240_
	);
	LUT2 #(
		.INIT('h1)
	) name11729 (
		_w22066_,
		_w22067_,
		_w22241_
	);
	LUT2 #(
		.INIT('h1)
	) name11730 (
		_w22068_,
		_w22069_,
		_w22242_
	);
	LUT2 #(
		.INIT('h1)
	) name11731 (
		_w22070_,
		_w22071_,
		_w22243_
	);
	LUT2 #(
		.INIT('h1)
	) name11732 (
		_w22072_,
		_w22073_,
		_w22244_
	);
	LUT2 #(
		.INIT('h1)
	) name11733 (
		_w22074_,
		_w22075_,
		_w22245_
	);
	LUT2 #(
		.INIT('h1)
	) name11734 (
		_w22076_,
		_w22077_,
		_w22246_
	);
	LUT2 #(
		.INIT('h1)
	) name11735 (
		_w22078_,
		_w22079_,
		_w22247_
	);
	LUT2 #(
		.INIT('h1)
	) name11736 (
		_w22080_,
		_w22081_,
		_w22248_
	);
	LUT2 #(
		.INIT('h1)
	) name11737 (
		_w22082_,
		_w22083_,
		_w22249_
	);
	LUT2 #(
		.INIT('h1)
	) name11738 (
		_w22084_,
		_w22085_,
		_w22250_
	);
	LUT2 #(
		.INIT('h1)
	) name11739 (
		_w22086_,
		_w22087_,
		_w22251_
	);
	LUT2 #(
		.INIT('h1)
	) name11740 (
		_w22088_,
		_w22089_,
		_w22252_
	);
	LUT2 #(
		.INIT('h1)
	) name11741 (
		_w22090_,
		_w22091_,
		_w22253_
	);
	LUT2 #(
		.INIT('h1)
	) name11742 (
		_w22092_,
		_w22093_,
		_w22254_
	);
	LUT2 #(
		.INIT('h1)
	) name11743 (
		_w22094_,
		_w22095_,
		_w22255_
	);
	LUT2 #(
		.INIT('h1)
	) name11744 (
		_w22096_,
		_w22097_,
		_w22256_
	);
	LUT2 #(
		.INIT('h1)
	) name11745 (
		_w22098_,
		_w22099_,
		_w22257_
	);
	LUT2 #(
		.INIT('h1)
	) name11746 (
		_w22100_,
		_w22101_,
		_w22258_
	);
	LUT2 #(
		.INIT('h1)
	) name11747 (
		_w22102_,
		_w22103_,
		_w22259_
	);
	LUT2 #(
		.INIT('h1)
	) name11748 (
		_w22104_,
		_w22105_,
		_w22260_
	);
	LUT2 #(
		.INIT('h1)
	) name11749 (
		_w22106_,
		_w22107_,
		_w22261_
	);
	LUT2 #(
		.INIT('h1)
	) name11750 (
		_w22108_,
		_w22109_,
		_w22262_
	);
	LUT2 #(
		.INIT('h1)
	) name11751 (
		_w22110_,
		_w22111_,
		_w22263_
	);
	LUT2 #(
		.INIT('h1)
	) name11752 (
		_w22112_,
		_w22113_,
		_w22264_
	);
	LUT2 #(
		.INIT('h1)
	) name11753 (
		_w22114_,
		_w22115_,
		_w22265_
	);
	LUT2 #(
		.INIT('h1)
	) name11754 (
		_w22116_,
		_w22117_,
		_w22266_
	);
	LUT2 #(
		.INIT('h1)
	) name11755 (
		_w22118_,
		_w22119_,
		_w22267_
	);
	LUT2 #(
		.INIT('h1)
	) name11756 (
		_w22120_,
		_w22121_,
		_w22268_
	);
	LUT2 #(
		.INIT('h1)
	) name11757 (
		_w22122_,
		_w22123_,
		_w22269_
	);
	LUT2 #(
		.INIT('h1)
	) name11758 (
		_w22124_,
		_w22125_,
		_w22270_
	);
	LUT2 #(
		.INIT('h1)
	) name11759 (
		_w22126_,
		_w22127_,
		_w22271_
	);
	LUT2 #(
		.INIT('h1)
	) name11760 (
		_w22128_,
		_w22129_,
		_w22272_
	);
	LUT2 #(
		.INIT('h1)
	) name11761 (
		_w22130_,
		_w22131_,
		_w22273_
	);
	LUT2 #(
		.INIT('h1)
	) name11762 (
		_w22132_,
		_w22133_,
		_w22274_
	);
	LUT2 #(
		.INIT('h1)
	) name11763 (
		_w22134_,
		_w22135_,
		_w22275_
	);
	LUT2 #(
		.INIT('h1)
	) name11764 (
		_w22136_,
		_w22137_,
		_w22276_
	);
	LUT2 #(
		.INIT('h1)
	) name11765 (
		_w22138_,
		_w22139_,
		_w22277_
	);
	LUT2 #(
		.INIT('h1)
	) name11766 (
		_w22140_,
		_w22141_,
		_w22278_
	);
	LUT2 #(
		.INIT('h1)
	) name11767 (
		_w22142_,
		_w22143_,
		_w22279_
	);
	LUT2 #(
		.INIT('h1)
	) name11768 (
		_w22144_,
		_w22145_,
		_w22280_
	);
	LUT2 #(
		.INIT('h1)
	) name11769 (
		_w22146_,
		_w22147_,
		_w22281_
	);
	LUT2 #(
		.INIT('h1)
	) name11770 (
		_w22148_,
		_w22149_,
		_w22282_
	);
	LUT2 #(
		.INIT('h1)
	) name11771 (
		_w22150_,
		_w22151_,
		_w22283_
	);
	LUT2 #(
		.INIT('h1)
	) name11772 (
		_w22152_,
		_w22153_,
		_w22284_
	);
	LUT2 #(
		.INIT('h1)
	) name11773 (
		_w22154_,
		_w22155_,
		_w22285_
	);
	LUT2 #(
		.INIT('h1)
	) name11774 (
		_w22156_,
		_w22157_,
		_w22286_
	);
	LUT2 #(
		.INIT('h1)
	) name11775 (
		_w22158_,
		_w22159_,
		_w22287_
	);
	LUT2 #(
		.INIT('h8)
	) name11776 (
		_w22286_,
		_w22287_,
		_w22288_
	);
	LUT2 #(
		.INIT('h8)
	) name11777 (
		_w22284_,
		_w22285_,
		_w22289_
	);
	LUT2 #(
		.INIT('h8)
	) name11778 (
		_w22282_,
		_w22283_,
		_w22290_
	);
	LUT2 #(
		.INIT('h8)
	) name11779 (
		_w22280_,
		_w22281_,
		_w22291_
	);
	LUT2 #(
		.INIT('h8)
	) name11780 (
		_w22278_,
		_w22279_,
		_w22292_
	);
	LUT2 #(
		.INIT('h8)
	) name11781 (
		_w22276_,
		_w22277_,
		_w22293_
	);
	LUT2 #(
		.INIT('h8)
	) name11782 (
		_w22274_,
		_w22275_,
		_w22294_
	);
	LUT2 #(
		.INIT('h8)
	) name11783 (
		_w22272_,
		_w22273_,
		_w22295_
	);
	LUT2 #(
		.INIT('h8)
	) name11784 (
		_w22270_,
		_w22271_,
		_w22296_
	);
	LUT2 #(
		.INIT('h8)
	) name11785 (
		_w22268_,
		_w22269_,
		_w22297_
	);
	LUT2 #(
		.INIT('h8)
	) name11786 (
		_w22266_,
		_w22267_,
		_w22298_
	);
	LUT2 #(
		.INIT('h8)
	) name11787 (
		_w22264_,
		_w22265_,
		_w22299_
	);
	LUT2 #(
		.INIT('h8)
	) name11788 (
		_w22262_,
		_w22263_,
		_w22300_
	);
	LUT2 #(
		.INIT('h8)
	) name11789 (
		_w22260_,
		_w22261_,
		_w22301_
	);
	LUT2 #(
		.INIT('h8)
	) name11790 (
		_w22258_,
		_w22259_,
		_w22302_
	);
	LUT2 #(
		.INIT('h8)
	) name11791 (
		_w22256_,
		_w22257_,
		_w22303_
	);
	LUT2 #(
		.INIT('h8)
	) name11792 (
		_w22254_,
		_w22255_,
		_w22304_
	);
	LUT2 #(
		.INIT('h8)
	) name11793 (
		_w22252_,
		_w22253_,
		_w22305_
	);
	LUT2 #(
		.INIT('h8)
	) name11794 (
		_w22250_,
		_w22251_,
		_w22306_
	);
	LUT2 #(
		.INIT('h8)
	) name11795 (
		_w22248_,
		_w22249_,
		_w22307_
	);
	LUT2 #(
		.INIT('h8)
	) name11796 (
		_w22246_,
		_w22247_,
		_w22308_
	);
	LUT2 #(
		.INIT('h8)
	) name11797 (
		_w22244_,
		_w22245_,
		_w22309_
	);
	LUT2 #(
		.INIT('h8)
	) name11798 (
		_w22242_,
		_w22243_,
		_w22310_
	);
	LUT2 #(
		.INIT('h8)
	) name11799 (
		_w22240_,
		_w22241_,
		_w22311_
	);
	LUT2 #(
		.INIT('h8)
	) name11800 (
		_w22238_,
		_w22239_,
		_w22312_
	);
	LUT2 #(
		.INIT('h8)
	) name11801 (
		_w22236_,
		_w22237_,
		_w22313_
	);
	LUT2 #(
		.INIT('h8)
	) name11802 (
		_w22234_,
		_w22235_,
		_w22314_
	);
	LUT2 #(
		.INIT('h8)
	) name11803 (
		_w22232_,
		_w22233_,
		_w22315_
	);
	LUT2 #(
		.INIT('h8)
	) name11804 (
		_w22230_,
		_w22231_,
		_w22316_
	);
	LUT2 #(
		.INIT('h8)
	) name11805 (
		_w22228_,
		_w22229_,
		_w22317_
	);
	LUT2 #(
		.INIT('h8)
	) name11806 (
		_w22226_,
		_w22227_,
		_w22318_
	);
	LUT2 #(
		.INIT('h8)
	) name11807 (
		_w22224_,
		_w22225_,
		_w22319_
	);
	LUT2 #(
		.INIT('h8)
	) name11808 (
		_w22222_,
		_w22223_,
		_w22320_
	);
	LUT2 #(
		.INIT('h8)
	) name11809 (
		_w22220_,
		_w22221_,
		_w22321_
	);
	LUT2 #(
		.INIT('h8)
	) name11810 (
		_w22218_,
		_w22219_,
		_w22322_
	);
	LUT2 #(
		.INIT('h8)
	) name11811 (
		_w22216_,
		_w22217_,
		_w22323_
	);
	LUT2 #(
		.INIT('h8)
	) name11812 (
		_w22214_,
		_w22215_,
		_w22324_
	);
	LUT2 #(
		.INIT('h8)
	) name11813 (
		_w22212_,
		_w22213_,
		_w22325_
	);
	LUT2 #(
		.INIT('h8)
	) name11814 (
		_w22210_,
		_w22211_,
		_w22326_
	);
	LUT2 #(
		.INIT('h8)
	) name11815 (
		_w22208_,
		_w22209_,
		_w22327_
	);
	LUT2 #(
		.INIT('h8)
	) name11816 (
		_w22206_,
		_w22207_,
		_w22328_
	);
	LUT2 #(
		.INIT('h8)
	) name11817 (
		_w22204_,
		_w22205_,
		_w22329_
	);
	LUT2 #(
		.INIT('h8)
	) name11818 (
		_w22202_,
		_w22203_,
		_w22330_
	);
	LUT2 #(
		.INIT('h8)
	) name11819 (
		_w22200_,
		_w22201_,
		_w22331_
	);
	LUT2 #(
		.INIT('h8)
	) name11820 (
		_w22198_,
		_w22199_,
		_w22332_
	);
	LUT2 #(
		.INIT('h8)
	) name11821 (
		_w22196_,
		_w22197_,
		_w22333_
	);
	LUT2 #(
		.INIT('h8)
	) name11822 (
		_w22194_,
		_w22195_,
		_w22334_
	);
	LUT2 #(
		.INIT('h8)
	) name11823 (
		_w22192_,
		_w22193_,
		_w22335_
	);
	LUT2 #(
		.INIT('h8)
	) name11824 (
		_w22190_,
		_w22191_,
		_w22336_
	);
	LUT2 #(
		.INIT('h8)
	) name11825 (
		_w22188_,
		_w22189_,
		_w22337_
	);
	LUT2 #(
		.INIT('h8)
	) name11826 (
		_w22186_,
		_w22187_,
		_w22338_
	);
	LUT2 #(
		.INIT('h8)
	) name11827 (
		_w22184_,
		_w22185_,
		_w22339_
	);
	LUT2 #(
		.INIT('h8)
	) name11828 (
		_w22182_,
		_w22183_,
		_w22340_
	);
	LUT2 #(
		.INIT('h8)
	) name11829 (
		_w22180_,
		_w22181_,
		_w22341_
	);
	LUT2 #(
		.INIT('h8)
	) name11830 (
		_w22178_,
		_w22179_,
		_w22342_
	);
	LUT2 #(
		.INIT('h8)
	) name11831 (
		_w22176_,
		_w22177_,
		_w22343_
	);
	LUT2 #(
		.INIT('h8)
	) name11832 (
		_w22174_,
		_w22175_,
		_w22344_
	);
	LUT2 #(
		.INIT('h8)
	) name11833 (
		_w22172_,
		_w22173_,
		_w22345_
	);
	LUT2 #(
		.INIT('h8)
	) name11834 (
		_w22170_,
		_w22171_,
		_w22346_
	);
	LUT2 #(
		.INIT('h8)
	) name11835 (
		_w22168_,
		_w22169_,
		_w22347_
	);
	LUT2 #(
		.INIT('h8)
	) name11836 (
		_w22166_,
		_w22167_,
		_w22348_
	);
	LUT2 #(
		.INIT('h8)
	) name11837 (
		_w22164_,
		_w22165_,
		_w22349_
	);
	LUT2 #(
		.INIT('h8)
	) name11838 (
		_w22162_,
		_w22163_,
		_w22350_
	);
	LUT2 #(
		.INIT('h8)
	) name11839 (
		_w22160_,
		_w22161_,
		_w22351_
	);
	LUT2 #(
		.INIT('h8)
	) name11840 (
		_w22350_,
		_w22351_,
		_w22352_
	);
	LUT2 #(
		.INIT('h8)
	) name11841 (
		_w22348_,
		_w22349_,
		_w22353_
	);
	LUT2 #(
		.INIT('h8)
	) name11842 (
		_w22346_,
		_w22347_,
		_w22354_
	);
	LUT2 #(
		.INIT('h8)
	) name11843 (
		_w22344_,
		_w22345_,
		_w22355_
	);
	LUT2 #(
		.INIT('h8)
	) name11844 (
		_w22342_,
		_w22343_,
		_w22356_
	);
	LUT2 #(
		.INIT('h8)
	) name11845 (
		_w22340_,
		_w22341_,
		_w22357_
	);
	LUT2 #(
		.INIT('h8)
	) name11846 (
		_w22338_,
		_w22339_,
		_w22358_
	);
	LUT2 #(
		.INIT('h8)
	) name11847 (
		_w22336_,
		_w22337_,
		_w22359_
	);
	LUT2 #(
		.INIT('h8)
	) name11848 (
		_w22334_,
		_w22335_,
		_w22360_
	);
	LUT2 #(
		.INIT('h8)
	) name11849 (
		_w22332_,
		_w22333_,
		_w22361_
	);
	LUT2 #(
		.INIT('h8)
	) name11850 (
		_w22330_,
		_w22331_,
		_w22362_
	);
	LUT2 #(
		.INIT('h8)
	) name11851 (
		_w22328_,
		_w22329_,
		_w22363_
	);
	LUT2 #(
		.INIT('h8)
	) name11852 (
		_w22326_,
		_w22327_,
		_w22364_
	);
	LUT2 #(
		.INIT('h8)
	) name11853 (
		_w22324_,
		_w22325_,
		_w22365_
	);
	LUT2 #(
		.INIT('h8)
	) name11854 (
		_w22322_,
		_w22323_,
		_w22366_
	);
	LUT2 #(
		.INIT('h8)
	) name11855 (
		_w22320_,
		_w22321_,
		_w22367_
	);
	LUT2 #(
		.INIT('h8)
	) name11856 (
		_w22318_,
		_w22319_,
		_w22368_
	);
	LUT2 #(
		.INIT('h8)
	) name11857 (
		_w22316_,
		_w22317_,
		_w22369_
	);
	LUT2 #(
		.INIT('h8)
	) name11858 (
		_w22314_,
		_w22315_,
		_w22370_
	);
	LUT2 #(
		.INIT('h8)
	) name11859 (
		_w22312_,
		_w22313_,
		_w22371_
	);
	LUT2 #(
		.INIT('h8)
	) name11860 (
		_w22310_,
		_w22311_,
		_w22372_
	);
	LUT2 #(
		.INIT('h8)
	) name11861 (
		_w22308_,
		_w22309_,
		_w22373_
	);
	LUT2 #(
		.INIT('h8)
	) name11862 (
		_w22306_,
		_w22307_,
		_w22374_
	);
	LUT2 #(
		.INIT('h8)
	) name11863 (
		_w22304_,
		_w22305_,
		_w22375_
	);
	LUT2 #(
		.INIT('h8)
	) name11864 (
		_w22302_,
		_w22303_,
		_w22376_
	);
	LUT2 #(
		.INIT('h8)
	) name11865 (
		_w22300_,
		_w22301_,
		_w22377_
	);
	LUT2 #(
		.INIT('h8)
	) name11866 (
		_w22298_,
		_w22299_,
		_w22378_
	);
	LUT2 #(
		.INIT('h8)
	) name11867 (
		_w22296_,
		_w22297_,
		_w22379_
	);
	LUT2 #(
		.INIT('h8)
	) name11868 (
		_w22294_,
		_w22295_,
		_w22380_
	);
	LUT2 #(
		.INIT('h8)
	) name11869 (
		_w22292_,
		_w22293_,
		_w22381_
	);
	LUT2 #(
		.INIT('h8)
	) name11870 (
		_w22290_,
		_w22291_,
		_w22382_
	);
	LUT2 #(
		.INIT('h8)
	) name11871 (
		_w22288_,
		_w22289_,
		_w22383_
	);
	LUT2 #(
		.INIT('h8)
	) name11872 (
		_w22382_,
		_w22383_,
		_w22384_
	);
	LUT2 #(
		.INIT('h8)
	) name11873 (
		_w22380_,
		_w22381_,
		_w22385_
	);
	LUT2 #(
		.INIT('h8)
	) name11874 (
		_w22378_,
		_w22379_,
		_w22386_
	);
	LUT2 #(
		.INIT('h8)
	) name11875 (
		_w22376_,
		_w22377_,
		_w22387_
	);
	LUT2 #(
		.INIT('h8)
	) name11876 (
		_w22374_,
		_w22375_,
		_w22388_
	);
	LUT2 #(
		.INIT('h8)
	) name11877 (
		_w22372_,
		_w22373_,
		_w22389_
	);
	LUT2 #(
		.INIT('h8)
	) name11878 (
		_w22370_,
		_w22371_,
		_w22390_
	);
	LUT2 #(
		.INIT('h8)
	) name11879 (
		_w22368_,
		_w22369_,
		_w22391_
	);
	LUT2 #(
		.INIT('h8)
	) name11880 (
		_w22366_,
		_w22367_,
		_w22392_
	);
	LUT2 #(
		.INIT('h8)
	) name11881 (
		_w22364_,
		_w22365_,
		_w22393_
	);
	LUT2 #(
		.INIT('h8)
	) name11882 (
		_w22362_,
		_w22363_,
		_w22394_
	);
	LUT2 #(
		.INIT('h8)
	) name11883 (
		_w22360_,
		_w22361_,
		_w22395_
	);
	LUT2 #(
		.INIT('h8)
	) name11884 (
		_w22358_,
		_w22359_,
		_w22396_
	);
	LUT2 #(
		.INIT('h8)
	) name11885 (
		_w22356_,
		_w22357_,
		_w22397_
	);
	LUT2 #(
		.INIT('h8)
	) name11886 (
		_w22354_,
		_w22355_,
		_w22398_
	);
	LUT2 #(
		.INIT('h8)
	) name11887 (
		_w22352_,
		_w22353_,
		_w22399_
	);
	LUT2 #(
		.INIT('h8)
	) name11888 (
		_w22398_,
		_w22399_,
		_w22400_
	);
	LUT2 #(
		.INIT('h8)
	) name11889 (
		_w22396_,
		_w22397_,
		_w22401_
	);
	LUT2 #(
		.INIT('h8)
	) name11890 (
		_w22394_,
		_w22395_,
		_w22402_
	);
	LUT2 #(
		.INIT('h8)
	) name11891 (
		_w22392_,
		_w22393_,
		_w22403_
	);
	LUT2 #(
		.INIT('h8)
	) name11892 (
		_w22390_,
		_w22391_,
		_w22404_
	);
	LUT2 #(
		.INIT('h8)
	) name11893 (
		_w22388_,
		_w22389_,
		_w22405_
	);
	LUT2 #(
		.INIT('h8)
	) name11894 (
		_w22386_,
		_w22387_,
		_w22406_
	);
	LUT2 #(
		.INIT('h8)
	) name11895 (
		_w22384_,
		_w22385_,
		_w22407_
	);
	LUT2 #(
		.INIT('h8)
	) name11896 (
		_w22406_,
		_w22407_,
		_w22408_
	);
	LUT2 #(
		.INIT('h8)
	) name11897 (
		_w22404_,
		_w22405_,
		_w22409_
	);
	LUT2 #(
		.INIT('h8)
	) name11898 (
		_w22402_,
		_w22403_,
		_w22410_
	);
	LUT2 #(
		.INIT('h8)
	) name11899 (
		_w22400_,
		_w22401_,
		_w22411_
	);
	LUT2 #(
		.INIT('h8)
	) name11900 (
		_w22410_,
		_w22411_,
		_w22412_
	);
	LUT2 #(
		.INIT('h8)
	) name11901 (
		_w22408_,
		_w22409_,
		_w22413_
	);
	LUT2 #(
		.INIT('h8)
	) name11902 (
		_w22412_,
		_w22413_,
		_w22414_
	);
	LUT2 #(
		.INIT('h1)
	) name11903 (
		wb_rst_i_pad,
		_w22414_,
		_w22415_
	);
	LUT2 #(
		.INIT('h8)
	) name11904 (
		_w12656_,
		_w22415_,
		_w22416_
	);
	LUT2 #(
		.INIT('h1)
	) name11905 (
		_w21903_,
		_w22416_,
		_w22417_
	);
	LUT2 #(
		.INIT('h2)
	) name11906 (
		\wishbone_LatchedTxLength_reg[8]/NET0131 ,
		_w12656_,
		_w22418_
	);
	LUT2 #(
		.INIT('h1)
	) name11907 (
		_w15111_,
		_w22418_,
		_w22419_
	);
	LUT2 #(
		.INIT('h2)
	) name11908 (
		\wishbone_LatchedTxLength_reg[6]/NET0131 ,
		_w12656_,
		_w22420_
	);
	LUT2 #(
		.INIT('h8)
	) name11909 (
		\wishbone_bd_ram_mem2_reg[189][22]/P0001 ,
		_w13042_,
		_w22421_
	);
	LUT2 #(
		.INIT('h8)
	) name11910 (
		\wishbone_bd_ram_mem2_reg[166][22]/P0001 ,
		_w13040_,
		_w22422_
	);
	LUT2 #(
		.INIT('h8)
	) name11911 (
		\wishbone_bd_ram_mem2_reg[44][22]/P0001 ,
		_w12896_,
		_w22423_
	);
	LUT2 #(
		.INIT('h8)
	) name11912 (
		\wishbone_bd_ram_mem2_reg[121][22]/P0001 ,
		_w13078_,
		_w22424_
	);
	LUT2 #(
		.INIT('h8)
	) name11913 (
		\wishbone_bd_ram_mem2_reg[56][22]/P0001 ,
		_w12778_,
		_w22425_
	);
	LUT2 #(
		.INIT('h8)
	) name11914 (
		\wishbone_bd_ram_mem2_reg[127][22]/P0001 ,
		_w13164_,
		_w22426_
	);
	LUT2 #(
		.INIT('h8)
	) name11915 (
		\wishbone_bd_ram_mem2_reg[49][22]/P0001 ,
		_w12994_,
		_w22427_
	);
	LUT2 #(
		.INIT('h8)
	) name11916 (
		\wishbone_bd_ram_mem2_reg[15][22]/P0001 ,
		_w13210_,
		_w22428_
	);
	LUT2 #(
		.INIT('h8)
	) name11917 (
		\wishbone_bd_ram_mem2_reg[156][22]/P0001 ,
		_w13190_,
		_w22429_
	);
	LUT2 #(
		.INIT('h8)
	) name11918 (
		\wishbone_bd_ram_mem2_reg[252][22]/P0001 ,
		_w13080_,
		_w22430_
	);
	LUT2 #(
		.INIT('h8)
	) name11919 (
		\wishbone_bd_ram_mem2_reg[175][22]/P0001 ,
		_w13126_,
		_w22431_
	);
	LUT2 #(
		.INIT('h8)
	) name11920 (
		\wishbone_bd_ram_mem2_reg[53][22]/P0001 ,
		_w13020_,
		_w22432_
	);
	LUT2 #(
		.INIT('h8)
	) name11921 (
		\wishbone_bd_ram_mem2_reg[38][22]/P0001 ,
		_w13182_,
		_w22433_
	);
	LUT2 #(
		.INIT('h8)
	) name11922 (
		\wishbone_bd_ram_mem2_reg[234][22]/P0001 ,
		_w13214_,
		_w22434_
	);
	LUT2 #(
		.INIT('h8)
	) name11923 (
		\wishbone_bd_ram_mem2_reg[20][22]/P0001 ,
		_w13174_,
		_w22435_
	);
	LUT2 #(
		.INIT('h8)
	) name11924 (
		\wishbone_bd_ram_mem2_reg[45][22]/P0001 ,
		_w12908_,
		_w22436_
	);
	LUT2 #(
		.INIT('h8)
	) name11925 (
		\wishbone_bd_ram_mem2_reg[200][22]/P0001 ,
		_w12988_,
		_w22437_
	);
	LUT2 #(
		.INIT('h8)
	) name11926 (
		\wishbone_bd_ram_mem2_reg[139][22]/P0001 ,
		_w12814_,
		_w22438_
	);
	LUT2 #(
		.INIT('h8)
	) name11927 (
		\wishbone_bd_ram_mem2_reg[61][22]/P0001 ,
		_w12725_,
		_w22439_
	);
	LUT2 #(
		.INIT('h8)
	) name11928 (
		\wishbone_bd_ram_mem2_reg[17][22]/P0001 ,
		_w12848_,
		_w22440_
	);
	LUT2 #(
		.INIT('h8)
	) name11929 (
		\wishbone_bd_ram_mem2_reg[160][22]/P0001 ,
		_w12872_,
		_w22441_
	);
	LUT2 #(
		.INIT('h8)
	) name11930 (
		\wishbone_bd_ram_mem2_reg[23][22]/P0001 ,
		_w13008_,
		_w22442_
	);
	LUT2 #(
		.INIT('h8)
	) name11931 (
		\wishbone_bd_ram_mem2_reg[191][22]/P0001 ,
		_w13034_,
		_w22443_
	);
	LUT2 #(
		.INIT('h8)
	) name11932 (
		\wishbone_bd_ram_mem2_reg[98][22]/P0001 ,
		_w12816_,
		_w22444_
	);
	LUT2 #(
		.INIT('h8)
	) name11933 (
		\wishbone_bd_ram_mem2_reg[75][22]/P0001 ,
		_w12826_,
		_w22445_
	);
	LUT2 #(
		.INIT('h8)
	) name11934 (
		\wishbone_bd_ram_mem2_reg[157][22]/P0001 ,
		_w12926_,
		_w22446_
	);
	LUT2 #(
		.INIT('h8)
	) name11935 (
		\wishbone_bd_ram_mem2_reg[145][22]/P0001 ,
		_w13106_,
		_w22447_
	);
	LUT2 #(
		.INIT('h8)
	) name11936 (
		\wishbone_bd_ram_mem2_reg[237][22]/P0001 ,
		_w12990_,
		_w22448_
	);
	LUT2 #(
		.INIT('h8)
	) name11937 (
		\wishbone_bd_ram_mem2_reg[112][22]/P0001 ,
		_w12733_,
		_w22449_
	);
	LUT2 #(
		.INIT('h8)
	) name11938 (
		\wishbone_bd_ram_mem2_reg[169][22]/P0001 ,
		_w12722_,
		_w22450_
	);
	LUT2 #(
		.INIT('h8)
	) name11939 (
		\wishbone_bd_ram_mem2_reg[105][22]/P0001 ,
		_w12751_,
		_w22451_
	);
	LUT2 #(
		.INIT('h8)
	) name11940 (
		\wishbone_bd_ram_mem2_reg[220][22]/P0001 ,
		_w13066_,
		_w22452_
	);
	LUT2 #(
		.INIT('h8)
	) name11941 (
		\wishbone_bd_ram_mem2_reg[100][22]/P0001 ,
		_w12960_,
		_w22453_
	);
	LUT2 #(
		.INIT('h8)
	) name11942 (
		\wishbone_bd_ram_mem2_reg[246][22]/P0001 ,
		_w13076_,
		_w22454_
	);
	LUT2 #(
		.INIT('h8)
	) name11943 (
		\wishbone_bd_ram_mem2_reg[10][22]/P0001 ,
		_w13172_,
		_w22455_
	);
	LUT2 #(
		.INIT('h8)
	) name11944 (
		\wishbone_bd_ram_mem2_reg[31][22]/P0001 ,
		_w13198_,
		_w22456_
	);
	LUT2 #(
		.INIT('h8)
	) name11945 (
		\wishbone_bd_ram_mem2_reg[18][22]/P0001 ,
		_w12679_,
		_w22457_
	);
	LUT2 #(
		.INIT('h8)
	) name11946 (
		\wishbone_bd_ram_mem2_reg[55][22]/P0001 ,
		_w12785_,
		_w22458_
	);
	LUT2 #(
		.INIT('h8)
	) name11947 (
		\wishbone_bd_ram_mem2_reg[77][22]/P0001 ,
		_w12982_,
		_w22459_
	);
	LUT2 #(
		.INIT('h8)
	) name11948 (
		\wishbone_bd_ram_mem2_reg[66][22]/P0001 ,
		_w12824_,
		_w22460_
	);
	LUT2 #(
		.INIT('h8)
	) name11949 (
		\wishbone_bd_ram_mem2_reg[114][22]/P0001 ,
		_w13202_,
		_w22461_
	);
	LUT2 #(
		.INIT('h8)
	) name11950 (
		\wishbone_bd_ram_mem2_reg[208][22]/P0001 ,
		_w13032_,
		_w22462_
	);
	LUT2 #(
		.INIT('h8)
	) name11951 (
		\wishbone_bd_ram_mem2_reg[95][22]/P0001 ,
		_w12844_,
		_w22463_
	);
	LUT2 #(
		.INIT('h8)
	) name11952 (
		\wishbone_bd_ram_mem2_reg[24][22]/P0001 ,
		_w13084_,
		_w22464_
	);
	LUT2 #(
		.INIT('h8)
	) name11953 (
		\wishbone_bd_ram_mem2_reg[203][22]/P0001 ,
		_w13158_,
		_w22465_
	);
	LUT2 #(
		.INIT('h8)
	) name11954 (
		\wishbone_bd_ram_mem2_reg[232][22]/P0001 ,
		_w12758_,
		_w22466_
	);
	LUT2 #(
		.INIT('h8)
	) name11955 (
		\wishbone_bd_ram_mem2_reg[159][22]/P0001 ,
		_w12774_,
		_w22467_
	);
	LUT2 #(
		.INIT('h8)
	) name11956 (
		\wishbone_bd_ram_mem2_reg[233][22]/P0001 ,
		_w12836_,
		_w22468_
	);
	LUT2 #(
		.INIT('h8)
	) name11957 (
		\wishbone_bd_ram_mem2_reg[244][22]/P0001 ,
		_w12747_,
		_w22469_
	);
	LUT2 #(
		.INIT('h8)
	) name11958 (
		\wishbone_bd_ram_mem2_reg[215][22]/P0001 ,
		_w12974_,
		_w22470_
	);
	LUT2 #(
		.INIT('h8)
	) name11959 (
		\wishbone_bd_ram_mem2_reg[217][22]/P0001 ,
		_w13188_,
		_w22471_
	);
	LUT2 #(
		.INIT('h8)
	) name11960 (
		\wishbone_bd_ram_mem2_reg[34][22]/P0001 ,
		_w12930_,
		_w22472_
	);
	LUT2 #(
		.INIT('h8)
	) name11961 (
		\wishbone_bd_ram_mem2_reg[35][22]/P0001 ,
		_w12703_,
		_w22473_
	);
	LUT2 #(
		.INIT('h8)
	) name11962 (
		\wishbone_bd_ram_mem2_reg[184][22]/P0001 ,
		_w13062_,
		_w22474_
	);
	LUT2 #(
		.INIT('h8)
	) name11963 (
		\wishbone_bd_ram_mem2_reg[16][22]/P0001 ,
		_w13140_,
		_w22475_
	);
	LUT2 #(
		.INIT('h8)
	) name11964 (
		\wishbone_bd_ram_mem2_reg[130][22]/P0001 ,
		_w12914_,
		_w22476_
	);
	LUT2 #(
		.INIT('h8)
	) name11965 (
		\wishbone_bd_ram_mem2_reg[143][22]/P0001 ,
		_w12922_,
		_w22477_
	);
	LUT2 #(
		.INIT('h8)
	) name11966 (
		\wishbone_bd_ram_mem2_reg[96][22]/P0001 ,
		_w12912_,
		_w22478_
	);
	LUT2 #(
		.INIT('h8)
	) name11967 (
		\wishbone_bd_ram_mem2_reg[136][22]/P0001 ,
		_w13064_,
		_w22479_
	);
	LUT2 #(
		.INIT('h8)
	) name11968 (
		\wishbone_bd_ram_mem2_reg[137][22]/P0001 ,
		_w13168_,
		_w22480_
	);
	LUT2 #(
		.INIT('h8)
	) name11969 (
		\wishbone_bd_ram_mem2_reg[207][22]/P0001 ,
		_w13180_,
		_w22481_
	);
	LUT2 #(
		.INIT('h8)
	) name11970 (
		\wishbone_bd_ram_mem2_reg[26][22]/P0001 ,
		_w12699_,
		_w22482_
	);
	LUT2 #(
		.INIT('h8)
	) name11971 (
		\wishbone_bd_ram_mem2_reg[154][22]/P0001 ,
		_w12962_,
		_w22483_
	);
	LUT2 #(
		.INIT('h8)
	) name11972 (
		\wishbone_bd_ram_mem2_reg[113][22]/P0001 ,
		_w13026_,
		_w22484_
	);
	LUT2 #(
		.INIT('h8)
	) name11973 (
		\wishbone_bd_ram_mem2_reg[248][22]/P0001 ,
		_w12789_,
		_w22485_
	);
	LUT2 #(
		.INIT('h8)
	) name11974 (
		\wishbone_bd_ram_mem2_reg[164][22]/P0001 ,
		_w12876_,
		_w22486_
	);
	LUT2 #(
		.INIT('h8)
	) name11975 (
		\wishbone_bd_ram_mem2_reg[251][22]/P0001 ,
		_w13054_,
		_w22487_
	);
	LUT2 #(
		.INIT('h8)
	) name11976 (
		\wishbone_bd_ram_mem2_reg[50][22]/P0001 ,
		_w13150_,
		_w22488_
	);
	LUT2 #(
		.INIT('h8)
	) name11977 (
		\wishbone_bd_ram_mem2_reg[42][22]/P0001 ,
		_w12842_,
		_w22489_
	);
	LUT2 #(
		.INIT('h8)
	) name11978 (
		\wishbone_bd_ram_mem2_reg[107][22]/P0001 ,
		_w12749_,
		_w22490_
	);
	LUT2 #(
		.INIT('h8)
	) name11979 (
		\wishbone_bd_ram_mem2_reg[2][22]/P0001 ,
		_w13088_,
		_w22491_
	);
	LUT2 #(
		.INIT('h8)
	) name11980 (
		\wishbone_bd_ram_mem2_reg[138][22]/P0001 ,
		_w12958_,
		_w22492_
	);
	LUT2 #(
		.INIT('h8)
	) name11981 (
		\wishbone_bd_ram_mem2_reg[30][22]/P0001 ,
		_w13104_,
		_w22493_
	);
	LUT2 #(
		.INIT('h8)
	) name11982 (
		\wishbone_bd_ram_mem2_reg[212][22]/P0001 ,
		_w12796_,
		_w22494_
	);
	LUT2 #(
		.INIT('h8)
	) name11983 (
		\wishbone_bd_ram_mem2_reg[146][22]/P0001 ,
		_w13060_,
		_w22495_
	);
	LUT2 #(
		.INIT('h8)
	) name11984 (
		\wishbone_bd_ram_mem2_reg[206][22]/P0001 ,
		_w12954_,
		_w22496_
	);
	LUT2 #(
		.INIT('h8)
	) name11985 (
		\wishbone_bd_ram_mem2_reg[174][22]/P0001 ,
		_w12972_,
		_w22497_
	);
	LUT2 #(
		.INIT('h8)
	) name11986 (
		\wishbone_bd_ram_mem2_reg[165][22]/P0001 ,
		_w13044_,
		_w22498_
	);
	LUT2 #(
		.INIT('h8)
	) name11987 (
		\wishbone_bd_ram_mem2_reg[226][22]/P0001 ,
		_w13138_,
		_w22499_
	);
	LUT2 #(
		.INIT('h8)
	) name11988 (
		\wishbone_bd_ram_mem2_reg[243][22]/P0001 ,
		_w12804_,
		_w22500_
	);
	LUT2 #(
		.INIT('h8)
	) name11989 (
		\wishbone_bd_ram_mem2_reg[202][22]/P0001 ,
		_w12870_,
		_w22501_
	);
	LUT2 #(
		.INIT('h8)
	) name11990 (
		\wishbone_bd_ram_mem2_reg[228][22]/P0001 ,
		_w12765_,
		_w22502_
	);
	LUT2 #(
		.INIT('h8)
	) name11991 (
		\wishbone_bd_ram_mem2_reg[64][22]/P0001 ,
		_w12976_,
		_w22503_
	);
	LUT2 #(
		.INIT('h8)
	) name11992 (
		\wishbone_bd_ram_mem2_reg[247][22]/P0001 ,
		_w12818_,
		_w22504_
	);
	LUT2 #(
		.INIT('h8)
	) name11993 (
		\wishbone_bd_ram_mem2_reg[86][22]/P0001 ,
		_w12735_,
		_w22505_
	);
	LUT2 #(
		.INIT('h8)
	) name11994 (
		\wishbone_bd_ram_mem2_reg[79][22]/P0001 ,
		_w13212_,
		_w22506_
	);
	LUT2 #(
		.INIT('h8)
	) name11995 (
		\wishbone_bd_ram_mem2_reg[52][22]/P0001 ,
		_w13082_,
		_w22507_
	);
	LUT2 #(
		.INIT('h8)
	) name11996 (
		\wishbone_bd_ram_mem2_reg[74][22]/P0001 ,
		_w12812_,
		_w22508_
	);
	LUT2 #(
		.INIT('h8)
	) name11997 (
		\wishbone_bd_ram_mem2_reg[32][22]/P0001 ,
		_w13120_,
		_w22509_
	);
	LUT2 #(
		.INIT('h8)
	) name11998 (
		\wishbone_bd_ram_mem2_reg[194][22]/P0001 ,
		_w12772_,
		_w22510_
	);
	LUT2 #(
		.INIT('h8)
	) name11999 (
		\wishbone_bd_ram_mem2_reg[51][22]/P0001 ,
		_w13024_,
		_w22511_
	);
	LUT2 #(
		.INIT('h8)
	) name12000 (
		\wishbone_bd_ram_mem2_reg[180][22]/P0001 ,
		_w12791_,
		_w22512_
	);
	LUT2 #(
		.INIT('h8)
	) name12001 (
		\wishbone_bd_ram_mem2_reg[133][22]/P0001 ,
		_w12761_,
		_w22513_
	);
	LUT2 #(
		.INIT('h8)
	) name12002 (
		\wishbone_bd_ram_mem2_reg[204][22]/P0001 ,
		_w13162_,
		_w22514_
	);
	LUT2 #(
		.INIT('h8)
	) name12003 (
		\wishbone_bd_ram_mem2_reg[135][22]/P0001 ,
		_w13124_,
		_w22515_
	);
	LUT2 #(
		.INIT('h8)
	) name12004 (
		\wishbone_bd_ram_mem2_reg[111][22]/P0001 ,
		_w12744_,
		_w22516_
	);
	LUT2 #(
		.INIT('h8)
	) name12005 (
		\wishbone_bd_ram_mem2_reg[214][22]/P0001 ,
		_w12984_,
		_w22517_
	);
	LUT2 #(
		.INIT('h8)
	) name12006 (
		\wishbone_bd_ram_mem2_reg[173][22]/P0001 ,
		_w12854_,
		_w22518_
	);
	LUT2 #(
		.INIT('h8)
	) name12007 (
		\wishbone_bd_ram_mem2_reg[60][22]/P0001 ,
		_w13204_,
		_w22519_
	);
	LUT2 #(
		.INIT('h8)
	) name12008 (
		\wishbone_bd_ram_mem2_reg[5][22]/P0001 ,
		_w12878_,
		_w22520_
	);
	LUT2 #(
		.INIT('h8)
	) name12009 (
		\wishbone_bd_ram_mem2_reg[116][22]/P0001 ,
		_w12998_,
		_w22521_
	);
	LUT2 #(
		.INIT('h8)
	) name12010 (
		\wishbone_bd_ram_mem2_reg[144][22]/P0001 ,
		_w12756_,
		_w22522_
	);
	LUT2 #(
		.INIT('h8)
	) name12011 (
		\wishbone_bd_ram_mem2_reg[80][22]/P0001 ,
		_w12689_,
		_w22523_
	);
	LUT2 #(
		.INIT('h8)
	) name12012 (
		\wishbone_bd_ram_mem2_reg[108][22]/P0001 ,
		_w13156_,
		_w22524_
	);
	LUT2 #(
		.INIT('h8)
	) name12013 (
		\wishbone_bd_ram_mem2_reg[76][22]/P0001 ,
		_w13184_,
		_w22525_
	);
	LUT2 #(
		.INIT('h8)
	) name12014 (
		\wishbone_bd_ram_mem2_reg[14][22]/P0001 ,
		_w13086_,
		_w22526_
	);
	LUT2 #(
		.INIT('h8)
	) name12015 (
		\wishbone_bd_ram_mem2_reg[57][22]/P0001 ,
		_w13116_,
		_w22527_
	);
	LUT2 #(
		.INIT('h8)
	) name12016 (
		\wishbone_bd_ram_mem2_reg[153][22]/P0001 ,
		_w12890_,
		_w22528_
	);
	LUT2 #(
		.INIT('h8)
	) name12017 (
		\wishbone_bd_ram_mem2_reg[97][22]/P0001 ,
		_w13096_,
		_w22529_
	);
	LUT2 #(
		.INIT('h8)
	) name12018 (
		\wishbone_bd_ram_mem2_reg[141][22]/P0001 ,
		_w13004_,
		_w22530_
	);
	LUT2 #(
		.INIT('h8)
	) name12019 (
		\wishbone_bd_ram_mem2_reg[58][22]/P0001 ,
		_w13070_,
		_w22531_
	);
	LUT2 #(
		.INIT('h8)
	) name12020 (
		\wishbone_bd_ram_mem2_reg[0][22]/P0001 ,
		_w12717_,
		_w22532_
	);
	LUT2 #(
		.INIT('h8)
	) name12021 (
		\wishbone_bd_ram_mem2_reg[106][22]/P0001 ,
		_w12713_,
		_w22533_
	);
	LUT2 #(
		.INIT('h8)
	) name12022 (
		\wishbone_bd_ram_mem2_reg[85][22]/P0001 ,
		_w13216_,
		_w22534_
	);
	LUT2 #(
		.INIT('h8)
	) name12023 (
		\wishbone_bd_ram_mem2_reg[221][22]/P0001 ,
		_w12802_,
		_w22535_
	);
	LUT2 #(
		.INIT('h8)
	) name12024 (
		\wishbone_bd_ram_mem2_reg[128][22]/P0001 ,
		_w12793_,
		_w22536_
	);
	LUT2 #(
		.INIT('h8)
	) name12025 (
		\wishbone_bd_ram_mem2_reg[140][22]/P0001 ,
		_w12894_,
		_w22537_
	);
	LUT2 #(
		.INIT('h8)
	) name12026 (
		\wishbone_bd_ram_mem2_reg[59][22]/P0001 ,
		_w12780_,
		_w22538_
	);
	LUT2 #(
		.INIT('h8)
	) name12027 (
		\wishbone_bd_ram_mem2_reg[176][22]/P0001 ,
		_w12868_,
		_w22539_
	);
	LUT2 #(
		.INIT('h8)
	) name12028 (
		\wishbone_bd_ram_mem2_reg[67][22]/P0001 ,
		_w13134_,
		_w22540_
	);
	LUT2 #(
		.INIT('h8)
	) name12029 (
		\wishbone_bd_ram_mem2_reg[222][22]/P0001 ,
		_w13094_,
		_w22541_
	);
	LUT2 #(
		.INIT('h8)
	) name12030 (
		\wishbone_bd_ram_mem2_reg[254][22]/P0001 ,
		_w12892_,
		_w22542_
	);
	LUT2 #(
		.INIT('h8)
	) name12031 (
		\wishbone_bd_ram_mem2_reg[148][22]/P0001 ,
		_w13000_,
		_w22543_
	);
	LUT2 #(
		.INIT('h8)
	) name12032 (
		\wishbone_bd_ram_mem2_reg[239][22]/P0001 ,
		_w12862_,
		_w22544_
	);
	LUT2 #(
		.INIT('h8)
	) name12033 (
		\wishbone_bd_ram_mem2_reg[104][22]/P0001 ,
		_w13148_,
		_w22545_
	);
	LUT2 #(
		.INIT('h8)
	) name12034 (
		\wishbone_bd_ram_mem2_reg[41][22]/P0001 ,
		_w13052_,
		_w22546_
	);
	LUT2 #(
		.INIT('h8)
	) name12035 (
		\wishbone_bd_ram_mem2_reg[63][22]/P0001 ,
		_w12850_,
		_w22547_
	);
	LUT2 #(
		.INIT('h8)
	) name12036 (
		\wishbone_bd_ram_mem2_reg[210][22]/P0001 ,
		_w12924_,
		_w22548_
	);
	LUT2 #(
		.INIT('h8)
	) name12037 (
		\wishbone_bd_ram_mem2_reg[192][22]/P0001 ,
		_w12938_,
		_w22549_
	);
	LUT2 #(
		.INIT('h8)
	) name12038 (
		\wishbone_bd_ram_mem2_reg[134][22]/P0001 ,
		_w12763_,
		_w22550_
	);
	LUT2 #(
		.INIT('h8)
	) name12039 (
		\wishbone_bd_ram_mem2_reg[225][22]/P0001 ,
		_w13092_,
		_w22551_
	);
	LUT2 #(
		.INIT('h8)
	) name12040 (
		\wishbone_bd_ram_mem2_reg[91][22]/P0001 ,
		_w13074_,
		_w22552_
	);
	LUT2 #(
		.INIT('h8)
	) name12041 (
		\wishbone_bd_ram_mem2_reg[151][22]/P0001 ,
		_w13142_,
		_w22553_
	);
	LUT2 #(
		.INIT('h8)
	) name12042 (
		\wishbone_bd_ram_mem2_reg[6][22]/P0001 ,
		_w12968_,
		_w22554_
	);
	LUT2 #(
		.INIT('h8)
	) name12043 (
		\wishbone_bd_ram_mem2_reg[230][22]/P0001 ,
		_w13036_,
		_w22555_
	);
	LUT2 #(
		.INIT('h8)
	) name12044 (
		\wishbone_bd_ram_mem2_reg[102][22]/P0001 ,
		_w12685_,
		_w22556_
	);
	LUT2 #(
		.INIT('h8)
	) name12045 (
		\wishbone_bd_ram_mem2_reg[40][22]/P0001 ,
		_w13132_,
		_w22557_
	);
	LUT2 #(
		.INIT('h8)
	) name12046 (
		\wishbone_bd_ram_mem2_reg[65][22]/P0001 ,
		_w13176_,
		_w22558_
	);
	LUT2 #(
		.INIT('h8)
	) name12047 (
		\wishbone_bd_ram_mem2_reg[213][22]/P0001 ,
		_w13002_,
		_w22559_
	);
	LUT2 #(
		.INIT('h8)
	) name12048 (
		\wishbone_bd_ram_mem2_reg[71][22]/P0001 ,
		_w12798_,
		_w22560_
	);
	LUT2 #(
		.INIT('h8)
	) name12049 (
		\wishbone_bd_ram_mem2_reg[224][22]/P0001 ,
		_w12902_,
		_w22561_
	);
	LUT2 #(
		.INIT('h8)
	) name12050 (
		\wishbone_bd_ram_mem2_reg[186][22]/P0001 ,
		_w12783_,
		_w22562_
	);
	LUT2 #(
		.INIT('h8)
	) name12051 (
		\wishbone_bd_ram_mem2_reg[193][22]/P0001 ,
		_w13056_,
		_w22563_
	);
	LUT2 #(
		.INIT('h8)
	) name12052 (
		\wishbone_bd_ram_mem2_reg[78][22]/P0001 ,
		_w12874_,
		_w22564_
	);
	LUT2 #(
		.INIT('h8)
	) name12053 (
		\wishbone_bd_ram_mem2_reg[170][22]/P0001 ,
		_w13030_,
		_w22565_
	);
	LUT2 #(
		.INIT('h8)
	) name12054 (
		\wishbone_bd_ram_mem2_reg[152][22]/P0001 ,
		_w12966_,
		_w22566_
	);
	LUT2 #(
		.INIT('h8)
	) name12055 (
		\wishbone_bd_ram_mem2_reg[62][22]/P0001 ,
		_w12673_,
		_w22567_
	);
	LUT2 #(
		.INIT('h8)
	) name12056 (
		\wishbone_bd_ram_mem2_reg[229][22]/P0001 ,
		_w12711_,
		_w22568_
	);
	LUT2 #(
		.INIT('h8)
	) name12057 (
		\wishbone_bd_ram_mem2_reg[70][22]/P0001 ,
		_w12840_,
		_w22569_
	);
	LUT2 #(
		.INIT('h8)
	) name12058 (
		\wishbone_bd_ram_mem2_reg[129][22]/P0001 ,
		_w12776_,
		_w22570_
	);
	LUT2 #(
		.INIT('h8)
	) name12059 (
		\wishbone_bd_ram_mem2_reg[54][22]/P0001 ,
		_w12770_,
		_w22571_
	);
	LUT2 #(
		.INIT('h8)
	) name12060 (
		\wishbone_bd_ram_mem2_reg[73][22]/P0001 ,
		_w12918_,
		_w22572_
	);
	LUT2 #(
		.INIT('h8)
	) name12061 (
		\wishbone_bd_ram_mem2_reg[163][22]/P0001 ,
		_w12882_,
		_w22573_
	);
	LUT2 #(
		.INIT('h8)
	) name12062 (
		\wishbone_bd_ram_mem2_reg[255][22]/P0001 ,
		_w13072_,
		_w22574_
	);
	LUT2 #(
		.INIT('h8)
	) name12063 (
		\wishbone_bd_ram_mem2_reg[99][22]/P0001 ,
		_w13038_,
		_w22575_
	);
	LUT2 #(
		.INIT('h8)
	) name12064 (
		\wishbone_bd_ram_mem2_reg[119][22]/P0001 ,
		_w13048_,
		_w22576_
	);
	LUT2 #(
		.INIT('h8)
	) name12065 (
		\wishbone_bd_ram_mem2_reg[81][22]/P0001 ,
		_w12950_,
		_w22577_
	);
	LUT2 #(
		.INIT('h8)
	) name12066 (
		\wishbone_bd_ram_mem2_reg[238][22]/P0001 ,
		_w13160_,
		_w22578_
	);
	LUT2 #(
		.INIT('h8)
	) name12067 (
		\wishbone_bd_ram_mem2_reg[28][22]/P0001 ,
		_w13170_,
		_w22579_
	);
	LUT2 #(
		.INIT('h8)
	) name12068 (
		\wishbone_bd_ram_mem2_reg[183][22]/P0001 ,
		_w12787_,
		_w22580_
	);
	LUT2 #(
		.INIT('h8)
	) name12069 (
		\wishbone_bd_ram_mem2_reg[245][22]/P0001 ,
		_w13022_,
		_w22581_
	);
	LUT2 #(
		.INIT('h8)
	) name12070 (
		\wishbone_bd_ram_mem2_reg[236][22]/P0001 ,
		_w12731_,
		_w22582_
	);
	LUT2 #(
		.INIT('h8)
	) name12071 (
		\wishbone_bd_ram_mem2_reg[218][22]/P0001 ,
		_w13206_,
		_w22583_
	);
	LUT2 #(
		.INIT('h8)
	) name12072 (
		\wishbone_bd_ram_mem2_reg[162][22]/P0001 ,
		_w13098_,
		_w22584_
	);
	LUT2 #(
		.INIT('h8)
	) name12073 (
		\wishbone_bd_ram_mem2_reg[231][22]/P0001 ,
		_w12856_,
		_w22585_
	);
	LUT2 #(
		.INIT('h8)
	) name12074 (
		\wishbone_bd_ram_mem2_reg[123][22]/P0001 ,
		_w13114_,
		_w22586_
	);
	LUT2 #(
		.INIT('h8)
	) name12075 (
		\wishbone_bd_ram_mem2_reg[171][22]/P0001 ,
		_w12910_,
		_w22587_
	);
	LUT2 #(
		.INIT('h8)
	) name12076 (
		\wishbone_bd_ram_mem2_reg[103][22]/P0001 ,
		_w12846_,
		_w22588_
	);
	LUT2 #(
		.INIT('h8)
	) name12077 (
		\wishbone_bd_ram_mem2_reg[93][22]/P0001 ,
		_w13016_,
		_w22589_
	);
	LUT2 #(
		.INIT('h8)
	) name12078 (
		\wishbone_bd_ram_mem2_reg[158][22]/P0001 ,
		_w12898_,
		_w22590_
	);
	LUT2 #(
		.INIT('h8)
	) name12079 (
		\wishbone_bd_ram_mem2_reg[33][22]/P0001 ,
		_w12980_,
		_w22591_
	);
	LUT2 #(
		.INIT('h8)
	) name12080 (
		\wishbone_bd_ram_mem2_reg[205][22]/P0001 ,
		_w13068_,
		_w22592_
	);
	LUT2 #(
		.INIT('h8)
	) name12081 (
		\wishbone_bd_ram_mem2_reg[46][22]/P0001 ,
		_w12884_,
		_w22593_
	);
	LUT2 #(
		.INIT('h8)
	) name12082 (
		\wishbone_bd_ram_mem2_reg[178][22]/P0001 ,
		_w12886_,
		_w22594_
	);
	LUT2 #(
		.INIT('h8)
	) name12083 (
		\wishbone_bd_ram_mem2_reg[198][22]/P0001 ,
		_w12832_,
		_w22595_
	);
	LUT2 #(
		.INIT('h8)
	) name12084 (
		\wishbone_bd_ram_mem2_reg[132][22]/P0001 ,
		_w12992_,
		_w22596_
	);
	LUT2 #(
		.INIT('h8)
	) name12085 (
		\wishbone_bd_ram_mem2_reg[92][22]/P0001 ,
		_w13010_,
		_w22597_
	);
	LUT2 #(
		.INIT('h8)
	) name12086 (
		\wishbone_bd_ram_mem2_reg[195][22]/P0001 ,
		_w13144_,
		_w22598_
	);
	LUT2 #(
		.INIT('h8)
	) name12087 (
		\wishbone_bd_ram_mem2_reg[150][22]/P0001 ,
		_w13136_,
		_w22599_
	);
	LUT2 #(
		.INIT('h8)
	) name12088 (
		\wishbone_bd_ram_mem2_reg[211][22]/P0001 ,
		_w13166_,
		_w22600_
	);
	LUT2 #(
		.INIT('h8)
	) name12089 (
		\wishbone_bd_ram_mem2_reg[199][22]/P0001 ,
		_w12768_,
		_w22601_
	);
	LUT2 #(
		.INIT('h8)
	) name12090 (
		\wishbone_bd_ram_mem2_reg[235][22]/P0001 ,
		_w12696_,
		_w22602_
	);
	LUT2 #(
		.INIT('h8)
	) name12091 (
		\wishbone_bd_ram_mem2_reg[185][22]/P0001 ,
		_w12940_,
		_w22603_
	);
	LUT2 #(
		.INIT('h8)
	) name12092 (
		\wishbone_bd_ram_mem2_reg[241][22]/P0001 ,
		_w13006_,
		_w22604_
	);
	LUT2 #(
		.INIT('h8)
	) name12093 (
		\wishbone_bd_ram_mem2_reg[227][22]/P0001 ,
		_w12936_,
		_w22605_
	);
	LUT2 #(
		.INIT('h8)
	) name12094 (
		\wishbone_bd_ram_mem2_reg[182][22]/P0001 ,
		_w12820_,
		_w22606_
	);
	LUT2 #(
		.INIT('h8)
	) name12095 (
		\wishbone_bd_ram_mem2_reg[219][22]/P0001 ,
		_w12806_,
		_w22607_
	);
	LUT2 #(
		.INIT('h8)
	) name12096 (
		\wishbone_bd_ram_mem2_reg[3][22]/P0001 ,
		_w12866_,
		_w22608_
	);
	LUT2 #(
		.INIT('h8)
	) name12097 (
		\wishbone_bd_ram_mem2_reg[13][22]/P0001 ,
		_w13178_,
		_w22609_
	);
	LUT2 #(
		.INIT('h8)
	) name12098 (
		\wishbone_bd_ram_mem2_reg[101][22]/P0001 ,
		_w13192_,
		_w22610_
	);
	LUT2 #(
		.INIT('h8)
	) name12099 (
		\wishbone_bd_ram_mem2_reg[43][22]/P0001 ,
		_w13200_,
		_w22611_
	);
	LUT2 #(
		.INIT('h8)
	) name12100 (
		\wishbone_bd_ram_mem2_reg[110][22]/P0001 ,
		_w13046_,
		_w22612_
	);
	LUT2 #(
		.INIT('h8)
	) name12101 (
		\wishbone_bd_ram_mem2_reg[187][22]/P0001 ,
		_w13196_,
		_w22613_
	);
	LUT2 #(
		.INIT('h8)
	) name12102 (
		\wishbone_bd_ram_mem2_reg[172][22]/P0001 ,
		_w12944_,
		_w22614_
	);
	LUT2 #(
		.INIT('h8)
	) name12103 (
		\wishbone_bd_ram_mem2_reg[109][22]/P0001 ,
		_w12888_,
		_w22615_
	);
	LUT2 #(
		.INIT('h8)
	) name12104 (
		\wishbone_bd_ram_mem2_reg[82][22]/P0001 ,
		_w12942_,
		_w22616_
	);
	LUT2 #(
		.INIT('h8)
	) name12105 (
		\wishbone_bd_ram_mem2_reg[250][22]/P0001 ,
		_w13128_,
		_w22617_
	);
	LUT2 #(
		.INIT('h8)
	) name12106 (
		\wishbone_bd_ram_mem2_reg[12][22]/P0001 ,
		_w13118_,
		_w22618_
	);
	LUT2 #(
		.INIT('h8)
	) name12107 (
		\wishbone_bd_ram_mem2_reg[27][22]/P0001 ,
		_w12880_,
		_w22619_
	);
	LUT2 #(
		.INIT('h8)
	) name12108 (
		\wishbone_bd_ram_mem2_reg[88][22]/P0001 ,
		_w12860_,
		_w22620_
	);
	LUT2 #(
		.INIT('h8)
	) name12109 (
		\wishbone_bd_ram_mem2_reg[11][22]/P0001 ,
		_w13194_,
		_w22621_
	);
	LUT2 #(
		.INIT('h8)
	) name12110 (
		\wishbone_bd_ram_mem2_reg[147][22]/P0001 ,
		_w13146_,
		_w22622_
	);
	LUT2 #(
		.INIT('h8)
	) name12111 (
		\wishbone_bd_ram_mem2_reg[36][22]/P0001 ,
		_w12800_,
		_w22623_
	);
	LUT2 #(
		.INIT('h8)
	) name12112 (
		\wishbone_bd_ram_mem2_reg[87][22]/P0001 ,
		_w13154_,
		_w22624_
	);
	LUT2 #(
		.INIT('h8)
	) name12113 (
		\wishbone_bd_ram_mem2_reg[131][22]/P0001 ,
		_w12852_,
		_w22625_
	);
	LUT2 #(
		.INIT('h8)
	) name12114 (
		\wishbone_bd_ram_mem2_reg[68][22]/P0001 ,
		_w12946_,
		_w22626_
	);
	LUT2 #(
		.INIT('h8)
	) name12115 (
		\wishbone_bd_ram_mem2_reg[196][22]/P0001 ,
		_w13090_,
		_w22627_
	);
	LUT2 #(
		.INIT('h8)
	) name12116 (
		\wishbone_bd_ram_mem2_reg[115][22]/P0001 ,
		_w13112_,
		_w22628_
	);
	LUT2 #(
		.INIT('h8)
	) name12117 (
		\wishbone_bd_ram_mem2_reg[149][22]/P0001 ,
		_w12741_,
		_w22629_
	);
	LUT2 #(
		.INIT('h8)
	) name12118 (
		\wishbone_bd_ram_mem2_reg[1][22]/P0001 ,
		_w13014_,
		_w22630_
	);
	LUT2 #(
		.INIT('h8)
	) name12119 (
		\wishbone_bd_ram_mem2_reg[201][22]/P0001 ,
		_w12822_,
		_w22631_
	);
	LUT2 #(
		.INIT('h8)
	) name12120 (
		\wishbone_bd_ram_mem2_reg[117][22]/P0001 ,
		_w12715_,
		_w22632_
	);
	LUT2 #(
		.INIT('h8)
	) name12121 (
		\wishbone_bd_ram_mem2_reg[4][22]/P0001 ,
		_w12666_,
		_w22633_
	);
	LUT2 #(
		.INIT('h8)
	) name12122 (
		\wishbone_bd_ram_mem2_reg[21][22]/P0001 ,
		_w12906_,
		_w22634_
	);
	LUT2 #(
		.INIT('h8)
	) name12123 (
		\wishbone_bd_ram_mem2_reg[167][22]/P0001 ,
		_w12986_,
		_w22635_
	);
	LUT2 #(
		.INIT('h8)
	) name12124 (
		\wishbone_bd_ram_mem2_reg[181][22]/P0001 ,
		_w12828_,
		_w22636_
	);
	LUT2 #(
		.INIT('h8)
	) name12125 (
		\wishbone_bd_ram_mem2_reg[47][22]/P0001 ,
		_w12904_,
		_w22637_
	);
	LUT2 #(
		.INIT('h8)
	) name12126 (
		\wishbone_bd_ram_mem2_reg[125][22]/P0001 ,
		_w12956_,
		_w22638_
	);
	LUT2 #(
		.INIT('h8)
	) name12127 (
		\wishbone_bd_ram_mem2_reg[216][22]/P0001 ,
		_w13028_,
		_w22639_
	);
	LUT2 #(
		.INIT('h8)
	) name12128 (
		\wishbone_bd_ram_mem2_reg[19][22]/P0001 ,
		_w13012_,
		_w22640_
	);
	LUT2 #(
		.INIT('h8)
	) name12129 (
		\wishbone_bd_ram_mem2_reg[72][22]/P0001 ,
		_w12810_,
		_w22641_
	);
	LUT2 #(
		.INIT('h8)
	) name12130 (
		\wishbone_bd_ram_mem2_reg[9][22]/P0001 ,
		_w12808_,
		_w22642_
	);
	LUT2 #(
		.INIT('h8)
	) name12131 (
		\wishbone_bd_ram_mem2_reg[90][22]/P0001 ,
		_w12978_,
		_w22643_
	);
	LUT2 #(
		.INIT('h8)
	) name12132 (
		\wishbone_bd_ram_mem2_reg[168][22]/P0001 ,
		_w13208_,
		_w22644_
	);
	LUT2 #(
		.INIT('h8)
	) name12133 (
		\wishbone_bd_ram_mem2_reg[120][22]/P0001 ,
		_w12707_,
		_w22645_
	);
	LUT2 #(
		.INIT('h8)
	) name12134 (
		\wishbone_bd_ram_mem2_reg[242][22]/P0001 ,
		_w12932_,
		_w22646_
	);
	LUT2 #(
		.INIT('h8)
	) name12135 (
		\wishbone_bd_ram_mem2_reg[249][22]/P0001 ,
		_w12900_,
		_w22647_
	);
	LUT2 #(
		.INIT('h8)
	) name12136 (
		\wishbone_bd_ram_mem2_reg[223][22]/P0001 ,
		_w12838_,
		_w22648_
	);
	LUT2 #(
		.INIT('h8)
	) name12137 (
		\wishbone_bd_ram_mem2_reg[179][22]/P0001 ,
		_w13050_,
		_w22649_
	);
	LUT2 #(
		.INIT('h8)
	) name12138 (
		\wishbone_bd_ram_mem2_reg[126][22]/P0001 ,
		_w13218_,
		_w22650_
	);
	LUT2 #(
		.INIT('h8)
	) name12139 (
		\wishbone_bd_ram_mem2_reg[7][22]/P0001 ,
		_w12728_,
		_w22651_
	);
	LUT2 #(
		.INIT('h8)
	) name12140 (
		\wishbone_bd_ram_mem2_reg[209][22]/P0001 ,
		_w13152_,
		_w22652_
	);
	LUT2 #(
		.INIT('h8)
	) name12141 (
		\wishbone_bd_ram_mem2_reg[253][22]/P0001 ,
		_w13100_,
		_w22653_
	);
	LUT2 #(
		.INIT('h8)
	) name12142 (
		\wishbone_bd_ram_mem2_reg[84][22]/P0001 ,
		_w12934_,
		_w22654_
	);
	LUT2 #(
		.INIT('h8)
	) name12143 (
		\wishbone_bd_ram_mem2_reg[8][22]/P0001 ,
		_w12920_,
		_w22655_
	);
	LUT2 #(
		.INIT('h8)
	) name12144 (
		\wishbone_bd_ram_mem2_reg[37][22]/P0001 ,
		_w13102_,
		_w22656_
	);
	LUT2 #(
		.INIT('h8)
	) name12145 (
		\wishbone_bd_ram_mem2_reg[240][22]/P0001 ,
		_w12864_,
		_w22657_
	);
	LUT2 #(
		.INIT('h8)
	) name12146 (
		\wishbone_bd_ram_mem2_reg[29][22]/P0001 ,
		_w12952_,
		_w22658_
	);
	LUT2 #(
		.INIT('h8)
	) name12147 (
		\wishbone_bd_ram_mem2_reg[25][22]/P0001 ,
		_w13108_,
		_w22659_
	);
	LUT2 #(
		.INIT('h8)
	) name12148 (
		\wishbone_bd_ram_mem2_reg[124][22]/P0001 ,
		_w13058_,
		_w22660_
	);
	LUT2 #(
		.INIT('h8)
	) name12149 (
		\wishbone_bd_ram_mem2_reg[94][22]/P0001 ,
		_w13186_,
		_w22661_
	);
	LUT2 #(
		.INIT('h8)
	) name12150 (
		\wishbone_bd_ram_mem2_reg[177][22]/P0001 ,
		_w12996_,
		_w22662_
	);
	LUT2 #(
		.INIT('h8)
	) name12151 (
		\wishbone_bd_ram_mem2_reg[155][22]/P0001 ,
		_w13122_,
		_w22663_
	);
	LUT2 #(
		.INIT('h8)
	) name12152 (
		\wishbone_bd_ram_mem2_reg[48][22]/P0001 ,
		_w12970_,
		_w22664_
	);
	LUT2 #(
		.INIT('h8)
	) name12153 (
		\wishbone_bd_ram_mem2_reg[190][22]/P0001 ,
		_w12858_,
		_w22665_
	);
	LUT2 #(
		.INIT('h8)
	) name12154 (
		\wishbone_bd_ram_mem2_reg[22][22]/P0001 ,
		_w13110_,
		_w22666_
	);
	LUT2 #(
		.INIT('h8)
	) name12155 (
		\wishbone_bd_ram_mem2_reg[89][22]/P0001 ,
		_w12964_,
		_w22667_
	);
	LUT2 #(
		.INIT('h8)
	) name12156 (
		\wishbone_bd_ram_mem2_reg[197][22]/P0001 ,
		_w12834_,
		_w22668_
	);
	LUT2 #(
		.INIT('h8)
	) name12157 (
		\wishbone_bd_ram_mem2_reg[39][22]/P0001 ,
		_w13018_,
		_w22669_
	);
	LUT2 #(
		.INIT('h8)
	) name12158 (
		\wishbone_bd_ram_mem2_reg[142][22]/P0001 ,
		_w12928_,
		_w22670_
	);
	LUT2 #(
		.INIT('h8)
	) name12159 (
		\wishbone_bd_ram_mem2_reg[122][22]/P0001 ,
		_w13130_,
		_w22671_
	);
	LUT2 #(
		.INIT('h8)
	) name12160 (
		\wishbone_bd_ram_mem2_reg[83][22]/P0001 ,
		_w12916_,
		_w22672_
	);
	LUT2 #(
		.INIT('h8)
	) name12161 (
		\wishbone_bd_ram_mem2_reg[69][22]/P0001 ,
		_w12738_,
		_w22673_
	);
	LUT2 #(
		.INIT('h8)
	) name12162 (
		\wishbone_bd_ram_mem2_reg[188][22]/P0001 ,
		_w12948_,
		_w22674_
	);
	LUT2 #(
		.INIT('h8)
	) name12163 (
		\wishbone_bd_ram_mem2_reg[118][22]/P0001 ,
		_w12830_,
		_w22675_
	);
	LUT2 #(
		.INIT('h8)
	) name12164 (
		\wishbone_bd_ram_mem2_reg[161][22]/P0001 ,
		_w12754_,
		_w22676_
	);
	LUT2 #(
		.INIT('h1)
	) name12165 (
		_w22421_,
		_w22422_,
		_w22677_
	);
	LUT2 #(
		.INIT('h1)
	) name12166 (
		_w22423_,
		_w22424_,
		_w22678_
	);
	LUT2 #(
		.INIT('h1)
	) name12167 (
		_w22425_,
		_w22426_,
		_w22679_
	);
	LUT2 #(
		.INIT('h1)
	) name12168 (
		_w22427_,
		_w22428_,
		_w22680_
	);
	LUT2 #(
		.INIT('h1)
	) name12169 (
		_w22429_,
		_w22430_,
		_w22681_
	);
	LUT2 #(
		.INIT('h1)
	) name12170 (
		_w22431_,
		_w22432_,
		_w22682_
	);
	LUT2 #(
		.INIT('h1)
	) name12171 (
		_w22433_,
		_w22434_,
		_w22683_
	);
	LUT2 #(
		.INIT('h1)
	) name12172 (
		_w22435_,
		_w22436_,
		_w22684_
	);
	LUT2 #(
		.INIT('h1)
	) name12173 (
		_w22437_,
		_w22438_,
		_w22685_
	);
	LUT2 #(
		.INIT('h1)
	) name12174 (
		_w22439_,
		_w22440_,
		_w22686_
	);
	LUT2 #(
		.INIT('h1)
	) name12175 (
		_w22441_,
		_w22442_,
		_w22687_
	);
	LUT2 #(
		.INIT('h1)
	) name12176 (
		_w22443_,
		_w22444_,
		_w22688_
	);
	LUT2 #(
		.INIT('h1)
	) name12177 (
		_w22445_,
		_w22446_,
		_w22689_
	);
	LUT2 #(
		.INIT('h1)
	) name12178 (
		_w22447_,
		_w22448_,
		_w22690_
	);
	LUT2 #(
		.INIT('h1)
	) name12179 (
		_w22449_,
		_w22450_,
		_w22691_
	);
	LUT2 #(
		.INIT('h1)
	) name12180 (
		_w22451_,
		_w22452_,
		_w22692_
	);
	LUT2 #(
		.INIT('h1)
	) name12181 (
		_w22453_,
		_w22454_,
		_w22693_
	);
	LUT2 #(
		.INIT('h1)
	) name12182 (
		_w22455_,
		_w22456_,
		_w22694_
	);
	LUT2 #(
		.INIT('h1)
	) name12183 (
		_w22457_,
		_w22458_,
		_w22695_
	);
	LUT2 #(
		.INIT('h1)
	) name12184 (
		_w22459_,
		_w22460_,
		_w22696_
	);
	LUT2 #(
		.INIT('h1)
	) name12185 (
		_w22461_,
		_w22462_,
		_w22697_
	);
	LUT2 #(
		.INIT('h1)
	) name12186 (
		_w22463_,
		_w22464_,
		_w22698_
	);
	LUT2 #(
		.INIT('h1)
	) name12187 (
		_w22465_,
		_w22466_,
		_w22699_
	);
	LUT2 #(
		.INIT('h1)
	) name12188 (
		_w22467_,
		_w22468_,
		_w22700_
	);
	LUT2 #(
		.INIT('h1)
	) name12189 (
		_w22469_,
		_w22470_,
		_w22701_
	);
	LUT2 #(
		.INIT('h1)
	) name12190 (
		_w22471_,
		_w22472_,
		_w22702_
	);
	LUT2 #(
		.INIT('h1)
	) name12191 (
		_w22473_,
		_w22474_,
		_w22703_
	);
	LUT2 #(
		.INIT('h1)
	) name12192 (
		_w22475_,
		_w22476_,
		_w22704_
	);
	LUT2 #(
		.INIT('h1)
	) name12193 (
		_w22477_,
		_w22478_,
		_w22705_
	);
	LUT2 #(
		.INIT('h1)
	) name12194 (
		_w22479_,
		_w22480_,
		_w22706_
	);
	LUT2 #(
		.INIT('h1)
	) name12195 (
		_w22481_,
		_w22482_,
		_w22707_
	);
	LUT2 #(
		.INIT('h1)
	) name12196 (
		_w22483_,
		_w22484_,
		_w22708_
	);
	LUT2 #(
		.INIT('h1)
	) name12197 (
		_w22485_,
		_w22486_,
		_w22709_
	);
	LUT2 #(
		.INIT('h1)
	) name12198 (
		_w22487_,
		_w22488_,
		_w22710_
	);
	LUT2 #(
		.INIT('h1)
	) name12199 (
		_w22489_,
		_w22490_,
		_w22711_
	);
	LUT2 #(
		.INIT('h1)
	) name12200 (
		_w22491_,
		_w22492_,
		_w22712_
	);
	LUT2 #(
		.INIT('h1)
	) name12201 (
		_w22493_,
		_w22494_,
		_w22713_
	);
	LUT2 #(
		.INIT('h1)
	) name12202 (
		_w22495_,
		_w22496_,
		_w22714_
	);
	LUT2 #(
		.INIT('h1)
	) name12203 (
		_w22497_,
		_w22498_,
		_w22715_
	);
	LUT2 #(
		.INIT('h1)
	) name12204 (
		_w22499_,
		_w22500_,
		_w22716_
	);
	LUT2 #(
		.INIT('h1)
	) name12205 (
		_w22501_,
		_w22502_,
		_w22717_
	);
	LUT2 #(
		.INIT('h1)
	) name12206 (
		_w22503_,
		_w22504_,
		_w22718_
	);
	LUT2 #(
		.INIT('h1)
	) name12207 (
		_w22505_,
		_w22506_,
		_w22719_
	);
	LUT2 #(
		.INIT('h1)
	) name12208 (
		_w22507_,
		_w22508_,
		_w22720_
	);
	LUT2 #(
		.INIT('h1)
	) name12209 (
		_w22509_,
		_w22510_,
		_w22721_
	);
	LUT2 #(
		.INIT('h1)
	) name12210 (
		_w22511_,
		_w22512_,
		_w22722_
	);
	LUT2 #(
		.INIT('h1)
	) name12211 (
		_w22513_,
		_w22514_,
		_w22723_
	);
	LUT2 #(
		.INIT('h1)
	) name12212 (
		_w22515_,
		_w22516_,
		_w22724_
	);
	LUT2 #(
		.INIT('h1)
	) name12213 (
		_w22517_,
		_w22518_,
		_w22725_
	);
	LUT2 #(
		.INIT('h1)
	) name12214 (
		_w22519_,
		_w22520_,
		_w22726_
	);
	LUT2 #(
		.INIT('h1)
	) name12215 (
		_w22521_,
		_w22522_,
		_w22727_
	);
	LUT2 #(
		.INIT('h1)
	) name12216 (
		_w22523_,
		_w22524_,
		_w22728_
	);
	LUT2 #(
		.INIT('h1)
	) name12217 (
		_w22525_,
		_w22526_,
		_w22729_
	);
	LUT2 #(
		.INIT('h1)
	) name12218 (
		_w22527_,
		_w22528_,
		_w22730_
	);
	LUT2 #(
		.INIT('h1)
	) name12219 (
		_w22529_,
		_w22530_,
		_w22731_
	);
	LUT2 #(
		.INIT('h1)
	) name12220 (
		_w22531_,
		_w22532_,
		_w22732_
	);
	LUT2 #(
		.INIT('h1)
	) name12221 (
		_w22533_,
		_w22534_,
		_w22733_
	);
	LUT2 #(
		.INIT('h1)
	) name12222 (
		_w22535_,
		_w22536_,
		_w22734_
	);
	LUT2 #(
		.INIT('h1)
	) name12223 (
		_w22537_,
		_w22538_,
		_w22735_
	);
	LUT2 #(
		.INIT('h1)
	) name12224 (
		_w22539_,
		_w22540_,
		_w22736_
	);
	LUT2 #(
		.INIT('h1)
	) name12225 (
		_w22541_,
		_w22542_,
		_w22737_
	);
	LUT2 #(
		.INIT('h1)
	) name12226 (
		_w22543_,
		_w22544_,
		_w22738_
	);
	LUT2 #(
		.INIT('h1)
	) name12227 (
		_w22545_,
		_w22546_,
		_w22739_
	);
	LUT2 #(
		.INIT('h1)
	) name12228 (
		_w22547_,
		_w22548_,
		_w22740_
	);
	LUT2 #(
		.INIT('h1)
	) name12229 (
		_w22549_,
		_w22550_,
		_w22741_
	);
	LUT2 #(
		.INIT('h1)
	) name12230 (
		_w22551_,
		_w22552_,
		_w22742_
	);
	LUT2 #(
		.INIT('h1)
	) name12231 (
		_w22553_,
		_w22554_,
		_w22743_
	);
	LUT2 #(
		.INIT('h1)
	) name12232 (
		_w22555_,
		_w22556_,
		_w22744_
	);
	LUT2 #(
		.INIT('h1)
	) name12233 (
		_w22557_,
		_w22558_,
		_w22745_
	);
	LUT2 #(
		.INIT('h1)
	) name12234 (
		_w22559_,
		_w22560_,
		_w22746_
	);
	LUT2 #(
		.INIT('h1)
	) name12235 (
		_w22561_,
		_w22562_,
		_w22747_
	);
	LUT2 #(
		.INIT('h1)
	) name12236 (
		_w22563_,
		_w22564_,
		_w22748_
	);
	LUT2 #(
		.INIT('h1)
	) name12237 (
		_w22565_,
		_w22566_,
		_w22749_
	);
	LUT2 #(
		.INIT('h1)
	) name12238 (
		_w22567_,
		_w22568_,
		_w22750_
	);
	LUT2 #(
		.INIT('h1)
	) name12239 (
		_w22569_,
		_w22570_,
		_w22751_
	);
	LUT2 #(
		.INIT('h1)
	) name12240 (
		_w22571_,
		_w22572_,
		_w22752_
	);
	LUT2 #(
		.INIT('h1)
	) name12241 (
		_w22573_,
		_w22574_,
		_w22753_
	);
	LUT2 #(
		.INIT('h1)
	) name12242 (
		_w22575_,
		_w22576_,
		_w22754_
	);
	LUT2 #(
		.INIT('h1)
	) name12243 (
		_w22577_,
		_w22578_,
		_w22755_
	);
	LUT2 #(
		.INIT('h1)
	) name12244 (
		_w22579_,
		_w22580_,
		_w22756_
	);
	LUT2 #(
		.INIT('h1)
	) name12245 (
		_w22581_,
		_w22582_,
		_w22757_
	);
	LUT2 #(
		.INIT('h1)
	) name12246 (
		_w22583_,
		_w22584_,
		_w22758_
	);
	LUT2 #(
		.INIT('h1)
	) name12247 (
		_w22585_,
		_w22586_,
		_w22759_
	);
	LUT2 #(
		.INIT('h1)
	) name12248 (
		_w22587_,
		_w22588_,
		_w22760_
	);
	LUT2 #(
		.INIT('h1)
	) name12249 (
		_w22589_,
		_w22590_,
		_w22761_
	);
	LUT2 #(
		.INIT('h1)
	) name12250 (
		_w22591_,
		_w22592_,
		_w22762_
	);
	LUT2 #(
		.INIT('h1)
	) name12251 (
		_w22593_,
		_w22594_,
		_w22763_
	);
	LUT2 #(
		.INIT('h1)
	) name12252 (
		_w22595_,
		_w22596_,
		_w22764_
	);
	LUT2 #(
		.INIT('h1)
	) name12253 (
		_w22597_,
		_w22598_,
		_w22765_
	);
	LUT2 #(
		.INIT('h1)
	) name12254 (
		_w22599_,
		_w22600_,
		_w22766_
	);
	LUT2 #(
		.INIT('h1)
	) name12255 (
		_w22601_,
		_w22602_,
		_w22767_
	);
	LUT2 #(
		.INIT('h1)
	) name12256 (
		_w22603_,
		_w22604_,
		_w22768_
	);
	LUT2 #(
		.INIT('h1)
	) name12257 (
		_w22605_,
		_w22606_,
		_w22769_
	);
	LUT2 #(
		.INIT('h1)
	) name12258 (
		_w22607_,
		_w22608_,
		_w22770_
	);
	LUT2 #(
		.INIT('h1)
	) name12259 (
		_w22609_,
		_w22610_,
		_w22771_
	);
	LUT2 #(
		.INIT('h1)
	) name12260 (
		_w22611_,
		_w22612_,
		_w22772_
	);
	LUT2 #(
		.INIT('h1)
	) name12261 (
		_w22613_,
		_w22614_,
		_w22773_
	);
	LUT2 #(
		.INIT('h1)
	) name12262 (
		_w22615_,
		_w22616_,
		_w22774_
	);
	LUT2 #(
		.INIT('h1)
	) name12263 (
		_w22617_,
		_w22618_,
		_w22775_
	);
	LUT2 #(
		.INIT('h1)
	) name12264 (
		_w22619_,
		_w22620_,
		_w22776_
	);
	LUT2 #(
		.INIT('h1)
	) name12265 (
		_w22621_,
		_w22622_,
		_w22777_
	);
	LUT2 #(
		.INIT('h1)
	) name12266 (
		_w22623_,
		_w22624_,
		_w22778_
	);
	LUT2 #(
		.INIT('h1)
	) name12267 (
		_w22625_,
		_w22626_,
		_w22779_
	);
	LUT2 #(
		.INIT('h1)
	) name12268 (
		_w22627_,
		_w22628_,
		_w22780_
	);
	LUT2 #(
		.INIT('h1)
	) name12269 (
		_w22629_,
		_w22630_,
		_w22781_
	);
	LUT2 #(
		.INIT('h1)
	) name12270 (
		_w22631_,
		_w22632_,
		_w22782_
	);
	LUT2 #(
		.INIT('h1)
	) name12271 (
		_w22633_,
		_w22634_,
		_w22783_
	);
	LUT2 #(
		.INIT('h1)
	) name12272 (
		_w22635_,
		_w22636_,
		_w22784_
	);
	LUT2 #(
		.INIT('h1)
	) name12273 (
		_w22637_,
		_w22638_,
		_w22785_
	);
	LUT2 #(
		.INIT('h1)
	) name12274 (
		_w22639_,
		_w22640_,
		_w22786_
	);
	LUT2 #(
		.INIT('h1)
	) name12275 (
		_w22641_,
		_w22642_,
		_w22787_
	);
	LUT2 #(
		.INIT('h1)
	) name12276 (
		_w22643_,
		_w22644_,
		_w22788_
	);
	LUT2 #(
		.INIT('h1)
	) name12277 (
		_w22645_,
		_w22646_,
		_w22789_
	);
	LUT2 #(
		.INIT('h1)
	) name12278 (
		_w22647_,
		_w22648_,
		_w22790_
	);
	LUT2 #(
		.INIT('h1)
	) name12279 (
		_w22649_,
		_w22650_,
		_w22791_
	);
	LUT2 #(
		.INIT('h1)
	) name12280 (
		_w22651_,
		_w22652_,
		_w22792_
	);
	LUT2 #(
		.INIT('h1)
	) name12281 (
		_w22653_,
		_w22654_,
		_w22793_
	);
	LUT2 #(
		.INIT('h1)
	) name12282 (
		_w22655_,
		_w22656_,
		_w22794_
	);
	LUT2 #(
		.INIT('h1)
	) name12283 (
		_w22657_,
		_w22658_,
		_w22795_
	);
	LUT2 #(
		.INIT('h1)
	) name12284 (
		_w22659_,
		_w22660_,
		_w22796_
	);
	LUT2 #(
		.INIT('h1)
	) name12285 (
		_w22661_,
		_w22662_,
		_w22797_
	);
	LUT2 #(
		.INIT('h1)
	) name12286 (
		_w22663_,
		_w22664_,
		_w22798_
	);
	LUT2 #(
		.INIT('h1)
	) name12287 (
		_w22665_,
		_w22666_,
		_w22799_
	);
	LUT2 #(
		.INIT('h1)
	) name12288 (
		_w22667_,
		_w22668_,
		_w22800_
	);
	LUT2 #(
		.INIT('h1)
	) name12289 (
		_w22669_,
		_w22670_,
		_w22801_
	);
	LUT2 #(
		.INIT('h1)
	) name12290 (
		_w22671_,
		_w22672_,
		_w22802_
	);
	LUT2 #(
		.INIT('h1)
	) name12291 (
		_w22673_,
		_w22674_,
		_w22803_
	);
	LUT2 #(
		.INIT('h1)
	) name12292 (
		_w22675_,
		_w22676_,
		_w22804_
	);
	LUT2 #(
		.INIT('h8)
	) name12293 (
		_w22803_,
		_w22804_,
		_w22805_
	);
	LUT2 #(
		.INIT('h8)
	) name12294 (
		_w22801_,
		_w22802_,
		_w22806_
	);
	LUT2 #(
		.INIT('h8)
	) name12295 (
		_w22799_,
		_w22800_,
		_w22807_
	);
	LUT2 #(
		.INIT('h8)
	) name12296 (
		_w22797_,
		_w22798_,
		_w22808_
	);
	LUT2 #(
		.INIT('h8)
	) name12297 (
		_w22795_,
		_w22796_,
		_w22809_
	);
	LUT2 #(
		.INIT('h8)
	) name12298 (
		_w22793_,
		_w22794_,
		_w22810_
	);
	LUT2 #(
		.INIT('h8)
	) name12299 (
		_w22791_,
		_w22792_,
		_w22811_
	);
	LUT2 #(
		.INIT('h8)
	) name12300 (
		_w22789_,
		_w22790_,
		_w22812_
	);
	LUT2 #(
		.INIT('h8)
	) name12301 (
		_w22787_,
		_w22788_,
		_w22813_
	);
	LUT2 #(
		.INIT('h8)
	) name12302 (
		_w22785_,
		_w22786_,
		_w22814_
	);
	LUT2 #(
		.INIT('h8)
	) name12303 (
		_w22783_,
		_w22784_,
		_w22815_
	);
	LUT2 #(
		.INIT('h8)
	) name12304 (
		_w22781_,
		_w22782_,
		_w22816_
	);
	LUT2 #(
		.INIT('h8)
	) name12305 (
		_w22779_,
		_w22780_,
		_w22817_
	);
	LUT2 #(
		.INIT('h8)
	) name12306 (
		_w22777_,
		_w22778_,
		_w22818_
	);
	LUT2 #(
		.INIT('h8)
	) name12307 (
		_w22775_,
		_w22776_,
		_w22819_
	);
	LUT2 #(
		.INIT('h8)
	) name12308 (
		_w22773_,
		_w22774_,
		_w22820_
	);
	LUT2 #(
		.INIT('h8)
	) name12309 (
		_w22771_,
		_w22772_,
		_w22821_
	);
	LUT2 #(
		.INIT('h8)
	) name12310 (
		_w22769_,
		_w22770_,
		_w22822_
	);
	LUT2 #(
		.INIT('h8)
	) name12311 (
		_w22767_,
		_w22768_,
		_w22823_
	);
	LUT2 #(
		.INIT('h8)
	) name12312 (
		_w22765_,
		_w22766_,
		_w22824_
	);
	LUT2 #(
		.INIT('h8)
	) name12313 (
		_w22763_,
		_w22764_,
		_w22825_
	);
	LUT2 #(
		.INIT('h8)
	) name12314 (
		_w22761_,
		_w22762_,
		_w22826_
	);
	LUT2 #(
		.INIT('h8)
	) name12315 (
		_w22759_,
		_w22760_,
		_w22827_
	);
	LUT2 #(
		.INIT('h8)
	) name12316 (
		_w22757_,
		_w22758_,
		_w22828_
	);
	LUT2 #(
		.INIT('h8)
	) name12317 (
		_w22755_,
		_w22756_,
		_w22829_
	);
	LUT2 #(
		.INIT('h8)
	) name12318 (
		_w22753_,
		_w22754_,
		_w22830_
	);
	LUT2 #(
		.INIT('h8)
	) name12319 (
		_w22751_,
		_w22752_,
		_w22831_
	);
	LUT2 #(
		.INIT('h8)
	) name12320 (
		_w22749_,
		_w22750_,
		_w22832_
	);
	LUT2 #(
		.INIT('h8)
	) name12321 (
		_w22747_,
		_w22748_,
		_w22833_
	);
	LUT2 #(
		.INIT('h8)
	) name12322 (
		_w22745_,
		_w22746_,
		_w22834_
	);
	LUT2 #(
		.INIT('h8)
	) name12323 (
		_w22743_,
		_w22744_,
		_w22835_
	);
	LUT2 #(
		.INIT('h8)
	) name12324 (
		_w22741_,
		_w22742_,
		_w22836_
	);
	LUT2 #(
		.INIT('h8)
	) name12325 (
		_w22739_,
		_w22740_,
		_w22837_
	);
	LUT2 #(
		.INIT('h8)
	) name12326 (
		_w22737_,
		_w22738_,
		_w22838_
	);
	LUT2 #(
		.INIT('h8)
	) name12327 (
		_w22735_,
		_w22736_,
		_w22839_
	);
	LUT2 #(
		.INIT('h8)
	) name12328 (
		_w22733_,
		_w22734_,
		_w22840_
	);
	LUT2 #(
		.INIT('h8)
	) name12329 (
		_w22731_,
		_w22732_,
		_w22841_
	);
	LUT2 #(
		.INIT('h8)
	) name12330 (
		_w22729_,
		_w22730_,
		_w22842_
	);
	LUT2 #(
		.INIT('h8)
	) name12331 (
		_w22727_,
		_w22728_,
		_w22843_
	);
	LUT2 #(
		.INIT('h8)
	) name12332 (
		_w22725_,
		_w22726_,
		_w22844_
	);
	LUT2 #(
		.INIT('h8)
	) name12333 (
		_w22723_,
		_w22724_,
		_w22845_
	);
	LUT2 #(
		.INIT('h8)
	) name12334 (
		_w22721_,
		_w22722_,
		_w22846_
	);
	LUT2 #(
		.INIT('h8)
	) name12335 (
		_w22719_,
		_w22720_,
		_w22847_
	);
	LUT2 #(
		.INIT('h8)
	) name12336 (
		_w22717_,
		_w22718_,
		_w22848_
	);
	LUT2 #(
		.INIT('h8)
	) name12337 (
		_w22715_,
		_w22716_,
		_w22849_
	);
	LUT2 #(
		.INIT('h8)
	) name12338 (
		_w22713_,
		_w22714_,
		_w22850_
	);
	LUT2 #(
		.INIT('h8)
	) name12339 (
		_w22711_,
		_w22712_,
		_w22851_
	);
	LUT2 #(
		.INIT('h8)
	) name12340 (
		_w22709_,
		_w22710_,
		_w22852_
	);
	LUT2 #(
		.INIT('h8)
	) name12341 (
		_w22707_,
		_w22708_,
		_w22853_
	);
	LUT2 #(
		.INIT('h8)
	) name12342 (
		_w22705_,
		_w22706_,
		_w22854_
	);
	LUT2 #(
		.INIT('h8)
	) name12343 (
		_w22703_,
		_w22704_,
		_w22855_
	);
	LUT2 #(
		.INIT('h8)
	) name12344 (
		_w22701_,
		_w22702_,
		_w22856_
	);
	LUT2 #(
		.INIT('h8)
	) name12345 (
		_w22699_,
		_w22700_,
		_w22857_
	);
	LUT2 #(
		.INIT('h8)
	) name12346 (
		_w22697_,
		_w22698_,
		_w22858_
	);
	LUT2 #(
		.INIT('h8)
	) name12347 (
		_w22695_,
		_w22696_,
		_w22859_
	);
	LUT2 #(
		.INIT('h8)
	) name12348 (
		_w22693_,
		_w22694_,
		_w22860_
	);
	LUT2 #(
		.INIT('h8)
	) name12349 (
		_w22691_,
		_w22692_,
		_w22861_
	);
	LUT2 #(
		.INIT('h8)
	) name12350 (
		_w22689_,
		_w22690_,
		_w22862_
	);
	LUT2 #(
		.INIT('h8)
	) name12351 (
		_w22687_,
		_w22688_,
		_w22863_
	);
	LUT2 #(
		.INIT('h8)
	) name12352 (
		_w22685_,
		_w22686_,
		_w22864_
	);
	LUT2 #(
		.INIT('h8)
	) name12353 (
		_w22683_,
		_w22684_,
		_w22865_
	);
	LUT2 #(
		.INIT('h8)
	) name12354 (
		_w22681_,
		_w22682_,
		_w22866_
	);
	LUT2 #(
		.INIT('h8)
	) name12355 (
		_w22679_,
		_w22680_,
		_w22867_
	);
	LUT2 #(
		.INIT('h8)
	) name12356 (
		_w22677_,
		_w22678_,
		_w22868_
	);
	LUT2 #(
		.INIT('h8)
	) name12357 (
		_w22867_,
		_w22868_,
		_w22869_
	);
	LUT2 #(
		.INIT('h8)
	) name12358 (
		_w22865_,
		_w22866_,
		_w22870_
	);
	LUT2 #(
		.INIT('h8)
	) name12359 (
		_w22863_,
		_w22864_,
		_w22871_
	);
	LUT2 #(
		.INIT('h8)
	) name12360 (
		_w22861_,
		_w22862_,
		_w22872_
	);
	LUT2 #(
		.INIT('h8)
	) name12361 (
		_w22859_,
		_w22860_,
		_w22873_
	);
	LUT2 #(
		.INIT('h8)
	) name12362 (
		_w22857_,
		_w22858_,
		_w22874_
	);
	LUT2 #(
		.INIT('h8)
	) name12363 (
		_w22855_,
		_w22856_,
		_w22875_
	);
	LUT2 #(
		.INIT('h8)
	) name12364 (
		_w22853_,
		_w22854_,
		_w22876_
	);
	LUT2 #(
		.INIT('h8)
	) name12365 (
		_w22851_,
		_w22852_,
		_w22877_
	);
	LUT2 #(
		.INIT('h8)
	) name12366 (
		_w22849_,
		_w22850_,
		_w22878_
	);
	LUT2 #(
		.INIT('h8)
	) name12367 (
		_w22847_,
		_w22848_,
		_w22879_
	);
	LUT2 #(
		.INIT('h8)
	) name12368 (
		_w22845_,
		_w22846_,
		_w22880_
	);
	LUT2 #(
		.INIT('h8)
	) name12369 (
		_w22843_,
		_w22844_,
		_w22881_
	);
	LUT2 #(
		.INIT('h8)
	) name12370 (
		_w22841_,
		_w22842_,
		_w22882_
	);
	LUT2 #(
		.INIT('h8)
	) name12371 (
		_w22839_,
		_w22840_,
		_w22883_
	);
	LUT2 #(
		.INIT('h8)
	) name12372 (
		_w22837_,
		_w22838_,
		_w22884_
	);
	LUT2 #(
		.INIT('h8)
	) name12373 (
		_w22835_,
		_w22836_,
		_w22885_
	);
	LUT2 #(
		.INIT('h8)
	) name12374 (
		_w22833_,
		_w22834_,
		_w22886_
	);
	LUT2 #(
		.INIT('h8)
	) name12375 (
		_w22831_,
		_w22832_,
		_w22887_
	);
	LUT2 #(
		.INIT('h8)
	) name12376 (
		_w22829_,
		_w22830_,
		_w22888_
	);
	LUT2 #(
		.INIT('h8)
	) name12377 (
		_w22827_,
		_w22828_,
		_w22889_
	);
	LUT2 #(
		.INIT('h8)
	) name12378 (
		_w22825_,
		_w22826_,
		_w22890_
	);
	LUT2 #(
		.INIT('h8)
	) name12379 (
		_w22823_,
		_w22824_,
		_w22891_
	);
	LUT2 #(
		.INIT('h8)
	) name12380 (
		_w22821_,
		_w22822_,
		_w22892_
	);
	LUT2 #(
		.INIT('h8)
	) name12381 (
		_w22819_,
		_w22820_,
		_w22893_
	);
	LUT2 #(
		.INIT('h8)
	) name12382 (
		_w22817_,
		_w22818_,
		_w22894_
	);
	LUT2 #(
		.INIT('h8)
	) name12383 (
		_w22815_,
		_w22816_,
		_w22895_
	);
	LUT2 #(
		.INIT('h8)
	) name12384 (
		_w22813_,
		_w22814_,
		_w22896_
	);
	LUT2 #(
		.INIT('h8)
	) name12385 (
		_w22811_,
		_w22812_,
		_w22897_
	);
	LUT2 #(
		.INIT('h8)
	) name12386 (
		_w22809_,
		_w22810_,
		_w22898_
	);
	LUT2 #(
		.INIT('h8)
	) name12387 (
		_w22807_,
		_w22808_,
		_w22899_
	);
	LUT2 #(
		.INIT('h8)
	) name12388 (
		_w22805_,
		_w22806_,
		_w22900_
	);
	LUT2 #(
		.INIT('h8)
	) name12389 (
		_w22899_,
		_w22900_,
		_w22901_
	);
	LUT2 #(
		.INIT('h8)
	) name12390 (
		_w22897_,
		_w22898_,
		_w22902_
	);
	LUT2 #(
		.INIT('h8)
	) name12391 (
		_w22895_,
		_w22896_,
		_w22903_
	);
	LUT2 #(
		.INIT('h8)
	) name12392 (
		_w22893_,
		_w22894_,
		_w22904_
	);
	LUT2 #(
		.INIT('h8)
	) name12393 (
		_w22891_,
		_w22892_,
		_w22905_
	);
	LUT2 #(
		.INIT('h8)
	) name12394 (
		_w22889_,
		_w22890_,
		_w22906_
	);
	LUT2 #(
		.INIT('h8)
	) name12395 (
		_w22887_,
		_w22888_,
		_w22907_
	);
	LUT2 #(
		.INIT('h8)
	) name12396 (
		_w22885_,
		_w22886_,
		_w22908_
	);
	LUT2 #(
		.INIT('h8)
	) name12397 (
		_w22883_,
		_w22884_,
		_w22909_
	);
	LUT2 #(
		.INIT('h8)
	) name12398 (
		_w22881_,
		_w22882_,
		_w22910_
	);
	LUT2 #(
		.INIT('h8)
	) name12399 (
		_w22879_,
		_w22880_,
		_w22911_
	);
	LUT2 #(
		.INIT('h8)
	) name12400 (
		_w22877_,
		_w22878_,
		_w22912_
	);
	LUT2 #(
		.INIT('h8)
	) name12401 (
		_w22875_,
		_w22876_,
		_w22913_
	);
	LUT2 #(
		.INIT('h8)
	) name12402 (
		_w22873_,
		_w22874_,
		_w22914_
	);
	LUT2 #(
		.INIT('h8)
	) name12403 (
		_w22871_,
		_w22872_,
		_w22915_
	);
	LUT2 #(
		.INIT('h8)
	) name12404 (
		_w22869_,
		_w22870_,
		_w22916_
	);
	LUT2 #(
		.INIT('h8)
	) name12405 (
		_w22915_,
		_w22916_,
		_w22917_
	);
	LUT2 #(
		.INIT('h8)
	) name12406 (
		_w22913_,
		_w22914_,
		_w22918_
	);
	LUT2 #(
		.INIT('h8)
	) name12407 (
		_w22911_,
		_w22912_,
		_w22919_
	);
	LUT2 #(
		.INIT('h8)
	) name12408 (
		_w22909_,
		_w22910_,
		_w22920_
	);
	LUT2 #(
		.INIT('h8)
	) name12409 (
		_w22907_,
		_w22908_,
		_w22921_
	);
	LUT2 #(
		.INIT('h8)
	) name12410 (
		_w22905_,
		_w22906_,
		_w22922_
	);
	LUT2 #(
		.INIT('h8)
	) name12411 (
		_w22903_,
		_w22904_,
		_w22923_
	);
	LUT2 #(
		.INIT('h8)
	) name12412 (
		_w22901_,
		_w22902_,
		_w22924_
	);
	LUT2 #(
		.INIT('h8)
	) name12413 (
		_w22923_,
		_w22924_,
		_w22925_
	);
	LUT2 #(
		.INIT('h8)
	) name12414 (
		_w22921_,
		_w22922_,
		_w22926_
	);
	LUT2 #(
		.INIT('h8)
	) name12415 (
		_w22919_,
		_w22920_,
		_w22927_
	);
	LUT2 #(
		.INIT('h8)
	) name12416 (
		_w22917_,
		_w22918_,
		_w22928_
	);
	LUT2 #(
		.INIT('h8)
	) name12417 (
		_w22927_,
		_w22928_,
		_w22929_
	);
	LUT2 #(
		.INIT('h8)
	) name12418 (
		_w22925_,
		_w22926_,
		_w22930_
	);
	LUT2 #(
		.INIT('h8)
	) name12419 (
		_w22929_,
		_w22930_,
		_w22931_
	);
	LUT2 #(
		.INIT('h1)
	) name12420 (
		wb_rst_i_pad,
		_w22931_,
		_w22932_
	);
	LUT2 #(
		.INIT('h8)
	) name12421 (
		_w12656_,
		_w22932_,
		_w22933_
	);
	LUT2 #(
		.INIT('h1)
	) name12422 (
		_w22420_,
		_w22933_,
		_w22934_
	);
	LUT2 #(
		.INIT('h2)
	) name12423 (
		\wishbone_LatchedTxLength_reg[9]/NET0131 ,
		_w12656_,
		_w22935_
	);
	LUT2 #(
		.INIT('h1)
	) name12424 (
		_w17811_,
		_w22935_,
		_w22936_
	);
	LUT2 #(
		.INIT('h8)
	) name12425 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w22937_
	);
	LUT2 #(
		.INIT('h1)
	) name12426 (
		\wb_sel_i[0]_pad ,
		\wb_sel_i[1]_pad ,
		_w22938_
	);
	LUT2 #(
		.INIT('h1)
	) name12427 (
		\wb_sel_i[2]_pad ,
		\wb_sel_i[3]_pad ,
		_w22939_
	);
	LUT2 #(
		.INIT('h8)
	) name12428 (
		_w22938_,
		_w22939_,
		_w22940_
	);
	LUT2 #(
		.INIT('h1)
	) name12429 (
		\wb_adr_i[11]_pad ,
		_w22940_,
		_w22941_
	);
	LUT2 #(
		.INIT('h8)
	) name12430 (
		_w22937_,
		_w22941_,
		_w22942_
	);
	LUT2 #(
		.INIT('h4)
	) name12431 (
		\wb_adr_i[10]_pad ,
		_w22942_,
		_w22943_
	);
	LUT2 #(
		.INIT('h4)
	) name12432 (
		wb_we_i_pad,
		_w22943_,
		_w22944_
	);
	LUT2 #(
		.INIT('h1)
	) name12433 (
		_w21900_,
		_w22944_,
		_w22945_
	);
	LUT2 #(
		.INIT('h1)
	) name12434 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w22946_
	);
	LUT2 #(
		.INIT('h8)
	) name12435 (
		\wb_adr_i[3]_pad ,
		_w22946_,
		_w22947_
	);
	LUT2 #(
		.INIT('h1)
	) name12436 (
		\wb_adr_i[7]_pad ,
		\wb_adr_i[9]_pad ,
		_w22948_
	);
	LUT2 #(
		.INIT('h8)
	) name12437 (
		\wb_adr_i[6]_pad ,
		_w22948_,
		_w22949_
	);
	LUT2 #(
		.INIT('h1)
	) name12438 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[8]_pad ,
		_w22950_
	);
	LUT2 #(
		.INIT('h8)
	) name12439 (
		_w22949_,
		_w22950_,
		_w22951_
	);
	LUT2 #(
		.INIT('h8)
	) name12440 (
		_w22947_,
		_w22951_,
		_w22952_
	);
	LUT2 #(
		.INIT('h8)
	) name12441 (
		\ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 ,
		_w22952_,
		_w22953_
	);
	LUT2 #(
		.INIT('h2)
	) name12442 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[8]_pad ,
		_w22954_
	);
	LUT2 #(
		.INIT('h8)
	) name12443 (
		_w22949_,
		_w22954_,
		_w22955_
	);
	LUT2 #(
		.INIT('h8)
	) name12444 (
		_w22947_,
		_w22955_,
		_w22956_
	);
	LUT2 #(
		.INIT('h8)
	) name12445 (
		\ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 ,
		_w22956_,
		_w22957_
	);
	LUT2 #(
		.INIT('h4)
	) name12446 (
		\wb_adr_i[3]_pad ,
		_w22946_,
		_w22958_
	);
	LUT2 #(
		.INIT('h8)
	) name12447 (
		_w22951_,
		_w22958_,
		_w22959_
	);
	LUT2 #(
		.INIT('h8)
	) name12448 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		_w22959_,
		_w22960_
	);
	LUT2 #(
		.INIT('h4)
	) name12449 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w22961_
	);
	LUT2 #(
		.INIT('h4)
	) name12450 (
		\wb_adr_i[8]_pad ,
		_w22948_,
		_w22962_
	);
	LUT2 #(
		.INIT('h4)
	) name12451 (
		\wb_adr_i[6]_pad ,
		_w22962_,
		_w22963_
	);
	LUT2 #(
		.INIT('h4)
	) name12452 (
		\wb_adr_i[5]_pad ,
		_w22963_,
		_w22964_
	);
	LUT2 #(
		.INIT('h8)
	) name12453 (
		_w22961_,
		_w22964_,
		_w22965_
	);
	LUT2 #(
		.INIT('h8)
	) name12454 (
		\wb_adr_i[4]_pad ,
		_w22965_,
		_w22966_
	);
	LUT2 #(
		.INIT('h8)
	) name12455 (
		\ethreg1_PACKETLEN_2_DataOut_reg[5]/NET0131 ,
		_w22966_,
		_w22967_
	);
	LUT2 #(
		.INIT('h1)
	) name12456 (
		_w22953_,
		_w22957_,
		_w22968_
	);
	LUT2 #(
		.INIT('h4)
	) name12457 (
		_w22960_,
		_w22968_,
		_w22969_
	);
	LUT2 #(
		.INIT('h8)
	) name12458 (
		_w22944_,
		_w22969_,
		_w22970_
	);
	LUT2 #(
		.INIT('h4)
	) name12459 (
		_w22967_,
		_w22970_,
		_w22971_
	);
	LUT2 #(
		.INIT('h1)
	) name12460 (
		_w22945_,
		_w22971_,
		_w22972_
	);
	LUT2 #(
		.INIT('h1)
	) name12461 (
		_w22932_,
		_w22944_,
		_w22973_
	);
	LUT2 #(
		.INIT('h8)
	) name12462 (
		\ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 ,
		_w22952_,
		_w22974_
	);
	LUT2 #(
		.INIT('h8)
	) name12463 (
		\ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 ,
		_w22956_,
		_w22975_
	);
	LUT2 #(
		.INIT('h8)
	) name12464 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		_w22959_,
		_w22976_
	);
	LUT2 #(
		.INIT('h8)
	) name12465 (
		\ethreg1_PACKETLEN_2_DataOut_reg[6]/NET0131 ,
		_w22966_,
		_w22977_
	);
	LUT2 #(
		.INIT('h1)
	) name12466 (
		_w22974_,
		_w22975_,
		_w22978_
	);
	LUT2 #(
		.INIT('h4)
	) name12467 (
		_w22976_,
		_w22978_,
		_w22979_
	);
	LUT2 #(
		.INIT('h8)
	) name12468 (
		_w22944_,
		_w22979_,
		_w22980_
	);
	LUT2 #(
		.INIT('h4)
	) name12469 (
		_w22977_,
		_w22980_,
		_w22981_
	);
	LUT2 #(
		.INIT('h1)
	) name12470 (
		_w22973_,
		_w22981_,
		_w22982_
	);
	LUT2 #(
		.INIT('h8)
	) name12471 (
		\wishbone_bd_ram_mem1_reg[17][12]/P0001 ,
		_w12848_,
		_w22983_
	);
	LUT2 #(
		.INIT('h8)
	) name12472 (
		\wishbone_bd_ram_mem1_reg[95][12]/P0001 ,
		_w12844_,
		_w22984_
	);
	LUT2 #(
		.INIT('h8)
	) name12473 (
		\wishbone_bd_ram_mem1_reg[189][12]/P0001 ,
		_w13042_,
		_w22985_
	);
	LUT2 #(
		.INIT('h8)
	) name12474 (
		\wishbone_bd_ram_mem1_reg[145][12]/P0001 ,
		_w13106_,
		_w22986_
	);
	LUT2 #(
		.INIT('h8)
	) name12475 (
		\wishbone_bd_ram_mem1_reg[236][12]/P0001 ,
		_w12731_,
		_w22987_
	);
	LUT2 #(
		.INIT('h8)
	) name12476 (
		\wishbone_bd_ram_mem1_reg[86][12]/P0001 ,
		_w12735_,
		_w22988_
	);
	LUT2 #(
		.INIT('h8)
	) name12477 (
		\wishbone_bd_ram_mem1_reg[161][12]/P0001 ,
		_w12754_,
		_w22989_
	);
	LUT2 #(
		.INIT('h8)
	) name12478 (
		\wishbone_bd_ram_mem1_reg[117][12]/P0001 ,
		_w12715_,
		_w22990_
	);
	LUT2 #(
		.INIT('h8)
	) name12479 (
		\wishbone_bd_ram_mem1_reg[211][12]/P0001 ,
		_w13166_,
		_w22991_
	);
	LUT2 #(
		.INIT('h8)
	) name12480 (
		\wishbone_bd_ram_mem1_reg[194][12]/P0001 ,
		_w12772_,
		_w22992_
	);
	LUT2 #(
		.INIT('h8)
	) name12481 (
		\wishbone_bd_ram_mem1_reg[166][12]/P0001 ,
		_w13040_,
		_w22993_
	);
	LUT2 #(
		.INIT('h8)
	) name12482 (
		\wishbone_bd_ram_mem1_reg[208][12]/P0001 ,
		_w13032_,
		_w22994_
	);
	LUT2 #(
		.INIT('h8)
	) name12483 (
		\wishbone_bd_ram_mem1_reg[13][12]/P0001 ,
		_w13178_,
		_w22995_
	);
	LUT2 #(
		.INIT('h8)
	) name12484 (
		\wishbone_bd_ram_mem1_reg[83][12]/P0001 ,
		_w12916_,
		_w22996_
	);
	LUT2 #(
		.INIT('h8)
	) name12485 (
		\wishbone_bd_ram_mem1_reg[125][12]/P0001 ,
		_w12956_,
		_w22997_
	);
	LUT2 #(
		.INIT('h8)
	) name12486 (
		\wishbone_bd_ram_mem1_reg[22][12]/P0001 ,
		_w13110_,
		_w22998_
	);
	LUT2 #(
		.INIT('h8)
	) name12487 (
		\wishbone_bd_ram_mem1_reg[212][12]/P0001 ,
		_w12796_,
		_w22999_
	);
	LUT2 #(
		.INIT('h8)
	) name12488 (
		\wishbone_bd_ram_mem1_reg[59][12]/P0001 ,
		_w12780_,
		_w23000_
	);
	LUT2 #(
		.INIT('h8)
	) name12489 (
		\wishbone_bd_ram_mem1_reg[85][12]/P0001 ,
		_w13216_,
		_w23001_
	);
	LUT2 #(
		.INIT('h8)
	) name12490 (
		\wishbone_bd_ram_mem1_reg[90][12]/P0001 ,
		_w12978_,
		_w23002_
	);
	LUT2 #(
		.INIT('h8)
	) name12491 (
		\wishbone_bd_ram_mem1_reg[33][12]/P0001 ,
		_w12980_,
		_w23003_
	);
	LUT2 #(
		.INIT('h8)
	) name12492 (
		\wishbone_bd_ram_mem1_reg[238][12]/P0001 ,
		_w13160_,
		_w23004_
	);
	LUT2 #(
		.INIT('h8)
	) name12493 (
		\wishbone_bd_ram_mem1_reg[153][12]/P0001 ,
		_w12890_,
		_w23005_
	);
	LUT2 #(
		.INIT('h8)
	) name12494 (
		\wishbone_bd_ram_mem1_reg[24][12]/P0001 ,
		_w13084_,
		_w23006_
	);
	LUT2 #(
		.INIT('h8)
	) name12495 (
		\wishbone_bd_ram_mem1_reg[165][12]/P0001 ,
		_w13044_,
		_w23007_
	);
	LUT2 #(
		.INIT('h8)
	) name12496 (
		\wishbone_bd_ram_mem1_reg[146][12]/P0001 ,
		_w13060_,
		_w23008_
	);
	LUT2 #(
		.INIT('h8)
	) name12497 (
		\wishbone_bd_ram_mem1_reg[128][12]/P0001 ,
		_w12793_,
		_w23009_
	);
	LUT2 #(
		.INIT('h8)
	) name12498 (
		\wishbone_bd_ram_mem1_reg[28][12]/P0001 ,
		_w13170_,
		_w23010_
	);
	LUT2 #(
		.INIT('h8)
	) name12499 (
		\wishbone_bd_ram_mem1_reg[139][12]/P0001 ,
		_w12814_,
		_w23011_
	);
	LUT2 #(
		.INIT('h8)
	) name12500 (
		\wishbone_bd_ram_mem1_reg[97][12]/P0001 ,
		_w13096_,
		_w23012_
	);
	LUT2 #(
		.INIT('h8)
	) name12501 (
		\wishbone_bd_ram_mem1_reg[232][12]/P0001 ,
		_w12758_,
		_w23013_
	);
	LUT2 #(
		.INIT('h8)
	) name12502 (
		\wishbone_bd_ram_mem1_reg[223][12]/P0001 ,
		_w12838_,
		_w23014_
	);
	LUT2 #(
		.INIT('h8)
	) name12503 (
		\wishbone_bd_ram_mem1_reg[250][12]/P0001 ,
		_w13128_,
		_w23015_
	);
	LUT2 #(
		.INIT('h8)
	) name12504 (
		\wishbone_bd_ram_mem1_reg[23][12]/P0001 ,
		_w13008_,
		_w23016_
	);
	LUT2 #(
		.INIT('h8)
	) name12505 (
		\wishbone_bd_ram_mem1_reg[66][12]/P0001 ,
		_w12824_,
		_w23017_
	);
	LUT2 #(
		.INIT('h8)
	) name12506 (
		\wishbone_bd_ram_mem1_reg[116][12]/P0001 ,
		_w12998_,
		_w23018_
	);
	LUT2 #(
		.INIT('h8)
	) name12507 (
		\wishbone_bd_ram_mem1_reg[20][12]/P0001 ,
		_w13174_,
		_w23019_
	);
	LUT2 #(
		.INIT('h8)
	) name12508 (
		\wishbone_bd_ram_mem1_reg[123][12]/P0001 ,
		_w13114_,
		_w23020_
	);
	LUT2 #(
		.INIT('h8)
	) name12509 (
		\wishbone_bd_ram_mem1_reg[63][12]/P0001 ,
		_w12850_,
		_w23021_
	);
	LUT2 #(
		.INIT('h8)
	) name12510 (
		\wishbone_bd_ram_mem1_reg[196][12]/P0001 ,
		_w13090_,
		_w23022_
	);
	LUT2 #(
		.INIT('h8)
	) name12511 (
		\wishbone_bd_ram_mem1_reg[38][12]/P0001 ,
		_w13182_,
		_w23023_
	);
	LUT2 #(
		.INIT('h8)
	) name12512 (
		\wishbone_bd_ram_mem1_reg[202][12]/P0001 ,
		_w12870_,
		_w23024_
	);
	LUT2 #(
		.INIT('h8)
	) name12513 (
		\wishbone_bd_ram_mem1_reg[131][12]/P0001 ,
		_w12852_,
		_w23025_
	);
	LUT2 #(
		.INIT('h8)
	) name12514 (
		\wishbone_bd_ram_mem1_reg[29][12]/P0001 ,
		_w12952_,
		_w23026_
	);
	LUT2 #(
		.INIT('h8)
	) name12515 (
		\wishbone_bd_ram_mem1_reg[235][12]/P0001 ,
		_w12696_,
		_w23027_
	);
	LUT2 #(
		.INIT('h8)
	) name12516 (
		\wishbone_bd_ram_mem1_reg[124][12]/P0001 ,
		_w13058_,
		_w23028_
	);
	LUT2 #(
		.INIT('h8)
	) name12517 (
		\wishbone_bd_ram_mem1_reg[110][12]/P0001 ,
		_w13046_,
		_w23029_
	);
	LUT2 #(
		.INIT('h8)
	) name12518 (
		\wishbone_bd_ram_mem1_reg[181][12]/P0001 ,
		_w12828_,
		_w23030_
	);
	LUT2 #(
		.INIT('h8)
	) name12519 (
		\wishbone_bd_ram_mem1_reg[141][12]/P0001 ,
		_w13004_,
		_w23031_
	);
	LUT2 #(
		.INIT('h8)
	) name12520 (
		\wishbone_bd_ram_mem1_reg[169][12]/P0001 ,
		_w12722_,
		_w23032_
	);
	LUT2 #(
		.INIT('h8)
	) name12521 (
		\wishbone_bd_ram_mem1_reg[4][12]/P0001 ,
		_w12666_,
		_w23033_
	);
	LUT2 #(
		.INIT('h8)
	) name12522 (
		\wishbone_bd_ram_mem1_reg[78][12]/P0001 ,
		_w12874_,
		_w23034_
	);
	LUT2 #(
		.INIT('h8)
	) name12523 (
		\wishbone_bd_ram_mem1_reg[76][12]/P0001 ,
		_w13184_,
		_w23035_
	);
	LUT2 #(
		.INIT('h8)
	) name12524 (
		\wishbone_bd_ram_mem1_reg[233][12]/P0001 ,
		_w12836_,
		_w23036_
	);
	LUT2 #(
		.INIT('h8)
	) name12525 (
		\wishbone_bd_ram_mem1_reg[200][12]/P0001 ,
		_w12988_,
		_w23037_
	);
	LUT2 #(
		.INIT('h8)
	) name12526 (
		\wishbone_bd_ram_mem1_reg[242][12]/P0001 ,
		_w12932_,
		_w23038_
	);
	LUT2 #(
		.INIT('h8)
	) name12527 (
		\wishbone_bd_ram_mem1_reg[247][12]/P0001 ,
		_w12818_,
		_w23039_
	);
	LUT2 #(
		.INIT('h8)
	) name12528 (
		\wishbone_bd_ram_mem1_reg[240][12]/P0001 ,
		_w12864_,
		_w23040_
	);
	LUT2 #(
		.INIT('h8)
	) name12529 (
		\wishbone_bd_ram_mem1_reg[6][12]/P0001 ,
		_w12968_,
		_w23041_
	);
	LUT2 #(
		.INIT('h8)
	) name12530 (
		\wishbone_bd_ram_mem1_reg[81][12]/P0001 ,
		_w12950_,
		_w23042_
	);
	LUT2 #(
		.INIT('h8)
	) name12531 (
		\wishbone_bd_ram_mem1_reg[218][12]/P0001 ,
		_w13206_,
		_w23043_
	);
	LUT2 #(
		.INIT('h8)
	) name12532 (
		\wishbone_bd_ram_mem1_reg[57][12]/P0001 ,
		_w13116_,
		_w23044_
	);
	LUT2 #(
		.INIT('h8)
	) name12533 (
		\wishbone_bd_ram_mem1_reg[134][12]/P0001 ,
		_w12763_,
		_w23045_
	);
	LUT2 #(
		.INIT('h8)
	) name12534 (
		\wishbone_bd_ram_mem1_reg[183][12]/P0001 ,
		_w12787_,
		_w23046_
	);
	LUT2 #(
		.INIT('h8)
	) name12535 (
		\wishbone_bd_ram_mem1_reg[193][12]/P0001 ,
		_w13056_,
		_w23047_
	);
	LUT2 #(
		.INIT('h8)
	) name12536 (
		\wishbone_bd_ram_mem1_reg[126][12]/P0001 ,
		_w13218_,
		_w23048_
	);
	LUT2 #(
		.INIT('h8)
	) name12537 (
		\wishbone_bd_ram_mem1_reg[35][12]/P0001 ,
		_w12703_,
		_w23049_
	);
	LUT2 #(
		.INIT('h8)
	) name12538 (
		\wishbone_bd_ram_mem1_reg[191][12]/P0001 ,
		_w13034_,
		_w23050_
	);
	LUT2 #(
		.INIT('h8)
	) name12539 (
		\wishbone_bd_ram_mem1_reg[118][12]/P0001 ,
		_w12830_,
		_w23051_
	);
	LUT2 #(
		.INIT('h8)
	) name12540 (
		\wishbone_bd_ram_mem1_reg[231][12]/P0001 ,
		_w12856_,
		_w23052_
	);
	LUT2 #(
		.INIT('h8)
	) name12541 (
		\wishbone_bd_ram_mem1_reg[121][12]/P0001 ,
		_w13078_,
		_w23053_
	);
	LUT2 #(
		.INIT('h8)
	) name12542 (
		\wishbone_bd_ram_mem1_reg[229][12]/P0001 ,
		_w12711_,
		_w23054_
	);
	LUT2 #(
		.INIT('h8)
	) name12543 (
		\wishbone_bd_ram_mem1_reg[144][12]/P0001 ,
		_w12756_,
		_w23055_
	);
	LUT2 #(
		.INIT('h8)
	) name12544 (
		\wishbone_bd_ram_mem1_reg[49][12]/P0001 ,
		_w12994_,
		_w23056_
	);
	LUT2 #(
		.INIT('h8)
	) name12545 (
		\wishbone_bd_ram_mem1_reg[220][12]/P0001 ,
		_w13066_,
		_w23057_
	);
	LUT2 #(
		.INIT('h8)
	) name12546 (
		\wishbone_bd_ram_mem1_reg[210][12]/P0001 ,
		_w12924_,
		_w23058_
	);
	LUT2 #(
		.INIT('h8)
	) name12547 (
		\wishbone_bd_ram_mem1_reg[104][12]/P0001 ,
		_w13148_,
		_w23059_
	);
	LUT2 #(
		.INIT('h8)
	) name12548 (
		\wishbone_bd_ram_mem1_reg[248][12]/P0001 ,
		_w12789_,
		_w23060_
	);
	LUT2 #(
		.INIT('h8)
	) name12549 (
		\wishbone_bd_ram_mem1_reg[241][12]/P0001 ,
		_w13006_,
		_w23061_
	);
	LUT2 #(
		.INIT('h8)
	) name12550 (
		\wishbone_bd_ram_mem1_reg[127][12]/P0001 ,
		_w13164_,
		_w23062_
	);
	LUT2 #(
		.INIT('h8)
	) name12551 (
		\wishbone_bd_ram_mem1_reg[82][12]/P0001 ,
		_w12942_,
		_w23063_
	);
	LUT2 #(
		.INIT('h8)
	) name12552 (
		\wishbone_bd_ram_mem1_reg[55][12]/P0001 ,
		_w12785_,
		_w23064_
	);
	LUT2 #(
		.INIT('h8)
	) name12553 (
		\wishbone_bd_ram_mem1_reg[205][12]/P0001 ,
		_w13068_,
		_w23065_
	);
	LUT2 #(
		.INIT('h8)
	) name12554 (
		\wishbone_bd_ram_mem1_reg[175][12]/P0001 ,
		_w13126_,
		_w23066_
	);
	LUT2 #(
		.INIT('h8)
	) name12555 (
		\wishbone_bd_ram_mem1_reg[43][12]/P0001 ,
		_w13200_,
		_w23067_
	);
	LUT2 #(
		.INIT('h8)
	) name12556 (
		\wishbone_bd_ram_mem1_reg[135][12]/P0001 ,
		_w13124_,
		_w23068_
	);
	LUT2 #(
		.INIT('h8)
	) name12557 (
		\wishbone_bd_ram_mem1_reg[103][12]/P0001 ,
		_w12846_,
		_w23069_
	);
	LUT2 #(
		.INIT('h8)
	) name12558 (
		\wishbone_bd_ram_mem1_reg[219][12]/P0001 ,
		_w12806_,
		_w23070_
	);
	LUT2 #(
		.INIT('h8)
	) name12559 (
		\wishbone_bd_ram_mem1_reg[112][12]/P0001 ,
		_w12733_,
		_w23071_
	);
	LUT2 #(
		.INIT('h8)
	) name12560 (
		\wishbone_bd_ram_mem1_reg[249][12]/P0001 ,
		_w12900_,
		_w23072_
	);
	LUT2 #(
		.INIT('h8)
	) name12561 (
		\wishbone_bd_ram_mem1_reg[201][12]/P0001 ,
		_w12822_,
		_w23073_
	);
	LUT2 #(
		.INIT('h8)
	) name12562 (
		\wishbone_bd_ram_mem1_reg[47][12]/P0001 ,
		_w12904_,
		_w23074_
	);
	LUT2 #(
		.INIT('h8)
	) name12563 (
		\wishbone_bd_ram_mem1_reg[252][12]/P0001 ,
		_w13080_,
		_w23075_
	);
	LUT2 #(
		.INIT('h8)
	) name12564 (
		\wishbone_bd_ram_mem1_reg[180][12]/P0001 ,
		_w12791_,
		_w23076_
	);
	LUT2 #(
		.INIT('h8)
	) name12565 (
		\wishbone_bd_ram_mem1_reg[1][12]/P0001 ,
		_w13014_,
		_w23077_
	);
	LUT2 #(
		.INIT('h8)
	) name12566 (
		\wishbone_bd_ram_mem1_reg[31][12]/P0001 ,
		_w13198_,
		_w23078_
	);
	LUT2 #(
		.INIT('h8)
	) name12567 (
		\wishbone_bd_ram_mem1_reg[227][12]/P0001 ,
		_w12936_,
		_w23079_
	);
	LUT2 #(
		.INIT('h8)
	) name12568 (
		\wishbone_bd_ram_mem1_reg[199][12]/P0001 ,
		_w12768_,
		_w23080_
	);
	LUT2 #(
		.INIT('h8)
	) name12569 (
		\wishbone_bd_ram_mem1_reg[244][12]/P0001 ,
		_w12747_,
		_w23081_
	);
	LUT2 #(
		.INIT('h8)
	) name12570 (
		\wishbone_bd_ram_mem1_reg[26][12]/P0001 ,
		_w12699_,
		_w23082_
	);
	LUT2 #(
		.INIT('h8)
	) name12571 (
		\wishbone_bd_ram_mem1_reg[216][12]/P0001 ,
		_w13028_,
		_w23083_
	);
	LUT2 #(
		.INIT('h8)
	) name12572 (
		\wishbone_bd_ram_mem1_reg[174][12]/P0001 ,
		_w12972_,
		_w23084_
	);
	LUT2 #(
		.INIT('h8)
	) name12573 (
		\wishbone_bd_ram_mem1_reg[77][12]/P0001 ,
		_w12982_,
		_w23085_
	);
	LUT2 #(
		.INIT('h8)
	) name12574 (
		\wishbone_bd_ram_mem1_reg[120][12]/P0001 ,
		_w12707_,
		_w23086_
	);
	LUT2 #(
		.INIT('h8)
	) name12575 (
		\wishbone_bd_ram_mem1_reg[217][12]/P0001 ,
		_w13188_,
		_w23087_
	);
	LUT2 #(
		.INIT('h8)
	) name12576 (
		\wishbone_bd_ram_mem1_reg[234][12]/P0001 ,
		_w13214_,
		_w23088_
	);
	LUT2 #(
		.INIT('h8)
	) name12577 (
		\wishbone_bd_ram_mem1_reg[5][12]/P0001 ,
		_w12878_,
		_w23089_
	);
	LUT2 #(
		.INIT('h8)
	) name12578 (
		\wishbone_bd_ram_mem1_reg[62][12]/P0001 ,
		_w12673_,
		_w23090_
	);
	LUT2 #(
		.INIT('h8)
	) name12579 (
		\wishbone_bd_ram_mem1_reg[155][12]/P0001 ,
		_w13122_,
		_w23091_
	);
	LUT2 #(
		.INIT('h8)
	) name12580 (
		\wishbone_bd_ram_mem1_reg[27][12]/P0001 ,
		_w12880_,
		_w23092_
	);
	LUT2 #(
		.INIT('h8)
	) name12581 (
		\wishbone_bd_ram_mem1_reg[111][12]/P0001 ,
		_w12744_,
		_w23093_
	);
	LUT2 #(
		.INIT('h8)
	) name12582 (
		\wishbone_bd_ram_mem1_reg[225][12]/P0001 ,
		_w13092_,
		_w23094_
	);
	LUT2 #(
		.INIT('h8)
	) name12583 (
		\wishbone_bd_ram_mem1_reg[243][12]/P0001 ,
		_w12804_,
		_w23095_
	);
	LUT2 #(
		.INIT('h8)
	) name12584 (
		\wishbone_bd_ram_mem1_reg[96][12]/P0001 ,
		_w12912_,
		_w23096_
	);
	LUT2 #(
		.INIT('h8)
	) name12585 (
		\wishbone_bd_ram_mem1_reg[239][12]/P0001 ,
		_w12862_,
		_w23097_
	);
	LUT2 #(
		.INIT('h8)
	) name12586 (
		\wishbone_bd_ram_mem1_reg[7][12]/P0001 ,
		_w12728_,
		_w23098_
	);
	LUT2 #(
		.INIT('h8)
	) name12587 (
		\wishbone_bd_ram_mem1_reg[8][12]/P0001 ,
		_w12920_,
		_w23099_
	);
	LUT2 #(
		.INIT('h8)
	) name12588 (
		\wishbone_bd_ram_mem1_reg[245][12]/P0001 ,
		_w13022_,
		_w23100_
	);
	LUT2 #(
		.INIT('h8)
	) name12589 (
		\wishbone_bd_ram_mem1_reg[105][12]/P0001 ,
		_w12751_,
		_w23101_
	);
	LUT2 #(
		.INIT('h8)
	) name12590 (
		\wishbone_bd_ram_mem1_reg[106][12]/P0001 ,
		_w12713_,
		_w23102_
	);
	LUT2 #(
		.INIT('h8)
	) name12591 (
		\wishbone_bd_ram_mem1_reg[129][12]/P0001 ,
		_w12776_,
		_w23103_
	);
	LUT2 #(
		.INIT('h8)
	) name12592 (
		\wishbone_bd_ram_mem1_reg[215][12]/P0001 ,
		_w12974_,
		_w23104_
	);
	LUT2 #(
		.INIT('h8)
	) name12593 (
		\wishbone_bd_ram_mem1_reg[52][12]/P0001 ,
		_w13082_,
		_w23105_
	);
	LUT2 #(
		.INIT('h8)
	) name12594 (
		\wishbone_bd_ram_mem1_reg[147][12]/P0001 ,
		_w13146_,
		_w23106_
	);
	LUT2 #(
		.INIT('h8)
	) name12595 (
		\wishbone_bd_ram_mem1_reg[230][12]/P0001 ,
		_w13036_,
		_w23107_
	);
	LUT2 #(
		.INIT('h8)
	) name12596 (
		\wishbone_bd_ram_mem1_reg[158][12]/P0001 ,
		_w12898_,
		_w23108_
	);
	LUT2 #(
		.INIT('h8)
	) name12597 (
		\wishbone_bd_ram_mem1_reg[187][12]/P0001 ,
		_w13196_,
		_w23109_
	);
	LUT2 #(
		.INIT('h8)
	) name12598 (
		\wishbone_bd_ram_mem1_reg[54][12]/P0001 ,
		_w12770_,
		_w23110_
	);
	LUT2 #(
		.INIT('h8)
	) name12599 (
		\wishbone_bd_ram_mem1_reg[72][12]/P0001 ,
		_w12810_,
		_w23111_
	);
	LUT2 #(
		.INIT('h8)
	) name12600 (
		\wishbone_bd_ram_mem1_reg[184][12]/P0001 ,
		_w13062_,
		_w23112_
	);
	LUT2 #(
		.INIT('h8)
	) name12601 (
		\wishbone_bd_ram_mem1_reg[11][12]/P0001 ,
		_w13194_,
		_w23113_
	);
	LUT2 #(
		.INIT('h8)
	) name12602 (
		\wishbone_bd_ram_mem1_reg[214][12]/P0001 ,
		_w12984_,
		_w23114_
	);
	LUT2 #(
		.INIT('h8)
	) name12603 (
		\wishbone_bd_ram_mem1_reg[80][12]/P0001 ,
		_w12689_,
		_w23115_
	);
	LUT2 #(
		.INIT('h8)
	) name12604 (
		\wishbone_bd_ram_mem1_reg[91][12]/P0001 ,
		_w13074_,
		_w23116_
	);
	LUT2 #(
		.INIT('h8)
	) name12605 (
		\wishbone_bd_ram_mem1_reg[102][12]/P0001 ,
		_w12685_,
		_w23117_
	);
	LUT2 #(
		.INIT('h8)
	) name12606 (
		\wishbone_bd_ram_mem1_reg[67][12]/P0001 ,
		_w13134_,
		_w23118_
	);
	LUT2 #(
		.INIT('h8)
	) name12607 (
		\wishbone_bd_ram_mem1_reg[50][12]/P0001 ,
		_w13150_,
		_w23119_
	);
	LUT2 #(
		.INIT('h8)
	) name12608 (
		\wishbone_bd_ram_mem1_reg[61][12]/P0001 ,
		_w12725_,
		_w23120_
	);
	LUT2 #(
		.INIT('h8)
	) name12609 (
		\wishbone_bd_ram_mem1_reg[53][12]/P0001 ,
		_w13020_,
		_w23121_
	);
	LUT2 #(
		.INIT('h8)
	) name12610 (
		\wishbone_bd_ram_mem1_reg[246][12]/P0001 ,
		_w13076_,
		_w23122_
	);
	LUT2 #(
		.INIT('h8)
	) name12611 (
		\wishbone_bd_ram_mem1_reg[133][12]/P0001 ,
		_w12761_,
		_w23123_
	);
	LUT2 #(
		.INIT('h8)
	) name12612 (
		\wishbone_bd_ram_mem1_reg[221][12]/P0001 ,
		_w12802_,
		_w23124_
	);
	LUT2 #(
		.INIT('h8)
	) name12613 (
		\wishbone_bd_ram_mem1_reg[226][12]/P0001 ,
		_w13138_,
		_w23125_
	);
	LUT2 #(
		.INIT('h8)
	) name12614 (
		\wishbone_bd_ram_mem1_reg[88][12]/P0001 ,
		_w12860_,
		_w23126_
	);
	LUT2 #(
		.INIT('h8)
	) name12615 (
		\wishbone_bd_ram_mem1_reg[3][12]/P0001 ,
		_w12866_,
		_w23127_
	);
	LUT2 #(
		.INIT('h8)
	) name12616 (
		\wishbone_bd_ram_mem1_reg[159][12]/P0001 ,
		_w12774_,
		_w23128_
	);
	LUT2 #(
		.INIT('h8)
	) name12617 (
		\wishbone_bd_ram_mem1_reg[156][12]/P0001 ,
		_w13190_,
		_w23129_
	);
	LUT2 #(
		.INIT('h8)
	) name12618 (
		\wishbone_bd_ram_mem1_reg[251][12]/P0001 ,
		_w13054_,
		_w23130_
	);
	LUT2 #(
		.INIT('h8)
	) name12619 (
		\wishbone_bd_ram_mem1_reg[98][12]/P0001 ,
		_w12816_,
		_w23131_
	);
	LUT2 #(
		.INIT('h8)
	) name12620 (
		\wishbone_bd_ram_mem1_reg[130][12]/P0001 ,
		_w12914_,
		_w23132_
	);
	LUT2 #(
		.INIT('h8)
	) name12621 (
		\wishbone_bd_ram_mem1_reg[100][12]/P0001 ,
		_w12960_,
		_w23133_
	);
	LUT2 #(
		.INIT('h8)
	) name12622 (
		\wishbone_bd_ram_mem1_reg[99][12]/P0001 ,
		_w13038_,
		_w23134_
	);
	LUT2 #(
		.INIT('h8)
	) name12623 (
		\wishbone_bd_ram_mem1_reg[71][12]/P0001 ,
		_w12798_,
		_w23135_
	);
	LUT2 #(
		.INIT('h8)
	) name12624 (
		\wishbone_bd_ram_mem1_reg[2][12]/P0001 ,
		_w13088_,
		_w23136_
	);
	LUT2 #(
		.INIT('h8)
	) name12625 (
		\wishbone_bd_ram_mem1_reg[168][12]/P0001 ,
		_w13208_,
		_w23137_
	);
	LUT2 #(
		.INIT('h8)
	) name12626 (
		\wishbone_bd_ram_mem1_reg[203][12]/P0001 ,
		_w13158_,
		_w23138_
	);
	LUT2 #(
		.INIT('h8)
	) name12627 (
		\wishbone_bd_ram_mem1_reg[172][12]/P0001 ,
		_w12944_,
		_w23139_
	);
	LUT2 #(
		.INIT('h8)
	) name12628 (
		\wishbone_bd_ram_mem1_reg[213][12]/P0001 ,
		_w13002_,
		_w23140_
	);
	LUT2 #(
		.INIT('h8)
	) name12629 (
		\wishbone_bd_ram_mem1_reg[150][12]/P0001 ,
		_w13136_,
		_w23141_
	);
	LUT2 #(
		.INIT('h8)
	) name12630 (
		\wishbone_bd_ram_mem1_reg[157][12]/P0001 ,
		_w12926_,
		_w23142_
	);
	LUT2 #(
		.INIT('h8)
	) name12631 (
		\wishbone_bd_ram_mem1_reg[87][12]/P0001 ,
		_w13154_,
		_w23143_
	);
	LUT2 #(
		.INIT('h8)
	) name12632 (
		\wishbone_bd_ram_mem1_reg[84][12]/P0001 ,
		_w12934_,
		_w23144_
	);
	LUT2 #(
		.INIT('h8)
	) name12633 (
		\wishbone_bd_ram_mem1_reg[186][12]/P0001 ,
		_w12783_,
		_w23145_
	);
	LUT2 #(
		.INIT('h8)
	) name12634 (
		\wishbone_bd_ram_mem1_reg[114][12]/P0001 ,
		_w13202_,
		_w23146_
	);
	LUT2 #(
		.INIT('h8)
	) name12635 (
		\wishbone_bd_ram_mem1_reg[9][12]/P0001 ,
		_w12808_,
		_w23147_
	);
	LUT2 #(
		.INIT('h8)
	) name12636 (
		\wishbone_bd_ram_mem1_reg[228][12]/P0001 ,
		_w12765_,
		_w23148_
	);
	LUT2 #(
		.INIT('h8)
	) name12637 (
		\wishbone_bd_ram_mem1_reg[79][12]/P0001 ,
		_w13212_,
		_w23149_
	);
	LUT2 #(
		.INIT('h8)
	) name12638 (
		\wishbone_bd_ram_mem1_reg[40][12]/P0001 ,
		_w13132_,
		_w23150_
	);
	LUT2 #(
		.INIT('h8)
	) name12639 (
		\wishbone_bd_ram_mem1_reg[48][12]/P0001 ,
		_w12970_,
		_w23151_
	);
	LUT2 #(
		.INIT('h8)
	) name12640 (
		\wishbone_bd_ram_mem1_reg[237][12]/P0001 ,
		_w12990_,
		_w23152_
	);
	LUT2 #(
		.INIT('h8)
	) name12641 (
		\wishbone_bd_ram_mem1_reg[107][12]/P0001 ,
		_w12749_,
		_w23153_
	);
	LUT2 #(
		.INIT('h8)
	) name12642 (
		\wishbone_bd_ram_mem1_reg[16][12]/P0001 ,
		_w13140_,
		_w23154_
	);
	LUT2 #(
		.INIT('h8)
	) name12643 (
		\wishbone_bd_ram_mem1_reg[51][12]/P0001 ,
		_w13024_,
		_w23155_
	);
	LUT2 #(
		.INIT('h8)
	) name12644 (
		\wishbone_bd_ram_mem1_reg[93][12]/P0001 ,
		_w13016_,
		_w23156_
	);
	LUT2 #(
		.INIT('h8)
	) name12645 (
		\wishbone_bd_ram_mem1_reg[254][12]/P0001 ,
		_w12892_,
		_w23157_
	);
	LUT2 #(
		.INIT('h8)
	) name12646 (
		\wishbone_bd_ram_mem1_reg[222][12]/P0001 ,
		_w13094_,
		_w23158_
	);
	LUT2 #(
		.INIT('h8)
	) name12647 (
		\wishbone_bd_ram_mem1_reg[39][12]/P0001 ,
		_w13018_,
		_w23159_
	);
	LUT2 #(
		.INIT('h8)
	) name12648 (
		\wishbone_bd_ram_mem1_reg[152][12]/P0001 ,
		_w12966_,
		_w23160_
	);
	LUT2 #(
		.INIT('h8)
	) name12649 (
		\wishbone_bd_ram_mem1_reg[195][12]/P0001 ,
		_w13144_,
		_w23161_
	);
	LUT2 #(
		.INIT('h8)
	) name12650 (
		\wishbone_bd_ram_mem1_reg[113][12]/P0001 ,
		_w13026_,
		_w23162_
	);
	LUT2 #(
		.INIT('h8)
	) name12651 (
		\wishbone_bd_ram_mem1_reg[34][12]/P0001 ,
		_w12930_,
		_w23163_
	);
	LUT2 #(
		.INIT('h8)
	) name12652 (
		\wishbone_bd_ram_mem1_reg[21][12]/P0001 ,
		_w12906_,
		_w23164_
	);
	LUT2 #(
		.INIT('h8)
	) name12653 (
		\wishbone_bd_ram_mem1_reg[140][12]/P0001 ,
		_w12894_,
		_w23165_
	);
	LUT2 #(
		.INIT('h8)
	) name12654 (
		\wishbone_bd_ram_mem1_reg[75][12]/P0001 ,
		_w12826_,
		_w23166_
	);
	LUT2 #(
		.INIT('h8)
	) name12655 (
		\wishbone_bd_ram_mem1_reg[137][12]/P0001 ,
		_w13168_,
		_w23167_
	);
	LUT2 #(
		.INIT('h8)
	) name12656 (
		\wishbone_bd_ram_mem1_reg[197][12]/P0001 ,
		_w12834_,
		_w23168_
	);
	LUT2 #(
		.INIT('h8)
	) name12657 (
		\wishbone_bd_ram_mem1_reg[253][12]/P0001 ,
		_w13100_,
		_w23169_
	);
	LUT2 #(
		.INIT('h8)
	) name12658 (
		\wishbone_bd_ram_mem1_reg[44][12]/P0001 ,
		_w12896_,
		_w23170_
	);
	LUT2 #(
		.INIT('h8)
	) name12659 (
		\wishbone_bd_ram_mem1_reg[68][12]/P0001 ,
		_w12946_,
		_w23171_
	);
	LUT2 #(
		.INIT('h8)
	) name12660 (
		\wishbone_bd_ram_mem1_reg[15][12]/P0001 ,
		_w13210_,
		_w23172_
	);
	LUT2 #(
		.INIT('h8)
	) name12661 (
		\wishbone_bd_ram_mem1_reg[42][12]/P0001 ,
		_w12842_,
		_w23173_
	);
	LUT2 #(
		.INIT('h8)
	) name12662 (
		\wishbone_bd_ram_mem1_reg[46][12]/P0001 ,
		_w12884_,
		_w23174_
	);
	LUT2 #(
		.INIT('h8)
	) name12663 (
		\wishbone_bd_ram_mem1_reg[190][12]/P0001 ,
		_w12858_,
		_w23175_
	);
	LUT2 #(
		.INIT('h8)
	) name12664 (
		\wishbone_bd_ram_mem1_reg[198][12]/P0001 ,
		_w12832_,
		_w23176_
	);
	LUT2 #(
		.INIT('h8)
	) name12665 (
		\wishbone_bd_ram_mem1_reg[122][12]/P0001 ,
		_w13130_,
		_w23177_
	);
	LUT2 #(
		.INIT('h8)
	) name12666 (
		\wishbone_bd_ram_mem1_reg[92][12]/P0001 ,
		_w13010_,
		_w23178_
	);
	LUT2 #(
		.INIT('h8)
	) name12667 (
		\wishbone_bd_ram_mem1_reg[142][12]/P0001 ,
		_w12928_,
		_w23179_
	);
	LUT2 #(
		.INIT('h8)
	) name12668 (
		\wishbone_bd_ram_mem1_reg[204][12]/P0001 ,
		_w13162_,
		_w23180_
	);
	LUT2 #(
		.INIT('h8)
	) name12669 (
		\wishbone_bd_ram_mem1_reg[12][12]/P0001 ,
		_w13118_,
		_w23181_
	);
	LUT2 #(
		.INIT('h8)
	) name12670 (
		\wishbone_bd_ram_mem1_reg[143][12]/P0001 ,
		_w12922_,
		_w23182_
	);
	LUT2 #(
		.INIT('h8)
	) name12671 (
		\wishbone_bd_ram_mem1_reg[132][12]/P0001 ,
		_w12992_,
		_w23183_
	);
	LUT2 #(
		.INIT('h8)
	) name12672 (
		\wishbone_bd_ram_mem1_reg[167][12]/P0001 ,
		_w12986_,
		_w23184_
	);
	LUT2 #(
		.INIT('h8)
	) name12673 (
		\wishbone_bd_ram_mem1_reg[19][12]/P0001 ,
		_w13012_,
		_w23185_
	);
	LUT2 #(
		.INIT('h8)
	) name12674 (
		\wishbone_bd_ram_mem1_reg[115][12]/P0001 ,
		_w13112_,
		_w23186_
	);
	LUT2 #(
		.INIT('h8)
	) name12675 (
		\wishbone_bd_ram_mem1_reg[119][12]/P0001 ,
		_w13048_,
		_w23187_
	);
	LUT2 #(
		.INIT('h8)
	) name12676 (
		\wishbone_bd_ram_mem1_reg[64][12]/P0001 ,
		_w12976_,
		_w23188_
	);
	LUT2 #(
		.INIT('h8)
	) name12677 (
		\wishbone_bd_ram_mem1_reg[25][12]/P0001 ,
		_w13108_,
		_w23189_
	);
	LUT2 #(
		.INIT('h8)
	) name12678 (
		\wishbone_bd_ram_mem1_reg[188][12]/P0001 ,
		_w12948_,
		_w23190_
	);
	LUT2 #(
		.INIT('h8)
	) name12679 (
		\wishbone_bd_ram_mem1_reg[177][12]/P0001 ,
		_w12996_,
		_w23191_
	);
	LUT2 #(
		.INIT('h8)
	) name12680 (
		\wishbone_bd_ram_mem1_reg[89][12]/P0001 ,
		_w12964_,
		_w23192_
	);
	LUT2 #(
		.INIT('h8)
	) name12681 (
		\wishbone_bd_ram_mem1_reg[154][12]/P0001 ,
		_w12962_,
		_w23193_
	);
	LUT2 #(
		.INIT('h8)
	) name12682 (
		\wishbone_bd_ram_mem1_reg[101][12]/P0001 ,
		_w13192_,
		_w23194_
	);
	LUT2 #(
		.INIT('h8)
	) name12683 (
		\wishbone_bd_ram_mem1_reg[108][12]/P0001 ,
		_w13156_,
		_w23195_
	);
	LUT2 #(
		.INIT('h8)
	) name12684 (
		\wishbone_bd_ram_mem1_reg[69][12]/P0001 ,
		_w12738_,
		_w23196_
	);
	LUT2 #(
		.INIT('h8)
	) name12685 (
		\wishbone_bd_ram_mem1_reg[41][12]/P0001 ,
		_w13052_,
		_w23197_
	);
	LUT2 #(
		.INIT('h8)
	) name12686 (
		\wishbone_bd_ram_mem1_reg[207][12]/P0001 ,
		_w13180_,
		_w23198_
	);
	LUT2 #(
		.INIT('h8)
	) name12687 (
		\wishbone_bd_ram_mem1_reg[60][12]/P0001 ,
		_w13204_,
		_w23199_
	);
	LUT2 #(
		.INIT('h8)
	) name12688 (
		\wishbone_bd_ram_mem1_reg[18][12]/P0001 ,
		_w12679_,
		_w23200_
	);
	LUT2 #(
		.INIT('h8)
	) name12689 (
		\wishbone_bd_ram_mem1_reg[10][12]/P0001 ,
		_w13172_,
		_w23201_
	);
	LUT2 #(
		.INIT('h8)
	) name12690 (
		\wishbone_bd_ram_mem1_reg[206][12]/P0001 ,
		_w12954_,
		_w23202_
	);
	LUT2 #(
		.INIT('h8)
	) name12691 (
		\wishbone_bd_ram_mem1_reg[164][12]/P0001 ,
		_w12876_,
		_w23203_
	);
	LUT2 #(
		.INIT('h8)
	) name12692 (
		\wishbone_bd_ram_mem1_reg[149][12]/P0001 ,
		_w12741_,
		_w23204_
	);
	LUT2 #(
		.INIT('h8)
	) name12693 (
		\wishbone_bd_ram_mem1_reg[58][12]/P0001 ,
		_w13070_,
		_w23205_
	);
	LUT2 #(
		.INIT('h8)
	) name12694 (
		\wishbone_bd_ram_mem1_reg[162][12]/P0001 ,
		_w13098_,
		_w23206_
	);
	LUT2 #(
		.INIT('h8)
	) name12695 (
		\wishbone_bd_ram_mem1_reg[56][12]/P0001 ,
		_w12778_,
		_w23207_
	);
	LUT2 #(
		.INIT('h8)
	) name12696 (
		\wishbone_bd_ram_mem1_reg[179][12]/P0001 ,
		_w13050_,
		_w23208_
	);
	LUT2 #(
		.INIT('h8)
	) name12697 (
		\wishbone_bd_ram_mem1_reg[255][12]/P0001 ,
		_w13072_,
		_w23209_
	);
	LUT2 #(
		.INIT('h8)
	) name12698 (
		\wishbone_bd_ram_mem1_reg[37][12]/P0001 ,
		_w13102_,
		_w23210_
	);
	LUT2 #(
		.INIT('h8)
	) name12699 (
		\wishbone_bd_ram_mem1_reg[224][12]/P0001 ,
		_w12902_,
		_w23211_
	);
	LUT2 #(
		.INIT('h8)
	) name12700 (
		\wishbone_bd_ram_mem1_reg[182][12]/P0001 ,
		_w12820_,
		_w23212_
	);
	LUT2 #(
		.INIT('h8)
	) name12701 (
		\wishbone_bd_ram_mem1_reg[0][12]/P0001 ,
		_w12717_,
		_w23213_
	);
	LUT2 #(
		.INIT('h8)
	) name12702 (
		\wishbone_bd_ram_mem1_reg[32][12]/P0001 ,
		_w13120_,
		_w23214_
	);
	LUT2 #(
		.INIT('h8)
	) name12703 (
		\wishbone_bd_ram_mem1_reg[178][12]/P0001 ,
		_w12886_,
		_w23215_
	);
	LUT2 #(
		.INIT('h8)
	) name12704 (
		\wishbone_bd_ram_mem1_reg[30][12]/P0001 ,
		_w13104_,
		_w23216_
	);
	LUT2 #(
		.INIT('h8)
	) name12705 (
		\wishbone_bd_ram_mem1_reg[171][12]/P0001 ,
		_w12910_,
		_w23217_
	);
	LUT2 #(
		.INIT('h8)
	) name12706 (
		\wishbone_bd_ram_mem1_reg[160][12]/P0001 ,
		_w12872_,
		_w23218_
	);
	LUT2 #(
		.INIT('h8)
	) name12707 (
		\wishbone_bd_ram_mem1_reg[45][12]/P0001 ,
		_w12908_,
		_w23219_
	);
	LUT2 #(
		.INIT('h8)
	) name12708 (
		\wishbone_bd_ram_mem1_reg[170][12]/P0001 ,
		_w13030_,
		_w23220_
	);
	LUT2 #(
		.INIT('h8)
	) name12709 (
		\wishbone_bd_ram_mem1_reg[94][12]/P0001 ,
		_w13186_,
		_w23221_
	);
	LUT2 #(
		.INIT('h8)
	) name12710 (
		\wishbone_bd_ram_mem1_reg[74][12]/P0001 ,
		_w12812_,
		_w23222_
	);
	LUT2 #(
		.INIT('h8)
	) name12711 (
		\wishbone_bd_ram_mem1_reg[70][12]/P0001 ,
		_w12840_,
		_w23223_
	);
	LUT2 #(
		.INIT('h8)
	) name12712 (
		\wishbone_bd_ram_mem1_reg[148][12]/P0001 ,
		_w13000_,
		_w23224_
	);
	LUT2 #(
		.INIT('h8)
	) name12713 (
		\wishbone_bd_ram_mem1_reg[138][12]/P0001 ,
		_w12958_,
		_w23225_
	);
	LUT2 #(
		.INIT('h8)
	) name12714 (
		\wishbone_bd_ram_mem1_reg[109][12]/P0001 ,
		_w12888_,
		_w23226_
	);
	LUT2 #(
		.INIT('h8)
	) name12715 (
		\wishbone_bd_ram_mem1_reg[14][12]/P0001 ,
		_w13086_,
		_w23227_
	);
	LUT2 #(
		.INIT('h8)
	) name12716 (
		\wishbone_bd_ram_mem1_reg[163][12]/P0001 ,
		_w12882_,
		_w23228_
	);
	LUT2 #(
		.INIT('h8)
	) name12717 (
		\wishbone_bd_ram_mem1_reg[173][12]/P0001 ,
		_w12854_,
		_w23229_
	);
	LUT2 #(
		.INIT('h8)
	) name12718 (
		\wishbone_bd_ram_mem1_reg[192][12]/P0001 ,
		_w12938_,
		_w23230_
	);
	LUT2 #(
		.INIT('h8)
	) name12719 (
		\wishbone_bd_ram_mem1_reg[185][12]/P0001 ,
		_w12940_,
		_w23231_
	);
	LUT2 #(
		.INIT('h8)
	) name12720 (
		\wishbone_bd_ram_mem1_reg[36][12]/P0001 ,
		_w12800_,
		_w23232_
	);
	LUT2 #(
		.INIT('h8)
	) name12721 (
		\wishbone_bd_ram_mem1_reg[73][12]/P0001 ,
		_w12918_,
		_w23233_
	);
	LUT2 #(
		.INIT('h8)
	) name12722 (
		\wishbone_bd_ram_mem1_reg[136][12]/P0001 ,
		_w13064_,
		_w23234_
	);
	LUT2 #(
		.INIT('h8)
	) name12723 (
		\wishbone_bd_ram_mem1_reg[209][12]/P0001 ,
		_w13152_,
		_w23235_
	);
	LUT2 #(
		.INIT('h8)
	) name12724 (
		\wishbone_bd_ram_mem1_reg[176][12]/P0001 ,
		_w12868_,
		_w23236_
	);
	LUT2 #(
		.INIT('h8)
	) name12725 (
		\wishbone_bd_ram_mem1_reg[65][12]/P0001 ,
		_w13176_,
		_w23237_
	);
	LUT2 #(
		.INIT('h8)
	) name12726 (
		\wishbone_bd_ram_mem1_reg[151][12]/P0001 ,
		_w13142_,
		_w23238_
	);
	LUT2 #(
		.INIT('h1)
	) name12727 (
		_w22983_,
		_w22984_,
		_w23239_
	);
	LUT2 #(
		.INIT('h1)
	) name12728 (
		_w22985_,
		_w22986_,
		_w23240_
	);
	LUT2 #(
		.INIT('h1)
	) name12729 (
		_w22987_,
		_w22988_,
		_w23241_
	);
	LUT2 #(
		.INIT('h1)
	) name12730 (
		_w22989_,
		_w22990_,
		_w23242_
	);
	LUT2 #(
		.INIT('h1)
	) name12731 (
		_w22991_,
		_w22992_,
		_w23243_
	);
	LUT2 #(
		.INIT('h1)
	) name12732 (
		_w22993_,
		_w22994_,
		_w23244_
	);
	LUT2 #(
		.INIT('h1)
	) name12733 (
		_w22995_,
		_w22996_,
		_w23245_
	);
	LUT2 #(
		.INIT('h1)
	) name12734 (
		_w22997_,
		_w22998_,
		_w23246_
	);
	LUT2 #(
		.INIT('h1)
	) name12735 (
		_w22999_,
		_w23000_,
		_w23247_
	);
	LUT2 #(
		.INIT('h1)
	) name12736 (
		_w23001_,
		_w23002_,
		_w23248_
	);
	LUT2 #(
		.INIT('h1)
	) name12737 (
		_w23003_,
		_w23004_,
		_w23249_
	);
	LUT2 #(
		.INIT('h1)
	) name12738 (
		_w23005_,
		_w23006_,
		_w23250_
	);
	LUT2 #(
		.INIT('h1)
	) name12739 (
		_w23007_,
		_w23008_,
		_w23251_
	);
	LUT2 #(
		.INIT('h1)
	) name12740 (
		_w23009_,
		_w23010_,
		_w23252_
	);
	LUT2 #(
		.INIT('h1)
	) name12741 (
		_w23011_,
		_w23012_,
		_w23253_
	);
	LUT2 #(
		.INIT('h1)
	) name12742 (
		_w23013_,
		_w23014_,
		_w23254_
	);
	LUT2 #(
		.INIT('h1)
	) name12743 (
		_w23015_,
		_w23016_,
		_w23255_
	);
	LUT2 #(
		.INIT('h1)
	) name12744 (
		_w23017_,
		_w23018_,
		_w23256_
	);
	LUT2 #(
		.INIT('h1)
	) name12745 (
		_w23019_,
		_w23020_,
		_w23257_
	);
	LUT2 #(
		.INIT('h1)
	) name12746 (
		_w23021_,
		_w23022_,
		_w23258_
	);
	LUT2 #(
		.INIT('h1)
	) name12747 (
		_w23023_,
		_w23024_,
		_w23259_
	);
	LUT2 #(
		.INIT('h1)
	) name12748 (
		_w23025_,
		_w23026_,
		_w23260_
	);
	LUT2 #(
		.INIT('h1)
	) name12749 (
		_w23027_,
		_w23028_,
		_w23261_
	);
	LUT2 #(
		.INIT('h1)
	) name12750 (
		_w23029_,
		_w23030_,
		_w23262_
	);
	LUT2 #(
		.INIT('h1)
	) name12751 (
		_w23031_,
		_w23032_,
		_w23263_
	);
	LUT2 #(
		.INIT('h1)
	) name12752 (
		_w23033_,
		_w23034_,
		_w23264_
	);
	LUT2 #(
		.INIT('h1)
	) name12753 (
		_w23035_,
		_w23036_,
		_w23265_
	);
	LUT2 #(
		.INIT('h1)
	) name12754 (
		_w23037_,
		_w23038_,
		_w23266_
	);
	LUT2 #(
		.INIT('h1)
	) name12755 (
		_w23039_,
		_w23040_,
		_w23267_
	);
	LUT2 #(
		.INIT('h1)
	) name12756 (
		_w23041_,
		_w23042_,
		_w23268_
	);
	LUT2 #(
		.INIT('h1)
	) name12757 (
		_w23043_,
		_w23044_,
		_w23269_
	);
	LUT2 #(
		.INIT('h1)
	) name12758 (
		_w23045_,
		_w23046_,
		_w23270_
	);
	LUT2 #(
		.INIT('h1)
	) name12759 (
		_w23047_,
		_w23048_,
		_w23271_
	);
	LUT2 #(
		.INIT('h1)
	) name12760 (
		_w23049_,
		_w23050_,
		_w23272_
	);
	LUT2 #(
		.INIT('h1)
	) name12761 (
		_w23051_,
		_w23052_,
		_w23273_
	);
	LUT2 #(
		.INIT('h1)
	) name12762 (
		_w23053_,
		_w23054_,
		_w23274_
	);
	LUT2 #(
		.INIT('h1)
	) name12763 (
		_w23055_,
		_w23056_,
		_w23275_
	);
	LUT2 #(
		.INIT('h1)
	) name12764 (
		_w23057_,
		_w23058_,
		_w23276_
	);
	LUT2 #(
		.INIT('h1)
	) name12765 (
		_w23059_,
		_w23060_,
		_w23277_
	);
	LUT2 #(
		.INIT('h1)
	) name12766 (
		_w23061_,
		_w23062_,
		_w23278_
	);
	LUT2 #(
		.INIT('h1)
	) name12767 (
		_w23063_,
		_w23064_,
		_w23279_
	);
	LUT2 #(
		.INIT('h1)
	) name12768 (
		_w23065_,
		_w23066_,
		_w23280_
	);
	LUT2 #(
		.INIT('h1)
	) name12769 (
		_w23067_,
		_w23068_,
		_w23281_
	);
	LUT2 #(
		.INIT('h1)
	) name12770 (
		_w23069_,
		_w23070_,
		_w23282_
	);
	LUT2 #(
		.INIT('h1)
	) name12771 (
		_w23071_,
		_w23072_,
		_w23283_
	);
	LUT2 #(
		.INIT('h1)
	) name12772 (
		_w23073_,
		_w23074_,
		_w23284_
	);
	LUT2 #(
		.INIT('h1)
	) name12773 (
		_w23075_,
		_w23076_,
		_w23285_
	);
	LUT2 #(
		.INIT('h1)
	) name12774 (
		_w23077_,
		_w23078_,
		_w23286_
	);
	LUT2 #(
		.INIT('h1)
	) name12775 (
		_w23079_,
		_w23080_,
		_w23287_
	);
	LUT2 #(
		.INIT('h1)
	) name12776 (
		_w23081_,
		_w23082_,
		_w23288_
	);
	LUT2 #(
		.INIT('h1)
	) name12777 (
		_w23083_,
		_w23084_,
		_w23289_
	);
	LUT2 #(
		.INIT('h1)
	) name12778 (
		_w23085_,
		_w23086_,
		_w23290_
	);
	LUT2 #(
		.INIT('h1)
	) name12779 (
		_w23087_,
		_w23088_,
		_w23291_
	);
	LUT2 #(
		.INIT('h1)
	) name12780 (
		_w23089_,
		_w23090_,
		_w23292_
	);
	LUT2 #(
		.INIT('h1)
	) name12781 (
		_w23091_,
		_w23092_,
		_w23293_
	);
	LUT2 #(
		.INIT('h1)
	) name12782 (
		_w23093_,
		_w23094_,
		_w23294_
	);
	LUT2 #(
		.INIT('h1)
	) name12783 (
		_w23095_,
		_w23096_,
		_w23295_
	);
	LUT2 #(
		.INIT('h1)
	) name12784 (
		_w23097_,
		_w23098_,
		_w23296_
	);
	LUT2 #(
		.INIT('h1)
	) name12785 (
		_w23099_,
		_w23100_,
		_w23297_
	);
	LUT2 #(
		.INIT('h1)
	) name12786 (
		_w23101_,
		_w23102_,
		_w23298_
	);
	LUT2 #(
		.INIT('h1)
	) name12787 (
		_w23103_,
		_w23104_,
		_w23299_
	);
	LUT2 #(
		.INIT('h1)
	) name12788 (
		_w23105_,
		_w23106_,
		_w23300_
	);
	LUT2 #(
		.INIT('h1)
	) name12789 (
		_w23107_,
		_w23108_,
		_w23301_
	);
	LUT2 #(
		.INIT('h1)
	) name12790 (
		_w23109_,
		_w23110_,
		_w23302_
	);
	LUT2 #(
		.INIT('h1)
	) name12791 (
		_w23111_,
		_w23112_,
		_w23303_
	);
	LUT2 #(
		.INIT('h1)
	) name12792 (
		_w23113_,
		_w23114_,
		_w23304_
	);
	LUT2 #(
		.INIT('h1)
	) name12793 (
		_w23115_,
		_w23116_,
		_w23305_
	);
	LUT2 #(
		.INIT('h1)
	) name12794 (
		_w23117_,
		_w23118_,
		_w23306_
	);
	LUT2 #(
		.INIT('h1)
	) name12795 (
		_w23119_,
		_w23120_,
		_w23307_
	);
	LUT2 #(
		.INIT('h1)
	) name12796 (
		_w23121_,
		_w23122_,
		_w23308_
	);
	LUT2 #(
		.INIT('h1)
	) name12797 (
		_w23123_,
		_w23124_,
		_w23309_
	);
	LUT2 #(
		.INIT('h1)
	) name12798 (
		_w23125_,
		_w23126_,
		_w23310_
	);
	LUT2 #(
		.INIT('h1)
	) name12799 (
		_w23127_,
		_w23128_,
		_w23311_
	);
	LUT2 #(
		.INIT('h1)
	) name12800 (
		_w23129_,
		_w23130_,
		_w23312_
	);
	LUT2 #(
		.INIT('h1)
	) name12801 (
		_w23131_,
		_w23132_,
		_w23313_
	);
	LUT2 #(
		.INIT('h1)
	) name12802 (
		_w23133_,
		_w23134_,
		_w23314_
	);
	LUT2 #(
		.INIT('h1)
	) name12803 (
		_w23135_,
		_w23136_,
		_w23315_
	);
	LUT2 #(
		.INIT('h1)
	) name12804 (
		_w23137_,
		_w23138_,
		_w23316_
	);
	LUT2 #(
		.INIT('h1)
	) name12805 (
		_w23139_,
		_w23140_,
		_w23317_
	);
	LUT2 #(
		.INIT('h1)
	) name12806 (
		_w23141_,
		_w23142_,
		_w23318_
	);
	LUT2 #(
		.INIT('h1)
	) name12807 (
		_w23143_,
		_w23144_,
		_w23319_
	);
	LUT2 #(
		.INIT('h1)
	) name12808 (
		_w23145_,
		_w23146_,
		_w23320_
	);
	LUT2 #(
		.INIT('h1)
	) name12809 (
		_w23147_,
		_w23148_,
		_w23321_
	);
	LUT2 #(
		.INIT('h1)
	) name12810 (
		_w23149_,
		_w23150_,
		_w23322_
	);
	LUT2 #(
		.INIT('h1)
	) name12811 (
		_w23151_,
		_w23152_,
		_w23323_
	);
	LUT2 #(
		.INIT('h1)
	) name12812 (
		_w23153_,
		_w23154_,
		_w23324_
	);
	LUT2 #(
		.INIT('h1)
	) name12813 (
		_w23155_,
		_w23156_,
		_w23325_
	);
	LUT2 #(
		.INIT('h1)
	) name12814 (
		_w23157_,
		_w23158_,
		_w23326_
	);
	LUT2 #(
		.INIT('h1)
	) name12815 (
		_w23159_,
		_w23160_,
		_w23327_
	);
	LUT2 #(
		.INIT('h1)
	) name12816 (
		_w23161_,
		_w23162_,
		_w23328_
	);
	LUT2 #(
		.INIT('h1)
	) name12817 (
		_w23163_,
		_w23164_,
		_w23329_
	);
	LUT2 #(
		.INIT('h1)
	) name12818 (
		_w23165_,
		_w23166_,
		_w23330_
	);
	LUT2 #(
		.INIT('h1)
	) name12819 (
		_w23167_,
		_w23168_,
		_w23331_
	);
	LUT2 #(
		.INIT('h1)
	) name12820 (
		_w23169_,
		_w23170_,
		_w23332_
	);
	LUT2 #(
		.INIT('h1)
	) name12821 (
		_w23171_,
		_w23172_,
		_w23333_
	);
	LUT2 #(
		.INIT('h1)
	) name12822 (
		_w23173_,
		_w23174_,
		_w23334_
	);
	LUT2 #(
		.INIT('h1)
	) name12823 (
		_w23175_,
		_w23176_,
		_w23335_
	);
	LUT2 #(
		.INIT('h1)
	) name12824 (
		_w23177_,
		_w23178_,
		_w23336_
	);
	LUT2 #(
		.INIT('h1)
	) name12825 (
		_w23179_,
		_w23180_,
		_w23337_
	);
	LUT2 #(
		.INIT('h1)
	) name12826 (
		_w23181_,
		_w23182_,
		_w23338_
	);
	LUT2 #(
		.INIT('h1)
	) name12827 (
		_w23183_,
		_w23184_,
		_w23339_
	);
	LUT2 #(
		.INIT('h1)
	) name12828 (
		_w23185_,
		_w23186_,
		_w23340_
	);
	LUT2 #(
		.INIT('h1)
	) name12829 (
		_w23187_,
		_w23188_,
		_w23341_
	);
	LUT2 #(
		.INIT('h1)
	) name12830 (
		_w23189_,
		_w23190_,
		_w23342_
	);
	LUT2 #(
		.INIT('h1)
	) name12831 (
		_w23191_,
		_w23192_,
		_w23343_
	);
	LUT2 #(
		.INIT('h1)
	) name12832 (
		_w23193_,
		_w23194_,
		_w23344_
	);
	LUT2 #(
		.INIT('h1)
	) name12833 (
		_w23195_,
		_w23196_,
		_w23345_
	);
	LUT2 #(
		.INIT('h1)
	) name12834 (
		_w23197_,
		_w23198_,
		_w23346_
	);
	LUT2 #(
		.INIT('h1)
	) name12835 (
		_w23199_,
		_w23200_,
		_w23347_
	);
	LUT2 #(
		.INIT('h1)
	) name12836 (
		_w23201_,
		_w23202_,
		_w23348_
	);
	LUT2 #(
		.INIT('h1)
	) name12837 (
		_w23203_,
		_w23204_,
		_w23349_
	);
	LUT2 #(
		.INIT('h1)
	) name12838 (
		_w23205_,
		_w23206_,
		_w23350_
	);
	LUT2 #(
		.INIT('h1)
	) name12839 (
		_w23207_,
		_w23208_,
		_w23351_
	);
	LUT2 #(
		.INIT('h1)
	) name12840 (
		_w23209_,
		_w23210_,
		_w23352_
	);
	LUT2 #(
		.INIT('h1)
	) name12841 (
		_w23211_,
		_w23212_,
		_w23353_
	);
	LUT2 #(
		.INIT('h1)
	) name12842 (
		_w23213_,
		_w23214_,
		_w23354_
	);
	LUT2 #(
		.INIT('h1)
	) name12843 (
		_w23215_,
		_w23216_,
		_w23355_
	);
	LUT2 #(
		.INIT('h1)
	) name12844 (
		_w23217_,
		_w23218_,
		_w23356_
	);
	LUT2 #(
		.INIT('h1)
	) name12845 (
		_w23219_,
		_w23220_,
		_w23357_
	);
	LUT2 #(
		.INIT('h1)
	) name12846 (
		_w23221_,
		_w23222_,
		_w23358_
	);
	LUT2 #(
		.INIT('h1)
	) name12847 (
		_w23223_,
		_w23224_,
		_w23359_
	);
	LUT2 #(
		.INIT('h1)
	) name12848 (
		_w23225_,
		_w23226_,
		_w23360_
	);
	LUT2 #(
		.INIT('h1)
	) name12849 (
		_w23227_,
		_w23228_,
		_w23361_
	);
	LUT2 #(
		.INIT('h1)
	) name12850 (
		_w23229_,
		_w23230_,
		_w23362_
	);
	LUT2 #(
		.INIT('h1)
	) name12851 (
		_w23231_,
		_w23232_,
		_w23363_
	);
	LUT2 #(
		.INIT('h1)
	) name12852 (
		_w23233_,
		_w23234_,
		_w23364_
	);
	LUT2 #(
		.INIT('h1)
	) name12853 (
		_w23235_,
		_w23236_,
		_w23365_
	);
	LUT2 #(
		.INIT('h1)
	) name12854 (
		_w23237_,
		_w23238_,
		_w23366_
	);
	LUT2 #(
		.INIT('h8)
	) name12855 (
		_w23365_,
		_w23366_,
		_w23367_
	);
	LUT2 #(
		.INIT('h8)
	) name12856 (
		_w23363_,
		_w23364_,
		_w23368_
	);
	LUT2 #(
		.INIT('h8)
	) name12857 (
		_w23361_,
		_w23362_,
		_w23369_
	);
	LUT2 #(
		.INIT('h8)
	) name12858 (
		_w23359_,
		_w23360_,
		_w23370_
	);
	LUT2 #(
		.INIT('h8)
	) name12859 (
		_w23357_,
		_w23358_,
		_w23371_
	);
	LUT2 #(
		.INIT('h8)
	) name12860 (
		_w23355_,
		_w23356_,
		_w23372_
	);
	LUT2 #(
		.INIT('h8)
	) name12861 (
		_w23353_,
		_w23354_,
		_w23373_
	);
	LUT2 #(
		.INIT('h8)
	) name12862 (
		_w23351_,
		_w23352_,
		_w23374_
	);
	LUT2 #(
		.INIT('h8)
	) name12863 (
		_w23349_,
		_w23350_,
		_w23375_
	);
	LUT2 #(
		.INIT('h8)
	) name12864 (
		_w23347_,
		_w23348_,
		_w23376_
	);
	LUT2 #(
		.INIT('h8)
	) name12865 (
		_w23345_,
		_w23346_,
		_w23377_
	);
	LUT2 #(
		.INIT('h8)
	) name12866 (
		_w23343_,
		_w23344_,
		_w23378_
	);
	LUT2 #(
		.INIT('h8)
	) name12867 (
		_w23341_,
		_w23342_,
		_w23379_
	);
	LUT2 #(
		.INIT('h8)
	) name12868 (
		_w23339_,
		_w23340_,
		_w23380_
	);
	LUT2 #(
		.INIT('h8)
	) name12869 (
		_w23337_,
		_w23338_,
		_w23381_
	);
	LUT2 #(
		.INIT('h8)
	) name12870 (
		_w23335_,
		_w23336_,
		_w23382_
	);
	LUT2 #(
		.INIT('h8)
	) name12871 (
		_w23333_,
		_w23334_,
		_w23383_
	);
	LUT2 #(
		.INIT('h8)
	) name12872 (
		_w23331_,
		_w23332_,
		_w23384_
	);
	LUT2 #(
		.INIT('h8)
	) name12873 (
		_w23329_,
		_w23330_,
		_w23385_
	);
	LUT2 #(
		.INIT('h8)
	) name12874 (
		_w23327_,
		_w23328_,
		_w23386_
	);
	LUT2 #(
		.INIT('h8)
	) name12875 (
		_w23325_,
		_w23326_,
		_w23387_
	);
	LUT2 #(
		.INIT('h8)
	) name12876 (
		_w23323_,
		_w23324_,
		_w23388_
	);
	LUT2 #(
		.INIT('h8)
	) name12877 (
		_w23321_,
		_w23322_,
		_w23389_
	);
	LUT2 #(
		.INIT('h8)
	) name12878 (
		_w23319_,
		_w23320_,
		_w23390_
	);
	LUT2 #(
		.INIT('h8)
	) name12879 (
		_w23317_,
		_w23318_,
		_w23391_
	);
	LUT2 #(
		.INIT('h8)
	) name12880 (
		_w23315_,
		_w23316_,
		_w23392_
	);
	LUT2 #(
		.INIT('h8)
	) name12881 (
		_w23313_,
		_w23314_,
		_w23393_
	);
	LUT2 #(
		.INIT('h8)
	) name12882 (
		_w23311_,
		_w23312_,
		_w23394_
	);
	LUT2 #(
		.INIT('h8)
	) name12883 (
		_w23309_,
		_w23310_,
		_w23395_
	);
	LUT2 #(
		.INIT('h8)
	) name12884 (
		_w23307_,
		_w23308_,
		_w23396_
	);
	LUT2 #(
		.INIT('h8)
	) name12885 (
		_w23305_,
		_w23306_,
		_w23397_
	);
	LUT2 #(
		.INIT('h8)
	) name12886 (
		_w23303_,
		_w23304_,
		_w23398_
	);
	LUT2 #(
		.INIT('h8)
	) name12887 (
		_w23301_,
		_w23302_,
		_w23399_
	);
	LUT2 #(
		.INIT('h8)
	) name12888 (
		_w23299_,
		_w23300_,
		_w23400_
	);
	LUT2 #(
		.INIT('h8)
	) name12889 (
		_w23297_,
		_w23298_,
		_w23401_
	);
	LUT2 #(
		.INIT('h8)
	) name12890 (
		_w23295_,
		_w23296_,
		_w23402_
	);
	LUT2 #(
		.INIT('h8)
	) name12891 (
		_w23293_,
		_w23294_,
		_w23403_
	);
	LUT2 #(
		.INIT('h8)
	) name12892 (
		_w23291_,
		_w23292_,
		_w23404_
	);
	LUT2 #(
		.INIT('h8)
	) name12893 (
		_w23289_,
		_w23290_,
		_w23405_
	);
	LUT2 #(
		.INIT('h8)
	) name12894 (
		_w23287_,
		_w23288_,
		_w23406_
	);
	LUT2 #(
		.INIT('h8)
	) name12895 (
		_w23285_,
		_w23286_,
		_w23407_
	);
	LUT2 #(
		.INIT('h8)
	) name12896 (
		_w23283_,
		_w23284_,
		_w23408_
	);
	LUT2 #(
		.INIT('h8)
	) name12897 (
		_w23281_,
		_w23282_,
		_w23409_
	);
	LUT2 #(
		.INIT('h8)
	) name12898 (
		_w23279_,
		_w23280_,
		_w23410_
	);
	LUT2 #(
		.INIT('h8)
	) name12899 (
		_w23277_,
		_w23278_,
		_w23411_
	);
	LUT2 #(
		.INIT('h8)
	) name12900 (
		_w23275_,
		_w23276_,
		_w23412_
	);
	LUT2 #(
		.INIT('h8)
	) name12901 (
		_w23273_,
		_w23274_,
		_w23413_
	);
	LUT2 #(
		.INIT('h8)
	) name12902 (
		_w23271_,
		_w23272_,
		_w23414_
	);
	LUT2 #(
		.INIT('h8)
	) name12903 (
		_w23269_,
		_w23270_,
		_w23415_
	);
	LUT2 #(
		.INIT('h8)
	) name12904 (
		_w23267_,
		_w23268_,
		_w23416_
	);
	LUT2 #(
		.INIT('h8)
	) name12905 (
		_w23265_,
		_w23266_,
		_w23417_
	);
	LUT2 #(
		.INIT('h8)
	) name12906 (
		_w23263_,
		_w23264_,
		_w23418_
	);
	LUT2 #(
		.INIT('h8)
	) name12907 (
		_w23261_,
		_w23262_,
		_w23419_
	);
	LUT2 #(
		.INIT('h8)
	) name12908 (
		_w23259_,
		_w23260_,
		_w23420_
	);
	LUT2 #(
		.INIT('h8)
	) name12909 (
		_w23257_,
		_w23258_,
		_w23421_
	);
	LUT2 #(
		.INIT('h8)
	) name12910 (
		_w23255_,
		_w23256_,
		_w23422_
	);
	LUT2 #(
		.INIT('h8)
	) name12911 (
		_w23253_,
		_w23254_,
		_w23423_
	);
	LUT2 #(
		.INIT('h8)
	) name12912 (
		_w23251_,
		_w23252_,
		_w23424_
	);
	LUT2 #(
		.INIT('h8)
	) name12913 (
		_w23249_,
		_w23250_,
		_w23425_
	);
	LUT2 #(
		.INIT('h8)
	) name12914 (
		_w23247_,
		_w23248_,
		_w23426_
	);
	LUT2 #(
		.INIT('h8)
	) name12915 (
		_w23245_,
		_w23246_,
		_w23427_
	);
	LUT2 #(
		.INIT('h8)
	) name12916 (
		_w23243_,
		_w23244_,
		_w23428_
	);
	LUT2 #(
		.INIT('h8)
	) name12917 (
		_w23241_,
		_w23242_,
		_w23429_
	);
	LUT2 #(
		.INIT('h8)
	) name12918 (
		_w23239_,
		_w23240_,
		_w23430_
	);
	LUT2 #(
		.INIT('h8)
	) name12919 (
		_w23429_,
		_w23430_,
		_w23431_
	);
	LUT2 #(
		.INIT('h8)
	) name12920 (
		_w23427_,
		_w23428_,
		_w23432_
	);
	LUT2 #(
		.INIT('h8)
	) name12921 (
		_w23425_,
		_w23426_,
		_w23433_
	);
	LUT2 #(
		.INIT('h8)
	) name12922 (
		_w23423_,
		_w23424_,
		_w23434_
	);
	LUT2 #(
		.INIT('h8)
	) name12923 (
		_w23421_,
		_w23422_,
		_w23435_
	);
	LUT2 #(
		.INIT('h8)
	) name12924 (
		_w23419_,
		_w23420_,
		_w23436_
	);
	LUT2 #(
		.INIT('h8)
	) name12925 (
		_w23417_,
		_w23418_,
		_w23437_
	);
	LUT2 #(
		.INIT('h8)
	) name12926 (
		_w23415_,
		_w23416_,
		_w23438_
	);
	LUT2 #(
		.INIT('h8)
	) name12927 (
		_w23413_,
		_w23414_,
		_w23439_
	);
	LUT2 #(
		.INIT('h8)
	) name12928 (
		_w23411_,
		_w23412_,
		_w23440_
	);
	LUT2 #(
		.INIT('h8)
	) name12929 (
		_w23409_,
		_w23410_,
		_w23441_
	);
	LUT2 #(
		.INIT('h8)
	) name12930 (
		_w23407_,
		_w23408_,
		_w23442_
	);
	LUT2 #(
		.INIT('h8)
	) name12931 (
		_w23405_,
		_w23406_,
		_w23443_
	);
	LUT2 #(
		.INIT('h8)
	) name12932 (
		_w23403_,
		_w23404_,
		_w23444_
	);
	LUT2 #(
		.INIT('h8)
	) name12933 (
		_w23401_,
		_w23402_,
		_w23445_
	);
	LUT2 #(
		.INIT('h8)
	) name12934 (
		_w23399_,
		_w23400_,
		_w23446_
	);
	LUT2 #(
		.INIT('h8)
	) name12935 (
		_w23397_,
		_w23398_,
		_w23447_
	);
	LUT2 #(
		.INIT('h8)
	) name12936 (
		_w23395_,
		_w23396_,
		_w23448_
	);
	LUT2 #(
		.INIT('h8)
	) name12937 (
		_w23393_,
		_w23394_,
		_w23449_
	);
	LUT2 #(
		.INIT('h8)
	) name12938 (
		_w23391_,
		_w23392_,
		_w23450_
	);
	LUT2 #(
		.INIT('h8)
	) name12939 (
		_w23389_,
		_w23390_,
		_w23451_
	);
	LUT2 #(
		.INIT('h8)
	) name12940 (
		_w23387_,
		_w23388_,
		_w23452_
	);
	LUT2 #(
		.INIT('h8)
	) name12941 (
		_w23385_,
		_w23386_,
		_w23453_
	);
	LUT2 #(
		.INIT('h8)
	) name12942 (
		_w23383_,
		_w23384_,
		_w23454_
	);
	LUT2 #(
		.INIT('h8)
	) name12943 (
		_w23381_,
		_w23382_,
		_w23455_
	);
	LUT2 #(
		.INIT('h8)
	) name12944 (
		_w23379_,
		_w23380_,
		_w23456_
	);
	LUT2 #(
		.INIT('h8)
	) name12945 (
		_w23377_,
		_w23378_,
		_w23457_
	);
	LUT2 #(
		.INIT('h8)
	) name12946 (
		_w23375_,
		_w23376_,
		_w23458_
	);
	LUT2 #(
		.INIT('h8)
	) name12947 (
		_w23373_,
		_w23374_,
		_w23459_
	);
	LUT2 #(
		.INIT('h8)
	) name12948 (
		_w23371_,
		_w23372_,
		_w23460_
	);
	LUT2 #(
		.INIT('h8)
	) name12949 (
		_w23369_,
		_w23370_,
		_w23461_
	);
	LUT2 #(
		.INIT('h8)
	) name12950 (
		_w23367_,
		_w23368_,
		_w23462_
	);
	LUT2 #(
		.INIT('h8)
	) name12951 (
		_w23461_,
		_w23462_,
		_w23463_
	);
	LUT2 #(
		.INIT('h8)
	) name12952 (
		_w23459_,
		_w23460_,
		_w23464_
	);
	LUT2 #(
		.INIT('h8)
	) name12953 (
		_w23457_,
		_w23458_,
		_w23465_
	);
	LUT2 #(
		.INIT('h8)
	) name12954 (
		_w23455_,
		_w23456_,
		_w23466_
	);
	LUT2 #(
		.INIT('h8)
	) name12955 (
		_w23453_,
		_w23454_,
		_w23467_
	);
	LUT2 #(
		.INIT('h8)
	) name12956 (
		_w23451_,
		_w23452_,
		_w23468_
	);
	LUT2 #(
		.INIT('h8)
	) name12957 (
		_w23449_,
		_w23450_,
		_w23469_
	);
	LUT2 #(
		.INIT('h8)
	) name12958 (
		_w23447_,
		_w23448_,
		_w23470_
	);
	LUT2 #(
		.INIT('h8)
	) name12959 (
		_w23445_,
		_w23446_,
		_w23471_
	);
	LUT2 #(
		.INIT('h8)
	) name12960 (
		_w23443_,
		_w23444_,
		_w23472_
	);
	LUT2 #(
		.INIT('h8)
	) name12961 (
		_w23441_,
		_w23442_,
		_w23473_
	);
	LUT2 #(
		.INIT('h8)
	) name12962 (
		_w23439_,
		_w23440_,
		_w23474_
	);
	LUT2 #(
		.INIT('h8)
	) name12963 (
		_w23437_,
		_w23438_,
		_w23475_
	);
	LUT2 #(
		.INIT('h8)
	) name12964 (
		_w23435_,
		_w23436_,
		_w23476_
	);
	LUT2 #(
		.INIT('h8)
	) name12965 (
		_w23433_,
		_w23434_,
		_w23477_
	);
	LUT2 #(
		.INIT('h8)
	) name12966 (
		_w23431_,
		_w23432_,
		_w23478_
	);
	LUT2 #(
		.INIT('h8)
	) name12967 (
		_w23477_,
		_w23478_,
		_w23479_
	);
	LUT2 #(
		.INIT('h8)
	) name12968 (
		_w23475_,
		_w23476_,
		_w23480_
	);
	LUT2 #(
		.INIT('h8)
	) name12969 (
		_w23473_,
		_w23474_,
		_w23481_
	);
	LUT2 #(
		.INIT('h8)
	) name12970 (
		_w23471_,
		_w23472_,
		_w23482_
	);
	LUT2 #(
		.INIT('h8)
	) name12971 (
		_w23469_,
		_w23470_,
		_w23483_
	);
	LUT2 #(
		.INIT('h8)
	) name12972 (
		_w23467_,
		_w23468_,
		_w23484_
	);
	LUT2 #(
		.INIT('h8)
	) name12973 (
		_w23465_,
		_w23466_,
		_w23485_
	);
	LUT2 #(
		.INIT('h8)
	) name12974 (
		_w23463_,
		_w23464_,
		_w23486_
	);
	LUT2 #(
		.INIT('h8)
	) name12975 (
		_w23485_,
		_w23486_,
		_w23487_
	);
	LUT2 #(
		.INIT('h8)
	) name12976 (
		_w23483_,
		_w23484_,
		_w23488_
	);
	LUT2 #(
		.INIT('h8)
	) name12977 (
		_w23481_,
		_w23482_,
		_w23489_
	);
	LUT2 #(
		.INIT('h8)
	) name12978 (
		_w23479_,
		_w23480_,
		_w23490_
	);
	LUT2 #(
		.INIT('h8)
	) name12979 (
		_w23489_,
		_w23490_,
		_w23491_
	);
	LUT2 #(
		.INIT('h8)
	) name12980 (
		_w23487_,
		_w23488_,
		_w23492_
	);
	LUT2 #(
		.INIT('h8)
	) name12981 (
		_w23491_,
		_w23492_,
		_w23493_
	);
	LUT2 #(
		.INIT('h1)
	) name12982 (
		wb_rst_i_pad,
		_w23493_,
		_w23494_
	);
	LUT2 #(
		.INIT('h1)
	) name12983 (
		_w22944_,
		_w23494_,
		_w23495_
	);
	LUT2 #(
		.INIT('h8)
	) name12984 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		_w22959_,
		_w23496_
	);
	LUT2 #(
		.INIT('h4)
	) name12985 (
		\wb_adr_i[3]_pad ,
		\wb_adr_i[4]_pad ,
		_w23497_
	);
	LUT2 #(
		.INIT('h4)
	) name12986 (
		\wb_adr_i[5]_pad ,
		_w23497_,
		_w23498_
	);
	LUT2 #(
		.INIT('h8)
	) name12987 (
		_w22951_,
		_w23498_,
		_w23499_
	);
	LUT2 #(
		.INIT('h8)
	) name12988 (
		\ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 ,
		_w23499_,
		_w23500_
	);
	LUT2 #(
		.INIT('h8)
	) name12989 (
		_w22955_,
		_w22958_,
		_w23501_
	);
	LUT2 #(
		.INIT('h8)
	) name12990 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		_w23501_,
		_w23502_
	);
	LUT2 #(
		.INIT('h2)
	) name12991 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		_w23503_
	);
	LUT2 #(
		.INIT('h8)
	) name12992 (
		_w22950_,
		_w23503_,
		_w23504_
	);
	LUT2 #(
		.INIT('h8)
	) name12993 (
		\wb_adr_i[3]_pad ,
		_w22948_,
		_w23505_
	);
	LUT2 #(
		.INIT('h8)
	) name12994 (
		\wb_adr_i[5]_pad ,
		_w23505_,
		_w23506_
	);
	LUT2 #(
		.INIT('h8)
	) name12995 (
		_w23504_,
		_w23506_,
		_w23507_
	);
	LUT2 #(
		.INIT('h8)
	) name12996 (
		\ethreg1_MIIRX_DATA_DataOut_reg[12]/NET0131 ,
		_w23507_,
		_w23508_
	);
	LUT2 #(
		.INIT('h8)
	) name12997 (
		\ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 ,
		_w22952_,
		_w23509_
	);
	LUT2 #(
		.INIT('h8)
	) name12998 (
		\ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 ,
		_w22956_,
		_w23510_
	);
	LUT2 #(
		.INIT('h4)
	) name12999 (
		\wb_adr_i[3]_pad ,
		_w22948_,
		_w23511_
	);
	LUT2 #(
		.INIT('h8)
	) name13000 (
		\wb_adr_i[5]_pad ,
		_w23511_,
		_w23512_
	);
	LUT2 #(
		.INIT('h8)
	) name13001 (
		_w23504_,
		_w23512_,
		_w23513_
	);
	LUT2 #(
		.INIT('h8)
	) name13002 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w23513_,
		_w23514_
	);
	LUT2 #(
		.INIT('h8)
	) name13003 (
		\ethreg1_PACKETLEN_1_DataOut_reg[4]/NET0131 ,
		_w22966_,
		_w23515_
	);
	LUT2 #(
		.INIT('h4)
	) name13004 (
		\wb_adr_i[5]_pad ,
		_w23511_,
		_w23516_
	);
	LUT2 #(
		.INIT('h1)
	) name13005 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[6]_pad ,
		_w23517_
	);
	LUT2 #(
		.INIT('h8)
	) name13006 (
		_w22950_,
		_w23517_,
		_w23518_
	);
	LUT2 #(
		.INIT('h8)
	) name13007 (
		_w23516_,
		_w23518_,
		_w23519_
	);
	LUT2 #(
		.INIT('h8)
	) name13008 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w23519_,
		_w23520_
	);
	LUT2 #(
		.INIT('h8)
	) name13009 (
		_w22954_,
		_w23503_,
		_w23521_
	);
	LUT2 #(
		.INIT('h8)
	) name13010 (
		_w23512_,
		_w23521_,
		_w23522_
	);
	LUT2 #(
		.INIT('h8)
	) name13011 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 ,
		_w23522_,
		_w23523_
	);
	LUT2 #(
		.INIT('h1)
	) name13012 (
		_w23496_,
		_w23500_,
		_w23524_
	);
	LUT2 #(
		.INIT('h1)
	) name13013 (
		_w23502_,
		_w23508_,
		_w23525_
	);
	LUT2 #(
		.INIT('h1)
	) name13014 (
		_w23509_,
		_w23510_,
		_w23526_
	);
	LUT2 #(
		.INIT('h1)
	) name13015 (
		_w23514_,
		_w23520_,
		_w23527_
	);
	LUT2 #(
		.INIT('h4)
	) name13016 (
		_w23523_,
		_w23527_,
		_w23528_
	);
	LUT2 #(
		.INIT('h8)
	) name13017 (
		_w23525_,
		_w23526_,
		_w23529_
	);
	LUT2 #(
		.INIT('h8)
	) name13018 (
		_w22944_,
		_w23524_,
		_w23530_
	);
	LUT2 #(
		.INIT('h8)
	) name13019 (
		_w23529_,
		_w23530_,
		_w23531_
	);
	LUT2 #(
		.INIT('h4)
	) name13020 (
		_w23515_,
		_w23528_,
		_w23532_
	);
	LUT2 #(
		.INIT('h8)
	) name13021 (
		_w23531_,
		_w23532_,
		_w23533_
	);
	LUT2 #(
		.INIT('h1)
	) name13022 (
		_w23495_,
		_w23533_,
		_w23534_
	);
	LUT2 #(
		.INIT('h2)
	) name13023 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w12657_,
		_w23535_
	);
	LUT2 #(
		.INIT('h4)
	) name13024 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w16763_,
		_w23536_
	);
	LUT2 #(
		.INIT('h2)
	) name13025 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w23536_,
		_w23537_
	);
	LUT2 #(
		.INIT('h2)
	) name13026 (
		_w16762_,
		_w16764_,
		_w23538_
	);
	LUT2 #(
		.INIT('h4)
	) name13027 (
		_w23537_,
		_w23538_,
		_w23539_
	);
	LUT2 #(
		.INIT('h1)
	) name13028 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w13485_,
		_w23540_
	);
	LUT2 #(
		.INIT('h2)
	) name13029 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w23540_,
		_w23541_
	);
	LUT2 #(
		.INIT('h1)
	) name13030 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w23541_,
		_w23542_
	);
	LUT2 #(
		.INIT('h2)
	) name13031 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w23542_,
		_w23543_
	);
	LUT2 #(
		.INIT('h4)
	) name13032 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w23542_,
		_w23544_
	);
	LUT2 #(
		.INIT('h1)
	) name13033 (
		_w16762_,
		_w23543_,
		_w23545_
	);
	LUT2 #(
		.INIT('h4)
	) name13034 (
		_w23544_,
		_w23545_,
		_w23546_
	);
	LUT2 #(
		.INIT('h2)
	) name13035 (
		_w13500_,
		_w23539_,
		_w23547_
	);
	LUT2 #(
		.INIT('h4)
	) name13036 (
		_w23546_,
		_w23547_,
		_w23548_
	);
	LUT2 #(
		.INIT('h1)
	) name13037 (
		_w23535_,
		_w23548_,
		_w23549_
	);
	LUT2 #(
		.INIT('h1)
	) name13038 (
		_w12656_,
		_w23549_,
		_w23550_
	);
	LUT2 #(
		.INIT('h1)
	) name13039 (
		_w21384_,
		_w23550_,
		_w23551_
	);
	LUT2 #(
		.INIT('h2)
	) name13040 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w12657_,
		_w23552_
	);
	LUT2 #(
		.INIT('h4)
	) name13041 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w13481_,
		_w23553_
	);
	LUT2 #(
		.INIT('h2)
	) name13042 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w23553_,
		_w23554_
	);
	LUT2 #(
		.INIT('h1)
	) name13043 (
		_w13483_,
		_w23554_,
		_w23555_
	);
	LUT2 #(
		.INIT('h2)
	) name13044 (
		_w16748_,
		_w23555_,
		_w23556_
	);
	LUT2 #(
		.INIT('h4)
	) name13045 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w16757_,
		_w23557_
	);
	LUT2 #(
		.INIT('h4)
	) name13046 (
		_w16757_,
		_w23555_,
		_w23558_
	);
	LUT2 #(
		.INIT('h2)
	) name13047 (
		_w16756_,
		_w23557_,
		_w23559_
	);
	LUT2 #(
		.INIT('h4)
	) name13048 (
		_w23558_,
		_w23559_,
		_w23560_
	);
	LUT2 #(
		.INIT('h4)
	) name13049 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w16753_,
		_w23561_
	);
	LUT2 #(
		.INIT('h8)
	) name13050 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w23561_,
		_w23562_
	);
	LUT2 #(
		.INIT('h4)
	) name13051 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		_w23562_,
		_w23563_
	);
	LUT2 #(
		.INIT('h8)
	) name13052 (
		_w16763_,
		_w23553_,
		_w23564_
	);
	LUT2 #(
		.INIT('h1)
	) name13053 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w23564_,
		_w23565_
	);
	LUT2 #(
		.INIT('h2)
	) name13054 (
		_w16762_,
		_w23565_,
		_w23566_
	);
	LUT2 #(
		.INIT('h4)
	) name13055 (
		_w23563_,
		_w23566_,
		_w23567_
	);
	LUT2 #(
		.INIT('h1)
	) name13056 (
		\wishbone_TxLength_reg[6]/NET0131 ,
		_w23561_,
		_w23568_
	);
	LUT2 #(
		.INIT('h2)
	) name13057 (
		_w16750_,
		_w23562_,
		_w23569_
	);
	LUT2 #(
		.INIT('h4)
	) name13058 (
		_w23568_,
		_w23569_,
		_w23570_
	);
	LUT2 #(
		.INIT('h1)
	) name13059 (
		_w23556_,
		_w23560_,
		_w23571_
	);
	LUT2 #(
		.INIT('h1)
	) name13060 (
		_w23567_,
		_w23570_,
		_w23572_
	);
	LUT2 #(
		.INIT('h8)
	) name13061 (
		_w23571_,
		_w23572_,
		_w23573_
	);
	LUT2 #(
		.INIT('h2)
	) name13062 (
		_w13500_,
		_w23573_,
		_w23574_
	);
	LUT2 #(
		.INIT('h1)
	) name13063 (
		_w23552_,
		_w23574_,
		_w23575_
	);
	LUT2 #(
		.INIT('h1)
	) name13064 (
		_w12656_,
		_w23575_,
		_w23576_
	);
	LUT2 #(
		.INIT('h1)
	) name13065 (
		_w22933_,
		_w23576_,
		_w23577_
	);
	LUT2 #(
		.INIT('h2)
	) name13066 (
		\wishbone_TxPointerLSB_reg[1]/NET0131 ,
		_w17883_,
		_w23578_
	);
	LUT2 #(
		.INIT('h8)
	) name13067 (
		_w16210_,
		_w17883_,
		_w23579_
	);
	LUT2 #(
		.INIT('h1)
	) name13068 (
		_w23578_,
		_w23579_,
		_w23580_
	);
	LUT2 #(
		.INIT('h1)
	) name13069 (
		_w12657_,
		_w17883_,
		_w23581_
	);
	LUT2 #(
		.INIT('h8)
	) name13070 (
		\wishbone_TxPointerLSB_rst_reg[0]/NET0131 ,
		_w23581_,
		_w23582_
	);
	LUT2 #(
		.INIT('h8)
	) name13071 (
		\wishbone_bd_ram_mem0_reg[185][0]/P0001 ,
		_w12940_,
		_w23583_
	);
	LUT2 #(
		.INIT('h8)
	) name13072 (
		\wishbone_bd_ram_mem0_reg[130][0]/P0001 ,
		_w12914_,
		_w23584_
	);
	LUT2 #(
		.INIT('h8)
	) name13073 (
		\wishbone_bd_ram_mem0_reg[235][0]/P0001 ,
		_w12696_,
		_w23585_
	);
	LUT2 #(
		.INIT('h8)
	) name13074 (
		\wishbone_bd_ram_mem0_reg[21][0]/P0001 ,
		_w12906_,
		_w23586_
	);
	LUT2 #(
		.INIT('h8)
	) name13075 (
		\wishbone_bd_ram_mem0_reg[183][0]/P0001 ,
		_w12787_,
		_w23587_
	);
	LUT2 #(
		.INIT('h8)
	) name13076 (
		\wishbone_bd_ram_mem0_reg[60][0]/P0001 ,
		_w13204_,
		_w23588_
	);
	LUT2 #(
		.INIT('h8)
	) name13077 (
		\wishbone_bd_ram_mem0_reg[86][0]/P0001 ,
		_w12735_,
		_w23589_
	);
	LUT2 #(
		.INIT('h8)
	) name13078 (
		\wishbone_bd_ram_mem0_reg[6][0]/P0001 ,
		_w12968_,
		_w23590_
	);
	LUT2 #(
		.INIT('h8)
	) name13079 (
		\wishbone_bd_ram_mem0_reg[197][0]/P0001 ,
		_w12834_,
		_w23591_
	);
	LUT2 #(
		.INIT('h8)
	) name13080 (
		\wishbone_bd_ram_mem0_reg[122][0]/P0001 ,
		_w13130_,
		_w23592_
	);
	LUT2 #(
		.INIT('h8)
	) name13081 (
		\wishbone_bd_ram_mem0_reg[244][0]/P0001 ,
		_w12747_,
		_w23593_
	);
	LUT2 #(
		.INIT('h8)
	) name13082 (
		\wishbone_bd_ram_mem0_reg[93][0]/P0001 ,
		_w13016_,
		_w23594_
	);
	LUT2 #(
		.INIT('h8)
	) name13083 (
		\wishbone_bd_ram_mem0_reg[175][0]/P0001 ,
		_w13126_,
		_w23595_
	);
	LUT2 #(
		.INIT('h8)
	) name13084 (
		\wishbone_bd_ram_mem0_reg[36][0]/P0001 ,
		_w12800_,
		_w23596_
	);
	LUT2 #(
		.INIT('h8)
	) name13085 (
		\wishbone_bd_ram_mem0_reg[247][0]/P0001 ,
		_w12818_,
		_w23597_
	);
	LUT2 #(
		.INIT('h8)
	) name13086 (
		\wishbone_bd_ram_mem0_reg[215][0]/P0001 ,
		_w12974_,
		_w23598_
	);
	LUT2 #(
		.INIT('h8)
	) name13087 (
		\wishbone_bd_ram_mem0_reg[223][0]/P0001 ,
		_w12838_,
		_w23599_
	);
	LUT2 #(
		.INIT('h8)
	) name13088 (
		\wishbone_bd_ram_mem0_reg[66][0]/P0001 ,
		_w12824_,
		_w23600_
	);
	LUT2 #(
		.INIT('h8)
	) name13089 (
		\wishbone_bd_ram_mem0_reg[12][0]/P0001 ,
		_w13118_,
		_w23601_
	);
	LUT2 #(
		.INIT('h8)
	) name13090 (
		\wishbone_bd_ram_mem0_reg[211][0]/P0001 ,
		_w13166_,
		_w23602_
	);
	LUT2 #(
		.INIT('h8)
	) name13091 (
		\wishbone_bd_ram_mem0_reg[68][0]/P0001 ,
		_w12946_,
		_w23603_
	);
	LUT2 #(
		.INIT('h8)
	) name13092 (
		\wishbone_bd_ram_mem0_reg[31][0]/P0001 ,
		_w13198_,
		_w23604_
	);
	LUT2 #(
		.INIT('h8)
	) name13093 (
		\wishbone_bd_ram_mem0_reg[209][0]/P0001 ,
		_w13152_,
		_w23605_
	);
	LUT2 #(
		.INIT('h8)
	) name13094 (
		\wishbone_bd_ram_mem0_reg[179][0]/P0001 ,
		_w13050_,
		_w23606_
	);
	LUT2 #(
		.INIT('h8)
	) name13095 (
		\wishbone_bd_ram_mem0_reg[237][0]/P0001 ,
		_w12990_,
		_w23607_
	);
	LUT2 #(
		.INIT('h8)
	) name13096 (
		\wishbone_bd_ram_mem0_reg[135][0]/P0001 ,
		_w13124_,
		_w23608_
	);
	LUT2 #(
		.INIT('h8)
	) name13097 (
		\wishbone_bd_ram_mem0_reg[192][0]/P0001 ,
		_w12938_,
		_w23609_
	);
	LUT2 #(
		.INIT('h8)
	) name13098 (
		\wishbone_bd_ram_mem0_reg[198][0]/P0001 ,
		_w12832_,
		_w23610_
	);
	LUT2 #(
		.INIT('h8)
	) name13099 (
		\wishbone_bd_ram_mem0_reg[91][0]/P0001 ,
		_w13074_,
		_w23611_
	);
	LUT2 #(
		.INIT('h8)
	) name13100 (
		\wishbone_bd_ram_mem0_reg[133][0]/P0001 ,
		_w12761_,
		_w23612_
	);
	LUT2 #(
		.INIT('h8)
	) name13101 (
		\wishbone_bd_ram_mem0_reg[234][0]/P0001 ,
		_w13214_,
		_w23613_
	);
	LUT2 #(
		.INIT('h8)
	) name13102 (
		\wishbone_bd_ram_mem0_reg[42][0]/P0001 ,
		_w12842_,
		_w23614_
	);
	LUT2 #(
		.INIT('h8)
	) name13103 (
		\wishbone_bd_ram_mem0_reg[87][0]/P0001 ,
		_w13154_,
		_w23615_
	);
	LUT2 #(
		.INIT('h8)
	) name13104 (
		\wishbone_bd_ram_mem0_reg[82][0]/P0001 ,
		_w12942_,
		_w23616_
	);
	LUT2 #(
		.INIT('h8)
	) name13105 (
		\wishbone_bd_ram_mem0_reg[11][0]/P0001 ,
		_w13194_,
		_w23617_
	);
	LUT2 #(
		.INIT('h8)
	) name13106 (
		\wishbone_bd_ram_mem0_reg[81][0]/P0001 ,
		_w12950_,
		_w23618_
	);
	LUT2 #(
		.INIT('h8)
	) name13107 (
		\wishbone_bd_ram_mem0_reg[144][0]/P0001 ,
		_w12756_,
		_w23619_
	);
	LUT2 #(
		.INIT('h8)
	) name13108 (
		\wishbone_bd_ram_mem0_reg[188][0]/P0001 ,
		_w12948_,
		_w23620_
	);
	LUT2 #(
		.INIT('h8)
	) name13109 (
		\wishbone_bd_ram_mem0_reg[249][0]/P0001 ,
		_w12900_,
		_w23621_
	);
	LUT2 #(
		.INIT('h8)
	) name13110 (
		\wishbone_bd_ram_mem0_reg[251][0]/P0001 ,
		_w13054_,
		_w23622_
	);
	LUT2 #(
		.INIT('h8)
	) name13111 (
		\wishbone_bd_ram_mem0_reg[18][0]/P0001 ,
		_w12679_,
		_w23623_
	);
	LUT2 #(
		.INIT('h8)
	) name13112 (
		\wishbone_bd_ram_mem0_reg[111][0]/P0001 ,
		_w12744_,
		_w23624_
	);
	LUT2 #(
		.INIT('h8)
	) name13113 (
		\wishbone_bd_ram_mem0_reg[242][0]/P0001 ,
		_w12932_,
		_w23625_
	);
	LUT2 #(
		.INIT('h8)
	) name13114 (
		\wishbone_bd_ram_mem0_reg[78][0]/P0001 ,
		_w12874_,
		_w23626_
	);
	LUT2 #(
		.INIT('h8)
	) name13115 (
		\wishbone_bd_ram_mem0_reg[160][0]/P0001 ,
		_w12872_,
		_w23627_
	);
	LUT2 #(
		.INIT('h8)
	) name13116 (
		\wishbone_bd_ram_mem0_reg[32][0]/P0001 ,
		_w13120_,
		_w23628_
	);
	LUT2 #(
		.INIT('h8)
	) name13117 (
		\wishbone_bd_ram_mem0_reg[169][0]/P0001 ,
		_w12722_,
		_w23629_
	);
	LUT2 #(
		.INIT('h8)
	) name13118 (
		\wishbone_bd_ram_mem0_reg[216][0]/P0001 ,
		_w13028_,
		_w23630_
	);
	LUT2 #(
		.INIT('h8)
	) name13119 (
		\wishbone_bd_ram_mem0_reg[199][0]/P0001 ,
		_w12768_,
		_w23631_
	);
	LUT2 #(
		.INIT('h8)
	) name13120 (
		\wishbone_bd_ram_mem0_reg[250][0]/P0001 ,
		_w13128_,
		_w23632_
	);
	LUT2 #(
		.INIT('h8)
	) name13121 (
		\wishbone_bd_ram_mem0_reg[5][0]/P0001 ,
		_w12878_,
		_w23633_
	);
	LUT2 #(
		.INIT('h8)
	) name13122 (
		\wishbone_bd_ram_mem0_reg[9][0]/P0001 ,
		_w12808_,
		_w23634_
	);
	LUT2 #(
		.INIT('h8)
	) name13123 (
		\wishbone_bd_ram_mem0_reg[195][0]/P0001 ,
		_w13144_,
		_w23635_
	);
	LUT2 #(
		.INIT('h8)
	) name13124 (
		\wishbone_bd_ram_mem0_reg[226][0]/P0001 ,
		_w13138_,
		_w23636_
	);
	LUT2 #(
		.INIT('h8)
	) name13125 (
		\wishbone_bd_ram_mem0_reg[24][0]/P0001 ,
		_w13084_,
		_w23637_
	);
	LUT2 #(
		.INIT('h8)
	) name13126 (
		\wishbone_bd_ram_mem0_reg[8][0]/P0001 ,
		_w12920_,
		_w23638_
	);
	LUT2 #(
		.INIT('h8)
	) name13127 (
		\wishbone_bd_ram_mem0_reg[64][0]/P0001 ,
		_w12976_,
		_w23639_
	);
	LUT2 #(
		.INIT('h8)
	) name13128 (
		\wishbone_bd_ram_mem0_reg[222][0]/P0001 ,
		_w13094_,
		_w23640_
	);
	LUT2 #(
		.INIT('h8)
	) name13129 (
		\wishbone_bd_ram_mem0_reg[10][0]/P0001 ,
		_w13172_,
		_w23641_
	);
	LUT2 #(
		.INIT('h8)
	) name13130 (
		\wishbone_bd_ram_mem0_reg[28][0]/P0001 ,
		_w13170_,
		_w23642_
	);
	LUT2 #(
		.INIT('h8)
	) name13131 (
		\wishbone_bd_ram_mem0_reg[214][0]/P0001 ,
		_w12984_,
		_w23643_
	);
	LUT2 #(
		.INIT('h8)
	) name13132 (
		\wishbone_bd_ram_mem0_reg[203][0]/P0001 ,
		_w13158_,
		_w23644_
	);
	LUT2 #(
		.INIT('h8)
	) name13133 (
		\wishbone_bd_ram_mem0_reg[232][0]/P0001 ,
		_w12758_,
		_w23645_
	);
	LUT2 #(
		.INIT('h8)
	) name13134 (
		\wishbone_bd_ram_mem0_reg[140][0]/P0001 ,
		_w12894_,
		_w23646_
	);
	LUT2 #(
		.INIT('h8)
	) name13135 (
		\wishbone_bd_ram_mem0_reg[228][0]/P0001 ,
		_w12765_,
		_w23647_
	);
	LUT2 #(
		.INIT('h8)
	) name13136 (
		\wishbone_bd_ram_mem0_reg[0][0]/P0001 ,
		_w12717_,
		_w23648_
	);
	LUT2 #(
		.INIT('h8)
	) name13137 (
		\wishbone_bd_ram_mem0_reg[184][0]/P0001 ,
		_w13062_,
		_w23649_
	);
	LUT2 #(
		.INIT('h8)
	) name13138 (
		\wishbone_bd_ram_mem0_reg[30][0]/P0001 ,
		_w13104_,
		_w23650_
	);
	LUT2 #(
		.INIT('h8)
	) name13139 (
		\wishbone_bd_ram_mem0_reg[114][0]/P0001 ,
		_w13202_,
		_w23651_
	);
	LUT2 #(
		.INIT('h8)
	) name13140 (
		\wishbone_bd_ram_mem0_reg[79][0]/P0001 ,
		_w13212_,
		_w23652_
	);
	LUT2 #(
		.INIT('h8)
	) name13141 (
		\wishbone_bd_ram_mem0_reg[151][0]/P0001 ,
		_w13142_,
		_w23653_
	);
	LUT2 #(
		.INIT('h8)
	) name13142 (
		\wishbone_bd_ram_mem0_reg[112][0]/P0001 ,
		_w12733_,
		_w23654_
	);
	LUT2 #(
		.INIT('h8)
	) name13143 (
		\wishbone_bd_ram_mem0_reg[126][0]/P0001 ,
		_w13218_,
		_w23655_
	);
	LUT2 #(
		.INIT('h8)
	) name13144 (
		\wishbone_bd_ram_mem0_reg[47][0]/P0001 ,
		_w12904_,
		_w23656_
	);
	LUT2 #(
		.INIT('h8)
	) name13145 (
		\wishbone_bd_ram_mem0_reg[58][0]/P0001 ,
		_w13070_,
		_w23657_
	);
	LUT2 #(
		.INIT('h8)
	) name13146 (
		\wishbone_bd_ram_mem0_reg[196][0]/P0001 ,
		_w13090_,
		_w23658_
	);
	LUT2 #(
		.INIT('h8)
	) name13147 (
		\wishbone_bd_ram_mem0_reg[103][0]/P0001 ,
		_w12846_,
		_w23659_
	);
	LUT2 #(
		.INIT('h8)
	) name13148 (
		\wishbone_bd_ram_mem0_reg[7][0]/P0001 ,
		_w12728_,
		_w23660_
	);
	LUT2 #(
		.INIT('h8)
	) name13149 (
		\wishbone_bd_ram_mem0_reg[45][0]/P0001 ,
		_w12908_,
		_w23661_
	);
	LUT2 #(
		.INIT('h8)
	) name13150 (
		\wishbone_bd_ram_mem0_reg[39][0]/P0001 ,
		_w13018_,
		_w23662_
	);
	LUT2 #(
		.INIT('h8)
	) name13151 (
		\wishbone_bd_ram_mem0_reg[159][0]/P0001 ,
		_w12774_,
		_w23663_
	);
	LUT2 #(
		.INIT('h8)
	) name13152 (
		\wishbone_bd_ram_mem0_reg[25][0]/P0001 ,
		_w13108_,
		_w23664_
	);
	LUT2 #(
		.INIT('h8)
	) name13153 (
		\wishbone_bd_ram_mem0_reg[26][0]/P0001 ,
		_w12699_,
		_w23665_
	);
	LUT2 #(
		.INIT('h8)
	) name13154 (
		\wishbone_bd_ram_mem0_reg[146][0]/P0001 ,
		_w13060_,
		_w23666_
	);
	LUT2 #(
		.INIT('h8)
	) name13155 (
		\wishbone_bd_ram_mem0_reg[153][0]/P0001 ,
		_w12890_,
		_w23667_
	);
	LUT2 #(
		.INIT('h8)
	) name13156 (
		\wishbone_bd_ram_mem0_reg[174][0]/P0001 ,
		_w12972_,
		_w23668_
	);
	LUT2 #(
		.INIT('h8)
	) name13157 (
		\wishbone_bd_ram_mem0_reg[166][0]/P0001 ,
		_w13040_,
		_w23669_
	);
	LUT2 #(
		.INIT('h8)
	) name13158 (
		\wishbone_bd_ram_mem0_reg[150][0]/P0001 ,
		_w13136_,
		_w23670_
	);
	LUT2 #(
		.INIT('h8)
	) name13159 (
		\wishbone_bd_ram_mem0_reg[101][0]/P0001 ,
		_w13192_,
		_w23671_
	);
	LUT2 #(
		.INIT('h8)
	) name13160 (
		\wishbone_bd_ram_mem0_reg[238][0]/P0001 ,
		_w13160_,
		_w23672_
	);
	LUT2 #(
		.INIT('h8)
	) name13161 (
		\wishbone_bd_ram_mem0_reg[115][0]/P0001 ,
		_w13112_,
		_w23673_
	);
	LUT2 #(
		.INIT('h8)
	) name13162 (
		\wishbone_bd_ram_mem0_reg[164][0]/P0001 ,
		_w12876_,
		_w23674_
	);
	LUT2 #(
		.INIT('h8)
	) name13163 (
		\wishbone_bd_ram_mem0_reg[14][0]/P0001 ,
		_w13086_,
		_w23675_
	);
	LUT2 #(
		.INIT('h8)
	) name13164 (
		\wishbone_bd_ram_mem0_reg[189][0]/P0001 ,
		_w13042_,
		_w23676_
	);
	LUT2 #(
		.INIT('h8)
	) name13165 (
		\wishbone_bd_ram_mem0_reg[3][0]/P0001 ,
		_w12866_,
		_w23677_
	);
	LUT2 #(
		.INIT('h8)
	) name13166 (
		\wishbone_bd_ram_mem0_reg[194][0]/P0001 ,
		_w12772_,
		_w23678_
	);
	LUT2 #(
		.INIT('h8)
	) name13167 (
		\wishbone_bd_ram_mem0_reg[213][0]/P0001 ,
		_w13002_,
		_w23679_
	);
	LUT2 #(
		.INIT('h8)
	) name13168 (
		\wishbone_bd_ram_mem0_reg[212][0]/P0001 ,
		_w12796_,
		_w23680_
	);
	LUT2 #(
		.INIT('h8)
	) name13169 (
		\wishbone_bd_ram_mem0_reg[84][0]/P0001 ,
		_w12934_,
		_w23681_
	);
	LUT2 #(
		.INIT('h8)
	) name13170 (
		\wishbone_bd_ram_mem0_reg[1][0]/P0001 ,
		_w13014_,
		_w23682_
	);
	LUT2 #(
		.INIT('h8)
	) name13171 (
		\wishbone_bd_ram_mem0_reg[155][0]/P0001 ,
		_w13122_,
		_w23683_
	);
	LUT2 #(
		.INIT('h8)
	) name13172 (
		\wishbone_bd_ram_mem0_reg[62][0]/P0001 ,
		_w12673_,
		_w23684_
	);
	LUT2 #(
		.INIT('h8)
	) name13173 (
		\wishbone_bd_ram_mem0_reg[148][0]/P0001 ,
		_w13000_,
		_w23685_
	);
	LUT2 #(
		.INIT('h8)
	) name13174 (
		\wishbone_bd_ram_mem0_reg[89][0]/P0001 ,
		_w12964_,
		_w23686_
	);
	LUT2 #(
		.INIT('h8)
	) name13175 (
		\wishbone_bd_ram_mem0_reg[41][0]/P0001 ,
		_w13052_,
		_w23687_
	);
	LUT2 #(
		.INIT('h8)
	) name13176 (
		\wishbone_bd_ram_mem0_reg[46][0]/P0001 ,
		_w12884_,
		_w23688_
	);
	LUT2 #(
		.INIT('h8)
	) name13177 (
		\wishbone_bd_ram_mem0_reg[61][0]/P0001 ,
		_w12725_,
		_w23689_
	);
	LUT2 #(
		.INIT('h8)
	) name13178 (
		\wishbone_bd_ram_mem0_reg[230][0]/P0001 ,
		_w13036_,
		_w23690_
	);
	LUT2 #(
		.INIT('h8)
	) name13179 (
		\wishbone_bd_ram_mem0_reg[252][0]/P0001 ,
		_w13080_,
		_w23691_
	);
	LUT2 #(
		.INIT('h8)
	) name13180 (
		\wishbone_bd_ram_mem0_reg[96][0]/P0001 ,
		_w12912_,
		_w23692_
	);
	LUT2 #(
		.INIT('h8)
	) name13181 (
		\wishbone_bd_ram_mem0_reg[123][0]/P0001 ,
		_w13114_,
		_w23693_
	);
	LUT2 #(
		.INIT('h8)
	) name13182 (
		\wishbone_bd_ram_mem0_reg[102][0]/P0001 ,
		_w12685_,
		_w23694_
	);
	LUT2 #(
		.INIT('h8)
	) name13183 (
		\wishbone_bd_ram_mem0_reg[236][0]/P0001 ,
		_w12731_,
		_w23695_
	);
	LUT2 #(
		.INIT('h8)
	) name13184 (
		\wishbone_bd_ram_mem0_reg[113][0]/P0001 ,
		_w13026_,
		_w23696_
	);
	LUT2 #(
		.INIT('h8)
	) name13185 (
		\wishbone_bd_ram_mem0_reg[109][0]/P0001 ,
		_w12888_,
		_w23697_
	);
	LUT2 #(
		.INIT('h8)
	) name13186 (
		\wishbone_bd_ram_mem0_reg[127][0]/P0001 ,
		_w13164_,
		_w23698_
	);
	LUT2 #(
		.INIT('h8)
	) name13187 (
		\wishbone_bd_ram_mem0_reg[205][0]/P0001 ,
		_w13068_,
		_w23699_
	);
	LUT2 #(
		.INIT('h8)
	) name13188 (
		\wishbone_bd_ram_mem0_reg[207][0]/P0001 ,
		_w13180_,
		_w23700_
	);
	LUT2 #(
		.INIT('h8)
	) name13189 (
		\wishbone_bd_ram_mem0_reg[110][0]/P0001 ,
		_w13046_,
		_w23701_
	);
	LUT2 #(
		.INIT('h8)
	) name13190 (
		\wishbone_bd_ram_mem0_reg[149][0]/P0001 ,
		_w12741_,
		_w23702_
	);
	LUT2 #(
		.INIT('h8)
	) name13191 (
		\wishbone_bd_ram_mem0_reg[241][0]/P0001 ,
		_w13006_,
		_w23703_
	);
	LUT2 #(
		.INIT('h8)
	) name13192 (
		\wishbone_bd_ram_mem0_reg[186][0]/P0001 ,
		_w12783_,
		_w23704_
	);
	LUT2 #(
		.INIT('h8)
	) name13193 (
		\wishbone_bd_ram_mem0_reg[119][0]/P0001 ,
		_w13048_,
		_w23705_
	);
	LUT2 #(
		.INIT('h8)
	) name13194 (
		\wishbone_bd_ram_mem0_reg[48][0]/P0001 ,
		_w12970_,
		_w23706_
	);
	LUT2 #(
		.INIT('h8)
	) name13195 (
		\wishbone_bd_ram_mem0_reg[171][0]/P0001 ,
		_w12910_,
		_w23707_
	);
	LUT2 #(
		.INIT('h8)
	) name13196 (
		\wishbone_bd_ram_mem0_reg[22][0]/P0001 ,
		_w13110_,
		_w23708_
	);
	LUT2 #(
		.INIT('h8)
	) name13197 (
		\wishbone_bd_ram_mem0_reg[132][0]/P0001 ,
		_w12992_,
		_w23709_
	);
	LUT2 #(
		.INIT('h8)
	) name13198 (
		\wishbone_bd_ram_mem0_reg[165][0]/P0001 ,
		_w13044_,
		_w23710_
	);
	LUT2 #(
		.INIT('h8)
	) name13199 (
		\wishbone_bd_ram_mem0_reg[141][0]/P0001 ,
		_w13004_,
		_w23711_
	);
	LUT2 #(
		.INIT('h8)
	) name13200 (
		\wishbone_bd_ram_mem0_reg[105][0]/P0001 ,
		_w12751_,
		_w23712_
	);
	LUT2 #(
		.INIT('h8)
	) name13201 (
		\wishbone_bd_ram_mem0_reg[59][0]/P0001 ,
		_w12780_,
		_w23713_
	);
	LUT2 #(
		.INIT('h8)
	) name13202 (
		\wishbone_bd_ram_mem0_reg[51][0]/P0001 ,
		_w13024_,
		_w23714_
	);
	LUT2 #(
		.INIT('h8)
	) name13203 (
		\wishbone_bd_ram_mem0_reg[52][0]/P0001 ,
		_w13082_,
		_w23715_
	);
	LUT2 #(
		.INIT('h8)
	) name13204 (
		\wishbone_bd_ram_mem0_reg[201][0]/P0001 ,
		_w12822_,
		_w23716_
	);
	LUT2 #(
		.INIT('h8)
	) name13205 (
		\wishbone_bd_ram_mem0_reg[4][0]/P0001 ,
		_w12666_,
		_w23717_
	);
	LUT2 #(
		.INIT('h8)
	) name13206 (
		\wishbone_bd_ram_mem0_reg[107][0]/P0001 ,
		_w12749_,
		_w23718_
	);
	LUT2 #(
		.INIT('h8)
	) name13207 (
		\wishbone_bd_ram_mem0_reg[88][0]/P0001 ,
		_w12860_,
		_w23719_
	);
	LUT2 #(
		.INIT('h8)
	) name13208 (
		\wishbone_bd_ram_mem0_reg[204][0]/P0001 ,
		_w13162_,
		_w23720_
	);
	LUT2 #(
		.INIT('h8)
	) name13209 (
		\wishbone_bd_ram_mem0_reg[54][0]/P0001 ,
		_w12770_,
		_w23721_
	);
	LUT2 #(
		.INIT('h8)
	) name13210 (
		\wishbone_bd_ram_mem0_reg[117][0]/P0001 ,
		_w12715_,
		_w23722_
	);
	LUT2 #(
		.INIT('h8)
	) name13211 (
		\wishbone_bd_ram_mem0_reg[34][0]/P0001 ,
		_w12930_,
		_w23723_
	);
	LUT2 #(
		.INIT('h8)
	) name13212 (
		\wishbone_bd_ram_mem0_reg[70][0]/P0001 ,
		_w12840_,
		_w23724_
	);
	LUT2 #(
		.INIT('h8)
	) name13213 (
		\wishbone_bd_ram_mem0_reg[73][0]/P0001 ,
		_w12918_,
		_w23725_
	);
	LUT2 #(
		.INIT('h8)
	) name13214 (
		\wishbone_bd_ram_mem0_reg[157][0]/P0001 ,
		_w12926_,
		_w23726_
	);
	LUT2 #(
		.INIT('h8)
	) name13215 (
		\wishbone_bd_ram_mem0_reg[255][0]/P0001 ,
		_w13072_,
		_w23727_
	);
	LUT2 #(
		.INIT('h8)
	) name13216 (
		\wishbone_bd_ram_mem0_reg[138][0]/P0001 ,
		_w12958_,
		_w23728_
	);
	LUT2 #(
		.INIT('h8)
	) name13217 (
		\wishbone_bd_ram_mem0_reg[104][0]/P0001 ,
		_w13148_,
		_w23729_
	);
	LUT2 #(
		.INIT('h8)
	) name13218 (
		\wishbone_bd_ram_mem0_reg[167][0]/P0001 ,
		_w12986_,
		_w23730_
	);
	LUT2 #(
		.INIT('h8)
	) name13219 (
		\wishbone_bd_ram_mem0_reg[20][0]/P0001 ,
		_w13174_,
		_w23731_
	);
	LUT2 #(
		.INIT('h8)
	) name13220 (
		\wishbone_bd_ram_mem0_reg[178][0]/P0001 ,
		_w12886_,
		_w23732_
	);
	LUT2 #(
		.INIT('h8)
	) name13221 (
		\wishbone_bd_ram_mem0_reg[139][0]/P0001 ,
		_w12814_,
		_w23733_
	);
	LUT2 #(
		.INIT('h8)
	) name13222 (
		\wishbone_bd_ram_mem0_reg[206][0]/P0001 ,
		_w12954_,
		_w23734_
	);
	LUT2 #(
		.INIT('h8)
	) name13223 (
		\wishbone_bd_ram_mem0_reg[129][0]/P0001 ,
		_w12776_,
		_w23735_
	);
	LUT2 #(
		.INIT('h8)
	) name13224 (
		\wishbone_bd_ram_mem0_reg[56][0]/P0001 ,
		_w12778_,
		_w23736_
	);
	LUT2 #(
		.INIT('h8)
	) name13225 (
		\wishbone_bd_ram_mem0_reg[19][0]/P0001 ,
		_w13012_,
		_w23737_
	);
	LUT2 #(
		.INIT('h8)
	) name13226 (
		\wishbone_bd_ram_mem0_reg[108][0]/P0001 ,
		_w13156_,
		_w23738_
	);
	LUT2 #(
		.INIT('h8)
	) name13227 (
		\wishbone_bd_ram_mem0_reg[218][0]/P0001 ,
		_w13206_,
		_w23739_
	);
	LUT2 #(
		.INIT('h8)
	) name13228 (
		\wishbone_bd_ram_mem0_reg[239][0]/P0001 ,
		_w12862_,
		_w23740_
	);
	LUT2 #(
		.INIT('h8)
	) name13229 (
		\wishbone_bd_ram_mem0_reg[92][0]/P0001 ,
		_w13010_,
		_w23741_
	);
	LUT2 #(
		.INIT('h8)
	) name13230 (
		\wishbone_bd_ram_mem0_reg[173][0]/P0001 ,
		_w12854_,
		_w23742_
	);
	LUT2 #(
		.INIT('h8)
	) name13231 (
		\wishbone_bd_ram_mem0_reg[221][0]/P0001 ,
		_w12802_,
		_w23743_
	);
	LUT2 #(
		.INIT('h8)
	) name13232 (
		\wishbone_bd_ram_mem0_reg[220][0]/P0001 ,
		_w13066_,
		_w23744_
	);
	LUT2 #(
		.INIT('h8)
	) name13233 (
		\wishbone_bd_ram_mem0_reg[136][0]/P0001 ,
		_w13064_,
		_w23745_
	);
	LUT2 #(
		.INIT('h8)
	) name13234 (
		\wishbone_bd_ram_mem0_reg[145][0]/P0001 ,
		_w13106_,
		_w23746_
	);
	LUT2 #(
		.INIT('h8)
	) name13235 (
		\wishbone_bd_ram_mem0_reg[143][0]/P0001 ,
		_w12922_,
		_w23747_
	);
	LUT2 #(
		.INIT('h8)
	) name13236 (
		\wishbone_bd_ram_mem0_reg[254][0]/P0001 ,
		_w12892_,
		_w23748_
	);
	LUT2 #(
		.INIT('h8)
	) name13237 (
		\wishbone_bd_ram_mem0_reg[27][0]/P0001 ,
		_w12880_,
		_w23749_
	);
	LUT2 #(
		.INIT('h8)
	) name13238 (
		\wishbone_bd_ram_mem0_reg[29][0]/P0001 ,
		_w12952_,
		_w23750_
	);
	LUT2 #(
		.INIT('h8)
	) name13239 (
		\wishbone_bd_ram_mem0_reg[154][0]/P0001 ,
		_w12962_,
		_w23751_
	);
	LUT2 #(
		.INIT('h8)
	) name13240 (
		\wishbone_bd_ram_mem0_reg[83][0]/P0001 ,
		_w12916_,
		_w23752_
	);
	LUT2 #(
		.INIT('h8)
	) name13241 (
		\wishbone_bd_ram_mem0_reg[13][0]/P0001 ,
		_w13178_,
		_w23753_
	);
	LUT2 #(
		.INIT('h8)
	) name13242 (
		\wishbone_bd_ram_mem0_reg[80][0]/P0001 ,
		_w12689_,
		_w23754_
	);
	LUT2 #(
		.INIT('h8)
	) name13243 (
		\wishbone_bd_ram_mem0_reg[172][0]/P0001 ,
		_w12944_,
		_w23755_
	);
	LUT2 #(
		.INIT('h8)
	) name13244 (
		\wishbone_bd_ram_mem0_reg[100][0]/P0001 ,
		_w12960_,
		_w23756_
	);
	LUT2 #(
		.INIT('h8)
	) name13245 (
		\wishbone_bd_ram_mem0_reg[71][0]/P0001 ,
		_w12798_,
		_w23757_
	);
	LUT2 #(
		.INIT('h8)
	) name13246 (
		\wishbone_bd_ram_mem0_reg[35][0]/P0001 ,
		_w12703_,
		_w23758_
	);
	LUT2 #(
		.INIT('h8)
	) name13247 (
		\wishbone_bd_ram_mem0_reg[224][0]/P0001 ,
		_w12902_,
		_w23759_
	);
	LUT2 #(
		.INIT('h8)
	) name13248 (
		\wishbone_bd_ram_mem0_reg[53][0]/P0001 ,
		_w13020_,
		_w23760_
	);
	LUT2 #(
		.INIT('h8)
	) name13249 (
		\wishbone_bd_ram_mem0_reg[253][0]/P0001 ,
		_w13100_,
		_w23761_
	);
	LUT2 #(
		.INIT('h8)
	) name13250 (
		\wishbone_bd_ram_mem0_reg[170][0]/P0001 ,
		_w13030_,
		_w23762_
	);
	LUT2 #(
		.INIT('h8)
	) name13251 (
		\wishbone_bd_ram_mem0_reg[95][0]/P0001 ,
		_w12844_,
		_w23763_
	);
	LUT2 #(
		.INIT('h8)
	) name13252 (
		\wishbone_bd_ram_mem0_reg[156][0]/P0001 ,
		_w13190_,
		_w23764_
	);
	LUT2 #(
		.INIT('h8)
	) name13253 (
		\wishbone_bd_ram_mem0_reg[72][0]/P0001 ,
		_w12810_,
		_w23765_
	);
	LUT2 #(
		.INIT('h8)
	) name13254 (
		\wishbone_bd_ram_mem0_reg[142][0]/P0001 ,
		_w12928_,
		_w23766_
	);
	LUT2 #(
		.INIT('h8)
	) name13255 (
		\wishbone_bd_ram_mem0_reg[97][0]/P0001 ,
		_w13096_,
		_w23767_
	);
	LUT2 #(
		.INIT('h8)
	) name13256 (
		\wishbone_bd_ram_mem0_reg[65][0]/P0001 ,
		_w13176_,
		_w23768_
	);
	LUT2 #(
		.INIT('h8)
	) name13257 (
		\wishbone_bd_ram_mem0_reg[245][0]/P0001 ,
		_w13022_,
		_w23769_
	);
	LUT2 #(
		.INIT('h8)
	) name13258 (
		\wishbone_bd_ram_mem0_reg[2][0]/P0001 ,
		_w13088_,
		_w23770_
	);
	LUT2 #(
		.INIT('h8)
	) name13259 (
		\wishbone_bd_ram_mem0_reg[182][0]/P0001 ,
		_w12820_,
		_w23771_
	);
	LUT2 #(
		.INIT('h8)
	) name13260 (
		\wishbone_bd_ram_mem0_reg[99][0]/P0001 ,
		_w13038_,
		_w23772_
	);
	LUT2 #(
		.INIT('h8)
	) name13261 (
		\wishbone_bd_ram_mem0_reg[67][0]/P0001 ,
		_w13134_,
		_w23773_
	);
	LUT2 #(
		.INIT('h8)
	) name13262 (
		\wishbone_bd_ram_mem0_reg[116][0]/P0001 ,
		_w12998_,
		_w23774_
	);
	LUT2 #(
		.INIT('h8)
	) name13263 (
		\wishbone_bd_ram_mem0_reg[75][0]/P0001 ,
		_w12826_,
		_w23775_
	);
	LUT2 #(
		.INIT('h8)
	) name13264 (
		\wishbone_bd_ram_mem0_reg[168][0]/P0001 ,
		_w13208_,
		_w23776_
	);
	LUT2 #(
		.INIT('h8)
	) name13265 (
		\wishbone_bd_ram_mem0_reg[240][0]/P0001 ,
		_w12864_,
		_w23777_
	);
	LUT2 #(
		.INIT('h8)
	) name13266 (
		\wishbone_bd_ram_mem0_reg[152][0]/P0001 ,
		_w12966_,
		_w23778_
	);
	LUT2 #(
		.INIT('h8)
	) name13267 (
		\wishbone_bd_ram_mem0_reg[227][0]/P0001 ,
		_w12936_,
		_w23779_
	);
	LUT2 #(
		.INIT('h8)
	) name13268 (
		\wishbone_bd_ram_mem0_reg[106][0]/P0001 ,
		_w12713_,
		_w23780_
	);
	LUT2 #(
		.INIT('h8)
	) name13269 (
		\wishbone_bd_ram_mem0_reg[161][0]/P0001 ,
		_w12754_,
		_w23781_
	);
	LUT2 #(
		.INIT('h8)
	) name13270 (
		\wishbone_bd_ram_mem0_reg[85][0]/P0001 ,
		_w13216_,
		_w23782_
	);
	LUT2 #(
		.INIT('h8)
	) name13271 (
		\wishbone_bd_ram_mem0_reg[202][0]/P0001 ,
		_w12870_,
		_w23783_
	);
	LUT2 #(
		.INIT('h8)
	) name13272 (
		\wishbone_bd_ram_mem0_reg[23][0]/P0001 ,
		_w13008_,
		_w23784_
	);
	LUT2 #(
		.INIT('h8)
	) name13273 (
		\wishbone_bd_ram_mem0_reg[208][0]/P0001 ,
		_w13032_,
		_w23785_
	);
	LUT2 #(
		.INIT('h8)
	) name13274 (
		\wishbone_bd_ram_mem0_reg[76][0]/P0001 ,
		_w13184_,
		_w23786_
	);
	LUT2 #(
		.INIT('h8)
	) name13275 (
		\wishbone_bd_ram_mem0_reg[90][0]/P0001 ,
		_w12978_,
		_w23787_
	);
	LUT2 #(
		.INIT('h8)
	) name13276 (
		\wishbone_bd_ram_mem0_reg[128][0]/P0001 ,
		_w12793_,
		_w23788_
	);
	LUT2 #(
		.INIT('h8)
	) name13277 (
		\wishbone_bd_ram_mem0_reg[187][0]/P0001 ,
		_w13196_,
		_w23789_
	);
	LUT2 #(
		.INIT('h8)
	) name13278 (
		\wishbone_bd_ram_mem0_reg[248][0]/P0001 ,
		_w12789_,
		_w23790_
	);
	LUT2 #(
		.INIT('h8)
	) name13279 (
		\wishbone_bd_ram_mem0_reg[243][0]/P0001 ,
		_w12804_,
		_w23791_
	);
	LUT2 #(
		.INIT('h8)
	) name13280 (
		\wishbone_bd_ram_mem0_reg[191][0]/P0001 ,
		_w13034_,
		_w23792_
	);
	LUT2 #(
		.INIT('h8)
	) name13281 (
		\wishbone_bd_ram_mem0_reg[217][0]/P0001 ,
		_w13188_,
		_w23793_
	);
	LUT2 #(
		.INIT('h8)
	) name13282 (
		\wishbone_bd_ram_mem0_reg[229][0]/P0001 ,
		_w12711_,
		_w23794_
	);
	LUT2 #(
		.INIT('h8)
	) name13283 (
		\wishbone_bd_ram_mem0_reg[57][0]/P0001 ,
		_w13116_,
		_w23795_
	);
	LUT2 #(
		.INIT('h8)
	) name13284 (
		\wishbone_bd_ram_mem0_reg[177][0]/P0001 ,
		_w12996_,
		_w23796_
	);
	LUT2 #(
		.INIT('h8)
	) name13285 (
		\wishbone_bd_ram_mem0_reg[163][0]/P0001 ,
		_w12882_,
		_w23797_
	);
	LUT2 #(
		.INIT('h8)
	) name13286 (
		\wishbone_bd_ram_mem0_reg[190][0]/P0001 ,
		_w12858_,
		_w23798_
	);
	LUT2 #(
		.INIT('h8)
	) name13287 (
		\wishbone_bd_ram_mem0_reg[120][0]/P0001 ,
		_w12707_,
		_w23799_
	);
	LUT2 #(
		.INIT('h8)
	) name13288 (
		\wishbone_bd_ram_mem0_reg[17][0]/P0001 ,
		_w12848_,
		_w23800_
	);
	LUT2 #(
		.INIT('h8)
	) name13289 (
		\wishbone_bd_ram_mem0_reg[225][0]/P0001 ,
		_w13092_,
		_w23801_
	);
	LUT2 #(
		.INIT('h8)
	) name13290 (
		\wishbone_bd_ram_mem0_reg[219][0]/P0001 ,
		_w12806_,
		_w23802_
	);
	LUT2 #(
		.INIT('h8)
	) name13291 (
		\wishbone_bd_ram_mem0_reg[231][0]/P0001 ,
		_w12856_,
		_w23803_
	);
	LUT2 #(
		.INIT('h8)
	) name13292 (
		\wishbone_bd_ram_mem0_reg[77][0]/P0001 ,
		_w12982_,
		_w23804_
	);
	LUT2 #(
		.INIT('h8)
	) name13293 (
		\wishbone_bd_ram_mem0_reg[37][0]/P0001 ,
		_w13102_,
		_w23805_
	);
	LUT2 #(
		.INIT('h8)
	) name13294 (
		\wishbone_bd_ram_mem0_reg[181][0]/P0001 ,
		_w12828_,
		_w23806_
	);
	LUT2 #(
		.INIT('h8)
	) name13295 (
		\wishbone_bd_ram_mem0_reg[44][0]/P0001 ,
		_w12896_,
		_w23807_
	);
	LUT2 #(
		.INIT('h8)
	) name13296 (
		\wishbone_bd_ram_mem0_reg[118][0]/P0001 ,
		_w12830_,
		_w23808_
	);
	LUT2 #(
		.INIT('h8)
	) name13297 (
		\wishbone_bd_ram_mem0_reg[137][0]/P0001 ,
		_w13168_,
		_w23809_
	);
	LUT2 #(
		.INIT('h8)
	) name13298 (
		\wishbone_bd_ram_mem0_reg[43][0]/P0001 ,
		_w13200_,
		_w23810_
	);
	LUT2 #(
		.INIT('h8)
	) name13299 (
		\wishbone_bd_ram_mem0_reg[200][0]/P0001 ,
		_w12988_,
		_w23811_
	);
	LUT2 #(
		.INIT('h8)
	) name13300 (
		\wishbone_bd_ram_mem0_reg[125][0]/P0001 ,
		_w12956_,
		_w23812_
	);
	LUT2 #(
		.INIT('h8)
	) name13301 (
		\wishbone_bd_ram_mem0_reg[124][0]/P0001 ,
		_w13058_,
		_w23813_
	);
	LUT2 #(
		.INIT('h8)
	) name13302 (
		\wishbone_bd_ram_mem0_reg[15][0]/P0001 ,
		_w13210_,
		_w23814_
	);
	LUT2 #(
		.INIT('h8)
	) name13303 (
		\wishbone_bd_ram_mem0_reg[63][0]/P0001 ,
		_w12850_,
		_w23815_
	);
	LUT2 #(
		.INIT('h8)
	) name13304 (
		\wishbone_bd_ram_mem0_reg[69][0]/P0001 ,
		_w12738_,
		_w23816_
	);
	LUT2 #(
		.INIT('h8)
	) name13305 (
		\wishbone_bd_ram_mem0_reg[40][0]/P0001 ,
		_w13132_,
		_w23817_
	);
	LUT2 #(
		.INIT('h8)
	) name13306 (
		\wishbone_bd_ram_mem0_reg[16][0]/P0001 ,
		_w13140_,
		_w23818_
	);
	LUT2 #(
		.INIT('h8)
	) name13307 (
		\wishbone_bd_ram_mem0_reg[55][0]/P0001 ,
		_w12785_,
		_w23819_
	);
	LUT2 #(
		.INIT('h8)
	) name13308 (
		\wishbone_bd_ram_mem0_reg[131][0]/P0001 ,
		_w12852_,
		_w23820_
	);
	LUT2 #(
		.INIT('h8)
	) name13309 (
		\wishbone_bd_ram_mem0_reg[233][0]/P0001 ,
		_w12836_,
		_w23821_
	);
	LUT2 #(
		.INIT('h8)
	) name13310 (
		\wishbone_bd_ram_mem0_reg[158][0]/P0001 ,
		_w12898_,
		_w23822_
	);
	LUT2 #(
		.INIT('h8)
	) name13311 (
		\wishbone_bd_ram_mem0_reg[147][0]/P0001 ,
		_w13146_,
		_w23823_
	);
	LUT2 #(
		.INIT('h8)
	) name13312 (
		\wishbone_bd_ram_mem0_reg[49][0]/P0001 ,
		_w12994_,
		_w23824_
	);
	LUT2 #(
		.INIT('h8)
	) name13313 (
		\wishbone_bd_ram_mem0_reg[94][0]/P0001 ,
		_w13186_,
		_w23825_
	);
	LUT2 #(
		.INIT('h8)
	) name13314 (
		\wishbone_bd_ram_mem0_reg[74][0]/P0001 ,
		_w12812_,
		_w23826_
	);
	LUT2 #(
		.INIT('h8)
	) name13315 (
		\wishbone_bd_ram_mem0_reg[246][0]/P0001 ,
		_w13076_,
		_w23827_
	);
	LUT2 #(
		.INIT('h8)
	) name13316 (
		\wishbone_bd_ram_mem0_reg[193][0]/P0001 ,
		_w13056_,
		_w23828_
	);
	LUT2 #(
		.INIT('h8)
	) name13317 (
		\wishbone_bd_ram_mem0_reg[50][0]/P0001 ,
		_w13150_,
		_w23829_
	);
	LUT2 #(
		.INIT('h8)
	) name13318 (
		\wishbone_bd_ram_mem0_reg[38][0]/P0001 ,
		_w13182_,
		_w23830_
	);
	LUT2 #(
		.INIT('h8)
	) name13319 (
		\wishbone_bd_ram_mem0_reg[121][0]/P0001 ,
		_w13078_,
		_w23831_
	);
	LUT2 #(
		.INIT('h8)
	) name13320 (
		\wishbone_bd_ram_mem0_reg[162][0]/P0001 ,
		_w13098_,
		_w23832_
	);
	LUT2 #(
		.INIT('h8)
	) name13321 (
		\wishbone_bd_ram_mem0_reg[210][0]/P0001 ,
		_w12924_,
		_w23833_
	);
	LUT2 #(
		.INIT('h8)
	) name13322 (
		\wishbone_bd_ram_mem0_reg[176][0]/P0001 ,
		_w12868_,
		_w23834_
	);
	LUT2 #(
		.INIT('h8)
	) name13323 (
		\wishbone_bd_ram_mem0_reg[33][0]/P0001 ,
		_w12980_,
		_w23835_
	);
	LUT2 #(
		.INIT('h8)
	) name13324 (
		\wishbone_bd_ram_mem0_reg[134][0]/P0001 ,
		_w12763_,
		_w23836_
	);
	LUT2 #(
		.INIT('h8)
	) name13325 (
		\wishbone_bd_ram_mem0_reg[180][0]/P0001 ,
		_w12791_,
		_w23837_
	);
	LUT2 #(
		.INIT('h8)
	) name13326 (
		\wishbone_bd_ram_mem0_reg[98][0]/P0001 ,
		_w12816_,
		_w23838_
	);
	LUT2 #(
		.INIT('h1)
	) name13327 (
		_w23583_,
		_w23584_,
		_w23839_
	);
	LUT2 #(
		.INIT('h1)
	) name13328 (
		_w23585_,
		_w23586_,
		_w23840_
	);
	LUT2 #(
		.INIT('h1)
	) name13329 (
		_w23587_,
		_w23588_,
		_w23841_
	);
	LUT2 #(
		.INIT('h1)
	) name13330 (
		_w23589_,
		_w23590_,
		_w23842_
	);
	LUT2 #(
		.INIT('h1)
	) name13331 (
		_w23591_,
		_w23592_,
		_w23843_
	);
	LUT2 #(
		.INIT('h1)
	) name13332 (
		_w23593_,
		_w23594_,
		_w23844_
	);
	LUT2 #(
		.INIT('h1)
	) name13333 (
		_w23595_,
		_w23596_,
		_w23845_
	);
	LUT2 #(
		.INIT('h1)
	) name13334 (
		_w23597_,
		_w23598_,
		_w23846_
	);
	LUT2 #(
		.INIT('h1)
	) name13335 (
		_w23599_,
		_w23600_,
		_w23847_
	);
	LUT2 #(
		.INIT('h1)
	) name13336 (
		_w23601_,
		_w23602_,
		_w23848_
	);
	LUT2 #(
		.INIT('h1)
	) name13337 (
		_w23603_,
		_w23604_,
		_w23849_
	);
	LUT2 #(
		.INIT('h1)
	) name13338 (
		_w23605_,
		_w23606_,
		_w23850_
	);
	LUT2 #(
		.INIT('h1)
	) name13339 (
		_w23607_,
		_w23608_,
		_w23851_
	);
	LUT2 #(
		.INIT('h1)
	) name13340 (
		_w23609_,
		_w23610_,
		_w23852_
	);
	LUT2 #(
		.INIT('h1)
	) name13341 (
		_w23611_,
		_w23612_,
		_w23853_
	);
	LUT2 #(
		.INIT('h1)
	) name13342 (
		_w23613_,
		_w23614_,
		_w23854_
	);
	LUT2 #(
		.INIT('h1)
	) name13343 (
		_w23615_,
		_w23616_,
		_w23855_
	);
	LUT2 #(
		.INIT('h1)
	) name13344 (
		_w23617_,
		_w23618_,
		_w23856_
	);
	LUT2 #(
		.INIT('h1)
	) name13345 (
		_w23619_,
		_w23620_,
		_w23857_
	);
	LUT2 #(
		.INIT('h1)
	) name13346 (
		_w23621_,
		_w23622_,
		_w23858_
	);
	LUT2 #(
		.INIT('h1)
	) name13347 (
		_w23623_,
		_w23624_,
		_w23859_
	);
	LUT2 #(
		.INIT('h1)
	) name13348 (
		_w23625_,
		_w23626_,
		_w23860_
	);
	LUT2 #(
		.INIT('h1)
	) name13349 (
		_w23627_,
		_w23628_,
		_w23861_
	);
	LUT2 #(
		.INIT('h1)
	) name13350 (
		_w23629_,
		_w23630_,
		_w23862_
	);
	LUT2 #(
		.INIT('h1)
	) name13351 (
		_w23631_,
		_w23632_,
		_w23863_
	);
	LUT2 #(
		.INIT('h1)
	) name13352 (
		_w23633_,
		_w23634_,
		_w23864_
	);
	LUT2 #(
		.INIT('h1)
	) name13353 (
		_w23635_,
		_w23636_,
		_w23865_
	);
	LUT2 #(
		.INIT('h1)
	) name13354 (
		_w23637_,
		_w23638_,
		_w23866_
	);
	LUT2 #(
		.INIT('h1)
	) name13355 (
		_w23639_,
		_w23640_,
		_w23867_
	);
	LUT2 #(
		.INIT('h1)
	) name13356 (
		_w23641_,
		_w23642_,
		_w23868_
	);
	LUT2 #(
		.INIT('h1)
	) name13357 (
		_w23643_,
		_w23644_,
		_w23869_
	);
	LUT2 #(
		.INIT('h1)
	) name13358 (
		_w23645_,
		_w23646_,
		_w23870_
	);
	LUT2 #(
		.INIT('h1)
	) name13359 (
		_w23647_,
		_w23648_,
		_w23871_
	);
	LUT2 #(
		.INIT('h1)
	) name13360 (
		_w23649_,
		_w23650_,
		_w23872_
	);
	LUT2 #(
		.INIT('h1)
	) name13361 (
		_w23651_,
		_w23652_,
		_w23873_
	);
	LUT2 #(
		.INIT('h1)
	) name13362 (
		_w23653_,
		_w23654_,
		_w23874_
	);
	LUT2 #(
		.INIT('h1)
	) name13363 (
		_w23655_,
		_w23656_,
		_w23875_
	);
	LUT2 #(
		.INIT('h1)
	) name13364 (
		_w23657_,
		_w23658_,
		_w23876_
	);
	LUT2 #(
		.INIT('h1)
	) name13365 (
		_w23659_,
		_w23660_,
		_w23877_
	);
	LUT2 #(
		.INIT('h1)
	) name13366 (
		_w23661_,
		_w23662_,
		_w23878_
	);
	LUT2 #(
		.INIT('h1)
	) name13367 (
		_w23663_,
		_w23664_,
		_w23879_
	);
	LUT2 #(
		.INIT('h1)
	) name13368 (
		_w23665_,
		_w23666_,
		_w23880_
	);
	LUT2 #(
		.INIT('h1)
	) name13369 (
		_w23667_,
		_w23668_,
		_w23881_
	);
	LUT2 #(
		.INIT('h1)
	) name13370 (
		_w23669_,
		_w23670_,
		_w23882_
	);
	LUT2 #(
		.INIT('h1)
	) name13371 (
		_w23671_,
		_w23672_,
		_w23883_
	);
	LUT2 #(
		.INIT('h1)
	) name13372 (
		_w23673_,
		_w23674_,
		_w23884_
	);
	LUT2 #(
		.INIT('h1)
	) name13373 (
		_w23675_,
		_w23676_,
		_w23885_
	);
	LUT2 #(
		.INIT('h1)
	) name13374 (
		_w23677_,
		_w23678_,
		_w23886_
	);
	LUT2 #(
		.INIT('h1)
	) name13375 (
		_w23679_,
		_w23680_,
		_w23887_
	);
	LUT2 #(
		.INIT('h1)
	) name13376 (
		_w23681_,
		_w23682_,
		_w23888_
	);
	LUT2 #(
		.INIT('h1)
	) name13377 (
		_w23683_,
		_w23684_,
		_w23889_
	);
	LUT2 #(
		.INIT('h1)
	) name13378 (
		_w23685_,
		_w23686_,
		_w23890_
	);
	LUT2 #(
		.INIT('h1)
	) name13379 (
		_w23687_,
		_w23688_,
		_w23891_
	);
	LUT2 #(
		.INIT('h1)
	) name13380 (
		_w23689_,
		_w23690_,
		_w23892_
	);
	LUT2 #(
		.INIT('h1)
	) name13381 (
		_w23691_,
		_w23692_,
		_w23893_
	);
	LUT2 #(
		.INIT('h1)
	) name13382 (
		_w23693_,
		_w23694_,
		_w23894_
	);
	LUT2 #(
		.INIT('h1)
	) name13383 (
		_w23695_,
		_w23696_,
		_w23895_
	);
	LUT2 #(
		.INIT('h1)
	) name13384 (
		_w23697_,
		_w23698_,
		_w23896_
	);
	LUT2 #(
		.INIT('h1)
	) name13385 (
		_w23699_,
		_w23700_,
		_w23897_
	);
	LUT2 #(
		.INIT('h1)
	) name13386 (
		_w23701_,
		_w23702_,
		_w23898_
	);
	LUT2 #(
		.INIT('h1)
	) name13387 (
		_w23703_,
		_w23704_,
		_w23899_
	);
	LUT2 #(
		.INIT('h1)
	) name13388 (
		_w23705_,
		_w23706_,
		_w23900_
	);
	LUT2 #(
		.INIT('h1)
	) name13389 (
		_w23707_,
		_w23708_,
		_w23901_
	);
	LUT2 #(
		.INIT('h1)
	) name13390 (
		_w23709_,
		_w23710_,
		_w23902_
	);
	LUT2 #(
		.INIT('h1)
	) name13391 (
		_w23711_,
		_w23712_,
		_w23903_
	);
	LUT2 #(
		.INIT('h1)
	) name13392 (
		_w23713_,
		_w23714_,
		_w23904_
	);
	LUT2 #(
		.INIT('h1)
	) name13393 (
		_w23715_,
		_w23716_,
		_w23905_
	);
	LUT2 #(
		.INIT('h1)
	) name13394 (
		_w23717_,
		_w23718_,
		_w23906_
	);
	LUT2 #(
		.INIT('h1)
	) name13395 (
		_w23719_,
		_w23720_,
		_w23907_
	);
	LUT2 #(
		.INIT('h1)
	) name13396 (
		_w23721_,
		_w23722_,
		_w23908_
	);
	LUT2 #(
		.INIT('h1)
	) name13397 (
		_w23723_,
		_w23724_,
		_w23909_
	);
	LUT2 #(
		.INIT('h1)
	) name13398 (
		_w23725_,
		_w23726_,
		_w23910_
	);
	LUT2 #(
		.INIT('h1)
	) name13399 (
		_w23727_,
		_w23728_,
		_w23911_
	);
	LUT2 #(
		.INIT('h1)
	) name13400 (
		_w23729_,
		_w23730_,
		_w23912_
	);
	LUT2 #(
		.INIT('h1)
	) name13401 (
		_w23731_,
		_w23732_,
		_w23913_
	);
	LUT2 #(
		.INIT('h1)
	) name13402 (
		_w23733_,
		_w23734_,
		_w23914_
	);
	LUT2 #(
		.INIT('h1)
	) name13403 (
		_w23735_,
		_w23736_,
		_w23915_
	);
	LUT2 #(
		.INIT('h1)
	) name13404 (
		_w23737_,
		_w23738_,
		_w23916_
	);
	LUT2 #(
		.INIT('h1)
	) name13405 (
		_w23739_,
		_w23740_,
		_w23917_
	);
	LUT2 #(
		.INIT('h1)
	) name13406 (
		_w23741_,
		_w23742_,
		_w23918_
	);
	LUT2 #(
		.INIT('h1)
	) name13407 (
		_w23743_,
		_w23744_,
		_w23919_
	);
	LUT2 #(
		.INIT('h1)
	) name13408 (
		_w23745_,
		_w23746_,
		_w23920_
	);
	LUT2 #(
		.INIT('h1)
	) name13409 (
		_w23747_,
		_w23748_,
		_w23921_
	);
	LUT2 #(
		.INIT('h1)
	) name13410 (
		_w23749_,
		_w23750_,
		_w23922_
	);
	LUT2 #(
		.INIT('h1)
	) name13411 (
		_w23751_,
		_w23752_,
		_w23923_
	);
	LUT2 #(
		.INIT('h1)
	) name13412 (
		_w23753_,
		_w23754_,
		_w23924_
	);
	LUT2 #(
		.INIT('h1)
	) name13413 (
		_w23755_,
		_w23756_,
		_w23925_
	);
	LUT2 #(
		.INIT('h1)
	) name13414 (
		_w23757_,
		_w23758_,
		_w23926_
	);
	LUT2 #(
		.INIT('h1)
	) name13415 (
		_w23759_,
		_w23760_,
		_w23927_
	);
	LUT2 #(
		.INIT('h1)
	) name13416 (
		_w23761_,
		_w23762_,
		_w23928_
	);
	LUT2 #(
		.INIT('h1)
	) name13417 (
		_w23763_,
		_w23764_,
		_w23929_
	);
	LUT2 #(
		.INIT('h1)
	) name13418 (
		_w23765_,
		_w23766_,
		_w23930_
	);
	LUT2 #(
		.INIT('h1)
	) name13419 (
		_w23767_,
		_w23768_,
		_w23931_
	);
	LUT2 #(
		.INIT('h1)
	) name13420 (
		_w23769_,
		_w23770_,
		_w23932_
	);
	LUT2 #(
		.INIT('h1)
	) name13421 (
		_w23771_,
		_w23772_,
		_w23933_
	);
	LUT2 #(
		.INIT('h1)
	) name13422 (
		_w23773_,
		_w23774_,
		_w23934_
	);
	LUT2 #(
		.INIT('h1)
	) name13423 (
		_w23775_,
		_w23776_,
		_w23935_
	);
	LUT2 #(
		.INIT('h1)
	) name13424 (
		_w23777_,
		_w23778_,
		_w23936_
	);
	LUT2 #(
		.INIT('h1)
	) name13425 (
		_w23779_,
		_w23780_,
		_w23937_
	);
	LUT2 #(
		.INIT('h1)
	) name13426 (
		_w23781_,
		_w23782_,
		_w23938_
	);
	LUT2 #(
		.INIT('h1)
	) name13427 (
		_w23783_,
		_w23784_,
		_w23939_
	);
	LUT2 #(
		.INIT('h1)
	) name13428 (
		_w23785_,
		_w23786_,
		_w23940_
	);
	LUT2 #(
		.INIT('h1)
	) name13429 (
		_w23787_,
		_w23788_,
		_w23941_
	);
	LUT2 #(
		.INIT('h1)
	) name13430 (
		_w23789_,
		_w23790_,
		_w23942_
	);
	LUT2 #(
		.INIT('h1)
	) name13431 (
		_w23791_,
		_w23792_,
		_w23943_
	);
	LUT2 #(
		.INIT('h1)
	) name13432 (
		_w23793_,
		_w23794_,
		_w23944_
	);
	LUT2 #(
		.INIT('h1)
	) name13433 (
		_w23795_,
		_w23796_,
		_w23945_
	);
	LUT2 #(
		.INIT('h1)
	) name13434 (
		_w23797_,
		_w23798_,
		_w23946_
	);
	LUT2 #(
		.INIT('h1)
	) name13435 (
		_w23799_,
		_w23800_,
		_w23947_
	);
	LUT2 #(
		.INIT('h1)
	) name13436 (
		_w23801_,
		_w23802_,
		_w23948_
	);
	LUT2 #(
		.INIT('h1)
	) name13437 (
		_w23803_,
		_w23804_,
		_w23949_
	);
	LUT2 #(
		.INIT('h1)
	) name13438 (
		_w23805_,
		_w23806_,
		_w23950_
	);
	LUT2 #(
		.INIT('h1)
	) name13439 (
		_w23807_,
		_w23808_,
		_w23951_
	);
	LUT2 #(
		.INIT('h1)
	) name13440 (
		_w23809_,
		_w23810_,
		_w23952_
	);
	LUT2 #(
		.INIT('h1)
	) name13441 (
		_w23811_,
		_w23812_,
		_w23953_
	);
	LUT2 #(
		.INIT('h1)
	) name13442 (
		_w23813_,
		_w23814_,
		_w23954_
	);
	LUT2 #(
		.INIT('h1)
	) name13443 (
		_w23815_,
		_w23816_,
		_w23955_
	);
	LUT2 #(
		.INIT('h1)
	) name13444 (
		_w23817_,
		_w23818_,
		_w23956_
	);
	LUT2 #(
		.INIT('h1)
	) name13445 (
		_w23819_,
		_w23820_,
		_w23957_
	);
	LUT2 #(
		.INIT('h1)
	) name13446 (
		_w23821_,
		_w23822_,
		_w23958_
	);
	LUT2 #(
		.INIT('h1)
	) name13447 (
		_w23823_,
		_w23824_,
		_w23959_
	);
	LUT2 #(
		.INIT('h1)
	) name13448 (
		_w23825_,
		_w23826_,
		_w23960_
	);
	LUT2 #(
		.INIT('h1)
	) name13449 (
		_w23827_,
		_w23828_,
		_w23961_
	);
	LUT2 #(
		.INIT('h1)
	) name13450 (
		_w23829_,
		_w23830_,
		_w23962_
	);
	LUT2 #(
		.INIT('h1)
	) name13451 (
		_w23831_,
		_w23832_,
		_w23963_
	);
	LUT2 #(
		.INIT('h1)
	) name13452 (
		_w23833_,
		_w23834_,
		_w23964_
	);
	LUT2 #(
		.INIT('h1)
	) name13453 (
		_w23835_,
		_w23836_,
		_w23965_
	);
	LUT2 #(
		.INIT('h1)
	) name13454 (
		_w23837_,
		_w23838_,
		_w23966_
	);
	LUT2 #(
		.INIT('h8)
	) name13455 (
		_w23965_,
		_w23966_,
		_w23967_
	);
	LUT2 #(
		.INIT('h8)
	) name13456 (
		_w23963_,
		_w23964_,
		_w23968_
	);
	LUT2 #(
		.INIT('h8)
	) name13457 (
		_w23961_,
		_w23962_,
		_w23969_
	);
	LUT2 #(
		.INIT('h8)
	) name13458 (
		_w23959_,
		_w23960_,
		_w23970_
	);
	LUT2 #(
		.INIT('h8)
	) name13459 (
		_w23957_,
		_w23958_,
		_w23971_
	);
	LUT2 #(
		.INIT('h8)
	) name13460 (
		_w23955_,
		_w23956_,
		_w23972_
	);
	LUT2 #(
		.INIT('h8)
	) name13461 (
		_w23953_,
		_w23954_,
		_w23973_
	);
	LUT2 #(
		.INIT('h8)
	) name13462 (
		_w23951_,
		_w23952_,
		_w23974_
	);
	LUT2 #(
		.INIT('h8)
	) name13463 (
		_w23949_,
		_w23950_,
		_w23975_
	);
	LUT2 #(
		.INIT('h8)
	) name13464 (
		_w23947_,
		_w23948_,
		_w23976_
	);
	LUT2 #(
		.INIT('h8)
	) name13465 (
		_w23945_,
		_w23946_,
		_w23977_
	);
	LUT2 #(
		.INIT('h8)
	) name13466 (
		_w23943_,
		_w23944_,
		_w23978_
	);
	LUT2 #(
		.INIT('h8)
	) name13467 (
		_w23941_,
		_w23942_,
		_w23979_
	);
	LUT2 #(
		.INIT('h8)
	) name13468 (
		_w23939_,
		_w23940_,
		_w23980_
	);
	LUT2 #(
		.INIT('h8)
	) name13469 (
		_w23937_,
		_w23938_,
		_w23981_
	);
	LUT2 #(
		.INIT('h8)
	) name13470 (
		_w23935_,
		_w23936_,
		_w23982_
	);
	LUT2 #(
		.INIT('h8)
	) name13471 (
		_w23933_,
		_w23934_,
		_w23983_
	);
	LUT2 #(
		.INIT('h8)
	) name13472 (
		_w23931_,
		_w23932_,
		_w23984_
	);
	LUT2 #(
		.INIT('h8)
	) name13473 (
		_w23929_,
		_w23930_,
		_w23985_
	);
	LUT2 #(
		.INIT('h8)
	) name13474 (
		_w23927_,
		_w23928_,
		_w23986_
	);
	LUT2 #(
		.INIT('h8)
	) name13475 (
		_w23925_,
		_w23926_,
		_w23987_
	);
	LUT2 #(
		.INIT('h8)
	) name13476 (
		_w23923_,
		_w23924_,
		_w23988_
	);
	LUT2 #(
		.INIT('h8)
	) name13477 (
		_w23921_,
		_w23922_,
		_w23989_
	);
	LUT2 #(
		.INIT('h8)
	) name13478 (
		_w23919_,
		_w23920_,
		_w23990_
	);
	LUT2 #(
		.INIT('h8)
	) name13479 (
		_w23917_,
		_w23918_,
		_w23991_
	);
	LUT2 #(
		.INIT('h8)
	) name13480 (
		_w23915_,
		_w23916_,
		_w23992_
	);
	LUT2 #(
		.INIT('h8)
	) name13481 (
		_w23913_,
		_w23914_,
		_w23993_
	);
	LUT2 #(
		.INIT('h8)
	) name13482 (
		_w23911_,
		_w23912_,
		_w23994_
	);
	LUT2 #(
		.INIT('h8)
	) name13483 (
		_w23909_,
		_w23910_,
		_w23995_
	);
	LUT2 #(
		.INIT('h8)
	) name13484 (
		_w23907_,
		_w23908_,
		_w23996_
	);
	LUT2 #(
		.INIT('h8)
	) name13485 (
		_w23905_,
		_w23906_,
		_w23997_
	);
	LUT2 #(
		.INIT('h8)
	) name13486 (
		_w23903_,
		_w23904_,
		_w23998_
	);
	LUT2 #(
		.INIT('h8)
	) name13487 (
		_w23901_,
		_w23902_,
		_w23999_
	);
	LUT2 #(
		.INIT('h8)
	) name13488 (
		_w23899_,
		_w23900_,
		_w24000_
	);
	LUT2 #(
		.INIT('h8)
	) name13489 (
		_w23897_,
		_w23898_,
		_w24001_
	);
	LUT2 #(
		.INIT('h8)
	) name13490 (
		_w23895_,
		_w23896_,
		_w24002_
	);
	LUT2 #(
		.INIT('h8)
	) name13491 (
		_w23893_,
		_w23894_,
		_w24003_
	);
	LUT2 #(
		.INIT('h8)
	) name13492 (
		_w23891_,
		_w23892_,
		_w24004_
	);
	LUT2 #(
		.INIT('h8)
	) name13493 (
		_w23889_,
		_w23890_,
		_w24005_
	);
	LUT2 #(
		.INIT('h8)
	) name13494 (
		_w23887_,
		_w23888_,
		_w24006_
	);
	LUT2 #(
		.INIT('h8)
	) name13495 (
		_w23885_,
		_w23886_,
		_w24007_
	);
	LUT2 #(
		.INIT('h8)
	) name13496 (
		_w23883_,
		_w23884_,
		_w24008_
	);
	LUT2 #(
		.INIT('h8)
	) name13497 (
		_w23881_,
		_w23882_,
		_w24009_
	);
	LUT2 #(
		.INIT('h8)
	) name13498 (
		_w23879_,
		_w23880_,
		_w24010_
	);
	LUT2 #(
		.INIT('h8)
	) name13499 (
		_w23877_,
		_w23878_,
		_w24011_
	);
	LUT2 #(
		.INIT('h8)
	) name13500 (
		_w23875_,
		_w23876_,
		_w24012_
	);
	LUT2 #(
		.INIT('h8)
	) name13501 (
		_w23873_,
		_w23874_,
		_w24013_
	);
	LUT2 #(
		.INIT('h8)
	) name13502 (
		_w23871_,
		_w23872_,
		_w24014_
	);
	LUT2 #(
		.INIT('h8)
	) name13503 (
		_w23869_,
		_w23870_,
		_w24015_
	);
	LUT2 #(
		.INIT('h8)
	) name13504 (
		_w23867_,
		_w23868_,
		_w24016_
	);
	LUT2 #(
		.INIT('h8)
	) name13505 (
		_w23865_,
		_w23866_,
		_w24017_
	);
	LUT2 #(
		.INIT('h8)
	) name13506 (
		_w23863_,
		_w23864_,
		_w24018_
	);
	LUT2 #(
		.INIT('h8)
	) name13507 (
		_w23861_,
		_w23862_,
		_w24019_
	);
	LUT2 #(
		.INIT('h8)
	) name13508 (
		_w23859_,
		_w23860_,
		_w24020_
	);
	LUT2 #(
		.INIT('h8)
	) name13509 (
		_w23857_,
		_w23858_,
		_w24021_
	);
	LUT2 #(
		.INIT('h8)
	) name13510 (
		_w23855_,
		_w23856_,
		_w24022_
	);
	LUT2 #(
		.INIT('h8)
	) name13511 (
		_w23853_,
		_w23854_,
		_w24023_
	);
	LUT2 #(
		.INIT('h8)
	) name13512 (
		_w23851_,
		_w23852_,
		_w24024_
	);
	LUT2 #(
		.INIT('h8)
	) name13513 (
		_w23849_,
		_w23850_,
		_w24025_
	);
	LUT2 #(
		.INIT('h8)
	) name13514 (
		_w23847_,
		_w23848_,
		_w24026_
	);
	LUT2 #(
		.INIT('h8)
	) name13515 (
		_w23845_,
		_w23846_,
		_w24027_
	);
	LUT2 #(
		.INIT('h8)
	) name13516 (
		_w23843_,
		_w23844_,
		_w24028_
	);
	LUT2 #(
		.INIT('h8)
	) name13517 (
		_w23841_,
		_w23842_,
		_w24029_
	);
	LUT2 #(
		.INIT('h8)
	) name13518 (
		_w23839_,
		_w23840_,
		_w24030_
	);
	LUT2 #(
		.INIT('h8)
	) name13519 (
		_w24029_,
		_w24030_,
		_w24031_
	);
	LUT2 #(
		.INIT('h8)
	) name13520 (
		_w24027_,
		_w24028_,
		_w24032_
	);
	LUT2 #(
		.INIT('h8)
	) name13521 (
		_w24025_,
		_w24026_,
		_w24033_
	);
	LUT2 #(
		.INIT('h8)
	) name13522 (
		_w24023_,
		_w24024_,
		_w24034_
	);
	LUT2 #(
		.INIT('h8)
	) name13523 (
		_w24021_,
		_w24022_,
		_w24035_
	);
	LUT2 #(
		.INIT('h8)
	) name13524 (
		_w24019_,
		_w24020_,
		_w24036_
	);
	LUT2 #(
		.INIT('h8)
	) name13525 (
		_w24017_,
		_w24018_,
		_w24037_
	);
	LUT2 #(
		.INIT('h8)
	) name13526 (
		_w24015_,
		_w24016_,
		_w24038_
	);
	LUT2 #(
		.INIT('h8)
	) name13527 (
		_w24013_,
		_w24014_,
		_w24039_
	);
	LUT2 #(
		.INIT('h8)
	) name13528 (
		_w24011_,
		_w24012_,
		_w24040_
	);
	LUT2 #(
		.INIT('h8)
	) name13529 (
		_w24009_,
		_w24010_,
		_w24041_
	);
	LUT2 #(
		.INIT('h8)
	) name13530 (
		_w24007_,
		_w24008_,
		_w24042_
	);
	LUT2 #(
		.INIT('h8)
	) name13531 (
		_w24005_,
		_w24006_,
		_w24043_
	);
	LUT2 #(
		.INIT('h8)
	) name13532 (
		_w24003_,
		_w24004_,
		_w24044_
	);
	LUT2 #(
		.INIT('h8)
	) name13533 (
		_w24001_,
		_w24002_,
		_w24045_
	);
	LUT2 #(
		.INIT('h8)
	) name13534 (
		_w23999_,
		_w24000_,
		_w24046_
	);
	LUT2 #(
		.INIT('h8)
	) name13535 (
		_w23997_,
		_w23998_,
		_w24047_
	);
	LUT2 #(
		.INIT('h8)
	) name13536 (
		_w23995_,
		_w23996_,
		_w24048_
	);
	LUT2 #(
		.INIT('h8)
	) name13537 (
		_w23993_,
		_w23994_,
		_w24049_
	);
	LUT2 #(
		.INIT('h8)
	) name13538 (
		_w23991_,
		_w23992_,
		_w24050_
	);
	LUT2 #(
		.INIT('h8)
	) name13539 (
		_w23989_,
		_w23990_,
		_w24051_
	);
	LUT2 #(
		.INIT('h8)
	) name13540 (
		_w23987_,
		_w23988_,
		_w24052_
	);
	LUT2 #(
		.INIT('h8)
	) name13541 (
		_w23985_,
		_w23986_,
		_w24053_
	);
	LUT2 #(
		.INIT('h8)
	) name13542 (
		_w23983_,
		_w23984_,
		_w24054_
	);
	LUT2 #(
		.INIT('h8)
	) name13543 (
		_w23981_,
		_w23982_,
		_w24055_
	);
	LUT2 #(
		.INIT('h8)
	) name13544 (
		_w23979_,
		_w23980_,
		_w24056_
	);
	LUT2 #(
		.INIT('h8)
	) name13545 (
		_w23977_,
		_w23978_,
		_w24057_
	);
	LUT2 #(
		.INIT('h8)
	) name13546 (
		_w23975_,
		_w23976_,
		_w24058_
	);
	LUT2 #(
		.INIT('h8)
	) name13547 (
		_w23973_,
		_w23974_,
		_w24059_
	);
	LUT2 #(
		.INIT('h8)
	) name13548 (
		_w23971_,
		_w23972_,
		_w24060_
	);
	LUT2 #(
		.INIT('h8)
	) name13549 (
		_w23969_,
		_w23970_,
		_w24061_
	);
	LUT2 #(
		.INIT('h8)
	) name13550 (
		_w23967_,
		_w23968_,
		_w24062_
	);
	LUT2 #(
		.INIT('h8)
	) name13551 (
		_w24061_,
		_w24062_,
		_w24063_
	);
	LUT2 #(
		.INIT('h8)
	) name13552 (
		_w24059_,
		_w24060_,
		_w24064_
	);
	LUT2 #(
		.INIT('h8)
	) name13553 (
		_w24057_,
		_w24058_,
		_w24065_
	);
	LUT2 #(
		.INIT('h8)
	) name13554 (
		_w24055_,
		_w24056_,
		_w24066_
	);
	LUT2 #(
		.INIT('h8)
	) name13555 (
		_w24053_,
		_w24054_,
		_w24067_
	);
	LUT2 #(
		.INIT('h8)
	) name13556 (
		_w24051_,
		_w24052_,
		_w24068_
	);
	LUT2 #(
		.INIT('h8)
	) name13557 (
		_w24049_,
		_w24050_,
		_w24069_
	);
	LUT2 #(
		.INIT('h8)
	) name13558 (
		_w24047_,
		_w24048_,
		_w24070_
	);
	LUT2 #(
		.INIT('h8)
	) name13559 (
		_w24045_,
		_w24046_,
		_w24071_
	);
	LUT2 #(
		.INIT('h8)
	) name13560 (
		_w24043_,
		_w24044_,
		_w24072_
	);
	LUT2 #(
		.INIT('h8)
	) name13561 (
		_w24041_,
		_w24042_,
		_w24073_
	);
	LUT2 #(
		.INIT('h8)
	) name13562 (
		_w24039_,
		_w24040_,
		_w24074_
	);
	LUT2 #(
		.INIT('h8)
	) name13563 (
		_w24037_,
		_w24038_,
		_w24075_
	);
	LUT2 #(
		.INIT('h8)
	) name13564 (
		_w24035_,
		_w24036_,
		_w24076_
	);
	LUT2 #(
		.INIT('h8)
	) name13565 (
		_w24033_,
		_w24034_,
		_w24077_
	);
	LUT2 #(
		.INIT('h8)
	) name13566 (
		_w24031_,
		_w24032_,
		_w24078_
	);
	LUT2 #(
		.INIT('h8)
	) name13567 (
		_w24077_,
		_w24078_,
		_w24079_
	);
	LUT2 #(
		.INIT('h8)
	) name13568 (
		_w24075_,
		_w24076_,
		_w24080_
	);
	LUT2 #(
		.INIT('h8)
	) name13569 (
		_w24073_,
		_w24074_,
		_w24081_
	);
	LUT2 #(
		.INIT('h8)
	) name13570 (
		_w24071_,
		_w24072_,
		_w24082_
	);
	LUT2 #(
		.INIT('h8)
	) name13571 (
		_w24069_,
		_w24070_,
		_w24083_
	);
	LUT2 #(
		.INIT('h8)
	) name13572 (
		_w24067_,
		_w24068_,
		_w24084_
	);
	LUT2 #(
		.INIT('h8)
	) name13573 (
		_w24065_,
		_w24066_,
		_w24085_
	);
	LUT2 #(
		.INIT('h8)
	) name13574 (
		_w24063_,
		_w24064_,
		_w24086_
	);
	LUT2 #(
		.INIT('h8)
	) name13575 (
		_w24085_,
		_w24086_,
		_w24087_
	);
	LUT2 #(
		.INIT('h8)
	) name13576 (
		_w24083_,
		_w24084_,
		_w24088_
	);
	LUT2 #(
		.INIT('h8)
	) name13577 (
		_w24081_,
		_w24082_,
		_w24089_
	);
	LUT2 #(
		.INIT('h8)
	) name13578 (
		_w24079_,
		_w24080_,
		_w24090_
	);
	LUT2 #(
		.INIT('h8)
	) name13579 (
		_w24089_,
		_w24090_,
		_w24091_
	);
	LUT2 #(
		.INIT('h8)
	) name13580 (
		_w24087_,
		_w24088_,
		_w24092_
	);
	LUT2 #(
		.INIT('h8)
	) name13581 (
		_w24091_,
		_w24092_,
		_w24093_
	);
	LUT2 #(
		.INIT('h1)
	) name13582 (
		wb_rst_i_pad,
		_w24093_,
		_w24094_
	);
	LUT2 #(
		.INIT('h8)
	) name13583 (
		_w17883_,
		_w24094_,
		_w24095_
	);
	LUT2 #(
		.INIT('h1)
	) name13584 (
		_w23582_,
		_w24095_,
		_w24096_
	);
	LUT2 #(
		.INIT('h2)
	) name13585 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		_w17883_,
		_w24097_
	);
	LUT2 #(
		.INIT('h1)
	) name13586 (
		_w24095_,
		_w24097_,
		_w24098_
	);
	LUT2 #(
		.INIT('h8)
	) name13587 (
		\wishbone_TxPointerLSB_rst_reg[1]/NET0131 ,
		_w23581_,
		_w24099_
	);
	LUT2 #(
		.INIT('h1)
	) name13588 (
		_w23579_,
		_w24099_,
		_w24100_
	);
	LUT2 #(
		.INIT('h1)
	) name13589 (
		_w22415_,
		_w22944_,
		_w24101_
	);
	LUT2 #(
		.INIT('h8)
	) name13590 (
		\ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 ,
		_w22952_,
		_w24102_
	);
	LUT2 #(
		.INIT('h8)
	) name13591 (
		\ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 ,
		_w22956_,
		_w24103_
	);
	LUT2 #(
		.INIT('h8)
	) name13592 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		_w22959_,
		_w24104_
	);
	LUT2 #(
		.INIT('h8)
	) name13593 (
		\ethreg1_PACKETLEN_2_DataOut_reg[7]/NET0131 ,
		_w22966_,
		_w24105_
	);
	LUT2 #(
		.INIT('h1)
	) name13594 (
		_w24102_,
		_w24103_,
		_w24106_
	);
	LUT2 #(
		.INIT('h4)
	) name13595 (
		_w24104_,
		_w24106_,
		_w24107_
	);
	LUT2 #(
		.INIT('h8)
	) name13596 (
		_w22944_,
		_w24107_,
		_w24108_
	);
	LUT2 #(
		.INIT('h4)
	) name13597 (
		_w24105_,
		_w24108_,
		_w24109_
	);
	LUT2 #(
		.INIT('h1)
	) name13598 (
		_w24101_,
		_w24109_,
		_w24110_
	);
	LUT2 #(
		.INIT('h1)
	) name13599 (
		_w15110_,
		_w22944_,
		_w24111_
	);
	LUT2 #(
		.INIT('h8)
	) name13600 (
		\ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 ,
		_w22952_,
		_w24112_
	);
	LUT2 #(
		.INIT('h8)
	) name13601 (
		\ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 ,
		_w22956_,
		_w24113_
	);
	LUT2 #(
		.INIT('h8)
	) name13602 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		_w22959_,
		_w24114_
	);
	LUT2 #(
		.INIT('h8)
	) name13603 (
		\ethreg1_PACKETLEN_3_DataOut_reg[0]/NET0131 ,
		_w22966_,
		_w24115_
	);
	LUT2 #(
		.INIT('h1)
	) name13604 (
		_w24112_,
		_w24113_,
		_w24116_
	);
	LUT2 #(
		.INIT('h4)
	) name13605 (
		_w24114_,
		_w24116_,
		_w24117_
	);
	LUT2 #(
		.INIT('h8)
	) name13606 (
		_w22944_,
		_w24117_,
		_w24118_
	);
	LUT2 #(
		.INIT('h4)
	) name13607 (
		_w24115_,
		_w24118_,
		_w24119_
	);
	LUT2 #(
		.INIT('h1)
	) name13608 (
		_w24111_,
		_w24119_,
		_w24120_
	);
	LUT2 #(
		.INIT('h1)
	) name13609 (
		_w17810_,
		_w22944_,
		_w24121_
	);
	LUT2 #(
		.INIT('h8)
	) name13610 (
		\ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 ,
		_w22952_,
		_w24122_
	);
	LUT2 #(
		.INIT('h8)
	) name13611 (
		\ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 ,
		_w22956_,
		_w24123_
	);
	LUT2 #(
		.INIT('h8)
	) name13612 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		_w22959_,
		_w24124_
	);
	LUT2 #(
		.INIT('h8)
	) name13613 (
		\ethreg1_PACKETLEN_3_DataOut_reg[1]/NET0131 ,
		_w22966_,
		_w24125_
	);
	LUT2 #(
		.INIT('h1)
	) name13614 (
		_w24122_,
		_w24123_,
		_w24126_
	);
	LUT2 #(
		.INIT('h4)
	) name13615 (
		_w24124_,
		_w24126_,
		_w24127_
	);
	LUT2 #(
		.INIT('h8)
	) name13616 (
		_w22944_,
		_w24127_,
		_w24128_
	);
	LUT2 #(
		.INIT('h4)
	) name13617 (
		_w24125_,
		_w24128_,
		_w24129_
	);
	LUT2 #(
		.INIT('h1)
	) name13618 (
		_w24121_,
		_w24129_,
		_w24130_
	);
	LUT2 #(
		.INIT('h1)
	) name13619 (
		_w17287_,
		_w22944_,
		_w24131_
	);
	LUT2 #(
		.INIT('h8)
	) name13620 (
		\ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 ,
		_w22952_,
		_w24132_
	);
	LUT2 #(
		.INIT('h8)
	) name13621 (
		\ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 ,
		_w22956_,
		_w24133_
	);
	LUT2 #(
		.INIT('h8)
	) name13622 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		_w22959_,
		_w24134_
	);
	LUT2 #(
		.INIT('h8)
	) name13623 (
		\ethreg1_PACKETLEN_3_DataOut_reg[2]/NET0131 ,
		_w22966_,
		_w24135_
	);
	LUT2 #(
		.INIT('h1)
	) name13624 (
		_w24132_,
		_w24133_,
		_w24136_
	);
	LUT2 #(
		.INIT('h4)
	) name13625 (
		_w24134_,
		_w24136_,
		_w24137_
	);
	LUT2 #(
		.INIT('h8)
	) name13626 (
		_w22944_,
		_w24137_,
		_w24138_
	);
	LUT2 #(
		.INIT('h4)
	) name13627 (
		_w24135_,
		_w24138_,
		_w24139_
	);
	LUT2 #(
		.INIT('h1)
	) name13628 (
		_w24131_,
		_w24139_,
		_w24140_
	);
	LUT2 #(
		.INIT('h1)
	) name13629 (
		_w20856_,
		_w22944_,
		_w24141_
	);
	LUT2 #(
		.INIT('h8)
	) name13630 (
		\ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 ,
		_w22952_,
		_w24142_
	);
	LUT2 #(
		.INIT('h8)
	) name13631 (
		\ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 ,
		_w22956_,
		_w24143_
	);
	LUT2 #(
		.INIT('h8)
	) name13632 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		_w22959_,
		_w24144_
	);
	LUT2 #(
		.INIT('h8)
	) name13633 (
		\ethreg1_PACKETLEN_3_DataOut_reg[3]/NET0131 ,
		_w22966_,
		_w24145_
	);
	LUT2 #(
		.INIT('h1)
	) name13634 (
		_w24142_,
		_w24143_,
		_w24146_
	);
	LUT2 #(
		.INIT('h4)
	) name13635 (
		_w24144_,
		_w24146_,
		_w24147_
	);
	LUT2 #(
		.INIT('h8)
	) name13636 (
		_w22944_,
		_w24147_,
		_w24148_
	);
	LUT2 #(
		.INIT('h4)
	) name13637 (
		_w24145_,
		_w24148_,
		_w24149_
	);
	LUT2 #(
		.INIT('h1)
	) name13638 (
		_w24141_,
		_w24149_,
		_w24150_
	);
	LUT2 #(
		.INIT('h1)
	) name13639 (
		_w13475_,
		_w22944_,
		_w24151_
	);
	LUT2 #(
		.INIT('h8)
	) name13640 (
		\ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 ,
		_w22952_,
		_w24152_
	);
	LUT2 #(
		.INIT('h8)
	) name13641 (
		\ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 ,
		_w22956_,
		_w24153_
	);
	LUT2 #(
		.INIT('h8)
	) name13642 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		_w22959_,
		_w24154_
	);
	LUT2 #(
		.INIT('h8)
	) name13643 (
		\ethreg1_PACKETLEN_3_DataOut_reg[4]/NET0131 ,
		_w22966_,
		_w24155_
	);
	LUT2 #(
		.INIT('h1)
	) name13644 (
		_w24152_,
		_w24153_,
		_w24156_
	);
	LUT2 #(
		.INIT('h4)
	) name13645 (
		_w24154_,
		_w24156_,
		_w24157_
	);
	LUT2 #(
		.INIT('h8)
	) name13646 (
		_w22944_,
		_w24157_,
		_w24158_
	);
	LUT2 #(
		.INIT('h4)
	) name13647 (
		_w24155_,
		_w24158_,
		_w24159_
	);
	LUT2 #(
		.INIT('h1)
	) name13648 (
		_w24151_,
		_w24159_,
		_w24160_
	);
	LUT2 #(
		.INIT('h1)
	) name13649 (
		_w14019_,
		_w22944_,
		_w24161_
	);
	LUT2 #(
		.INIT('h8)
	) name13650 (
		\ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 ,
		_w22952_,
		_w24162_
	);
	LUT2 #(
		.INIT('h8)
	) name13651 (
		\ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 ,
		_w22956_,
		_w24163_
	);
	LUT2 #(
		.INIT('h8)
	) name13652 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		_w22959_,
		_w24164_
	);
	LUT2 #(
		.INIT('h8)
	) name13653 (
		\ethreg1_PACKETLEN_3_DataOut_reg[5]/NET0131 ,
		_w22966_,
		_w24165_
	);
	LUT2 #(
		.INIT('h1)
	) name13654 (
		_w24162_,
		_w24163_,
		_w24166_
	);
	LUT2 #(
		.INIT('h4)
	) name13655 (
		_w24164_,
		_w24166_,
		_w24167_
	);
	LUT2 #(
		.INIT('h8)
	) name13656 (
		_w22944_,
		_w24167_,
		_w24168_
	);
	LUT2 #(
		.INIT('h4)
	) name13657 (
		_w24165_,
		_w24168_,
		_w24169_
	);
	LUT2 #(
		.INIT('h1)
	) name13658 (
		_w24161_,
		_w24169_,
		_w24170_
	);
	LUT2 #(
		.INIT('h8)
	) name13659 (
		m_wb_we_o_pad,
		_w12573_,
		_w24171_
	);
	LUT2 #(
		.INIT('h2)
	) name13660 (
		_w12632_,
		_w24171_,
		_w24172_
	);
	LUT2 #(
		.INIT('h1)
	) name13661 (
		_w14536_,
		_w22944_,
		_w24173_
	);
	LUT2 #(
		.INIT('h8)
	) name13662 (
		\ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 ,
		_w22952_,
		_w24174_
	);
	LUT2 #(
		.INIT('h8)
	) name13663 (
		\ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 ,
		_w22956_,
		_w24175_
	);
	LUT2 #(
		.INIT('h8)
	) name13664 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		_w22959_,
		_w24176_
	);
	LUT2 #(
		.INIT('h8)
	) name13665 (
		\ethreg1_PACKETLEN_3_DataOut_reg[6]/NET0131 ,
		_w22966_,
		_w24177_
	);
	LUT2 #(
		.INIT('h1)
	) name13666 (
		_w24174_,
		_w24175_,
		_w24178_
	);
	LUT2 #(
		.INIT('h4)
	) name13667 (
		_w24176_,
		_w24178_,
		_w24179_
	);
	LUT2 #(
		.INIT('h8)
	) name13668 (
		_w22944_,
		_w24179_,
		_w24180_
	);
	LUT2 #(
		.INIT('h4)
	) name13669 (
		_w24177_,
		_w24180_,
		_w24181_
	);
	LUT2 #(
		.INIT('h1)
	) name13670 (
		_w24173_,
		_w24181_,
		_w24182_
	);
	LUT2 #(
		.INIT('h1)
	) name13671 (
		_w19604_,
		_w22944_,
		_w24183_
	);
	LUT2 #(
		.INIT('h8)
	) name13672 (
		\ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 ,
		_w22952_,
		_w24184_
	);
	LUT2 #(
		.INIT('h8)
	) name13673 (
		\ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 ,
		_w22956_,
		_w24185_
	);
	LUT2 #(
		.INIT('h8)
	) name13674 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		_w22959_,
		_w24186_
	);
	LUT2 #(
		.INIT('h8)
	) name13675 (
		\ethreg1_PACKETLEN_3_DataOut_reg[7]/NET0131 ,
		_w22966_,
		_w24187_
	);
	LUT2 #(
		.INIT('h1)
	) name13676 (
		_w24184_,
		_w24185_,
		_w24188_
	);
	LUT2 #(
		.INIT('h4)
	) name13677 (
		_w24186_,
		_w24188_,
		_w24189_
	);
	LUT2 #(
		.INIT('h8)
	) name13678 (
		_w22944_,
		_w24189_,
		_w24190_
	);
	LUT2 #(
		.INIT('h4)
	) name13679 (
		_w24187_,
		_w24190_,
		_w24191_
	);
	LUT2 #(
		.INIT('h1)
	) name13680 (
		_w24183_,
		_w24191_,
		_w24192_
	);
	LUT2 #(
		.INIT('h8)
	) name13681 (
		\wishbone_bd_ram_mem0_reg[17][3]/P0001 ,
		_w12848_,
		_w24193_
	);
	LUT2 #(
		.INIT('h8)
	) name13682 (
		\wishbone_bd_ram_mem0_reg[57][3]/P0001 ,
		_w13116_,
		_w24194_
	);
	LUT2 #(
		.INIT('h8)
	) name13683 (
		\wishbone_bd_ram_mem0_reg[40][3]/P0001 ,
		_w13132_,
		_w24195_
	);
	LUT2 #(
		.INIT('h8)
	) name13684 (
		\wishbone_bd_ram_mem0_reg[182][3]/P0001 ,
		_w12820_,
		_w24196_
	);
	LUT2 #(
		.INIT('h8)
	) name13685 (
		\wishbone_bd_ram_mem0_reg[86][3]/P0001 ,
		_w12735_,
		_w24197_
	);
	LUT2 #(
		.INIT('h8)
	) name13686 (
		\wishbone_bd_ram_mem0_reg[236][3]/P0001 ,
		_w12731_,
		_w24198_
	);
	LUT2 #(
		.INIT('h8)
	) name13687 (
		\wishbone_bd_ram_mem0_reg[160][3]/P0001 ,
		_w12872_,
		_w24199_
	);
	LUT2 #(
		.INIT('h8)
	) name13688 (
		\wishbone_bd_ram_mem0_reg[32][3]/P0001 ,
		_w13120_,
		_w24200_
	);
	LUT2 #(
		.INIT('h8)
	) name13689 (
		\wishbone_bd_ram_mem0_reg[189][3]/P0001 ,
		_w13042_,
		_w24201_
	);
	LUT2 #(
		.INIT('h8)
	) name13690 (
		\wishbone_bd_ram_mem0_reg[248][3]/P0001 ,
		_w12789_,
		_w24202_
	);
	LUT2 #(
		.INIT('h8)
	) name13691 (
		\wishbone_bd_ram_mem0_reg[79][3]/P0001 ,
		_w13212_,
		_w24203_
	);
	LUT2 #(
		.INIT('h8)
	) name13692 (
		\wishbone_bd_ram_mem0_reg[167][3]/P0001 ,
		_w12986_,
		_w24204_
	);
	LUT2 #(
		.INIT('h8)
	) name13693 (
		\wishbone_bd_ram_mem0_reg[9][3]/P0001 ,
		_w12808_,
		_w24205_
	);
	LUT2 #(
		.INIT('h8)
	) name13694 (
		\wishbone_bd_ram_mem0_reg[92][3]/P0001 ,
		_w13010_,
		_w24206_
	);
	LUT2 #(
		.INIT('h8)
	) name13695 (
		\wishbone_bd_ram_mem0_reg[39][3]/P0001 ,
		_w13018_,
		_w24207_
	);
	LUT2 #(
		.INIT('h8)
	) name13696 (
		\wishbone_bd_ram_mem0_reg[28][3]/P0001 ,
		_w13170_,
		_w24208_
	);
	LUT2 #(
		.INIT('h8)
	) name13697 (
		\wishbone_bd_ram_mem0_reg[212][3]/P0001 ,
		_w12796_,
		_w24209_
	);
	LUT2 #(
		.INIT('h8)
	) name13698 (
		\wishbone_bd_ram_mem0_reg[241][3]/P0001 ,
		_w13006_,
		_w24210_
	);
	LUT2 #(
		.INIT('h8)
	) name13699 (
		\wishbone_bd_ram_mem0_reg[85][3]/P0001 ,
		_w13216_,
		_w24211_
	);
	LUT2 #(
		.INIT('h8)
	) name13700 (
		\wishbone_bd_ram_mem0_reg[65][3]/P0001 ,
		_w13176_,
		_w24212_
	);
	LUT2 #(
		.INIT('h8)
	) name13701 (
		\wishbone_bd_ram_mem0_reg[148][3]/P0001 ,
		_w13000_,
		_w24213_
	);
	LUT2 #(
		.INIT('h8)
	) name13702 (
		\wishbone_bd_ram_mem0_reg[202][3]/P0001 ,
		_w12870_,
		_w24214_
	);
	LUT2 #(
		.INIT('h8)
	) name13703 (
		\wishbone_bd_ram_mem0_reg[244][3]/P0001 ,
		_w12747_,
		_w24215_
	);
	LUT2 #(
		.INIT('h8)
	) name13704 (
		\wishbone_bd_ram_mem0_reg[125][3]/P0001 ,
		_w12956_,
		_w24216_
	);
	LUT2 #(
		.INIT('h8)
	) name13705 (
		\wishbone_bd_ram_mem0_reg[87][3]/P0001 ,
		_w13154_,
		_w24217_
	);
	LUT2 #(
		.INIT('h8)
	) name13706 (
		\wishbone_bd_ram_mem0_reg[135][3]/P0001 ,
		_w13124_,
		_w24218_
	);
	LUT2 #(
		.INIT('h8)
	) name13707 (
		\wishbone_bd_ram_mem0_reg[98][3]/P0001 ,
		_w12816_,
		_w24219_
	);
	LUT2 #(
		.INIT('h8)
	) name13708 (
		\wishbone_bd_ram_mem0_reg[198][3]/P0001 ,
		_w12832_,
		_w24220_
	);
	LUT2 #(
		.INIT('h8)
	) name13709 (
		\wishbone_bd_ram_mem0_reg[186][3]/P0001 ,
		_w12783_,
		_w24221_
	);
	LUT2 #(
		.INIT('h8)
	) name13710 (
		\wishbone_bd_ram_mem0_reg[101][3]/P0001 ,
		_w13192_,
		_w24222_
	);
	LUT2 #(
		.INIT('h8)
	) name13711 (
		\wishbone_bd_ram_mem0_reg[210][3]/P0001 ,
		_w12924_,
		_w24223_
	);
	LUT2 #(
		.INIT('h8)
	) name13712 (
		\wishbone_bd_ram_mem0_reg[140][3]/P0001 ,
		_w12894_,
		_w24224_
	);
	LUT2 #(
		.INIT('h8)
	) name13713 (
		\wishbone_bd_ram_mem0_reg[150][3]/P0001 ,
		_w13136_,
		_w24225_
	);
	LUT2 #(
		.INIT('h8)
	) name13714 (
		\wishbone_bd_ram_mem0_reg[207][3]/P0001 ,
		_w13180_,
		_w24226_
	);
	LUT2 #(
		.INIT('h8)
	) name13715 (
		\wishbone_bd_ram_mem0_reg[7][3]/P0001 ,
		_w12728_,
		_w24227_
	);
	LUT2 #(
		.INIT('h8)
	) name13716 (
		\wishbone_bd_ram_mem0_reg[142][3]/P0001 ,
		_w12928_,
		_w24228_
	);
	LUT2 #(
		.INIT('h8)
	) name13717 (
		\wishbone_bd_ram_mem0_reg[131][3]/P0001 ,
		_w12852_,
		_w24229_
	);
	LUT2 #(
		.INIT('h8)
	) name13718 (
		\wishbone_bd_ram_mem0_reg[155][3]/P0001 ,
		_w13122_,
		_w24230_
	);
	LUT2 #(
		.INIT('h8)
	) name13719 (
		\wishbone_bd_ram_mem0_reg[222][3]/P0001 ,
		_w13094_,
		_w24231_
	);
	LUT2 #(
		.INIT('h8)
	) name13720 (
		\wishbone_bd_ram_mem0_reg[46][3]/P0001 ,
		_w12884_,
		_w24232_
	);
	LUT2 #(
		.INIT('h8)
	) name13721 (
		\wishbone_bd_ram_mem0_reg[242][3]/P0001 ,
		_w12932_,
		_w24233_
	);
	LUT2 #(
		.INIT('h8)
	) name13722 (
		\wishbone_bd_ram_mem0_reg[238][3]/P0001 ,
		_w13160_,
		_w24234_
	);
	LUT2 #(
		.INIT('h8)
	) name13723 (
		\wishbone_bd_ram_mem0_reg[130][3]/P0001 ,
		_w12914_,
		_w24235_
	);
	LUT2 #(
		.INIT('h8)
	) name13724 (
		\wishbone_bd_ram_mem0_reg[141][3]/P0001 ,
		_w13004_,
		_w24236_
	);
	LUT2 #(
		.INIT('h8)
	) name13725 (
		\wishbone_bd_ram_mem0_reg[235][3]/P0001 ,
		_w12696_,
		_w24237_
	);
	LUT2 #(
		.INIT('h8)
	) name13726 (
		\wishbone_bd_ram_mem0_reg[99][3]/P0001 ,
		_w13038_,
		_w24238_
	);
	LUT2 #(
		.INIT('h8)
	) name13727 (
		\wishbone_bd_ram_mem0_reg[147][3]/P0001 ,
		_w13146_,
		_w24239_
	);
	LUT2 #(
		.INIT('h8)
	) name13728 (
		\wishbone_bd_ram_mem0_reg[206][3]/P0001 ,
		_w12954_,
		_w24240_
	);
	LUT2 #(
		.INIT('h8)
	) name13729 (
		\wishbone_bd_ram_mem0_reg[199][3]/P0001 ,
		_w12768_,
		_w24241_
	);
	LUT2 #(
		.INIT('h8)
	) name13730 (
		\wishbone_bd_ram_mem0_reg[83][3]/P0001 ,
		_w12916_,
		_w24242_
	);
	LUT2 #(
		.INIT('h8)
	) name13731 (
		\wishbone_bd_ram_mem0_reg[5][3]/P0001 ,
		_w12878_,
		_w24243_
	);
	LUT2 #(
		.INIT('h8)
	) name13732 (
		\wishbone_bd_ram_mem0_reg[78][3]/P0001 ,
		_w12874_,
		_w24244_
	);
	LUT2 #(
		.INIT('h8)
	) name13733 (
		\wishbone_bd_ram_mem0_reg[76][3]/P0001 ,
		_w13184_,
		_w24245_
	);
	LUT2 #(
		.INIT('h8)
	) name13734 (
		\wishbone_bd_ram_mem0_reg[196][3]/P0001 ,
		_w13090_,
		_w24246_
	);
	LUT2 #(
		.INIT('h8)
	) name13735 (
		\wishbone_bd_ram_mem0_reg[151][3]/P0001 ,
		_w13142_,
		_w24247_
	);
	LUT2 #(
		.INIT('h8)
	) name13736 (
		\wishbone_bd_ram_mem0_reg[185][3]/P0001 ,
		_w12940_,
		_w24248_
	);
	LUT2 #(
		.INIT('h8)
	) name13737 (
		\wishbone_bd_ram_mem0_reg[59][3]/P0001 ,
		_w12780_,
		_w24249_
	);
	LUT2 #(
		.INIT('h8)
	) name13738 (
		\wishbone_bd_ram_mem0_reg[249][3]/P0001 ,
		_w12900_,
		_w24250_
	);
	LUT2 #(
		.INIT('h8)
	) name13739 (
		\wishbone_bd_ram_mem0_reg[8][3]/P0001 ,
		_w12920_,
		_w24251_
	);
	LUT2 #(
		.INIT('h8)
	) name13740 (
		\wishbone_bd_ram_mem0_reg[81][3]/P0001 ,
		_w12950_,
		_w24252_
	);
	LUT2 #(
		.INIT('h8)
	) name13741 (
		\wishbone_bd_ram_mem0_reg[221][3]/P0001 ,
		_w12802_,
		_w24253_
	);
	LUT2 #(
		.INIT('h8)
	) name13742 (
		\wishbone_bd_ram_mem0_reg[64][3]/P0001 ,
		_w12976_,
		_w24254_
	);
	LUT2 #(
		.INIT('h8)
	) name13743 (
		\wishbone_bd_ram_mem0_reg[139][3]/P0001 ,
		_w12814_,
		_w24255_
	);
	LUT2 #(
		.INIT('h8)
	) name13744 (
		\wishbone_bd_ram_mem0_reg[243][3]/P0001 ,
		_w12804_,
		_w24256_
	);
	LUT2 #(
		.INIT('h8)
	) name13745 (
		\wishbone_bd_ram_mem0_reg[225][3]/P0001 ,
		_w13092_,
		_w24257_
	);
	LUT2 #(
		.INIT('h8)
	) name13746 (
		\wishbone_bd_ram_mem0_reg[179][3]/P0001 ,
		_w13050_,
		_w24258_
	);
	LUT2 #(
		.INIT('h8)
	) name13747 (
		\wishbone_bd_ram_mem0_reg[216][3]/P0001 ,
		_w13028_,
		_w24259_
	);
	LUT2 #(
		.INIT('h8)
	) name13748 (
		\wishbone_bd_ram_mem0_reg[30][3]/P0001 ,
		_w13104_,
		_w24260_
	);
	LUT2 #(
		.INIT('h8)
	) name13749 (
		\wishbone_bd_ram_mem0_reg[144][3]/P0001 ,
		_w12756_,
		_w24261_
	);
	LUT2 #(
		.INIT('h8)
	) name13750 (
		\wishbone_bd_ram_mem0_reg[153][3]/P0001 ,
		_w12890_,
		_w24262_
	);
	LUT2 #(
		.INIT('h8)
	) name13751 (
		\wishbone_bd_ram_mem0_reg[3][3]/P0001 ,
		_w12866_,
		_w24263_
	);
	LUT2 #(
		.INIT('h8)
	) name13752 (
		\wishbone_bd_ram_mem0_reg[122][3]/P0001 ,
		_w13130_,
		_w24264_
	);
	LUT2 #(
		.INIT('h8)
	) name13753 (
		\wishbone_bd_ram_mem0_reg[14][3]/P0001 ,
		_w13086_,
		_w24265_
	);
	LUT2 #(
		.INIT('h8)
	) name13754 (
		\wishbone_bd_ram_mem0_reg[49][3]/P0001 ,
		_w12994_,
		_w24266_
	);
	LUT2 #(
		.INIT('h8)
	) name13755 (
		\wishbone_bd_ram_mem0_reg[231][3]/P0001 ,
		_w12856_,
		_w24267_
	);
	LUT2 #(
		.INIT('h8)
	) name13756 (
		\wishbone_bd_ram_mem0_reg[226][3]/P0001 ,
		_w13138_,
		_w24268_
	);
	LUT2 #(
		.INIT('h8)
	) name13757 (
		\wishbone_bd_ram_mem0_reg[43][3]/P0001 ,
		_w13200_,
		_w24269_
	);
	LUT2 #(
		.INIT('h8)
	) name13758 (
		\wishbone_bd_ram_mem0_reg[194][3]/P0001 ,
		_w12772_,
		_w24270_
	);
	LUT2 #(
		.INIT('h8)
	) name13759 (
		\wishbone_bd_ram_mem0_reg[229][3]/P0001 ,
		_w12711_,
		_w24271_
	);
	LUT2 #(
		.INIT('h8)
	) name13760 (
		\wishbone_bd_ram_mem0_reg[21][3]/P0001 ,
		_w12906_,
		_w24272_
	);
	LUT2 #(
		.INIT('h8)
	) name13761 (
		\wishbone_bd_ram_mem0_reg[94][3]/P0001 ,
		_w13186_,
		_w24273_
	);
	LUT2 #(
		.INIT('h8)
	) name13762 (
		\wishbone_bd_ram_mem0_reg[97][3]/P0001 ,
		_w13096_,
		_w24274_
	);
	LUT2 #(
		.INIT('h8)
	) name13763 (
		\wishbone_bd_ram_mem0_reg[128][3]/P0001 ,
		_w12793_,
		_w24275_
	);
	LUT2 #(
		.INIT('h8)
	) name13764 (
		\wishbone_bd_ram_mem0_reg[175][3]/P0001 ,
		_w13126_,
		_w24276_
	);
	LUT2 #(
		.INIT('h8)
	) name13765 (
		\wishbone_bd_ram_mem0_reg[209][3]/P0001 ,
		_w13152_,
		_w24277_
	);
	LUT2 #(
		.INIT('h8)
	) name13766 (
		\wishbone_bd_ram_mem0_reg[12][3]/P0001 ,
		_w13118_,
		_w24278_
	);
	LUT2 #(
		.INIT('h8)
	) name13767 (
		\wishbone_bd_ram_mem0_reg[37][3]/P0001 ,
		_w13102_,
		_w24279_
	);
	LUT2 #(
		.INIT('h8)
	) name13768 (
		\wishbone_bd_ram_mem0_reg[162][3]/P0001 ,
		_w13098_,
		_w24280_
	);
	LUT2 #(
		.INIT('h8)
	) name13769 (
		\wishbone_bd_ram_mem0_reg[11][3]/P0001 ,
		_w13194_,
		_w24281_
	);
	LUT2 #(
		.INIT('h8)
	) name13770 (
		\wishbone_bd_ram_mem0_reg[246][3]/P0001 ,
		_w13076_,
		_w24282_
	);
	LUT2 #(
		.INIT('h8)
	) name13771 (
		\wishbone_bd_ram_mem0_reg[115][3]/P0001 ,
		_w13112_,
		_w24283_
	);
	LUT2 #(
		.INIT('h8)
	) name13772 (
		\wishbone_bd_ram_mem0_reg[156][3]/P0001 ,
		_w13190_,
		_w24284_
	);
	LUT2 #(
		.INIT('h8)
	) name13773 (
		\wishbone_bd_ram_mem0_reg[187][3]/P0001 ,
		_w13196_,
		_w24285_
	);
	LUT2 #(
		.INIT('h8)
	) name13774 (
		\wishbone_bd_ram_mem0_reg[197][3]/P0001 ,
		_w12834_,
		_w24286_
	);
	LUT2 #(
		.INIT('h8)
	) name13775 (
		\wishbone_bd_ram_mem0_reg[102][3]/P0001 ,
		_w12685_,
		_w24287_
	);
	LUT2 #(
		.INIT('h8)
	) name13776 (
		\wishbone_bd_ram_mem0_reg[228][3]/P0001 ,
		_w12765_,
		_w24288_
	);
	LUT2 #(
		.INIT('h8)
	) name13777 (
		\wishbone_bd_ram_mem0_reg[239][3]/P0001 ,
		_w12862_,
		_w24289_
	);
	LUT2 #(
		.INIT('h8)
	) name13778 (
		\wishbone_bd_ram_mem0_reg[223][3]/P0001 ,
		_w12838_,
		_w24290_
	);
	LUT2 #(
		.INIT('h8)
	) name13779 (
		\wishbone_bd_ram_mem0_reg[149][3]/P0001 ,
		_w12741_,
		_w24291_
	);
	LUT2 #(
		.INIT('h8)
	) name13780 (
		\wishbone_bd_ram_mem0_reg[4][3]/P0001 ,
		_w12666_,
		_w24292_
	);
	LUT2 #(
		.INIT('h8)
	) name13781 (
		\wishbone_bd_ram_mem0_reg[137][3]/P0001 ,
		_w13168_,
		_w24293_
	);
	LUT2 #(
		.INIT('h8)
	) name13782 (
		\wishbone_bd_ram_mem0_reg[174][3]/P0001 ,
		_w12972_,
		_w24294_
	);
	LUT2 #(
		.INIT('h8)
	) name13783 (
		\wishbone_bd_ram_mem0_reg[164][3]/P0001 ,
		_w12876_,
		_w24295_
	);
	LUT2 #(
		.INIT('h8)
	) name13784 (
		\wishbone_bd_ram_mem0_reg[146][3]/P0001 ,
		_w13060_,
		_w24296_
	);
	LUT2 #(
		.INIT('h8)
	) name13785 (
		\wishbone_bd_ram_mem0_reg[105][3]/P0001 ,
		_w12751_,
		_w24297_
	);
	LUT2 #(
		.INIT('h8)
	) name13786 (
		\wishbone_bd_ram_mem0_reg[74][3]/P0001 ,
		_w12812_,
		_w24298_
	);
	LUT2 #(
		.INIT('h8)
	) name13787 (
		\wishbone_bd_ram_mem0_reg[44][3]/P0001 ,
		_w12896_,
		_w24299_
	);
	LUT2 #(
		.INIT('h8)
	) name13788 (
		\wishbone_bd_ram_mem0_reg[120][3]/P0001 ,
		_w12707_,
		_w24300_
	);
	LUT2 #(
		.INIT('h8)
	) name13789 (
		\wishbone_bd_ram_mem0_reg[133][3]/P0001 ,
		_w12761_,
		_w24301_
	);
	LUT2 #(
		.INIT('h8)
	) name13790 (
		\wishbone_bd_ram_mem0_reg[157][3]/P0001 ,
		_w12926_,
		_w24302_
	);
	LUT2 #(
		.INIT('h8)
	) name13791 (
		\wishbone_bd_ram_mem0_reg[123][3]/P0001 ,
		_w13114_,
		_w24303_
	);
	LUT2 #(
		.INIT('h8)
	) name13792 (
		\wishbone_bd_ram_mem0_reg[38][3]/P0001 ,
		_w13182_,
		_w24304_
	);
	LUT2 #(
		.INIT('h8)
	) name13793 (
		\wishbone_bd_ram_mem0_reg[211][3]/P0001 ,
		_w13166_,
		_w24305_
	);
	LUT2 #(
		.INIT('h8)
	) name13794 (
		\wishbone_bd_ram_mem0_reg[106][3]/P0001 ,
		_w12713_,
		_w24306_
	);
	LUT2 #(
		.INIT('h8)
	) name13795 (
		\wishbone_bd_ram_mem0_reg[190][3]/P0001 ,
		_w12858_,
		_w24307_
	);
	LUT2 #(
		.INIT('h8)
	) name13796 (
		\wishbone_bd_ram_mem0_reg[108][3]/P0001 ,
		_w13156_,
		_w24308_
	);
	LUT2 #(
		.INIT('h8)
	) name13797 (
		\wishbone_bd_ram_mem0_reg[247][3]/P0001 ,
		_w12818_,
		_w24309_
	);
	LUT2 #(
		.INIT('h8)
	) name13798 (
		\wishbone_bd_ram_mem0_reg[93][3]/P0001 ,
		_w13016_,
		_w24310_
	);
	LUT2 #(
		.INIT('h8)
	) name13799 (
		\wishbone_bd_ram_mem0_reg[48][3]/P0001 ,
		_w12970_,
		_w24311_
	);
	LUT2 #(
		.INIT('h8)
	) name13800 (
		\wishbone_bd_ram_mem0_reg[96][3]/P0001 ,
		_w12912_,
		_w24312_
	);
	LUT2 #(
		.INIT('h8)
	) name13801 (
		\wishbone_bd_ram_mem0_reg[111][3]/P0001 ,
		_w12744_,
		_w24313_
	);
	LUT2 #(
		.INIT('h8)
	) name13802 (
		\wishbone_bd_ram_mem0_reg[215][3]/P0001 ,
		_w12974_,
		_w24314_
	);
	LUT2 #(
		.INIT('h8)
	) name13803 (
		\wishbone_bd_ram_mem0_reg[119][3]/P0001 ,
		_w13048_,
		_w24315_
	);
	LUT2 #(
		.INIT('h8)
	) name13804 (
		\wishbone_bd_ram_mem0_reg[181][3]/P0001 ,
		_w12828_,
		_w24316_
	);
	LUT2 #(
		.INIT('h8)
	) name13805 (
		\wishbone_bd_ram_mem0_reg[180][3]/P0001 ,
		_w12791_,
		_w24317_
	);
	LUT2 #(
		.INIT('h8)
	) name13806 (
		\wishbone_bd_ram_mem0_reg[109][3]/P0001 ,
		_w12888_,
		_w24318_
	);
	LUT2 #(
		.INIT('h8)
	) name13807 (
		\wishbone_bd_ram_mem0_reg[117][3]/P0001 ,
		_w12715_,
		_w24319_
	);
	LUT2 #(
		.INIT('h8)
	) name13808 (
		\wishbone_bd_ram_mem0_reg[184][3]/P0001 ,
		_w13062_,
		_w24320_
	);
	LUT2 #(
		.INIT('h8)
	) name13809 (
		\wishbone_bd_ram_mem0_reg[89][3]/P0001 ,
		_w12964_,
		_w24321_
	);
	LUT2 #(
		.INIT('h8)
	) name13810 (
		\wishbone_bd_ram_mem0_reg[54][3]/P0001 ,
		_w12770_,
		_w24322_
	);
	LUT2 #(
		.INIT('h8)
	) name13811 (
		\wishbone_bd_ram_mem0_reg[31][3]/P0001 ,
		_w13198_,
		_w24323_
	);
	LUT2 #(
		.INIT('h8)
	) name13812 (
		\wishbone_bd_ram_mem0_reg[172][3]/P0001 ,
		_w12944_,
		_w24324_
	);
	LUT2 #(
		.INIT('h8)
	) name13813 (
		\wishbone_bd_ram_mem0_reg[90][3]/P0001 ,
		_w12978_,
		_w24325_
	);
	LUT2 #(
		.INIT('h8)
	) name13814 (
		\wishbone_bd_ram_mem0_reg[75][3]/P0001 ,
		_w12826_,
		_w24326_
	);
	LUT2 #(
		.INIT('h8)
	) name13815 (
		\wishbone_bd_ram_mem0_reg[61][3]/P0001 ,
		_w12725_,
		_w24327_
	);
	LUT2 #(
		.INIT('h8)
	) name13816 (
		\wishbone_bd_ram_mem0_reg[171][3]/P0001 ,
		_w12910_,
		_w24328_
	);
	LUT2 #(
		.INIT('h8)
	) name13817 (
		\wishbone_bd_ram_mem0_reg[27][3]/P0001 ,
		_w12880_,
		_w24329_
	);
	LUT2 #(
		.INIT('h8)
	) name13818 (
		\wishbone_bd_ram_mem0_reg[166][3]/P0001 ,
		_w13040_,
		_w24330_
	);
	LUT2 #(
		.INIT('h8)
	) name13819 (
		\wishbone_bd_ram_mem0_reg[53][3]/P0001 ,
		_w13020_,
		_w24331_
	);
	LUT2 #(
		.INIT('h8)
	) name13820 (
		\wishbone_bd_ram_mem0_reg[129][3]/P0001 ,
		_w12776_,
		_w24332_
	);
	LUT2 #(
		.INIT('h8)
	) name13821 (
		\wishbone_bd_ram_mem0_reg[114][3]/P0001 ,
		_w13202_,
		_w24333_
	);
	LUT2 #(
		.INIT('h8)
	) name13822 (
		\wishbone_bd_ram_mem0_reg[237][3]/P0001 ,
		_w12990_,
		_w24334_
	);
	LUT2 #(
		.INIT('h8)
	) name13823 (
		\wishbone_bd_ram_mem0_reg[158][3]/P0001 ,
		_w12898_,
		_w24335_
	);
	LUT2 #(
		.INIT('h8)
	) name13824 (
		\wishbone_bd_ram_mem0_reg[173][3]/P0001 ,
		_w12854_,
		_w24336_
	);
	LUT2 #(
		.INIT('h8)
	) name13825 (
		\wishbone_bd_ram_mem0_reg[121][3]/P0001 ,
		_w13078_,
		_w24337_
	);
	LUT2 #(
		.INIT('h8)
	) name13826 (
		\wishbone_bd_ram_mem0_reg[138][3]/P0001 ,
		_w12958_,
		_w24338_
	);
	LUT2 #(
		.INIT('h8)
	) name13827 (
		\wishbone_bd_ram_mem0_reg[47][3]/P0001 ,
		_w12904_,
		_w24339_
	);
	LUT2 #(
		.INIT('h8)
	) name13828 (
		\wishbone_bd_ram_mem0_reg[251][3]/P0001 ,
		_w13054_,
		_w24340_
	);
	LUT2 #(
		.INIT('h8)
	) name13829 (
		\wishbone_bd_ram_mem0_reg[20][3]/P0001 ,
		_w13174_,
		_w24341_
	);
	LUT2 #(
		.INIT('h8)
	) name13830 (
		\wishbone_bd_ram_mem0_reg[112][3]/P0001 ,
		_w12733_,
		_w24342_
	);
	LUT2 #(
		.INIT('h8)
	) name13831 (
		\wishbone_bd_ram_mem0_reg[208][3]/P0001 ,
		_w13032_,
		_w24343_
	);
	LUT2 #(
		.INIT('h8)
	) name13832 (
		\wishbone_bd_ram_mem0_reg[169][3]/P0001 ,
		_w12722_,
		_w24344_
	);
	LUT2 #(
		.INIT('h8)
	) name13833 (
		\wishbone_bd_ram_mem0_reg[55][3]/P0001 ,
		_w12785_,
		_w24345_
	);
	LUT2 #(
		.INIT('h8)
	) name13834 (
		\wishbone_bd_ram_mem0_reg[24][3]/P0001 ,
		_w13084_,
		_w24346_
	);
	LUT2 #(
		.INIT('h8)
	) name13835 (
		\wishbone_bd_ram_mem0_reg[168][3]/P0001 ,
		_w13208_,
		_w24347_
	);
	LUT2 #(
		.INIT('h8)
	) name13836 (
		\wishbone_bd_ram_mem0_reg[118][3]/P0001 ,
		_w12830_,
		_w24348_
	);
	LUT2 #(
		.INIT('h8)
	) name13837 (
		\wishbone_bd_ram_mem0_reg[214][3]/P0001 ,
		_w12984_,
		_w24349_
	);
	LUT2 #(
		.INIT('h8)
	) name13838 (
		\wishbone_bd_ram_mem0_reg[213][3]/P0001 ,
		_w13002_,
		_w24350_
	);
	LUT2 #(
		.INIT('h8)
	) name13839 (
		\wishbone_bd_ram_mem0_reg[51][3]/P0001 ,
		_w13024_,
		_w24351_
	);
	LUT2 #(
		.INIT('h8)
	) name13840 (
		\wishbone_bd_ram_mem0_reg[220][3]/P0001 ,
		_w13066_,
		_w24352_
	);
	LUT2 #(
		.INIT('h8)
	) name13841 (
		\wishbone_bd_ram_mem0_reg[70][3]/P0001 ,
		_w12840_,
		_w24353_
	);
	LUT2 #(
		.INIT('h8)
	) name13842 (
		\wishbone_bd_ram_mem0_reg[58][3]/P0001 ,
		_w13070_,
		_w24354_
	);
	LUT2 #(
		.INIT('h8)
	) name13843 (
		\wishbone_bd_ram_mem0_reg[136][3]/P0001 ,
		_w13064_,
		_w24355_
	);
	LUT2 #(
		.INIT('h8)
	) name13844 (
		\wishbone_bd_ram_mem0_reg[224][3]/P0001 ,
		_w12902_,
		_w24356_
	);
	LUT2 #(
		.INIT('h8)
	) name13845 (
		\wishbone_bd_ram_mem0_reg[143][3]/P0001 ,
		_w12922_,
		_w24357_
	);
	LUT2 #(
		.INIT('h8)
	) name13846 (
		\wishbone_bd_ram_mem0_reg[63][3]/P0001 ,
		_w12850_,
		_w24358_
	);
	LUT2 #(
		.INIT('h8)
	) name13847 (
		\wishbone_bd_ram_mem0_reg[77][3]/P0001 ,
		_w12982_,
		_w24359_
	);
	LUT2 #(
		.INIT('h8)
	) name13848 (
		\wishbone_bd_ram_mem0_reg[230][3]/P0001 ,
		_w13036_,
		_w24360_
	);
	LUT2 #(
		.INIT('h8)
	) name13849 (
		\wishbone_bd_ram_mem0_reg[217][3]/P0001 ,
		_w13188_,
		_w24361_
	);
	LUT2 #(
		.INIT('h8)
	) name13850 (
		\wishbone_bd_ram_mem0_reg[154][3]/P0001 ,
		_w12962_,
		_w24362_
	);
	LUT2 #(
		.INIT('h8)
	) name13851 (
		\wishbone_bd_ram_mem0_reg[42][3]/P0001 ,
		_w12842_,
		_w24363_
	);
	LUT2 #(
		.INIT('h8)
	) name13852 (
		\wishbone_bd_ram_mem0_reg[183][3]/P0001 ,
		_w12787_,
		_w24364_
	);
	LUT2 #(
		.INIT('h8)
	) name13853 (
		\wishbone_bd_ram_mem0_reg[36][3]/P0001 ,
		_w12800_,
		_w24365_
	);
	LUT2 #(
		.INIT('h8)
	) name13854 (
		\wishbone_bd_ram_mem0_reg[245][3]/P0001 ,
		_w13022_,
		_w24366_
	);
	LUT2 #(
		.INIT('h8)
	) name13855 (
		\wishbone_bd_ram_mem0_reg[56][3]/P0001 ,
		_w12778_,
		_w24367_
	);
	LUT2 #(
		.INIT('h8)
	) name13856 (
		\wishbone_bd_ram_mem0_reg[193][3]/P0001 ,
		_w13056_,
		_w24368_
	);
	LUT2 #(
		.INIT('h8)
	) name13857 (
		\wishbone_bd_ram_mem0_reg[145][3]/P0001 ,
		_w13106_,
		_w24369_
	);
	LUT2 #(
		.INIT('h8)
	) name13858 (
		\wishbone_bd_ram_mem0_reg[110][3]/P0001 ,
		_w13046_,
		_w24370_
	);
	LUT2 #(
		.INIT('h8)
	) name13859 (
		\wishbone_bd_ram_mem0_reg[116][3]/P0001 ,
		_w12998_,
		_w24371_
	);
	LUT2 #(
		.INIT('h8)
	) name13860 (
		\wishbone_bd_ram_mem0_reg[204][3]/P0001 ,
		_w13162_,
		_w24372_
	);
	LUT2 #(
		.INIT('h8)
	) name13861 (
		\wishbone_bd_ram_mem0_reg[178][3]/P0001 ,
		_w12886_,
		_w24373_
	);
	LUT2 #(
		.INIT('h8)
	) name13862 (
		\wishbone_bd_ram_mem0_reg[170][3]/P0001 ,
		_w13030_,
		_w24374_
	);
	LUT2 #(
		.INIT('h8)
	) name13863 (
		\wishbone_bd_ram_mem0_reg[191][3]/P0001 ,
		_w13034_,
		_w24375_
	);
	LUT2 #(
		.INIT('h8)
	) name13864 (
		\wishbone_bd_ram_mem0_reg[91][3]/P0001 ,
		_w13074_,
		_w24376_
	);
	LUT2 #(
		.INIT('h8)
	) name13865 (
		\wishbone_bd_ram_mem0_reg[127][3]/P0001 ,
		_w13164_,
		_w24377_
	);
	LUT2 #(
		.INIT('h8)
	) name13866 (
		\wishbone_bd_ram_mem0_reg[107][3]/P0001 ,
		_w12749_,
		_w24378_
	);
	LUT2 #(
		.INIT('h8)
	) name13867 (
		\wishbone_bd_ram_mem0_reg[233][3]/P0001 ,
		_w12836_,
		_w24379_
	);
	LUT2 #(
		.INIT('h8)
	) name13868 (
		\wishbone_bd_ram_mem0_reg[0][3]/P0001 ,
		_w12717_,
		_w24380_
	);
	LUT2 #(
		.INIT('h8)
	) name13869 (
		\wishbone_bd_ram_mem0_reg[1][3]/P0001 ,
		_w13014_,
		_w24381_
	);
	LUT2 #(
		.INIT('h8)
	) name13870 (
		\wishbone_bd_ram_mem0_reg[66][3]/P0001 ,
		_w12824_,
		_w24382_
	);
	LUT2 #(
		.INIT('h8)
	) name13871 (
		\wishbone_bd_ram_mem0_reg[52][3]/P0001 ,
		_w13082_,
		_w24383_
	);
	LUT2 #(
		.INIT('h8)
	) name13872 (
		\wishbone_bd_ram_mem0_reg[232][3]/P0001 ,
		_w12758_,
		_w24384_
	);
	LUT2 #(
		.INIT('h8)
	) name13873 (
		\wishbone_bd_ram_mem0_reg[201][3]/P0001 ,
		_w12822_,
		_w24385_
	);
	LUT2 #(
		.INIT('h8)
	) name13874 (
		\wishbone_bd_ram_mem0_reg[195][3]/P0001 ,
		_w13144_,
		_w24386_
	);
	LUT2 #(
		.INIT('h8)
	) name13875 (
		\wishbone_bd_ram_mem0_reg[188][3]/P0001 ,
		_w12948_,
		_w24387_
	);
	LUT2 #(
		.INIT('h8)
	) name13876 (
		\wishbone_bd_ram_mem0_reg[165][3]/P0001 ,
		_w13044_,
		_w24388_
	);
	LUT2 #(
		.INIT('h8)
	) name13877 (
		\wishbone_bd_ram_mem0_reg[227][3]/P0001 ,
		_w12936_,
		_w24389_
	);
	LUT2 #(
		.INIT('h8)
	) name13878 (
		\wishbone_bd_ram_mem0_reg[33][3]/P0001 ,
		_w12980_,
		_w24390_
	);
	LUT2 #(
		.INIT('h8)
	) name13879 (
		\wishbone_bd_ram_mem0_reg[13][3]/P0001 ,
		_w13178_,
		_w24391_
	);
	LUT2 #(
		.INIT('h8)
	) name13880 (
		\wishbone_bd_ram_mem0_reg[177][3]/P0001 ,
		_w12996_,
		_w24392_
	);
	LUT2 #(
		.INIT('h8)
	) name13881 (
		\wishbone_bd_ram_mem0_reg[10][3]/P0001 ,
		_w13172_,
		_w24393_
	);
	LUT2 #(
		.INIT('h8)
	) name13882 (
		\wishbone_bd_ram_mem0_reg[23][3]/P0001 ,
		_w13008_,
		_w24394_
	);
	LUT2 #(
		.INIT('h8)
	) name13883 (
		\wishbone_bd_ram_mem0_reg[22][3]/P0001 ,
		_w13110_,
		_w24395_
	);
	LUT2 #(
		.INIT('h8)
	) name13884 (
		\wishbone_bd_ram_mem0_reg[134][3]/P0001 ,
		_w12763_,
		_w24396_
	);
	LUT2 #(
		.INIT('h8)
	) name13885 (
		\wishbone_bd_ram_mem0_reg[60][3]/P0001 ,
		_w13204_,
		_w24397_
	);
	LUT2 #(
		.INIT('h8)
	) name13886 (
		\wishbone_bd_ram_mem0_reg[18][3]/P0001 ,
		_w12679_,
		_w24398_
	);
	LUT2 #(
		.INIT('h8)
	) name13887 (
		\wishbone_bd_ram_mem0_reg[25][3]/P0001 ,
		_w13108_,
		_w24399_
	);
	LUT2 #(
		.INIT('h8)
	) name13888 (
		\wishbone_bd_ram_mem0_reg[124][3]/P0001 ,
		_w13058_,
		_w24400_
	);
	LUT2 #(
		.INIT('h8)
	) name13889 (
		\wishbone_bd_ram_mem0_reg[29][3]/P0001 ,
		_w12952_,
		_w24401_
	);
	LUT2 #(
		.INIT('h8)
	) name13890 (
		\wishbone_bd_ram_mem0_reg[72][3]/P0001 ,
		_w12810_,
		_w24402_
	);
	LUT2 #(
		.INIT('h8)
	) name13891 (
		\wishbone_bd_ram_mem0_reg[250][3]/P0001 ,
		_w13128_,
		_w24403_
	);
	LUT2 #(
		.INIT('h8)
	) name13892 (
		\wishbone_bd_ram_mem0_reg[71][3]/P0001 ,
		_w12798_,
		_w24404_
	);
	LUT2 #(
		.INIT('h8)
	) name13893 (
		\wishbone_bd_ram_mem0_reg[2][3]/P0001 ,
		_w13088_,
		_w24405_
	);
	LUT2 #(
		.INIT('h8)
	) name13894 (
		\wishbone_bd_ram_mem0_reg[69][3]/P0001 ,
		_w12738_,
		_w24406_
	);
	LUT2 #(
		.INIT('h8)
	) name13895 (
		\wishbone_bd_ram_mem0_reg[152][3]/P0001 ,
		_w12966_,
		_w24407_
	);
	LUT2 #(
		.INIT('h8)
	) name13896 (
		\wishbone_bd_ram_mem0_reg[253][3]/P0001 ,
		_w13100_,
		_w24408_
	);
	LUT2 #(
		.INIT('h8)
	) name13897 (
		\wishbone_bd_ram_mem0_reg[161][3]/P0001 ,
		_w12754_,
		_w24409_
	);
	LUT2 #(
		.INIT('h8)
	) name13898 (
		\wishbone_bd_ram_mem0_reg[95][3]/P0001 ,
		_w12844_,
		_w24410_
	);
	LUT2 #(
		.INIT('h8)
	) name13899 (
		\wishbone_bd_ram_mem0_reg[132][3]/P0001 ,
		_w12992_,
		_w24411_
	);
	LUT2 #(
		.INIT('h8)
	) name13900 (
		\wishbone_bd_ram_mem0_reg[41][3]/P0001 ,
		_w13052_,
		_w24412_
	);
	LUT2 #(
		.INIT('h8)
	) name13901 (
		\wishbone_bd_ram_mem0_reg[84][3]/P0001 ,
		_w12934_,
		_w24413_
	);
	LUT2 #(
		.INIT('h8)
	) name13902 (
		\wishbone_bd_ram_mem0_reg[50][3]/P0001 ,
		_w13150_,
		_w24414_
	);
	LUT2 #(
		.INIT('h8)
	) name13903 (
		\wishbone_bd_ram_mem0_reg[68][3]/P0001 ,
		_w12946_,
		_w24415_
	);
	LUT2 #(
		.INIT('h8)
	) name13904 (
		\wishbone_bd_ram_mem0_reg[219][3]/P0001 ,
		_w12806_,
		_w24416_
	);
	LUT2 #(
		.INIT('h8)
	) name13905 (
		\wishbone_bd_ram_mem0_reg[192][3]/P0001 ,
		_w12938_,
		_w24417_
	);
	LUT2 #(
		.INIT('h8)
	) name13906 (
		\wishbone_bd_ram_mem0_reg[126][3]/P0001 ,
		_w13218_,
		_w24418_
	);
	LUT2 #(
		.INIT('h8)
	) name13907 (
		\wishbone_bd_ram_mem0_reg[240][3]/P0001 ,
		_w12864_,
		_w24419_
	);
	LUT2 #(
		.INIT('h8)
	) name13908 (
		\wishbone_bd_ram_mem0_reg[113][3]/P0001 ,
		_w13026_,
		_w24420_
	);
	LUT2 #(
		.INIT('h8)
	) name13909 (
		\wishbone_bd_ram_mem0_reg[205][3]/P0001 ,
		_w13068_,
		_w24421_
	);
	LUT2 #(
		.INIT('h8)
	) name13910 (
		\wishbone_bd_ram_mem0_reg[255][3]/P0001 ,
		_w13072_,
		_w24422_
	);
	LUT2 #(
		.INIT('h8)
	) name13911 (
		\wishbone_bd_ram_mem0_reg[45][3]/P0001 ,
		_w12908_,
		_w24423_
	);
	LUT2 #(
		.INIT('h8)
	) name13912 (
		\wishbone_bd_ram_mem0_reg[15][3]/P0001 ,
		_w13210_,
		_w24424_
	);
	LUT2 #(
		.INIT('h8)
	) name13913 (
		\wishbone_bd_ram_mem0_reg[35][3]/P0001 ,
		_w12703_,
		_w24425_
	);
	LUT2 #(
		.INIT('h8)
	) name13914 (
		\wishbone_bd_ram_mem0_reg[62][3]/P0001 ,
		_w12673_,
		_w24426_
	);
	LUT2 #(
		.INIT('h8)
	) name13915 (
		\wishbone_bd_ram_mem0_reg[67][3]/P0001 ,
		_w13134_,
		_w24427_
	);
	LUT2 #(
		.INIT('h8)
	) name13916 (
		\wishbone_bd_ram_mem0_reg[16][3]/P0001 ,
		_w13140_,
		_w24428_
	);
	LUT2 #(
		.INIT('h8)
	) name13917 (
		\wishbone_bd_ram_mem0_reg[252][3]/P0001 ,
		_w13080_,
		_w24429_
	);
	LUT2 #(
		.INIT('h8)
	) name13918 (
		\wishbone_bd_ram_mem0_reg[34][3]/P0001 ,
		_w12930_,
		_w24430_
	);
	LUT2 #(
		.INIT('h8)
	) name13919 (
		\wishbone_bd_ram_mem0_reg[73][3]/P0001 ,
		_w12918_,
		_w24431_
	);
	LUT2 #(
		.INIT('h8)
	) name13920 (
		\wishbone_bd_ram_mem0_reg[234][3]/P0001 ,
		_w13214_,
		_w24432_
	);
	LUT2 #(
		.INIT('h8)
	) name13921 (
		\wishbone_bd_ram_mem0_reg[163][3]/P0001 ,
		_w12882_,
		_w24433_
	);
	LUT2 #(
		.INIT('h8)
	) name13922 (
		\wishbone_bd_ram_mem0_reg[103][3]/P0001 ,
		_w12846_,
		_w24434_
	);
	LUT2 #(
		.INIT('h8)
	) name13923 (
		\wishbone_bd_ram_mem0_reg[100][3]/P0001 ,
		_w12960_,
		_w24435_
	);
	LUT2 #(
		.INIT('h8)
	) name13924 (
		\wishbone_bd_ram_mem0_reg[159][3]/P0001 ,
		_w12774_,
		_w24436_
	);
	LUT2 #(
		.INIT('h8)
	) name13925 (
		\wishbone_bd_ram_mem0_reg[254][3]/P0001 ,
		_w12892_,
		_w24437_
	);
	LUT2 #(
		.INIT('h8)
	) name13926 (
		\wishbone_bd_ram_mem0_reg[6][3]/P0001 ,
		_w12968_,
		_w24438_
	);
	LUT2 #(
		.INIT('h8)
	) name13927 (
		\wishbone_bd_ram_mem0_reg[88][3]/P0001 ,
		_w12860_,
		_w24439_
	);
	LUT2 #(
		.INIT('h8)
	) name13928 (
		\wishbone_bd_ram_mem0_reg[203][3]/P0001 ,
		_w13158_,
		_w24440_
	);
	LUT2 #(
		.INIT('h8)
	) name13929 (
		\wishbone_bd_ram_mem0_reg[26][3]/P0001 ,
		_w12699_,
		_w24441_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		\wishbone_bd_ram_mem0_reg[218][3]/P0001 ,
		_w13206_,
		_w24442_
	);
	LUT2 #(
		.INIT('h8)
	) name13931 (
		\wishbone_bd_ram_mem0_reg[82][3]/P0001 ,
		_w12942_,
		_w24443_
	);
	LUT2 #(
		.INIT('h8)
	) name13932 (
		\wishbone_bd_ram_mem0_reg[19][3]/P0001 ,
		_w13012_,
		_w24444_
	);
	LUT2 #(
		.INIT('h8)
	) name13933 (
		\wishbone_bd_ram_mem0_reg[104][3]/P0001 ,
		_w13148_,
		_w24445_
	);
	LUT2 #(
		.INIT('h8)
	) name13934 (
		\wishbone_bd_ram_mem0_reg[176][3]/P0001 ,
		_w12868_,
		_w24446_
	);
	LUT2 #(
		.INIT('h8)
	) name13935 (
		\wishbone_bd_ram_mem0_reg[80][3]/P0001 ,
		_w12689_,
		_w24447_
	);
	LUT2 #(
		.INIT('h8)
	) name13936 (
		\wishbone_bd_ram_mem0_reg[200][3]/P0001 ,
		_w12988_,
		_w24448_
	);
	LUT2 #(
		.INIT('h1)
	) name13937 (
		_w24193_,
		_w24194_,
		_w24449_
	);
	LUT2 #(
		.INIT('h1)
	) name13938 (
		_w24195_,
		_w24196_,
		_w24450_
	);
	LUT2 #(
		.INIT('h1)
	) name13939 (
		_w24197_,
		_w24198_,
		_w24451_
	);
	LUT2 #(
		.INIT('h1)
	) name13940 (
		_w24199_,
		_w24200_,
		_w24452_
	);
	LUT2 #(
		.INIT('h1)
	) name13941 (
		_w24201_,
		_w24202_,
		_w24453_
	);
	LUT2 #(
		.INIT('h1)
	) name13942 (
		_w24203_,
		_w24204_,
		_w24454_
	);
	LUT2 #(
		.INIT('h1)
	) name13943 (
		_w24205_,
		_w24206_,
		_w24455_
	);
	LUT2 #(
		.INIT('h1)
	) name13944 (
		_w24207_,
		_w24208_,
		_w24456_
	);
	LUT2 #(
		.INIT('h1)
	) name13945 (
		_w24209_,
		_w24210_,
		_w24457_
	);
	LUT2 #(
		.INIT('h1)
	) name13946 (
		_w24211_,
		_w24212_,
		_w24458_
	);
	LUT2 #(
		.INIT('h1)
	) name13947 (
		_w24213_,
		_w24214_,
		_w24459_
	);
	LUT2 #(
		.INIT('h1)
	) name13948 (
		_w24215_,
		_w24216_,
		_w24460_
	);
	LUT2 #(
		.INIT('h1)
	) name13949 (
		_w24217_,
		_w24218_,
		_w24461_
	);
	LUT2 #(
		.INIT('h1)
	) name13950 (
		_w24219_,
		_w24220_,
		_w24462_
	);
	LUT2 #(
		.INIT('h1)
	) name13951 (
		_w24221_,
		_w24222_,
		_w24463_
	);
	LUT2 #(
		.INIT('h1)
	) name13952 (
		_w24223_,
		_w24224_,
		_w24464_
	);
	LUT2 #(
		.INIT('h1)
	) name13953 (
		_w24225_,
		_w24226_,
		_w24465_
	);
	LUT2 #(
		.INIT('h1)
	) name13954 (
		_w24227_,
		_w24228_,
		_w24466_
	);
	LUT2 #(
		.INIT('h1)
	) name13955 (
		_w24229_,
		_w24230_,
		_w24467_
	);
	LUT2 #(
		.INIT('h1)
	) name13956 (
		_w24231_,
		_w24232_,
		_w24468_
	);
	LUT2 #(
		.INIT('h1)
	) name13957 (
		_w24233_,
		_w24234_,
		_w24469_
	);
	LUT2 #(
		.INIT('h1)
	) name13958 (
		_w24235_,
		_w24236_,
		_w24470_
	);
	LUT2 #(
		.INIT('h1)
	) name13959 (
		_w24237_,
		_w24238_,
		_w24471_
	);
	LUT2 #(
		.INIT('h1)
	) name13960 (
		_w24239_,
		_w24240_,
		_w24472_
	);
	LUT2 #(
		.INIT('h1)
	) name13961 (
		_w24241_,
		_w24242_,
		_w24473_
	);
	LUT2 #(
		.INIT('h1)
	) name13962 (
		_w24243_,
		_w24244_,
		_w24474_
	);
	LUT2 #(
		.INIT('h1)
	) name13963 (
		_w24245_,
		_w24246_,
		_w24475_
	);
	LUT2 #(
		.INIT('h1)
	) name13964 (
		_w24247_,
		_w24248_,
		_w24476_
	);
	LUT2 #(
		.INIT('h1)
	) name13965 (
		_w24249_,
		_w24250_,
		_w24477_
	);
	LUT2 #(
		.INIT('h1)
	) name13966 (
		_w24251_,
		_w24252_,
		_w24478_
	);
	LUT2 #(
		.INIT('h1)
	) name13967 (
		_w24253_,
		_w24254_,
		_w24479_
	);
	LUT2 #(
		.INIT('h1)
	) name13968 (
		_w24255_,
		_w24256_,
		_w24480_
	);
	LUT2 #(
		.INIT('h1)
	) name13969 (
		_w24257_,
		_w24258_,
		_w24481_
	);
	LUT2 #(
		.INIT('h1)
	) name13970 (
		_w24259_,
		_w24260_,
		_w24482_
	);
	LUT2 #(
		.INIT('h1)
	) name13971 (
		_w24261_,
		_w24262_,
		_w24483_
	);
	LUT2 #(
		.INIT('h1)
	) name13972 (
		_w24263_,
		_w24264_,
		_w24484_
	);
	LUT2 #(
		.INIT('h1)
	) name13973 (
		_w24265_,
		_w24266_,
		_w24485_
	);
	LUT2 #(
		.INIT('h1)
	) name13974 (
		_w24267_,
		_w24268_,
		_w24486_
	);
	LUT2 #(
		.INIT('h1)
	) name13975 (
		_w24269_,
		_w24270_,
		_w24487_
	);
	LUT2 #(
		.INIT('h1)
	) name13976 (
		_w24271_,
		_w24272_,
		_w24488_
	);
	LUT2 #(
		.INIT('h1)
	) name13977 (
		_w24273_,
		_w24274_,
		_w24489_
	);
	LUT2 #(
		.INIT('h1)
	) name13978 (
		_w24275_,
		_w24276_,
		_w24490_
	);
	LUT2 #(
		.INIT('h1)
	) name13979 (
		_w24277_,
		_w24278_,
		_w24491_
	);
	LUT2 #(
		.INIT('h1)
	) name13980 (
		_w24279_,
		_w24280_,
		_w24492_
	);
	LUT2 #(
		.INIT('h1)
	) name13981 (
		_w24281_,
		_w24282_,
		_w24493_
	);
	LUT2 #(
		.INIT('h1)
	) name13982 (
		_w24283_,
		_w24284_,
		_w24494_
	);
	LUT2 #(
		.INIT('h1)
	) name13983 (
		_w24285_,
		_w24286_,
		_w24495_
	);
	LUT2 #(
		.INIT('h1)
	) name13984 (
		_w24287_,
		_w24288_,
		_w24496_
	);
	LUT2 #(
		.INIT('h1)
	) name13985 (
		_w24289_,
		_w24290_,
		_w24497_
	);
	LUT2 #(
		.INIT('h1)
	) name13986 (
		_w24291_,
		_w24292_,
		_w24498_
	);
	LUT2 #(
		.INIT('h1)
	) name13987 (
		_w24293_,
		_w24294_,
		_w24499_
	);
	LUT2 #(
		.INIT('h1)
	) name13988 (
		_w24295_,
		_w24296_,
		_w24500_
	);
	LUT2 #(
		.INIT('h1)
	) name13989 (
		_w24297_,
		_w24298_,
		_w24501_
	);
	LUT2 #(
		.INIT('h1)
	) name13990 (
		_w24299_,
		_w24300_,
		_w24502_
	);
	LUT2 #(
		.INIT('h1)
	) name13991 (
		_w24301_,
		_w24302_,
		_w24503_
	);
	LUT2 #(
		.INIT('h1)
	) name13992 (
		_w24303_,
		_w24304_,
		_w24504_
	);
	LUT2 #(
		.INIT('h1)
	) name13993 (
		_w24305_,
		_w24306_,
		_w24505_
	);
	LUT2 #(
		.INIT('h1)
	) name13994 (
		_w24307_,
		_w24308_,
		_w24506_
	);
	LUT2 #(
		.INIT('h1)
	) name13995 (
		_w24309_,
		_w24310_,
		_w24507_
	);
	LUT2 #(
		.INIT('h1)
	) name13996 (
		_w24311_,
		_w24312_,
		_w24508_
	);
	LUT2 #(
		.INIT('h1)
	) name13997 (
		_w24313_,
		_w24314_,
		_w24509_
	);
	LUT2 #(
		.INIT('h1)
	) name13998 (
		_w24315_,
		_w24316_,
		_w24510_
	);
	LUT2 #(
		.INIT('h1)
	) name13999 (
		_w24317_,
		_w24318_,
		_w24511_
	);
	LUT2 #(
		.INIT('h1)
	) name14000 (
		_w24319_,
		_w24320_,
		_w24512_
	);
	LUT2 #(
		.INIT('h1)
	) name14001 (
		_w24321_,
		_w24322_,
		_w24513_
	);
	LUT2 #(
		.INIT('h1)
	) name14002 (
		_w24323_,
		_w24324_,
		_w24514_
	);
	LUT2 #(
		.INIT('h1)
	) name14003 (
		_w24325_,
		_w24326_,
		_w24515_
	);
	LUT2 #(
		.INIT('h1)
	) name14004 (
		_w24327_,
		_w24328_,
		_w24516_
	);
	LUT2 #(
		.INIT('h1)
	) name14005 (
		_w24329_,
		_w24330_,
		_w24517_
	);
	LUT2 #(
		.INIT('h1)
	) name14006 (
		_w24331_,
		_w24332_,
		_w24518_
	);
	LUT2 #(
		.INIT('h1)
	) name14007 (
		_w24333_,
		_w24334_,
		_w24519_
	);
	LUT2 #(
		.INIT('h1)
	) name14008 (
		_w24335_,
		_w24336_,
		_w24520_
	);
	LUT2 #(
		.INIT('h1)
	) name14009 (
		_w24337_,
		_w24338_,
		_w24521_
	);
	LUT2 #(
		.INIT('h1)
	) name14010 (
		_w24339_,
		_w24340_,
		_w24522_
	);
	LUT2 #(
		.INIT('h1)
	) name14011 (
		_w24341_,
		_w24342_,
		_w24523_
	);
	LUT2 #(
		.INIT('h1)
	) name14012 (
		_w24343_,
		_w24344_,
		_w24524_
	);
	LUT2 #(
		.INIT('h1)
	) name14013 (
		_w24345_,
		_w24346_,
		_w24525_
	);
	LUT2 #(
		.INIT('h1)
	) name14014 (
		_w24347_,
		_w24348_,
		_w24526_
	);
	LUT2 #(
		.INIT('h1)
	) name14015 (
		_w24349_,
		_w24350_,
		_w24527_
	);
	LUT2 #(
		.INIT('h1)
	) name14016 (
		_w24351_,
		_w24352_,
		_w24528_
	);
	LUT2 #(
		.INIT('h1)
	) name14017 (
		_w24353_,
		_w24354_,
		_w24529_
	);
	LUT2 #(
		.INIT('h1)
	) name14018 (
		_w24355_,
		_w24356_,
		_w24530_
	);
	LUT2 #(
		.INIT('h1)
	) name14019 (
		_w24357_,
		_w24358_,
		_w24531_
	);
	LUT2 #(
		.INIT('h1)
	) name14020 (
		_w24359_,
		_w24360_,
		_w24532_
	);
	LUT2 #(
		.INIT('h1)
	) name14021 (
		_w24361_,
		_w24362_,
		_w24533_
	);
	LUT2 #(
		.INIT('h1)
	) name14022 (
		_w24363_,
		_w24364_,
		_w24534_
	);
	LUT2 #(
		.INIT('h1)
	) name14023 (
		_w24365_,
		_w24366_,
		_w24535_
	);
	LUT2 #(
		.INIT('h1)
	) name14024 (
		_w24367_,
		_w24368_,
		_w24536_
	);
	LUT2 #(
		.INIT('h1)
	) name14025 (
		_w24369_,
		_w24370_,
		_w24537_
	);
	LUT2 #(
		.INIT('h1)
	) name14026 (
		_w24371_,
		_w24372_,
		_w24538_
	);
	LUT2 #(
		.INIT('h1)
	) name14027 (
		_w24373_,
		_w24374_,
		_w24539_
	);
	LUT2 #(
		.INIT('h1)
	) name14028 (
		_w24375_,
		_w24376_,
		_w24540_
	);
	LUT2 #(
		.INIT('h1)
	) name14029 (
		_w24377_,
		_w24378_,
		_w24541_
	);
	LUT2 #(
		.INIT('h1)
	) name14030 (
		_w24379_,
		_w24380_,
		_w24542_
	);
	LUT2 #(
		.INIT('h1)
	) name14031 (
		_w24381_,
		_w24382_,
		_w24543_
	);
	LUT2 #(
		.INIT('h1)
	) name14032 (
		_w24383_,
		_w24384_,
		_w24544_
	);
	LUT2 #(
		.INIT('h1)
	) name14033 (
		_w24385_,
		_w24386_,
		_w24545_
	);
	LUT2 #(
		.INIT('h1)
	) name14034 (
		_w24387_,
		_w24388_,
		_w24546_
	);
	LUT2 #(
		.INIT('h1)
	) name14035 (
		_w24389_,
		_w24390_,
		_w24547_
	);
	LUT2 #(
		.INIT('h1)
	) name14036 (
		_w24391_,
		_w24392_,
		_w24548_
	);
	LUT2 #(
		.INIT('h1)
	) name14037 (
		_w24393_,
		_w24394_,
		_w24549_
	);
	LUT2 #(
		.INIT('h1)
	) name14038 (
		_w24395_,
		_w24396_,
		_w24550_
	);
	LUT2 #(
		.INIT('h1)
	) name14039 (
		_w24397_,
		_w24398_,
		_w24551_
	);
	LUT2 #(
		.INIT('h1)
	) name14040 (
		_w24399_,
		_w24400_,
		_w24552_
	);
	LUT2 #(
		.INIT('h1)
	) name14041 (
		_w24401_,
		_w24402_,
		_w24553_
	);
	LUT2 #(
		.INIT('h1)
	) name14042 (
		_w24403_,
		_w24404_,
		_w24554_
	);
	LUT2 #(
		.INIT('h1)
	) name14043 (
		_w24405_,
		_w24406_,
		_w24555_
	);
	LUT2 #(
		.INIT('h1)
	) name14044 (
		_w24407_,
		_w24408_,
		_w24556_
	);
	LUT2 #(
		.INIT('h1)
	) name14045 (
		_w24409_,
		_w24410_,
		_w24557_
	);
	LUT2 #(
		.INIT('h1)
	) name14046 (
		_w24411_,
		_w24412_,
		_w24558_
	);
	LUT2 #(
		.INIT('h1)
	) name14047 (
		_w24413_,
		_w24414_,
		_w24559_
	);
	LUT2 #(
		.INIT('h1)
	) name14048 (
		_w24415_,
		_w24416_,
		_w24560_
	);
	LUT2 #(
		.INIT('h1)
	) name14049 (
		_w24417_,
		_w24418_,
		_w24561_
	);
	LUT2 #(
		.INIT('h1)
	) name14050 (
		_w24419_,
		_w24420_,
		_w24562_
	);
	LUT2 #(
		.INIT('h1)
	) name14051 (
		_w24421_,
		_w24422_,
		_w24563_
	);
	LUT2 #(
		.INIT('h1)
	) name14052 (
		_w24423_,
		_w24424_,
		_w24564_
	);
	LUT2 #(
		.INIT('h1)
	) name14053 (
		_w24425_,
		_w24426_,
		_w24565_
	);
	LUT2 #(
		.INIT('h1)
	) name14054 (
		_w24427_,
		_w24428_,
		_w24566_
	);
	LUT2 #(
		.INIT('h1)
	) name14055 (
		_w24429_,
		_w24430_,
		_w24567_
	);
	LUT2 #(
		.INIT('h1)
	) name14056 (
		_w24431_,
		_w24432_,
		_w24568_
	);
	LUT2 #(
		.INIT('h1)
	) name14057 (
		_w24433_,
		_w24434_,
		_w24569_
	);
	LUT2 #(
		.INIT('h1)
	) name14058 (
		_w24435_,
		_w24436_,
		_w24570_
	);
	LUT2 #(
		.INIT('h1)
	) name14059 (
		_w24437_,
		_w24438_,
		_w24571_
	);
	LUT2 #(
		.INIT('h1)
	) name14060 (
		_w24439_,
		_w24440_,
		_w24572_
	);
	LUT2 #(
		.INIT('h1)
	) name14061 (
		_w24441_,
		_w24442_,
		_w24573_
	);
	LUT2 #(
		.INIT('h1)
	) name14062 (
		_w24443_,
		_w24444_,
		_w24574_
	);
	LUT2 #(
		.INIT('h1)
	) name14063 (
		_w24445_,
		_w24446_,
		_w24575_
	);
	LUT2 #(
		.INIT('h1)
	) name14064 (
		_w24447_,
		_w24448_,
		_w24576_
	);
	LUT2 #(
		.INIT('h8)
	) name14065 (
		_w24575_,
		_w24576_,
		_w24577_
	);
	LUT2 #(
		.INIT('h8)
	) name14066 (
		_w24573_,
		_w24574_,
		_w24578_
	);
	LUT2 #(
		.INIT('h8)
	) name14067 (
		_w24571_,
		_w24572_,
		_w24579_
	);
	LUT2 #(
		.INIT('h8)
	) name14068 (
		_w24569_,
		_w24570_,
		_w24580_
	);
	LUT2 #(
		.INIT('h8)
	) name14069 (
		_w24567_,
		_w24568_,
		_w24581_
	);
	LUT2 #(
		.INIT('h8)
	) name14070 (
		_w24565_,
		_w24566_,
		_w24582_
	);
	LUT2 #(
		.INIT('h8)
	) name14071 (
		_w24563_,
		_w24564_,
		_w24583_
	);
	LUT2 #(
		.INIT('h8)
	) name14072 (
		_w24561_,
		_w24562_,
		_w24584_
	);
	LUT2 #(
		.INIT('h8)
	) name14073 (
		_w24559_,
		_w24560_,
		_w24585_
	);
	LUT2 #(
		.INIT('h8)
	) name14074 (
		_w24557_,
		_w24558_,
		_w24586_
	);
	LUT2 #(
		.INIT('h8)
	) name14075 (
		_w24555_,
		_w24556_,
		_w24587_
	);
	LUT2 #(
		.INIT('h8)
	) name14076 (
		_w24553_,
		_w24554_,
		_w24588_
	);
	LUT2 #(
		.INIT('h8)
	) name14077 (
		_w24551_,
		_w24552_,
		_w24589_
	);
	LUT2 #(
		.INIT('h8)
	) name14078 (
		_w24549_,
		_w24550_,
		_w24590_
	);
	LUT2 #(
		.INIT('h8)
	) name14079 (
		_w24547_,
		_w24548_,
		_w24591_
	);
	LUT2 #(
		.INIT('h8)
	) name14080 (
		_w24545_,
		_w24546_,
		_w24592_
	);
	LUT2 #(
		.INIT('h8)
	) name14081 (
		_w24543_,
		_w24544_,
		_w24593_
	);
	LUT2 #(
		.INIT('h8)
	) name14082 (
		_w24541_,
		_w24542_,
		_w24594_
	);
	LUT2 #(
		.INIT('h8)
	) name14083 (
		_w24539_,
		_w24540_,
		_w24595_
	);
	LUT2 #(
		.INIT('h8)
	) name14084 (
		_w24537_,
		_w24538_,
		_w24596_
	);
	LUT2 #(
		.INIT('h8)
	) name14085 (
		_w24535_,
		_w24536_,
		_w24597_
	);
	LUT2 #(
		.INIT('h8)
	) name14086 (
		_w24533_,
		_w24534_,
		_w24598_
	);
	LUT2 #(
		.INIT('h8)
	) name14087 (
		_w24531_,
		_w24532_,
		_w24599_
	);
	LUT2 #(
		.INIT('h8)
	) name14088 (
		_w24529_,
		_w24530_,
		_w24600_
	);
	LUT2 #(
		.INIT('h8)
	) name14089 (
		_w24527_,
		_w24528_,
		_w24601_
	);
	LUT2 #(
		.INIT('h8)
	) name14090 (
		_w24525_,
		_w24526_,
		_w24602_
	);
	LUT2 #(
		.INIT('h8)
	) name14091 (
		_w24523_,
		_w24524_,
		_w24603_
	);
	LUT2 #(
		.INIT('h8)
	) name14092 (
		_w24521_,
		_w24522_,
		_w24604_
	);
	LUT2 #(
		.INIT('h8)
	) name14093 (
		_w24519_,
		_w24520_,
		_w24605_
	);
	LUT2 #(
		.INIT('h8)
	) name14094 (
		_w24517_,
		_w24518_,
		_w24606_
	);
	LUT2 #(
		.INIT('h8)
	) name14095 (
		_w24515_,
		_w24516_,
		_w24607_
	);
	LUT2 #(
		.INIT('h8)
	) name14096 (
		_w24513_,
		_w24514_,
		_w24608_
	);
	LUT2 #(
		.INIT('h8)
	) name14097 (
		_w24511_,
		_w24512_,
		_w24609_
	);
	LUT2 #(
		.INIT('h8)
	) name14098 (
		_w24509_,
		_w24510_,
		_w24610_
	);
	LUT2 #(
		.INIT('h8)
	) name14099 (
		_w24507_,
		_w24508_,
		_w24611_
	);
	LUT2 #(
		.INIT('h8)
	) name14100 (
		_w24505_,
		_w24506_,
		_w24612_
	);
	LUT2 #(
		.INIT('h8)
	) name14101 (
		_w24503_,
		_w24504_,
		_w24613_
	);
	LUT2 #(
		.INIT('h8)
	) name14102 (
		_w24501_,
		_w24502_,
		_w24614_
	);
	LUT2 #(
		.INIT('h8)
	) name14103 (
		_w24499_,
		_w24500_,
		_w24615_
	);
	LUT2 #(
		.INIT('h8)
	) name14104 (
		_w24497_,
		_w24498_,
		_w24616_
	);
	LUT2 #(
		.INIT('h8)
	) name14105 (
		_w24495_,
		_w24496_,
		_w24617_
	);
	LUT2 #(
		.INIT('h8)
	) name14106 (
		_w24493_,
		_w24494_,
		_w24618_
	);
	LUT2 #(
		.INIT('h8)
	) name14107 (
		_w24491_,
		_w24492_,
		_w24619_
	);
	LUT2 #(
		.INIT('h8)
	) name14108 (
		_w24489_,
		_w24490_,
		_w24620_
	);
	LUT2 #(
		.INIT('h8)
	) name14109 (
		_w24487_,
		_w24488_,
		_w24621_
	);
	LUT2 #(
		.INIT('h8)
	) name14110 (
		_w24485_,
		_w24486_,
		_w24622_
	);
	LUT2 #(
		.INIT('h8)
	) name14111 (
		_w24483_,
		_w24484_,
		_w24623_
	);
	LUT2 #(
		.INIT('h8)
	) name14112 (
		_w24481_,
		_w24482_,
		_w24624_
	);
	LUT2 #(
		.INIT('h8)
	) name14113 (
		_w24479_,
		_w24480_,
		_w24625_
	);
	LUT2 #(
		.INIT('h8)
	) name14114 (
		_w24477_,
		_w24478_,
		_w24626_
	);
	LUT2 #(
		.INIT('h8)
	) name14115 (
		_w24475_,
		_w24476_,
		_w24627_
	);
	LUT2 #(
		.INIT('h8)
	) name14116 (
		_w24473_,
		_w24474_,
		_w24628_
	);
	LUT2 #(
		.INIT('h8)
	) name14117 (
		_w24471_,
		_w24472_,
		_w24629_
	);
	LUT2 #(
		.INIT('h8)
	) name14118 (
		_w24469_,
		_w24470_,
		_w24630_
	);
	LUT2 #(
		.INIT('h8)
	) name14119 (
		_w24467_,
		_w24468_,
		_w24631_
	);
	LUT2 #(
		.INIT('h8)
	) name14120 (
		_w24465_,
		_w24466_,
		_w24632_
	);
	LUT2 #(
		.INIT('h8)
	) name14121 (
		_w24463_,
		_w24464_,
		_w24633_
	);
	LUT2 #(
		.INIT('h8)
	) name14122 (
		_w24461_,
		_w24462_,
		_w24634_
	);
	LUT2 #(
		.INIT('h8)
	) name14123 (
		_w24459_,
		_w24460_,
		_w24635_
	);
	LUT2 #(
		.INIT('h8)
	) name14124 (
		_w24457_,
		_w24458_,
		_w24636_
	);
	LUT2 #(
		.INIT('h8)
	) name14125 (
		_w24455_,
		_w24456_,
		_w24637_
	);
	LUT2 #(
		.INIT('h8)
	) name14126 (
		_w24453_,
		_w24454_,
		_w24638_
	);
	LUT2 #(
		.INIT('h8)
	) name14127 (
		_w24451_,
		_w24452_,
		_w24639_
	);
	LUT2 #(
		.INIT('h8)
	) name14128 (
		_w24449_,
		_w24450_,
		_w24640_
	);
	LUT2 #(
		.INIT('h8)
	) name14129 (
		_w24639_,
		_w24640_,
		_w24641_
	);
	LUT2 #(
		.INIT('h8)
	) name14130 (
		_w24637_,
		_w24638_,
		_w24642_
	);
	LUT2 #(
		.INIT('h8)
	) name14131 (
		_w24635_,
		_w24636_,
		_w24643_
	);
	LUT2 #(
		.INIT('h8)
	) name14132 (
		_w24633_,
		_w24634_,
		_w24644_
	);
	LUT2 #(
		.INIT('h8)
	) name14133 (
		_w24631_,
		_w24632_,
		_w24645_
	);
	LUT2 #(
		.INIT('h8)
	) name14134 (
		_w24629_,
		_w24630_,
		_w24646_
	);
	LUT2 #(
		.INIT('h8)
	) name14135 (
		_w24627_,
		_w24628_,
		_w24647_
	);
	LUT2 #(
		.INIT('h8)
	) name14136 (
		_w24625_,
		_w24626_,
		_w24648_
	);
	LUT2 #(
		.INIT('h8)
	) name14137 (
		_w24623_,
		_w24624_,
		_w24649_
	);
	LUT2 #(
		.INIT('h8)
	) name14138 (
		_w24621_,
		_w24622_,
		_w24650_
	);
	LUT2 #(
		.INIT('h8)
	) name14139 (
		_w24619_,
		_w24620_,
		_w24651_
	);
	LUT2 #(
		.INIT('h8)
	) name14140 (
		_w24617_,
		_w24618_,
		_w24652_
	);
	LUT2 #(
		.INIT('h8)
	) name14141 (
		_w24615_,
		_w24616_,
		_w24653_
	);
	LUT2 #(
		.INIT('h8)
	) name14142 (
		_w24613_,
		_w24614_,
		_w24654_
	);
	LUT2 #(
		.INIT('h8)
	) name14143 (
		_w24611_,
		_w24612_,
		_w24655_
	);
	LUT2 #(
		.INIT('h8)
	) name14144 (
		_w24609_,
		_w24610_,
		_w24656_
	);
	LUT2 #(
		.INIT('h8)
	) name14145 (
		_w24607_,
		_w24608_,
		_w24657_
	);
	LUT2 #(
		.INIT('h8)
	) name14146 (
		_w24605_,
		_w24606_,
		_w24658_
	);
	LUT2 #(
		.INIT('h8)
	) name14147 (
		_w24603_,
		_w24604_,
		_w24659_
	);
	LUT2 #(
		.INIT('h8)
	) name14148 (
		_w24601_,
		_w24602_,
		_w24660_
	);
	LUT2 #(
		.INIT('h8)
	) name14149 (
		_w24599_,
		_w24600_,
		_w24661_
	);
	LUT2 #(
		.INIT('h8)
	) name14150 (
		_w24597_,
		_w24598_,
		_w24662_
	);
	LUT2 #(
		.INIT('h8)
	) name14151 (
		_w24595_,
		_w24596_,
		_w24663_
	);
	LUT2 #(
		.INIT('h8)
	) name14152 (
		_w24593_,
		_w24594_,
		_w24664_
	);
	LUT2 #(
		.INIT('h8)
	) name14153 (
		_w24591_,
		_w24592_,
		_w24665_
	);
	LUT2 #(
		.INIT('h8)
	) name14154 (
		_w24589_,
		_w24590_,
		_w24666_
	);
	LUT2 #(
		.INIT('h8)
	) name14155 (
		_w24587_,
		_w24588_,
		_w24667_
	);
	LUT2 #(
		.INIT('h8)
	) name14156 (
		_w24585_,
		_w24586_,
		_w24668_
	);
	LUT2 #(
		.INIT('h8)
	) name14157 (
		_w24583_,
		_w24584_,
		_w24669_
	);
	LUT2 #(
		.INIT('h8)
	) name14158 (
		_w24581_,
		_w24582_,
		_w24670_
	);
	LUT2 #(
		.INIT('h8)
	) name14159 (
		_w24579_,
		_w24580_,
		_w24671_
	);
	LUT2 #(
		.INIT('h8)
	) name14160 (
		_w24577_,
		_w24578_,
		_w24672_
	);
	LUT2 #(
		.INIT('h8)
	) name14161 (
		_w24671_,
		_w24672_,
		_w24673_
	);
	LUT2 #(
		.INIT('h8)
	) name14162 (
		_w24669_,
		_w24670_,
		_w24674_
	);
	LUT2 #(
		.INIT('h8)
	) name14163 (
		_w24667_,
		_w24668_,
		_w24675_
	);
	LUT2 #(
		.INIT('h8)
	) name14164 (
		_w24665_,
		_w24666_,
		_w24676_
	);
	LUT2 #(
		.INIT('h8)
	) name14165 (
		_w24663_,
		_w24664_,
		_w24677_
	);
	LUT2 #(
		.INIT('h8)
	) name14166 (
		_w24661_,
		_w24662_,
		_w24678_
	);
	LUT2 #(
		.INIT('h8)
	) name14167 (
		_w24659_,
		_w24660_,
		_w24679_
	);
	LUT2 #(
		.INIT('h8)
	) name14168 (
		_w24657_,
		_w24658_,
		_w24680_
	);
	LUT2 #(
		.INIT('h8)
	) name14169 (
		_w24655_,
		_w24656_,
		_w24681_
	);
	LUT2 #(
		.INIT('h8)
	) name14170 (
		_w24653_,
		_w24654_,
		_w24682_
	);
	LUT2 #(
		.INIT('h8)
	) name14171 (
		_w24651_,
		_w24652_,
		_w24683_
	);
	LUT2 #(
		.INIT('h8)
	) name14172 (
		_w24649_,
		_w24650_,
		_w24684_
	);
	LUT2 #(
		.INIT('h8)
	) name14173 (
		_w24647_,
		_w24648_,
		_w24685_
	);
	LUT2 #(
		.INIT('h8)
	) name14174 (
		_w24645_,
		_w24646_,
		_w24686_
	);
	LUT2 #(
		.INIT('h8)
	) name14175 (
		_w24643_,
		_w24644_,
		_w24687_
	);
	LUT2 #(
		.INIT('h8)
	) name14176 (
		_w24641_,
		_w24642_,
		_w24688_
	);
	LUT2 #(
		.INIT('h8)
	) name14177 (
		_w24687_,
		_w24688_,
		_w24689_
	);
	LUT2 #(
		.INIT('h8)
	) name14178 (
		_w24685_,
		_w24686_,
		_w24690_
	);
	LUT2 #(
		.INIT('h8)
	) name14179 (
		_w24683_,
		_w24684_,
		_w24691_
	);
	LUT2 #(
		.INIT('h8)
	) name14180 (
		_w24681_,
		_w24682_,
		_w24692_
	);
	LUT2 #(
		.INIT('h8)
	) name14181 (
		_w24679_,
		_w24680_,
		_w24693_
	);
	LUT2 #(
		.INIT('h8)
	) name14182 (
		_w24677_,
		_w24678_,
		_w24694_
	);
	LUT2 #(
		.INIT('h8)
	) name14183 (
		_w24675_,
		_w24676_,
		_w24695_
	);
	LUT2 #(
		.INIT('h8)
	) name14184 (
		_w24673_,
		_w24674_,
		_w24696_
	);
	LUT2 #(
		.INIT('h8)
	) name14185 (
		_w24695_,
		_w24696_,
		_w24697_
	);
	LUT2 #(
		.INIT('h8)
	) name14186 (
		_w24693_,
		_w24694_,
		_w24698_
	);
	LUT2 #(
		.INIT('h8)
	) name14187 (
		_w24691_,
		_w24692_,
		_w24699_
	);
	LUT2 #(
		.INIT('h8)
	) name14188 (
		_w24689_,
		_w24690_,
		_w24700_
	);
	LUT2 #(
		.INIT('h8)
	) name14189 (
		_w24699_,
		_w24700_,
		_w24701_
	);
	LUT2 #(
		.INIT('h8)
	) name14190 (
		_w24697_,
		_w24698_,
		_w24702_
	);
	LUT2 #(
		.INIT('h8)
	) name14191 (
		_w24701_,
		_w24702_,
		_w24703_
	);
	LUT2 #(
		.INIT('h1)
	) name14192 (
		wb_rst_i_pad,
		_w24703_,
		_w24704_
	);
	LUT2 #(
		.INIT('h1)
	) name14193 (
		_w22944_,
		_w24704_,
		_w24705_
	);
	LUT2 #(
		.INIT('h8)
	) name14194 (
		_w22954_,
		_w23517_,
		_w24706_
	);
	LUT2 #(
		.INIT('h8)
	) name14195 (
		_w23516_,
		_w24706_,
		_w24707_
	);
	LUT2 #(
		.INIT('h8)
	) name14196 (
		\ethreg1_irq_rxe_reg/NET0131 ,
		_w24707_,
		_w24708_
	);
	LUT2 #(
		.INIT('h8)
	) name14197 (
		\ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 ,
		_w23499_,
		_w24709_
	);
	LUT2 #(
		.INIT('h8)
	) name14198 (
		_w23504_,
		_w23516_,
		_w24710_
	);
	LUT2 #(
		.INIT('h8)
	) name14199 (
		\ethreg1_IPGR1_0_DataOut_reg[3]/NET0131 ,
		_w24710_,
		_w24711_
	);
	LUT2 #(
		.INIT('h8)
	) name14200 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 ,
		_w23513_,
		_w24712_
	);
	LUT2 #(
		.INIT('h8)
	) name14201 (
		_w23512_,
		_w23518_,
		_w24713_
	);
	LUT2 #(
		.INIT('h8)
	) name14202 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w24713_,
		_w24714_
	);
	LUT2 #(
		.INIT('h8)
	) name14203 (
		\ethreg1_PACKETLEN_0_DataOut_reg[3]/NET0131 ,
		_w22966_,
		_w24715_
	);
	LUT2 #(
		.INIT('h4)
	) name14204 (
		\wb_adr_i[5]_pad ,
		_w23505_,
		_w24716_
	);
	LUT2 #(
		.INIT('h8)
	) name14205 (
		_w24706_,
		_w24716_,
		_w24717_
	);
	LUT2 #(
		.INIT('h8)
	) name14206 (
		\ethreg1_IPGT_0_DataOut_reg[3]/NET0131 ,
		_w24717_,
		_w24718_
	);
	LUT2 #(
		.INIT('h8)
	) name14207 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 ,
		_w23522_,
		_w24719_
	);
	LUT2 #(
		.INIT('h8)
	) name14208 (
		\ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 ,
		_w22952_,
		_w24720_
	);
	LUT2 #(
		.INIT('h8)
	) name14209 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		_w23501_,
		_w24721_
	);
	LUT2 #(
		.INIT('h8)
	) name14210 (
		_w23518_,
		_w24716_,
		_w24722_
	);
	LUT2 #(
		.INIT('h8)
	) name14211 (
		\ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 ,
		_w24722_,
		_w24723_
	);
	LUT2 #(
		.INIT('h8)
	) name14212 (
		_w23516_,
		_w23521_,
		_w24724_
	);
	LUT2 #(
		.INIT('h8)
	) name14213 (
		\ethreg1_IPGR2_0_DataOut_reg[3]/NET0131 ,
		_w24724_,
		_w24725_
	);
	LUT2 #(
		.INIT('h8)
	) name14214 (
		_w23506_,
		_w23518_,
		_w24726_
	);
	LUT2 #(
		.INIT('h8)
	) name14215 (
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w24726_,
		_w24727_
	);
	LUT2 #(
		.INIT('h8)
	) name14216 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w24728_
	);
	LUT2 #(
		.INIT('h8)
	) name14217 (
		_w22964_,
		_w24728_,
		_w24729_
	);
	LUT2 #(
		.INIT('h8)
	) name14218 (
		\wb_adr_i[4]_pad ,
		_w24729_,
		_w24730_
	);
	LUT2 #(
		.INIT('h8)
	) name14219 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		_w24730_,
		_w24731_
	);
	LUT2 #(
		.INIT('h8)
	) name14220 (
		\ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 ,
		_w22956_,
		_w24732_
	);
	LUT2 #(
		.INIT('h8)
	) name14221 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		_w22959_,
		_w24733_
	);
	LUT2 #(
		.INIT('h8)
	) name14222 (
		\ethreg1_MIIRX_DATA_DataOut_reg[3]/NET0131 ,
		_w23507_,
		_w24734_
	);
	LUT2 #(
		.INIT('h8)
	) name14223 (
		\ethreg1_MODER_0_DataOut_reg[3]/NET0131 ,
		_w23519_,
		_w24735_
	);
	LUT2 #(
		.INIT('h1)
	) name14224 (
		_w24708_,
		_w24709_,
		_w24736_
	);
	LUT2 #(
		.INIT('h1)
	) name14225 (
		_w24711_,
		_w24712_,
		_w24737_
	);
	LUT2 #(
		.INIT('h1)
	) name14226 (
		_w24714_,
		_w24718_,
		_w24738_
	);
	LUT2 #(
		.INIT('h1)
	) name14227 (
		_w24719_,
		_w24720_,
		_w24739_
	);
	LUT2 #(
		.INIT('h1)
	) name14228 (
		_w24721_,
		_w24723_,
		_w24740_
	);
	LUT2 #(
		.INIT('h1)
	) name14229 (
		_w24725_,
		_w24727_,
		_w24741_
	);
	LUT2 #(
		.INIT('h1)
	) name14230 (
		_w24732_,
		_w24733_,
		_w24742_
	);
	LUT2 #(
		.INIT('h1)
	) name14231 (
		_w24734_,
		_w24735_,
		_w24743_
	);
	LUT2 #(
		.INIT('h8)
	) name14232 (
		_w24742_,
		_w24743_,
		_w24744_
	);
	LUT2 #(
		.INIT('h8)
	) name14233 (
		_w24740_,
		_w24741_,
		_w24745_
	);
	LUT2 #(
		.INIT('h8)
	) name14234 (
		_w24738_,
		_w24739_,
		_w24746_
	);
	LUT2 #(
		.INIT('h8)
	) name14235 (
		_w24736_,
		_w24737_,
		_w24747_
	);
	LUT2 #(
		.INIT('h8)
	) name14236 (
		_w22944_,
		_w24747_,
		_w24748_
	);
	LUT2 #(
		.INIT('h8)
	) name14237 (
		_w24745_,
		_w24746_,
		_w24749_
	);
	LUT2 #(
		.INIT('h4)
	) name14238 (
		_w24715_,
		_w24744_,
		_w24750_
	);
	LUT2 #(
		.INIT('h4)
	) name14239 (
		_w24731_,
		_w24750_,
		_w24751_
	);
	LUT2 #(
		.INIT('h8)
	) name14240 (
		_w24748_,
		_w24749_,
		_w24752_
	);
	LUT2 #(
		.INIT('h8)
	) name14241 (
		_w24751_,
		_w24752_,
		_w24753_
	);
	LUT2 #(
		.INIT('h1)
	) name14242 (
		_w24705_,
		_w24753_,
		_w24754_
	);
	LUT2 #(
		.INIT('h8)
	) name14243 (
		\wishbone_bd_ram_mem0_reg[0][4]/P0001 ,
		_w12717_,
		_w24755_
	);
	LUT2 #(
		.INIT('h8)
	) name14244 (
		\wishbone_bd_ram_mem0_reg[161][4]/P0001 ,
		_w12754_,
		_w24756_
	);
	LUT2 #(
		.INIT('h8)
	) name14245 (
		\wishbone_bd_ram_mem0_reg[212][4]/P0001 ,
		_w12796_,
		_w24757_
	);
	LUT2 #(
		.INIT('h8)
	) name14246 (
		\wishbone_bd_ram_mem0_reg[108][4]/P0001 ,
		_w13156_,
		_w24758_
	);
	LUT2 #(
		.INIT('h8)
	) name14247 (
		\wishbone_bd_ram_mem0_reg[156][4]/P0001 ,
		_w13190_,
		_w24759_
	);
	LUT2 #(
		.INIT('h8)
	) name14248 (
		\wishbone_bd_ram_mem0_reg[66][4]/P0001 ,
		_w12824_,
		_w24760_
	);
	LUT2 #(
		.INIT('h8)
	) name14249 (
		\wishbone_bd_ram_mem0_reg[171][4]/P0001 ,
		_w12910_,
		_w24761_
	);
	LUT2 #(
		.INIT('h8)
	) name14250 (
		\wishbone_bd_ram_mem0_reg[182][4]/P0001 ,
		_w12820_,
		_w24762_
	);
	LUT2 #(
		.INIT('h8)
	) name14251 (
		\wishbone_bd_ram_mem0_reg[3][4]/P0001 ,
		_w12866_,
		_w24763_
	);
	LUT2 #(
		.INIT('h8)
	) name14252 (
		\wishbone_bd_ram_mem0_reg[83][4]/P0001 ,
		_w12916_,
		_w24764_
	);
	LUT2 #(
		.INIT('h8)
	) name14253 (
		\wishbone_bd_ram_mem0_reg[242][4]/P0001 ,
		_w12932_,
		_w24765_
	);
	LUT2 #(
		.INIT('h8)
	) name14254 (
		\wishbone_bd_ram_mem0_reg[234][4]/P0001 ,
		_w13214_,
		_w24766_
	);
	LUT2 #(
		.INIT('h8)
	) name14255 (
		\wishbone_bd_ram_mem0_reg[1][4]/P0001 ,
		_w13014_,
		_w24767_
	);
	LUT2 #(
		.INIT('h8)
	) name14256 (
		\wishbone_bd_ram_mem0_reg[188][4]/P0001 ,
		_w12948_,
		_w24768_
	);
	LUT2 #(
		.INIT('h8)
	) name14257 (
		\wishbone_bd_ram_mem0_reg[246][4]/P0001 ,
		_w13076_,
		_w24769_
	);
	LUT2 #(
		.INIT('h8)
	) name14258 (
		\wishbone_bd_ram_mem0_reg[6][4]/P0001 ,
		_w12968_,
		_w24770_
	);
	LUT2 #(
		.INIT('h8)
	) name14259 (
		\wishbone_bd_ram_mem0_reg[58][4]/P0001 ,
		_w13070_,
		_w24771_
	);
	LUT2 #(
		.INIT('h8)
	) name14260 (
		\wishbone_bd_ram_mem0_reg[101][4]/P0001 ,
		_w13192_,
		_w24772_
	);
	LUT2 #(
		.INIT('h8)
	) name14261 (
		\wishbone_bd_ram_mem0_reg[4][4]/P0001 ,
		_w12666_,
		_w24773_
	);
	LUT2 #(
		.INIT('h8)
	) name14262 (
		\wishbone_bd_ram_mem0_reg[209][4]/P0001 ,
		_w13152_,
		_w24774_
	);
	LUT2 #(
		.INIT('h8)
	) name14263 (
		\wishbone_bd_ram_mem0_reg[141][4]/P0001 ,
		_w13004_,
		_w24775_
	);
	LUT2 #(
		.INIT('h8)
	) name14264 (
		\wishbone_bd_ram_mem0_reg[133][4]/P0001 ,
		_w12761_,
		_w24776_
	);
	LUT2 #(
		.INIT('h8)
	) name14265 (
		\wishbone_bd_ram_mem0_reg[199][4]/P0001 ,
		_w12768_,
		_w24777_
	);
	LUT2 #(
		.INIT('h8)
	) name14266 (
		\wishbone_bd_ram_mem0_reg[120][4]/P0001 ,
		_w12707_,
		_w24778_
	);
	LUT2 #(
		.INIT('h8)
	) name14267 (
		\wishbone_bd_ram_mem0_reg[228][4]/P0001 ,
		_w12765_,
		_w24779_
	);
	LUT2 #(
		.INIT('h8)
	) name14268 (
		\wishbone_bd_ram_mem0_reg[118][4]/P0001 ,
		_w12830_,
		_w24780_
	);
	LUT2 #(
		.INIT('h8)
	) name14269 (
		\wishbone_bd_ram_mem0_reg[164][4]/P0001 ,
		_w12876_,
		_w24781_
	);
	LUT2 #(
		.INIT('h8)
	) name14270 (
		\wishbone_bd_ram_mem0_reg[202][4]/P0001 ,
		_w12870_,
		_w24782_
	);
	LUT2 #(
		.INIT('h8)
	) name14271 (
		\wishbone_bd_ram_mem0_reg[241][4]/P0001 ,
		_w13006_,
		_w24783_
	);
	LUT2 #(
		.INIT('h8)
	) name14272 (
		\wishbone_bd_ram_mem0_reg[208][4]/P0001 ,
		_w13032_,
		_w24784_
	);
	LUT2 #(
		.INIT('h8)
	) name14273 (
		\wishbone_bd_ram_mem0_reg[93][4]/P0001 ,
		_w13016_,
		_w24785_
	);
	LUT2 #(
		.INIT('h8)
	) name14274 (
		\wishbone_bd_ram_mem0_reg[98][4]/P0001 ,
		_w12816_,
		_w24786_
	);
	LUT2 #(
		.INIT('h8)
	) name14275 (
		\wishbone_bd_ram_mem0_reg[100][4]/P0001 ,
		_w12960_,
		_w24787_
	);
	LUT2 #(
		.INIT('h8)
	) name14276 (
		\wishbone_bd_ram_mem0_reg[168][4]/P0001 ,
		_w13208_,
		_w24788_
	);
	LUT2 #(
		.INIT('h8)
	) name14277 (
		\wishbone_bd_ram_mem0_reg[23][4]/P0001 ,
		_w13008_,
		_w24789_
	);
	LUT2 #(
		.INIT('h8)
	) name14278 (
		\wishbone_bd_ram_mem0_reg[137][4]/P0001 ,
		_w13168_,
		_w24790_
	);
	LUT2 #(
		.INIT('h8)
	) name14279 (
		\wishbone_bd_ram_mem0_reg[88][4]/P0001 ,
		_w12860_,
		_w24791_
	);
	LUT2 #(
		.INIT('h8)
	) name14280 (
		\wishbone_bd_ram_mem0_reg[172][4]/P0001 ,
		_w12944_,
		_w24792_
	);
	LUT2 #(
		.INIT('h8)
	) name14281 (
		\wishbone_bd_ram_mem0_reg[94][4]/P0001 ,
		_w13186_,
		_w24793_
	);
	LUT2 #(
		.INIT('h8)
	) name14282 (
		\wishbone_bd_ram_mem0_reg[213][4]/P0001 ,
		_w13002_,
		_w24794_
	);
	LUT2 #(
		.INIT('h8)
	) name14283 (
		\wishbone_bd_ram_mem0_reg[140][4]/P0001 ,
		_w12894_,
		_w24795_
	);
	LUT2 #(
		.INIT('h8)
	) name14284 (
		\wishbone_bd_ram_mem0_reg[249][4]/P0001 ,
		_w12900_,
		_w24796_
	);
	LUT2 #(
		.INIT('h8)
	) name14285 (
		\wishbone_bd_ram_mem0_reg[189][4]/P0001 ,
		_w13042_,
		_w24797_
	);
	LUT2 #(
		.INIT('h8)
	) name14286 (
		\wishbone_bd_ram_mem0_reg[34][4]/P0001 ,
		_w12930_,
		_w24798_
	);
	LUT2 #(
		.INIT('h8)
	) name14287 (
		\wishbone_bd_ram_mem0_reg[33][4]/P0001 ,
		_w12980_,
		_w24799_
	);
	LUT2 #(
		.INIT('h8)
	) name14288 (
		\wishbone_bd_ram_mem0_reg[123][4]/P0001 ,
		_w13114_,
		_w24800_
	);
	LUT2 #(
		.INIT('h8)
	) name14289 (
		\wishbone_bd_ram_mem0_reg[28][4]/P0001 ,
		_w13170_,
		_w24801_
	);
	LUT2 #(
		.INIT('h8)
	) name14290 (
		\wishbone_bd_ram_mem0_reg[201][4]/P0001 ,
		_w12822_,
		_w24802_
	);
	LUT2 #(
		.INIT('h8)
	) name14291 (
		\wishbone_bd_ram_mem0_reg[203][4]/P0001 ,
		_w13158_,
		_w24803_
	);
	LUT2 #(
		.INIT('h8)
	) name14292 (
		\wishbone_bd_ram_mem0_reg[252][4]/P0001 ,
		_w13080_,
		_w24804_
	);
	LUT2 #(
		.INIT('h8)
	) name14293 (
		\wishbone_bd_ram_mem0_reg[65][4]/P0001 ,
		_w13176_,
		_w24805_
	);
	LUT2 #(
		.INIT('h8)
	) name14294 (
		\wishbone_bd_ram_mem0_reg[103][4]/P0001 ,
		_w12846_,
		_w24806_
	);
	LUT2 #(
		.INIT('h8)
	) name14295 (
		\wishbone_bd_ram_mem0_reg[240][4]/P0001 ,
		_w12864_,
		_w24807_
	);
	LUT2 #(
		.INIT('h8)
	) name14296 (
		\wishbone_bd_ram_mem0_reg[10][4]/P0001 ,
		_w13172_,
		_w24808_
	);
	LUT2 #(
		.INIT('h8)
	) name14297 (
		\wishbone_bd_ram_mem0_reg[130][4]/P0001 ,
		_w12914_,
		_w24809_
	);
	LUT2 #(
		.INIT('h8)
	) name14298 (
		\wishbone_bd_ram_mem0_reg[43][4]/P0001 ,
		_w13200_,
		_w24810_
	);
	LUT2 #(
		.INIT('h8)
	) name14299 (
		\wishbone_bd_ram_mem0_reg[177][4]/P0001 ,
		_w12996_,
		_w24811_
	);
	LUT2 #(
		.INIT('h8)
	) name14300 (
		\wishbone_bd_ram_mem0_reg[251][4]/P0001 ,
		_w13054_,
		_w24812_
	);
	LUT2 #(
		.INIT('h8)
	) name14301 (
		\wishbone_bd_ram_mem0_reg[134][4]/P0001 ,
		_w12763_,
		_w24813_
	);
	LUT2 #(
		.INIT('h8)
	) name14302 (
		\wishbone_bd_ram_mem0_reg[110][4]/P0001 ,
		_w13046_,
		_w24814_
	);
	LUT2 #(
		.INIT('h8)
	) name14303 (
		\wishbone_bd_ram_mem0_reg[207][4]/P0001 ,
		_w13180_,
		_w24815_
	);
	LUT2 #(
		.INIT('h8)
	) name14304 (
		\wishbone_bd_ram_mem0_reg[104][4]/P0001 ,
		_w13148_,
		_w24816_
	);
	LUT2 #(
		.INIT('h8)
	) name14305 (
		\wishbone_bd_ram_mem0_reg[63][4]/P0001 ,
		_w12850_,
		_w24817_
	);
	LUT2 #(
		.INIT('h8)
	) name14306 (
		\wishbone_bd_ram_mem0_reg[127][4]/P0001 ,
		_w13164_,
		_w24818_
	);
	LUT2 #(
		.INIT('h8)
	) name14307 (
		\wishbone_bd_ram_mem0_reg[226][4]/P0001 ,
		_w13138_,
		_w24819_
	);
	LUT2 #(
		.INIT('h8)
	) name14308 (
		\wishbone_bd_ram_mem0_reg[243][4]/P0001 ,
		_w12804_,
		_w24820_
	);
	LUT2 #(
		.INIT('h8)
	) name14309 (
		\wishbone_bd_ram_mem0_reg[36][4]/P0001 ,
		_w12800_,
		_w24821_
	);
	LUT2 #(
		.INIT('h8)
	) name14310 (
		\wishbone_bd_ram_mem0_reg[17][4]/P0001 ,
		_w12848_,
		_w24822_
	);
	LUT2 #(
		.INIT('h8)
	) name14311 (
		\wishbone_bd_ram_mem0_reg[145][4]/P0001 ,
		_w13106_,
		_w24823_
	);
	LUT2 #(
		.INIT('h8)
	) name14312 (
		\wishbone_bd_ram_mem0_reg[107][4]/P0001 ,
		_w12749_,
		_w24824_
	);
	LUT2 #(
		.INIT('h8)
	) name14313 (
		\wishbone_bd_ram_mem0_reg[106][4]/P0001 ,
		_w12713_,
		_w24825_
	);
	LUT2 #(
		.INIT('h8)
	) name14314 (
		\wishbone_bd_ram_mem0_reg[129][4]/P0001 ,
		_w12776_,
		_w24826_
	);
	LUT2 #(
		.INIT('h8)
	) name14315 (
		\wishbone_bd_ram_mem0_reg[12][4]/P0001 ,
		_w13118_,
		_w24827_
	);
	LUT2 #(
		.INIT('h8)
	) name14316 (
		\wishbone_bd_ram_mem0_reg[244][4]/P0001 ,
		_w12747_,
		_w24828_
	);
	LUT2 #(
		.INIT('h8)
	) name14317 (
		\wishbone_bd_ram_mem0_reg[143][4]/P0001 ,
		_w12922_,
		_w24829_
	);
	LUT2 #(
		.INIT('h8)
	) name14318 (
		\wishbone_bd_ram_mem0_reg[97][4]/P0001 ,
		_w13096_,
		_w24830_
	);
	LUT2 #(
		.INIT('h8)
	) name14319 (
		\wishbone_bd_ram_mem0_reg[231][4]/P0001 ,
		_w12856_,
		_w24831_
	);
	LUT2 #(
		.INIT('h8)
	) name14320 (
		\wishbone_bd_ram_mem0_reg[253][4]/P0001 ,
		_w13100_,
		_w24832_
	);
	LUT2 #(
		.INIT('h8)
	) name14321 (
		\wishbone_bd_ram_mem0_reg[225][4]/P0001 ,
		_w13092_,
		_w24833_
	);
	LUT2 #(
		.INIT('h8)
	) name14322 (
		\wishbone_bd_ram_mem0_reg[5][4]/P0001 ,
		_w12878_,
		_w24834_
	);
	LUT2 #(
		.INIT('h8)
	) name14323 (
		\wishbone_bd_ram_mem0_reg[54][4]/P0001 ,
		_w12770_,
		_w24835_
	);
	LUT2 #(
		.INIT('h8)
	) name14324 (
		\wishbone_bd_ram_mem0_reg[87][4]/P0001 ,
		_w13154_,
		_w24836_
	);
	LUT2 #(
		.INIT('h8)
	) name14325 (
		\wishbone_bd_ram_mem0_reg[119][4]/P0001 ,
		_w13048_,
		_w24837_
	);
	LUT2 #(
		.INIT('h8)
	) name14326 (
		\wishbone_bd_ram_mem0_reg[37][4]/P0001 ,
		_w13102_,
		_w24838_
	);
	LUT2 #(
		.INIT('h8)
	) name14327 (
		\wishbone_bd_ram_mem0_reg[61][4]/P0001 ,
		_w12725_,
		_w24839_
	);
	LUT2 #(
		.INIT('h8)
	) name14328 (
		\wishbone_bd_ram_mem0_reg[72][4]/P0001 ,
		_w12810_,
		_w24840_
	);
	LUT2 #(
		.INIT('h8)
	) name14329 (
		\wishbone_bd_ram_mem0_reg[9][4]/P0001 ,
		_w12808_,
		_w24841_
	);
	LUT2 #(
		.INIT('h8)
	) name14330 (
		\wishbone_bd_ram_mem0_reg[35][4]/P0001 ,
		_w12703_,
		_w24842_
	);
	LUT2 #(
		.INIT('h8)
	) name14331 (
		\wishbone_bd_ram_mem0_reg[22][4]/P0001 ,
		_w13110_,
		_w24843_
	);
	LUT2 #(
		.INIT('h8)
	) name14332 (
		\wishbone_bd_ram_mem0_reg[187][4]/P0001 ,
		_w13196_,
		_w24844_
	);
	LUT2 #(
		.INIT('h8)
	) name14333 (
		\wishbone_bd_ram_mem0_reg[25][4]/P0001 ,
		_w13108_,
		_w24845_
	);
	LUT2 #(
		.INIT('h8)
	) name14334 (
		\wishbone_bd_ram_mem0_reg[146][4]/P0001 ,
		_w13060_,
		_w24846_
	);
	LUT2 #(
		.INIT('h8)
	) name14335 (
		\wishbone_bd_ram_mem0_reg[48][4]/P0001 ,
		_w12970_,
		_w24847_
	);
	LUT2 #(
		.INIT('h8)
	) name14336 (
		\wishbone_bd_ram_mem0_reg[95][4]/P0001 ,
		_w12844_,
		_w24848_
	);
	LUT2 #(
		.INIT('h8)
	) name14337 (
		\wishbone_bd_ram_mem0_reg[62][4]/P0001 ,
		_w12673_,
		_w24849_
	);
	LUT2 #(
		.INIT('h8)
	) name14338 (
		\wishbone_bd_ram_mem0_reg[139][4]/P0001 ,
		_w12814_,
		_w24850_
	);
	LUT2 #(
		.INIT('h8)
	) name14339 (
		\wishbone_bd_ram_mem0_reg[215][4]/P0001 ,
		_w12974_,
		_w24851_
	);
	LUT2 #(
		.INIT('h8)
	) name14340 (
		\wishbone_bd_ram_mem0_reg[175][4]/P0001 ,
		_w13126_,
		_w24852_
	);
	LUT2 #(
		.INIT('h8)
	) name14341 (
		\wishbone_bd_ram_mem0_reg[60][4]/P0001 ,
		_w13204_,
		_w24853_
	);
	LUT2 #(
		.INIT('h8)
	) name14342 (
		\wishbone_bd_ram_mem0_reg[193][4]/P0001 ,
		_w13056_,
		_w24854_
	);
	LUT2 #(
		.INIT('h8)
	) name14343 (
		\wishbone_bd_ram_mem0_reg[55][4]/P0001 ,
		_w12785_,
		_w24855_
	);
	LUT2 #(
		.INIT('h8)
	) name14344 (
		\wishbone_bd_ram_mem0_reg[77][4]/P0001 ,
		_w12982_,
		_w24856_
	);
	LUT2 #(
		.INIT('h8)
	) name14345 (
		\wishbone_bd_ram_mem0_reg[153][4]/P0001 ,
		_w12890_,
		_w24857_
	);
	LUT2 #(
		.INIT('h8)
	) name14346 (
		\wishbone_bd_ram_mem0_reg[192][4]/P0001 ,
		_w12938_,
		_w24858_
	);
	LUT2 #(
		.INIT('h8)
	) name14347 (
		\wishbone_bd_ram_mem0_reg[51][4]/P0001 ,
		_w13024_,
		_w24859_
	);
	LUT2 #(
		.INIT('h8)
	) name14348 (
		\wishbone_bd_ram_mem0_reg[206][4]/P0001 ,
		_w12954_,
		_w24860_
	);
	LUT2 #(
		.INIT('h8)
	) name14349 (
		\wishbone_bd_ram_mem0_reg[173][4]/P0001 ,
		_w12854_,
		_w24861_
	);
	LUT2 #(
		.INIT('h8)
	) name14350 (
		\wishbone_bd_ram_mem0_reg[39][4]/P0001 ,
		_w13018_,
		_w24862_
	);
	LUT2 #(
		.INIT('h8)
	) name14351 (
		\wishbone_bd_ram_mem0_reg[196][4]/P0001 ,
		_w13090_,
		_w24863_
	);
	LUT2 #(
		.INIT('h8)
	) name14352 (
		\wishbone_bd_ram_mem0_reg[135][4]/P0001 ,
		_w13124_,
		_w24864_
	);
	LUT2 #(
		.INIT('h8)
	) name14353 (
		\wishbone_bd_ram_mem0_reg[82][4]/P0001 ,
		_w12942_,
		_w24865_
	);
	LUT2 #(
		.INIT('h8)
	) name14354 (
		\wishbone_bd_ram_mem0_reg[166][4]/P0001 ,
		_w13040_,
		_w24866_
	);
	LUT2 #(
		.INIT('h8)
	) name14355 (
		\wishbone_bd_ram_mem0_reg[236][4]/P0001 ,
		_w12731_,
		_w24867_
	);
	LUT2 #(
		.INIT('h8)
	) name14356 (
		\wishbone_bd_ram_mem0_reg[157][4]/P0001 ,
		_w12926_,
		_w24868_
	);
	LUT2 #(
		.INIT('h8)
	) name14357 (
		\wishbone_bd_ram_mem0_reg[111][4]/P0001 ,
		_w12744_,
		_w24869_
	);
	LUT2 #(
		.INIT('h8)
	) name14358 (
		\wishbone_bd_ram_mem0_reg[49][4]/P0001 ,
		_w12994_,
		_w24870_
	);
	LUT2 #(
		.INIT('h8)
	) name14359 (
		\wishbone_bd_ram_mem0_reg[179][4]/P0001 ,
		_w13050_,
		_w24871_
	);
	LUT2 #(
		.INIT('h8)
	) name14360 (
		\wishbone_bd_ram_mem0_reg[184][4]/P0001 ,
		_w13062_,
		_w24872_
	);
	LUT2 #(
		.INIT('h8)
	) name14361 (
		\wishbone_bd_ram_mem0_reg[237][4]/P0001 ,
		_w12990_,
		_w24873_
	);
	LUT2 #(
		.INIT('h8)
	) name14362 (
		\wishbone_bd_ram_mem0_reg[21][4]/P0001 ,
		_w12906_,
		_w24874_
	);
	LUT2 #(
		.INIT('h8)
	) name14363 (
		\wishbone_bd_ram_mem0_reg[165][4]/P0001 ,
		_w13044_,
		_w24875_
	);
	LUT2 #(
		.INIT('h8)
	) name14364 (
		\wishbone_bd_ram_mem0_reg[147][4]/P0001 ,
		_w13146_,
		_w24876_
	);
	LUT2 #(
		.INIT('h8)
	) name14365 (
		\wishbone_bd_ram_mem0_reg[38][4]/P0001 ,
		_w13182_,
		_w24877_
	);
	LUT2 #(
		.INIT('h8)
	) name14366 (
		\wishbone_bd_ram_mem0_reg[233][4]/P0001 ,
		_w12836_,
		_w24878_
	);
	LUT2 #(
		.INIT('h8)
	) name14367 (
		\wishbone_bd_ram_mem0_reg[86][4]/P0001 ,
		_w12735_,
		_w24879_
	);
	LUT2 #(
		.INIT('h8)
	) name14368 (
		\wishbone_bd_ram_mem0_reg[14][4]/P0001 ,
		_w13086_,
		_w24880_
	);
	LUT2 #(
		.INIT('h8)
	) name14369 (
		\wishbone_bd_ram_mem0_reg[116][4]/P0001 ,
		_w12998_,
		_w24881_
	);
	LUT2 #(
		.INIT('h8)
	) name14370 (
		\wishbone_bd_ram_mem0_reg[186][4]/P0001 ,
		_w12783_,
		_w24882_
	);
	LUT2 #(
		.INIT('h8)
	) name14371 (
		\wishbone_bd_ram_mem0_reg[148][4]/P0001 ,
		_w13000_,
		_w24883_
	);
	LUT2 #(
		.INIT('h8)
	) name14372 (
		\wishbone_bd_ram_mem0_reg[167][4]/P0001 ,
		_w12986_,
		_w24884_
	);
	LUT2 #(
		.INIT('h8)
	) name14373 (
		\wishbone_bd_ram_mem0_reg[216][4]/P0001 ,
		_w13028_,
		_w24885_
	);
	LUT2 #(
		.INIT('h8)
	) name14374 (
		\wishbone_bd_ram_mem0_reg[11][4]/P0001 ,
		_w13194_,
		_w24886_
	);
	LUT2 #(
		.INIT('h8)
	) name14375 (
		\wishbone_bd_ram_mem0_reg[47][4]/P0001 ,
		_w12904_,
		_w24887_
	);
	LUT2 #(
		.INIT('h8)
	) name14376 (
		\wishbone_bd_ram_mem0_reg[181][4]/P0001 ,
		_w12828_,
		_w24888_
	);
	LUT2 #(
		.INIT('h8)
	) name14377 (
		\wishbone_bd_ram_mem0_reg[20][4]/P0001 ,
		_w13174_,
		_w24889_
	);
	LUT2 #(
		.INIT('h8)
	) name14378 (
		\wishbone_bd_ram_mem0_reg[155][4]/P0001 ,
		_w13122_,
		_w24890_
	);
	LUT2 #(
		.INIT('h8)
	) name14379 (
		\wishbone_bd_ram_mem0_reg[40][4]/P0001 ,
		_w13132_,
		_w24891_
	);
	LUT2 #(
		.INIT('h8)
	) name14380 (
		\wishbone_bd_ram_mem0_reg[149][4]/P0001 ,
		_w12741_,
		_w24892_
	);
	LUT2 #(
		.INIT('h8)
	) name14381 (
		\wishbone_bd_ram_mem0_reg[250][4]/P0001 ,
		_w13128_,
		_w24893_
	);
	LUT2 #(
		.INIT('h8)
	) name14382 (
		\wishbone_bd_ram_mem0_reg[138][4]/P0001 ,
		_w12958_,
		_w24894_
	);
	LUT2 #(
		.INIT('h8)
	) name14383 (
		\wishbone_bd_ram_mem0_reg[68][4]/P0001 ,
		_w12946_,
		_w24895_
	);
	LUT2 #(
		.INIT('h8)
	) name14384 (
		\wishbone_bd_ram_mem0_reg[198][4]/P0001 ,
		_w12832_,
		_w24896_
	);
	LUT2 #(
		.INIT('h8)
	) name14385 (
		\wishbone_bd_ram_mem0_reg[176][4]/P0001 ,
		_w12868_,
		_w24897_
	);
	LUT2 #(
		.INIT('h8)
	) name14386 (
		\wishbone_bd_ram_mem0_reg[26][4]/P0001 ,
		_w12699_,
		_w24898_
	);
	LUT2 #(
		.INIT('h8)
	) name14387 (
		\wishbone_bd_ram_mem0_reg[230][4]/P0001 ,
		_w13036_,
		_w24899_
	);
	LUT2 #(
		.INIT('h8)
	) name14388 (
		\wishbone_bd_ram_mem0_reg[45][4]/P0001 ,
		_w12908_,
		_w24900_
	);
	LUT2 #(
		.INIT('h8)
	) name14389 (
		\wishbone_bd_ram_mem0_reg[160][4]/P0001 ,
		_w12872_,
		_w24901_
	);
	LUT2 #(
		.INIT('h8)
	) name14390 (
		\wishbone_bd_ram_mem0_reg[41][4]/P0001 ,
		_w13052_,
		_w24902_
	);
	LUT2 #(
		.INIT('h8)
	) name14391 (
		\wishbone_bd_ram_mem0_reg[80][4]/P0001 ,
		_w12689_,
		_w24903_
	);
	LUT2 #(
		.INIT('h8)
	) name14392 (
		\wishbone_bd_ram_mem0_reg[53][4]/P0001 ,
		_w13020_,
		_w24904_
	);
	LUT2 #(
		.INIT('h8)
	) name14393 (
		\wishbone_bd_ram_mem0_reg[59][4]/P0001 ,
		_w12780_,
		_w24905_
	);
	LUT2 #(
		.INIT('h8)
	) name14394 (
		\wishbone_bd_ram_mem0_reg[150][4]/P0001 ,
		_w13136_,
		_w24906_
	);
	LUT2 #(
		.INIT('h8)
	) name14395 (
		\wishbone_bd_ram_mem0_reg[109][4]/P0001 ,
		_w12888_,
		_w24907_
	);
	LUT2 #(
		.INIT('h8)
	) name14396 (
		\wishbone_bd_ram_mem0_reg[170][4]/P0001 ,
		_w13030_,
		_w24908_
	);
	LUT2 #(
		.INIT('h8)
	) name14397 (
		\wishbone_bd_ram_mem0_reg[32][4]/P0001 ,
		_w13120_,
		_w24909_
	);
	LUT2 #(
		.INIT('h8)
	) name14398 (
		\wishbone_bd_ram_mem0_reg[128][4]/P0001 ,
		_w12793_,
		_w24910_
	);
	LUT2 #(
		.INIT('h8)
	) name14399 (
		\wishbone_bd_ram_mem0_reg[117][4]/P0001 ,
		_w12715_,
		_w24911_
	);
	LUT2 #(
		.INIT('h8)
	) name14400 (
		\wishbone_bd_ram_mem0_reg[70][4]/P0001 ,
		_w12840_,
		_w24912_
	);
	LUT2 #(
		.INIT('h8)
	) name14401 (
		\wishbone_bd_ram_mem0_reg[115][4]/P0001 ,
		_w13112_,
		_w24913_
	);
	LUT2 #(
		.INIT('h8)
	) name14402 (
		\wishbone_bd_ram_mem0_reg[183][4]/P0001 ,
		_w12787_,
		_w24914_
	);
	LUT2 #(
		.INIT('h8)
	) name14403 (
		\wishbone_bd_ram_mem0_reg[238][4]/P0001 ,
		_w13160_,
		_w24915_
	);
	LUT2 #(
		.INIT('h8)
	) name14404 (
		\wishbone_bd_ram_mem0_reg[200][4]/P0001 ,
		_w12988_,
		_w24916_
	);
	LUT2 #(
		.INIT('h8)
	) name14405 (
		\wishbone_bd_ram_mem0_reg[122][4]/P0001 ,
		_w13130_,
		_w24917_
	);
	LUT2 #(
		.INIT('h8)
	) name14406 (
		\wishbone_bd_ram_mem0_reg[235][4]/P0001 ,
		_w12696_,
		_w24918_
	);
	LUT2 #(
		.INIT('h8)
	) name14407 (
		\wishbone_bd_ram_mem0_reg[151][4]/P0001 ,
		_w13142_,
		_w24919_
	);
	LUT2 #(
		.INIT('h8)
	) name14408 (
		\wishbone_bd_ram_mem0_reg[131][4]/P0001 ,
		_w12852_,
		_w24920_
	);
	LUT2 #(
		.INIT('h8)
	) name14409 (
		\wishbone_bd_ram_mem0_reg[144][4]/P0001 ,
		_w12756_,
		_w24921_
	);
	LUT2 #(
		.INIT('h8)
	) name14410 (
		\wishbone_bd_ram_mem0_reg[102][4]/P0001 ,
		_w12685_,
		_w24922_
	);
	LUT2 #(
		.INIT('h8)
	) name14411 (
		\wishbone_bd_ram_mem0_reg[99][4]/P0001 ,
		_w13038_,
		_w24923_
	);
	LUT2 #(
		.INIT('h8)
	) name14412 (
		\wishbone_bd_ram_mem0_reg[158][4]/P0001 ,
		_w12898_,
		_w24924_
	);
	LUT2 #(
		.INIT('h8)
	) name14413 (
		\wishbone_bd_ram_mem0_reg[8][4]/P0001 ,
		_w12920_,
		_w24925_
	);
	LUT2 #(
		.INIT('h8)
	) name14414 (
		\wishbone_bd_ram_mem0_reg[85][4]/P0001 ,
		_w13216_,
		_w24926_
	);
	LUT2 #(
		.INIT('h8)
	) name14415 (
		\wishbone_bd_ram_mem0_reg[46][4]/P0001 ,
		_w12884_,
		_w24927_
	);
	LUT2 #(
		.INIT('h8)
	) name14416 (
		\wishbone_bd_ram_mem0_reg[44][4]/P0001 ,
		_w12896_,
		_w24928_
	);
	LUT2 #(
		.INIT('h8)
	) name14417 (
		\wishbone_bd_ram_mem0_reg[195][4]/P0001 ,
		_w13144_,
		_w24929_
	);
	LUT2 #(
		.INIT('h8)
	) name14418 (
		\wishbone_bd_ram_mem0_reg[112][4]/P0001 ,
		_w12733_,
		_w24930_
	);
	LUT2 #(
		.INIT('h8)
	) name14419 (
		\wishbone_bd_ram_mem0_reg[90][4]/P0001 ,
		_w12978_,
		_w24931_
	);
	LUT2 #(
		.INIT('h8)
	) name14420 (
		\wishbone_bd_ram_mem0_reg[210][4]/P0001 ,
		_w12924_,
		_w24932_
	);
	LUT2 #(
		.INIT('h8)
	) name14421 (
		\wishbone_bd_ram_mem0_reg[71][4]/P0001 ,
		_w12798_,
		_w24933_
	);
	LUT2 #(
		.INIT('h8)
	) name14422 (
		\wishbone_bd_ram_mem0_reg[191][4]/P0001 ,
		_w13034_,
		_w24934_
	);
	LUT2 #(
		.INIT('h8)
	) name14423 (
		\wishbone_bd_ram_mem0_reg[223][4]/P0001 ,
		_w12838_,
		_w24935_
	);
	LUT2 #(
		.INIT('h8)
	) name14424 (
		\wishbone_bd_ram_mem0_reg[27][4]/P0001 ,
		_w12880_,
		_w24936_
	);
	LUT2 #(
		.INIT('h8)
	) name14425 (
		\wishbone_bd_ram_mem0_reg[247][4]/P0001 ,
		_w12818_,
		_w24937_
	);
	LUT2 #(
		.INIT('h8)
	) name14426 (
		\wishbone_bd_ram_mem0_reg[152][4]/P0001 ,
		_w12966_,
		_w24938_
	);
	LUT2 #(
		.INIT('h8)
	) name14427 (
		\wishbone_bd_ram_mem0_reg[239][4]/P0001 ,
		_w12862_,
		_w24939_
	);
	LUT2 #(
		.INIT('h8)
	) name14428 (
		\wishbone_bd_ram_mem0_reg[174][4]/P0001 ,
		_w12972_,
		_w24940_
	);
	LUT2 #(
		.INIT('h8)
	) name14429 (
		\wishbone_bd_ram_mem0_reg[245][4]/P0001 ,
		_w13022_,
		_w24941_
	);
	LUT2 #(
		.INIT('h8)
	) name14430 (
		\wishbone_bd_ram_mem0_reg[16][4]/P0001 ,
		_w13140_,
		_w24942_
	);
	LUT2 #(
		.INIT('h8)
	) name14431 (
		\wishbone_bd_ram_mem0_reg[121][4]/P0001 ,
		_w13078_,
		_w24943_
	);
	LUT2 #(
		.INIT('h8)
	) name14432 (
		\wishbone_bd_ram_mem0_reg[214][4]/P0001 ,
		_w12984_,
		_w24944_
	);
	LUT2 #(
		.INIT('h8)
	) name14433 (
		\wishbone_bd_ram_mem0_reg[67][4]/P0001 ,
		_w13134_,
		_w24945_
	);
	LUT2 #(
		.INIT('h8)
	) name14434 (
		\wishbone_bd_ram_mem0_reg[124][4]/P0001 ,
		_w13058_,
		_w24946_
	);
	LUT2 #(
		.INIT('h8)
	) name14435 (
		\wishbone_bd_ram_mem0_reg[254][4]/P0001 ,
		_w12892_,
		_w24947_
	);
	LUT2 #(
		.INIT('h8)
	) name14436 (
		\wishbone_bd_ram_mem0_reg[91][4]/P0001 ,
		_w13074_,
		_w24948_
	);
	LUT2 #(
		.INIT('h8)
	) name14437 (
		\wishbone_bd_ram_mem0_reg[222][4]/P0001 ,
		_w13094_,
		_w24949_
	);
	LUT2 #(
		.INIT('h8)
	) name14438 (
		\wishbone_bd_ram_mem0_reg[154][4]/P0001 ,
		_w12962_,
		_w24950_
	);
	LUT2 #(
		.INIT('h8)
	) name14439 (
		\wishbone_bd_ram_mem0_reg[229][4]/P0001 ,
		_w12711_,
		_w24951_
	);
	LUT2 #(
		.INIT('h8)
	) name14440 (
		\wishbone_bd_ram_mem0_reg[52][4]/P0001 ,
		_w13082_,
		_w24952_
	);
	LUT2 #(
		.INIT('h8)
	) name14441 (
		\wishbone_bd_ram_mem0_reg[126][4]/P0001 ,
		_w13218_,
		_w24953_
	);
	LUT2 #(
		.INIT('h8)
	) name14442 (
		\wishbone_bd_ram_mem0_reg[89][4]/P0001 ,
		_w12964_,
		_w24954_
	);
	LUT2 #(
		.INIT('h8)
	) name14443 (
		\wishbone_bd_ram_mem0_reg[219][4]/P0001 ,
		_w12806_,
		_w24955_
	);
	LUT2 #(
		.INIT('h8)
	) name14444 (
		\wishbone_bd_ram_mem0_reg[31][4]/P0001 ,
		_w13198_,
		_w24956_
	);
	LUT2 #(
		.INIT('h8)
	) name14445 (
		\wishbone_bd_ram_mem0_reg[248][4]/P0001 ,
		_w12789_,
		_w24957_
	);
	LUT2 #(
		.INIT('h8)
	) name14446 (
		\wishbone_bd_ram_mem0_reg[81][4]/P0001 ,
		_w12950_,
		_w24958_
	);
	LUT2 #(
		.INIT('h8)
	) name14447 (
		\wishbone_bd_ram_mem0_reg[69][4]/P0001 ,
		_w12738_,
		_w24959_
	);
	LUT2 #(
		.INIT('h8)
	) name14448 (
		\wishbone_bd_ram_mem0_reg[42][4]/P0001 ,
		_w12842_,
		_w24960_
	);
	LUT2 #(
		.INIT('h8)
	) name14449 (
		\wishbone_bd_ram_mem0_reg[7][4]/P0001 ,
		_w12728_,
		_w24961_
	);
	LUT2 #(
		.INIT('h8)
	) name14450 (
		\wishbone_bd_ram_mem0_reg[19][4]/P0001 ,
		_w13012_,
		_w24962_
	);
	LUT2 #(
		.INIT('h8)
	) name14451 (
		\wishbone_bd_ram_mem0_reg[64][4]/P0001 ,
		_w12976_,
		_w24963_
	);
	LUT2 #(
		.INIT('h8)
	) name14452 (
		\wishbone_bd_ram_mem0_reg[113][4]/P0001 ,
		_w13026_,
		_w24964_
	);
	LUT2 #(
		.INIT('h8)
	) name14453 (
		\wishbone_bd_ram_mem0_reg[227][4]/P0001 ,
		_w12936_,
		_w24965_
	);
	LUT2 #(
		.INIT('h8)
	) name14454 (
		\wishbone_bd_ram_mem0_reg[105][4]/P0001 ,
		_w12751_,
		_w24966_
	);
	LUT2 #(
		.INIT('h8)
	) name14455 (
		\wishbone_bd_ram_mem0_reg[13][4]/P0001 ,
		_w13178_,
		_w24967_
	);
	LUT2 #(
		.INIT('h8)
	) name14456 (
		\wishbone_bd_ram_mem0_reg[114][4]/P0001 ,
		_w13202_,
		_w24968_
	);
	LUT2 #(
		.INIT('h8)
	) name14457 (
		\wishbone_bd_ram_mem0_reg[142][4]/P0001 ,
		_w12928_,
		_w24969_
	);
	LUT2 #(
		.INIT('h8)
	) name14458 (
		\wishbone_bd_ram_mem0_reg[178][4]/P0001 ,
		_w12886_,
		_w24970_
	);
	LUT2 #(
		.INIT('h8)
	) name14459 (
		\wishbone_bd_ram_mem0_reg[56][4]/P0001 ,
		_w12778_,
		_w24971_
	);
	LUT2 #(
		.INIT('h8)
	) name14460 (
		\wishbone_bd_ram_mem0_reg[84][4]/P0001 ,
		_w12934_,
		_w24972_
	);
	LUT2 #(
		.INIT('h8)
	) name14461 (
		\wishbone_bd_ram_mem0_reg[232][4]/P0001 ,
		_w12758_,
		_w24973_
	);
	LUT2 #(
		.INIT('h8)
	) name14462 (
		\wishbone_bd_ram_mem0_reg[159][4]/P0001 ,
		_w12774_,
		_w24974_
	);
	LUT2 #(
		.INIT('h8)
	) name14463 (
		\wishbone_bd_ram_mem0_reg[125][4]/P0001 ,
		_w12956_,
		_w24975_
	);
	LUT2 #(
		.INIT('h8)
	) name14464 (
		\wishbone_bd_ram_mem0_reg[30][4]/P0001 ,
		_w13104_,
		_w24976_
	);
	LUT2 #(
		.INIT('h8)
	) name14465 (
		\wishbone_bd_ram_mem0_reg[220][4]/P0001 ,
		_w13066_,
		_w24977_
	);
	LUT2 #(
		.INIT('h8)
	) name14466 (
		\wishbone_bd_ram_mem0_reg[218][4]/P0001 ,
		_w13206_,
		_w24978_
	);
	LUT2 #(
		.INIT('h8)
	) name14467 (
		\wishbone_bd_ram_mem0_reg[57][4]/P0001 ,
		_w13116_,
		_w24979_
	);
	LUT2 #(
		.INIT('h8)
	) name14468 (
		\wishbone_bd_ram_mem0_reg[79][4]/P0001 ,
		_w13212_,
		_w24980_
	);
	LUT2 #(
		.INIT('h8)
	) name14469 (
		\wishbone_bd_ram_mem0_reg[163][4]/P0001 ,
		_w12882_,
		_w24981_
	);
	LUT2 #(
		.INIT('h8)
	) name14470 (
		\wishbone_bd_ram_mem0_reg[211][4]/P0001 ,
		_w13166_,
		_w24982_
	);
	LUT2 #(
		.INIT('h8)
	) name14471 (
		\wishbone_bd_ram_mem0_reg[185][4]/P0001 ,
		_w12940_,
		_w24983_
	);
	LUT2 #(
		.INIT('h8)
	) name14472 (
		\wishbone_bd_ram_mem0_reg[197][4]/P0001 ,
		_w12834_,
		_w24984_
	);
	LUT2 #(
		.INIT('h8)
	) name14473 (
		\wishbone_bd_ram_mem0_reg[169][4]/P0001 ,
		_w12722_,
		_w24985_
	);
	LUT2 #(
		.INIT('h8)
	) name14474 (
		\wishbone_bd_ram_mem0_reg[73][4]/P0001 ,
		_w12918_,
		_w24986_
	);
	LUT2 #(
		.INIT('h8)
	) name14475 (
		\wishbone_bd_ram_mem0_reg[15][4]/P0001 ,
		_w13210_,
		_w24987_
	);
	LUT2 #(
		.INIT('h8)
	) name14476 (
		\wishbone_bd_ram_mem0_reg[78][4]/P0001 ,
		_w12874_,
		_w24988_
	);
	LUT2 #(
		.INIT('h8)
	) name14477 (
		\wishbone_bd_ram_mem0_reg[204][4]/P0001 ,
		_w13162_,
		_w24989_
	);
	LUT2 #(
		.INIT('h8)
	) name14478 (
		\wishbone_bd_ram_mem0_reg[24][4]/P0001 ,
		_w13084_,
		_w24990_
	);
	LUT2 #(
		.INIT('h8)
	) name14479 (
		\wishbone_bd_ram_mem0_reg[190][4]/P0001 ,
		_w12858_,
		_w24991_
	);
	LUT2 #(
		.INIT('h8)
	) name14480 (
		\wishbone_bd_ram_mem0_reg[18][4]/P0001 ,
		_w12679_,
		_w24992_
	);
	LUT2 #(
		.INIT('h8)
	) name14481 (
		\wishbone_bd_ram_mem0_reg[217][4]/P0001 ,
		_w13188_,
		_w24993_
	);
	LUT2 #(
		.INIT('h8)
	) name14482 (
		\wishbone_bd_ram_mem0_reg[205][4]/P0001 ,
		_w13068_,
		_w24994_
	);
	LUT2 #(
		.INIT('h8)
	) name14483 (
		\wishbone_bd_ram_mem0_reg[221][4]/P0001 ,
		_w12802_,
		_w24995_
	);
	LUT2 #(
		.INIT('h8)
	) name14484 (
		\wishbone_bd_ram_mem0_reg[180][4]/P0001 ,
		_w12791_,
		_w24996_
	);
	LUT2 #(
		.INIT('h8)
	) name14485 (
		\wishbone_bd_ram_mem0_reg[76][4]/P0001 ,
		_w13184_,
		_w24997_
	);
	LUT2 #(
		.INIT('h8)
	) name14486 (
		\wishbone_bd_ram_mem0_reg[74][4]/P0001 ,
		_w12812_,
		_w24998_
	);
	LUT2 #(
		.INIT('h8)
	) name14487 (
		\wishbone_bd_ram_mem0_reg[194][4]/P0001 ,
		_w12772_,
		_w24999_
	);
	LUT2 #(
		.INIT('h8)
	) name14488 (
		\wishbone_bd_ram_mem0_reg[132][4]/P0001 ,
		_w12992_,
		_w25000_
	);
	LUT2 #(
		.INIT('h8)
	) name14489 (
		\wishbone_bd_ram_mem0_reg[2][4]/P0001 ,
		_w13088_,
		_w25001_
	);
	LUT2 #(
		.INIT('h8)
	) name14490 (
		\wishbone_bd_ram_mem0_reg[255][4]/P0001 ,
		_w13072_,
		_w25002_
	);
	LUT2 #(
		.INIT('h8)
	) name14491 (
		\wishbone_bd_ram_mem0_reg[29][4]/P0001 ,
		_w12952_,
		_w25003_
	);
	LUT2 #(
		.INIT('h8)
	) name14492 (
		\wishbone_bd_ram_mem0_reg[136][4]/P0001 ,
		_w13064_,
		_w25004_
	);
	LUT2 #(
		.INIT('h8)
	) name14493 (
		\wishbone_bd_ram_mem0_reg[162][4]/P0001 ,
		_w13098_,
		_w25005_
	);
	LUT2 #(
		.INIT('h8)
	) name14494 (
		\wishbone_bd_ram_mem0_reg[75][4]/P0001 ,
		_w12826_,
		_w25006_
	);
	LUT2 #(
		.INIT('h8)
	) name14495 (
		\wishbone_bd_ram_mem0_reg[50][4]/P0001 ,
		_w13150_,
		_w25007_
	);
	LUT2 #(
		.INIT('h8)
	) name14496 (
		\wishbone_bd_ram_mem0_reg[92][4]/P0001 ,
		_w13010_,
		_w25008_
	);
	LUT2 #(
		.INIT('h8)
	) name14497 (
		\wishbone_bd_ram_mem0_reg[96][4]/P0001 ,
		_w12912_,
		_w25009_
	);
	LUT2 #(
		.INIT('h8)
	) name14498 (
		\wishbone_bd_ram_mem0_reg[224][4]/P0001 ,
		_w12902_,
		_w25010_
	);
	LUT2 #(
		.INIT('h1)
	) name14499 (
		_w24755_,
		_w24756_,
		_w25011_
	);
	LUT2 #(
		.INIT('h1)
	) name14500 (
		_w24757_,
		_w24758_,
		_w25012_
	);
	LUT2 #(
		.INIT('h1)
	) name14501 (
		_w24759_,
		_w24760_,
		_w25013_
	);
	LUT2 #(
		.INIT('h1)
	) name14502 (
		_w24761_,
		_w24762_,
		_w25014_
	);
	LUT2 #(
		.INIT('h1)
	) name14503 (
		_w24763_,
		_w24764_,
		_w25015_
	);
	LUT2 #(
		.INIT('h1)
	) name14504 (
		_w24765_,
		_w24766_,
		_w25016_
	);
	LUT2 #(
		.INIT('h1)
	) name14505 (
		_w24767_,
		_w24768_,
		_w25017_
	);
	LUT2 #(
		.INIT('h1)
	) name14506 (
		_w24769_,
		_w24770_,
		_w25018_
	);
	LUT2 #(
		.INIT('h1)
	) name14507 (
		_w24771_,
		_w24772_,
		_w25019_
	);
	LUT2 #(
		.INIT('h1)
	) name14508 (
		_w24773_,
		_w24774_,
		_w25020_
	);
	LUT2 #(
		.INIT('h1)
	) name14509 (
		_w24775_,
		_w24776_,
		_w25021_
	);
	LUT2 #(
		.INIT('h1)
	) name14510 (
		_w24777_,
		_w24778_,
		_w25022_
	);
	LUT2 #(
		.INIT('h1)
	) name14511 (
		_w24779_,
		_w24780_,
		_w25023_
	);
	LUT2 #(
		.INIT('h1)
	) name14512 (
		_w24781_,
		_w24782_,
		_w25024_
	);
	LUT2 #(
		.INIT('h1)
	) name14513 (
		_w24783_,
		_w24784_,
		_w25025_
	);
	LUT2 #(
		.INIT('h1)
	) name14514 (
		_w24785_,
		_w24786_,
		_w25026_
	);
	LUT2 #(
		.INIT('h1)
	) name14515 (
		_w24787_,
		_w24788_,
		_w25027_
	);
	LUT2 #(
		.INIT('h1)
	) name14516 (
		_w24789_,
		_w24790_,
		_w25028_
	);
	LUT2 #(
		.INIT('h1)
	) name14517 (
		_w24791_,
		_w24792_,
		_w25029_
	);
	LUT2 #(
		.INIT('h1)
	) name14518 (
		_w24793_,
		_w24794_,
		_w25030_
	);
	LUT2 #(
		.INIT('h1)
	) name14519 (
		_w24795_,
		_w24796_,
		_w25031_
	);
	LUT2 #(
		.INIT('h1)
	) name14520 (
		_w24797_,
		_w24798_,
		_w25032_
	);
	LUT2 #(
		.INIT('h1)
	) name14521 (
		_w24799_,
		_w24800_,
		_w25033_
	);
	LUT2 #(
		.INIT('h1)
	) name14522 (
		_w24801_,
		_w24802_,
		_w25034_
	);
	LUT2 #(
		.INIT('h1)
	) name14523 (
		_w24803_,
		_w24804_,
		_w25035_
	);
	LUT2 #(
		.INIT('h1)
	) name14524 (
		_w24805_,
		_w24806_,
		_w25036_
	);
	LUT2 #(
		.INIT('h1)
	) name14525 (
		_w24807_,
		_w24808_,
		_w25037_
	);
	LUT2 #(
		.INIT('h1)
	) name14526 (
		_w24809_,
		_w24810_,
		_w25038_
	);
	LUT2 #(
		.INIT('h1)
	) name14527 (
		_w24811_,
		_w24812_,
		_w25039_
	);
	LUT2 #(
		.INIT('h1)
	) name14528 (
		_w24813_,
		_w24814_,
		_w25040_
	);
	LUT2 #(
		.INIT('h1)
	) name14529 (
		_w24815_,
		_w24816_,
		_w25041_
	);
	LUT2 #(
		.INIT('h1)
	) name14530 (
		_w24817_,
		_w24818_,
		_w25042_
	);
	LUT2 #(
		.INIT('h1)
	) name14531 (
		_w24819_,
		_w24820_,
		_w25043_
	);
	LUT2 #(
		.INIT('h1)
	) name14532 (
		_w24821_,
		_w24822_,
		_w25044_
	);
	LUT2 #(
		.INIT('h1)
	) name14533 (
		_w24823_,
		_w24824_,
		_w25045_
	);
	LUT2 #(
		.INIT('h1)
	) name14534 (
		_w24825_,
		_w24826_,
		_w25046_
	);
	LUT2 #(
		.INIT('h1)
	) name14535 (
		_w24827_,
		_w24828_,
		_w25047_
	);
	LUT2 #(
		.INIT('h1)
	) name14536 (
		_w24829_,
		_w24830_,
		_w25048_
	);
	LUT2 #(
		.INIT('h1)
	) name14537 (
		_w24831_,
		_w24832_,
		_w25049_
	);
	LUT2 #(
		.INIT('h1)
	) name14538 (
		_w24833_,
		_w24834_,
		_w25050_
	);
	LUT2 #(
		.INIT('h1)
	) name14539 (
		_w24835_,
		_w24836_,
		_w25051_
	);
	LUT2 #(
		.INIT('h1)
	) name14540 (
		_w24837_,
		_w24838_,
		_w25052_
	);
	LUT2 #(
		.INIT('h1)
	) name14541 (
		_w24839_,
		_w24840_,
		_w25053_
	);
	LUT2 #(
		.INIT('h1)
	) name14542 (
		_w24841_,
		_w24842_,
		_w25054_
	);
	LUT2 #(
		.INIT('h1)
	) name14543 (
		_w24843_,
		_w24844_,
		_w25055_
	);
	LUT2 #(
		.INIT('h1)
	) name14544 (
		_w24845_,
		_w24846_,
		_w25056_
	);
	LUT2 #(
		.INIT('h1)
	) name14545 (
		_w24847_,
		_w24848_,
		_w25057_
	);
	LUT2 #(
		.INIT('h1)
	) name14546 (
		_w24849_,
		_w24850_,
		_w25058_
	);
	LUT2 #(
		.INIT('h1)
	) name14547 (
		_w24851_,
		_w24852_,
		_w25059_
	);
	LUT2 #(
		.INIT('h1)
	) name14548 (
		_w24853_,
		_w24854_,
		_w25060_
	);
	LUT2 #(
		.INIT('h1)
	) name14549 (
		_w24855_,
		_w24856_,
		_w25061_
	);
	LUT2 #(
		.INIT('h1)
	) name14550 (
		_w24857_,
		_w24858_,
		_w25062_
	);
	LUT2 #(
		.INIT('h1)
	) name14551 (
		_w24859_,
		_w24860_,
		_w25063_
	);
	LUT2 #(
		.INIT('h1)
	) name14552 (
		_w24861_,
		_w24862_,
		_w25064_
	);
	LUT2 #(
		.INIT('h1)
	) name14553 (
		_w24863_,
		_w24864_,
		_w25065_
	);
	LUT2 #(
		.INIT('h1)
	) name14554 (
		_w24865_,
		_w24866_,
		_w25066_
	);
	LUT2 #(
		.INIT('h1)
	) name14555 (
		_w24867_,
		_w24868_,
		_w25067_
	);
	LUT2 #(
		.INIT('h1)
	) name14556 (
		_w24869_,
		_w24870_,
		_w25068_
	);
	LUT2 #(
		.INIT('h1)
	) name14557 (
		_w24871_,
		_w24872_,
		_w25069_
	);
	LUT2 #(
		.INIT('h1)
	) name14558 (
		_w24873_,
		_w24874_,
		_w25070_
	);
	LUT2 #(
		.INIT('h1)
	) name14559 (
		_w24875_,
		_w24876_,
		_w25071_
	);
	LUT2 #(
		.INIT('h1)
	) name14560 (
		_w24877_,
		_w24878_,
		_w25072_
	);
	LUT2 #(
		.INIT('h1)
	) name14561 (
		_w24879_,
		_w24880_,
		_w25073_
	);
	LUT2 #(
		.INIT('h1)
	) name14562 (
		_w24881_,
		_w24882_,
		_w25074_
	);
	LUT2 #(
		.INIT('h1)
	) name14563 (
		_w24883_,
		_w24884_,
		_w25075_
	);
	LUT2 #(
		.INIT('h1)
	) name14564 (
		_w24885_,
		_w24886_,
		_w25076_
	);
	LUT2 #(
		.INIT('h1)
	) name14565 (
		_w24887_,
		_w24888_,
		_w25077_
	);
	LUT2 #(
		.INIT('h1)
	) name14566 (
		_w24889_,
		_w24890_,
		_w25078_
	);
	LUT2 #(
		.INIT('h1)
	) name14567 (
		_w24891_,
		_w24892_,
		_w25079_
	);
	LUT2 #(
		.INIT('h1)
	) name14568 (
		_w24893_,
		_w24894_,
		_w25080_
	);
	LUT2 #(
		.INIT('h1)
	) name14569 (
		_w24895_,
		_w24896_,
		_w25081_
	);
	LUT2 #(
		.INIT('h1)
	) name14570 (
		_w24897_,
		_w24898_,
		_w25082_
	);
	LUT2 #(
		.INIT('h1)
	) name14571 (
		_w24899_,
		_w24900_,
		_w25083_
	);
	LUT2 #(
		.INIT('h1)
	) name14572 (
		_w24901_,
		_w24902_,
		_w25084_
	);
	LUT2 #(
		.INIT('h1)
	) name14573 (
		_w24903_,
		_w24904_,
		_w25085_
	);
	LUT2 #(
		.INIT('h1)
	) name14574 (
		_w24905_,
		_w24906_,
		_w25086_
	);
	LUT2 #(
		.INIT('h1)
	) name14575 (
		_w24907_,
		_w24908_,
		_w25087_
	);
	LUT2 #(
		.INIT('h1)
	) name14576 (
		_w24909_,
		_w24910_,
		_w25088_
	);
	LUT2 #(
		.INIT('h1)
	) name14577 (
		_w24911_,
		_w24912_,
		_w25089_
	);
	LUT2 #(
		.INIT('h1)
	) name14578 (
		_w24913_,
		_w24914_,
		_w25090_
	);
	LUT2 #(
		.INIT('h1)
	) name14579 (
		_w24915_,
		_w24916_,
		_w25091_
	);
	LUT2 #(
		.INIT('h1)
	) name14580 (
		_w24917_,
		_w24918_,
		_w25092_
	);
	LUT2 #(
		.INIT('h1)
	) name14581 (
		_w24919_,
		_w24920_,
		_w25093_
	);
	LUT2 #(
		.INIT('h1)
	) name14582 (
		_w24921_,
		_w24922_,
		_w25094_
	);
	LUT2 #(
		.INIT('h1)
	) name14583 (
		_w24923_,
		_w24924_,
		_w25095_
	);
	LUT2 #(
		.INIT('h1)
	) name14584 (
		_w24925_,
		_w24926_,
		_w25096_
	);
	LUT2 #(
		.INIT('h1)
	) name14585 (
		_w24927_,
		_w24928_,
		_w25097_
	);
	LUT2 #(
		.INIT('h1)
	) name14586 (
		_w24929_,
		_w24930_,
		_w25098_
	);
	LUT2 #(
		.INIT('h1)
	) name14587 (
		_w24931_,
		_w24932_,
		_w25099_
	);
	LUT2 #(
		.INIT('h1)
	) name14588 (
		_w24933_,
		_w24934_,
		_w25100_
	);
	LUT2 #(
		.INIT('h1)
	) name14589 (
		_w24935_,
		_w24936_,
		_w25101_
	);
	LUT2 #(
		.INIT('h1)
	) name14590 (
		_w24937_,
		_w24938_,
		_w25102_
	);
	LUT2 #(
		.INIT('h1)
	) name14591 (
		_w24939_,
		_w24940_,
		_w25103_
	);
	LUT2 #(
		.INIT('h1)
	) name14592 (
		_w24941_,
		_w24942_,
		_w25104_
	);
	LUT2 #(
		.INIT('h1)
	) name14593 (
		_w24943_,
		_w24944_,
		_w25105_
	);
	LUT2 #(
		.INIT('h1)
	) name14594 (
		_w24945_,
		_w24946_,
		_w25106_
	);
	LUT2 #(
		.INIT('h1)
	) name14595 (
		_w24947_,
		_w24948_,
		_w25107_
	);
	LUT2 #(
		.INIT('h1)
	) name14596 (
		_w24949_,
		_w24950_,
		_w25108_
	);
	LUT2 #(
		.INIT('h1)
	) name14597 (
		_w24951_,
		_w24952_,
		_w25109_
	);
	LUT2 #(
		.INIT('h1)
	) name14598 (
		_w24953_,
		_w24954_,
		_w25110_
	);
	LUT2 #(
		.INIT('h1)
	) name14599 (
		_w24955_,
		_w24956_,
		_w25111_
	);
	LUT2 #(
		.INIT('h1)
	) name14600 (
		_w24957_,
		_w24958_,
		_w25112_
	);
	LUT2 #(
		.INIT('h1)
	) name14601 (
		_w24959_,
		_w24960_,
		_w25113_
	);
	LUT2 #(
		.INIT('h1)
	) name14602 (
		_w24961_,
		_w24962_,
		_w25114_
	);
	LUT2 #(
		.INIT('h1)
	) name14603 (
		_w24963_,
		_w24964_,
		_w25115_
	);
	LUT2 #(
		.INIT('h1)
	) name14604 (
		_w24965_,
		_w24966_,
		_w25116_
	);
	LUT2 #(
		.INIT('h1)
	) name14605 (
		_w24967_,
		_w24968_,
		_w25117_
	);
	LUT2 #(
		.INIT('h1)
	) name14606 (
		_w24969_,
		_w24970_,
		_w25118_
	);
	LUT2 #(
		.INIT('h1)
	) name14607 (
		_w24971_,
		_w24972_,
		_w25119_
	);
	LUT2 #(
		.INIT('h1)
	) name14608 (
		_w24973_,
		_w24974_,
		_w25120_
	);
	LUT2 #(
		.INIT('h1)
	) name14609 (
		_w24975_,
		_w24976_,
		_w25121_
	);
	LUT2 #(
		.INIT('h1)
	) name14610 (
		_w24977_,
		_w24978_,
		_w25122_
	);
	LUT2 #(
		.INIT('h1)
	) name14611 (
		_w24979_,
		_w24980_,
		_w25123_
	);
	LUT2 #(
		.INIT('h1)
	) name14612 (
		_w24981_,
		_w24982_,
		_w25124_
	);
	LUT2 #(
		.INIT('h1)
	) name14613 (
		_w24983_,
		_w24984_,
		_w25125_
	);
	LUT2 #(
		.INIT('h1)
	) name14614 (
		_w24985_,
		_w24986_,
		_w25126_
	);
	LUT2 #(
		.INIT('h1)
	) name14615 (
		_w24987_,
		_w24988_,
		_w25127_
	);
	LUT2 #(
		.INIT('h1)
	) name14616 (
		_w24989_,
		_w24990_,
		_w25128_
	);
	LUT2 #(
		.INIT('h1)
	) name14617 (
		_w24991_,
		_w24992_,
		_w25129_
	);
	LUT2 #(
		.INIT('h1)
	) name14618 (
		_w24993_,
		_w24994_,
		_w25130_
	);
	LUT2 #(
		.INIT('h1)
	) name14619 (
		_w24995_,
		_w24996_,
		_w25131_
	);
	LUT2 #(
		.INIT('h1)
	) name14620 (
		_w24997_,
		_w24998_,
		_w25132_
	);
	LUT2 #(
		.INIT('h1)
	) name14621 (
		_w24999_,
		_w25000_,
		_w25133_
	);
	LUT2 #(
		.INIT('h1)
	) name14622 (
		_w25001_,
		_w25002_,
		_w25134_
	);
	LUT2 #(
		.INIT('h1)
	) name14623 (
		_w25003_,
		_w25004_,
		_w25135_
	);
	LUT2 #(
		.INIT('h1)
	) name14624 (
		_w25005_,
		_w25006_,
		_w25136_
	);
	LUT2 #(
		.INIT('h1)
	) name14625 (
		_w25007_,
		_w25008_,
		_w25137_
	);
	LUT2 #(
		.INIT('h1)
	) name14626 (
		_w25009_,
		_w25010_,
		_w25138_
	);
	LUT2 #(
		.INIT('h8)
	) name14627 (
		_w25137_,
		_w25138_,
		_w25139_
	);
	LUT2 #(
		.INIT('h8)
	) name14628 (
		_w25135_,
		_w25136_,
		_w25140_
	);
	LUT2 #(
		.INIT('h8)
	) name14629 (
		_w25133_,
		_w25134_,
		_w25141_
	);
	LUT2 #(
		.INIT('h8)
	) name14630 (
		_w25131_,
		_w25132_,
		_w25142_
	);
	LUT2 #(
		.INIT('h8)
	) name14631 (
		_w25129_,
		_w25130_,
		_w25143_
	);
	LUT2 #(
		.INIT('h8)
	) name14632 (
		_w25127_,
		_w25128_,
		_w25144_
	);
	LUT2 #(
		.INIT('h8)
	) name14633 (
		_w25125_,
		_w25126_,
		_w25145_
	);
	LUT2 #(
		.INIT('h8)
	) name14634 (
		_w25123_,
		_w25124_,
		_w25146_
	);
	LUT2 #(
		.INIT('h8)
	) name14635 (
		_w25121_,
		_w25122_,
		_w25147_
	);
	LUT2 #(
		.INIT('h8)
	) name14636 (
		_w25119_,
		_w25120_,
		_w25148_
	);
	LUT2 #(
		.INIT('h8)
	) name14637 (
		_w25117_,
		_w25118_,
		_w25149_
	);
	LUT2 #(
		.INIT('h8)
	) name14638 (
		_w25115_,
		_w25116_,
		_w25150_
	);
	LUT2 #(
		.INIT('h8)
	) name14639 (
		_w25113_,
		_w25114_,
		_w25151_
	);
	LUT2 #(
		.INIT('h8)
	) name14640 (
		_w25111_,
		_w25112_,
		_w25152_
	);
	LUT2 #(
		.INIT('h8)
	) name14641 (
		_w25109_,
		_w25110_,
		_w25153_
	);
	LUT2 #(
		.INIT('h8)
	) name14642 (
		_w25107_,
		_w25108_,
		_w25154_
	);
	LUT2 #(
		.INIT('h8)
	) name14643 (
		_w25105_,
		_w25106_,
		_w25155_
	);
	LUT2 #(
		.INIT('h8)
	) name14644 (
		_w25103_,
		_w25104_,
		_w25156_
	);
	LUT2 #(
		.INIT('h8)
	) name14645 (
		_w25101_,
		_w25102_,
		_w25157_
	);
	LUT2 #(
		.INIT('h8)
	) name14646 (
		_w25099_,
		_w25100_,
		_w25158_
	);
	LUT2 #(
		.INIT('h8)
	) name14647 (
		_w25097_,
		_w25098_,
		_w25159_
	);
	LUT2 #(
		.INIT('h8)
	) name14648 (
		_w25095_,
		_w25096_,
		_w25160_
	);
	LUT2 #(
		.INIT('h8)
	) name14649 (
		_w25093_,
		_w25094_,
		_w25161_
	);
	LUT2 #(
		.INIT('h8)
	) name14650 (
		_w25091_,
		_w25092_,
		_w25162_
	);
	LUT2 #(
		.INIT('h8)
	) name14651 (
		_w25089_,
		_w25090_,
		_w25163_
	);
	LUT2 #(
		.INIT('h8)
	) name14652 (
		_w25087_,
		_w25088_,
		_w25164_
	);
	LUT2 #(
		.INIT('h8)
	) name14653 (
		_w25085_,
		_w25086_,
		_w25165_
	);
	LUT2 #(
		.INIT('h8)
	) name14654 (
		_w25083_,
		_w25084_,
		_w25166_
	);
	LUT2 #(
		.INIT('h8)
	) name14655 (
		_w25081_,
		_w25082_,
		_w25167_
	);
	LUT2 #(
		.INIT('h8)
	) name14656 (
		_w25079_,
		_w25080_,
		_w25168_
	);
	LUT2 #(
		.INIT('h8)
	) name14657 (
		_w25077_,
		_w25078_,
		_w25169_
	);
	LUT2 #(
		.INIT('h8)
	) name14658 (
		_w25075_,
		_w25076_,
		_w25170_
	);
	LUT2 #(
		.INIT('h8)
	) name14659 (
		_w25073_,
		_w25074_,
		_w25171_
	);
	LUT2 #(
		.INIT('h8)
	) name14660 (
		_w25071_,
		_w25072_,
		_w25172_
	);
	LUT2 #(
		.INIT('h8)
	) name14661 (
		_w25069_,
		_w25070_,
		_w25173_
	);
	LUT2 #(
		.INIT('h8)
	) name14662 (
		_w25067_,
		_w25068_,
		_w25174_
	);
	LUT2 #(
		.INIT('h8)
	) name14663 (
		_w25065_,
		_w25066_,
		_w25175_
	);
	LUT2 #(
		.INIT('h8)
	) name14664 (
		_w25063_,
		_w25064_,
		_w25176_
	);
	LUT2 #(
		.INIT('h8)
	) name14665 (
		_w25061_,
		_w25062_,
		_w25177_
	);
	LUT2 #(
		.INIT('h8)
	) name14666 (
		_w25059_,
		_w25060_,
		_w25178_
	);
	LUT2 #(
		.INIT('h8)
	) name14667 (
		_w25057_,
		_w25058_,
		_w25179_
	);
	LUT2 #(
		.INIT('h8)
	) name14668 (
		_w25055_,
		_w25056_,
		_w25180_
	);
	LUT2 #(
		.INIT('h8)
	) name14669 (
		_w25053_,
		_w25054_,
		_w25181_
	);
	LUT2 #(
		.INIT('h8)
	) name14670 (
		_w25051_,
		_w25052_,
		_w25182_
	);
	LUT2 #(
		.INIT('h8)
	) name14671 (
		_w25049_,
		_w25050_,
		_w25183_
	);
	LUT2 #(
		.INIT('h8)
	) name14672 (
		_w25047_,
		_w25048_,
		_w25184_
	);
	LUT2 #(
		.INIT('h8)
	) name14673 (
		_w25045_,
		_w25046_,
		_w25185_
	);
	LUT2 #(
		.INIT('h8)
	) name14674 (
		_w25043_,
		_w25044_,
		_w25186_
	);
	LUT2 #(
		.INIT('h8)
	) name14675 (
		_w25041_,
		_w25042_,
		_w25187_
	);
	LUT2 #(
		.INIT('h8)
	) name14676 (
		_w25039_,
		_w25040_,
		_w25188_
	);
	LUT2 #(
		.INIT('h8)
	) name14677 (
		_w25037_,
		_w25038_,
		_w25189_
	);
	LUT2 #(
		.INIT('h8)
	) name14678 (
		_w25035_,
		_w25036_,
		_w25190_
	);
	LUT2 #(
		.INIT('h8)
	) name14679 (
		_w25033_,
		_w25034_,
		_w25191_
	);
	LUT2 #(
		.INIT('h8)
	) name14680 (
		_w25031_,
		_w25032_,
		_w25192_
	);
	LUT2 #(
		.INIT('h8)
	) name14681 (
		_w25029_,
		_w25030_,
		_w25193_
	);
	LUT2 #(
		.INIT('h8)
	) name14682 (
		_w25027_,
		_w25028_,
		_w25194_
	);
	LUT2 #(
		.INIT('h8)
	) name14683 (
		_w25025_,
		_w25026_,
		_w25195_
	);
	LUT2 #(
		.INIT('h8)
	) name14684 (
		_w25023_,
		_w25024_,
		_w25196_
	);
	LUT2 #(
		.INIT('h8)
	) name14685 (
		_w25021_,
		_w25022_,
		_w25197_
	);
	LUT2 #(
		.INIT('h8)
	) name14686 (
		_w25019_,
		_w25020_,
		_w25198_
	);
	LUT2 #(
		.INIT('h8)
	) name14687 (
		_w25017_,
		_w25018_,
		_w25199_
	);
	LUT2 #(
		.INIT('h8)
	) name14688 (
		_w25015_,
		_w25016_,
		_w25200_
	);
	LUT2 #(
		.INIT('h8)
	) name14689 (
		_w25013_,
		_w25014_,
		_w25201_
	);
	LUT2 #(
		.INIT('h8)
	) name14690 (
		_w25011_,
		_w25012_,
		_w25202_
	);
	LUT2 #(
		.INIT('h8)
	) name14691 (
		_w25201_,
		_w25202_,
		_w25203_
	);
	LUT2 #(
		.INIT('h8)
	) name14692 (
		_w25199_,
		_w25200_,
		_w25204_
	);
	LUT2 #(
		.INIT('h8)
	) name14693 (
		_w25197_,
		_w25198_,
		_w25205_
	);
	LUT2 #(
		.INIT('h8)
	) name14694 (
		_w25195_,
		_w25196_,
		_w25206_
	);
	LUT2 #(
		.INIT('h8)
	) name14695 (
		_w25193_,
		_w25194_,
		_w25207_
	);
	LUT2 #(
		.INIT('h8)
	) name14696 (
		_w25191_,
		_w25192_,
		_w25208_
	);
	LUT2 #(
		.INIT('h8)
	) name14697 (
		_w25189_,
		_w25190_,
		_w25209_
	);
	LUT2 #(
		.INIT('h8)
	) name14698 (
		_w25187_,
		_w25188_,
		_w25210_
	);
	LUT2 #(
		.INIT('h8)
	) name14699 (
		_w25185_,
		_w25186_,
		_w25211_
	);
	LUT2 #(
		.INIT('h8)
	) name14700 (
		_w25183_,
		_w25184_,
		_w25212_
	);
	LUT2 #(
		.INIT('h8)
	) name14701 (
		_w25181_,
		_w25182_,
		_w25213_
	);
	LUT2 #(
		.INIT('h8)
	) name14702 (
		_w25179_,
		_w25180_,
		_w25214_
	);
	LUT2 #(
		.INIT('h8)
	) name14703 (
		_w25177_,
		_w25178_,
		_w25215_
	);
	LUT2 #(
		.INIT('h8)
	) name14704 (
		_w25175_,
		_w25176_,
		_w25216_
	);
	LUT2 #(
		.INIT('h8)
	) name14705 (
		_w25173_,
		_w25174_,
		_w25217_
	);
	LUT2 #(
		.INIT('h8)
	) name14706 (
		_w25171_,
		_w25172_,
		_w25218_
	);
	LUT2 #(
		.INIT('h8)
	) name14707 (
		_w25169_,
		_w25170_,
		_w25219_
	);
	LUT2 #(
		.INIT('h8)
	) name14708 (
		_w25167_,
		_w25168_,
		_w25220_
	);
	LUT2 #(
		.INIT('h8)
	) name14709 (
		_w25165_,
		_w25166_,
		_w25221_
	);
	LUT2 #(
		.INIT('h8)
	) name14710 (
		_w25163_,
		_w25164_,
		_w25222_
	);
	LUT2 #(
		.INIT('h8)
	) name14711 (
		_w25161_,
		_w25162_,
		_w25223_
	);
	LUT2 #(
		.INIT('h8)
	) name14712 (
		_w25159_,
		_w25160_,
		_w25224_
	);
	LUT2 #(
		.INIT('h8)
	) name14713 (
		_w25157_,
		_w25158_,
		_w25225_
	);
	LUT2 #(
		.INIT('h8)
	) name14714 (
		_w25155_,
		_w25156_,
		_w25226_
	);
	LUT2 #(
		.INIT('h8)
	) name14715 (
		_w25153_,
		_w25154_,
		_w25227_
	);
	LUT2 #(
		.INIT('h8)
	) name14716 (
		_w25151_,
		_w25152_,
		_w25228_
	);
	LUT2 #(
		.INIT('h8)
	) name14717 (
		_w25149_,
		_w25150_,
		_w25229_
	);
	LUT2 #(
		.INIT('h8)
	) name14718 (
		_w25147_,
		_w25148_,
		_w25230_
	);
	LUT2 #(
		.INIT('h8)
	) name14719 (
		_w25145_,
		_w25146_,
		_w25231_
	);
	LUT2 #(
		.INIT('h8)
	) name14720 (
		_w25143_,
		_w25144_,
		_w25232_
	);
	LUT2 #(
		.INIT('h8)
	) name14721 (
		_w25141_,
		_w25142_,
		_w25233_
	);
	LUT2 #(
		.INIT('h8)
	) name14722 (
		_w25139_,
		_w25140_,
		_w25234_
	);
	LUT2 #(
		.INIT('h8)
	) name14723 (
		_w25233_,
		_w25234_,
		_w25235_
	);
	LUT2 #(
		.INIT('h8)
	) name14724 (
		_w25231_,
		_w25232_,
		_w25236_
	);
	LUT2 #(
		.INIT('h8)
	) name14725 (
		_w25229_,
		_w25230_,
		_w25237_
	);
	LUT2 #(
		.INIT('h8)
	) name14726 (
		_w25227_,
		_w25228_,
		_w25238_
	);
	LUT2 #(
		.INIT('h8)
	) name14727 (
		_w25225_,
		_w25226_,
		_w25239_
	);
	LUT2 #(
		.INIT('h8)
	) name14728 (
		_w25223_,
		_w25224_,
		_w25240_
	);
	LUT2 #(
		.INIT('h8)
	) name14729 (
		_w25221_,
		_w25222_,
		_w25241_
	);
	LUT2 #(
		.INIT('h8)
	) name14730 (
		_w25219_,
		_w25220_,
		_w25242_
	);
	LUT2 #(
		.INIT('h8)
	) name14731 (
		_w25217_,
		_w25218_,
		_w25243_
	);
	LUT2 #(
		.INIT('h8)
	) name14732 (
		_w25215_,
		_w25216_,
		_w25244_
	);
	LUT2 #(
		.INIT('h8)
	) name14733 (
		_w25213_,
		_w25214_,
		_w25245_
	);
	LUT2 #(
		.INIT('h8)
	) name14734 (
		_w25211_,
		_w25212_,
		_w25246_
	);
	LUT2 #(
		.INIT('h8)
	) name14735 (
		_w25209_,
		_w25210_,
		_w25247_
	);
	LUT2 #(
		.INIT('h8)
	) name14736 (
		_w25207_,
		_w25208_,
		_w25248_
	);
	LUT2 #(
		.INIT('h8)
	) name14737 (
		_w25205_,
		_w25206_,
		_w25249_
	);
	LUT2 #(
		.INIT('h8)
	) name14738 (
		_w25203_,
		_w25204_,
		_w25250_
	);
	LUT2 #(
		.INIT('h8)
	) name14739 (
		_w25249_,
		_w25250_,
		_w25251_
	);
	LUT2 #(
		.INIT('h8)
	) name14740 (
		_w25247_,
		_w25248_,
		_w25252_
	);
	LUT2 #(
		.INIT('h8)
	) name14741 (
		_w25245_,
		_w25246_,
		_w25253_
	);
	LUT2 #(
		.INIT('h8)
	) name14742 (
		_w25243_,
		_w25244_,
		_w25254_
	);
	LUT2 #(
		.INIT('h8)
	) name14743 (
		_w25241_,
		_w25242_,
		_w25255_
	);
	LUT2 #(
		.INIT('h8)
	) name14744 (
		_w25239_,
		_w25240_,
		_w25256_
	);
	LUT2 #(
		.INIT('h8)
	) name14745 (
		_w25237_,
		_w25238_,
		_w25257_
	);
	LUT2 #(
		.INIT('h8)
	) name14746 (
		_w25235_,
		_w25236_,
		_w25258_
	);
	LUT2 #(
		.INIT('h8)
	) name14747 (
		_w25257_,
		_w25258_,
		_w25259_
	);
	LUT2 #(
		.INIT('h8)
	) name14748 (
		_w25255_,
		_w25256_,
		_w25260_
	);
	LUT2 #(
		.INIT('h8)
	) name14749 (
		_w25253_,
		_w25254_,
		_w25261_
	);
	LUT2 #(
		.INIT('h8)
	) name14750 (
		_w25251_,
		_w25252_,
		_w25262_
	);
	LUT2 #(
		.INIT('h8)
	) name14751 (
		_w25261_,
		_w25262_,
		_w25263_
	);
	LUT2 #(
		.INIT('h8)
	) name14752 (
		_w25259_,
		_w25260_,
		_w25264_
	);
	LUT2 #(
		.INIT('h8)
	) name14753 (
		_w25263_,
		_w25264_,
		_w25265_
	);
	LUT2 #(
		.INIT('h1)
	) name14754 (
		wb_rst_i_pad,
		_w25265_,
		_w25266_
	);
	LUT2 #(
		.INIT('h1)
	) name14755 (
		_w22944_,
		_w25266_,
		_w25267_
	);
	LUT2 #(
		.INIT('h8)
	) name14756 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 ,
		_w23522_,
		_w25268_
	);
	LUT2 #(
		.INIT('h8)
	) name14757 (
		\ethreg1_IPGR1_0_DataOut_reg[4]/NET0131 ,
		_w24710_,
		_w25269_
	);
	LUT2 #(
		.INIT('h8)
	) name14758 (
		\ethreg1_IPGT_0_DataOut_reg[4]/NET0131 ,
		_w24717_,
		_w25270_
	);
	LUT2 #(
		.INIT('h8)
	) name14759 (
		\ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 ,
		_w24722_,
		_w25271_
	);
	LUT2 #(
		.INIT('h8)
	) name14760 (
		\ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 ,
		_w23499_,
		_w25272_
	);
	LUT2 #(
		.INIT('h8)
	) name14761 (
		\ethreg1_PACKETLEN_0_DataOut_reg[4]/NET0131 ,
		_w22966_,
		_w25273_
	);
	LUT2 #(
		.INIT('h8)
	) name14762 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		_w24726_,
		_w25274_
	);
	LUT2 #(
		.INIT('h8)
	) name14763 (
		\ethreg1_irq_busy_reg/NET0131 ,
		_w24707_,
		_w25275_
	);
	LUT2 #(
		.INIT('h8)
	) name14764 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 ,
		_w23513_,
		_w25276_
	);
	LUT2 #(
		.INIT('h8)
	) name14765 (
		\ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 ,
		_w22956_,
		_w25277_
	);
	LUT2 #(
		.INIT('h8)
	) name14766 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		_w22959_,
		_w25278_
	);
	LUT2 #(
		.INIT('h8)
	) name14767 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		_w23501_,
		_w25279_
	);
	LUT2 #(
		.INIT('h8)
	) name14768 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		_w24713_,
		_w25280_
	);
	LUT2 #(
		.INIT('h8)
	) name14769 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		_w24730_,
		_w25281_
	);
	LUT2 #(
		.INIT('h8)
	) name14770 (
		\ethreg1_IPGR2_0_DataOut_reg[4]/NET0131 ,
		_w24724_,
		_w25282_
	);
	LUT2 #(
		.INIT('h8)
	) name14771 (
		\ethreg1_MIIRX_DATA_DataOut_reg[4]/NET0131 ,
		_w23507_,
		_w25283_
	);
	LUT2 #(
		.INIT('h8)
	) name14772 (
		\ethreg1_MODER_0_DataOut_reg[4]/NET0131 ,
		_w23519_,
		_w25284_
	);
	LUT2 #(
		.INIT('h8)
	) name14773 (
		\ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 ,
		_w22952_,
		_w25285_
	);
	LUT2 #(
		.INIT('h1)
	) name14774 (
		_w25268_,
		_w25269_,
		_w25286_
	);
	LUT2 #(
		.INIT('h1)
	) name14775 (
		_w25270_,
		_w25271_,
		_w25287_
	);
	LUT2 #(
		.INIT('h1)
	) name14776 (
		_w25272_,
		_w25274_,
		_w25288_
	);
	LUT2 #(
		.INIT('h1)
	) name14777 (
		_w25275_,
		_w25276_,
		_w25289_
	);
	LUT2 #(
		.INIT('h1)
	) name14778 (
		_w25277_,
		_w25278_,
		_w25290_
	);
	LUT2 #(
		.INIT('h1)
	) name14779 (
		_w25279_,
		_w25280_,
		_w25291_
	);
	LUT2 #(
		.INIT('h1)
	) name14780 (
		_w25282_,
		_w25283_,
		_w25292_
	);
	LUT2 #(
		.INIT('h1)
	) name14781 (
		_w25284_,
		_w25285_,
		_w25293_
	);
	LUT2 #(
		.INIT('h8)
	) name14782 (
		_w25292_,
		_w25293_,
		_w25294_
	);
	LUT2 #(
		.INIT('h8)
	) name14783 (
		_w25290_,
		_w25291_,
		_w25295_
	);
	LUT2 #(
		.INIT('h8)
	) name14784 (
		_w25288_,
		_w25289_,
		_w25296_
	);
	LUT2 #(
		.INIT('h8)
	) name14785 (
		_w25286_,
		_w25287_,
		_w25297_
	);
	LUT2 #(
		.INIT('h8)
	) name14786 (
		_w22944_,
		_w25297_,
		_w25298_
	);
	LUT2 #(
		.INIT('h8)
	) name14787 (
		_w25295_,
		_w25296_,
		_w25299_
	);
	LUT2 #(
		.INIT('h4)
	) name14788 (
		_w25273_,
		_w25294_,
		_w25300_
	);
	LUT2 #(
		.INIT('h4)
	) name14789 (
		_w25281_,
		_w25300_,
		_w25301_
	);
	LUT2 #(
		.INIT('h8)
	) name14790 (
		_w25298_,
		_w25299_,
		_w25302_
	);
	LUT2 #(
		.INIT('h8)
	) name14791 (
		_w25301_,
		_w25302_,
		_w25303_
	);
	LUT2 #(
		.INIT('h1)
	) name14792 (
		_w25267_,
		_w25303_,
		_w25304_
	);
	LUT2 #(
		.INIT('h8)
	) name14793 (
		\wishbone_bd_ram_mem0_reg[30][5]/P0001 ,
		_w13104_,
		_w25305_
	);
	LUT2 #(
		.INIT('h8)
	) name14794 (
		\wishbone_bd_ram_mem0_reg[60][5]/P0001 ,
		_w13204_,
		_w25306_
	);
	LUT2 #(
		.INIT('h8)
	) name14795 (
		\wishbone_bd_ram_mem0_reg[33][5]/P0001 ,
		_w12980_,
		_w25307_
	);
	LUT2 #(
		.INIT('h8)
	) name14796 (
		\wishbone_bd_ram_mem0_reg[95][5]/P0001 ,
		_w12844_,
		_w25308_
	);
	LUT2 #(
		.INIT('h8)
	) name14797 (
		\wishbone_bd_ram_mem0_reg[61][5]/P0001 ,
		_w12725_,
		_w25309_
	);
	LUT2 #(
		.INIT('h8)
	) name14798 (
		\wishbone_bd_ram_mem0_reg[200][5]/P0001 ,
		_w12988_,
		_w25310_
	);
	LUT2 #(
		.INIT('h8)
	) name14799 (
		\wishbone_bd_ram_mem0_reg[149][5]/P0001 ,
		_w12741_,
		_w25311_
	);
	LUT2 #(
		.INIT('h8)
	) name14800 (
		\wishbone_bd_ram_mem0_reg[32][5]/P0001 ,
		_w13120_,
		_w25312_
	);
	LUT2 #(
		.INIT('h8)
	) name14801 (
		\wishbone_bd_ram_mem0_reg[166][5]/P0001 ,
		_w13040_,
		_w25313_
	);
	LUT2 #(
		.INIT('h8)
	) name14802 (
		\wishbone_bd_ram_mem0_reg[246][5]/P0001 ,
		_w13076_,
		_w25314_
	);
	LUT2 #(
		.INIT('h8)
	) name14803 (
		\wishbone_bd_ram_mem0_reg[175][5]/P0001 ,
		_w13126_,
		_w25315_
	);
	LUT2 #(
		.INIT('h8)
	) name14804 (
		\wishbone_bd_ram_mem0_reg[150][5]/P0001 ,
		_w13136_,
		_w25316_
	);
	LUT2 #(
		.INIT('h8)
	) name14805 (
		\wishbone_bd_ram_mem0_reg[50][5]/P0001 ,
		_w13150_,
		_w25317_
	);
	LUT2 #(
		.INIT('h8)
	) name14806 (
		\wishbone_bd_ram_mem0_reg[94][5]/P0001 ,
		_w13186_,
		_w25318_
	);
	LUT2 #(
		.INIT('h8)
	) name14807 (
		\wishbone_bd_ram_mem0_reg[39][5]/P0001 ,
		_w13018_,
		_w25319_
	);
	LUT2 #(
		.INIT('h8)
	) name14808 (
		\wishbone_bd_ram_mem0_reg[51][5]/P0001 ,
		_w13024_,
		_w25320_
	);
	LUT2 #(
		.INIT('h8)
	) name14809 (
		\wishbone_bd_ram_mem0_reg[127][5]/P0001 ,
		_w13164_,
		_w25321_
	);
	LUT2 #(
		.INIT('h8)
	) name14810 (
		\wishbone_bd_ram_mem0_reg[232][5]/P0001 ,
		_w12758_,
		_w25322_
	);
	LUT2 #(
		.INIT('h8)
	) name14811 (
		\wishbone_bd_ram_mem0_reg[56][5]/P0001 ,
		_w12778_,
		_w25323_
	);
	LUT2 #(
		.INIT('h8)
	) name14812 (
		\wishbone_bd_ram_mem0_reg[1][5]/P0001 ,
		_w13014_,
		_w25324_
	);
	LUT2 #(
		.INIT('h8)
	) name14813 (
		\wishbone_bd_ram_mem0_reg[57][5]/P0001 ,
		_w13116_,
		_w25325_
	);
	LUT2 #(
		.INIT('h8)
	) name14814 (
		\wishbone_bd_ram_mem0_reg[198][5]/P0001 ,
		_w12832_,
		_w25326_
	);
	LUT2 #(
		.INIT('h8)
	) name14815 (
		\wishbone_bd_ram_mem0_reg[242][5]/P0001 ,
		_w12932_,
		_w25327_
	);
	LUT2 #(
		.INIT('h8)
	) name14816 (
		\wishbone_bd_ram_mem0_reg[180][5]/P0001 ,
		_w12791_,
		_w25328_
	);
	LUT2 #(
		.INIT('h8)
	) name14817 (
		\wishbone_bd_ram_mem0_reg[91][5]/P0001 ,
		_w13074_,
		_w25329_
	);
	LUT2 #(
		.INIT('h8)
	) name14818 (
		\wishbone_bd_ram_mem0_reg[49][5]/P0001 ,
		_w12994_,
		_w25330_
	);
	LUT2 #(
		.INIT('h8)
	) name14819 (
		\wishbone_bd_ram_mem0_reg[98][5]/P0001 ,
		_w12816_,
		_w25331_
	);
	LUT2 #(
		.INIT('h8)
	) name14820 (
		\wishbone_bd_ram_mem0_reg[105][5]/P0001 ,
		_w12751_,
		_w25332_
	);
	LUT2 #(
		.INIT('h8)
	) name14821 (
		\wishbone_bd_ram_mem0_reg[237][5]/P0001 ,
		_w12990_,
		_w25333_
	);
	LUT2 #(
		.INIT('h8)
	) name14822 (
		\wishbone_bd_ram_mem0_reg[100][5]/P0001 ,
		_w12960_,
		_w25334_
	);
	LUT2 #(
		.INIT('h8)
	) name14823 (
		\wishbone_bd_ram_mem0_reg[154][5]/P0001 ,
		_w12962_,
		_w25335_
	);
	LUT2 #(
		.INIT('h8)
	) name14824 (
		\wishbone_bd_ram_mem0_reg[173][5]/P0001 ,
		_w12854_,
		_w25336_
	);
	LUT2 #(
		.INIT('h8)
	) name14825 (
		\wishbone_bd_ram_mem0_reg[123][5]/P0001 ,
		_w13114_,
		_w25337_
	);
	LUT2 #(
		.INIT('h8)
	) name14826 (
		\wishbone_bd_ram_mem0_reg[181][5]/P0001 ,
		_w12828_,
		_w25338_
	);
	LUT2 #(
		.INIT('h8)
	) name14827 (
		\wishbone_bd_ram_mem0_reg[28][5]/P0001 ,
		_w13170_,
		_w25339_
	);
	LUT2 #(
		.INIT('h8)
	) name14828 (
		\wishbone_bd_ram_mem0_reg[218][5]/P0001 ,
		_w13206_,
		_w25340_
	);
	LUT2 #(
		.INIT('h8)
	) name14829 (
		\wishbone_bd_ram_mem0_reg[64][5]/P0001 ,
		_w12976_,
		_w25341_
	);
	LUT2 #(
		.INIT('h8)
	) name14830 (
		\wishbone_bd_ram_mem0_reg[71][5]/P0001 ,
		_w12798_,
		_w25342_
	);
	LUT2 #(
		.INIT('h8)
	) name14831 (
		\wishbone_bd_ram_mem0_reg[195][5]/P0001 ,
		_w13144_,
		_w25343_
	);
	LUT2 #(
		.INIT('h8)
	) name14832 (
		\wishbone_bd_ram_mem0_reg[41][5]/P0001 ,
		_w13052_,
		_w25344_
	);
	LUT2 #(
		.INIT('h8)
	) name14833 (
		\wishbone_bd_ram_mem0_reg[211][5]/P0001 ,
		_w13166_,
		_w25345_
	);
	LUT2 #(
		.INIT('h8)
	) name14834 (
		\wishbone_bd_ram_mem0_reg[189][5]/P0001 ,
		_w13042_,
		_w25346_
	);
	LUT2 #(
		.INIT('h8)
	) name14835 (
		\wishbone_bd_ram_mem0_reg[146][5]/P0001 ,
		_w13060_,
		_w25347_
	);
	LUT2 #(
		.INIT('h8)
	) name14836 (
		\wishbone_bd_ram_mem0_reg[157][5]/P0001 ,
		_w12926_,
		_w25348_
	);
	LUT2 #(
		.INIT('h8)
	) name14837 (
		\wishbone_bd_ram_mem0_reg[247][5]/P0001 ,
		_w12818_,
		_w25349_
	);
	LUT2 #(
		.INIT('h8)
	) name14838 (
		\wishbone_bd_ram_mem0_reg[197][5]/P0001 ,
		_w12834_,
		_w25350_
	);
	LUT2 #(
		.INIT('h8)
	) name14839 (
		\wishbone_bd_ram_mem0_reg[55][5]/P0001 ,
		_w12785_,
		_w25351_
	);
	LUT2 #(
		.INIT('h8)
	) name14840 (
		\wishbone_bd_ram_mem0_reg[194][5]/P0001 ,
		_w12772_,
		_w25352_
	);
	LUT2 #(
		.INIT('h8)
	) name14841 (
		\wishbone_bd_ram_mem0_reg[106][5]/P0001 ,
		_w12713_,
		_w25353_
	);
	LUT2 #(
		.INIT('h8)
	) name14842 (
		\wishbone_bd_ram_mem0_reg[215][5]/P0001 ,
		_w12974_,
		_w25354_
	);
	LUT2 #(
		.INIT('h8)
	) name14843 (
		\wishbone_bd_ram_mem0_reg[12][5]/P0001 ,
		_w13118_,
		_w25355_
	);
	LUT2 #(
		.INIT('h8)
	) name14844 (
		\wishbone_bd_ram_mem0_reg[118][5]/P0001 ,
		_w12830_,
		_w25356_
	);
	LUT2 #(
		.INIT('h8)
	) name14845 (
		\wishbone_bd_ram_mem0_reg[14][5]/P0001 ,
		_w13086_,
		_w25357_
	);
	LUT2 #(
		.INIT('h8)
	) name14846 (
		\wishbone_bd_ram_mem0_reg[169][5]/P0001 ,
		_w12722_,
		_w25358_
	);
	LUT2 #(
		.INIT('h8)
	) name14847 (
		\wishbone_bd_ram_mem0_reg[143][5]/P0001 ,
		_w12922_,
		_w25359_
	);
	LUT2 #(
		.INIT('h8)
	) name14848 (
		\wishbone_bd_ram_mem0_reg[185][5]/P0001 ,
		_w12940_,
		_w25360_
	);
	LUT2 #(
		.INIT('h8)
	) name14849 (
		\wishbone_bd_ram_mem0_reg[120][5]/P0001 ,
		_w12707_,
		_w25361_
	);
	LUT2 #(
		.INIT('h8)
	) name14850 (
		\wishbone_bd_ram_mem0_reg[239][5]/P0001 ,
		_w12862_,
		_w25362_
	);
	LUT2 #(
		.INIT('h8)
	) name14851 (
		\wishbone_bd_ram_mem0_reg[116][5]/P0001 ,
		_w12998_,
		_w25363_
	);
	LUT2 #(
		.INIT('h8)
	) name14852 (
		\wishbone_bd_ram_mem0_reg[122][5]/P0001 ,
		_w13130_,
		_w25364_
	);
	LUT2 #(
		.INIT('h8)
	) name14853 (
		\wishbone_bd_ram_mem0_reg[15][5]/P0001 ,
		_w13210_,
		_w25365_
	);
	LUT2 #(
		.INIT('h8)
	) name14854 (
		\wishbone_bd_ram_mem0_reg[131][5]/P0001 ,
		_w12852_,
		_w25366_
	);
	LUT2 #(
		.INIT('h8)
	) name14855 (
		\wishbone_bd_ram_mem0_reg[172][5]/P0001 ,
		_w12944_,
		_w25367_
	);
	LUT2 #(
		.INIT('h8)
	) name14856 (
		\wishbone_bd_ram_mem0_reg[209][5]/P0001 ,
		_w13152_,
		_w25368_
	);
	LUT2 #(
		.INIT('h8)
	) name14857 (
		\wishbone_bd_ram_mem0_reg[201][5]/P0001 ,
		_w12822_,
		_w25369_
	);
	LUT2 #(
		.INIT('h8)
	) name14858 (
		\wishbone_bd_ram_mem0_reg[183][5]/P0001 ,
		_w12787_,
		_w25370_
	);
	LUT2 #(
		.INIT('h8)
	) name14859 (
		\wishbone_bd_ram_mem0_reg[76][5]/P0001 ,
		_w13184_,
		_w25371_
	);
	LUT2 #(
		.INIT('h8)
	) name14860 (
		\wishbone_bd_ram_mem0_reg[43][5]/P0001 ,
		_w13200_,
		_w25372_
	);
	LUT2 #(
		.INIT('h8)
	) name14861 (
		\wishbone_bd_ram_mem0_reg[23][5]/P0001 ,
		_w13008_,
		_w25373_
	);
	LUT2 #(
		.INIT('h8)
	) name14862 (
		\wishbone_bd_ram_mem0_reg[145][5]/P0001 ,
		_w13106_,
		_w25374_
	);
	LUT2 #(
		.INIT('h8)
	) name14863 (
		\wishbone_bd_ram_mem0_reg[44][5]/P0001 ,
		_w12896_,
		_w25375_
	);
	LUT2 #(
		.INIT('h8)
	) name14864 (
		\wishbone_bd_ram_mem0_reg[136][5]/P0001 ,
		_w13064_,
		_w25376_
	);
	LUT2 #(
		.INIT('h8)
	) name14865 (
		\wishbone_bd_ram_mem0_reg[13][5]/P0001 ,
		_w13178_,
		_w25377_
	);
	LUT2 #(
		.INIT('h8)
	) name14866 (
		\wishbone_bd_ram_mem0_reg[74][5]/P0001 ,
		_w12812_,
		_w25378_
	);
	LUT2 #(
		.INIT('h8)
	) name14867 (
		\wishbone_bd_ram_mem0_reg[125][5]/P0001 ,
		_w12956_,
		_w25379_
	);
	LUT2 #(
		.INIT('h8)
	) name14868 (
		\wishbone_bd_ram_mem0_reg[216][5]/P0001 ,
		_w13028_,
		_w25380_
	);
	LUT2 #(
		.INIT('h8)
	) name14869 (
		\wishbone_bd_ram_mem0_reg[236][5]/P0001 ,
		_w12731_,
		_w25381_
	);
	LUT2 #(
		.INIT('h8)
	) name14870 (
		\wishbone_bd_ram_mem0_reg[207][5]/P0001 ,
		_w13180_,
		_w25382_
	);
	LUT2 #(
		.INIT('h8)
	) name14871 (
		\wishbone_bd_ram_mem0_reg[227][5]/P0001 ,
		_w12936_,
		_w25383_
	);
	LUT2 #(
		.INIT('h8)
	) name14872 (
		\wishbone_bd_ram_mem0_reg[138][5]/P0001 ,
		_w12958_,
		_w25384_
	);
	LUT2 #(
		.INIT('h8)
	) name14873 (
		\wishbone_bd_ram_mem0_reg[241][5]/P0001 ,
		_w13006_,
		_w25385_
	);
	LUT2 #(
		.INIT('h8)
	) name14874 (
		\wishbone_bd_ram_mem0_reg[193][5]/P0001 ,
		_w13056_,
		_w25386_
	);
	LUT2 #(
		.INIT('h8)
	) name14875 (
		\wishbone_bd_ram_mem0_reg[141][5]/P0001 ,
		_w13004_,
		_w25387_
	);
	LUT2 #(
		.INIT('h8)
	) name14876 (
		\wishbone_bd_ram_mem0_reg[203][5]/P0001 ,
		_w13158_,
		_w25388_
	);
	LUT2 #(
		.INIT('h8)
	) name14877 (
		\wishbone_bd_ram_mem0_reg[80][5]/P0001 ,
		_w12689_,
		_w25389_
	);
	LUT2 #(
		.INIT('h8)
	) name14878 (
		\wishbone_bd_ram_mem0_reg[37][5]/P0001 ,
		_w13102_,
		_w25390_
	);
	LUT2 #(
		.INIT('h8)
	) name14879 (
		\wishbone_bd_ram_mem0_reg[18][5]/P0001 ,
		_w12679_,
		_w25391_
	);
	LUT2 #(
		.INIT('h8)
	) name14880 (
		\wishbone_bd_ram_mem0_reg[73][5]/P0001 ,
		_w12918_,
		_w25392_
	);
	LUT2 #(
		.INIT('h8)
	) name14881 (
		\wishbone_bd_ram_mem0_reg[159][5]/P0001 ,
		_w12774_,
		_w25393_
	);
	LUT2 #(
		.INIT('h8)
	) name14882 (
		\wishbone_bd_ram_mem0_reg[248][5]/P0001 ,
		_w12789_,
		_w25394_
	);
	LUT2 #(
		.INIT('h8)
	) name14883 (
		\wishbone_bd_ram_mem0_reg[48][5]/P0001 ,
		_w12970_,
		_w25395_
	);
	LUT2 #(
		.INIT('h8)
	) name14884 (
		\wishbone_bd_ram_mem0_reg[121][5]/P0001 ,
		_w13078_,
		_w25396_
	);
	LUT2 #(
		.INIT('h8)
	) name14885 (
		\wishbone_bd_ram_mem0_reg[187][5]/P0001 ,
		_w13196_,
		_w25397_
	);
	LUT2 #(
		.INIT('h8)
	) name14886 (
		\wishbone_bd_ram_mem0_reg[170][5]/P0001 ,
		_w13030_,
		_w25398_
	);
	LUT2 #(
		.INIT('h8)
	) name14887 (
		\wishbone_bd_ram_mem0_reg[29][5]/P0001 ,
		_w12952_,
		_w25399_
	);
	LUT2 #(
		.INIT('h8)
	) name14888 (
		\wishbone_bd_ram_mem0_reg[210][5]/P0001 ,
		_w12924_,
		_w25400_
	);
	LUT2 #(
		.INIT('h8)
	) name14889 (
		\wishbone_bd_ram_mem0_reg[206][5]/P0001 ,
		_w12954_,
		_w25401_
	);
	LUT2 #(
		.INIT('h8)
	) name14890 (
		\wishbone_bd_ram_mem0_reg[204][5]/P0001 ,
		_w13162_,
		_w25402_
	);
	LUT2 #(
		.INIT('h8)
	) name14891 (
		\wishbone_bd_ram_mem0_reg[20][5]/P0001 ,
		_w13174_,
		_w25403_
	);
	LUT2 #(
		.INIT('h8)
	) name14892 (
		\wishbone_bd_ram_mem0_reg[4][5]/P0001 ,
		_w12666_,
		_w25404_
	);
	LUT2 #(
		.INIT('h8)
	) name14893 (
		\wishbone_bd_ram_mem0_reg[208][5]/P0001 ,
		_w13032_,
		_w25405_
	);
	LUT2 #(
		.INIT('h8)
	) name14894 (
		\wishbone_bd_ram_mem0_reg[102][5]/P0001 ,
		_w12685_,
		_w25406_
	);
	LUT2 #(
		.INIT('h8)
	) name14895 (
		\wishbone_bd_ram_mem0_reg[174][5]/P0001 ,
		_w12972_,
		_w25407_
	);
	LUT2 #(
		.INIT('h8)
	) name14896 (
		\wishbone_bd_ram_mem0_reg[231][5]/P0001 ,
		_w12856_,
		_w25408_
	);
	LUT2 #(
		.INIT('h8)
	) name14897 (
		\wishbone_bd_ram_mem0_reg[171][5]/P0001 ,
		_w12910_,
		_w25409_
	);
	LUT2 #(
		.INIT('h8)
	) name14898 (
		\wishbone_bd_ram_mem0_reg[35][5]/P0001 ,
		_w12703_,
		_w25410_
	);
	LUT2 #(
		.INIT('h8)
	) name14899 (
		\wishbone_bd_ram_mem0_reg[3][5]/P0001 ,
		_w12866_,
		_w25411_
	);
	LUT2 #(
		.INIT('h8)
	) name14900 (
		\wishbone_bd_ram_mem0_reg[88][5]/P0001 ,
		_w12860_,
		_w25412_
	);
	LUT2 #(
		.INIT('h8)
	) name14901 (
		\wishbone_bd_ram_mem0_reg[186][5]/P0001 ,
		_w12783_,
		_w25413_
	);
	LUT2 #(
		.INIT('h8)
	) name14902 (
		\wishbone_bd_ram_mem0_reg[26][5]/P0001 ,
		_w12699_,
		_w25414_
	);
	LUT2 #(
		.INIT('h8)
	) name14903 (
		\wishbone_bd_ram_mem0_reg[134][5]/P0001 ,
		_w12763_,
		_w25415_
	);
	LUT2 #(
		.INIT('h8)
	) name14904 (
		\wishbone_bd_ram_mem0_reg[38][5]/P0001 ,
		_w13182_,
		_w25416_
	);
	LUT2 #(
		.INIT('h8)
	) name14905 (
		\wishbone_bd_ram_mem0_reg[220][5]/P0001 ,
		_w13066_,
		_w25417_
	);
	LUT2 #(
		.INIT('h8)
	) name14906 (
		\wishbone_bd_ram_mem0_reg[245][5]/P0001 ,
		_w13022_,
		_w25418_
	);
	LUT2 #(
		.INIT('h8)
	) name14907 (
		\wishbone_bd_ram_mem0_reg[214][5]/P0001 ,
		_w12984_,
		_w25419_
	);
	LUT2 #(
		.INIT('h8)
	) name14908 (
		\wishbone_bd_ram_mem0_reg[108][5]/P0001 ,
		_w13156_,
		_w25420_
	);
	LUT2 #(
		.INIT('h8)
	) name14909 (
		\wishbone_bd_ram_mem0_reg[243][5]/P0001 ,
		_w12804_,
		_w25421_
	);
	LUT2 #(
		.INIT('h8)
	) name14910 (
		\wishbone_bd_ram_mem0_reg[99][5]/P0001 ,
		_w13038_,
		_w25422_
	);
	LUT2 #(
		.INIT('h8)
	) name14911 (
		\wishbone_bd_ram_mem0_reg[93][5]/P0001 ,
		_w13016_,
		_w25423_
	);
	LUT2 #(
		.INIT('h8)
	) name14912 (
		\wishbone_bd_ram_mem0_reg[65][5]/P0001 ,
		_w13176_,
		_w25424_
	);
	LUT2 #(
		.INIT('h8)
	) name14913 (
		\wishbone_bd_ram_mem0_reg[111][5]/P0001 ,
		_w12744_,
		_w25425_
	);
	LUT2 #(
		.INIT('h8)
	) name14914 (
		\wishbone_bd_ram_mem0_reg[229][5]/P0001 ,
		_w12711_,
		_w25426_
	);
	LUT2 #(
		.INIT('h8)
	) name14915 (
		\wishbone_bd_ram_mem0_reg[164][5]/P0001 ,
		_w12876_,
		_w25427_
	);
	LUT2 #(
		.INIT('h8)
	) name14916 (
		\wishbone_bd_ram_mem0_reg[225][5]/P0001 ,
		_w13092_,
		_w25428_
	);
	LUT2 #(
		.INIT('h8)
	) name14917 (
		\wishbone_bd_ram_mem0_reg[153][5]/P0001 ,
		_w12890_,
		_w25429_
	);
	LUT2 #(
		.INIT('h8)
	) name14918 (
		\wishbone_bd_ram_mem0_reg[70][5]/P0001 ,
		_w12840_,
		_w25430_
	);
	LUT2 #(
		.INIT('h8)
	) name14919 (
		\wishbone_bd_ram_mem0_reg[167][5]/P0001 ,
		_w12986_,
		_w25431_
	);
	LUT2 #(
		.INIT('h8)
	) name14920 (
		\wishbone_bd_ram_mem0_reg[132][5]/P0001 ,
		_w12992_,
		_w25432_
	);
	LUT2 #(
		.INIT('h8)
	) name14921 (
		\wishbone_bd_ram_mem0_reg[151][5]/P0001 ,
		_w13142_,
		_w25433_
	);
	LUT2 #(
		.INIT('h8)
	) name14922 (
		\wishbone_bd_ram_mem0_reg[129][5]/P0001 ,
		_w12776_,
		_w25434_
	);
	LUT2 #(
		.INIT('h8)
	) name14923 (
		\wishbone_bd_ram_mem0_reg[31][5]/P0001 ,
		_w13198_,
		_w25435_
	);
	LUT2 #(
		.INIT('h8)
	) name14924 (
		\wishbone_bd_ram_mem0_reg[75][5]/P0001 ,
		_w12826_,
		_w25436_
	);
	LUT2 #(
		.INIT('h8)
	) name14925 (
		\wishbone_bd_ram_mem0_reg[192][5]/P0001 ,
		_w12938_,
		_w25437_
	);
	LUT2 #(
		.INIT('h8)
	) name14926 (
		\wishbone_bd_ram_mem0_reg[25][5]/P0001 ,
		_w13108_,
		_w25438_
	);
	LUT2 #(
		.INIT('h8)
	) name14927 (
		\wishbone_bd_ram_mem0_reg[226][5]/P0001 ,
		_w13138_,
		_w25439_
	);
	LUT2 #(
		.INIT('h8)
	) name14928 (
		\wishbone_bd_ram_mem0_reg[144][5]/P0001 ,
		_w12756_,
		_w25440_
	);
	LUT2 #(
		.INIT('h8)
	) name14929 (
		\wishbone_bd_ram_mem0_reg[224][5]/P0001 ,
		_w12902_,
		_w25441_
	);
	LUT2 #(
		.INIT('h8)
	) name14930 (
		\wishbone_bd_ram_mem0_reg[85][5]/P0001 ,
		_w13216_,
		_w25442_
	);
	LUT2 #(
		.INIT('h8)
	) name14931 (
		\wishbone_bd_ram_mem0_reg[67][5]/P0001 ,
		_w13134_,
		_w25443_
	);
	LUT2 #(
		.INIT('h8)
	) name14932 (
		\wishbone_bd_ram_mem0_reg[142][5]/P0001 ,
		_w12928_,
		_w25444_
	);
	LUT2 #(
		.INIT('h8)
	) name14933 (
		\wishbone_bd_ram_mem0_reg[114][5]/P0001 ,
		_w13202_,
		_w25445_
	);
	LUT2 #(
		.INIT('h8)
	) name14934 (
		\wishbone_bd_ram_mem0_reg[228][5]/P0001 ,
		_w12765_,
		_w25446_
	);
	LUT2 #(
		.INIT('h8)
	) name14935 (
		\wishbone_bd_ram_mem0_reg[110][5]/P0001 ,
		_w13046_,
		_w25447_
	);
	LUT2 #(
		.INIT('h8)
	) name14936 (
		\wishbone_bd_ram_mem0_reg[78][5]/P0001 ,
		_w12874_,
		_w25448_
	);
	LUT2 #(
		.INIT('h8)
	) name14937 (
		\wishbone_bd_ram_mem0_reg[107][5]/P0001 ,
		_w12749_,
		_w25449_
	);
	LUT2 #(
		.INIT('h8)
	) name14938 (
		\wishbone_bd_ram_mem0_reg[165][5]/P0001 ,
		_w13044_,
		_w25450_
	);
	LUT2 #(
		.INIT('h8)
	) name14939 (
		\wishbone_bd_ram_mem0_reg[128][5]/P0001 ,
		_w12793_,
		_w25451_
	);
	LUT2 #(
		.INIT('h8)
	) name14940 (
		\wishbone_bd_ram_mem0_reg[254][5]/P0001 ,
		_w12892_,
		_w25452_
	);
	LUT2 #(
		.INIT('h8)
	) name14941 (
		\wishbone_bd_ram_mem0_reg[62][5]/P0001 ,
		_w12673_,
		_w25453_
	);
	LUT2 #(
		.INIT('h8)
	) name14942 (
		\wishbone_bd_ram_mem0_reg[112][5]/P0001 ,
		_w12733_,
		_w25454_
	);
	LUT2 #(
		.INIT('h8)
	) name14943 (
		\wishbone_bd_ram_mem0_reg[92][5]/P0001 ,
		_w13010_,
		_w25455_
	);
	LUT2 #(
		.INIT('h8)
	) name14944 (
		\wishbone_bd_ram_mem0_reg[168][5]/P0001 ,
		_w13208_,
		_w25456_
	);
	LUT2 #(
		.INIT('h8)
	) name14945 (
		\wishbone_bd_ram_mem0_reg[46][5]/P0001 ,
		_w12884_,
		_w25457_
	);
	LUT2 #(
		.INIT('h8)
	) name14946 (
		\wishbone_bd_ram_mem0_reg[24][5]/P0001 ,
		_w13084_,
		_w25458_
	);
	LUT2 #(
		.INIT('h8)
	) name14947 (
		\wishbone_bd_ram_mem0_reg[59][5]/P0001 ,
		_w12780_,
		_w25459_
	);
	LUT2 #(
		.INIT('h8)
	) name14948 (
		\wishbone_bd_ram_mem0_reg[135][5]/P0001 ,
		_w13124_,
		_w25460_
	);
	LUT2 #(
		.INIT('h8)
	) name14949 (
		\wishbone_bd_ram_mem0_reg[81][5]/P0001 ,
		_w12950_,
		_w25461_
	);
	LUT2 #(
		.INIT('h8)
	) name14950 (
		\wishbone_bd_ram_mem0_reg[178][5]/P0001 ,
		_w12886_,
		_w25462_
	);
	LUT2 #(
		.INIT('h8)
	) name14951 (
		\wishbone_bd_ram_mem0_reg[11][5]/P0001 ,
		_w13194_,
		_w25463_
	);
	LUT2 #(
		.INIT('h8)
	) name14952 (
		\wishbone_bd_ram_mem0_reg[5][5]/P0001 ,
		_w12878_,
		_w25464_
	);
	LUT2 #(
		.INIT('h8)
	) name14953 (
		\wishbone_bd_ram_mem0_reg[251][5]/P0001 ,
		_w13054_,
		_w25465_
	);
	LUT2 #(
		.INIT('h8)
	) name14954 (
		\wishbone_bd_ram_mem0_reg[235][5]/P0001 ,
		_w12696_,
		_w25466_
	);
	LUT2 #(
		.INIT('h8)
	) name14955 (
		\wishbone_bd_ram_mem0_reg[53][5]/P0001 ,
		_w13020_,
		_w25467_
	);
	LUT2 #(
		.INIT('h8)
	) name14956 (
		\wishbone_bd_ram_mem0_reg[223][5]/P0001 ,
		_w12838_,
		_w25468_
	);
	LUT2 #(
		.INIT('h8)
	) name14957 (
		\wishbone_bd_ram_mem0_reg[104][5]/P0001 ,
		_w13148_,
		_w25469_
	);
	LUT2 #(
		.INIT('h8)
	) name14958 (
		\wishbone_bd_ram_mem0_reg[63][5]/P0001 ,
		_w12850_,
		_w25470_
	);
	LUT2 #(
		.INIT('h8)
	) name14959 (
		\wishbone_bd_ram_mem0_reg[90][5]/P0001 ,
		_w12978_,
		_w25471_
	);
	LUT2 #(
		.INIT('h8)
	) name14960 (
		\wishbone_bd_ram_mem0_reg[96][5]/P0001 ,
		_w12912_,
		_w25472_
	);
	LUT2 #(
		.INIT('h8)
	) name14961 (
		\wishbone_bd_ram_mem0_reg[82][5]/P0001 ,
		_w12942_,
		_w25473_
	);
	LUT2 #(
		.INIT('h8)
	) name14962 (
		\wishbone_bd_ram_mem0_reg[222][5]/P0001 ,
		_w13094_,
		_w25474_
	);
	LUT2 #(
		.INIT('h8)
	) name14963 (
		\wishbone_bd_ram_mem0_reg[58][5]/P0001 ,
		_w13070_,
		_w25475_
	);
	LUT2 #(
		.INIT('h8)
	) name14964 (
		\wishbone_bd_ram_mem0_reg[113][5]/P0001 ,
		_w13026_,
		_w25476_
	);
	LUT2 #(
		.INIT('h8)
	) name14965 (
		\wishbone_bd_ram_mem0_reg[249][5]/P0001 ,
		_w12900_,
		_w25477_
	);
	LUT2 #(
		.INIT('h8)
	) name14966 (
		\wishbone_bd_ram_mem0_reg[238][5]/P0001 ,
		_w13160_,
		_w25478_
	);
	LUT2 #(
		.INIT('h8)
	) name14967 (
		\wishbone_bd_ram_mem0_reg[139][5]/P0001 ,
		_w12814_,
		_w25479_
	);
	LUT2 #(
		.INIT('h8)
	) name14968 (
		\wishbone_bd_ram_mem0_reg[97][5]/P0001 ,
		_w13096_,
		_w25480_
	);
	LUT2 #(
		.INIT('h8)
	) name14969 (
		\wishbone_bd_ram_mem0_reg[177][5]/P0001 ,
		_w12996_,
		_w25481_
	);
	LUT2 #(
		.INIT('h8)
	) name14970 (
		\wishbone_bd_ram_mem0_reg[133][5]/P0001 ,
		_w12761_,
		_w25482_
	);
	LUT2 #(
		.INIT('h8)
	) name14971 (
		\wishbone_bd_ram_mem0_reg[87][5]/P0001 ,
		_w13154_,
		_w25483_
	);
	LUT2 #(
		.INIT('h8)
	) name14972 (
		\wishbone_bd_ram_mem0_reg[179][5]/P0001 ,
		_w13050_,
		_w25484_
	);
	LUT2 #(
		.INIT('h8)
	) name14973 (
		\wishbone_bd_ram_mem0_reg[140][5]/P0001 ,
		_w12894_,
		_w25485_
	);
	LUT2 #(
		.INIT('h8)
	) name14974 (
		\wishbone_bd_ram_mem0_reg[69][5]/P0001 ,
		_w12738_,
		_w25486_
	);
	LUT2 #(
		.INIT('h8)
	) name14975 (
		\wishbone_bd_ram_mem0_reg[244][5]/P0001 ,
		_w12747_,
		_w25487_
	);
	LUT2 #(
		.INIT('h8)
	) name14976 (
		\wishbone_bd_ram_mem0_reg[202][5]/P0001 ,
		_w12870_,
		_w25488_
	);
	LUT2 #(
		.INIT('h8)
	) name14977 (
		\wishbone_bd_ram_mem0_reg[190][5]/P0001 ,
		_w12858_,
		_w25489_
	);
	LUT2 #(
		.INIT('h8)
	) name14978 (
		\wishbone_bd_ram_mem0_reg[103][5]/P0001 ,
		_w12846_,
		_w25490_
	);
	LUT2 #(
		.INIT('h8)
	) name14979 (
		\wishbone_bd_ram_mem0_reg[221][5]/P0001 ,
		_w12802_,
		_w25491_
	);
	LUT2 #(
		.INIT('h8)
	) name14980 (
		\wishbone_bd_ram_mem0_reg[9][5]/P0001 ,
		_w12808_,
		_w25492_
	);
	LUT2 #(
		.INIT('h8)
	) name14981 (
		\wishbone_bd_ram_mem0_reg[42][5]/P0001 ,
		_w12842_,
		_w25493_
	);
	LUT2 #(
		.INIT('h8)
	) name14982 (
		\wishbone_bd_ram_mem0_reg[10][5]/P0001 ,
		_w13172_,
		_w25494_
	);
	LUT2 #(
		.INIT('h8)
	) name14983 (
		\wishbone_bd_ram_mem0_reg[27][5]/P0001 ,
		_w12880_,
		_w25495_
	);
	LUT2 #(
		.INIT('h8)
	) name14984 (
		\wishbone_bd_ram_mem0_reg[162][5]/P0001 ,
		_w13098_,
		_w25496_
	);
	LUT2 #(
		.INIT('h8)
	) name14985 (
		\wishbone_bd_ram_mem0_reg[250][5]/P0001 ,
		_w13128_,
		_w25497_
	);
	LUT2 #(
		.INIT('h8)
	) name14986 (
		\wishbone_bd_ram_mem0_reg[184][5]/P0001 ,
		_w13062_,
		_w25498_
	);
	LUT2 #(
		.INIT('h8)
	) name14987 (
		\wishbone_bd_ram_mem0_reg[16][5]/P0001 ,
		_w13140_,
		_w25499_
	);
	LUT2 #(
		.INIT('h8)
	) name14988 (
		\wishbone_bd_ram_mem0_reg[176][5]/P0001 ,
		_w12868_,
		_w25500_
	);
	LUT2 #(
		.INIT('h8)
	) name14989 (
		\wishbone_bd_ram_mem0_reg[219][5]/P0001 ,
		_w12806_,
		_w25501_
	);
	LUT2 #(
		.INIT('h8)
	) name14990 (
		\wishbone_bd_ram_mem0_reg[0][5]/P0001 ,
		_w12717_,
		_w25502_
	);
	LUT2 #(
		.INIT('h8)
	) name14991 (
		\wishbone_bd_ram_mem0_reg[79][5]/P0001 ,
		_w13212_,
		_w25503_
	);
	LUT2 #(
		.INIT('h8)
	) name14992 (
		\wishbone_bd_ram_mem0_reg[156][5]/P0001 ,
		_w13190_,
		_w25504_
	);
	LUT2 #(
		.INIT('h8)
	) name14993 (
		\wishbone_bd_ram_mem0_reg[66][5]/P0001 ,
		_w12824_,
		_w25505_
	);
	LUT2 #(
		.INIT('h8)
	) name14994 (
		\wishbone_bd_ram_mem0_reg[163][5]/P0001 ,
		_w12882_,
		_w25506_
	);
	LUT2 #(
		.INIT('h8)
	) name14995 (
		\wishbone_bd_ram_mem0_reg[83][5]/P0001 ,
		_w12916_,
		_w25507_
	);
	LUT2 #(
		.INIT('h8)
	) name14996 (
		\wishbone_bd_ram_mem0_reg[152][5]/P0001 ,
		_w12966_,
		_w25508_
	);
	LUT2 #(
		.INIT('h8)
	) name14997 (
		\wishbone_bd_ram_mem0_reg[47][5]/P0001 ,
		_w12904_,
		_w25509_
	);
	LUT2 #(
		.INIT('h8)
	) name14998 (
		\wishbone_bd_ram_mem0_reg[40][5]/P0001 ,
		_w13132_,
		_w25510_
	);
	LUT2 #(
		.INIT('h8)
	) name14999 (
		\wishbone_bd_ram_mem0_reg[115][5]/P0001 ,
		_w13112_,
		_w25511_
	);
	LUT2 #(
		.INIT('h8)
	) name15000 (
		\wishbone_bd_ram_mem0_reg[22][5]/P0001 ,
		_w13110_,
		_w25512_
	);
	LUT2 #(
		.INIT('h8)
	) name15001 (
		\wishbone_bd_ram_mem0_reg[84][5]/P0001 ,
		_w12934_,
		_w25513_
	);
	LUT2 #(
		.INIT('h8)
	) name15002 (
		\wishbone_bd_ram_mem0_reg[17][5]/P0001 ,
		_w12848_,
		_w25514_
	);
	LUT2 #(
		.INIT('h8)
	) name15003 (
		\wishbone_bd_ram_mem0_reg[252][5]/P0001 ,
		_w13080_,
		_w25515_
	);
	LUT2 #(
		.INIT('h8)
	) name15004 (
		\wishbone_bd_ram_mem0_reg[155][5]/P0001 ,
		_w13122_,
		_w25516_
	);
	LUT2 #(
		.INIT('h8)
	) name15005 (
		\wishbone_bd_ram_mem0_reg[52][5]/P0001 ,
		_w13082_,
		_w25517_
	);
	LUT2 #(
		.INIT('h8)
	) name15006 (
		\wishbone_bd_ram_mem0_reg[8][5]/P0001 ,
		_w12920_,
		_w25518_
	);
	LUT2 #(
		.INIT('h8)
	) name15007 (
		\wishbone_bd_ram_mem0_reg[101][5]/P0001 ,
		_w13192_,
		_w25519_
	);
	LUT2 #(
		.INIT('h8)
	) name15008 (
		\wishbone_bd_ram_mem0_reg[217][5]/P0001 ,
		_w13188_,
		_w25520_
	);
	LUT2 #(
		.INIT('h8)
	) name15009 (
		\wishbone_bd_ram_mem0_reg[77][5]/P0001 ,
		_w12982_,
		_w25521_
	);
	LUT2 #(
		.INIT('h8)
	) name15010 (
		\wishbone_bd_ram_mem0_reg[182][5]/P0001 ,
		_w12820_,
		_w25522_
	);
	LUT2 #(
		.INIT('h8)
	) name15011 (
		\wishbone_bd_ram_mem0_reg[158][5]/P0001 ,
		_w12898_,
		_w25523_
	);
	LUT2 #(
		.INIT('h8)
	) name15012 (
		\wishbone_bd_ram_mem0_reg[7][5]/P0001 ,
		_w12728_,
		_w25524_
	);
	LUT2 #(
		.INIT('h8)
	) name15013 (
		\wishbone_bd_ram_mem0_reg[89][5]/P0001 ,
		_w12964_,
		_w25525_
	);
	LUT2 #(
		.INIT('h8)
	) name15014 (
		\wishbone_bd_ram_mem0_reg[2][5]/P0001 ,
		_w13088_,
		_w25526_
	);
	LUT2 #(
		.INIT('h8)
	) name15015 (
		\wishbone_bd_ram_mem0_reg[212][5]/P0001 ,
		_w12796_,
		_w25527_
	);
	LUT2 #(
		.INIT('h8)
	) name15016 (
		\wishbone_bd_ram_mem0_reg[86][5]/P0001 ,
		_w12735_,
		_w25528_
	);
	LUT2 #(
		.INIT('h8)
	) name15017 (
		\wishbone_bd_ram_mem0_reg[230][5]/P0001 ,
		_w13036_,
		_w25529_
	);
	LUT2 #(
		.INIT('h8)
	) name15018 (
		\wishbone_bd_ram_mem0_reg[205][5]/P0001 ,
		_w13068_,
		_w25530_
	);
	LUT2 #(
		.INIT('h8)
	) name15019 (
		\wishbone_bd_ram_mem0_reg[240][5]/P0001 ,
		_w12864_,
		_w25531_
	);
	LUT2 #(
		.INIT('h8)
	) name15020 (
		\wishbone_bd_ram_mem0_reg[255][5]/P0001 ,
		_w13072_,
		_w25532_
	);
	LUT2 #(
		.INIT('h8)
	) name15021 (
		\wishbone_bd_ram_mem0_reg[126][5]/P0001 ,
		_w13218_,
		_w25533_
	);
	LUT2 #(
		.INIT('h8)
	) name15022 (
		\wishbone_bd_ram_mem0_reg[191][5]/P0001 ,
		_w13034_,
		_w25534_
	);
	LUT2 #(
		.INIT('h8)
	) name15023 (
		\wishbone_bd_ram_mem0_reg[45][5]/P0001 ,
		_w12908_,
		_w25535_
	);
	LUT2 #(
		.INIT('h8)
	) name15024 (
		\wishbone_bd_ram_mem0_reg[19][5]/P0001 ,
		_w13012_,
		_w25536_
	);
	LUT2 #(
		.INIT('h8)
	) name15025 (
		\wishbone_bd_ram_mem0_reg[119][5]/P0001 ,
		_w13048_,
		_w25537_
	);
	LUT2 #(
		.INIT('h8)
	) name15026 (
		\wishbone_bd_ram_mem0_reg[148][5]/P0001 ,
		_w13000_,
		_w25538_
	);
	LUT2 #(
		.INIT('h8)
	) name15027 (
		\wishbone_bd_ram_mem0_reg[21][5]/P0001 ,
		_w12906_,
		_w25539_
	);
	LUT2 #(
		.INIT('h8)
	) name15028 (
		\wishbone_bd_ram_mem0_reg[68][5]/P0001 ,
		_w12946_,
		_w25540_
	);
	LUT2 #(
		.INIT('h8)
	) name15029 (
		\wishbone_bd_ram_mem0_reg[233][5]/P0001 ,
		_w12836_,
		_w25541_
	);
	LUT2 #(
		.INIT('h8)
	) name15030 (
		\wishbone_bd_ram_mem0_reg[161][5]/P0001 ,
		_w12754_,
		_w25542_
	);
	LUT2 #(
		.INIT('h8)
	) name15031 (
		\wishbone_bd_ram_mem0_reg[6][5]/P0001 ,
		_w12968_,
		_w25543_
	);
	LUT2 #(
		.INIT('h8)
	) name15032 (
		\wishbone_bd_ram_mem0_reg[188][5]/P0001 ,
		_w12948_,
		_w25544_
	);
	LUT2 #(
		.INIT('h8)
	) name15033 (
		\wishbone_bd_ram_mem0_reg[213][5]/P0001 ,
		_w13002_,
		_w25545_
	);
	LUT2 #(
		.INIT('h8)
	) name15034 (
		\wishbone_bd_ram_mem0_reg[130][5]/P0001 ,
		_w12914_,
		_w25546_
	);
	LUT2 #(
		.INIT('h8)
	) name15035 (
		\wishbone_bd_ram_mem0_reg[54][5]/P0001 ,
		_w12770_,
		_w25547_
	);
	LUT2 #(
		.INIT('h8)
	) name15036 (
		\wishbone_bd_ram_mem0_reg[36][5]/P0001 ,
		_w12800_,
		_w25548_
	);
	LUT2 #(
		.INIT('h8)
	) name15037 (
		\wishbone_bd_ram_mem0_reg[253][5]/P0001 ,
		_w13100_,
		_w25549_
	);
	LUT2 #(
		.INIT('h8)
	) name15038 (
		\wishbone_bd_ram_mem0_reg[109][5]/P0001 ,
		_w12888_,
		_w25550_
	);
	LUT2 #(
		.INIT('h8)
	) name15039 (
		\wishbone_bd_ram_mem0_reg[72][5]/P0001 ,
		_w12810_,
		_w25551_
	);
	LUT2 #(
		.INIT('h8)
	) name15040 (
		\wishbone_bd_ram_mem0_reg[199][5]/P0001 ,
		_w12768_,
		_w25552_
	);
	LUT2 #(
		.INIT('h8)
	) name15041 (
		\wishbone_bd_ram_mem0_reg[160][5]/P0001 ,
		_w12872_,
		_w25553_
	);
	LUT2 #(
		.INIT('h8)
	) name15042 (
		\wishbone_bd_ram_mem0_reg[117][5]/P0001 ,
		_w12715_,
		_w25554_
	);
	LUT2 #(
		.INIT('h8)
	) name15043 (
		\wishbone_bd_ram_mem0_reg[137][5]/P0001 ,
		_w13168_,
		_w25555_
	);
	LUT2 #(
		.INIT('h8)
	) name15044 (
		\wishbone_bd_ram_mem0_reg[147][5]/P0001 ,
		_w13146_,
		_w25556_
	);
	LUT2 #(
		.INIT('h8)
	) name15045 (
		\wishbone_bd_ram_mem0_reg[234][5]/P0001 ,
		_w13214_,
		_w25557_
	);
	LUT2 #(
		.INIT('h8)
	) name15046 (
		\wishbone_bd_ram_mem0_reg[124][5]/P0001 ,
		_w13058_,
		_w25558_
	);
	LUT2 #(
		.INIT('h8)
	) name15047 (
		\wishbone_bd_ram_mem0_reg[34][5]/P0001 ,
		_w12930_,
		_w25559_
	);
	LUT2 #(
		.INIT('h8)
	) name15048 (
		\wishbone_bd_ram_mem0_reg[196][5]/P0001 ,
		_w13090_,
		_w25560_
	);
	LUT2 #(
		.INIT('h1)
	) name15049 (
		_w25305_,
		_w25306_,
		_w25561_
	);
	LUT2 #(
		.INIT('h1)
	) name15050 (
		_w25307_,
		_w25308_,
		_w25562_
	);
	LUT2 #(
		.INIT('h1)
	) name15051 (
		_w25309_,
		_w25310_,
		_w25563_
	);
	LUT2 #(
		.INIT('h1)
	) name15052 (
		_w25311_,
		_w25312_,
		_w25564_
	);
	LUT2 #(
		.INIT('h1)
	) name15053 (
		_w25313_,
		_w25314_,
		_w25565_
	);
	LUT2 #(
		.INIT('h1)
	) name15054 (
		_w25315_,
		_w25316_,
		_w25566_
	);
	LUT2 #(
		.INIT('h1)
	) name15055 (
		_w25317_,
		_w25318_,
		_w25567_
	);
	LUT2 #(
		.INIT('h1)
	) name15056 (
		_w25319_,
		_w25320_,
		_w25568_
	);
	LUT2 #(
		.INIT('h1)
	) name15057 (
		_w25321_,
		_w25322_,
		_w25569_
	);
	LUT2 #(
		.INIT('h1)
	) name15058 (
		_w25323_,
		_w25324_,
		_w25570_
	);
	LUT2 #(
		.INIT('h1)
	) name15059 (
		_w25325_,
		_w25326_,
		_w25571_
	);
	LUT2 #(
		.INIT('h1)
	) name15060 (
		_w25327_,
		_w25328_,
		_w25572_
	);
	LUT2 #(
		.INIT('h1)
	) name15061 (
		_w25329_,
		_w25330_,
		_w25573_
	);
	LUT2 #(
		.INIT('h1)
	) name15062 (
		_w25331_,
		_w25332_,
		_w25574_
	);
	LUT2 #(
		.INIT('h1)
	) name15063 (
		_w25333_,
		_w25334_,
		_w25575_
	);
	LUT2 #(
		.INIT('h1)
	) name15064 (
		_w25335_,
		_w25336_,
		_w25576_
	);
	LUT2 #(
		.INIT('h1)
	) name15065 (
		_w25337_,
		_w25338_,
		_w25577_
	);
	LUT2 #(
		.INIT('h1)
	) name15066 (
		_w25339_,
		_w25340_,
		_w25578_
	);
	LUT2 #(
		.INIT('h1)
	) name15067 (
		_w25341_,
		_w25342_,
		_w25579_
	);
	LUT2 #(
		.INIT('h1)
	) name15068 (
		_w25343_,
		_w25344_,
		_w25580_
	);
	LUT2 #(
		.INIT('h1)
	) name15069 (
		_w25345_,
		_w25346_,
		_w25581_
	);
	LUT2 #(
		.INIT('h1)
	) name15070 (
		_w25347_,
		_w25348_,
		_w25582_
	);
	LUT2 #(
		.INIT('h1)
	) name15071 (
		_w25349_,
		_w25350_,
		_w25583_
	);
	LUT2 #(
		.INIT('h1)
	) name15072 (
		_w25351_,
		_w25352_,
		_w25584_
	);
	LUT2 #(
		.INIT('h1)
	) name15073 (
		_w25353_,
		_w25354_,
		_w25585_
	);
	LUT2 #(
		.INIT('h1)
	) name15074 (
		_w25355_,
		_w25356_,
		_w25586_
	);
	LUT2 #(
		.INIT('h1)
	) name15075 (
		_w25357_,
		_w25358_,
		_w25587_
	);
	LUT2 #(
		.INIT('h1)
	) name15076 (
		_w25359_,
		_w25360_,
		_w25588_
	);
	LUT2 #(
		.INIT('h1)
	) name15077 (
		_w25361_,
		_w25362_,
		_w25589_
	);
	LUT2 #(
		.INIT('h1)
	) name15078 (
		_w25363_,
		_w25364_,
		_w25590_
	);
	LUT2 #(
		.INIT('h1)
	) name15079 (
		_w25365_,
		_w25366_,
		_w25591_
	);
	LUT2 #(
		.INIT('h1)
	) name15080 (
		_w25367_,
		_w25368_,
		_w25592_
	);
	LUT2 #(
		.INIT('h1)
	) name15081 (
		_w25369_,
		_w25370_,
		_w25593_
	);
	LUT2 #(
		.INIT('h1)
	) name15082 (
		_w25371_,
		_w25372_,
		_w25594_
	);
	LUT2 #(
		.INIT('h1)
	) name15083 (
		_w25373_,
		_w25374_,
		_w25595_
	);
	LUT2 #(
		.INIT('h1)
	) name15084 (
		_w25375_,
		_w25376_,
		_w25596_
	);
	LUT2 #(
		.INIT('h1)
	) name15085 (
		_w25377_,
		_w25378_,
		_w25597_
	);
	LUT2 #(
		.INIT('h1)
	) name15086 (
		_w25379_,
		_w25380_,
		_w25598_
	);
	LUT2 #(
		.INIT('h1)
	) name15087 (
		_w25381_,
		_w25382_,
		_w25599_
	);
	LUT2 #(
		.INIT('h1)
	) name15088 (
		_w25383_,
		_w25384_,
		_w25600_
	);
	LUT2 #(
		.INIT('h1)
	) name15089 (
		_w25385_,
		_w25386_,
		_w25601_
	);
	LUT2 #(
		.INIT('h1)
	) name15090 (
		_w25387_,
		_w25388_,
		_w25602_
	);
	LUT2 #(
		.INIT('h1)
	) name15091 (
		_w25389_,
		_w25390_,
		_w25603_
	);
	LUT2 #(
		.INIT('h1)
	) name15092 (
		_w25391_,
		_w25392_,
		_w25604_
	);
	LUT2 #(
		.INIT('h1)
	) name15093 (
		_w25393_,
		_w25394_,
		_w25605_
	);
	LUT2 #(
		.INIT('h1)
	) name15094 (
		_w25395_,
		_w25396_,
		_w25606_
	);
	LUT2 #(
		.INIT('h1)
	) name15095 (
		_w25397_,
		_w25398_,
		_w25607_
	);
	LUT2 #(
		.INIT('h1)
	) name15096 (
		_w25399_,
		_w25400_,
		_w25608_
	);
	LUT2 #(
		.INIT('h1)
	) name15097 (
		_w25401_,
		_w25402_,
		_w25609_
	);
	LUT2 #(
		.INIT('h1)
	) name15098 (
		_w25403_,
		_w25404_,
		_w25610_
	);
	LUT2 #(
		.INIT('h1)
	) name15099 (
		_w25405_,
		_w25406_,
		_w25611_
	);
	LUT2 #(
		.INIT('h1)
	) name15100 (
		_w25407_,
		_w25408_,
		_w25612_
	);
	LUT2 #(
		.INIT('h1)
	) name15101 (
		_w25409_,
		_w25410_,
		_w25613_
	);
	LUT2 #(
		.INIT('h1)
	) name15102 (
		_w25411_,
		_w25412_,
		_w25614_
	);
	LUT2 #(
		.INIT('h1)
	) name15103 (
		_w25413_,
		_w25414_,
		_w25615_
	);
	LUT2 #(
		.INIT('h1)
	) name15104 (
		_w25415_,
		_w25416_,
		_w25616_
	);
	LUT2 #(
		.INIT('h1)
	) name15105 (
		_w25417_,
		_w25418_,
		_w25617_
	);
	LUT2 #(
		.INIT('h1)
	) name15106 (
		_w25419_,
		_w25420_,
		_w25618_
	);
	LUT2 #(
		.INIT('h1)
	) name15107 (
		_w25421_,
		_w25422_,
		_w25619_
	);
	LUT2 #(
		.INIT('h1)
	) name15108 (
		_w25423_,
		_w25424_,
		_w25620_
	);
	LUT2 #(
		.INIT('h1)
	) name15109 (
		_w25425_,
		_w25426_,
		_w25621_
	);
	LUT2 #(
		.INIT('h1)
	) name15110 (
		_w25427_,
		_w25428_,
		_w25622_
	);
	LUT2 #(
		.INIT('h1)
	) name15111 (
		_w25429_,
		_w25430_,
		_w25623_
	);
	LUT2 #(
		.INIT('h1)
	) name15112 (
		_w25431_,
		_w25432_,
		_w25624_
	);
	LUT2 #(
		.INIT('h1)
	) name15113 (
		_w25433_,
		_w25434_,
		_w25625_
	);
	LUT2 #(
		.INIT('h1)
	) name15114 (
		_w25435_,
		_w25436_,
		_w25626_
	);
	LUT2 #(
		.INIT('h1)
	) name15115 (
		_w25437_,
		_w25438_,
		_w25627_
	);
	LUT2 #(
		.INIT('h1)
	) name15116 (
		_w25439_,
		_w25440_,
		_w25628_
	);
	LUT2 #(
		.INIT('h1)
	) name15117 (
		_w25441_,
		_w25442_,
		_w25629_
	);
	LUT2 #(
		.INIT('h1)
	) name15118 (
		_w25443_,
		_w25444_,
		_w25630_
	);
	LUT2 #(
		.INIT('h1)
	) name15119 (
		_w25445_,
		_w25446_,
		_w25631_
	);
	LUT2 #(
		.INIT('h1)
	) name15120 (
		_w25447_,
		_w25448_,
		_w25632_
	);
	LUT2 #(
		.INIT('h1)
	) name15121 (
		_w25449_,
		_w25450_,
		_w25633_
	);
	LUT2 #(
		.INIT('h1)
	) name15122 (
		_w25451_,
		_w25452_,
		_w25634_
	);
	LUT2 #(
		.INIT('h1)
	) name15123 (
		_w25453_,
		_w25454_,
		_w25635_
	);
	LUT2 #(
		.INIT('h1)
	) name15124 (
		_w25455_,
		_w25456_,
		_w25636_
	);
	LUT2 #(
		.INIT('h1)
	) name15125 (
		_w25457_,
		_w25458_,
		_w25637_
	);
	LUT2 #(
		.INIT('h1)
	) name15126 (
		_w25459_,
		_w25460_,
		_w25638_
	);
	LUT2 #(
		.INIT('h1)
	) name15127 (
		_w25461_,
		_w25462_,
		_w25639_
	);
	LUT2 #(
		.INIT('h1)
	) name15128 (
		_w25463_,
		_w25464_,
		_w25640_
	);
	LUT2 #(
		.INIT('h1)
	) name15129 (
		_w25465_,
		_w25466_,
		_w25641_
	);
	LUT2 #(
		.INIT('h1)
	) name15130 (
		_w25467_,
		_w25468_,
		_w25642_
	);
	LUT2 #(
		.INIT('h1)
	) name15131 (
		_w25469_,
		_w25470_,
		_w25643_
	);
	LUT2 #(
		.INIT('h1)
	) name15132 (
		_w25471_,
		_w25472_,
		_w25644_
	);
	LUT2 #(
		.INIT('h1)
	) name15133 (
		_w25473_,
		_w25474_,
		_w25645_
	);
	LUT2 #(
		.INIT('h1)
	) name15134 (
		_w25475_,
		_w25476_,
		_w25646_
	);
	LUT2 #(
		.INIT('h1)
	) name15135 (
		_w25477_,
		_w25478_,
		_w25647_
	);
	LUT2 #(
		.INIT('h1)
	) name15136 (
		_w25479_,
		_w25480_,
		_w25648_
	);
	LUT2 #(
		.INIT('h1)
	) name15137 (
		_w25481_,
		_w25482_,
		_w25649_
	);
	LUT2 #(
		.INIT('h1)
	) name15138 (
		_w25483_,
		_w25484_,
		_w25650_
	);
	LUT2 #(
		.INIT('h1)
	) name15139 (
		_w25485_,
		_w25486_,
		_w25651_
	);
	LUT2 #(
		.INIT('h1)
	) name15140 (
		_w25487_,
		_w25488_,
		_w25652_
	);
	LUT2 #(
		.INIT('h1)
	) name15141 (
		_w25489_,
		_w25490_,
		_w25653_
	);
	LUT2 #(
		.INIT('h1)
	) name15142 (
		_w25491_,
		_w25492_,
		_w25654_
	);
	LUT2 #(
		.INIT('h1)
	) name15143 (
		_w25493_,
		_w25494_,
		_w25655_
	);
	LUT2 #(
		.INIT('h1)
	) name15144 (
		_w25495_,
		_w25496_,
		_w25656_
	);
	LUT2 #(
		.INIT('h1)
	) name15145 (
		_w25497_,
		_w25498_,
		_w25657_
	);
	LUT2 #(
		.INIT('h1)
	) name15146 (
		_w25499_,
		_w25500_,
		_w25658_
	);
	LUT2 #(
		.INIT('h1)
	) name15147 (
		_w25501_,
		_w25502_,
		_w25659_
	);
	LUT2 #(
		.INIT('h1)
	) name15148 (
		_w25503_,
		_w25504_,
		_w25660_
	);
	LUT2 #(
		.INIT('h1)
	) name15149 (
		_w25505_,
		_w25506_,
		_w25661_
	);
	LUT2 #(
		.INIT('h1)
	) name15150 (
		_w25507_,
		_w25508_,
		_w25662_
	);
	LUT2 #(
		.INIT('h1)
	) name15151 (
		_w25509_,
		_w25510_,
		_w25663_
	);
	LUT2 #(
		.INIT('h1)
	) name15152 (
		_w25511_,
		_w25512_,
		_w25664_
	);
	LUT2 #(
		.INIT('h1)
	) name15153 (
		_w25513_,
		_w25514_,
		_w25665_
	);
	LUT2 #(
		.INIT('h1)
	) name15154 (
		_w25515_,
		_w25516_,
		_w25666_
	);
	LUT2 #(
		.INIT('h1)
	) name15155 (
		_w25517_,
		_w25518_,
		_w25667_
	);
	LUT2 #(
		.INIT('h1)
	) name15156 (
		_w25519_,
		_w25520_,
		_w25668_
	);
	LUT2 #(
		.INIT('h1)
	) name15157 (
		_w25521_,
		_w25522_,
		_w25669_
	);
	LUT2 #(
		.INIT('h1)
	) name15158 (
		_w25523_,
		_w25524_,
		_w25670_
	);
	LUT2 #(
		.INIT('h1)
	) name15159 (
		_w25525_,
		_w25526_,
		_w25671_
	);
	LUT2 #(
		.INIT('h1)
	) name15160 (
		_w25527_,
		_w25528_,
		_w25672_
	);
	LUT2 #(
		.INIT('h1)
	) name15161 (
		_w25529_,
		_w25530_,
		_w25673_
	);
	LUT2 #(
		.INIT('h1)
	) name15162 (
		_w25531_,
		_w25532_,
		_w25674_
	);
	LUT2 #(
		.INIT('h1)
	) name15163 (
		_w25533_,
		_w25534_,
		_w25675_
	);
	LUT2 #(
		.INIT('h1)
	) name15164 (
		_w25535_,
		_w25536_,
		_w25676_
	);
	LUT2 #(
		.INIT('h1)
	) name15165 (
		_w25537_,
		_w25538_,
		_w25677_
	);
	LUT2 #(
		.INIT('h1)
	) name15166 (
		_w25539_,
		_w25540_,
		_w25678_
	);
	LUT2 #(
		.INIT('h1)
	) name15167 (
		_w25541_,
		_w25542_,
		_w25679_
	);
	LUT2 #(
		.INIT('h1)
	) name15168 (
		_w25543_,
		_w25544_,
		_w25680_
	);
	LUT2 #(
		.INIT('h1)
	) name15169 (
		_w25545_,
		_w25546_,
		_w25681_
	);
	LUT2 #(
		.INIT('h1)
	) name15170 (
		_w25547_,
		_w25548_,
		_w25682_
	);
	LUT2 #(
		.INIT('h1)
	) name15171 (
		_w25549_,
		_w25550_,
		_w25683_
	);
	LUT2 #(
		.INIT('h1)
	) name15172 (
		_w25551_,
		_w25552_,
		_w25684_
	);
	LUT2 #(
		.INIT('h1)
	) name15173 (
		_w25553_,
		_w25554_,
		_w25685_
	);
	LUT2 #(
		.INIT('h1)
	) name15174 (
		_w25555_,
		_w25556_,
		_w25686_
	);
	LUT2 #(
		.INIT('h1)
	) name15175 (
		_w25557_,
		_w25558_,
		_w25687_
	);
	LUT2 #(
		.INIT('h1)
	) name15176 (
		_w25559_,
		_w25560_,
		_w25688_
	);
	LUT2 #(
		.INIT('h8)
	) name15177 (
		_w25687_,
		_w25688_,
		_w25689_
	);
	LUT2 #(
		.INIT('h8)
	) name15178 (
		_w25685_,
		_w25686_,
		_w25690_
	);
	LUT2 #(
		.INIT('h8)
	) name15179 (
		_w25683_,
		_w25684_,
		_w25691_
	);
	LUT2 #(
		.INIT('h8)
	) name15180 (
		_w25681_,
		_w25682_,
		_w25692_
	);
	LUT2 #(
		.INIT('h8)
	) name15181 (
		_w25679_,
		_w25680_,
		_w25693_
	);
	LUT2 #(
		.INIT('h8)
	) name15182 (
		_w25677_,
		_w25678_,
		_w25694_
	);
	LUT2 #(
		.INIT('h8)
	) name15183 (
		_w25675_,
		_w25676_,
		_w25695_
	);
	LUT2 #(
		.INIT('h8)
	) name15184 (
		_w25673_,
		_w25674_,
		_w25696_
	);
	LUT2 #(
		.INIT('h8)
	) name15185 (
		_w25671_,
		_w25672_,
		_w25697_
	);
	LUT2 #(
		.INIT('h8)
	) name15186 (
		_w25669_,
		_w25670_,
		_w25698_
	);
	LUT2 #(
		.INIT('h8)
	) name15187 (
		_w25667_,
		_w25668_,
		_w25699_
	);
	LUT2 #(
		.INIT('h8)
	) name15188 (
		_w25665_,
		_w25666_,
		_w25700_
	);
	LUT2 #(
		.INIT('h8)
	) name15189 (
		_w25663_,
		_w25664_,
		_w25701_
	);
	LUT2 #(
		.INIT('h8)
	) name15190 (
		_w25661_,
		_w25662_,
		_w25702_
	);
	LUT2 #(
		.INIT('h8)
	) name15191 (
		_w25659_,
		_w25660_,
		_w25703_
	);
	LUT2 #(
		.INIT('h8)
	) name15192 (
		_w25657_,
		_w25658_,
		_w25704_
	);
	LUT2 #(
		.INIT('h8)
	) name15193 (
		_w25655_,
		_w25656_,
		_w25705_
	);
	LUT2 #(
		.INIT('h8)
	) name15194 (
		_w25653_,
		_w25654_,
		_w25706_
	);
	LUT2 #(
		.INIT('h8)
	) name15195 (
		_w25651_,
		_w25652_,
		_w25707_
	);
	LUT2 #(
		.INIT('h8)
	) name15196 (
		_w25649_,
		_w25650_,
		_w25708_
	);
	LUT2 #(
		.INIT('h8)
	) name15197 (
		_w25647_,
		_w25648_,
		_w25709_
	);
	LUT2 #(
		.INIT('h8)
	) name15198 (
		_w25645_,
		_w25646_,
		_w25710_
	);
	LUT2 #(
		.INIT('h8)
	) name15199 (
		_w25643_,
		_w25644_,
		_w25711_
	);
	LUT2 #(
		.INIT('h8)
	) name15200 (
		_w25641_,
		_w25642_,
		_w25712_
	);
	LUT2 #(
		.INIT('h8)
	) name15201 (
		_w25639_,
		_w25640_,
		_w25713_
	);
	LUT2 #(
		.INIT('h8)
	) name15202 (
		_w25637_,
		_w25638_,
		_w25714_
	);
	LUT2 #(
		.INIT('h8)
	) name15203 (
		_w25635_,
		_w25636_,
		_w25715_
	);
	LUT2 #(
		.INIT('h8)
	) name15204 (
		_w25633_,
		_w25634_,
		_w25716_
	);
	LUT2 #(
		.INIT('h8)
	) name15205 (
		_w25631_,
		_w25632_,
		_w25717_
	);
	LUT2 #(
		.INIT('h8)
	) name15206 (
		_w25629_,
		_w25630_,
		_w25718_
	);
	LUT2 #(
		.INIT('h8)
	) name15207 (
		_w25627_,
		_w25628_,
		_w25719_
	);
	LUT2 #(
		.INIT('h8)
	) name15208 (
		_w25625_,
		_w25626_,
		_w25720_
	);
	LUT2 #(
		.INIT('h8)
	) name15209 (
		_w25623_,
		_w25624_,
		_w25721_
	);
	LUT2 #(
		.INIT('h8)
	) name15210 (
		_w25621_,
		_w25622_,
		_w25722_
	);
	LUT2 #(
		.INIT('h8)
	) name15211 (
		_w25619_,
		_w25620_,
		_w25723_
	);
	LUT2 #(
		.INIT('h8)
	) name15212 (
		_w25617_,
		_w25618_,
		_w25724_
	);
	LUT2 #(
		.INIT('h8)
	) name15213 (
		_w25615_,
		_w25616_,
		_w25725_
	);
	LUT2 #(
		.INIT('h8)
	) name15214 (
		_w25613_,
		_w25614_,
		_w25726_
	);
	LUT2 #(
		.INIT('h8)
	) name15215 (
		_w25611_,
		_w25612_,
		_w25727_
	);
	LUT2 #(
		.INIT('h8)
	) name15216 (
		_w25609_,
		_w25610_,
		_w25728_
	);
	LUT2 #(
		.INIT('h8)
	) name15217 (
		_w25607_,
		_w25608_,
		_w25729_
	);
	LUT2 #(
		.INIT('h8)
	) name15218 (
		_w25605_,
		_w25606_,
		_w25730_
	);
	LUT2 #(
		.INIT('h8)
	) name15219 (
		_w25603_,
		_w25604_,
		_w25731_
	);
	LUT2 #(
		.INIT('h8)
	) name15220 (
		_w25601_,
		_w25602_,
		_w25732_
	);
	LUT2 #(
		.INIT('h8)
	) name15221 (
		_w25599_,
		_w25600_,
		_w25733_
	);
	LUT2 #(
		.INIT('h8)
	) name15222 (
		_w25597_,
		_w25598_,
		_w25734_
	);
	LUT2 #(
		.INIT('h8)
	) name15223 (
		_w25595_,
		_w25596_,
		_w25735_
	);
	LUT2 #(
		.INIT('h8)
	) name15224 (
		_w25593_,
		_w25594_,
		_w25736_
	);
	LUT2 #(
		.INIT('h8)
	) name15225 (
		_w25591_,
		_w25592_,
		_w25737_
	);
	LUT2 #(
		.INIT('h8)
	) name15226 (
		_w25589_,
		_w25590_,
		_w25738_
	);
	LUT2 #(
		.INIT('h8)
	) name15227 (
		_w25587_,
		_w25588_,
		_w25739_
	);
	LUT2 #(
		.INIT('h8)
	) name15228 (
		_w25585_,
		_w25586_,
		_w25740_
	);
	LUT2 #(
		.INIT('h8)
	) name15229 (
		_w25583_,
		_w25584_,
		_w25741_
	);
	LUT2 #(
		.INIT('h8)
	) name15230 (
		_w25581_,
		_w25582_,
		_w25742_
	);
	LUT2 #(
		.INIT('h8)
	) name15231 (
		_w25579_,
		_w25580_,
		_w25743_
	);
	LUT2 #(
		.INIT('h8)
	) name15232 (
		_w25577_,
		_w25578_,
		_w25744_
	);
	LUT2 #(
		.INIT('h8)
	) name15233 (
		_w25575_,
		_w25576_,
		_w25745_
	);
	LUT2 #(
		.INIT('h8)
	) name15234 (
		_w25573_,
		_w25574_,
		_w25746_
	);
	LUT2 #(
		.INIT('h8)
	) name15235 (
		_w25571_,
		_w25572_,
		_w25747_
	);
	LUT2 #(
		.INIT('h8)
	) name15236 (
		_w25569_,
		_w25570_,
		_w25748_
	);
	LUT2 #(
		.INIT('h8)
	) name15237 (
		_w25567_,
		_w25568_,
		_w25749_
	);
	LUT2 #(
		.INIT('h8)
	) name15238 (
		_w25565_,
		_w25566_,
		_w25750_
	);
	LUT2 #(
		.INIT('h8)
	) name15239 (
		_w25563_,
		_w25564_,
		_w25751_
	);
	LUT2 #(
		.INIT('h8)
	) name15240 (
		_w25561_,
		_w25562_,
		_w25752_
	);
	LUT2 #(
		.INIT('h8)
	) name15241 (
		_w25751_,
		_w25752_,
		_w25753_
	);
	LUT2 #(
		.INIT('h8)
	) name15242 (
		_w25749_,
		_w25750_,
		_w25754_
	);
	LUT2 #(
		.INIT('h8)
	) name15243 (
		_w25747_,
		_w25748_,
		_w25755_
	);
	LUT2 #(
		.INIT('h8)
	) name15244 (
		_w25745_,
		_w25746_,
		_w25756_
	);
	LUT2 #(
		.INIT('h8)
	) name15245 (
		_w25743_,
		_w25744_,
		_w25757_
	);
	LUT2 #(
		.INIT('h8)
	) name15246 (
		_w25741_,
		_w25742_,
		_w25758_
	);
	LUT2 #(
		.INIT('h8)
	) name15247 (
		_w25739_,
		_w25740_,
		_w25759_
	);
	LUT2 #(
		.INIT('h8)
	) name15248 (
		_w25737_,
		_w25738_,
		_w25760_
	);
	LUT2 #(
		.INIT('h8)
	) name15249 (
		_w25735_,
		_w25736_,
		_w25761_
	);
	LUT2 #(
		.INIT('h8)
	) name15250 (
		_w25733_,
		_w25734_,
		_w25762_
	);
	LUT2 #(
		.INIT('h8)
	) name15251 (
		_w25731_,
		_w25732_,
		_w25763_
	);
	LUT2 #(
		.INIT('h8)
	) name15252 (
		_w25729_,
		_w25730_,
		_w25764_
	);
	LUT2 #(
		.INIT('h8)
	) name15253 (
		_w25727_,
		_w25728_,
		_w25765_
	);
	LUT2 #(
		.INIT('h8)
	) name15254 (
		_w25725_,
		_w25726_,
		_w25766_
	);
	LUT2 #(
		.INIT('h8)
	) name15255 (
		_w25723_,
		_w25724_,
		_w25767_
	);
	LUT2 #(
		.INIT('h8)
	) name15256 (
		_w25721_,
		_w25722_,
		_w25768_
	);
	LUT2 #(
		.INIT('h8)
	) name15257 (
		_w25719_,
		_w25720_,
		_w25769_
	);
	LUT2 #(
		.INIT('h8)
	) name15258 (
		_w25717_,
		_w25718_,
		_w25770_
	);
	LUT2 #(
		.INIT('h8)
	) name15259 (
		_w25715_,
		_w25716_,
		_w25771_
	);
	LUT2 #(
		.INIT('h8)
	) name15260 (
		_w25713_,
		_w25714_,
		_w25772_
	);
	LUT2 #(
		.INIT('h8)
	) name15261 (
		_w25711_,
		_w25712_,
		_w25773_
	);
	LUT2 #(
		.INIT('h8)
	) name15262 (
		_w25709_,
		_w25710_,
		_w25774_
	);
	LUT2 #(
		.INIT('h8)
	) name15263 (
		_w25707_,
		_w25708_,
		_w25775_
	);
	LUT2 #(
		.INIT('h8)
	) name15264 (
		_w25705_,
		_w25706_,
		_w25776_
	);
	LUT2 #(
		.INIT('h8)
	) name15265 (
		_w25703_,
		_w25704_,
		_w25777_
	);
	LUT2 #(
		.INIT('h8)
	) name15266 (
		_w25701_,
		_w25702_,
		_w25778_
	);
	LUT2 #(
		.INIT('h8)
	) name15267 (
		_w25699_,
		_w25700_,
		_w25779_
	);
	LUT2 #(
		.INIT('h8)
	) name15268 (
		_w25697_,
		_w25698_,
		_w25780_
	);
	LUT2 #(
		.INIT('h8)
	) name15269 (
		_w25695_,
		_w25696_,
		_w25781_
	);
	LUT2 #(
		.INIT('h8)
	) name15270 (
		_w25693_,
		_w25694_,
		_w25782_
	);
	LUT2 #(
		.INIT('h8)
	) name15271 (
		_w25691_,
		_w25692_,
		_w25783_
	);
	LUT2 #(
		.INIT('h8)
	) name15272 (
		_w25689_,
		_w25690_,
		_w25784_
	);
	LUT2 #(
		.INIT('h8)
	) name15273 (
		_w25783_,
		_w25784_,
		_w25785_
	);
	LUT2 #(
		.INIT('h8)
	) name15274 (
		_w25781_,
		_w25782_,
		_w25786_
	);
	LUT2 #(
		.INIT('h8)
	) name15275 (
		_w25779_,
		_w25780_,
		_w25787_
	);
	LUT2 #(
		.INIT('h8)
	) name15276 (
		_w25777_,
		_w25778_,
		_w25788_
	);
	LUT2 #(
		.INIT('h8)
	) name15277 (
		_w25775_,
		_w25776_,
		_w25789_
	);
	LUT2 #(
		.INIT('h8)
	) name15278 (
		_w25773_,
		_w25774_,
		_w25790_
	);
	LUT2 #(
		.INIT('h8)
	) name15279 (
		_w25771_,
		_w25772_,
		_w25791_
	);
	LUT2 #(
		.INIT('h8)
	) name15280 (
		_w25769_,
		_w25770_,
		_w25792_
	);
	LUT2 #(
		.INIT('h8)
	) name15281 (
		_w25767_,
		_w25768_,
		_w25793_
	);
	LUT2 #(
		.INIT('h8)
	) name15282 (
		_w25765_,
		_w25766_,
		_w25794_
	);
	LUT2 #(
		.INIT('h8)
	) name15283 (
		_w25763_,
		_w25764_,
		_w25795_
	);
	LUT2 #(
		.INIT('h8)
	) name15284 (
		_w25761_,
		_w25762_,
		_w25796_
	);
	LUT2 #(
		.INIT('h8)
	) name15285 (
		_w25759_,
		_w25760_,
		_w25797_
	);
	LUT2 #(
		.INIT('h8)
	) name15286 (
		_w25757_,
		_w25758_,
		_w25798_
	);
	LUT2 #(
		.INIT('h8)
	) name15287 (
		_w25755_,
		_w25756_,
		_w25799_
	);
	LUT2 #(
		.INIT('h8)
	) name15288 (
		_w25753_,
		_w25754_,
		_w25800_
	);
	LUT2 #(
		.INIT('h8)
	) name15289 (
		_w25799_,
		_w25800_,
		_w25801_
	);
	LUT2 #(
		.INIT('h8)
	) name15290 (
		_w25797_,
		_w25798_,
		_w25802_
	);
	LUT2 #(
		.INIT('h8)
	) name15291 (
		_w25795_,
		_w25796_,
		_w25803_
	);
	LUT2 #(
		.INIT('h8)
	) name15292 (
		_w25793_,
		_w25794_,
		_w25804_
	);
	LUT2 #(
		.INIT('h8)
	) name15293 (
		_w25791_,
		_w25792_,
		_w25805_
	);
	LUT2 #(
		.INIT('h8)
	) name15294 (
		_w25789_,
		_w25790_,
		_w25806_
	);
	LUT2 #(
		.INIT('h8)
	) name15295 (
		_w25787_,
		_w25788_,
		_w25807_
	);
	LUT2 #(
		.INIT('h8)
	) name15296 (
		_w25785_,
		_w25786_,
		_w25808_
	);
	LUT2 #(
		.INIT('h8)
	) name15297 (
		_w25807_,
		_w25808_,
		_w25809_
	);
	LUT2 #(
		.INIT('h8)
	) name15298 (
		_w25805_,
		_w25806_,
		_w25810_
	);
	LUT2 #(
		.INIT('h8)
	) name15299 (
		_w25803_,
		_w25804_,
		_w25811_
	);
	LUT2 #(
		.INIT('h8)
	) name15300 (
		_w25801_,
		_w25802_,
		_w25812_
	);
	LUT2 #(
		.INIT('h8)
	) name15301 (
		_w25811_,
		_w25812_,
		_w25813_
	);
	LUT2 #(
		.INIT('h8)
	) name15302 (
		_w25809_,
		_w25810_,
		_w25814_
	);
	LUT2 #(
		.INIT('h8)
	) name15303 (
		_w25813_,
		_w25814_,
		_w25815_
	);
	LUT2 #(
		.INIT('h1)
	) name15304 (
		wb_rst_i_pad,
		_w25815_,
		_w25816_
	);
	LUT2 #(
		.INIT('h1)
	) name15305 (
		_w22944_,
		_w25816_,
		_w25817_
	);
	LUT2 #(
		.INIT('h8)
	) name15306 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 ,
		_w23522_,
		_w25818_
	);
	LUT2 #(
		.INIT('h8)
	) name15307 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		_w23501_,
		_w25819_
	);
	LUT2 #(
		.INIT('h8)
	) name15308 (
		\ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 ,
		_w22956_,
		_w25820_
	);
	LUT2 #(
		.INIT('h8)
	) name15309 (
		\ethreg1_IPGR1_0_DataOut_reg[5]/NET0131 ,
		_w24710_,
		_w25821_
	);
	LUT2 #(
		.INIT('h8)
	) name15310 (
		\ethreg1_MODER_0_DataOut_reg[5]/NET0131 ,
		_w23519_,
		_w25822_
	);
	LUT2 #(
		.INIT('h8)
	) name15311 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		_w22959_,
		_w25823_
	);
	LUT2 #(
		.INIT('h8)
	) name15312 (
		\ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 ,
		_w23499_,
		_w25824_
	);
	LUT2 #(
		.INIT('h8)
	) name15313 (
		\ethreg1_IPGR2_0_DataOut_reg[5]/NET0131 ,
		_w24724_,
		_w25825_
	);
	LUT2 #(
		.INIT('h8)
	) name15314 (
		\ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 ,
		_w22952_,
		_w25826_
	);
	LUT2 #(
		.INIT('h8)
	) name15315 (
		\ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 ,
		_w24722_,
		_w25827_
	);
	LUT2 #(
		.INIT('h8)
	) name15316 (
		\ethreg1_IPGT_0_DataOut_reg[5]/NET0131 ,
		_w24717_,
		_w25828_
	);
	LUT2 #(
		.INIT('h8)
	) name15317 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		_w24713_,
		_w25829_
	);
	LUT2 #(
		.INIT('h8)
	) name15318 (
		\ethreg1_irq_txc_reg/NET0131 ,
		_w24707_,
		_w25830_
	);
	LUT2 #(
		.INIT('h8)
	) name15319 (
		\ethreg1_PACKETLEN_0_DataOut_reg[5]/NET0131 ,
		_w22966_,
		_w25831_
	);
	LUT2 #(
		.INIT('h8)
	) name15320 (
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w24726_,
		_w25832_
	);
	LUT2 #(
		.INIT('h8)
	) name15321 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		_w24730_,
		_w25833_
	);
	LUT2 #(
		.INIT('h8)
	) name15322 (
		\ethreg1_MIIRX_DATA_DataOut_reg[5]/NET0131 ,
		_w23507_,
		_w25834_
	);
	LUT2 #(
		.INIT('h1)
	) name15323 (
		_w25818_,
		_w25819_,
		_w25835_
	);
	LUT2 #(
		.INIT('h1)
	) name15324 (
		_w25820_,
		_w25821_,
		_w25836_
	);
	LUT2 #(
		.INIT('h1)
	) name15325 (
		_w25822_,
		_w25823_,
		_w25837_
	);
	LUT2 #(
		.INIT('h1)
	) name15326 (
		_w25824_,
		_w25825_,
		_w25838_
	);
	LUT2 #(
		.INIT('h1)
	) name15327 (
		_w25826_,
		_w25827_,
		_w25839_
	);
	LUT2 #(
		.INIT('h1)
	) name15328 (
		_w25828_,
		_w25829_,
		_w25840_
	);
	LUT2 #(
		.INIT('h1)
	) name15329 (
		_w25830_,
		_w25832_,
		_w25841_
	);
	LUT2 #(
		.INIT('h4)
	) name15330 (
		_w25834_,
		_w25841_,
		_w25842_
	);
	LUT2 #(
		.INIT('h8)
	) name15331 (
		_w25839_,
		_w25840_,
		_w25843_
	);
	LUT2 #(
		.INIT('h8)
	) name15332 (
		_w25837_,
		_w25838_,
		_w25844_
	);
	LUT2 #(
		.INIT('h8)
	) name15333 (
		_w25835_,
		_w25836_,
		_w25845_
	);
	LUT2 #(
		.INIT('h8)
	) name15334 (
		_w22944_,
		_w25845_,
		_w25846_
	);
	LUT2 #(
		.INIT('h8)
	) name15335 (
		_w25843_,
		_w25844_,
		_w25847_
	);
	LUT2 #(
		.INIT('h4)
	) name15336 (
		_w25831_,
		_w25842_,
		_w25848_
	);
	LUT2 #(
		.INIT('h4)
	) name15337 (
		_w25833_,
		_w25848_,
		_w25849_
	);
	LUT2 #(
		.INIT('h8)
	) name15338 (
		_w25846_,
		_w25847_,
		_w25850_
	);
	LUT2 #(
		.INIT('h8)
	) name15339 (
		_w25849_,
		_w25850_,
		_w25851_
	);
	LUT2 #(
		.INIT('h1)
	) name15340 (
		_w25817_,
		_w25851_,
		_w25852_
	);
	LUT2 #(
		.INIT('h8)
	) name15341 (
		\wishbone_bd_ram_mem0_reg[8][7]/P0001 ,
		_w12920_,
		_w25853_
	);
	LUT2 #(
		.INIT('h8)
	) name15342 (
		\wishbone_bd_ram_mem0_reg[80][7]/P0001 ,
		_w12689_,
		_w25854_
	);
	LUT2 #(
		.INIT('h8)
	) name15343 (
		\wishbone_bd_ram_mem0_reg[230][7]/P0001 ,
		_w13036_,
		_w25855_
	);
	LUT2 #(
		.INIT('h8)
	) name15344 (
		\wishbone_bd_ram_mem0_reg[64][7]/P0001 ,
		_w12976_,
		_w25856_
	);
	LUT2 #(
		.INIT('h8)
	) name15345 (
		\wishbone_bd_ram_mem0_reg[57][7]/P0001 ,
		_w13116_,
		_w25857_
	);
	LUT2 #(
		.INIT('h8)
	) name15346 (
		\wishbone_bd_ram_mem0_reg[179][7]/P0001 ,
		_w13050_,
		_w25858_
	);
	LUT2 #(
		.INIT('h8)
	) name15347 (
		\wishbone_bd_ram_mem0_reg[42][7]/P0001 ,
		_w12842_,
		_w25859_
	);
	LUT2 #(
		.INIT('h8)
	) name15348 (
		\wishbone_bd_ram_mem0_reg[31][7]/P0001 ,
		_w13198_,
		_w25860_
	);
	LUT2 #(
		.INIT('h8)
	) name15349 (
		\wishbone_bd_ram_mem0_reg[107][7]/P0001 ,
		_w12749_,
		_w25861_
	);
	LUT2 #(
		.INIT('h8)
	) name15350 (
		\wishbone_bd_ram_mem0_reg[246][7]/P0001 ,
		_w13076_,
		_w25862_
	);
	LUT2 #(
		.INIT('h8)
	) name15351 (
		\wishbone_bd_ram_mem0_reg[77][7]/P0001 ,
		_w12982_,
		_w25863_
	);
	LUT2 #(
		.INIT('h8)
	) name15352 (
		\wishbone_bd_ram_mem0_reg[109][7]/P0001 ,
		_w12888_,
		_w25864_
	);
	LUT2 #(
		.INIT('h8)
	) name15353 (
		\wishbone_bd_ram_mem0_reg[16][7]/P0001 ,
		_w13140_,
		_w25865_
	);
	LUT2 #(
		.INIT('h8)
	) name15354 (
		\wishbone_bd_ram_mem0_reg[219][7]/P0001 ,
		_w12806_,
		_w25866_
	);
	LUT2 #(
		.INIT('h8)
	) name15355 (
		\wishbone_bd_ram_mem0_reg[38][7]/P0001 ,
		_w13182_,
		_w25867_
	);
	LUT2 #(
		.INIT('h8)
	) name15356 (
		\wishbone_bd_ram_mem0_reg[23][7]/P0001 ,
		_w13008_,
		_w25868_
	);
	LUT2 #(
		.INIT('h8)
	) name15357 (
		\wishbone_bd_ram_mem0_reg[255][7]/P0001 ,
		_w13072_,
		_w25869_
	);
	LUT2 #(
		.INIT('h8)
	) name15358 (
		\wishbone_bd_ram_mem0_reg[237][7]/P0001 ,
		_w12990_,
		_w25870_
	);
	LUT2 #(
		.INIT('h8)
	) name15359 (
		\wishbone_bd_ram_mem0_reg[128][7]/P0001 ,
		_w12793_,
		_w25871_
	);
	LUT2 #(
		.INIT('h8)
	) name15360 (
		\wishbone_bd_ram_mem0_reg[5][7]/P0001 ,
		_w12878_,
		_w25872_
	);
	LUT2 #(
		.INIT('h8)
	) name15361 (
		\wishbone_bd_ram_mem0_reg[61][7]/P0001 ,
		_w12725_,
		_w25873_
	);
	LUT2 #(
		.INIT('h8)
	) name15362 (
		\wishbone_bd_ram_mem0_reg[124][7]/P0001 ,
		_w13058_,
		_w25874_
	);
	LUT2 #(
		.INIT('h8)
	) name15363 (
		\wishbone_bd_ram_mem0_reg[247][7]/P0001 ,
		_w12818_,
		_w25875_
	);
	LUT2 #(
		.INIT('h8)
	) name15364 (
		\wishbone_bd_ram_mem0_reg[212][7]/P0001 ,
		_w12796_,
		_w25876_
	);
	LUT2 #(
		.INIT('h8)
	) name15365 (
		\wishbone_bd_ram_mem0_reg[70][7]/P0001 ,
		_w12840_,
		_w25877_
	);
	LUT2 #(
		.INIT('h8)
	) name15366 (
		\wishbone_bd_ram_mem0_reg[141][7]/P0001 ,
		_w13004_,
		_w25878_
	);
	LUT2 #(
		.INIT('h8)
	) name15367 (
		\wishbone_bd_ram_mem0_reg[108][7]/P0001 ,
		_w13156_,
		_w25879_
	);
	LUT2 #(
		.INIT('h8)
	) name15368 (
		\wishbone_bd_ram_mem0_reg[186][7]/P0001 ,
		_w12783_,
		_w25880_
	);
	LUT2 #(
		.INIT('h8)
	) name15369 (
		\wishbone_bd_ram_mem0_reg[196][7]/P0001 ,
		_w13090_,
		_w25881_
	);
	LUT2 #(
		.INIT('h8)
	) name15370 (
		\wishbone_bd_ram_mem0_reg[82][7]/P0001 ,
		_w12942_,
		_w25882_
	);
	LUT2 #(
		.INIT('h8)
	) name15371 (
		\wishbone_bd_ram_mem0_reg[253][7]/P0001 ,
		_w13100_,
		_w25883_
	);
	LUT2 #(
		.INIT('h8)
	) name15372 (
		\wishbone_bd_ram_mem0_reg[211][7]/P0001 ,
		_w13166_,
		_w25884_
	);
	LUT2 #(
		.INIT('h8)
	) name15373 (
		\wishbone_bd_ram_mem0_reg[150][7]/P0001 ,
		_w13136_,
		_w25885_
	);
	LUT2 #(
		.INIT('h8)
	) name15374 (
		\wishbone_bd_ram_mem0_reg[245][7]/P0001 ,
		_w13022_,
		_w25886_
	);
	LUT2 #(
		.INIT('h8)
	) name15375 (
		\wishbone_bd_ram_mem0_reg[74][7]/P0001 ,
		_w12812_,
		_w25887_
	);
	LUT2 #(
		.INIT('h8)
	) name15376 (
		\wishbone_bd_ram_mem0_reg[138][7]/P0001 ,
		_w12958_,
		_w25888_
	);
	LUT2 #(
		.INIT('h8)
	) name15377 (
		\wishbone_bd_ram_mem0_reg[3][7]/P0001 ,
		_w12866_,
		_w25889_
	);
	LUT2 #(
		.INIT('h8)
	) name15378 (
		\wishbone_bd_ram_mem0_reg[10][7]/P0001 ,
		_w13172_,
		_w25890_
	);
	LUT2 #(
		.INIT('h8)
	) name15379 (
		\wishbone_bd_ram_mem0_reg[198][7]/P0001 ,
		_w12832_,
		_w25891_
	);
	LUT2 #(
		.INIT('h8)
	) name15380 (
		\wishbone_bd_ram_mem0_reg[232][7]/P0001 ,
		_w12758_,
		_w25892_
	);
	LUT2 #(
		.INIT('h8)
	) name15381 (
		\wishbone_bd_ram_mem0_reg[120][7]/P0001 ,
		_w12707_,
		_w25893_
	);
	LUT2 #(
		.INIT('h8)
	) name15382 (
		\wishbone_bd_ram_mem0_reg[206][7]/P0001 ,
		_w12954_,
		_w25894_
	);
	LUT2 #(
		.INIT('h8)
	) name15383 (
		\wishbone_bd_ram_mem0_reg[13][7]/P0001 ,
		_w13178_,
		_w25895_
	);
	LUT2 #(
		.INIT('h8)
	) name15384 (
		\wishbone_bd_ram_mem0_reg[119][7]/P0001 ,
		_w13048_,
		_w25896_
	);
	LUT2 #(
		.INIT('h8)
	) name15385 (
		\wishbone_bd_ram_mem0_reg[224][7]/P0001 ,
		_w12902_,
		_w25897_
	);
	LUT2 #(
		.INIT('h8)
	) name15386 (
		\wishbone_bd_ram_mem0_reg[152][7]/P0001 ,
		_w12966_,
		_w25898_
	);
	LUT2 #(
		.INIT('h8)
	) name15387 (
		\wishbone_bd_ram_mem0_reg[35][7]/P0001 ,
		_w12703_,
		_w25899_
	);
	LUT2 #(
		.INIT('h8)
	) name15388 (
		\wishbone_bd_ram_mem0_reg[238][7]/P0001 ,
		_w13160_,
		_w25900_
	);
	LUT2 #(
		.INIT('h8)
	) name15389 (
		\wishbone_bd_ram_mem0_reg[191][7]/P0001 ,
		_w13034_,
		_w25901_
	);
	LUT2 #(
		.INIT('h8)
	) name15390 (
		\wishbone_bd_ram_mem0_reg[92][7]/P0001 ,
		_w13010_,
		_w25902_
	);
	LUT2 #(
		.INIT('h8)
	) name15391 (
		\wishbone_bd_ram_mem0_reg[30][7]/P0001 ,
		_w13104_,
		_w25903_
	);
	LUT2 #(
		.INIT('h8)
	) name15392 (
		\wishbone_bd_ram_mem0_reg[26][7]/P0001 ,
		_w12699_,
		_w25904_
	);
	LUT2 #(
		.INIT('h8)
	) name15393 (
		\wishbone_bd_ram_mem0_reg[7][7]/P0001 ,
		_w12728_,
		_w25905_
	);
	LUT2 #(
		.INIT('h8)
	) name15394 (
		\wishbone_bd_ram_mem0_reg[158][7]/P0001 ,
		_w12898_,
		_w25906_
	);
	LUT2 #(
		.INIT('h8)
	) name15395 (
		\wishbone_bd_ram_mem0_reg[102][7]/P0001 ,
		_w12685_,
		_w25907_
	);
	LUT2 #(
		.INIT('h8)
	) name15396 (
		\wishbone_bd_ram_mem0_reg[114][7]/P0001 ,
		_w13202_,
		_w25908_
	);
	LUT2 #(
		.INIT('h8)
	) name15397 (
		\wishbone_bd_ram_mem0_reg[151][7]/P0001 ,
		_w13142_,
		_w25909_
	);
	LUT2 #(
		.INIT('h8)
	) name15398 (
		\wishbone_bd_ram_mem0_reg[227][7]/P0001 ,
		_w12936_,
		_w25910_
	);
	LUT2 #(
		.INIT('h8)
	) name15399 (
		\wishbone_bd_ram_mem0_reg[122][7]/P0001 ,
		_w13130_,
		_w25911_
	);
	LUT2 #(
		.INIT('h8)
	) name15400 (
		\wishbone_bd_ram_mem0_reg[117][7]/P0001 ,
		_w12715_,
		_w25912_
	);
	LUT2 #(
		.INIT('h8)
	) name15401 (
		\wishbone_bd_ram_mem0_reg[221][7]/P0001 ,
		_w12802_,
		_w25913_
	);
	LUT2 #(
		.INIT('h8)
	) name15402 (
		\wishbone_bd_ram_mem0_reg[131][7]/P0001 ,
		_w12852_,
		_w25914_
	);
	LUT2 #(
		.INIT('h8)
	) name15403 (
		\wishbone_bd_ram_mem0_reg[210][7]/P0001 ,
		_w12924_,
		_w25915_
	);
	LUT2 #(
		.INIT('h8)
	) name15404 (
		\wishbone_bd_ram_mem0_reg[223][7]/P0001 ,
		_w12838_,
		_w25916_
	);
	LUT2 #(
		.INIT('h8)
	) name15405 (
		\wishbone_bd_ram_mem0_reg[176][7]/P0001 ,
		_w12868_,
		_w25917_
	);
	LUT2 #(
		.INIT('h8)
	) name15406 (
		\wishbone_bd_ram_mem0_reg[235][7]/P0001 ,
		_w12696_,
		_w25918_
	);
	LUT2 #(
		.INIT('h8)
	) name15407 (
		\wishbone_bd_ram_mem0_reg[163][7]/P0001 ,
		_w12882_,
		_w25919_
	);
	LUT2 #(
		.INIT('h8)
	) name15408 (
		\wishbone_bd_ram_mem0_reg[9][7]/P0001 ,
		_w12808_,
		_w25920_
	);
	LUT2 #(
		.INIT('h8)
	) name15409 (
		\wishbone_bd_ram_mem0_reg[156][7]/P0001 ,
		_w13190_,
		_w25921_
	);
	LUT2 #(
		.INIT('h8)
	) name15410 (
		\wishbone_bd_ram_mem0_reg[153][7]/P0001 ,
		_w12890_,
		_w25922_
	);
	LUT2 #(
		.INIT('h8)
	) name15411 (
		\wishbone_bd_ram_mem0_reg[44][7]/P0001 ,
		_w12896_,
		_w25923_
	);
	LUT2 #(
		.INIT('h8)
	) name15412 (
		\wishbone_bd_ram_mem0_reg[59][7]/P0001 ,
		_w12780_,
		_w25924_
	);
	LUT2 #(
		.INIT('h8)
	) name15413 (
		\wishbone_bd_ram_mem0_reg[17][7]/P0001 ,
		_w12848_,
		_w25925_
	);
	LUT2 #(
		.INIT('h8)
	) name15414 (
		\wishbone_bd_ram_mem0_reg[170][7]/P0001 ,
		_w13030_,
		_w25926_
	);
	LUT2 #(
		.INIT('h8)
	) name15415 (
		\wishbone_bd_ram_mem0_reg[192][7]/P0001 ,
		_w12938_,
		_w25927_
	);
	LUT2 #(
		.INIT('h8)
	) name15416 (
		\wishbone_bd_ram_mem0_reg[207][7]/P0001 ,
		_w13180_,
		_w25928_
	);
	LUT2 #(
		.INIT('h8)
	) name15417 (
		\wishbone_bd_ram_mem0_reg[166][7]/P0001 ,
		_w13040_,
		_w25929_
	);
	LUT2 #(
		.INIT('h8)
	) name15418 (
		\wishbone_bd_ram_mem0_reg[251][7]/P0001 ,
		_w13054_,
		_w25930_
	);
	LUT2 #(
		.INIT('h8)
	) name15419 (
		\wishbone_bd_ram_mem0_reg[178][7]/P0001 ,
		_w12886_,
		_w25931_
	);
	LUT2 #(
		.INIT('h8)
	) name15420 (
		\wishbone_bd_ram_mem0_reg[37][7]/P0001 ,
		_w13102_,
		_w25932_
	);
	LUT2 #(
		.INIT('h8)
	) name15421 (
		\wishbone_bd_ram_mem0_reg[222][7]/P0001 ,
		_w13094_,
		_w25933_
	);
	LUT2 #(
		.INIT('h8)
	) name15422 (
		\wishbone_bd_ram_mem0_reg[193][7]/P0001 ,
		_w13056_,
		_w25934_
	);
	LUT2 #(
		.INIT('h8)
	) name15423 (
		\wishbone_bd_ram_mem0_reg[85][7]/P0001 ,
		_w13216_,
		_w25935_
	);
	LUT2 #(
		.INIT('h8)
	) name15424 (
		\wishbone_bd_ram_mem0_reg[242][7]/P0001 ,
		_w12932_,
		_w25936_
	);
	LUT2 #(
		.INIT('h8)
	) name15425 (
		\wishbone_bd_ram_mem0_reg[49][7]/P0001 ,
		_w12994_,
		_w25937_
	);
	LUT2 #(
		.INIT('h8)
	) name15426 (
		\wishbone_bd_ram_mem0_reg[69][7]/P0001 ,
		_w12738_,
		_w25938_
	);
	LUT2 #(
		.INIT('h8)
	) name15427 (
		\wishbone_bd_ram_mem0_reg[21][7]/P0001 ,
		_w12906_,
		_w25939_
	);
	LUT2 #(
		.INIT('h8)
	) name15428 (
		\wishbone_bd_ram_mem0_reg[105][7]/P0001 ,
		_w12751_,
		_w25940_
	);
	LUT2 #(
		.INIT('h8)
	) name15429 (
		\wishbone_bd_ram_mem0_reg[116][7]/P0001 ,
		_w12998_,
		_w25941_
	);
	LUT2 #(
		.INIT('h8)
	) name15430 (
		\wishbone_bd_ram_mem0_reg[248][7]/P0001 ,
		_w12789_,
		_w25942_
	);
	LUT2 #(
		.INIT('h8)
	) name15431 (
		\wishbone_bd_ram_mem0_reg[28][7]/P0001 ,
		_w13170_,
		_w25943_
	);
	LUT2 #(
		.INIT('h8)
	) name15432 (
		\wishbone_bd_ram_mem0_reg[144][7]/P0001 ,
		_w12756_,
		_w25944_
	);
	LUT2 #(
		.INIT('h8)
	) name15433 (
		\wishbone_bd_ram_mem0_reg[240][7]/P0001 ,
		_w12864_,
		_w25945_
	);
	LUT2 #(
		.INIT('h8)
	) name15434 (
		\wishbone_bd_ram_mem0_reg[183][7]/P0001 ,
		_w12787_,
		_w25946_
	);
	LUT2 #(
		.INIT('h8)
	) name15435 (
		\wishbone_bd_ram_mem0_reg[118][7]/P0001 ,
		_w12830_,
		_w25947_
	);
	LUT2 #(
		.INIT('h8)
	) name15436 (
		\wishbone_bd_ram_mem0_reg[213][7]/P0001 ,
		_w13002_,
		_w25948_
	);
	LUT2 #(
		.INIT('h8)
	) name15437 (
		\wishbone_bd_ram_mem0_reg[91][7]/P0001 ,
		_w13074_,
		_w25949_
	);
	LUT2 #(
		.INIT('h8)
	) name15438 (
		\wishbone_bd_ram_mem0_reg[72][7]/P0001 ,
		_w12810_,
		_w25950_
	);
	LUT2 #(
		.INIT('h8)
	) name15439 (
		\wishbone_bd_ram_mem0_reg[149][7]/P0001 ,
		_w12741_,
		_w25951_
	);
	LUT2 #(
		.INIT('h8)
	) name15440 (
		\wishbone_bd_ram_mem0_reg[24][7]/P0001 ,
		_w13084_,
		_w25952_
	);
	LUT2 #(
		.INIT('h8)
	) name15441 (
		\wishbone_bd_ram_mem0_reg[218][7]/P0001 ,
		_w13206_,
		_w25953_
	);
	LUT2 #(
		.INIT('h8)
	) name15442 (
		\wishbone_bd_ram_mem0_reg[130][7]/P0001 ,
		_w12914_,
		_w25954_
	);
	LUT2 #(
		.INIT('h8)
	) name15443 (
		\wishbone_bd_ram_mem0_reg[79][7]/P0001 ,
		_w13212_,
		_w25955_
	);
	LUT2 #(
		.INIT('h8)
	) name15444 (
		\wishbone_bd_ram_mem0_reg[189][7]/P0001 ,
		_w13042_,
		_w25956_
	);
	LUT2 #(
		.INIT('h8)
	) name15445 (
		\wishbone_bd_ram_mem0_reg[172][7]/P0001 ,
		_w12944_,
		_w25957_
	);
	LUT2 #(
		.INIT('h8)
	) name15446 (
		\wishbone_bd_ram_mem0_reg[55][7]/P0001 ,
		_w12785_,
		_w25958_
	);
	LUT2 #(
		.INIT('h8)
	) name15447 (
		\wishbone_bd_ram_mem0_reg[95][7]/P0001 ,
		_w12844_,
		_w25959_
	);
	LUT2 #(
		.INIT('h8)
	) name15448 (
		\wishbone_bd_ram_mem0_reg[180][7]/P0001 ,
		_w12791_,
		_w25960_
	);
	LUT2 #(
		.INIT('h8)
	) name15449 (
		\wishbone_bd_ram_mem0_reg[22][7]/P0001 ,
		_w13110_,
		_w25961_
	);
	LUT2 #(
		.INIT('h8)
	) name15450 (
		\wishbone_bd_ram_mem0_reg[34][7]/P0001 ,
		_w12930_,
		_w25962_
	);
	LUT2 #(
		.INIT('h8)
	) name15451 (
		\wishbone_bd_ram_mem0_reg[136][7]/P0001 ,
		_w13064_,
		_w25963_
	);
	LUT2 #(
		.INIT('h8)
	) name15452 (
		\wishbone_bd_ram_mem0_reg[39][7]/P0001 ,
		_w13018_,
		_w25964_
	);
	LUT2 #(
		.INIT('h8)
	) name15453 (
		\wishbone_bd_ram_mem0_reg[161][7]/P0001 ,
		_w12754_,
		_w25965_
	);
	LUT2 #(
		.INIT('h8)
	) name15454 (
		\wishbone_bd_ram_mem0_reg[173][7]/P0001 ,
		_w12854_,
		_w25966_
	);
	LUT2 #(
		.INIT('h8)
	) name15455 (
		\wishbone_bd_ram_mem0_reg[233][7]/P0001 ,
		_w12836_,
		_w25967_
	);
	LUT2 #(
		.INIT('h8)
	) name15456 (
		\wishbone_bd_ram_mem0_reg[98][7]/P0001 ,
		_w12816_,
		_w25968_
	);
	LUT2 #(
		.INIT('h8)
	) name15457 (
		\wishbone_bd_ram_mem0_reg[244][7]/P0001 ,
		_w12747_,
		_w25969_
	);
	LUT2 #(
		.INIT('h8)
	) name15458 (
		\wishbone_bd_ram_mem0_reg[101][7]/P0001 ,
		_w13192_,
		_w25970_
	);
	LUT2 #(
		.INIT('h8)
	) name15459 (
		\wishbone_bd_ram_mem0_reg[169][7]/P0001 ,
		_w12722_,
		_w25971_
	);
	LUT2 #(
		.INIT('h8)
	) name15460 (
		\wishbone_bd_ram_mem0_reg[104][7]/P0001 ,
		_w13148_,
		_w25972_
	);
	LUT2 #(
		.INIT('h8)
	) name15461 (
		\wishbone_bd_ram_mem0_reg[112][7]/P0001 ,
		_w12733_,
		_w25973_
	);
	LUT2 #(
		.INIT('h8)
	) name15462 (
		\wishbone_bd_ram_mem0_reg[252][7]/P0001 ,
		_w13080_,
		_w25974_
	);
	LUT2 #(
		.INIT('h8)
	) name15463 (
		\wishbone_bd_ram_mem0_reg[60][7]/P0001 ,
		_w13204_,
		_w25975_
	);
	LUT2 #(
		.INIT('h8)
	) name15464 (
		\wishbone_bd_ram_mem0_reg[181][7]/P0001 ,
		_w12828_,
		_w25976_
	);
	LUT2 #(
		.INIT('h8)
	) name15465 (
		\wishbone_bd_ram_mem0_reg[243][7]/P0001 ,
		_w12804_,
		_w25977_
	);
	LUT2 #(
		.INIT('h8)
	) name15466 (
		\wishbone_bd_ram_mem0_reg[19][7]/P0001 ,
		_w13012_,
		_w25978_
	);
	LUT2 #(
		.INIT('h8)
	) name15467 (
		\wishbone_bd_ram_mem0_reg[190][7]/P0001 ,
		_w12858_,
		_w25979_
	);
	LUT2 #(
		.INIT('h8)
	) name15468 (
		\wishbone_bd_ram_mem0_reg[188][7]/P0001 ,
		_w12948_,
		_w25980_
	);
	LUT2 #(
		.INIT('h8)
	) name15469 (
		\wishbone_bd_ram_mem0_reg[125][7]/P0001 ,
		_w12956_,
		_w25981_
	);
	LUT2 #(
		.INIT('h8)
	) name15470 (
		\wishbone_bd_ram_mem0_reg[54][7]/P0001 ,
		_w12770_,
		_w25982_
	);
	LUT2 #(
		.INIT('h8)
	) name15471 (
		\wishbone_bd_ram_mem0_reg[32][7]/P0001 ,
		_w13120_,
		_w25983_
	);
	LUT2 #(
		.INIT('h8)
	) name15472 (
		\wishbone_bd_ram_mem0_reg[96][7]/P0001 ,
		_w12912_,
		_w25984_
	);
	LUT2 #(
		.INIT('h8)
	) name15473 (
		\wishbone_bd_ram_mem0_reg[145][7]/P0001 ,
		_w13106_,
		_w25985_
	);
	LUT2 #(
		.INIT('h8)
	) name15474 (
		\wishbone_bd_ram_mem0_reg[11][7]/P0001 ,
		_w13194_,
		_w25986_
	);
	LUT2 #(
		.INIT('h8)
	) name15475 (
		\wishbone_bd_ram_mem0_reg[148][7]/P0001 ,
		_w13000_,
		_w25987_
	);
	LUT2 #(
		.INIT('h8)
	) name15476 (
		\wishbone_bd_ram_mem0_reg[121][7]/P0001 ,
		_w13078_,
		_w25988_
	);
	LUT2 #(
		.INIT('h8)
	) name15477 (
		\wishbone_bd_ram_mem0_reg[27][7]/P0001 ,
		_w12880_,
		_w25989_
	);
	LUT2 #(
		.INIT('h8)
	) name15478 (
		\wishbone_bd_ram_mem0_reg[164][7]/P0001 ,
		_w12876_,
		_w25990_
	);
	LUT2 #(
		.INIT('h8)
	) name15479 (
		\wishbone_bd_ram_mem0_reg[216][7]/P0001 ,
		_w13028_,
		_w25991_
	);
	LUT2 #(
		.INIT('h8)
	) name15480 (
		\wishbone_bd_ram_mem0_reg[168][7]/P0001 ,
		_w13208_,
		_w25992_
	);
	LUT2 #(
		.INIT('h8)
	) name15481 (
		\wishbone_bd_ram_mem0_reg[185][7]/P0001 ,
		_w12940_,
		_w25993_
	);
	LUT2 #(
		.INIT('h8)
	) name15482 (
		\wishbone_bd_ram_mem0_reg[241][7]/P0001 ,
		_w13006_,
		_w25994_
	);
	LUT2 #(
		.INIT('h8)
	) name15483 (
		\wishbone_bd_ram_mem0_reg[93][7]/P0001 ,
		_w13016_,
		_w25995_
	);
	LUT2 #(
		.INIT('h8)
	) name15484 (
		\wishbone_bd_ram_mem0_reg[58][7]/P0001 ,
		_w13070_,
		_w25996_
	);
	LUT2 #(
		.INIT('h8)
	) name15485 (
		\wishbone_bd_ram_mem0_reg[90][7]/P0001 ,
		_w12978_,
		_w25997_
	);
	LUT2 #(
		.INIT('h8)
	) name15486 (
		\wishbone_bd_ram_mem0_reg[100][7]/P0001 ,
		_w12960_,
		_w25998_
	);
	LUT2 #(
		.INIT('h8)
	) name15487 (
		\wishbone_bd_ram_mem0_reg[47][7]/P0001 ,
		_w12904_,
		_w25999_
	);
	LUT2 #(
		.INIT('h8)
	) name15488 (
		\wishbone_bd_ram_mem0_reg[249][7]/P0001 ,
		_w12900_,
		_w26000_
	);
	LUT2 #(
		.INIT('h8)
	) name15489 (
		\wishbone_bd_ram_mem0_reg[135][7]/P0001 ,
		_w13124_,
		_w26001_
	);
	LUT2 #(
		.INIT('h8)
	) name15490 (
		\wishbone_bd_ram_mem0_reg[111][7]/P0001 ,
		_w12744_,
		_w26002_
	);
	LUT2 #(
		.INIT('h8)
	) name15491 (
		\wishbone_bd_ram_mem0_reg[134][7]/P0001 ,
		_w12763_,
		_w26003_
	);
	LUT2 #(
		.INIT('h8)
	) name15492 (
		\wishbone_bd_ram_mem0_reg[165][7]/P0001 ,
		_w13044_,
		_w26004_
	);
	LUT2 #(
		.INIT('h8)
	) name15493 (
		\wishbone_bd_ram_mem0_reg[73][7]/P0001 ,
		_w12918_,
		_w26005_
	);
	LUT2 #(
		.INIT('h8)
	) name15494 (
		\wishbone_bd_ram_mem0_reg[4][7]/P0001 ,
		_w12666_,
		_w26006_
	);
	LUT2 #(
		.INIT('h8)
	) name15495 (
		\wishbone_bd_ram_mem0_reg[129][7]/P0001 ,
		_w12776_,
		_w26007_
	);
	LUT2 #(
		.INIT('h8)
	) name15496 (
		\wishbone_bd_ram_mem0_reg[56][7]/P0001 ,
		_w12778_,
		_w26008_
	);
	LUT2 #(
		.INIT('h8)
	) name15497 (
		\wishbone_bd_ram_mem0_reg[162][7]/P0001 ,
		_w13098_,
		_w26009_
	);
	LUT2 #(
		.INIT('h8)
	) name15498 (
		\wishbone_bd_ram_mem0_reg[225][7]/P0001 ,
		_w13092_,
		_w26010_
	);
	LUT2 #(
		.INIT('h8)
	) name15499 (
		\wishbone_bd_ram_mem0_reg[6][7]/P0001 ,
		_w12968_,
		_w26011_
	);
	LUT2 #(
		.INIT('h8)
	) name15500 (
		\wishbone_bd_ram_mem0_reg[220][7]/P0001 ,
		_w13066_,
		_w26012_
	);
	LUT2 #(
		.INIT('h8)
	) name15501 (
		\wishbone_bd_ram_mem0_reg[48][7]/P0001 ,
		_w12970_,
		_w26013_
	);
	LUT2 #(
		.INIT('h8)
	) name15502 (
		\wishbone_bd_ram_mem0_reg[43][7]/P0001 ,
		_w13200_,
		_w26014_
	);
	LUT2 #(
		.INIT('h8)
	) name15503 (
		\wishbone_bd_ram_mem0_reg[142][7]/P0001 ,
		_w12928_,
		_w26015_
	);
	LUT2 #(
		.INIT('h8)
	) name15504 (
		\wishbone_bd_ram_mem0_reg[199][7]/P0001 ,
		_w12768_,
		_w26016_
	);
	LUT2 #(
		.INIT('h8)
	) name15505 (
		\wishbone_bd_ram_mem0_reg[146][7]/P0001 ,
		_w13060_,
		_w26017_
	);
	LUT2 #(
		.INIT('h8)
	) name15506 (
		\wishbone_bd_ram_mem0_reg[45][7]/P0001 ,
		_w12908_,
		_w26018_
	);
	LUT2 #(
		.INIT('h8)
	) name15507 (
		\wishbone_bd_ram_mem0_reg[106][7]/P0001 ,
		_w12713_,
		_w26019_
	);
	LUT2 #(
		.INIT('h8)
	) name15508 (
		\wishbone_bd_ram_mem0_reg[177][7]/P0001 ,
		_w12996_,
		_w26020_
	);
	LUT2 #(
		.INIT('h8)
	) name15509 (
		\wishbone_bd_ram_mem0_reg[53][7]/P0001 ,
		_w13020_,
		_w26021_
	);
	LUT2 #(
		.INIT('h8)
	) name15510 (
		\wishbone_bd_ram_mem0_reg[154][7]/P0001 ,
		_w12962_,
		_w26022_
	);
	LUT2 #(
		.INIT('h8)
	) name15511 (
		\wishbone_bd_ram_mem0_reg[12][7]/P0001 ,
		_w13118_,
		_w26023_
	);
	LUT2 #(
		.INIT('h8)
	) name15512 (
		\wishbone_bd_ram_mem0_reg[236][7]/P0001 ,
		_w12731_,
		_w26024_
	);
	LUT2 #(
		.INIT('h8)
	) name15513 (
		\wishbone_bd_ram_mem0_reg[36][7]/P0001 ,
		_w12800_,
		_w26025_
	);
	LUT2 #(
		.INIT('h8)
	) name15514 (
		\wishbone_bd_ram_mem0_reg[194][7]/P0001 ,
		_w12772_,
		_w26026_
	);
	LUT2 #(
		.INIT('h8)
	) name15515 (
		\wishbone_bd_ram_mem0_reg[202][7]/P0001 ,
		_w12870_,
		_w26027_
	);
	LUT2 #(
		.INIT('h8)
	) name15516 (
		\wishbone_bd_ram_mem0_reg[71][7]/P0001 ,
		_w12798_,
		_w26028_
	);
	LUT2 #(
		.INIT('h8)
	) name15517 (
		\wishbone_bd_ram_mem0_reg[143][7]/P0001 ,
		_w12922_,
		_w26029_
	);
	LUT2 #(
		.INIT('h8)
	) name15518 (
		\wishbone_bd_ram_mem0_reg[110][7]/P0001 ,
		_w13046_,
		_w26030_
	);
	LUT2 #(
		.INIT('h8)
	) name15519 (
		\wishbone_bd_ram_mem0_reg[167][7]/P0001 ,
		_w12986_,
		_w26031_
	);
	LUT2 #(
		.INIT('h8)
	) name15520 (
		\wishbone_bd_ram_mem0_reg[200][7]/P0001 ,
		_w12988_,
		_w26032_
	);
	LUT2 #(
		.INIT('h8)
	) name15521 (
		\wishbone_bd_ram_mem0_reg[203][7]/P0001 ,
		_w13158_,
		_w26033_
	);
	LUT2 #(
		.INIT('h8)
	) name15522 (
		\wishbone_bd_ram_mem0_reg[68][7]/P0001 ,
		_w12946_,
		_w26034_
	);
	LUT2 #(
		.INIT('h8)
	) name15523 (
		\wishbone_bd_ram_mem0_reg[197][7]/P0001 ,
		_w12834_,
		_w26035_
	);
	LUT2 #(
		.INIT('h8)
	) name15524 (
		\wishbone_bd_ram_mem0_reg[228][7]/P0001 ,
		_w12765_,
		_w26036_
	);
	LUT2 #(
		.INIT('h8)
	) name15525 (
		\wishbone_bd_ram_mem0_reg[229][7]/P0001 ,
		_w12711_,
		_w26037_
	);
	LUT2 #(
		.INIT('h8)
	) name15526 (
		\wishbone_bd_ram_mem0_reg[86][7]/P0001 ,
		_w12735_,
		_w26038_
	);
	LUT2 #(
		.INIT('h8)
	) name15527 (
		\wishbone_bd_ram_mem0_reg[208][7]/P0001 ,
		_w13032_,
		_w26039_
	);
	LUT2 #(
		.INIT('h8)
	) name15528 (
		\wishbone_bd_ram_mem0_reg[67][7]/P0001 ,
		_w13134_,
		_w26040_
	);
	LUT2 #(
		.INIT('h8)
	) name15529 (
		\wishbone_bd_ram_mem0_reg[50][7]/P0001 ,
		_w13150_,
		_w26041_
	);
	LUT2 #(
		.INIT('h8)
	) name15530 (
		\wishbone_bd_ram_mem0_reg[97][7]/P0001 ,
		_w13096_,
		_w26042_
	);
	LUT2 #(
		.INIT('h8)
	) name15531 (
		\wishbone_bd_ram_mem0_reg[175][7]/P0001 ,
		_w13126_,
		_w26043_
	);
	LUT2 #(
		.INIT('h8)
	) name15532 (
		\wishbone_bd_ram_mem0_reg[195][7]/P0001 ,
		_w13144_,
		_w26044_
	);
	LUT2 #(
		.INIT('h8)
	) name15533 (
		\wishbone_bd_ram_mem0_reg[226][7]/P0001 ,
		_w13138_,
		_w26045_
	);
	LUT2 #(
		.INIT('h8)
	) name15534 (
		\wishbone_bd_ram_mem0_reg[215][7]/P0001 ,
		_w12974_,
		_w26046_
	);
	LUT2 #(
		.INIT('h8)
	) name15535 (
		\wishbone_bd_ram_mem0_reg[184][7]/P0001 ,
		_w13062_,
		_w26047_
	);
	LUT2 #(
		.INIT('h8)
	) name15536 (
		\wishbone_bd_ram_mem0_reg[83][7]/P0001 ,
		_w12916_,
		_w26048_
	);
	LUT2 #(
		.INIT('h8)
	) name15537 (
		\wishbone_bd_ram_mem0_reg[201][7]/P0001 ,
		_w12822_,
		_w26049_
	);
	LUT2 #(
		.INIT('h8)
	) name15538 (
		\wishbone_bd_ram_mem0_reg[33][7]/P0001 ,
		_w12980_,
		_w26050_
	);
	LUT2 #(
		.INIT('h8)
	) name15539 (
		\wishbone_bd_ram_mem0_reg[52][7]/P0001 ,
		_w13082_,
		_w26051_
	);
	LUT2 #(
		.INIT('h8)
	) name15540 (
		\wishbone_bd_ram_mem0_reg[78][7]/P0001 ,
		_w12874_,
		_w26052_
	);
	LUT2 #(
		.INIT('h8)
	) name15541 (
		\wishbone_bd_ram_mem0_reg[66][7]/P0001 ,
		_w12824_,
		_w26053_
	);
	LUT2 #(
		.INIT('h8)
	) name15542 (
		\wishbone_bd_ram_mem0_reg[46][7]/P0001 ,
		_w12884_,
		_w26054_
	);
	LUT2 #(
		.INIT('h8)
	) name15543 (
		\wishbone_bd_ram_mem0_reg[159][7]/P0001 ,
		_w12774_,
		_w26055_
	);
	LUT2 #(
		.INIT('h8)
	) name15544 (
		\wishbone_bd_ram_mem0_reg[89][7]/P0001 ,
		_w12964_,
		_w26056_
	);
	LUT2 #(
		.INIT('h8)
	) name15545 (
		\wishbone_bd_ram_mem0_reg[171][7]/P0001 ,
		_w12910_,
		_w26057_
	);
	LUT2 #(
		.INIT('h8)
	) name15546 (
		\wishbone_bd_ram_mem0_reg[65][7]/P0001 ,
		_w13176_,
		_w26058_
	);
	LUT2 #(
		.INIT('h8)
	) name15547 (
		\wishbone_bd_ram_mem0_reg[14][7]/P0001 ,
		_w13086_,
		_w26059_
	);
	LUT2 #(
		.INIT('h8)
	) name15548 (
		\wishbone_bd_ram_mem0_reg[25][7]/P0001 ,
		_w13108_,
		_w26060_
	);
	LUT2 #(
		.INIT('h8)
	) name15549 (
		\wishbone_bd_ram_mem0_reg[160][7]/P0001 ,
		_w12872_,
		_w26061_
	);
	LUT2 #(
		.INIT('h8)
	) name15550 (
		\wishbone_bd_ram_mem0_reg[2][7]/P0001 ,
		_w13088_,
		_w26062_
	);
	LUT2 #(
		.INIT('h8)
	) name15551 (
		\wishbone_bd_ram_mem0_reg[254][7]/P0001 ,
		_w12892_,
		_w26063_
	);
	LUT2 #(
		.INIT('h8)
	) name15552 (
		\wishbone_bd_ram_mem0_reg[155][7]/P0001 ,
		_w13122_,
		_w26064_
	);
	LUT2 #(
		.INIT('h8)
	) name15553 (
		\wishbone_bd_ram_mem0_reg[29][7]/P0001 ,
		_w12952_,
		_w26065_
	);
	LUT2 #(
		.INIT('h8)
	) name15554 (
		\wishbone_bd_ram_mem0_reg[0][7]/P0001 ,
		_w12717_,
		_w26066_
	);
	LUT2 #(
		.INIT('h8)
	) name15555 (
		\wishbone_bd_ram_mem0_reg[99][7]/P0001 ,
		_w13038_,
		_w26067_
	);
	LUT2 #(
		.INIT('h8)
	) name15556 (
		\wishbone_bd_ram_mem0_reg[239][7]/P0001 ,
		_w12862_,
		_w26068_
	);
	LUT2 #(
		.INIT('h8)
	) name15557 (
		\wishbone_bd_ram_mem0_reg[62][7]/P0001 ,
		_w12673_,
		_w26069_
	);
	LUT2 #(
		.INIT('h8)
	) name15558 (
		\wishbone_bd_ram_mem0_reg[182][7]/P0001 ,
		_w12820_,
		_w26070_
	);
	LUT2 #(
		.INIT('h8)
	) name15559 (
		\wishbone_bd_ram_mem0_reg[94][7]/P0001 ,
		_w13186_,
		_w26071_
	);
	LUT2 #(
		.INIT('h8)
	) name15560 (
		\wishbone_bd_ram_mem0_reg[41][7]/P0001 ,
		_w13052_,
		_w26072_
	);
	LUT2 #(
		.INIT('h8)
	) name15561 (
		\wishbone_bd_ram_mem0_reg[217][7]/P0001 ,
		_w13188_,
		_w26073_
	);
	LUT2 #(
		.INIT('h8)
	) name15562 (
		\wishbone_bd_ram_mem0_reg[1][7]/P0001 ,
		_w13014_,
		_w26074_
	);
	LUT2 #(
		.INIT('h8)
	) name15563 (
		\wishbone_bd_ram_mem0_reg[84][7]/P0001 ,
		_w12934_,
		_w26075_
	);
	LUT2 #(
		.INIT('h8)
	) name15564 (
		\wishbone_bd_ram_mem0_reg[214][7]/P0001 ,
		_w12984_,
		_w26076_
	);
	LUT2 #(
		.INIT('h8)
	) name15565 (
		\wishbone_bd_ram_mem0_reg[231][7]/P0001 ,
		_w12856_,
		_w26077_
	);
	LUT2 #(
		.INIT('h8)
	) name15566 (
		\wishbone_bd_ram_mem0_reg[205][7]/P0001 ,
		_w13068_,
		_w26078_
	);
	LUT2 #(
		.INIT('h8)
	) name15567 (
		\wishbone_bd_ram_mem0_reg[187][7]/P0001 ,
		_w13196_,
		_w26079_
	);
	LUT2 #(
		.INIT('h8)
	) name15568 (
		\wishbone_bd_ram_mem0_reg[113][7]/P0001 ,
		_w13026_,
		_w26080_
	);
	LUT2 #(
		.INIT('h8)
	) name15569 (
		\wishbone_bd_ram_mem0_reg[126][7]/P0001 ,
		_w13218_,
		_w26081_
	);
	LUT2 #(
		.INIT('h8)
	) name15570 (
		\wishbone_bd_ram_mem0_reg[174][7]/P0001 ,
		_w12972_,
		_w26082_
	);
	LUT2 #(
		.INIT('h8)
	) name15571 (
		\wishbone_bd_ram_mem0_reg[63][7]/P0001 ,
		_w12850_,
		_w26083_
	);
	LUT2 #(
		.INIT('h8)
	) name15572 (
		\wishbone_bd_ram_mem0_reg[115][7]/P0001 ,
		_w13112_,
		_w26084_
	);
	LUT2 #(
		.INIT('h8)
	) name15573 (
		\wishbone_bd_ram_mem0_reg[147][7]/P0001 ,
		_w13146_,
		_w26085_
	);
	LUT2 #(
		.INIT('h8)
	) name15574 (
		\wishbone_bd_ram_mem0_reg[75][7]/P0001 ,
		_w12826_,
		_w26086_
	);
	LUT2 #(
		.INIT('h8)
	) name15575 (
		\wishbone_bd_ram_mem0_reg[18][7]/P0001 ,
		_w12679_,
		_w26087_
	);
	LUT2 #(
		.INIT('h8)
	) name15576 (
		\wishbone_bd_ram_mem0_reg[40][7]/P0001 ,
		_w13132_,
		_w26088_
	);
	LUT2 #(
		.INIT('h8)
	) name15577 (
		\wishbone_bd_ram_mem0_reg[139][7]/P0001 ,
		_w12814_,
		_w26089_
	);
	LUT2 #(
		.INIT('h8)
	) name15578 (
		\wishbone_bd_ram_mem0_reg[157][7]/P0001 ,
		_w12926_,
		_w26090_
	);
	LUT2 #(
		.INIT('h8)
	) name15579 (
		\wishbone_bd_ram_mem0_reg[15][7]/P0001 ,
		_w13210_,
		_w26091_
	);
	LUT2 #(
		.INIT('h8)
	) name15580 (
		\wishbone_bd_ram_mem0_reg[132][7]/P0001 ,
		_w12992_,
		_w26092_
	);
	LUT2 #(
		.INIT('h8)
	) name15581 (
		\wishbone_bd_ram_mem0_reg[87][7]/P0001 ,
		_w13154_,
		_w26093_
	);
	LUT2 #(
		.INIT('h8)
	) name15582 (
		\wishbone_bd_ram_mem0_reg[103][7]/P0001 ,
		_w12846_,
		_w26094_
	);
	LUT2 #(
		.INIT('h8)
	) name15583 (
		\wishbone_bd_ram_mem0_reg[234][7]/P0001 ,
		_w13214_,
		_w26095_
	);
	LUT2 #(
		.INIT('h8)
	) name15584 (
		\wishbone_bd_ram_mem0_reg[81][7]/P0001 ,
		_w12950_,
		_w26096_
	);
	LUT2 #(
		.INIT('h8)
	) name15585 (
		\wishbone_bd_ram_mem0_reg[250][7]/P0001 ,
		_w13128_,
		_w26097_
	);
	LUT2 #(
		.INIT('h8)
	) name15586 (
		\wishbone_bd_ram_mem0_reg[51][7]/P0001 ,
		_w13024_,
		_w26098_
	);
	LUT2 #(
		.INIT('h8)
	) name15587 (
		\wishbone_bd_ram_mem0_reg[209][7]/P0001 ,
		_w13152_,
		_w26099_
	);
	LUT2 #(
		.INIT('h8)
	) name15588 (
		\wishbone_bd_ram_mem0_reg[127][7]/P0001 ,
		_w13164_,
		_w26100_
	);
	LUT2 #(
		.INIT('h8)
	) name15589 (
		\wishbone_bd_ram_mem0_reg[140][7]/P0001 ,
		_w12894_,
		_w26101_
	);
	LUT2 #(
		.INIT('h8)
	) name15590 (
		\wishbone_bd_ram_mem0_reg[137][7]/P0001 ,
		_w13168_,
		_w26102_
	);
	LUT2 #(
		.INIT('h8)
	) name15591 (
		\wishbone_bd_ram_mem0_reg[123][7]/P0001 ,
		_w13114_,
		_w26103_
	);
	LUT2 #(
		.INIT('h8)
	) name15592 (
		\wishbone_bd_ram_mem0_reg[76][7]/P0001 ,
		_w13184_,
		_w26104_
	);
	LUT2 #(
		.INIT('h8)
	) name15593 (
		\wishbone_bd_ram_mem0_reg[88][7]/P0001 ,
		_w12860_,
		_w26105_
	);
	LUT2 #(
		.INIT('h8)
	) name15594 (
		\wishbone_bd_ram_mem0_reg[133][7]/P0001 ,
		_w12761_,
		_w26106_
	);
	LUT2 #(
		.INIT('h8)
	) name15595 (
		\wishbone_bd_ram_mem0_reg[20][7]/P0001 ,
		_w13174_,
		_w26107_
	);
	LUT2 #(
		.INIT('h8)
	) name15596 (
		\wishbone_bd_ram_mem0_reg[204][7]/P0001 ,
		_w13162_,
		_w26108_
	);
	LUT2 #(
		.INIT('h1)
	) name15597 (
		_w25853_,
		_w25854_,
		_w26109_
	);
	LUT2 #(
		.INIT('h1)
	) name15598 (
		_w25855_,
		_w25856_,
		_w26110_
	);
	LUT2 #(
		.INIT('h1)
	) name15599 (
		_w25857_,
		_w25858_,
		_w26111_
	);
	LUT2 #(
		.INIT('h1)
	) name15600 (
		_w25859_,
		_w25860_,
		_w26112_
	);
	LUT2 #(
		.INIT('h1)
	) name15601 (
		_w25861_,
		_w25862_,
		_w26113_
	);
	LUT2 #(
		.INIT('h1)
	) name15602 (
		_w25863_,
		_w25864_,
		_w26114_
	);
	LUT2 #(
		.INIT('h1)
	) name15603 (
		_w25865_,
		_w25866_,
		_w26115_
	);
	LUT2 #(
		.INIT('h1)
	) name15604 (
		_w25867_,
		_w25868_,
		_w26116_
	);
	LUT2 #(
		.INIT('h1)
	) name15605 (
		_w25869_,
		_w25870_,
		_w26117_
	);
	LUT2 #(
		.INIT('h1)
	) name15606 (
		_w25871_,
		_w25872_,
		_w26118_
	);
	LUT2 #(
		.INIT('h1)
	) name15607 (
		_w25873_,
		_w25874_,
		_w26119_
	);
	LUT2 #(
		.INIT('h1)
	) name15608 (
		_w25875_,
		_w25876_,
		_w26120_
	);
	LUT2 #(
		.INIT('h1)
	) name15609 (
		_w25877_,
		_w25878_,
		_w26121_
	);
	LUT2 #(
		.INIT('h1)
	) name15610 (
		_w25879_,
		_w25880_,
		_w26122_
	);
	LUT2 #(
		.INIT('h1)
	) name15611 (
		_w25881_,
		_w25882_,
		_w26123_
	);
	LUT2 #(
		.INIT('h1)
	) name15612 (
		_w25883_,
		_w25884_,
		_w26124_
	);
	LUT2 #(
		.INIT('h1)
	) name15613 (
		_w25885_,
		_w25886_,
		_w26125_
	);
	LUT2 #(
		.INIT('h1)
	) name15614 (
		_w25887_,
		_w25888_,
		_w26126_
	);
	LUT2 #(
		.INIT('h1)
	) name15615 (
		_w25889_,
		_w25890_,
		_w26127_
	);
	LUT2 #(
		.INIT('h1)
	) name15616 (
		_w25891_,
		_w25892_,
		_w26128_
	);
	LUT2 #(
		.INIT('h1)
	) name15617 (
		_w25893_,
		_w25894_,
		_w26129_
	);
	LUT2 #(
		.INIT('h1)
	) name15618 (
		_w25895_,
		_w25896_,
		_w26130_
	);
	LUT2 #(
		.INIT('h1)
	) name15619 (
		_w25897_,
		_w25898_,
		_w26131_
	);
	LUT2 #(
		.INIT('h1)
	) name15620 (
		_w25899_,
		_w25900_,
		_w26132_
	);
	LUT2 #(
		.INIT('h1)
	) name15621 (
		_w25901_,
		_w25902_,
		_w26133_
	);
	LUT2 #(
		.INIT('h1)
	) name15622 (
		_w25903_,
		_w25904_,
		_w26134_
	);
	LUT2 #(
		.INIT('h1)
	) name15623 (
		_w25905_,
		_w25906_,
		_w26135_
	);
	LUT2 #(
		.INIT('h1)
	) name15624 (
		_w25907_,
		_w25908_,
		_w26136_
	);
	LUT2 #(
		.INIT('h1)
	) name15625 (
		_w25909_,
		_w25910_,
		_w26137_
	);
	LUT2 #(
		.INIT('h1)
	) name15626 (
		_w25911_,
		_w25912_,
		_w26138_
	);
	LUT2 #(
		.INIT('h1)
	) name15627 (
		_w25913_,
		_w25914_,
		_w26139_
	);
	LUT2 #(
		.INIT('h1)
	) name15628 (
		_w25915_,
		_w25916_,
		_w26140_
	);
	LUT2 #(
		.INIT('h1)
	) name15629 (
		_w25917_,
		_w25918_,
		_w26141_
	);
	LUT2 #(
		.INIT('h1)
	) name15630 (
		_w25919_,
		_w25920_,
		_w26142_
	);
	LUT2 #(
		.INIT('h1)
	) name15631 (
		_w25921_,
		_w25922_,
		_w26143_
	);
	LUT2 #(
		.INIT('h1)
	) name15632 (
		_w25923_,
		_w25924_,
		_w26144_
	);
	LUT2 #(
		.INIT('h1)
	) name15633 (
		_w25925_,
		_w25926_,
		_w26145_
	);
	LUT2 #(
		.INIT('h1)
	) name15634 (
		_w25927_,
		_w25928_,
		_w26146_
	);
	LUT2 #(
		.INIT('h1)
	) name15635 (
		_w25929_,
		_w25930_,
		_w26147_
	);
	LUT2 #(
		.INIT('h1)
	) name15636 (
		_w25931_,
		_w25932_,
		_w26148_
	);
	LUT2 #(
		.INIT('h1)
	) name15637 (
		_w25933_,
		_w25934_,
		_w26149_
	);
	LUT2 #(
		.INIT('h1)
	) name15638 (
		_w25935_,
		_w25936_,
		_w26150_
	);
	LUT2 #(
		.INIT('h1)
	) name15639 (
		_w25937_,
		_w25938_,
		_w26151_
	);
	LUT2 #(
		.INIT('h1)
	) name15640 (
		_w25939_,
		_w25940_,
		_w26152_
	);
	LUT2 #(
		.INIT('h1)
	) name15641 (
		_w25941_,
		_w25942_,
		_w26153_
	);
	LUT2 #(
		.INIT('h1)
	) name15642 (
		_w25943_,
		_w25944_,
		_w26154_
	);
	LUT2 #(
		.INIT('h1)
	) name15643 (
		_w25945_,
		_w25946_,
		_w26155_
	);
	LUT2 #(
		.INIT('h1)
	) name15644 (
		_w25947_,
		_w25948_,
		_w26156_
	);
	LUT2 #(
		.INIT('h1)
	) name15645 (
		_w25949_,
		_w25950_,
		_w26157_
	);
	LUT2 #(
		.INIT('h1)
	) name15646 (
		_w25951_,
		_w25952_,
		_w26158_
	);
	LUT2 #(
		.INIT('h1)
	) name15647 (
		_w25953_,
		_w25954_,
		_w26159_
	);
	LUT2 #(
		.INIT('h1)
	) name15648 (
		_w25955_,
		_w25956_,
		_w26160_
	);
	LUT2 #(
		.INIT('h1)
	) name15649 (
		_w25957_,
		_w25958_,
		_w26161_
	);
	LUT2 #(
		.INIT('h1)
	) name15650 (
		_w25959_,
		_w25960_,
		_w26162_
	);
	LUT2 #(
		.INIT('h1)
	) name15651 (
		_w25961_,
		_w25962_,
		_w26163_
	);
	LUT2 #(
		.INIT('h1)
	) name15652 (
		_w25963_,
		_w25964_,
		_w26164_
	);
	LUT2 #(
		.INIT('h1)
	) name15653 (
		_w25965_,
		_w25966_,
		_w26165_
	);
	LUT2 #(
		.INIT('h1)
	) name15654 (
		_w25967_,
		_w25968_,
		_w26166_
	);
	LUT2 #(
		.INIT('h1)
	) name15655 (
		_w25969_,
		_w25970_,
		_w26167_
	);
	LUT2 #(
		.INIT('h1)
	) name15656 (
		_w25971_,
		_w25972_,
		_w26168_
	);
	LUT2 #(
		.INIT('h1)
	) name15657 (
		_w25973_,
		_w25974_,
		_w26169_
	);
	LUT2 #(
		.INIT('h1)
	) name15658 (
		_w25975_,
		_w25976_,
		_w26170_
	);
	LUT2 #(
		.INIT('h1)
	) name15659 (
		_w25977_,
		_w25978_,
		_w26171_
	);
	LUT2 #(
		.INIT('h1)
	) name15660 (
		_w25979_,
		_w25980_,
		_w26172_
	);
	LUT2 #(
		.INIT('h1)
	) name15661 (
		_w25981_,
		_w25982_,
		_w26173_
	);
	LUT2 #(
		.INIT('h1)
	) name15662 (
		_w25983_,
		_w25984_,
		_w26174_
	);
	LUT2 #(
		.INIT('h1)
	) name15663 (
		_w25985_,
		_w25986_,
		_w26175_
	);
	LUT2 #(
		.INIT('h1)
	) name15664 (
		_w25987_,
		_w25988_,
		_w26176_
	);
	LUT2 #(
		.INIT('h1)
	) name15665 (
		_w25989_,
		_w25990_,
		_w26177_
	);
	LUT2 #(
		.INIT('h1)
	) name15666 (
		_w25991_,
		_w25992_,
		_w26178_
	);
	LUT2 #(
		.INIT('h1)
	) name15667 (
		_w25993_,
		_w25994_,
		_w26179_
	);
	LUT2 #(
		.INIT('h1)
	) name15668 (
		_w25995_,
		_w25996_,
		_w26180_
	);
	LUT2 #(
		.INIT('h1)
	) name15669 (
		_w25997_,
		_w25998_,
		_w26181_
	);
	LUT2 #(
		.INIT('h1)
	) name15670 (
		_w25999_,
		_w26000_,
		_w26182_
	);
	LUT2 #(
		.INIT('h1)
	) name15671 (
		_w26001_,
		_w26002_,
		_w26183_
	);
	LUT2 #(
		.INIT('h1)
	) name15672 (
		_w26003_,
		_w26004_,
		_w26184_
	);
	LUT2 #(
		.INIT('h1)
	) name15673 (
		_w26005_,
		_w26006_,
		_w26185_
	);
	LUT2 #(
		.INIT('h1)
	) name15674 (
		_w26007_,
		_w26008_,
		_w26186_
	);
	LUT2 #(
		.INIT('h1)
	) name15675 (
		_w26009_,
		_w26010_,
		_w26187_
	);
	LUT2 #(
		.INIT('h1)
	) name15676 (
		_w26011_,
		_w26012_,
		_w26188_
	);
	LUT2 #(
		.INIT('h1)
	) name15677 (
		_w26013_,
		_w26014_,
		_w26189_
	);
	LUT2 #(
		.INIT('h1)
	) name15678 (
		_w26015_,
		_w26016_,
		_w26190_
	);
	LUT2 #(
		.INIT('h1)
	) name15679 (
		_w26017_,
		_w26018_,
		_w26191_
	);
	LUT2 #(
		.INIT('h1)
	) name15680 (
		_w26019_,
		_w26020_,
		_w26192_
	);
	LUT2 #(
		.INIT('h1)
	) name15681 (
		_w26021_,
		_w26022_,
		_w26193_
	);
	LUT2 #(
		.INIT('h1)
	) name15682 (
		_w26023_,
		_w26024_,
		_w26194_
	);
	LUT2 #(
		.INIT('h1)
	) name15683 (
		_w26025_,
		_w26026_,
		_w26195_
	);
	LUT2 #(
		.INIT('h1)
	) name15684 (
		_w26027_,
		_w26028_,
		_w26196_
	);
	LUT2 #(
		.INIT('h1)
	) name15685 (
		_w26029_,
		_w26030_,
		_w26197_
	);
	LUT2 #(
		.INIT('h1)
	) name15686 (
		_w26031_,
		_w26032_,
		_w26198_
	);
	LUT2 #(
		.INIT('h1)
	) name15687 (
		_w26033_,
		_w26034_,
		_w26199_
	);
	LUT2 #(
		.INIT('h1)
	) name15688 (
		_w26035_,
		_w26036_,
		_w26200_
	);
	LUT2 #(
		.INIT('h1)
	) name15689 (
		_w26037_,
		_w26038_,
		_w26201_
	);
	LUT2 #(
		.INIT('h1)
	) name15690 (
		_w26039_,
		_w26040_,
		_w26202_
	);
	LUT2 #(
		.INIT('h1)
	) name15691 (
		_w26041_,
		_w26042_,
		_w26203_
	);
	LUT2 #(
		.INIT('h1)
	) name15692 (
		_w26043_,
		_w26044_,
		_w26204_
	);
	LUT2 #(
		.INIT('h1)
	) name15693 (
		_w26045_,
		_w26046_,
		_w26205_
	);
	LUT2 #(
		.INIT('h1)
	) name15694 (
		_w26047_,
		_w26048_,
		_w26206_
	);
	LUT2 #(
		.INIT('h1)
	) name15695 (
		_w26049_,
		_w26050_,
		_w26207_
	);
	LUT2 #(
		.INIT('h1)
	) name15696 (
		_w26051_,
		_w26052_,
		_w26208_
	);
	LUT2 #(
		.INIT('h1)
	) name15697 (
		_w26053_,
		_w26054_,
		_w26209_
	);
	LUT2 #(
		.INIT('h1)
	) name15698 (
		_w26055_,
		_w26056_,
		_w26210_
	);
	LUT2 #(
		.INIT('h1)
	) name15699 (
		_w26057_,
		_w26058_,
		_w26211_
	);
	LUT2 #(
		.INIT('h1)
	) name15700 (
		_w26059_,
		_w26060_,
		_w26212_
	);
	LUT2 #(
		.INIT('h1)
	) name15701 (
		_w26061_,
		_w26062_,
		_w26213_
	);
	LUT2 #(
		.INIT('h1)
	) name15702 (
		_w26063_,
		_w26064_,
		_w26214_
	);
	LUT2 #(
		.INIT('h1)
	) name15703 (
		_w26065_,
		_w26066_,
		_w26215_
	);
	LUT2 #(
		.INIT('h1)
	) name15704 (
		_w26067_,
		_w26068_,
		_w26216_
	);
	LUT2 #(
		.INIT('h1)
	) name15705 (
		_w26069_,
		_w26070_,
		_w26217_
	);
	LUT2 #(
		.INIT('h1)
	) name15706 (
		_w26071_,
		_w26072_,
		_w26218_
	);
	LUT2 #(
		.INIT('h1)
	) name15707 (
		_w26073_,
		_w26074_,
		_w26219_
	);
	LUT2 #(
		.INIT('h1)
	) name15708 (
		_w26075_,
		_w26076_,
		_w26220_
	);
	LUT2 #(
		.INIT('h1)
	) name15709 (
		_w26077_,
		_w26078_,
		_w26221_
	);
	LUT2 #(
		.INIT('h1)
	) name15710 (
		_w26079_,
		_w26080_,
		_w26222_
	);
	LUT2 #(
		.INIT('h1)
	) name15711 (
		_w26081_,
		_w26082_,
		_w26223_
	);
	LUT2 #(
		.INIT('h1)
	) name15712 (
		_w26083_,
		_w26084_,
		_w26224_
	);
	LUT2 #(
		.INIT('h1)
	) name15713 (
		_w26085_,
		_w26086_,
		_w26225_
	);
	LUT2 #(
		.INIT('h1)
	) name15714 (
		_w26087_,
		_w26088_,
		_w26226_
	);
	LUT2 #(
		.INIT('h1)
	) name15715 (
		_w26089_,
		_w26090_,
		_w26227_
	);
	LUT2 #(
		.INIT('h1)
	) name15716 (
		_w26091_,
		_w26092_,
		_w26228_
	);
	LUT2 #(
		.INIT('h1)
	) name15717 (
		_w26093_,
		_w26094_,
		_w26229_
	);
	LUT2 #(
		.INIT('h1)
	) name15718 (
		_w26095_,
		_w26096_,
		_w26230_
	);
	LUT2 #(
		.INIT('h1)
	) name15719 (
		_w26097_,
		_w26098_,
		_w26231_
	);
	LUT2 #(
		.INIT('h1)
	) name15720 (
		_w26099_,
		_w26100_,
		_w26232_
	);
	LUT2 #(
		.INIT('h1)
	) name15721 (
		_w26101_,
		_w26102_,
		_w26233_
	);
	LUT2 #(
		.INIT('h1)
	) name15722 (
		_w26103_,
		_w26104_,
		_w26234_
	);
	LUT2 #(
		.INIT('h1)
	) name15723 (
		_w26105_,
		_w26106_,
		_w26235_
	);
	LUT2 #(
		.INIT('h1)
	) name15724 (
		_w26107_,
		_w26108_,
		_w26236_
	);
	LUT2 #(
		.INIT('h8)
	) name15725 (
		_w26235_,
		_w26236_,
		_w26237_
	);
	LUT2 #(
		.INIT('h8)
	) name15726 (
		_w26233_,
		_w26234_,
		_w26238_
	);
	LUT2 #(
		.INIT('h8)
	) name15727 (
		_w26231_,
		_w26232_,
		_w26239_
	);
	LUT2 #(
		.INIT('h8)
	) name15728 (
		_w26229_,
		_w26230_,
		_w26240_
	);
	LUT2 #(
		.INIT('h8)
	) name15729 (
		_w26227_,
		_w26228_,
		_w26241_
	);
	LUT2 #(
		.INIT('h8)
	) name15730 (
		_w26225_,
		_w26226_,
		_w26242_
	);
	LUT2 #(
		.INIT('h8)
	) name15731 (
		_w26223_,
		_w26224_,
		_w26243_
	);
	LUT2 #(
		.INIT('h8)
	) name15732 (
		_w26221_,
		_w26222_,
		_w26244_
	);
	LUT2 #(
		.INIT('h8)
	) name15733 (
		_w26219_,
		_w26220_,
		_w26245_
	);
	LUT2 #(
		.INIT('h8)
	) name15734 (
		_w26217_,
		_w26218_,
		_w26246_
	);
	LUT2 #(
		.INIT('h8)
	) name15735 (
		_w26215_,
		_w26216_,
		_w26247_
	);
	LUT2 #(
		.INIT('h8)
	) name15736 (
		_w26213_,
		_w26214_,
		_w26248_
	);
	LUT2 #(
		.INIT('h8)
	) name15737 (
		_w26211_,
		_w26212_,
		_w26249_
	);
	LUT2 #(
		.INIT('h8)
	) name15738 (
		_w26209_,
		_w26210_,
		_w26250_
	);
	LUT2 #(
		.INIT('h8)
	) name15739 (
		_w26207_,
		_w26208_,
		_w26251_
	);
	LUT2 #(
		.INIT('h8)
	) name15740 (
		_w26205_,
		_w26206_,
		_w26252_
	);
	LUT2 #(
		.INIT('h8)
	) name15741 (
		_w26203_,
		_w26204_,
		_w26253_
	);
	LUT2 #(
		.INIT('h8)
	) name15742 (
		_w26201_,
		_w26202_,
		_w26254_
	);
	LUT2 #(
		.INIT('h8)
	) name15743 (
		_w26199_,
		_w26200_,
		_w26255_
	);
	LUT2 #(
		.INIT('h8)
	) name15744 (
		_w26197_,
		_w26198_,
		_w26256_
	);
	LUT2 #(
		.INIT('h8)
	) name15745 (
		_w26195_,
		_w26196_,
		_w26257_
	);
	LUT2 #(
		.INIT('h8)
	) name15746 (
		_w26193_,
		_w26194_,
		_w26258_
	);
	LUT2 #(
		.INIT('h8)
	) name15747 (
		_w26191_,
		_w26192_,
		_w26259_
	);
	LUT2 #(
		.INIT('h8)
	) name15748 (
		_w26189_,
		_w26190_,
		_w26260_
	);
	LUT2 #(
		.INIT('h8)
	) name15749 (
		_w26187_,
		_w26188_,
		_w26261_
	);
	LUT2 #(
		.INIT('h8)
	) name15750 (
		_w26185_,
		_w26186_,
		_w26262_
	);
	LUT2 #(
		.INIT('h8)
	) name15751 (
		_w26183_,
		_w26184_,
		_w26263_
	);
	LUT2 #(
		.INIT('h8)
	) name15752 (
		_w26181_,
		_w26182_,
		_w26264_
	);
	LUT2 #(
		.INIT('h8)
	) name15753 (
		_w26179_,
		_w26180_,
		_w26265_
	);
	LUT2 #(
		.INIT('h8)
	) name15754 (
		_w26177_,
		_w26178_,
		_w26266_
	);
	LUT2 #(
		.INIT('h8)
	) name15755 (
		_w26175_,
		_w26176_,
		_w26267_
	);
	LUT2 #(
		.INIT('h8)
	) name15756 (
		_w26173_,
		_w26174_,
		_w26268_
	);
	LUT2 #(
		.INIT('h8)
	) name15757 (
		_w26171_,
		_w26172_,
		_w26269_
	);
	LUT2 #(
		.INIT('h8)
	) name15758 (
		_w26169_,
		_w26170_,
		_w26270_
	);
	LUT2 #(
		.INIT('h8)
	) name15759 (
		_w26167_,
		_w26168_,
		_w26271_
	);
	LUT2 #(
		.INIT('h8)
	) name15760 (
		_w26165_,
		_w26166_,
		_w26272_
	);
	LUT2 #(
		.INIT('h8)
	) name15761 (
		_w26163_,
		_w26164_,
		_w26273_
	);
	LUT2 #(
		.INIT('h8)
	) name15762 (
		_w26161_,
		_w26162_,
		_w26274_
	);
	LUT2 #(
		.INIT('h8)
	) name15763 (
		_w26159_,
		_w26160_,
		_w26275_
	);
	LUT2 #(
		.INIT('h8)
	) name15764 (
		_w26157_,
		_w26158_,
		_w26276_
	);
	LUT2 #(
		.INIT('h8)
	) name15765 (
		_w26155_,
		_w26156_,
		_w26277_
	);
	LUT2 #(
		.INIT('h8)
	) name15766 (
		_w26153_,
		_w26154_,
		_w26278_
	);
	LUT2 #(
		.INIT('h8)
	) name15767 (
		_w26151_,
		_w26152_,
		_w26279_
	);
	LUT2 #(
		.INIT('h8)
	) name15768 (
		_w26149_,
		_w26150_,
		_w26280_
	);
	LUT2 #(
		.INIT('h8)
	) name15769 (
		_w26147_,
		_w26148_,
		_w26281_
	);
	LUT2 #(
		.INIT('h8)
	) name15770 (
		_w26145_,
		_w26146_,
		_w26282_
	);
	LUT2 #(
		.INIT('h8)
	) name15771 (
		_w26143_,
		_w26144_,
		_w26283_
	);
	LUT2 #(
		.INIT('h8)
	) name15772 (
		_w26141_,
		_w26142_,
		_w26284_
	);
	LUT2 #(
		.INIT('h8)
	) name15773 (
		_w26139_,
		_w26140_,
		_w26285_
	);
	LUT2 #(
		.INIT('h8)
	) name15774 (
		_w26137_,
		_w26138_,
		_w26286_
	);
	LUT2 #(
		.INIT('h8)
	) name15775 (
		_w26135_,
		_w26136_,
		_w26287_
	);
	LUT2 #(
		.INIT('h8)
	) name15776 (
		_w26133_,
		_w26134_,
		_w26288_
	);
	LUT2 #(
		.INIT('h8)
	) name15777 (
		_w26131_,
		_w26132_,
		_w26289_
	);
	LUT2 #(
		.INIT('h8)
	) name15778 (
		_w26129_,
		_w26130_,
		_w26290_
	);
	LUT2 #(
		.INIT('h8)
	) name15779 (
		_w26127_,
		_w26128_,
		_w26291_
	);
	LUT2 #(
		.INIT('h8)
	) name15780 (
		_w26125_,
		_w26126_,
		_w26292_
	);
	LUT2 #(
		.INIT('h8)
	) name15781 (
		_w26123_,
		_w26124_,
		_w26293_
	);
	LUT2 #(
		.INIT('h8)
	) name15782 (
		_w26121_,
		_w26122_,
		_w26294_
	);
	LUT2 #(
		.INIT('h8)
	) name15783 (
		_w26119_,
		_w26120_,
		_w26295_
	);
	LUT2 #(
		.INIT('h8)
	) name15784 (
		_w26117_,
		_w26118_,
		_w26296_
	);
	LUT2 #(
		.INIT('h8)
	) name15785 (
		_w26115_,
		_w26116_,
		_w26297_
	);
	LUT2 #(
		.INIT('h8)
	) name15786 (
		_w26113_,
		_w26114_,
		_w26298_
	);
	LUT2 #(
		.INIT('h8)
	) name15787 (
		_w26111_,
		_w26112_,
		_w26299_
	);
	LUT2 #(
		.INIT('h8)
	) name15788 (
		_w26109_,
		_w26110_,
		_w26300_
	);
	LUT2 #(
		.INIT('h8)
	) name15789 (
		_w26299_,
		_w26300_,
		_w26301_
	);
	LUT2 #(
		.INIT('h8)
	) name15790 (
		_w26297_,
		_w26298_,
		_w26302_
	);
	LUT2 #(
		.INIT('h8)
	) name15791 (
		_w26295_,
		_w26296_,
		_w26303_
	);
	LUT2 #(
		.INIT('h8)
	) name15792 (
		_w26293_,
		_w26294_,
		_w26304_
	);
	LUT2 #(
		.INIT('h8)
	) name15793 (
		_w26291_,
		_w26292_,
		_w26305_
	);
	LUT2 #(
		.INIT('h8)
	) name15794 (
		_w26289_,
		_w26290_,
		_w26306_
	);
	LUT2 #(
		.INIT('h8)
	) name15795 (
		_w26287_,
		_w26288_,
		_w26307_
	);
	LUT2 #(
		.INIT('h8)
	) name15796 (
		_w26285_,
		_w26286_,
		_w26308_
	);
	LUT2 #(
		.INIT('h8)
	) name15797 (
		_w26283_,
		_w26284_,
		_w26309_
	);
	LUT2 #(
		.INIT('h8)
	) name15798 (
		_w26281_,
		_w26282_,
		_w26310_
	);
	LUT2 #(
		.INIT('h8)
	) name15799 (
		_w26279_,
		_w26280_,
		_w26311_
	);
	LUT2 #(
		.INIT('h8)
	) name15800 (
		_w26277_,
		_w26278_,
		_w26312_
	);
	LUT2 #(
		.INIT('h8)
	) name15801 (
		_w26275_,
		_w26276_,
		_w26313_
	);
	LUT2 #(
		.INIT('h8)
	) name15802 (
		_w26273_,
		_w26274_,
		_w26314_
	);
	LUT2 #(
		.INIT('h8)
	) name15803 (
		_w26271_,
		_w26272_,
		_w26315_
	);
	LUT2 #(
		.INIT('h8)
	) name15804 (
		_w26269_,
		_w26270_,
		_w26316_
	);
	LUT2 #(
		.INIT('h8)
	) name15805 (
		_w26267_,
		_w26268_,
		_w26317_
	);
	LUT2 #(
		.INIT('h8)
	) name15806 (
		_w26265_,
		_w26266_,
		_w26318_
	);
	LUT2 #(
		.INIT('h8)
	) name15807 (
		_w26263_,
		_w26264_,
		_w26319_
	);
	LUT2 #(
		.INIT('h8)
	) name15808 (
		_w26261_,
		_w26262_,
		_w26320_
	);
	LUT2 #(
		.INIT('h8)
	) name15809 (
		_w26259_,
		_w26260_,
		_w26321_
	);
	LUT2 #(
		.INIT('h8)
	) name15810 (
		_w26257_,
		_w26258_,
		_w26322_
	);
	LUT2 #(
		.INIT('h8)
	) name15811 (
		_w26255_,
		_w26256_,
		_w26323_
	);
	LUT2 #(
		.INIT('h8)
	) name15812 (
		_w26253_,
		_w26254_,
		_w26324_
	);
	LUT2 #(
		.INIT('h8)
	) name15813 (
		_w26251_,
		_w26252_,
		_w26325_
	);
	LUT2 #(
		.INIT('h8)
	) name15814 (
		_w26249_,
		_w26250_,
		_w26326_
	);
	LUT2 #(
		.INIT('h8)
	) name15815 (
		_w26247_,
		_w26248_,
		_w26327_
	);
	LUT2 #(
		.INIT('h8)
	) name15816 (
		_w26245_,
		_w26246_,
		_w26328_
	);
	LUT2 #(
		.INIT('h8)
	) name15817 (
		_w26243_,
		_w26244_,
		_w26329_
	);
	LUT2 #(
		.INIT('h8)
	) name15818 (
		_w26241_,
		_w26242_,
		_w26330_
	);
	LUT2 #(
		.INIT('h8)
	) name15819 (
		_w26239_,
		_w26240_,
		_w26331_
	);
	LUT2 #(
		.INIT('h8)
	) name15820 (
		_w26237_,
		_w26238_,
		_w26332_
	);
	LUT2 #(
		.INIT('h8)
	) name15821 (
		_w26331_,
		_w26332_,
		_w26333_
	);
	LUT2 #(
		.INIT('h8)
	) name15822 (
		_w26329_,
		_w26330_,
		_w26334_
	);
	LUT2 #(
		.INIT('h8)
	) name15823 (
		_w26327_,
		_w26328_,
		_w26335_
	);
	LUT2 #(
		.INIT('h8)
	) name15824 (
		_w26325_,
		_w26326_,
		_w26336_
	);
	LUT2 #(
		.INIT('h8)
	) name15825 (
		_w26323_,
		_w26324_,
		_w26337_
	);
	LUT2 #(
		.INIT('h8)
	) name15826 (
		_w26321_,
		_w26322_,
		_w26338_
	);
	LUT2 #(
		.INIT('h8)
	) name15827 (
		_w26319_,
		_w26320_,
		_w26339_
	);
	LUT2 #(
		.INIT('h8)
	) name15828 (
		_w26317_,
		_w26318_,
		_w26340_
	);
	LUT2 #(
		.INIT('h8)
	) name15829 (
		_w26315_,
		_w26316_,
		_w26341_
	);
	LUT2 #(
		.INIT('h8)
	) name15830 (
		_w26313_,
		_w26314_,
		_w26342_
	);
	LUT2 #(
		.INIT('h8)
	) name15831 (
		_w26311_,
		_w26312_,
		_w26343_
	);
	LUT2 #(
		.INIT('h8)
	) name15832 (
		_w26309_,
		_w26310_,
		_w26344_
	);
	LUT2 #(
		.INIT('h8)
	) name15833 (
		_w26307_,
		_w26308_,
		_w26345_
	);
	LUT2 #(
		.INIT('h8)
	) name15834 (
		_w26305_,
		_w26306_,
		_w26346_
	);
	LUT2 #(
		.INIT('h8)
	) name15835 (
		_w26303_,
		_w26304_,
		_w26347_
	);
	LUT2 #(
		.INIT('h8)
	) name15836 (
		_w26301_,
		_w26302_,
		_w26348_
	);
	LUT2 #(
		.INIT('h8)
	) name15837 (
		_w26347_,
		_w26348_,
		_w26349_
	);
	LUT2 #(
		.INIT('h8)
	) name15838 (
		_w26345_,
		_w26346_,
		_w26350_
	);
	LUT2 #(
		.INIT('h8)
	) name15839 (
		_w26343_,
		_w26344_,
		_w26351_
	);
	LUT2 #(
		.INIT('h8)
	) name15840 (
		_w26341_,
		_w26342_,
		_w26352_
	);
	LUT2 #(
		.INIT('h8)
	) name15841 (
		_w26339_,
		_w26340_,
		_w26353_
	);
	LUT2 #(
		.INIT('h8)
	) name15842 (
		_w26337_,
		_w26338_,
		_w26354_
	);
	LUT2 #(
		.INIT('h8)
	) name15843 (
		_w26335_,
		_w26336_,
		_w26355_
	);
	LUT2 #(
		.INIT('h8)
	) name15844 (
		_w26333_,
		_w26334_,
		_w26356_
	);
	LUT2 #(
		.INIT('h8)
	) name15845 (
		_w26355_,
		_w26356_,
		_w26357_
	);
	LUT2 #(
		.INIT('h8)
	) name15846 (
		_w26353_,
		_w26354_,
		_w26358_
	);
	LUT2 #(
		.INIT('h8)
	) name15847 (
		_w26351_,
		_w26352_,
		_w26359_
	);
	LUT2 #(
		.INIT('h8)
	) name15848 (
		_w26349_,
		_w26350_,
		_w26360_
	);
	LUT2 #(
		.INIT('h8)
	) name15849 (
		_w26359_,
		_w26360_,
		_w26361_
	);
	LUT2 #(
		.INIT('h8)
	) name15850 (
		_w26357_,
		_w26358_,
		_w26362_
	);
	LUT2 #(
		.INIT('h8)
	) name15851 (
		_w26361_,
		_w26362_,
		_w26363_
	);
	LUT2 #(
		.INIT('h1)
	) name15852 (
		wb_rst_i_pad,
		_w26363_,
		_w26364_
	);
	LUT2 #(
		.INIT('h1)
	) name15853 (
		_w22944_,
		_w26364_,
		_w26365_
	);
	LUT2 #(
		.INIT('h8)
	) name15854 (
		\ethreg1_PACKETLEN_0_DataOut_reg[7]/NET0131 ,
		_w22966_,
		_w26366_
	);
	LUT2 #(
		.INIT('h8)
	) name15855 (
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w24726_,
		_w26367_
	);
	LUT2 #(
		.INIT('h8)
	) name15856 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		_w23519_,
		_w26368_
	);
	LUT2 #(
		.INIT('h8)
	) name15857 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		_w22959_,
		_w26369_
	);
	LUT2 #(
		.INIT('h8)
	) name15858 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w24713_,
		_w26370_
	);
	LUT2 #(
		.INIT('h8)
	) name15859 (
		\ethreg1_MIIRX_DATA_DataOut_reg[7]/NET0131 ,
		_w23507_,
		_w26371_
	);
	LUT2 #(
		.INIT('h8)
	) name15860 (
		\ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 ,
		_w22952_,
		_w26372_
	);
	LUT2 #(
		.INIT('h8)
	) name15861 (
		\ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 ,
		_w22956_,
		_w26373_
	);
	LUT2 #(
		.INIT('h8)
	) name15862 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		_w23501_,
		_w26374_
	);
	LUT2 #(
		.INIT('h8)
	) name15863 (
		\ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 ,
		_w23499_,
		_w26375_
	);
	LUT2 #(
		.INIT('h8)
	) name15864 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 ,
		_w23522_,
		_w26376_
	);
	LUT2 #(
		.INIT('h1)
	) name15865 (
		_w26367_,
		_w26368_,
		_w26377_
	);
	LUT2 #(
		.INIT('h1)
	) name15866 (
		_w26369_,
		_w26370_,
		_w26378_
	);
	LUT2 #(
		.INIT('h1)
	) name15867 (
		_w26371_,
		_w26372_,
		_w26379_
	);
	LUT2 #(
		.INIT('h1)
	) name15868 (
		_w26373_,
		_w26374_,
		_w26380_
	);
	LUT2 #(
		.INIT('h1)
	) name15869 (
		_w26375_,
		_w26376_,
		_w26381_
	);
	LUT2 #(
		.INIT('h8)
	) name15870 (
		_w26380_,
		_w26381_,
		_w26382_
	);
	LUT2 #(
		.INIT('h8)
	) name15871 (
		_w26378_,
		_w26379_,
		_w26383_
	);
	LUT2 #(
		.INIT('h8)
	) name15872 (
		_w22944_,
		_w26377_,
		_w26384_
	);
	LUT2 #(
		.INIT('h8)
	) name15873 (
		_w26383_,
		_w26384_,
		_w26385_
	);
	LUT2 #(
		.INIT('h4)
	) name15874 (
		_w26366_,
		_w26382_,
		_w26386_
	);
	LUT2 #(
		.INIT('h8)
	) name15875 (
		_w26385_,
		_w26386_,
		_w26387_
	);
	LUT2 #(
		.INIT('h1)
	) name15876 (
		_w26365_,
		_w26387_,
		_w26388_
	);
	LUT2 #(
		.INIT('h8)
	) name15877 (
		\wishbone_bd_ram_mem1_reg[2][8]/P0001 ,
		_w13088_,
		_w26389_
	);
	LUT2 #(
		.INIT('h8)
	) name15878 (
		\wishbone_bd_ram_mem1_reg[56][8]/P0001 ,
		_w12778_,
		_w26390_
	);
	LUT2 #(
		.INIT('h8)
	) name15879 (
		\wishbone_bd_ram_mem1_reg[27][8]/P0001 ,
		_w12880_,
		_w26391_
	);
	LUT2 #(
		.INIT('h8)
	) name15880 (
		\wishbone_bd_ram_mem1_reg[189][8]/P0001 ,
		_w13042_,
		_w26392_
	);
	LUT2 #(
		.INIT('h8)
	) name15881 (
		\wishbone_bd_ram_mem1_reg[98][8]/P0001 ,
		_w12816_,
		_w26393_
	);
	LUT2 #(
		.INIT('h8)
	) name15882 (
		\wishbone_bd_ram_mem1_reg[84][8]/P0001 ,
		_w12934_,
		_w26394_
	);
	LUT2 #(
		.INIT('h8)
	) name15883 (
		\wishbone_bd_ram_mem1_reg[148][8]/P0001 ,
		_w13000_,
		_w26395_
	);
	LUT2 #(
		.INIT('h8)
	) name15884 (
		\wishbone_bd_ram_mem1_reg[115][8]/P0001 ,
		_w13112_,
		_w26396_
	);
	LUT2 #(
		.INIT('h8)
	) name15885 (
		\wishbone_bd_ram_mem1_reg[3][8]/P0001 ,
		_w12866_,
		_w26397_
	);
	LUT2 #(
		.INIT('h8)
	) name15886 (
		\wishbone_bd_ram_mem1_reg[253][8]/P0001 ,
		_w13100_,
		_w26398_
	);
	LUT2 #(
		.INIT('h8)
	) name15887 (
		\wishbone_bd_ram_mem1_reg[191][8]/P0001 ,
		_w13034_,
		_w26399_
	);
	LUT2 #(
		.INIT('h8)
	) name15888 (
		\wishbone_bd_ram_mem1_reg[152][8]/P0001 ,
		_w12966_,
		_w26400_
	);
	LUT2 #(
		.INIT('h8)
	) name15889 (
		\wishbone_bd_ram_mem1_reg[50][8]/P0001 ,
		_w13150_,
		_w26401_
	);
	LUT2 #(
		.INIT('h8)
	) name15890 (
		\wishbone_bd_ram_mem1_reg[177][8]/P0001 ,
		_w12996_,
		_w26402_
	);
	LUT2 #(
		.INIT('h8)
	) name15891 (
		\wishbone_bd_ram_mem1_reg[135][8]/P0001 ,
		_w13124_,
		_w26403_
	);
	LUT2 #(
		.INIT('h8)
	) name15892 (
		\wishbone_bd_ram_mem1_reg[51][8]/P0001 ,
		_w13024_,
		_w26404_
	);
	LUT2 #(
		.INIT('h8)
	) name15893 (
		\wishbone_bd_ram_mem1_reg[166][8]/P0001 ,
		_w13040_,
		_w26405_
	);
	LUT2 #(
		.INIT('h8)
	) name15894 (
		\wishbone_bd_ram_mem1_reg[133][8]/P0001 ,
		_w12761_,
		_w26406_
	);
	LUT2 #(
		.INIT('h8)
	) name15895 (
		\wishbone_bd_ram_mem1_reg[170][8]/P0001 ,
		_w13030_,
		_w26407_
	);
	LUT2 #(
		.INIT('h8)
	) name15896 (
		\wishbone_bd_ram_mem1_reg[173][8]/P0001 ,
		_w12854_,
		_w26408_
	);
	LUT2 #(
		.INIT('h8)
	) name15897 (
		\wishbone_bd_ram_mem1_reg[78][8]/P0001 ,
		_w12874_,
		_w26409_
	);
	LUT2 #(
		.INIT('h8)
	) name15898 (
		\wishbone_bd_ram_mem1_reg[228][8]/P0001 ,
		_w12765_,
		_w26410_
	);
	LUT2 #(
		.INIT('h8)
	) name15899 (
		\wishbone_bd_ram_mem1_reg[236][8]/P0001 ,
		_w12731_,
		_w26411_
	);
	LUT2 #(
		.INIT('h8)
	) name15900 (
		\wishbone_bd_ram_mem1_reg[144][8]/P0001 ,
		_w12756_,
		_w26412_
	);
	LUT2 #(
		.INIT('h8)
	) name15901 (
		\wishbone_bd_ram_mem1_reg[186][8]/P0001 ,
		_w12783_,
		_w26413_
	);
	LUT2 #(
		.INIT('h8)
	) name15902 (
		\wishbone_bd_ram_mem1_reg[131][8]/P0001 ,
		_w12852_,
		_w26414_
	);
	LUT2 #(
		.INIT('h8)
	) name15903 (
		\wishbone_bd_ram_mem1_reg[143][8]/P0001 ,
		_w12922_,
		_w26415_
	);
	LUT2 #(
		.INIT('h8)
	) name15904 (
		\wishbone_bd_ram_mem1_reg[193][8]/P0001 ,
		_w13056_,
		_w26416_
	);
	LUT2 #(
		.INIT('h8)
	) name15905 (
		\wishbone_bd_ram_mem1_reg[237][8]/P0001 ,
		_w12990_,
		_w26417_
	);
	LUT2 #(
		.INIT('h8)
	) name15906 (
		\wishbone_bd_ram_mem1_reg[59][8]/P0001 ,
		_w12780_,
		_w26418_
	);
	LUT2 #(
		.INIT('h8)
	) name15907 (
		\wishbone_bd_ram_mem1_reg[184][8]/P0001 ,
		_w13062_,
		_w26419_
	);
	LUT2 #(
		.INIT('h8)
	) name15908 (
		\wishbone_bd_ram_mem1_reg[95][8]/P0001 ,
		_w12844_,
		_w26420_
	);
	LUT2 #(
		.INIT('h8)
	) name15909 (
		\wishbone_bd_ram_mem1_reg[168][8]/P0001 ,
		_w13208_,
		_w26421_
	);
	LUT2 #(
		.INIT('h8)
	) name15910 (
		\wishbone_bd_ram_mem1_reg[221][8]/P0001 ,
		_w12802_,
		_w26422_
	);
	LUT2 #(
		.INIT('h8)
	) name15911 (
		\wishbone_bd_ram_mem1_reg[25][8]/P0001 ,
		_w13108_,
		_w26423_
	);
	LUT2 #(
		.INIT('h8)
	) name15912 (
		\wishbone_bd_ram_mem1_reg[218][8]/P0001 ,
		_w13206_,
		_w26424_
	);
	LUT2 #(
		.INIT('h8)
	) name15913 (
		\wishbone_bd_ram_mem1_reg[119][8]/P0001 ,
		_w13048_,
		_w26425_
	);
	LUT2 #(
		.INIT('h8)
	) name15914 (
		\wishbone_bd_ram_mem1_reg[138][8]/P0001 ,
		_w12958_,
		_w26426_
	);
	LUT2 #(
		.INIT('h8)
	) name15915 (
		\wishbone_bd_ram_mem1_reg[241][8]/P0001 ,
		_w13006_,
		_w26427_
	);
	LUT2 #(
		.INIT('h8)
	) name15916 (
		\wishbone_bd_ram_mem1_reg[36][8]/P0001 ,
		_w12800_,
		_w26428_
	);
	LUT2 #(
		.INIT('h8)
	) name15917 (
		\wishbone_bd_ram_mem1_reg[200][8]/P0001 ,
		_w12988_,
		_w26429_
	);
	LUT2 #(
		.INIT('h8)
	) name15918 (
		\wishbone_bd_ram_mem1_reg[249][8]/P0001 ,
		_w12900_,
		_w26430_
	);
	LUT2 #(
		.INIT('h8)
	) name15919 (
		\wishbone_bd_ram_mem1_reg[151][8]/P0001 ,
		_w13142_,
		_w26431_
	);
	LUT2 #(
		.INIT('h8)
	) name15920 (
		\wishbone_bd_ram_mem1_reg[157][8]/P0001 ,
		_w12926_,
		_w26432_
	);
	LUT2 #(
		.INIT('h8)
	) name15921 (
		\wishbone_bd_ram_mem1_reg[58][8]/P0001 ,
		_w13070_,
		_w26433_
	);
	LUT2 #(
		.INIT('h8)
	) name15922 (
		\wishbone_bd_ram_mem1_reg[123][8]/P0001 ,
		_w13114_,
		_w26434_
	);
	LUT2 #(
		.INIT('h8)
	) name15923 (
		\wishbone_bd_ram_mem1_reg[75][8]/P0001 ,
		_w12826_,
		_w26435_
	);
	LUT2 #(
		.INIT('h8)
	) name15924 (
		\wishbone_bd_ram_mem1_reg[215][8]/P0001 ,
		_w12974_,
		_w26436_
	);
	LUT2 #(
		.INIT('h8)
	) name15925 (
		\wishbone_bd_ram_mem1_reg[205][8]/P0001 ,
		_w13068_,
		_w26437_
	);
	LUT2 #(
		.INIT('h8)
	) name15926 (
		\wishbone_bd_ram_mem1_reg[201][8]/P0001 ,
		_w12822_,
		_w26438_
	);
	LUT2 #(
		.INIT('h8)
	) name15927 (
		\wishbone_bd_ram_mem1_reg[1][8]/P0001 ,
		_w13014_,
		_w26439_
	);
	LUT2 #(
		.INIT('h8)
	) name15928 (
		\wishbone_bd_ram_mem1_reg[96][8]/P0001 ,
		_w12912_,
		_w26440_
	);
	LUT2 #(
		.INIT('h8)
	) name15929 (
		\wishbone_bd_ram_mem1_reg[165][8]/P0001 ,
		_w13044_,
		_w26441_
	);
	LUT2 #(
		.INIT('h8)
	) name15930 (
		\wishbone_bd_ram_mem1_reg[10][8]/P0001 ,
		_w13172_,
		_w26442_
	);
	LUT2 #(
		.INIT('h8)
	) name15931 (
		\wishbone_bd_ram_mem1_reg[125][8]/P0001 ,
		_w12956_,
		_w26443_
	);
	LUT2 #(
		.INIT('h8)
	) name15932 (
		\wishbone_bd_ram_mem1_reg[140][8]/P0001 ,
		_w12894_,
		_w26444_
	);
	LUT2 #(
		.INIT('h8)
	) name15933 (
		\wishbone_bd_ram_mem1_reg[121][8]/P0001 ,
		_w13078_,
		_w26445_
	);
	LUT2 #(
		.INIT('h8)
	) name15934 (
		\wishbone_bd_ram_mem1_reg[254][8]/P0001 ,
		_w12892_,
		_w26446_
	);
	LUT2 #(
		.INIT('h8)
	) name15935 (
		\wishbone_bd_ram_mem1_reg[101][8]/P0001 ,
		_w13192_,
		_w26447_
	);
	LUT2 #(
		.INIT('h8)
	) name15936 (
		\wishbone_bd_ram_mem1_reg[162][8]/P0001 ,
		_w13098_,
		_w26448_
	);
	LUT2 #(
		.INIT('h8)
	) name15937 (
		\wishbone_bd_ram_mem1_reg[213][8]/P0001 ,
		_w13002_,
		_w26449_
	);
	LUT2 #(
		.INIT('h8)
	) name15938 (
		\wishbone_bd_ram_mem1_reg[161][8]/P0001 ,
		_w12754_,
		_w26450_
	);
	LUT2 #(
		.INIT('h8)
	) name15939 (
		\wishbone_bd_ram_mem1_reg[163][8]/P0001 ,
		_w12882_,
		_w26451_
	);
	LUT2 #(
		.INIT('h8)
	) name15940 (
		\wishbone_bd_ram_mem1_reg[185][8]/P0001 ,
		_w12940_,
		_w26452_
	);
	LUT2 #(
		.INIT('h8)
	) name15941 (
		\wishbone_bd_ram_mem1_reg[229][8]/P0001 ,
		_w12711_,
		_w26453_
	);
	LUT2 #(
		.INIT('h8)
	) name15942 (
		\wishbone_bd_ram_mem1_reg[127][8]/P0001 ,
		_w13164_,
		_w26454_
	);
	LUT2 #(
		.INIT('h8)
	) name15943 (
		\wishbone_bd_ram_mem1_reg[46][8]/P0001 ,
		_w12884_,
		_w26455_
	);
	LUT2 #(
		.INIT('h8)
	) name15944 (
		\wishbone_bd_ram_mem1_reg[44][8]/P0001 ,
		_w12896_,
		_w26456_
	);
	LUT2 #(
		.INIT('h8)
	) name15945 (
		\wishbone_bd_ram_mem1_reg[145][8]/P0001 ,
		_w13106_,
		_w26457_
	);
	LUT2 #(
		.INIT('h8)
	) name15946 (
		\wishbone_bd_ram_mem1_reg[174][8]/P0001 ,
		_w12972_,
		_w26458_
	);
	LUT2 #(
		.INIT('h8)
	) name15947 (
		\wishbone_bd_ram_mem1_reg[42][8]/P0001 ,
		_w12842_,
		_w26459_
	);
	LUT2 #(
		.INIT('h8)
	) name15948 (
		\wishbone_bd_ram_mem1_reg[117][8]/P0001 ,
		_w12715_,
		_w26460_
	);
	LUT2 #(
		.INIT('h8)
	) name15949 (
		\wishbone_bd_ram_mem1_reg[18][8]/P0001 ,
		_w12679_,
		_w26461_
	);
	LUT2 #(
		.INIT('h8)
	) name15950 (
		\wishbone_bd_ram_mem1_reg[211][8]/P0001 ,
		_w13166_,
		_w26462_
	);
	LUT2 #(
		.INIT('h8)
	) name15951 (
		\wishbone_bd_ram_mem1_reg[171][8]/P0001 ,
		_w12910_,
		_w26463_
	);
	LUT2 #(
		.INIT('h8)
	) name15952 (
		\wishbone_bd_ram_mem1_reg[48][8]/P0001 ,
		_w12970_,
		_w26464_
	);
	LUT2 #(
		.INIT('h8)
	) name15953 (
		\wishbone_bd_ram_mem1_reg[180][8]/P0001 ,
		_w12791_,
		_w26465_
	);
	LUT2 #(
		.INIT('h8)
	) name15954 (
		\wishbone_bd_ram_mem1_reg[178][8]/P0001 ,
		_w12886_,
		_w26466_
	);
	LUT2 #(
		.INIT('h8)
	) name15955 (
		\wishbone_bd_ram_mem1_reg[252][8]/P0001 ,
		_w13080_,
		_w26467_
	);
	LUT2 #(
		.INIT('h8)
	) name15956 (
		\wishbone_bd_ram_mem1_reg[5][8]/P0001 ,
		_w12878_,
		_w26468_
	);
	LUT2 #(
		.INIT('h8)
	) name15957 (
		\wishbone_bd_ram_mem1_reg[92][8]/P0001 ,
		_w13010_,
		_w26469_
	);
	LUT2 #(
		.INIT('h8)
	) name15958 (
		\wishbone_bd_ram_mem1_reg[232][8]/P0001 ,
		_w12758_,
		_w26470_
	);
	LUT2 #(
		.INIT('h8)
	) name15959 (
		\wishbone_bd_ram_mem1_reg[118][8]/P0001 ,
		_w12830_,
		_w26471_
	);
	LUT2 #(
		.INIT('h8)
	) name15960 (
		\wishbone_bd_ram_mem1_reg[4][8]/P0001 ,
		_w12666_,
		_w26472_
	);
	LUT2 #(
		.INIT('h8)
	) name15961 (
		\wishbone_bd_ram_mem1_reg[239][8]/P0001 ,
		_w12862_,
		_w26473_
	);
	LUT2 #(
		.INIT('h8)
	) name15962 (
		\wishbone_bd_ram_mem1_reg[33][8]/P0001 ,
		_w12980_,
		_w26474_
	);
	LUT2 #(
		.INIT('h8)
	) name15963 (
		\wishbone_bd_ram_mem1_reg[72][8]/P0001 ,
		_w12810_,
		_w26475_
	);
	LUT2 #(
		.INIT('h8)
	) name15964 (
		\wishbone_bd_ram_mem1_reg[223][8]/P0001 ,
		_w12838_,
		_w26476_
	);
	LUT2 #(
		.INIT('h8)
	) name15965 (
		\wishbone_bd_ram_mem1_reg[35][8]/P0001 ,
		_w12703_,
		_w26477_
	);
	LUT2 #(
		.INIT('h8)
	) name15966 (
		\wishbone_bd_ram_mem1_reg[226][8]/P0001 ,
		_w13138_,
		_w26478_
	);
	LUT2 #(
		.INIT('h8)
	) name15967 (
		\wishbone_bd_ram_mem1_reg[66][8]/P0001 ,
		_w12824_,
		_w26479_
	);
	LUT2 #(
		.INIT('h8)
	) name15968 (
		\wishbone_bd_ram_mem1_reg[89][8]/P0001 ,
		_w12964_,
		_w26480_
	);
	LUT2 #(
		.INIT('h8)
	) name15969 (
		\wishbone_bd_ram_mem1_reg[190][8]/P0001 ,
		_w12858_,
		_w26481_
	);
	LUT2 #(
		.INIT('h8)
	) name15970 (
		\wishbone_bd_ram_mem1_reg[43][8]/P0001 ,
		_w13200_,
		_w26482_
	);
	LUT2 #(
		.INIT('h8)
	) name15971 (
		\wishbone_bd_ram_mem1_reg[57][8]/P0001 ,
		_w13116_,
		_w26483_
	);
	LUT2 #(
		.INIT('h8)
	) name15972 (
		\wishbone_bd_ram_mem1_reg[188][8]/P0001 ,
		_w12948_,
		_w26484_
	);
	LUT2 #(
		.INIT('h8)
	) name15973 (
		\wishbone_bd_ram_mem1_reg[181][8]/P0001 ,
		_w12828_,
		_w26485_
	);
	LUT2 #(
		.INIT('h8)
	) name15974 (
		\wishbone_bd_ram_mem1_reg[113][8]/P0001 ,
		_w13026_,
		_w26486_
	);
	LUT2 #(
		.INIT('h8)
	) name15975 (
		\wishbone_bd_ram_mem1_reg[85][8]/P0001 ,
		_w13216_,
		_w26487_
	);
	LUT2 #(
		.INIT('h8)
	) name15976 (
		\wishbone_bd_ram_mem1_reg[30][8]/P0001 ,
		_w13104_,
		_w26488_
	);
	LUT2 #(
		.INIT('h8)
	) name15977 (
		\wishbone_bd_ram_mem1_reg[129][8]/P0001 ,
		_w12776_,
		_w26489_
	);
	LUT2 #(
		.INIT('h8)
	) name15978 (
		\wishbone_bd_ram_mem1_reg[104][8]/P0001 ,
		_w13148_,
		_w26490_
	);
	LUT2 #(
		.INIT('h8)
	) name15979 (
		\wishbone_bd_ram_mem1_reg[107][8]/P0001 ,
		_w12749_,
		_w26491_
	);
	LUT2 #(
		.INIT('h8)
	) name15980 (
		\wishbone_bd_ram_mem1_reg[231][8]/P0001 ,
		_w12856_,
		_w26492_
	);
	LUT2 #(
		.INIT('h8)
	) name15981 (
		\wishbone_bd_ram_mem1_reg[159][8]/P0001 ,
		_w12774_,
		_w26493_
	);
	LUT2 #(
		.INIT('h8)
	) name15982 (
		\wishbone_bd_ram_mem1_reg[240][8]/P0001 ,
		_w12864_,
		_w26494_
	);
	LUT2 #(
		.INIT('h8)
	) name15983 (
		\wishbone_bd_ram_mem1_reg[16][8]/P0001 ,
		_w13140_,
		_w26495_
	);
	LUT2 #(
		.INIT('h8)
	) name15984 (
		\wishbone_bd_ram_mem1_reg[68][8]/P0001 ,
		_w12946_,
		_w26496_
	);
	LUT2 #(
		.INIT('h8)
	) name15985 (
		\wishbone_bd_ram_mem1_reg[202][8]/P0001 ,
		_w12870_,
		_w26497_
	);
	LUT2 #(
		.INIT('h8)
	) name15986 (
		\wishbone_bd_ram_mem1_reg[86][8]/P0001 ,
		_w12735_,
		_w26498_
	);
	LUT2 #(
		.INIT('h8)
	) name15987 (
		\wishbone_bd_ram_mem1_reg[137][8]/P0001 ,
		_w13168_,
		_w26499_
	);
	LUT2 #(
		.INIT('h8)
	) name15988 (
		\wishbone_bd_ram_mem1_reg[29][8]/P0001 ,
		_w12952_,
		_w26500_
	);
	LUT2 #(
		.INIT('h8)
	) name15989 (
		\wishbone_bd_ram_mem1_reg[204][8]/P0001 ,
		_w13162_,
		_w26501_
	);
	LUT2 #(
		.INIT('h8)
	) name15990 (
		\wishbone_bd_ram_mem1_reg[160][8]/P0001 ,
		_w12872_,
		_w26502_
	);
	LUT2 #(
		.INIT('h8)
	) name15991 (
		\wishbone_bd_ram_mem1_reg[97][8]/P0001 ,
		_w13096_,
		_w26503_
	);
	LUT2 #(
		.INIT('h8)
	) name15992 (
		\wishbone_bd_ram_mem1_reg[120][8]/P0001 ,
		_w12707_,
		_w26504_
	);
	LUT2 #(
		.INIT('h8)
	) name15993 (
		\wishbone_bd_ram_mem1_reg[255][8]/P0001 ,
		_w13072_,
		_w26505_
	);
	LUT2 #(
		.INIT('h8)
	) name15994 (
		\wishbone_bd_ram_mem1_reg[111][8]/P0001 ,
		_w12744_,
		_w26506_
	);
	LUT2 #(
		.INIT('h8)
	) name15995 (
		\wishbone_bd_ram_mem1_reg[210][8]/P0001 ,
		_w12924_,
		_w26507_
	);
	LUT2 #(
		.INIT('h8)
	) name15996 (
		\wishbone_bd_ram_mem1_reg[19][8]/P0001 ,
		_w13012_,
		_w26508_
	);
	LUT2 #(
		.INIT('h8)
	) name15997 (
		\wishbone_bd_ram_mem1_reg[198][8]/P0001 ,
		_w12832_,
		_w26509_
	);
	LUT2 #(
		.INIT('h8)
	) name15998 (
		\wishbone_bd_ram_mem1_reg[32][8]/P0001 ,
		_w13120_,
		_w26510_
	);
	LUT2 #(
		.INIT('h8)
	) name15999 (
		\wishbone_bd_ram_mem1_reg[49][8]/P0001 ,
		_w12994_,
		_w26511_
	);
	LUT2 #(
		.INIT('h8)
	) name16000 (
		\wishbone_bd_ram_mem1_reg[251][8]/P0001 ,
		_w13054_,
		_w26512_
	);
	LUT2 #(
		.INIT('h8)
	) name16001 (
		\wishbone_bd_ram_mem1_reg[156][8]/P0001 ,
		_w13190_,
		_w26513_
	);
	LUT2 #(
		.INIT('h8)
	) name16002 (
		\wishbone_bd_ram_mem1_reg[31][8]/P0001 ,
		_w13198_,
		_w26514_
	);
	LUT2 #(
		.INIT('h8)
	) name16003 (
		\wishbone_bd_ram_mem1_reg[99][8]/P0001 ,
		_w13038_,
		_w26515_
	);
	LUT2 #(
		.INIT('h8)
	) name16004 (
		\wishbone_bd_ram_mem1_reg[91][8]/P0001 ,
		_w13074_,
		_w26516_
	);
	LUT2 #(
		.INIT('h8)
	) name16005 (
		\wishbone_bd_ram_mem1_reg[39][8]/P0001 ,
		_w13018_,
		_w26517_
	);
	LUT2 #(
		.INIT('h8)
	) name16006 (
		\wishbone_bd_ram_mem1_reg[82][8]/P0001 ,
		_w12942_,
		_w26518_
	);
	LUT2 #(
		.INIT('h8)
	) name16007 (
		\wishbone_bd_ram_mem1_reg[22][8]/P0001 ,
		_w13110_,
		_w26519_
	);
	LUT2 #(
		.INIT('h8)
	) name16008 (
		\wishbone_bd_ram_mem1_reg[28][8]/P0001 ,
		_w13170_,
		_w26520_
	);
	LUT2 #(
		.INIT('h8)
	) name16009 (
		\wishbone_bd_ram_mem1_reg[77][8]/P0001 ,
		_w12982_,
		_w26521_
	);
	LUT2 #(
		.INIT('h8)
	) name16010 (
		\wishbone_bd_ram_mem1_reg[217][8]/P0001 ,
		_w13188_,
		_w26522_
	);
	LUT2 #(
		.INIT('h8)
	) name16011 (
		\wishbone_bd_ram_mem1_reg[20][8]/P0001 ,
		_w13174_,
		_w26523_
	);
	LUT2 #(
		.INIT('h8)
	) name16012 (
		\wishbone_bd_ram_mem1_reg[88][8]/P0001 ,
		_w12860_,
		_w26524_
	);
	LUT2 #(
		.INIT('h8)
	) name16013 (
		\wishbone_bd_ram_mem1_reg[69][8]/P0001 ,
		_w12738_,
		_w26525_
	);
	LUT2 #(
		.INIT('h8)
	) name16014 (
		\wishbone_bd_ram_mem1_reg[60][8]/P0001 ,
		_w13204_,
		_w26526_
	);
	LUT2 #(
		.INIT('h8)
	) name16015 (
		\wishbone_bd_ram_mem1_reg[233][8]/P0001 ,
		_w12836_,
		_w26527_
	);
	LUT2 #(
		.INIT('h8)
	) name16016 (
		\wishbone_bd_ram_mem1_reg[122][8]/P0001 ,
		_w13130_,
		_w26528_
	);
	LUT2 #(
		.INIT('h8)
	) name16017 (
		\wishbone_bd_ram_mem1_reg[199][8]/P0001 ,
		_w12768_,
		_w26529_
	);
	LUT2 #(
		.INIT('h8)
	) name16018 (
		\wishbone_bd_ram_mem1_reg[234][8]/P0001 ,
		_w13214_,
		_w26530_
	);
	LUT2 #(
		.INIT('h8)
	) name16019 (
		\wishbone_bd_ram_mem1_reg[154][8]/P0001 ,
		_w12962_,
		_w26531_
	);
	LUT2 #(
		.INIT('h8)
	) name16020 (
		\wishbone_bd_ram_mem1_reg[141][8]/P0001 ,
		_w13004_,
		_w26532_
	);
	LUT2 #(
		.INIT('h8)
	) name16021 (
		\wishbone_bd_ram_mem1_reg[102][8]/P0001 ,
		_w12685_,
		_w26533_
	);
	LUT2 #(
		.INIT('h8)
	) name16022 (
		\wishbone_bd_ram_mem1_reg[53][8]/P0001 ,
		_w13020_,
		_w26534_
	);
	LUT2 #(
		.INIT('h8)
	) name16023 (
		\wishbone_bd_ram_mem1_reg[80][8]/P0001 ,
		_w12689_,
		_w26535_
	);
	LUT2 #(
		.INIT('h8)
	) name16024 (
		\wishbone_bd_ram_mem1_reg[70][8]/P0001 ,
		_w12840_,
		_w26536_
	);
	LUT2 #(
		.INIT('h8)
	) name16025 (
		\wishbone_bd_ram_mem1_reg[34][8]/P0001 ,
		_w12930_,
		_w26537_
	);
	LUT2 #(
		.INIT('h8)
	) name16026 (
		\wishbone_bd_ram_mem1_reg[139][8]/P0001 ,
		_w12814_,
		_w26538_
	);
	LUT2 #(
		.INIT('h8)
	) name16027 (
		\wishbone_bd_ram_mem1_reg[45][8]/P0001 ,
		_w12908_,
		_w26539_
	);
	LUT2 #(
		.INIT('h8)
	) name16028 (
		\wishbone_bd_ram_mem1_reg[100][8]/P0001 ,
		_w12960_,
		_w26540_
	);
	LUT2 #(
		.INIT('h8)
	) name16029 (
		\wishbone_bd_ram_mem1_reg[14][8]/P0001 ,
		_w13086_,
		_w26541_
	);
	LUT2 #(
		.INIT('h8)
	) name16030 (
		\wishbone_bd_ram_mem1_reg[13][8]/P0001 ,
		_w13178_,
		_w26542_
	);
	LUT2 #(
		.INIT('h8)
	) name16031 (
		\wishbone_bd_ram_mem1_reg[216][8]/P0001 ,
		_w13028_,
		_w26543_
	);
	LUT2 #(
		.INIT('h8)
	) name16032 (
		\wishbone_bd_ram_mem1_reg[26][8]/P0001 ,
		_w12699_,
		_w26544_
	);
	LUT2 #(
		.INIT('h8)
	) name16033 (
		\wishbone_bd_ram_mem1_reg[142][8]/P0001 ,
		_w12928_,
		_w26545_
	);
	LUT2 #(
		.INIT('h8)
	) name16034 (
		\wishbone_bd_ram_mem1_reg[169][8]/P0001 ,
		_w12722_,
		_w26546_
	);
	LUT2 #(
		.INIT('h8)
	) name16035 (
		\wishbone_bd_ram_mem1_reg[74][8]/P0001 ,
		_w12812_,
		_w26547_
	);
	LUT2 #(
		.INIT('h8)
	) name16036 (
		\wishbone_bd_ram_mem1_reg[212][8]/P0001 ,
		_w12796_,
		_w26548_
	);
	LUT2 #(
		.INIT('h8)
	) name16037 (
		\wishbone_bd_ram_mem1_reg[12][8]/P0001 ,
		_w13118_,
		_w26549_
	);
	LUT2 #(
		.INIT('h8)
	) name16038 (
		\wishbone_bd_ram_mem1_reg[62][8]/P0001 ,
		_w12673_,
		_w26550_
	);
	LUT2 #(
		.INIT('h8)
	) name16039 (
		\wishbone_bd_ram_mem1_reg[155][8]/P0001 ,
		_w13122_,
		_w26551_
	);
	LUT2 #(
		.INIT('h8)
	) name16040 (
		\wishbone_bd_ram_mem1_reg[247][8]/P0001 ,
		_w12818_,
		_w26552_
	);
	LUT2 #(
		.INIT('h8)
	) name16041 (
		\wishbone_bd_ram_mem1_reg[182][8]/P0001 ,
		_w12820_,
		_w26553_
	);
	LUT2 #(
		.INIT('h8)
	) name16042 (
		\wishbone_bd_ram_mem1_reg[136][8]/P0001 ,
		_w13064_,
		_w26554_
	);
	LUT2 #(
		.INIT('h8)
	) name16043 (
		\wishbone_bd_ram_mem1_reg[195][8]/P0001 ,
		_w13144_,
		_w26555_
	);
	LUT2 #(
		.INIT('h8)
	) name16044 (
		\wishbone_bd_ram_mem1_reg[108][8]/P0001 ,
		_w13156_,
		_w26556_
	);
	LUT2 #(
		.INIT('h8)
	) name16045 (
		\wishbone_bd_ram_mem1_reg[134][8]/P0001 ,
		_w12763_,
		_w26557_
	);
	LUT2 #(
		.INIT('h8)
	) name16046 (
		\wishbone_bd_ram_mem1_reg[176][8]/P0001 ,
		_w12868_,
		_w26558_
	);
	LUT2 #(
		.INIT('h8)
	) name16047 (
		\wishbone_bd_ram_mem1_reg[24][8]/P0001 ,
		_w13084_,
		_w26559_
	);
	LUT2 #(
		.INIT('h8)
	) name16048 (
		\wishbone_bd_ram_mem1_reg[220][8]/P0001 ,
		_w13066_,
		_w26560_
	);
	LUT2 #(
		.INIT('h8)
	) name16049 (
		\wishbone_bd_ram_mem1_reg[76][8]/P0001 ,
		_w13184_,
		_w26561_
	);
	LUT2 #(
		.INIT('h8)
	) name16050 (
		\wishbone_bd_ram_mem1_reg[87][8]/P0001 ,
		_w13154_,
		_w26562_
	);
	LUT2 #(
		.INIT('h8)
	) name16051 (
		\wishbone_bd_ram_mem1_reg[132][8]/P0001 ,
		_w12992_,
		_w26563_
	);
	LUT2 #(
		.INIT('h8)
	) name16052 (
		\wishbone_bd_ram_mem1_reg[196][8]/P0001 ,
		_w13090_,
		_w26564_
	);
	LUT2 #(
		.INIT('h8)
	) name16053 (
		\wishbone_bd_ram_mem1_reg[192][8]/P0001 ,
		_w12938_,
		_w26565_
	);
	LUT2 #(
		.INIT('h8)
	) name16054 (
		\wishbone_bd_ram_mem1_reg[94][8]/P0001 ,
		_w13186_,
		_w26566_
	);
	LUT2 #(
		.INIT('h8)
	) name16055 (
		\wishbone_bd_ram_mem1_reg[248][8]/P0001 ,
		_w12789_,
		_w26567_
	);
	LUT2 #(
		.INIT('h8)
	) name16056 (
		\wishbone_bd_ram_mem1_reg[175][8]/P0001 ,
		_w13126_,
		_w26568_
	);
	LUT2 #(
		.INIT('h8)
	) name16057 (
		\wishbone_bd_ram_mem1_reg[179][8]/P0001 ,
		_w13050_,
		_w26569_
	);
	LUT2 #(
		.INIT('h8)
	) name16058 (
		\wishbone_bd_ram_mem1_reg[40][8]/P0001 ,
		_w13132_,
		_w26570_
	);
	LUT2 #(
		.INIT('h8)
	) name16059 (
		\wishbone_bd_ram_mem1_reg[244][8]/P0001 ,
		_w12747_,
		_w26571_
	);
	LUT2 #(
		.INIT('h8)
	) name16060 (
		\wishbone_bd_ram_mem1_reg[63][8]/P0001 ,
		_w12850_,
		_w26572_
	);
	LUT2 #(
		.INIT('h8)
	) name16061 (
		\wishbone_bd_ram_mem1_reg[194][8]/P0001 ,
		_w12772_,
		_w26573_
	);
	LUT2 #(
		.INIT('h8)
	) name16062 (
		\wishbone_bd_ram_mem1_reg[153][8]/P0001 ,
		_w12890_,
		_w26574_
	);
	LUT2 #(
		.INIT('h8)
	) name16063 (
		\wishbone_bd_ram_mem1_reg[206][8]/P0001 ,
		_w12954_,
		_w26575_
	);
	LUT2 #(
		.INIT('h8)
	) name16064 (
		\wishbone_bd_ram_mem1_reg[17][8]/P0001 ,
		_w12848_,
		_w26576_
	);
	LUT2 #(
		.INIT('h8)
	) name16065 (
		\wishbone_bd_ram_mem1_reg[0][8]/P0001 ,
		_w12717_,
		_w26577_
	);
	LUT2 #(
		.INIT('h8)
	) name16066 (
		\wishbone_bd_ram_mem1_reg[23][8]/P0001 ,
		_w13008_,
		_w26578_
	);
	LUT2 #(
		.INIT('h8)
	) name16067 (
		\wishbone_bd_ram_mem1_reg[37][8]/P0001 ,
		_w13102_,
		_w26579_
	);
	LUT2 #(
		.INIT('h8)
	) name16068 (
		\wishbone_bd_ram_mem1_reg[112][8]/P0001 ,
		_w12733_,
		_w26580_
	);
	LUT2 #(
		.INIT('h8)
	) name16069 (
		\wishbone_bd_ram_mem1_reg[250][8]/P0001 ,
		_w13128_,
		_w26581_
	);
	LUT2 #(
		.INIT('h8)
	) name16070 (
		\wishbone_bd_ram_mem1_reg[110][8]/P0001 ,
		_w13046_,
		_w26582_
	);
	LUT2 #(
		.INIT('h8)
	) name16071 (
		\wishbone_bd_ram_mem1_reg[222][8]/P0001 ,
		_w13094_,
		_w26583_
	);
	LUT2 #(
		.INIT('h8)
	) name16072 (
		\wishbone_bd_ram_mem1_reg[158][8]/P0001 ,
		_w12898_,
		_w26584_
	);
	LUT2 #(
		.INIT('h8)
	) name16073 (
		\wishbone_bd_ram_mem1_reg[246][8]/P0001 ,
		_w13076_,
		_w26585_
	);
	LUT2 #(
		.INIT('h8)
	) name16074 (
		\wishbone_bd_ram_mem1_reg[65][8]/P0001 ,
		_w13176_,
		_w26586_
	);
	LUT2 #(
		.INIT('h8)
	) name16075 (
		\wishbone_bd_ram_mem1_reg[64][8]/P0001 ,
		_w12976_,
		_w26587_
	);
	LUT2 #(
		.INIT('h8)
	) name16076 (
		\wishbone_bd_ram_mem1_reg[103][8]/P0001 ,
		_w12846_,
		_w26588_
	);
	LUT2 #(
		.INIT('h8)
	) name16077 (
		\wishbone_bd_ram_mem1_reg[109][8]/P0001 ,
		_w12888_,
		_w26589_
	);
	LUT2 #(
		.INIT('h8)
	) name16078 (
		\wishbone_bd_ram_mem1_reg[219][8]/P0001 ,
		_w12806_,
		_w26590_
	);
	LUT2 #(
		.INIT('h8)
	) name16079 (
		\wishbone_bd_ram_mem1_reg[71][8]/P0001 ,
		_w12798_,
		_w26591_
	);
	LUT2 #(
		.INIT('h8)
	) name16080 (
		\wishbone_bd_ram_mem1_reg[54][8]/P0001 ,
		_w12770_,
		_w26592_
	);
	LUT2 #(
		.INIT('h8)
	) name16081 (
		\wishbone_bd_ram_mem1_reg[149][8]/P0001 ,
		_w12741_,
		_w26593_
	);
	LUT2 #(
		.INIT('h8)
	) name16082 (
		\wishbone_bd_ram_mem1_reg[8][8]/P0001 ,
		_w12920_,
		_w26594_
	);
	LUT2 #(
		.INIT('h8)
	) name16083 (
		\wishbone_bd_ram_mem1_reg[11][8]/P0001 ,
		_w13194_,
		_w26595_
	);
	LUT2 #(
		.INIT('h8)
	) name16084 (
		\wishbone_bd_ram_mem1_reg[55][8]/P0001 ,
		_w12785_,
		_w26596_
	);
	LUT2 #(
		.INIT('h8)
	) name16085 (
		\wishbone_bd_ram_mem1_reg[126][8]/P0001 ,
		_w13218_,
		_w26597_
	);
	LUT2 #(
		.INIT('h8)
	) name16086 (
		\wishbone_bd_ram_mem1_reg[209][8]/P0001 ,
		_w13152_,
		_w26598_
	);
	LUT2 #(
		.INIT('h8)
	) name16087 (
		\wishbone_bd_ram_mem1_reg[245][8]/P0001 ,
		_w13022_,
		_w26599_
	);
	LUT2 #(
		.INIT('h8)
	) name16088 (
		\wishbone_bd_ram_mem1_reg[208][8]/P0001 ,
		_w13032_,
		_w26600_
	);
	LUT2 #(
		.INIT('h8)
	) name16089 (
		\wishbone_bd_ram_mem1_reg[21][8]/P0001 ,
		_w12906_,
		_w26601_
	);
	LUT2 #(
		.INIT('h8)
	) name16090 (
		\wishbone_bd_ram_mem1_reg[164][8]/P0001 ,
		_w12876_,
		_w26602_
	);
	LUT2 #(
		.INIT('h8)
	) name16091 (
		\wishbone_bd_ram_mem1_reg[81][8]/P0001 ,
		_w12950_,
		_w26603_
	);
	LUT2 #(
		.INIT('h8)
	) name16092 (
		\wishbone_bd_ram_mem1_reg[187][8]/P0001 ,
		_w13196_,
		_w26604_
	);
	LUT2 #(
		.INIT('h8)
	) name16093 (
		\wishbone_bd_ram_mem1_reg[38][8]/P0001 ,
		_w13182_,
		_w26605_
	);
	LUT2 #(
		.INIT('h8)
	) name16094 (
		\wishbone_bd_ram_mem1_reg[230][8]/P0001 ,
		_w13036_,
		_w26606_
	);
	LUT2 #(
		.INIT('h8)
	) name16095 (
		\wishbone_bd_ram_mem1_reg[124][8]/P0001 ,
		_w13058_,
		_w26607_
	);
	LUT2 #(
		.INIT('h8)
	) name16096 (
		\wishbone_bd_ram_mem1_reg[73][8]/P0001 ,
		_w12918_,
		_w26608_
	);
	LUT2 #(
		.INIT('h8)
	) name16097 (
		\wishbone_bd_ram_mem1_reg[146][8]/P0001 ,
		_w13060_,
		_w26609_
	);
	LUT2 #(
		.INIT('h8)
	) name16098 (
		\wishbone_bd_ram_mem1_reg[67][8]/P0001 ,
		_w13134_,
		_w26610_
	);
	LUT2 #(
		.INIT('h8)
	) name16099 (
		\wishbone_bd_ram_mem1_reg[183][8]/P0001 ,
		_w12787_,
		_w26611_
	);
	LUT2 #(
		.INIT('h8)
	) name16100 (
		\wishbone_bd_ram_mem1_reg[167][8]/P0001 ,
		_w12986_,
		_w26612_
	);
	LUT2 #(
		.INIT('h8)
	) name16101 (
		\wishbone_bd_ram_mem1_reg[130][8]/P0001 ,
		_w12914_,
		_w26613_
	);
	LUT2 #(
		.INIT('h8)
	) name16102 (
		\wishbone_bd_ram_mem1_reg[243][8]/P0001 ,
		_w12804_,
		_w26614_
	);
	LUT2 #(
		.INIT('h8)
	) name16103 (
		\wishbone_bd_ram_mem1_reg[227][8]/P0001 ,
		_w12936_,
		_w26615_
	);
	LUT2 #(
		.INIT('h8)
	) name16104 (
		\wishbone_bd_ram_mem1_reg[235][8]/P0001 ,
		_w12696_,
		_w26616_
	);
	LUT2 #(
		.INIT('h8)
	) name16105 (
		\wishbone_bd_ram_mem1_reg[197][8]/P0001 ,
		_w12834_,
		_w26617_
	);
	LUT2 #(
		.INIT('h8)
	) name16106 (
		\wishbone_bd_ram_mem1_reg[203][8]/P0001 ,
		_w13158_,
		_w26618_
	);
	LUT2 #(
		.INIT('h8)
	) name16107 (
		\wishbone_bd_ram_mem1_reg[116][8]/P0001 ,
		_w12998_,
		_w26619_
	);
	LUT2 #(
		.INIT('h8)
	) name16108 (
		\wishbone_bd_ram_mem1_reg[6][8]/P0001 ,
		_w12968_,
		_w26620_
	);
	LUT2 #(
		.INIT('h8)
	) name16109 (
		\wishbone_bd_ram_mem1_reg[15][8]/P0001 ,
		_w13210_,
		_w26621_
	);
	LUT2 #(
		.INIT('h8)
	) name16110 (
		\wishbone_bd_ram_mem1_reg[47][8]/P0001 ,
		_w12904_,
		_w26622_
	);
	LUT2 #(
		.INIT('h8)
	) name16111 (
		\wishbone_bd_ram_mem1_reg[114][8]/P0001 ,
		_w13202_,
		_w26623_
	);
	LUT2 #(
		.INIT('h8)
	) name16112 (
		\wishbone_bd_ram_mem1_reg[106][8]/P0001 ,
		_w12713_,
		_w26624_
	);
	LUT2 #(
		.INIT('h8)
	) name16113 (
		\wishbone_bd_ram_mem1_reg[238][8]/P0001 ,
		_w13160_,
		_w26625_
	);
	LUT2 #(
		.INIT('h8)
	) name16114 (
		\wishbone_bd_ram_mem1_reg[128][8]/P0001 ,
		_w12793_,
		_w26626_
	);
	LUT2 #(
		.INIT('h8)
	) name16115 (
		\wishbone_bd_ram_mem1_reg[214][8]/P0001 ,
		_w12984_,
		_w26627_
	);
	LUT2 #(
		.INIT('h8)
	) name16116 (
		\wishbone_bd_ram_mem1_reg[172][8]/P0001 ,
		_w12944_,
		_w26628_
	);
	LUT2 #(
		.INIT('h8)
	) name16117 (
		\wishbone_bd_ram_mem1_reg[207][8]/P0001 ,
		_w13180_,
		_w26629_
	);
	LUT2 #(
		.INIT('h8)
	) name16118 (
		\wishbone_bd_ram_mem1_reg[90][8]/P0001 ,
		_w12978_,
		_w26630_
	);
	LUT2 #(
		.INIT('h8)
	) name16119 (
		\wishbone_bd_ram_mem1_reg[150][8]/P0001 ,
		_w13136_,
		_w26631_
	);
	LUT2 #(
		.INIT('h8)
	) name16120 (
		\wishbone_bd_ram_mem1_reg[147][8]/P0001 ,
		_w13146_,
		_w26632_
	);
	LUT2 #(
		.INIT('h8)
	) name16121 (
		\wishbone_bd_ram_mem1_reg[225][8]/P0001 ,
		_w13092_,
		_w26633_
	);
	LUT2 #(
		.INIT('h8)
	) name16122 (
		\wishbone_bd_ram_mem1_reg[7][8]/P0001 ,
		_w12728_,
		_w26634_
	);
	LUT2 #(
		.INIT('h8)
	) name16123 (
		\wishbone_bd_ram_mem1_reg[9][8]/P0001 ,
		_w12808_,
		_w26635_
	);
	LUT2 #(
		.INIT('h8)
	) name16124 (
		\wishbone_bd_ram_mem1_reg[242][8]/P0001 ,
		_w12932_,
		_w26636_
	);
	LUT2 #(
		.INIT('h8)
	) name16125 (
		\wishbone_bd_ram_mem1_reg[61][8]/P0001 ,
		_w12725_,
		_w26637_
	);
	LUT2 #(
		.INIT('h8)
	) name16126 (
		\wishbone_bd_ram_mem1_reg[93][8]/P0001 ,
		_w13016_,
		_w26638_
	);
	LUT2 #(
		.INIT('h8)
	) name16127 (
		\wishbone_bd_ram_mem1_reg[83][8]/P0001 ,
		_w12916_,
		_w26639_
	);
	LUT2 #(
		.INIT('h8)
	) name16128 (
		\wishbone_bd_ram_mem1_reg[41][8]/P0001 ,
		_w13052_,
		_w26640_
	);
	LUT2 #(
		.INIT('h8)
	) name16129 (
		\wishbone_bd_ram_mem1_reg[52][8]/P0001 ,
		_w13082_,
		_w26641_
	);
	LUT2 #(
		.INIT('h8)
	) name16130 (
		\wishbone_bd_ram_mem1_reg[105][8]/P0001 ,
		_w12751_,
		_w26642_
	);
	LUT2 #(
		.INIT('h8)
	) name16131 (
		\wishbone_bd_ram_mem1_reg[79][8]/P0001 ,
		_w13212_,
		_w26643_
	);
	LUT2 #(
		.INIT('h8)
	) name16132 (
		\wishbone_bd_ram_mem1_reg[224][8]/P0001 ,
		_w12902_,
		_w26644_
	);
	LUT2 #(
		.INIT('h1)
	) name16133 (
		_w26389_,
		_w26390_,
		_w26645_
	);
	LUT2 #(
		.INIT('h1)
	) name16134 (
		_w26391_,
		_w26392_,
		_w26646_
	);
	LUT2 #(
		.INIT('h1)
	) name16135 (
		_w26393_,
		_w26394_,
		_w26647_
	);
	LUT2 #(
		.INIT('h1)
	) name16136 (
		_w26395_,
		_w26396_,
		_w26648_
	);
	LUT2 #(
		.INIT('h1)
	) name16137 (
		_w26397_,
		_w26398_,
		_w26649_
	);
	LUT2 #(
		.INIT('h1)
	) name16138 (
		_w26399_,
		_w26400_,
		_w26650_
	);
	LUT2 #(
		.INIT('h1)
	) name16139 (
		_w26401_,
		_w26402_,
		_w26651_
	);
	LUT2 #(
		.INIT('h1)
	) name16140 (
		_w26403_,
		_w26404_,
		_w26652_
	);
	LUT2 #(
		.INIT('h1)
	) name16141 (
		_w26405_,
		_w26406_,
		_w26653_
	);
	LUT2 #(
		.INIT('h1)
	) name16142 (
		_w26407_,
		_w26408_,
		_w26654_
	);
	LUT2 #(
		.INIT('h1)
	) name16143 (
		_w26409_,
		_w26410_,
		_w26655_
	);
	LUT2 #(
		.INIT('h1)
	) name16144 (
		_w26411_,
		_w26412_,
		_w26656_
	);
	LUT2 #(
		.INIT('h1)
	) name16145 (
		_w26413_,
		_w26414_,
		_w26657_
	);
	LUT2 #(
		.INIT('h1)
	) name16146 (
		_w26415_,
		_w26416_,
		_w26658_
	);
	LUT2 #(
		.INIT('h1)
	) name16147 (
		_w26417_,
		_w26418_,
		_w26659_
	);
	LUT2 #(
		.INIT('h1)
	) name16148 (
		_w26419_,
		_w26420_,
		_w26660_
	);
	LUT2 #(
		.INIT('h1)
	) name16149 (
		_w26421_,
		_w26422_,
		_w26661_
	);
	LUT2 #(
		.INIT('h1)
	) name16150 (
		_w26423_,
		_w26424_,
		_w26662_
	);
	LUT2 #(
		.INIT('h1)
	) name16151 (
		_w26425_,
		_w26426_,
		_w26663_
	);
	LUT2 #(
		.INIT('h1)
	) name16152 (
		_w26427_,
		_w26428_,
		_w26664_
	);
	LUT2 #(
		.INIT('h1)
	) name16153 (
		_w26429_,
		_w26430_,
		_w26665_
	);
	LUT2 #(
		.INIT('h1)
	) name16154 (
		_w26431_,
		_w26432_,
		_w26666_
	);
	LUT2 #(
		.INIT('h1)
	) name16155 (
		_w26433_,
		_w26434_,
		_w26667_
	);
	LUT2 #(
		.INIT('h1)
	) name16156 (
		_w26435_,
		_w26436_,
		_w26668_
	);
	LUT2 #(
		.INIT('h1)
	) name16157 (
		_w26437_,
		_w26438_,
		_w26669_
	);
	LUT2 #(
		.INIT('h1)
	) name16158 (
		_w26439_,
		_w26440_,
		_w26670_
	);
	LUT2 #(
		.INIT('h1)
	) name16159 (
		_w26441_,
		_w26442_,
		_w26671_
	);
	LUT2 #(
		.INIT('h1)
	) name16160 (
		_w26443_,
		_w26444_,
		_w26672_
	);
	LUT2 #(
		.INIT('h1)
	) name16161 (
		_w26445_,
		_w26446_,
		_w26673_
	);
	LUT2 #(
		.INIT('h1)
	) name16162 (
		_w26447_,
		_w26448_,
		_w26674_
	);
	LUT2 #(
		.INIT('h1)
	) name16163 (
		_w26449_,
		_w26450_,
		_w26675_
	);
	LUT2 #(
		.INIT('h1)
	) name16164 (
		_w26451_,
		_w26452_,
		_w26676_
	);
	LUT2 #(
		.INIT('h1)
	) name16165 (
		_w26453_,
		_w26454_,
		_w26677_
	);
	LUT2 #(
		.INIT('h1)
	) name16166 (
		_w26455_,
		_w26456_,
		_w26678_
	);
	LUT2 #(
		.INIT('h1)
	) name16167 (
		_w26457_,
		_w26458_,
		_w26679_
	);
	LUT2 #(
		.INIT('h1)
	) name16168 (
		_w26459_,
		_w26460_,
		_w26680_
	);
	LUT2 #(
		.INIT('h1)
	) name16169 (
		_w26461_,
		_w26462_,
		_w26681_
	);
	LUT2 #(
		.INIT('h1)
	) name16170 (
		_w26463_,
		_w26464_,
		_w26682_
	);
	LUT2 #(
		.INIT('h1)
	) name16171 (
		_w26465_,
		_w26466_,
		_w26683_
	);
	LUT2 #(
		.INIT('h1)
	) name16172 (
		_w26467_,
		_w26468_,
		_w26684_
	);
	LUT2 #(
		.INIT('h1)
	) name16173 (
		_w26469_,
		_w26470_,
		_w26685_
	);
	LUT2 #(
		.INIT('h1)
	) name16174 (
		_w26471_,
		_w26472_,
		_w26686_
	);
	LUT2 #(
		.INIT('h1)
	) name16175 (
		_w26473_,
		_w26474_,
		_w26687_
	);
	LUT2 #(
		.INIT('h1)
	) name16176 (
		_w26475_,
		_w26476_,
		_w26688_
	);
	LUT2 #(
		.INIT('h1)
	) name16177 (
		_w26477_,
		_w26478_,
		_w26689_
	);
	LUT2 #(
		.INIT('h1)
	) name16178 (
		_w26479_,
		_w26480_,
		_w26690_
	);
	LUT2 #(
		.INIT('h1)
	) name16179 (
		_w26481_,
		_w26482_,
		_w26691_
	);
	LUT2 #(
		.INIT('h1)
	) name16180 (
		_w26483_,
		_w26484_,
		_w26692_
	);
	LUT2 #(
		.INIT('h1)
	) name16181 (
		_w26485_,
		_w26486_,
		_w26693_
	);
	LUT2 #(
		.INIT('h1)
	) name16182 (
		_w26487_,
		_w26488_,
		_w26694_
	);
	LUT2 #(
		.INIT('h1)
	) name16183 (
		_w26489_,
		_w26490_,
		_w26695_
	);
	LUT2 #(
		.INIT('h1)
	) name16184 (
		_w26491_,
		_w26492_,
		_w26696_
	);
	LUT2 #(
		.INIT('h1)
	) name16185 (
		_w26493_,
		_w26494_,
		_w26697_
	);
	LUT2 #(
		.INIT('h1)
	) name16186 (
		_w26495_,
		_w26496_,
		_w26698_
	);
	LUT2 #(
		.INIT('h1)
	) name16187 (
		_w26497_,
		_w26498_,
		_w26699_
	);
	LUT2 #(
		.INIT('h1)
	) name16188 (
		_w26499_,
		_w26500_,
		_w26700_
	);
	LUT2 #(
		.INIT('h1)
	) name16189 (
		_w26501_,
		_w26502_,
		_w26701_
	);
	LUT2 #(
		.INIT('h1)
	) name16190 (
		_w26503_,
		_w26504_,
		_w26702_
	);
	LUT2 #(
		.INIT('h1)
	) name16191 (
		_w26505_,
		_w26506_,
		_w26703_
	);
	LUT2 #(
		.INIT('h1)
	) name16192 (
		_w26507_,
		_w26508_,
		_w26704_
	);
	LUT2 #(
		.INIT('h1)
	) name16193 (
		_w26509_,
		_w26510_,
		_w26705_
	);
	LUT2 #(
		.INIT('h1)
	) name16194 (
		_w26511_,
		_w26512_,
		_w26706_
	);
	LUT2 #(
		.INIT('h1)
	) name16195 (
		_w26513_,
		_w26514_,
		_w26707_
	);
	LUT2 #(
		.INIT('h1)
	) name16196 (
		_w26515_,
		_w26516_,
		_w26708_
	);
	LUT2 #(
		.INIT('h1)
	) name16197 (
		_w26517_,
		_w26518_,
		_w26709_
	);
	LUT2 #(
		.INIT('h1)
	) name16198 (
		_w26519_,
		_w26520_,
		_w26710_
	);
	LUT2 #(
		.INIT('h1)
	) name16199 (
		_w26521_,
		_w26522_,
		_w26711_
	);
	LUT2 #(
		.INIT('h1)
	) name16200 (
		_w26523_,
		_w26524_,
		_w26712_
	);
	LUT2 #(
		.INIT('h1)
	) name16201 (
		_w26525_,
		_w26526_,
		_w26713_
	);
	LUT2 #(
		.INIT('h1)
	) name16202 (
		_w26527_,
		_w26528_,
		_w26714_
	);
	LUT2 #(
		.INIT('h1)
	) name16203 (
		_w26529_,
		_w26530_,
		_w26715_
	);
	LUT2 #(
		.INIT('h1)
	) name16204 (
		_w26531_,
		_w26532_,
		_w26716_
	);
	LUT2 #(
		.INIT('h1)
	) name16205 (
		_w26533_,
		_w26534_,
		_w26717_
	);
	LUT2 #(
		.INIT('h1)
	) name16206 (
		_w26535_,
		_w26536_,
		_w26718_
	);
	LUT2 #(
		.INIT('h1)
	) name16207 (
		_w26537_,
		_w26538_,
		_w26719_
	);
	LUT2 #(
		.INIT('h1)
	) name16208 (
		_w26539_,
		_w26540_,
		_w26720_
	);
	LUT2 #(
		.INIT('h1)
	) name16209 (
		_w26541_,
		_w26542_,
		_w26721_
	);
	LUT2 #(
		.INIT('h1)
	) name16210 (
		_w26543_,
		_w26544_,
		_w26722_
	);
	LUT2 #(
		.INIT('h1)
	) name16211 (
		_w26545_,
		_w26546_,
		_w26723_
	);
	LUT2 #(
		.INIT('h1)
	) name16212 (
		_w26547_,
		_w26548_,
		_w26724_
	);
	LUT2 #(
		.INIT('h1)
	) name16213 (
		_w26549_,
		_w26550_,
		_w26725_
	);
	LUT2 #(
		.INIT('h1)
	) name16214 (
		_w26551_,
		_w26552_,
		_w26726_
	);
	LUT2 #(
		.INIT('h1)
	) name16215 (
		_w26553_,
		_w26554_,
		_w26727_
	);
	LUT2 #(
		.INIT('h1)
	) name16216 (
		_w26555_,
		_w26556_,
		_w26728_
	);
	LUT2 #(
		.INIT('h1)
	) name16217 (
		_w26557_,
		_w26558_,
		_w26729_
	);
	LUT2 #(
		.INIT('h1)
	) name16218 (
		_w26559_,
		_w26560_,
		_w26730_
	);
	LUT2 #(
		.INIT('h1)
	) name16219 (
		_w26561_,
		_w26562_,
		_w26731_
	);
	LUT2 #(
		.INIT('h1)
	) name16220 (
		_w26563_,
		_w26564_,
		_w26732_
	);
	LUT2 #(
		.INIT('h1)
	) name16221 (
		_w26565_,
		_w26566_,
		_w26733_
	);
	LUT2 #(
		.INIT('h1)
	) name16222 (
		_w26567_,
		_w26568_,
		_w26734_
	);
	LUT2 #(
		.INIT('h1)
	) name16223 (
		_w26569_,
		_w26570_,
		_w26735_
	);
	LUT2 #(
		.INIT('h1)
	) name16224 (
		_w26571_,
		_w26572_,
		_w26736_
	);
	LUT2 #(
		.INIT('h1)
	) name16225 (
		_w26573_,
		_w26574_,
		_w26737_
	);
	LUT2 #(
		.INIT('h1)
	) name16226 (
		_w26575_,
		_w26576_,
		_w26738_
	);
	LUT2 #(
		.INIT('h1)
	) name16227 (
		_w26577_,
		_w26578_,
		_w26739_
	);
	LUT2 #(
		.INIT('h1)
	) name16228 (
		_w26579_,
		_w26580_,
		_w26740_
	);
	LUT2 #(
		.INIT('h1)
	) name16229 (
		_w26581_,
		_w26582_,
		_w26741_
	);
	LUT2 #(
		.INIT('h1)
	) name16230 (
		_w26583_,
		_w26584_,
		_w26742_
	);
	LUT2 #(
		.INIT('h1)
	) name16231 (
		_w26585_,
		_w26586_,
		_w26743_
	);
	LUT2 #(
		.INIT('h1)
	) name16232 (
		_w26587_,
		_w26588_,
		_w26744_
	);
	LUT2 #(
		.INIT('h1)
	) name16233 (
		_w26589_,
		_w26590_,
		_w26745_
	);
	LUT2 #(
		.INIT('h1)
	) name16234 (
		_w26591_,
		_w26592_,
		_w26746_
	);
	LUT2 #(
		.INIT('h1)
	) name16235 (
		_w26593_,
		_w26594_,
		_w26747_
	);
	LUT2 #(
		.INIT('h1)
	) name16236 (
		_w26595_,
		_w26596_,
		_w26748_
	);
	LUT2 #(
		.INIT('h1)
	) name16237 (
		_w26597_,
		_w26598_,
		_w26749_
	);
	LUT2 #(
		.INIT('h1)
	) name16238 (
		_w26599_,
		_w26600_,
		_w26750_
	);
	LUT2 #(
		.INIT('h1)
	) name16239 (
		_w26601_,
		_w26602_,
		_w26751_
	);
	LUT2 #(
		.INIT('h1)
	) name16240 (
		_w26603_,
		_w26604_,
		_w26752_
	);
	LUT2 #(
		.INIT('h1)
	) name16241 (
		_w26605_,
		_w26606_,
		_w26753_
	);
	LUT2 #(
		.INIT('h1)
	) name16242 (
		_w26607_,
		_w26608_,
		_w26754_
	);
	LUT2 #(
		.INIT('h1)
	) name16243 (
		_w26609_,
		_w26610_,
		_w26755_
	);
	LUT2 #(
		.INIT('h1)
	) name16244 (
		_w26611_,
		_w26612_,
		_w26756_
	);
	LUT2 #(
		.INIT('h1)
	) name16245 (
		_w26613_,
		_w26614_,
		_w26757_
	);
	LUT2 #(
		.INIT('h1)
	) name16246 (
		_w26615_,
		_w26616_,
		_w26758_
	);
	LUT2 #(
		.INIT('h1)
	) name16247 (
		_w26617_,
		_w26618_,
		_w26759_
	);
	LUT2 #(
		.INIT('h1)
	) name16248 (
		_w26619_,
		_w26620_,
		_w26760_
	);
	LUT2 #(
		.INIT('h1)
	) name16249 (
		_w26621_,
		_w26622_,
		_w26761_
	);
	LUT2 #(
		.INIT('h1)
	) name16250 (
		_w26623_,
		_w26624_,
		_w26762_
	);
	LUT2 #(
		.INIT('h1)
	) name16251 (
		_w26625_,
		_w26626_,
		_w26763_
	);
	LUT2 #(
		.INIT('h1)
	) name16252 (
		_w26627_,
		_w26628_,
		_w26764_
	);
	LUT2 #(
		.INIT('h1)
	) name16253 (
		_w26629_,
		_w26630_,
		_w26765_
	);
	LUT2 #(
		.INIT('h1)
	) name16254 (
		_w26631_,
		_w26632_,
		_w26766_
	);
	LUT2 #(
		.INIT('h1)
	) name16255 (
		_w26633_,
		_w26634_,
		_w26767_
	);
	LUT2 #(
		.INIT('h1)
	) name16256 (
		_w26635_,
		_w26636_,
		_w26768_
	);
	LUT2 #(
		.INIT('h1)
	) name16257 (
		_w26637_,
		_w26638_,
		_w26769_
	);
	LUT2 #(
		.INIT('h1)
	) name16258 (
		_w26639_,
		_w26640_,
		_w26770_
	);
	LUT2 #(
		.INIT('h1)
	) name16259 (
		_w26641_,
		_w26642_,
		_w26771_
	);
	LUT2 #(
		.INIT('h1)
	) name16260 (
		_w26643_,
		_w26644_,
		_w26772_
	);
	LUT2 #(
		.INIT('h8)
	) name16261 (
		_w26771_,
		_w26772_,
		_w26773_
	);
	LUT2 #(
		.INIT('h8)
	) name16262 (
		_w26769_,
		_w26770_,
		_w26774_
	);
	LUT2 #(
		.INIT('h8)
	) name16263 (
		_w26767_,
		_w26768_,
		_w26775_
	);
	LUT2 #(
		.INIT('h8)
	) name16264 (
		_w26765_,
		_w26766_,
		_w26776_
	);
	LUT2 #(
		.INIT('h8)
	) name16265 (
		_w26763_,
		_w26764_,
		_w26777_
	);
	LUT2 #(
		.INIT('h8)
	) name16266 (
		_w26761_,
		_w26762_,
		_w26778_
	);
	LUT2 #(
		.INIT('h8)
	) name16267 (
		_w26759_,
		_w26760_,
		_w26779_
	);
	LUT2 #(
		.INIT('h8)
	) name16268 (
		_w26757_,
		_w26758_,
		_w26780_
	);
	LUT2 #(
		.INIT('h8)
	) name16269 (
		_w26755_,
		_w26756_,
		_w26781_
	);
	LUT2 #(
		.INIT('h8)
	) name16270 (
		_w26753_,
		_w26754_,
		_w26782_
	);
	LUT2 #(
		.INIT('h8)
	) name16271 (
		_w26751_,
		_w26752_,
		_w26783_
	);
	LUT2 #(
		.INIT('h8)
	) name16272 (
		_w26749_,
		_w26750_,
		_w26784_
	);
	LUT2 #(
		.INIT('h8)
	) name16273 (
		_w26747_,
		_w26748_,
		_w26785_
	);
	LUT2 #(
		.INIT('h8)
	) name16274 (
		_w26745_,
		_w26746_,
		_w26786_
	);
	LUT2 #(
		.INIT('h8)
	) name16275 (
		_w26743_,
		_w26744_,
		_w26787_
	);
	LUT2 #(
		.INIT('h8)
	) name16276 (
		_w26741_,
		_w26742_,
		_w26788_
	);
	LUT2 #(
		.INIT('h8)
	) name16277 (
		_w26739_,
		_w26740_,
		_w26789_
	);
	LUT2 #(
		.INIT('h8)
	) name16278 (
		_w26737_,
		_w26738_,
		_w26790_
	);
	LUT2 #(
		.INIT('h8)
	) name16279 (
		_w26735_,
		_w26736_,
		_w26791_
	);
	LUT2 #(
		.INIT('h8)
	) name16280 (
		_w26733_,
		_w26734_,
		_w26792_
	);
	LUT2 #(
		.INIT('h8)
	) name16281 (
		_w26731_,
		_w26732_,
		_w26793_
	);
	LUT2 #(
		.INIT('h8)
	) name16282 (
		_w26729_,
		_w26730_,
		_w26794_
	);
	LUT2 #(
		.INIT('h8)
	) name16283 (
		_w26727_,
		_w26728_,
		_w26795_
	);
	LUT2 #(
		.INIT('h8)
	) name16284 (
		_w26725_,
		_w26726_,
		_w26796_
	);
	LUT2 #(
		.INIT('h8)
	) name16285 (
		_w26723_,
		_w26724_,
		_w26797_
	);
	LUT2 #(
		.INIT('h8)
	) name16286 (
		_w26721_,
		_w26722_,
		_w26798_
	);
	LUT2 #(
		.INIT('h8)
	) name16287 (
		_w26719_,
		_w26720_,
		_w26799_
	);
	LUT2 #(
		.INIT('h8)
	) name16288 (
		_w26717_,
		_w26718_,
		_w26800_
	);
	LUT2 #(
		.INIT('h8)
	) name16289 (
		_w26715_,
		_w26716_,
		_w26801_
	);
	LUT2 #(
		.INIT('h8)
	) name16290 (
		_w26713_,
		_w26714_,
		_w26802_
	);
	LUT2 #(
		.INIT('h8)
	) name16291 (
		_w26711_,
		_w26712_,
		_w26803_
	);
	LUT2 #(
		.INIT('h8)
	) name16292 (
		_w26709_,
		_w26710_,
		_w26804_
	);
	LUT2 #(
		.INIT('h8)
	) name16293 (
		_w26707_,
		_w26708_,
		_w26805_
	);
	LUT2 #(
		.INIT('h8)
	) name16294 (
		_w26705_,
		_w26706_,
		_w26806_
	);
	LUT2 #(
		.INIT('h8)
	) name16295 (
		_w26703_,
		_w26704_,
		_w26807_
	);
	LUT2 #(
		.INIT('h8)
	) name16296 (
		_w26701_,
		_w26702_,
		_w26808_
	);
	LUT2 #(
		.INIT('h8)
	) name16297 (
		_w26699_,
		_w26700_,
		_w26809_
	);
	LUT2 #(
		.INIT('h8)
	) name16298 (
		_w26697_,
		_w26698_,
		_w26810_
	);
	LUT2 #(
		.INIT('h8)
	) name16299 (
		_w26695_,
		_w26696_,
		_w26811_
	);
	LUT2 #(
		.INIT('h8)
	) name16300 (
		_w26693_,
		_w26694_,
		_w26812_
	);
	LUT2 #(
		.INIT('h8)
	) name16301 (
		_w26691_,
		_w26692_,
		_w26813_
	);
	LUT2 #(
		.INIT('h8)
	) name16302 (
		_w26689_,
		_w26690_,
		_w26814_
	);
	LUT2 #(
		.INIT('h8)
	) name16303 (
		_w26687_,
		_w26688_,
		_w26815_
	);
	LUT2 #(
		.INIT('h8)
	) name16304 (
		_w26685_,
		_w26686_,
		_w26816_
	);
	LUT2 #(
		.INIT('h8)
	) name16305 (
		_w26683_,
		_w26684_,
		_w26817_
	);
	LUT2 #(
		.INIT('h8)
	) name16306 (
		_w26681_,
		_w26682_,
		_w26818_
	);
	LUT2 #(
		.INIT('h8)
	) name16307 (
		_w26679_,
		_w26680_,
		_w26819_
	);
	LUT2 #(
		.INIT('h8)
	) name16308 (
		_w26677_,
		_w26678_,
		_w26820_
	);
	LUT2 #(
		.INIT('h8)
	) name16309 (
		_w26675_,
		_w26676_,
		_w26821_
	);
	LUT2 #(
		.INIT('h8)
	) name16310 (
		_w26673_,
		_w26674_,
		_w26822_
	);
	LUT2 #(
		.INIT('h8)
	) name16311 (
		_w26671_,
		_w26672_,
		_w26823_
	);
	LUT2 #(
		.INIT('h8)
	) name16312 (
		_w26669_,
		_w26670_,
		_w26824_
	);
	LUT2 #(
		.INIT('h8)
	) name16313 (
		_w26667_,
		_w26668_,
		_w26825_
	);
	LUT2 #(
		.INIT('h8)
	) name16314 (
		_w26665_,
		_w26666_,
		_w26826_
	);
	LUT2 #(
		.INIT('h8)
	) name16315 (
		_w26663_,
		_w26664_,
		_w26827_
	);
	LUT2 #(
		.INIT('h8)
	) name16316 (
		_w26661_,
		_w26662_,
		_w26828_
	);
	LUT2 #(
		.INIT('h8)
	) name16317 (
		_w26659_,
		_w26660_,
		_w26829_
	);
	LUT2 #(
		.INIT('h8)
	) name16318 (
		_w26657_,
		_w26658_,
		_w26830_
	);
	LUT2 #(
		.INIT('h8)
	) name16319 (
		_w26655_,
		_w26656_,
		_w26831_
	);
	LUT2 #(
		.INIT('h8)
	) name16320 (
		_w26653_,
		_w26654_,
		_w26832_
	);
	LUT2 #(
		.INIT('h8)
	) name16321 (
		_w26651_,
		_w26652_,
		_w26833_
	);
	LUT2 #(
		.INIT('h8)
	) name16322 (
		_w26649_,
		_w26650_,
		_w26834_
	);
	LUT2 #(
		.INIT('h8)
	) name16323 (
		_w26647_,
		_w26648_,
		_w26835_
	);
	LUT2 #(
		.INIT('h8)
	) name16324 (
		_w26645_,
		_w26646_,
		_w26836_
	);
	LUT2 #(
		.INIT('h8)
	) name16325 (
		_w26835_,
		_w26836_,
		_w26837_
	);
	LUT2 #(
		.INIT('h8)
	) name16326 (
		_w26833_,
		_w26834_,
		_w26838_
	);
	LUT2 #(
		.INIT('h8)
	) name16327 (
		_w26831_,
		_w26832_,
		_w26839_
	);
	LUT2 #(
		.INIT('h8)
	) name16328 (
		_w26829_,
		_w26830_,
		_w26840_
	);
	LUT2 #(
		.INIT('h8)
	) name16329 (
		_w26827_,
		_w26828_,
		_w26841_
	);
	LUT2 #(
		.INIT('h8)
	) name16330 (
		_w26825_,
		_w26826_,
		_w26842_
	);
	LUT2 #(
		.INIT('h8)
	) name16331 (
		_w26823_,
		_w26824_,
		_w26843_
	);
	LUT2 #(
		.INIT('h8)
	) name16332 (
		_w26821_,
		_w26822_,
		_w26844_
	);
	LUT2 #(
		.INIT('h8)
	) name16333 (
		_w26819_,
		_w26820_,
		_w26845_
	);
	LUT2 #(
		.INIT('h8)
	) name16334 (
		_w26817_,
		_w26818_,
		_w26846_
	);
	LUT2 #(
		.INIT('h8)
	) name16335 (
		_w26815_,
		_w26816_,
		_w26847_
	);
	LUT2 #(
		.INIT('h8)
	) name16336 (
		_w26813_,
		_w26814_,
		_w26848_
	);
	LUT2 #(
		.INIT('h8)
	) name16337 (
		_w26811_,
		_w26812_,
		_w26849_
	);
	LUT2 #(
		.INIT('h8)
	) name16338 (
		_w26809_,
		_w26810_,
		_w26850_
	);
	LUT2 #(
		.INIT('h8)
	) name16339 (
		_w26807_,
		_w26808_,
		_w26851_
	);
	LUT2 #(
		.INIT('h8)
	) name16340 (
		_w26805_,
		_w26806_,
		_w26852_
	);
	LUT2 #(
		.INIT('h8)
	) name16341 (
		_w26803_,
		_w26804_,
		_w26853_
	);
	LUT2 #(
		.INIT('h8)
	) name16342 (
		_w26801_,
		_w26802_,
		_w26854_
	);
	LUT2 #(
		.INIT('h8)
	) name16343 (
		_w26799_,
		_w26800_,
		_w26855_
	);
	LUT2 #(
		.INIT('h8)
	) name16344 (
		_w26797_,
		_w26798_,
		_w26856_
	);
	LUT2 #(
		.INIT('h8)
	) name16345 (
		_w26795_,
		_w26796_,
		_w26857_
	);
	LUT2 #(
		.INIT('h8)
	) name16346 (
		_w26793_,
		_w26794_,
		_w26858_
	);
	LUT2 #(
		.INIT('h8)
	) name16347 (
		_w26791_,
		_w26792_,
		_w26859_
	);
	LUT2 #(
		.INIT('h8)
	) name16348 (
		_w26789_,
		_w26790_,
		_w26860_
	);
	LUT2 #(
		.INIT('h8)
	) name16349 (
		_w26787_,
		_w26788_,
		_w26861_
	);
	LUT2 #(
		.INIT('h8)
	) name16350 (
		_w26785_,
		_w26786_,
		_w26862_
	);
	LUT2 #(
		.INIT('h8)
	) name16351 (
		_w26783_,
		_w26784_,
		_w26863_
	);
	LUT2 #(
		.INIT('h8)
	) name16352 (
		_w26781_,
		_w26782_,
		_w26864_
	);
	LUT2 #(
		.INIT('h8)
	) name16353 (
		_w26779_,
		_w26780_,
		_w26865_
	);
	LUT2 #(
		.INIT('h8)
	) name16354 (
		_w26777_,
		_w26778_,
		_w26866_
	);
	LUT2 #(
		.INIT('h8)
	) name16355 (
		_w26775_,
		_w26776_,
		_w26867_
	);
	LUT2 #(
		.INIT('h8)
	) name16356 (
		_w26773_,
		_w26774_,
		_w26868_
	);
	LUT2 #(
		.INIT('h8)
	) name16357 (
		_w26867_,
		_w26868_,
		_w26869_
	);
	LUT2 #(
		.INIT('h8)
	) name16358 (
		_w26865_,
		_w26866_,
		_w26870_
	);
	LUT2 #(
		.INIT('h8)
	) name16359 (
		_w26863_,
		_w26864_,
		_w26871_
	);
	LUT2 #(
		.INIT('h8)
	) name16360 (
		_w26861_,
		_w26862_,
		_w26872_
	);
	LUT2 #(
		.INIT('h8)
	) name16361 (
		_w26859_,
		_w26860_,
		_w26873_
	);
	LUT2 #(
		.INIT('h8)
	) name16362 (
		_w26857_,
		_w26858_,
		_w26874_
	);
	LUT2 #(
		.INIT('h8)
	) name16363 (
		_w26855_,
		_w26856_,
		_w26875_
	);
	LUT2 #(
		.INIT('h8)
	) name16364 (
		_w26853_,
		_w26854_,
		_w26876_
	);
	LUT2 #(
		.INIT('h8)
	) name16365 (
		_w26851_,
		_w26852_,
		_w26877_
	);
	LUT2 #(
		.INIT('h8)
	) name16366 (
		_w26849_,
		_w26850_,
		_w26878_
	);
	LUT2 #(
		.INIT('h8)
	) name16367 (
		_w26847_,
		_w26848_,
		_w26879_
	);
	LUT2 #(
		.INIT('h8)
	) name16368 (
		_w26845_,
		_w26846_,
		_w26880_
	);
	LUT2 #(
		.INIT('h8)
	) name16369 (
		_w26843_,
		_w26844_,
		_w26881_
	);
	LUT2 #(
		.INIT('h8)
	) name16370 (
		_w26841_,
		_w26842_,
		_w26882_
	);
	LUT2 #(
		.INIT('h8)
	) name16371 (
		_w26839_,
		_w26840_,
		_w26883_
	);
	LUT2 #(
		.INIT('h8)
	) name16372 (
		_w26837_,
		_w26838_,
		_w26884_
	);
	LUT2 #(
		.INIT('h8)
	) name16373 (
		_w26883_,
		_w26884_,
		_w26885_
	);
	LUT2 #(
		.INIT('h8)
	) name16374 (
		_w26881_,
		_w26882_,
		_w26886_
	);
	LUT2 #(
		.INIT('h8)
	) name16375 (
		_w26879_,
		_w26880_,
		_w26887_
	);
	LUT2 #(
		.INIT('h8)
	) name16376 (
		_w26877_,
		_w26878_,
		_w26888_
	);
	LUT2 #(
		.INIT('h8)
	) name16377 (
		_w26875_,
		_w26876_,
		_w26889_
	);
	LUT2 #(
		.INIT('h8)
	) name16378 (
		_w26873_,
		_w26874_,
		_w26890_
	);
	LUT2 #(
		.INIT('h8)
	) name16379 (
		_w26871_,
		_w26872_,
		_w26891_
	);
	LUT2 #(
		.INIT('h8)
	) name16380 (
		_w26869_,
		_w26870_,
		_w26892_
	);
	LUT2 #(
		.INIT('h8)
	) name16381 (
		_w26891_,
		_w26892_,
		_w26893_
	);
	LUT2 #(
		.INIT('h8)
	) name16382 (
		_w26889_,
		_w26890_,
		_w26894_
	);
	LUT2 #(
		.INIT('h8)
	) name16383 (
		_w26887_,
		_w26888_,
		_w26895_
	);
	LUT2 #(
		.INIT('h8)
	) name16384 (
		_w26885_,
		_w26886_,
		_w26896_
	);
	LUT2 #(
		.INIT('h8)
	) name16385 (
		_w26895_,
		_w26896_,
		_w26897_
	);
	LUT2 #(
		.INIT('h8)
	) name16386 (
		_w26893_,
		_w26894_,
		_w26898_
	);
	LUT2 #(
		.INIT('h8)
	) name16387 (
		_w26897_,
		_w26898_,
		_w26899_
	);
	LUT2 #(
		.INIT('h1)
	) name16388 (
		wb_rst_i_pad,
		_w26899_,
		_w26900_
	);
	LUT2 #(
		.INIT('h1)
	) name16389 (
		_w22944_,
		_w26900_,
		_w26901_
	);
	LUT2 #(
		.INIT('h8)
	) name16390 (
		\ethreg1_PACKETLEN_1_DataOut_reg[0]/NET0131 ,
		_w22966_,
		_w26902_
	);
	LUT2 #(
		.INIT('h8)
	) name16391 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 ,
		_w23522_,
		_w26903_
	);
	LUT2 #(
		.INIT('h8)
	) name16392 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		_w24726_,
		_w26904_
	);
	LUT2 #(
		.INIT('h8)
	) name16393 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		_w22959_,
		_w26905_
	);
	LUT2 #(
		.INIT('h8)
	) name16394 (
		\ethreg1_MODER_1_DataOut_reg[0]/NET0131 ,
		_w23519_,
		_w26906_
	);
	LUT2 #(
		.INIT('h8)
	) name16395 (
		\ethreg1_MIIRX_DATA_DataOut_reg[8]/NET0131 ,
		_w23507_,
		_w26907_
	);
	LUT2 #(
		.INIT('h8)
	) name16396 (
		\ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 ,
		_w22952_,
		_w26908_
	);
	LUT2 #(
		.INIT('h8)
	) name16397 (
		\ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 ,
		_w22956_,
		_w26909_
	);
	LUT2 #(
		.INIT('h8)
	) name16398 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		_w23501_,
		_w26910_
	);
	LUT2 #(
		.INIT('h8)
	) name16399 (
		\ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 ,
		_w23499_,
		_w26911_
	);
	LUT2 #(
		.INIT('h8)
	) name16400 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		_w23513_,
		_w26912_
	);
	LUT2 #(
		.INIT('h1)
	) name16401 (
		_w26903_,
		_w26904_,
		_w26913_
	);
	LUT2 #(
		.INIT('h1)
	) name16402 (
		_w26905_,
		_w26906_,
		_w26914_
	);
	LUT2 #(
		.INIT('h1)
	) name16403 (
		_w26907_,
		_w26908_,
		_w26915_
	);
	LUT2 #(
		.INIT('h1)
	) name16404 (
		_w26909_,
		_w26910_,
		_w26916_
	);
	LUT2 #(
		.INIT('h1)
	) name16405 (
		_w26911_,
		_w26912_,
		_w26917_
	);
	LUT2 #(
		.INIT('h8)
	) name16406 (
		_w26916_,
		_w26917_,
		_w26918_
	);
	LUT2 #(
		.INIT('h8)
	) name16407 (
		_w26914_,
		_w26915_,
		_w26919_
	);
	LUT2 #(
		.INIT('h8)
	) name16408 (
		_w22944_,
		_w26913_,
		_w26920_
	);
	LUT2 #(
		.INIT('h8)
	) name16409 (
		_w26919_,
		_w26920_,
		_w26921_
	);
	LUT2 #(
		.INIT('h4)
	) name16410 (
		_w26902_,
		_w26918_,
		_w26922_
	);
	LUT2 #(
		.INIT('h8)
	) name16411 (
		_w26921_,
		_w26922_,
		_w26923_
	);
	LUT2 #(
		.INIT('h1)
	) name16412 (
		_w26901_,
		_w26923_,
		_w26924_
	);
	LUT2 #(
		.INIT('h8)
	) name16413 (
		\wishbone_bd_ram_mem1_reg[9][9]/P0001 ,
		_w12808_,
		_w26925_
	);
	LUT2 #(
		.INIT('h8)
	) name16414 (
		\wishbone_bd_ram_mem1_reg[20][9]/P0001 ,
		_w13174_,
		_w26926_
	);
	LUT2 #(
		.INIT('h8)
	) name16415 (
		\wishbone_bd_ram_mem1_reg[30][9]/P0001 ,
		_w13104_,
		_w26927_
	);
	LUT2 #(
		.INIT('h8)
	) name16416 (
		\wishbone_bd_ram_mem1_reg[144][9]/P0001 ,
		_w12756_,
		_w26928_
	);
	LUT2 #(
		.INIT('h8)
	) name16417 (
		\wishbone_bd_ram_mem1_reg[84][9]/P0001 ,
		_w12934_,
		_w26929_
	);
	LUT2 #(
		.INIT('h8)
	) name16418 (
		\wishbone_bd_ram_mem1_reg[173][9]/P0001 ,
		_w12854_,
		_w26930_
	);
	LUT2 #(
		.INIT('h8)
	) name16419 (
		\wishbone_bd_ram_mem1_reg[119][9]/P0001 ,
		_w13048_,
		_w26931_
	);
	LUT2 #(
		.INIT('h8)
	) name16420 (
		\wishbone_bd_ram_mem1_reg[25][9]/P0001 ,
		_w13108_,
		_w26932_
	);
	LUT2 #(
		.INIT('h8)
	) name16421 (
		\wishbone_bd_ram_mem1_reg[231][9]/P0001 ,
		_w12856_,
		_w26933_
	);
	LUT2 #(
		.INIT('h8)
	) name16422 (
		\wishbone_bd_ram_mem1_reg[254][9]/P0001 ,
		_w12892_,
		_w26934_
	);
	LUT2 #(
		.INIT('h8)
	) name16423 (
		\wishbone_bd_ram_mem1_reg[205][9]/P0001 ,
		_w13068_,
		_w26935_
	);
	LUT2 #(
		.INIT('h8)
	) name16424 (
		\wishbone_bd_ram_mem1_reg[138][9]/P0001 ,
		_w12958_,
		_w26936_
	);
	LUT2 #(
		.INIT('h8)
	) name16425 (
		\wishbone_bd_ram_mem1_reg[13][9]/P0001 ,
		_w13178_,
		_w26937_
	);
	LUT2 #(
		.INIT('h8)
	) name16426 (
		\wishbone_bd_ram_mem1_reg[111][9]/P0001 ,
		_w12744_,
		_w26938_
	);
	LUT2 #(
		.INIT('h8)
	) name16427 (
		\wishbone_bd_ram_mem1_reg[118][9]/P0001 ,
		_w12830_,
		_w26939_
	);
	LUT2 #(
		.INIT('h8)
	) name16428 (
		\wishbone_bd_ram_mem1_reg[22][9]/P0001 ,
		_w13110_,
		_w26940_
	);
	LUT2 #(
		.INIT('h8)
	) name16429 (
		\wishbone_bd_ram_mem1_reg[68][9]/P0001 ,
		_w12946_,
		_w26941_
	);
	LUT2 #(
		.INIT('h8)
	) name16430 (
		\wishbone_bd_ram_mem1_reg[195][9]/P0001 ,
		_w13144_,
		_w26942_
	);
	LUT2 #(
		.INIT('h8)
	) name16431 (
		\wishbone_bd_ram_mem1_reg[166][9]/P0001 ,
		_w13040_,
		_w26943_
	);
	LUT2 #(
		.INIT('h8)
	) name16432 (
		\wishbone_bd_ram_mem1_reg[106][9]/P0001 ,
		_w12713_,
		_w26944_
	);
	LUT2 #(
		.INIT('h8)
	) name16433 (
		\wishbone_bd_ram_mem1_reg[73][9]/P0001 ,
		_w12918_,
		_w26945_
	);
	LUT2 #(
		.INIT('h8)
	) name16434 (
		\wishbone_bd_ram_mem1_reg[186][9]/P0001 ,
		_w12783_,
		_w26946_
	);
	LUT2 #(
		.INIT('h8)
	) name16435 (
		\wishbone_bd_ram_mem1_reg[236][9]/P0001 ,
		_w12731_,
		_w26947_
	);
	LUT2 #(
		.INIT('h8)
	) name16436 (
		\wishbone_bd_ram_mem1_reg[130][9]/P0001 ,
		_w12914_,
		_w26948_
	);
	LUT2 #(
		.INIT('h8)
	) name16437 (
		\wishbone_bd_ram_mem1_reg[193][9]/P0001 ,
		_w13056_,
		_w26949_
	);
	LUT2 #(
		.INIT('h8)
	) name16438 (
		\wishbone_bd_ram_mem1_reg[149][9]/P0001 ,
		_w12741_,
		_w26950_
	);
	LUT2 #(
		.INIT('h8)
	) name16439 (
		\wishbone_bd_ram_mem1_reg[151][9]/P0001 ,
		_w13142_,
		_w26951_
	);
	LUT2 #(
		.INIT('h8)
	) name16440 (
		\wishbone_bd_ram_mem1_reg[154][9]/P0001 ,
		_w12962_,
		_w26952_
	);
	LUT2 #(
		.INIT('h8)
	) name16441 (
		\wishbone_bd_ram_mem1_reg[139][9]/P0001 ,
		_w12814_,
		_w26953_
	);
	LUT2 #(
		.INIT('h8)
	) name16442 (
		\wishbone_bd_ram_mem1_reg[123][9]/P0001 ,
		_w13114_,
		_w26954_
	);
	LUT2 #(
		.INIT('h8)
	) name16443 (
		\wishbone_bd_ram_mem1_reg[196][9]/P0001 ,
		_w13090_,
		_w26955_
	);
	LUT2 #(
		.INIT('h8)
	) name16444 (
		\wishbone_bd_ram_mem1_reg[204][9]/P0001 ,
		_w13162_,
		_w26956_
	);
	LUT2 #(
		.INIT('h8)
	) name16445 (
		\wishbone_bd_ram_mem1_reg[168][9]/P0001 ,
		_w13208_,
		_w26957_
	);
	LUT2 #(
		.INIT('h8)
	) name16446 (
		\wishbone_bd_ram_mem1_reg[227][9]/P0001 ,
		_w12936_,
		_w26958_
	);
	LUT2 #(
		.INIT('h8)
	) name16447 (
		\wishbone_bd_ram_mem1_reg[55][9]/P0001 ,
		_w12785_,
		_w26959_
	);
	LUT2 #(
		.INIT('h8)
	) name16448 (
		\wishbone_bd_ram_mem1_reg[116][9]/P0001 ,
		_w12998_,
		_w26960_
	);
	LUT2 #(
		.INIT('h8)
	) name16449 (
		\wishbone_bd_ram_mem1_reg[61][9]/P0001 ,
		_w12725_,
		_w26961_
	);
	LUT2 #(
		.INIT('h8)
	) name16450 (
		\wishbone_bd_ram_mem1_reg[99][9]/P0001 ,
		_w13038_,
		_w26962_
	);
	LUT2 #(
		.INIT('h8)
	) name16451 (
		\wishbone_bd_ram_mem1_reg[228][9]/P0001 ,
		_w12765_,
		_w26963_
	);
	LUT2 #(
		.INIT('h8)
	) name16452 (
		\wishbone_bd_ram_mem1_reg[115][9]/P0001 ,
		_w13112_,
		_w26964_
	);
	LUT2 #(
		.INIT('h8)
	) name16453 (
		\wishbone_bd_ram_mem1_reg[255][9]/P0001 ,
		_w13072_,
		_w26965_
	);
	LUT2 #(
		.INIT('h8)
	) name16454 (
		\wishbone_bd_ram_mem1_reg[207][9]/P0001 ,
		_w13180_,
		_w26966_
	);
	LUT2 #(
		.INIT('h8)
	) name16455 (
		\wishbone_bd_ram_mem1_reg[121][9]/P0001 ,
		_w13078_,
		_w26967_
	);
	LUT2 #(
		.INIT('h8)
	) name16456 (
		\wishbone_bd_ram_mem1_reg[29][9]/P0001 ,
		_w12952_,
		_w26968_
	);
	LUT2 #(
		.INIT('h8)
	) name16457 (
		\wishbone_bd_ram_mem1_reg[49][9]/P0001 ,
		_w12994_,
		_w26969_
	);
	LUT2 #(
		.INIT('h8)
	) name16458 (
		\wishbone_bd_ram_mem1_reg[100][9]/P0001 ,
		_w12960_,
		_w26970_
	);
	LUT2 #(
		.INIT('h8)
	) name16459 (
		\wishbone_bd_ram_mem1_reg[80][9]/P0001 ,
		_w12689_,
		_w26971_
	);
	LUT2 #(
		.INIT('h8)
	) name16460 (
		\wishbone_bd_ram_mem1_reg[90][9]/P0001 ,
		_w12978_,
		_w26972_
	);
	LUT2 #(
		.INIT('h8)
	) name16461 (
		\wishbone_bd_ram_mem1_reg[220][9]/P0001 ,
		_w13066_,
		_w26973_
	);
	LUT2 #(
		.INIT('h8)
	) name16462 (
		\wishbone_bd_ram_mem1_reg[246][9]/P0001 ,
		_w13076_,
		_w26974_
	);
	LUT2 #(
		.INIT('h8)
	) name16463 (
		\wishbone_bd_ram_mem1_reg[2][9]/P0001 ,
		_w13088_,
		_w26975_
	);
	LUT2 #(
		.INIT('h8)
	) name16464 (
		\wishbone_bd_ram_mem1_reg[77][9]/P0001 ,
		_w12982_,
		_w26976_
	);
	LUT2 #(
		.INIT('h8)
	) name16465 (
		\wishbone_bd_ram_mem1_reg[165][9]/P0001 ,
		_w13044_,
		_w26977_
	);
	LUT2 #(
		.INIT('h8)
	) name16466 (
		\wishbone_bd_ram_mem1_reg[237][9]/P0001 ,
		_w12990_,
		_w26978_
	);
	LUT2 #(
		.INIT('h8)
	) name16467 (
		\wishbone_bd_ram_mem1_reg[146][9]/P0001 ,
		_w13060_,
		_w26979_
	);
	LUT2 #(
		.INIT('h8)
	) name16468 (
		\wishbone_bd_ram_mem1_reg[127][9]/P0001 ,
		_w13164_,
		_w26980_
	);
	LUT2 #(
		.INIT('h8)
	) name16469 (
		\wishbone_bd_ram_mem1_reg[180][9]/P0001 ,
		_w12791_,
		_w26981_
	);
	LUT2 #(
		.INIT('h8)
	) name16470 (
		\wishbone_bd_ram_mem1_reg[252][9]/P0001 ,
		_w13080_,
		_w26982_
	);
	LUT2 #(
		.INIT('h8)
	) name16471 (
		\wishbone_bd_ram_mem1_reg[167][9]/P0001 ,
		_w12986_,
		_w26983_
	);
	LUT2 #(
		.INIT('h8)
	) name16472 (
		\wishbone_bd_ram_mem1_reg[92][9]/P0001 ,
		_w13010_,
		_w26984_
	);
	LUT2 #(
		.INIT('h8)
	) name16473 (
		\wishbone_bd_ram_mem1_reg[213][9]/P0001 ,
		_w13002_,
		_w26985_
	);
	LUT2 #(
		.INIT('h8)
	) name16474 (
		\wishbone_bd_ram_mem1_reg[34][9]/P0001 ,
		_w12930_,
		_w26986_
	);
	LUT2 #(
		.INIT('h8)
	) name16475 (
		\wishbone_bd_ram_mem1_reg[184][9]/P0001 ,
		_w13062_,
		_w26987_
	);
	LUT2 #(
		.INIT('h8)
	) name16476 (
		\wishbone_bd_ram_mem1_reg[54][9]/P0001 ,
		_w12770_,
		_w26988_
	);
	LUT2 #(
		.INIT('h8)
	) name16477 (
		\wishbone_bd_ram_mem1_reg[194][9]/P0001 ,
		_w12772_,
		_w26989_
	);
	LUT2 #(
		.INIT('h8)
	) name16478 (
		\wishbone_bd_ram_mem1_reg[224][9]/P0001 ,
		_w12902_,
		_w26990_
	);
	LUT2 #(
		.INIT('h8)
	) name16479 (
		\wishbone_bd_ram_mem1_reg[185][9]/P0001 ,
		_w12940_,
		_w26991_
	);
	LUT2 #(
		.INIT('h8)
	) name16480 (
		\wishbone_bd_ram_mem1_reg[27][9]/P0001 ,
		_w12880_,
		_w26992_
	);
	LUT2 #(
		.INIT('h8)
	) name16481 (
		\wishbone_bd_ram_mem1_reg[107][9]/P0001 ,
		_w12749_,
		_w26993_
	);
	LUT2 #(
		.INIT('h8)
	) name16482 (
		\wishbone_bd_ram_mem1_reg[174][9]/P0001 ,
		_w12972_,
		_w26994_
	);
	LUT2 #(
		.INIT('h8)
	) name16483 (
		\wishbone_bd_ram_mem1_reg[1][9]/P0001 ,
		_w13014_,
		_w26995_
	);
	LUT2 #(
		.INIT('h8)
	) name16484 (
		\wishbone_bd_ram_mem1_reg[142][9]/P0001 ,
		_w12928_,
		_w26996_
	);
	LUT2 #(
		.INIT('h8)
	) name16485 (
		\wishbone_bd_ram_mem1_reg[52][9]/P0001 ,
		_w13082_,
		_w26997_
	);
	LUT2 #(
		.INIT('h8)
	) name16486 (
		\wishbone_bd_ram_mem1_reg[126][9]/P0001 ,
		_w13218_,
		_w26998_
	);
	LUT2 #(
		.INIT('h8)
	) name16487 (
		\wishbone_bd_ram_mem1_reg[171][9]/P0001 ,
		_w12910_,
		_w26999_
	);
	LUT2 #(
		.INIT('h8)
	) name16488 (
		\wishbone_bd_ram_mem1_reg[250][9]/P0001 ,
		_w13128_,
		_w27000_
	);
	LUT2 #(
		.INIT('h8)
	) name16489 (
		\wishbone_bd_ram_mem1_reg[95][9]/P0001 ,
		_w12844_,
		_w27001_
	);
	LUT2 #(
		.INIT('h8)
	) name16490 (
		\wishbone_bd_ram_mem1_reg[249][9]/P0001 ,
		_w12900_,
		_w27002_
	);
	LUT2 #(
		.INIT('h8)
	) name16491 (
		\wishbone_bd_ram_mem1_reg[201][9]/P0001 ,
		_w12822_,
		_w27003_
	);
	LUT2 #(
		.INIT('h8)
	) name16492 (
		\wishbone_bd_ram_mem1_reg[40][9]/P0001 ,
		_w13132_,
		_w27004_
	);
	LUT2 #(
		.INIT('h8)
	) name16493 (
		\wishbone_bd_ram_mem1_reg[48][9]/P0001 ,
		_w12970_,
		_w27005_
	);
	LUT2 #(
		.INIT('h8)
	) name16494 (
		\wishbone_bd_ram_mem1_reg[241][9]/P0001 ,
		_w13006_,
		_w27006_
	);
	LUT2 #(
		.INIT('h8)
	) name16495 (
		\wishbone_bd_ram_mem1_reg[57][9]/P0001 ,
		_w13116_,
		_w27007_
	);
	LUT2 #(
		.INIT('h8)
	) name16496 (
		\wishbone_bd_ram_mem1_reg[209][9]/P0001 ,
		_w13152_,
		_w27008_
	);
	LUT2 #(
		.INIT('h8)
	) name16497 (
		\wishbone_bd_ram_mem1_reg[39][9]/P0001 ,
		_w13018_,
		_w27009_
	);
	LUT2 #(
		.INIT('h8)
	) name16498 (
		\wishbone_bd_ram_mem1_reg[109][9]/P0001 ,
		_w12888_,
		_w27010_
	);
	LUT2 #(
		.INIT('h8)
	) name16499 (
		\wishbone_bd_ram_mem1_reg[82][9]/P0001 ,
		_w12942_,
		_w27011_
	);
	LUT2 #(
		.INIT('h8)
	) name16500 (
		\wishbone_bd_ram_mem1_reg[32][9]/P0001 ,
		_w13120_,
		_w27012_
	);
	LUT2 #(
		.INIT('h8)
	) name16501 (
		\wishbone_bd_ram_mem1_reg[7][9]/P0001 ,
		_w12728_,
		_w27013_
	);
	LUT2 #(
		.INIT('h8)
	) name16502 (
		\wishbone_bd_ram_mem1_reg[238][9]/P0001 ,
		_w13160_,
		_w27014_
	);
	LUT2 #(
		.INIT('h8)
	) name16503 (
		\wishbone_bd_ram_mem1_reg[36][9]/P0001 ,
		_w12800_,
		_w27015_
	);
	LUT2 #(
		.INIT('h8)
	) name16504 (
		\wishbone_bd_ram_mem1_reg[251][9]/P0001 ,
		_w13054_,
		_w27016_
	);
	LUT2 #(
		.INIT('h8)
	) name16505 (
		\wishbone_bd_ram_mem1_reg[178][9]/P0001 ,
		_w12886_,
		_w27017_
	);
	LUT2 #(
		.INIT('h8)
	) name16506 (
		\wishbone_bd_ram_mem1_reg[244][9]/P0001 ,
		_w12747_,
		_w27018_
	);
	LUT2 #(
		.INIT('h8)
	) name16507 (
		\wishbone_bd_ram_mem1_reg[160][9]/P0001 ,
		_w12872_,
		_w27019_
	);
	LUT2 #(
		.INIT('h8)
	) name16508 (
		\wishbone_bd_ram_mem1_reg[133][9]/P0001 ,
		_w12761_,
		_w27020_
	);
	LUT2 #(
		.INIT('h8)
	) name16509 (
		\wishbone_bd_ram_mem1_reg[42][9]/P0001 ,
		_w12842_,
		_w27021_
	);
	LUT2 #(
		.INIT('h8)
	) name16510 (
		\wishbone_bd_ram_mem1_reg[208][9]/P0001 ,
		_w13032_,
		_w27022_
	);
	LUT2 #(
		.INIT('h8)
	) name16511 (
		\wishbone_bd_ram_mem1_reg[85][9]/P0001 ,
		_w13216_,
		_w27023_
	);
	LUT2 #(
		.INIT('h8)
	) name16512 (
		\wishbone_bd_ram_mem1_reg[17][9]/P0001 ,
		_w12848_,
		_w27024_
	);
	LUT2 #(
		.INIT('h8)
	) name16513 (
		\wishbone_bd_ram_mem1_reg[134][9]/P0001 ,
		_w12763_,
		_w27025_
	);
	LUT2 #(
		.INIT('h8)
	) name16514 (
		\wishbone_bd_ram_mem1_reg[170][9]/P0001 ,
		_w13030_,
		_w27026_
	);
	LUT2 #(
		.INIT('h8)
	) name16515 (
		\wishbone_bd_ram_mem1_reg[45][9]/P0001 ,
		_w12908_,
		_w27027_
	);
	LUT2 #(
		.INIT('h8)
	) name16516 (
		\wishbone_bd_ram_mem1_reg[120][9]/P0001 ,
		_w12707_,
		_w27028_
	);
	LUT2 #(
		.INIT('h8)
	) name16517 (
		\wishbone_bd_ram_mem1_reg[10][9]/P0001 ,
		_w13172_,
		_w27029_
	);
	LUT2 #(
		.INIT('h8)
	) name16518 (
		\wishbone_bd_ram_mem1_reg[83][9]/P0001 ,
		_w12916_,
		_w27030_
	);
	LUT2 #(
		.INIT('h8)
	) name16519 (
		\wishbone_bd_ram_mem1_reg[21][9]/P0001 ,
		_w12906_,
		_w27031_
	);
	LUT2 #(
		.INIT('h8)
	) name16520 (
		\wishbone_bd_ram_mem1_reg[156][9]/P0001 ,
		_w13190_,
		_w27032_
	);
	LUT2 #(
		.INIT('h8)
	) name16521 (
		\wishbone_bd_ram_mem1_reg[132][9]/P0001 ,
		_w12992_,
		_w27033_
	);
	LUT2 #(
		.INIT('h8)
	) name16522 (
		\wishbone_bd_ram_mem1_reg[86][9]/P0001 ,
		_w12735_,
		_w27034_
	);
	LUT2 #(
		.INIT('h8)
	) name16523 (
		\wishbone_bd_ram_mem1_reg[117][9]/P0001 ,
		_w12715_,
		_w27035_
	);
	LUT2 #(
		.INIT('h8)
	) name16524 (
		\wishbone_bd_ram_mem1_reg[56][9]/P0001 ,
		_w12778_,
		_w27036_
	);
	LUT2 #(
		.INIT('h8)
	) name16525 (
		\wishbone_bd_ram_mem1_reg[197][9]/P0001 ,
		_w12834_,
		_w27037_
	);
	LUT2 #(
		.INIT('h8)
	) name16526 (
		\wishbone_bd_ram_mem1_reg[64][9]/P0001 ,
		_w12976_,
		_w27038_
	);
	LUT2 #(
		.INIT('h8)
	) name16527 (
		\wishbone_bd_ram_mem1_reg[206][9]/P0001 ,
		_w12954_,
		_w27039_
	);
	LUT2 #(
		.INIT('h8)
	) name16528 (
		\wishbone_bd_ram_mem1_reg[102][9]/P0001 ,
		_w12685_,
		_w27040_
	);
	LUT2 #(
		.INIT('h8)
	) name16529 (
		\wishbone_bd_ram_mem1_reg[223][9]/P0001 ,
		_w12838_,
		_w27041_
	);
	LUT2 #(
		.INIT('h8)
	) name16530 (
		\wishbone_bd_ram_mem1_reg[87][9]/P0001 ,
		_w13154_,
		_w27042_
	);
	LUT2 #(
		.INIT('h8)
	) name16531 (
		\wishbone_bd_ram_mem1_reg[97][9]/P0001 ,
		_w13096_,
		_w27043_
	);
	LUT2 #(
		.INIT('h8)
	) name16532 (
		\wishbone_bd_ram_mem1_reg[4][9]/P0001 ,
		_w12666_,
		_w27044_
	);
	LUT2 #(
		.INIT('h8)
	) name16533 (
		\wishbone_bd_ram_mem1_reg[202][9]/P0001 ,
		_w12870_,
		_w27045_
	);
	LUT2 #(
		.INIT('h8)
	) name16534 (
		\wishbone_bd_ram_mem1_reg[217][9]/P0001 ,
		_w13188_,
		_w27046_
	);
	LUT2 #(
		.INIT('h8)
	) name16535 (
		\wishbone_bd_ram_mem1_reg[157][9]/P0001 ,
		_w12926_,
		_w27047_
	);
	LUT2 #(
		.INIT('h8)
	) name16536 (
		\wishbone_bd_ram_mem1_reg[215][9]/P0001 ,
		_w12974_,
		_w27048_
	);
	LUT2 #(
		.INIT('h8)
	) name16537 (
		\wishbone_bd_ram_mem1_reg[189][9]/P0001 ,
		_w13042_,
		_w27049_
	);
	LUT2 #(
		.INIT('h8)
	) name16538 (
		\wishbone_bd_ram_mem1_reg[181][9]/P0001 ,
		_w12828_,
		_w27050_
	);
	LUT2 #(
		.INIT('h8)
	) name16539 (
		\wishbone_bd_ram_mem1_reg[129][9]/P0001 ,
		_w12776_,
		_w27051_
	);
	LUT2 #(
		.INIT('h8)
	) name16540 (
		\wishbone_bd_ram_mem1_reg[235][9]/P0001 ,
		_w12696_,
		_w27052_
	);
	LUT2 #(
		.INIT('h8)
	) name16541 (
		\wishbone_bd_ram_mem1_reg[96][9]/P0001 ,
		_w12912_,
		_w27053_
	);
	LUT2 #(
		.INIT('h8)
	) name16542 (
		\wishbone_bd_ram_mem1_reg[81][9]/P0001 ,
		_w12950_,
		_w27054_
	);
	LUT2 #(
		.INIT('h8)
	) name16543 (
		\wishbone_bd_ram_mem1_reg[14][9]/P0001 ,
		_w13086_,
		_w27055_
	);
	LUT2 #(
		.INIT('h8)
	) name16544 (
		\wishbone_bd_ram_mem1_reg[66][9]/P0001 ,
		_w12824_,
		_w27056_
	);
	LUT2 #(
		.INIT('h8)
	) name16545 (
		\wishbone_bd_ram_mem1_reg[43][9]/P0001 ,
		_w13200_,
		_w27057_
	);
	LUT2 #(
		.INIT('h8)
	) name16546 (
		\wishbone_bd_ram_mem1_reg[70][9]/P0001 ,
		_w12840_,
		_w27058_
	);
	LUT2 #(
		.INIT('h8)
	) name16547 (
		\wishbone_bd_ram_mem1_reg[60][9]/P0001 ,
		_w13204_,
		_w27059_
	);
	LUT2 #(
		.INIT('h8)
	) name16548 (
		\wishbone_bd_ram_mem1_reg[88][9]/P0001 ,
		_w12860_,
		_w27060_
	);
	LUT2 #(
		.INIT('h8)
	) name16549 (
		\wishbone_bd_ram_mem1_reg[69][9]/P0001 ,
		_w12738_,
		_w27061_
	);
	LUT2 #(
		.INIT('h8)
	) name16550 (
		\wishbone_bd_ram_mem1_reg[108][9]/P0001 ,
		_w13156_,
		_w27062_
	);
	LUT2 #(
		.INIT('h8)
	) name16551 (
		\wishbone_bd_ram_mem1_reg[248][9]/P0001 ,
		_w12789_,
		_w27063_
	);
	LUT2 #(
		.INIT('h8)
	) name16552 (
		\wishbone_bd_ram_mem1_reg[101][9]/P0001 ,
		_w13192_,
		_w27064_
	);
	LUT2 #(
		.INIT('h8)
	) name16553 (
		\wishbone_bd_ram_mem1_reg[203][9]/P0001 ,
		_w13158_,
		_w27065_
	);
	LUT2 #(
		.INIT('h8)
	) name16554 (
		\wishbone_bd_ram_mem1_reg[234][9]/P0001 ,
		_w13214_,
		_w27066_
	);
	LUT2 #(
		.INIT('h8)
	) name16555 (
		\wishbone_bd_ram_mem1_reg[198][9]/P0001 ,
		_w12832_,
		_w27067_
	);
	LUT2 #(
		.INIT('h8)
	) name16556 (
		\wishbone_bd_ram_mem1_reg[131][9]/P0001 ,
		_w12852_,
		_w27068_
	);
	LUT2 #(
		.INIT('h8)
	) name16557 (
		\wishbone_bd_ram_mem1_reg[145][9]/P0001 ,
		_w13106_,
		_w27069_
	);
	LUT2 #(
		.INIT('h8)
	) name16558 (
		\wishbone_bd_ram_mem1_reg[218][9]/P0001 ,
		_w13206_,
		_w27070_
	);
	LUT2 #(
		.INIT('h8)
	) name16559 (
		\wishbone_bd_ram_mem1_reg[78][9]/P0001 ,
		_w12874_,
		_w27071_
	);
	LUT2 #(
		.INIT('h8)
	) name16560 (
		\wishbone_bd_ram_mem1_reg[53][9]/P0001 ,
		_w13020_,
		_w27072_
	);
	LUT2 #(
		.INIT('h8)
	) name16561 (
		\wishbone_bd_ram_mem1_reg[26][9]/P0001 ,
		_w12699_,
		_w27073_
	);
	LUT2 #(
		.INIT('h8)
	) name16562 (
		\wishbone_bd_ram_mem1_reg[124][9]/P0001 ,
		_w13058_,
		_w27074_
	);
	LUT2 #(
		.INIT('h8)
	) name16563 (
		\wishbone_bd_ram_mem1_reg[33][9]/P0001 ,
		_w12980_,
		_w27075_
	);
	LUT2 #(
		.INIT('h8)
	) name16564 (
		\wishbone_bd_ram_mem1_reg[112][9]/P0001 ,
		_w12733_,
		_w27076_
	);
	LUT2 #(
		.INIT('h8)
	) name16565 (
		\wishbone_bd_ram_mem1_reg[15][9]/P0001 ,
		_w13210_,
		_w27077_
	);
	LUT2 #(
		.INIT('h8)
	) name16566 (
		\wishbone_bd_ram_mem1_reg[8][9]/P0001 ,
		_w12920_,
		_w27078_
	);
	LUT2 #(
		.INIT('h8)
	) name16567 (
		\wishbone_bd_ram_mem1_reg[169][9]/P0001 ,
		_w12722_,
		_w27079_
	);
	LUT2 #(
		.INIT('h8)
	) name16568 (
		\wishbone_bd_ram_mem1_reg[141][9]/P0001 ,
		_w13004_,
		_w27080_
	);
	LUT2 #(
		.INIT('h8)
	) name16569 (
		\wishbone_bd_ram_mem1_reg[155][9]/P0001 ,
		_w13122_,
		_w27081_
	);
	LUT2 #(
		.INIT('h8)
	) name16570 (
		\wishbone_bd_ram_mem1_reg[163][9]/P0001 ,
		_w12882_,
		_w27082_
	);
	LUT2 #(
		.INIT('h8)
	) name16571 (
		\wishbone_bd_ram_mem1_reg[74][9]/P0001 ,
		_w12812_,
		_w27083_
	);
	LUT2 #(
		.INIT('h8)
	) name16572 (
		\wishbone_bd_ram_mem1_reg[212][9]/P0001 ,
		_w12796_,
		_w27084_
	);
	LUT2 #(
		.INIT('h8)
	) name16573 (
		\wishbone_bd_ram_mem1_reg[240][9]/P0001 ,
		_w12864_,
		_w27085_
	);
	LUT2 #(
		.INIT('h8)
	) name16574 (
		\wishbone_bd_ram_mem1_reg[114][9]/P0001 ,
		_w13202_,
		_w27086_
	);
	LUT2 #(
		.INIT('h8)
	) name16575 (
		\wishbone_bd_ram_mem1_reg[150][9]/P0001 ,
		_w13136_,
		_w27087_
	);
	LUT2 #(
		.INIT('h8)
	) name16576 (
		\wishbone_bd_ram_mem1_reg[242][9]/P0001 ,
		_w12932_,
		_w27088_
	);
	LUT2 #(
		.INIT('h8)
	) name16577 (
		\wishbone_bd_ram_mem1_reg[153][9]/P0001 ,
		_w12890_,
		_w27089_
	);
	LUT2 #(
		.INIT('h8)
	) name16578 (
		\wishbone_bd_ram_mem1_reg[122][9]/P0001 ,
		_w13130_,
		_w27090_
	);
	LUT2 #(
		.INIT('h8)
	) name16579 (
		\wishbone_bd_ram_mem1_reg[98][9]/P0001 ,
		_w12816_,
		_w27091_
	);
	LUT2 #(
		.INIT('h8)
	) name16580 (
		\wishbone_bd_ram_mem1_reg[110][9]/P0001 ,
		_w13046_,
		_w27092_
	);
	LUT2 #(
		.INIT('h8)
	) name16581 (
		\wishbone_bd_ram_mem1_reg[63][9]/P0001 ,
		_w12850_,
		_w27093_
	);
	LUT2 #(
		.INIT('h8)
	) name16582 (
		\wishbone_bd_ram_mem1_reg[176][9]/P0001 ,
		_w12868_,
		_w27094_
	);
	LUT2 #(
		.INIT('h8)
	) name16583 (
		\wishbone_bd_ram_mem1_reg[41][9]/P0001 ,
		_w13052_,
		_w27095_
	);
	LUT2 #(
		.INIT('h8)
	) name16584 (
		\wishbone_bd_ram_mem1_reg[199][9]/P0001 ,
		_w12768_,
		_w27096_
	);
	LUT2 #(
		.INIT('h8)
	) name16585 (
		\wishbone_bd_ram_mem1_reg[76][9]/P0001 ,
		_w13184_,
		_w27097_
	);
	LUT2 #(
		.INIT('h8)
	) name16586 (
		\wishbone_bd_ram_mem1_reg[214][9]/P0001 ,
		_w12984_,
		_w27098_
	);
	LUT2 #(
		.INIT('h8)
	) name16587 (
		\wishbone_bd_ram_mem1_reg[210][9]/P0001 ,
		_w12924_,
		_w27099_
	);
	LUT2 #(
		.INIT('h8)
	) name16588 (
		\wishbone_bd_ram_mem1_reg[188][9]/P0001 ,
		_w12948_,
		_w27100_
	);
	LUT2 #(
		.INIT('h8)
	) name16589 (
		\wishbone_bd_ram_mem1_reg[125][9]/P0001 ,
		_w12956_,
		_w27101_
	);
	LUT2 #(
		.INIT('h8)
	) name16590 (
		\wishbone_bd_ram_mem1_reg[91][9]/P0001 ,
		_w13074_,
		_w27102_
	);
	LUT2 #(
		.INIT('h8)
	) name16591 (
		\wishbone_bd_ram_mem1_reg[152][9]/P0001 ,
		_w12966_,
		_w27103_
	);
	LUT2 #(
		.INIT('h8)
	) name16592 (
		\wishbone_bd_ram_mem1_reg[94][9]/P0001 ,
		_w13186_,
		_w27104_
	);
	LUT2 #(
		.INIT('h8)
	) name16593 (
		\wishbone_bd_ram_mem1_reg[211][9]/P0001 ,
		_w13166_,
		_w27105_
	);
	LUT2 #(
		.INIT('h8)
	) name16594 (
		\wishbone_bd_ram_mem1_reg[187][9]/P0001 ,
		_w13196_,
		_w27106_
	);
	LUT2 #(
		.INIT('h8)
	) name16595 (
		\wishbone_bd_ram_mem1_reg[140][9]/P0001 ,
		_w12894_,
		_w27107_
	);
	LUT2 #(
		.INIT('h8)
	) name16596 (
		\wishbone_bd_ram_mem1_reg[162][9]/P0001 ,
		_w13098_,
		_w27108_
	);
	LUT2 #(
		.INIT('h8)
	) name16597 (
		\wishbone_bd_ram_mem1_reg[233][9]/P0001 ,
		_w12836_,
		_w27109_
	);
	LUT2 #(
		.INIT('h8)
	) name16598 (
		\wishbone_bd_ram_mem1_reg[143][9]/P0001 ,
		_w12922_,
		_w27110_
	);
	LUT2 #(
		.INIT('h8)
	) name16599 (
		\wishbone_bd_ram_mem1_reg[226][9]/P0001 ,
		_w13138_,
		_w27111_
	);
	LUT2 #(
		.INIT('h8)
	) name16600 (
		\wishbone_bd_ram_mem1_reg[18][9]/P0001 ,
		_w12679_,
		_w27112_
	);
	LUT2 #(
		.INIT('h8)
	) name16601 (
		\wishbone_bd_ram_mem1_reg[12][9]/P0001 ,
		_w13118_,
		_w27113_
	);
	LUT2 #(
		.INIT('h8)
	) name16602 (
		\wishbone_bd_ram_mem1_reg[35][9]/P0001 ,
		_w12703_,
		_w27114_
	);
	LUT2 #(
		.INIT('h8)
	) name16603 (
		\wishbone_bd_ram_mem1_reg[16][9]/P0001 ,
		_w13140_,
		_w27115_
	);
	LUT2 #(
		.INIT('h8)
	) name16604 (
		\wishbone_bd_ram_mem1_reg[103][9]/P0001 ,
		_w12846_,
		_w27116_
	);
	LUT2 #(
		.INIT('h8)
	) name16605 (
		\wishbone_bd_ram_mem1_reg[190][9]/P0001 ,
		_w12858_,
		_w27117_
	);
	LUT2 #(
		.INIT('h8)
	) name16606 (
		\wishbone_bd_ram_mem1_reg[253][9]/P0001 ,
		_w13100_,
		_w27118_
	);
	LUT2 #(
		.INIT('h8)
	) name16607 (
		\wishbone_bd_ram_mem1_reg[158][9]/P0001 ,
		_w12898_,
		_w27119_
	);
	LUT2 #(
		.INIT('h8)
	) name16608 (
		\wishbone_bd_ram_mem1_reg[38][9]/P0001 ,
		_w13182_,
		_w27120_
	);
	LUT2 #(
		.INIT('h8)
	) name16609 (
		\wishbone_bd_ram_mem1_reg[221][9]/P0001 ,
		_w12802_,
		_w27121_
	);
	LUT2 #(
		.INIT('h8)
	) name16610 (
		\wishbone_bd_ram_mem1_reg[72][9]/P0001 ,
		_w12810_,
		_w27122_
	);
	LUT2 #(
		.INIT('h8)
	) name16611 (
		\wishbone_bd_ram_mem1_reg[37][9]/P0001 ,
		_w13102_,
		_w27123_
	);
	LUT2 #(
		.INIT('h8)
	) name16612 (
		\wishbone_bd_ram_mem1_reg[161][9]/P0001 ,
		_w12754_,
		_w27124_
	);
	LUT2 #(
		.INIT('h8)
	) name16613 (
		\wishbone_bd_ram_mem1_reg[6][9]/P0001 ,
		_w12968_,
		_w27125_
	);
	LUT2 #(
		.INIT('h8)
	) name16614 (
		\wishbone_bd_ram_mem1_reg[51][9]/P0001 ,
		_w13024_,
		_w27126_
	);
	LUT2 #(
		.INIT('h8)
	) name16615 (
		\wishbone_bd_ram_mem1_reg[147][9]/P0001 ,
		_w13146_,
		_w27127_
	);
	LUT2 #(
		.INIT('h8)
	) name16616 (
		\wishbone_bd_ram_mem1_reg[230][9]/P0001 ,
		_w13036_,
		_w27128_
	);
	LUT2 #(
		.INIT('h8)
	) name16617 (
		\wishbone_bd_ram_mem1_reg[135][9]/P0001 ,
		_w13124_,
		_w27129_
	);
	LUT2 #(
		.INIT('h8)
	) name16618 (
		\wishbone_bd_ram_mem1_reg[5][9]/P0001 ,
		_w12878_,
		_w27130_
	);
	LUT2 #(
		.INIT('h8)
	) name16619 (
		\wishbone_bd_ram_mem1_reg[28][9]/P0001 ,
		_w13170_,
		_w27131_
	);
	LUT2 #(
		.INIT('h8)
	) name16620 (
		\wishbone_bd_ram_mem1_reg[159][9]/P0001 ,
		_w12774_,
		_w27132_
	);
	LUT2 #(
		.INIT('h8)
	) name16621 (
		\wishbone_bd_ram_mem1_reg[148][9]/P0001 ,
		_w13000_,
		_w27133_
	);
	LUT2 #(
		.INIT('h8)
	) name16622 (
		\wishbone_bd_ram_mem1_reg[58][9]/P0001 ,
		_w13070_,
		_w27134_
	);
	LUT2 #(
		.INIT('h8)
	) name16623 (
		\wishbone_bd_ram_mem1_reg[245][9]/P0001 ,
		_w13022_,
		_w27135_
	);
	LUT2 #(
		.INIT('h8)
	) name16624 (
		\wishbone_bd_ram_mem1_reg[137][9]/P0001 ,
		_w13168_,
		_w27136_
	);
	LUT2 #(
		.INIT('h8)
	) name16625 (
		\wishbone_bd_ram_mem1_reg[0][9]/P0001 ,
		_w12717_,
		_w27137_
	);
	LUT2 #(
		.INIT('h8)
	) name16626 (
		\wishbone_bd_ram_mem1_reg[164][9]/P0001 ,
		_w12876_,
		_w27138_
	);
	LUT2 #(
		.INIT('h8)
	) name16627 (
		\wishbone_bd_ram_mem1_reg[65][9]/P0001 ,
		_w13176_,
		_w27139_
	);
	LUT2 #(
		.INIT('h8)
	) name16628 (
		\wishbone_bd_ram_mem1_reg[47][9]/P0001 ,
		_w12904_,
		_w27140_
	);
	LUT2 #(
		.INIT('h8)
	) name16629 (
		\wishbone_bd_ram_mem1_reg[113][9]/P0001 ,
		_w13026_,
		_w27141_
	);
	LUT2 #(
		.INIT('h8)
	) name16630 (
		\wishbone_bd_ram_mem1_reg[192][9]/P0001 ,
		_w12938_,
		_w27142_
	);
	LUT2 #(
		.INIT('h8)
	) name16631 (
		\wishbone_bd_ram_mem1_reg[222][9]/P0001 ,
		_w13094_,
		_w27143_
	);
	LUT2 #(
		.INIT('h8)
	) name16632 (
		\wishbone_bd_ram_mem1_reg[75][9]/P0001 ,
		_w12826_,
		_w27144_
	);
	LUT2 #(
		.INIT('h8)
	) name16633 (
		\wishbone_bd_ram_mem1_reg[182][9]/P0001 ,
		_w12820_,
		_w27145_
	);
	LUT2 #(
		.INIT('h8)
	) name16634 (
		\wishbone_bd_ram_mem1_reg[67][9]/P0001 ,
		_w13134_,
		_w27146_
	);
	LUT2 #(
		.INIT('h8)
	) name16635 (
		\wishbone_bd_ram_mem1_reg[24][9]/P0001 ,
		_w13084_,
		_w27147_
	);
	LUT2 #(
		.INIT('h8)
	) name16636 (
		\wishbone_bd_ram_mem1_reg[71][9]/P0001 ,
		_w12798_,
		_w27148_
	);
	LUT2 #(
		.INIT('h8)
	) name16637 (
		\wishbone_bd_ram_mem1_reg[177][9]/P0001 ,
		_w12996_,
		_w27149_
	);
	LUT2 #(
		.INIT('h8)
	) name16638 (
		\wishbone_bd_ram_mem1_reg[247][9]/P0001 ,
		_w12818_,
		_w27150_
	);
	LUT2 #(
		.INIT('h8)
	) name16639 (
		\wishbone_bd_ram_mem1_reg[229][9]/P0001 ,
		_w12711_,
		_w27151_
	);
	LUT2 #(
		.INIT('h8)
	) name16640 (
		\wishbone_bd_ram_mem1_reg[175][9]/P0001 ,
		_w13126_,
		_w27152_
	);
	LUT2 #(
		.INIT('h8)
	) name16641 (
		\wishbone_bd_ram_mem1_reg[200][9]/P0001 ,
		_w12988_,
		_w27153_
	);
	LUT2 #(
		.INIT('h8)
	) name16642 (
		\wishbone_bd_ram_mem1_reg[179][9]/P0001 ,
		_w13050_,
		_w27154_
	);
	LUT2 #(
		.INIT('h8)
	) name16643 (
		\wishbone_bd_ram_mem1_reg[59][9]/P0001 ,
		_w12780_,
		_w27155_
	);
	LUT2 #(
		.INIT('h8)
	) name16644 (
		\wishbone_bd_ram_mem1_reg[11][9]/P0001 ,
		_w13194_,
		_w27156_
	);
	LUT2 #(
		.INIT('h8)
	) name16645 (
		\wishbone_bd_ram_mem1_reg[46][9]/P0001 ,
		_w12884_,
		_w27157_
	);
	LUT2 #(
		.INIT('h8)
	) name16646 (
		\wishbone_bd_ram_mem1_reg[232][9]/P0001 ,
		_w12758_,
		_w27158_
	);
	LUT2 #(
		.INIT('h8)
	) name16647 (
		\wishbone_bd_ram_mem1_reg[79][9]/P0001 ,
		_w13212_,
		_w27159_
	);
	LUT2 #(
		.INIT('h8)
	) name16648 (
		\wishbone_bd_ram_mem1_reg[50][9]/P0001 ,
		_w13150_,
		_w27160_
	);
	LUT2 #(
		.INIT('h8)
	) name16649 (
		\wishbone_bd_ram_mem1_reg[225][9]/P0001 ,
		_w13092_,
		_w27161_
	);
	LUT2 #(
		.INIT('h8)
	) name16650 (
		\wishbone_bd_ram_mem1_reg[62][9]/P0001 ,
		_w12673_,
		_w27162_
	);
	LUT2 #(
		.INIT('h8)
	) name16651 (
		\wishbone_bd_ram_mem1_reg[219][9]/P0001 ,
		_w12806_,
		_w27163_
	);
	LUT2 #(
		.INIT('h8)
	) name16652 (
		\wishbone_bd_ram_mem1_reg[172][9]/P0001 ,
		_w12944_,
		_w27164_
	);
	LUT2 #(
		.INIT('h8)
	) name16653 (
		\wishbone_bd_ram_mem1_reg[31][9]/P0001 ,
		_w13198_,
		_w27165_
	);
	LUT2 #(
		.INIT('h8)
	) name16654 (
		\wishbone_bd_ram_mem1_reg[89][9]/P0001 ,
		_w12964_,
		_w27166_
	);
	LUT2 #(
		.INIT('h8)
	) name16655 (
		\wishbone_bd_ram_mem1_reg[136][9]/P0001 ,
		_w13064_,
		_w27167_
	);
	LUT2 #(
		.INIT('h8)
	) name16656 (
		\wishbone_bd_ram_mem1_reg[23][9]/P0001 ,
		_w13008_,
		_w27168_
	);
	LUT2 #(
		.INIT('h8)
	) name16657 (
		\wishbone_bd_ram_mem1_reg[239][9]/P0001 ,
		_w12862_,
		_w27169_
	);
	LUT2 #(
		.INIT('h8)
	) name16658 (
		\wishbone_bd_ram_mem1_reg[19][9]/P0001 ,
		_w13012_,
		_w27170_
	);
	LUT2 #(
		.INIT('h8)
	) name16659 (
		\wishbone_bd_ram_mem1_reg[44][9]/P0001 ,
		_w12896_,
		_w27171_
	);
	LUT2 #(
		.INIT('h8)
	) name16660 (
		\wishbone_bd_ram_mem1_reg[191][9]/P0001 ,
		_w13034_,
		_w27172_
	);
	LUT2 #(
		.INIT('h8)
	) name16661 (
		\wishbone_bd_ram_mem1_reg[128][9]/P0001 ,
		_w12793_,
		_w27173_
	);
	LUT2 #(
		.INIT('h8)
	) name16662 (
		\wishbone_bd_ram_mem1_reg[93][9]/P0001 ,
		_w13016_,
		_w27174_
	);
	LUT2 #(
		.INIT('h8)
	) name16663 (
		\wishbone_bd_ram_mem1_reg[105][9]/P0001 ,
		_w12751_,
		_w27175_
	);
	LUT2 #(
		.INIT('h8)
	) name16664 (
		\wishbone_bd_ram_mem1_reg[243][9]/P0001 ,
		_w12804_,
		_w27176_
	);
	LUT2 #(
		.INIT('h8)
	) name16665 (
		\wishbone_bd_ram_mem1_reg[3][9]/P0001 ,
		_w12866_,
		_w27177_
	);
	LUT2 #(
		.INIT('h8)
	) name16666 (
		\wishbone_bd_ram_mem1_reg[216][9]/P0001 ,
		_w13028_,
		_w27178_
	);
	LUT2 #(
		.INIT('h8)
	) name16667 (
		\wishbone_bd_ram_mem1_reg[104][9]/P0001 ,
		_w13148_,
		_w27179_
	);
	LUT2 #(
		.INIT('h8)
	) name16668 (
		\wishbone_bd_ram_mem1_reg[183][9]/P0001 ,
		_w12787_,
		_w27180_
	);
	LUT2 #(
		.INIT('h1)
	) name16669 (
		_w26925_,
		_w26926_,
		_w27181_
	);
	LUT2 #(
		.INIT('h1)
	) name16670 (
		_w26927_,
		_w26928_,
		_w27182_
	);
	LUT2 #(
		.INIT('h1)
	) name16671 (
		_w26929_,
		_w26930_,
		_w27183_
	);
	LUT2 #(
		.INIT('h1)
	) name16672 (
		_w26931_,
		_w26932_,
		_w27184_
	);
	LUT2 #(
		.INIT('h1)
	) name16673 (
		_w26933_,
		_w26934_,
		_w27185_
	);
	LUT2 #(
		.INIT('h1)
	) name16674 (
		_w26935_,
		_w26936_,
		_w27186_
	);
	LUT2 #(
		.INIT('h1)
	) name16675 (
		_w26937_,
		_w26938_,
		_w27187_
	);
	LUT2 #(
		.INIT('h1)
	) name16676 (
		_w26939_,
		_w26940_,
		_w27188_
	);
	LUT2 #(
		.INIT('h1)
	) name16677 (
		_w26941_,
		_w26942_,
		_w27189_
	);
	LUT2 #(
		.INIT('h1)
	) name16678 (
		_w26943_,
		_w26944_,
		_w27190_
	);
	LUT2 #(
		.INIT('h1)
	) name16679 (
		_w26945_,
		_w26946_,
		_w27191_
	);
	LUT2 #(
		.INIT('h1)
	) name16680 (
		_w26947_,
		_w26948_,
		_w27192_
	);
	LUT2 #(
		.INIT('h1)
	) name16681 (
		_w26949_,
		_w26950_,
		_w27193_
	);
	LUT2 #(
		.INIT('h1)
	) name16682 (
		_w26951_,
		_w26952_,
		_w27194_
	);
	LUT2 #(
		.INIT('h1)
	) name16683 (
		_w26953_,
		_w26954_,
		_w27195_
	);
	LUT2 #(
		.INIT('h1)
	) name16684 (
		_w26955_,
		_w26956_,
		_w27196_
	);
	LUT2 #(
		.INIT('h1)
	) name16685 (
		_w26957_,
		_w26958_,
		_w27197_
	);
	LUT2 #(
		.INIT('h1)
	) name16686 (
		_w26959_,
		_w26960_,
		_w27198_
	);
	LUT2 #(
		.INIT('h1)
	) name16687 (
		_w26961_,
		_w26962_,
		_w27199_
	);
	LUT2 #(
		.INIT('h1)
	) name16688 (
		_w26963_,
		_w26964_,
		_w27200_
	);
	LUT2 #(
		.INIT('h1)
	) name16689 (
		_w26965_,
		_w26966_,
		_w27201_
	);
	LUT2 #(
		.INIT('h1)
	) name16690 (
		_w26967_,
		_w26968_,
		_w27202_
	);
	LUT2 #(
		.INIT('h1)
	) name16691 (
		_w26969_,
		_w26970_,
		_w27203_
	);
	LUT2 #(
		.INIT('h1)
	) name16692 (
		_w26971_,
		_w26972_,
		_w27204_
	);
	LUT2 #(
		.INIT('h1)
	) name16693 (
		_w26973_,
		_w26974_,
		_w27205_
	);
	LUT2 #(
		.INIT('h1)
	) name16694 (
		_w26975_,
		_w26976_,
		_w27206_
	);
	LUT2 #(
		.INIT('h1)
	) name16695 (
		_w26977_,
		_w26978_,
		_w27207_
	);
	LUT2 #(
		.INIT('h1)
	) name16696 (
		_w26979_,
		_w26980_,
		_w27208_
	);
	LUT2 #(
		.INIT('h1)
	) name16697 (
		_w26981_,
		_w26982_,
		_w27209_
	);
	LUT2 #(
		.INIT('h1)
	) name16698 (
		_w26983_,
		_w26984_,
		_w27210_
	);
	LUT2 #(
		.INIT('h1)
	) name16699 (
		_w26985_,
		_w26986_,
		_w27211_
	);
	LUT2 #(
		.INIT('h1)
	) name16700 (
		_w26987_,
		_w26988_,
		_w27212_
	);
	LUT2 #(
		.INIT('h1)
	) name16701 (
		_w26989_,
		_w26990_,
		_w27213_
	);
	LUT2 #(
		.INIT('h1)
	) name16702 (
		_w26991_,
		_w26992_,
		_w27214_
	);
	LUT2 #(
		.INIT('h1)
	) name16703 (
		_w26993_,
		_w26994_,
		_w27215_
	);
	LUT2 #(
		.INIT('h1)
	) name16704 (
		_w26995_,
		_w26996_,
		_w27216_
	);
	LUT2 #(
		.INIT('h1)
	) name16705 (
		_w26997_,
		_w26998_,
		_w27217_
	);
	LUT2 #(
		.INIT('h1)
	) name16706 (
		_w26999_,
		_w27000_,
		_w27218_
	);
	LUT2 #(
		.INIT('h1)
	) name16707 (
		_w27001_,
		_w27002_,
		_w27219_
	);
	LUT2 #(
		.INIT('h1)
	) name16708 (
		_w27003_,
		_w27004_,
		_w27220_
	);
	LUT2 #(
		.INIT('h1)
	) name16709 (
		_w27005_,
		_w27006_,
		_w27221_
	);
	LUT2 #(
		.INIT('h1)
	) name16710 (
		_w27007_,
		_w27008_,
		_w27222_
	);
	LUT2 #(
		.INIT('h1)
	) name16711 (
		_w27009_,
		_w27010_,
		_w27223_
	);
	LUT2 #(
		.INIT('h1)
	) name16712 (
		_w27011_,
		_w27012_,
		_w27224_
	);
	LUT2 #(
		.INIT('h1)
	) name16713 (
		_w27013_,
		_w27014_,
		_w27225_
	);
	LUT2 #(
		.INIT('h1)
	) name16714 (
		_w27015_,
		_w27016_,
		_w27226_
	);
	LUT2 #(
		.INIT('h1)
	) name16715 (
		_w27017_,
		_w27018_,
		_w27227_
	);
	LUT2 #(
		.INIT('h1)
	) name16716 (
		_w27019_,
		_w27020_,
		_w27228_
	);
	LUT2 #(
		.INIT('h1)
	) name16717 (
		_w27021_,
		_w27022_,
		_w27229_
	);
	LUT2 #(
		.INIT('h1)
	) name16718 (
		_w27023_,
		_w27024_,
		_w27230_
	);
	LUT2 #(
		.INIT('h1)
	) name16719 (
		_w27025_,
		_w27026_,
		_w27231_
	);
	LUT2 #(
		.INIT('h1)
	) name16720 (
		_w27027_,
		_w27028_,
		_w27232_
	);
	LUT2 #(
		.INIT('h1)
	) name16721 (
		_w27029_,
		_w27030_,
		_w27233_
	);
	LUT2 #(
		.INIT('h1)
	) name16722 (
		_w27031_,
		_w27032_,
		_w27234_
	);
	LUT2 #(
		.INIT('h1)
	) name16723 (
		_w27033_,
		_w27034_,
		_w27235_
	);
	LUT2 #(
		.INIT('h1)
	) name16724 (
		_w27035_,
		_w27036_,
		_w27236_
	);
	LUT2 #(
		.INIT('h1)
	) name16725 (
		_w27037_,
		_w27038_,
		_w27237_
	);
	LUT2 #(
		.INIT('h1)
	) name16726 (
		_w27039_,
		_w27040_,
		_w27238_
	);
	LUT2 #(
		.INIT('h1)
	) name16727 (
		_w27041_,
		_w27042_,
		_w27239_
	);
	LUT2 #(
		.INIT('h1)
	) name16728 (
		_w27043_,
		_w27044_,
		_w27240_
	);
	LUT2 #(
		.INIT('h1)
	) name16729 (
		_w27045_,
		_w27046_,
		_w27241_
	);
	LUT2 #(
		.INIT('h1)
	) name16730 (
		_w27047_,
		_w27048_,
		_w27242_
	);
	LUT2 #(
		.INIT('h1)
	) name16731 (
		_w27049_,
		_w27050_,
		_w27243_
	);
	LUT2 #(
		.INIT('h1)
	) name16732 (
		_w27051_,
		_w27052_,
		_w27244_
	);
	LUT2 #(
		.INIT('h1)
	) name16733 (
		_w27053_,
		_w27054_,
		_w27245_
	);
	LUT2 #(
		.INIT('h1)
	) name16734 (
		_w27055_,
		_w27056_,
		_w27246_
	);
	LUT2 #(
		.INIT('h1)
	) name16735 (
		_w27057_,
		_w27058_,
		_w27247_
	);
	LUT2 #(
		.INIT('h1)
	) name16736 (
		_w27059_,
		_w27060_,
		_w27248_
	);
	LUT2 #(
		.INIT('h1)
	) name16737 (
		_w27061_,
		_w27062_,
		_w27249_
	);
	LUT2 #(
		.INIT('h1)
	) name16738 (
		_w27063_,
		_w27064_,
		_w27250_
	);
	LUT2 #(
		.INIT('h1)
	) name16739 (
		_w27065_,
		_w27066_,
		_w27251_
	);
	LUT2 #(
		.INIT('h1)
	) name16740 (
		_w27067_,
		_w27068_,
		_w27252_
	);
	LUT2 #(
		.INIT('h1)
	) name16741 (
		_w27069_,
		_w27070_,
		_w27253_
	);
	LUT2 #(
		.INIT('h1)
	) name16742 (
		_w27071_,
		_w27072_,
		_w27254_
	);
	LUT2 #(
		.INIT('h1)
	) name16743 (
		_w27073_,
		_w27074_,
		_w27255_
	);
	LUT2 #(
		.INIT('h1)
	) name16744 (
		_w27075_,
		_w27076_,
		_w27256_
	);
	LUT2 #(
		.INIT('h1)
	) name16745 (
		_w27077_,
		_w27078_,
		_w27257_
	);
	LUT2 #(
		.INIT('h1)
	) name16746 (
		_w27079_,
		_w27080_,
		_w27258_
	);
	LUT2 #(
		.INIT('h1)
	) name16747 (
		_w27081_,
		_w27082_,
		_w27259_
	);
	LUT2 #(
		.INIT('h1)
	) name16748 (
		_w27083_,
		_w27084_,
		_w27260_
	);
	LUT2 #(
		.INIT('h1)
	) name16749 (
		_w27085_,
		_w27086_,
		_w27261_
	);
	LUT2 #(
		.INIT('h1)
	) name16750 (
		_w27087_,
		_w27088_,
		_w27262_
	);
	LUT2 #(
		.INIT('h1)
	) name16751 (
		_w27089_,
		_w27090_,
		_w27263_
	);
	LUT2 #(
		.INIT('h1)
	) name16752 (
		_w27091_,
		_w27092_,
		_w27264_
	);
	LUT2 #(
		.INIT('h1)
	) name16753 (
		_w27093_,
		_w27094_,
		_w27265_
	);
	LUT2 #(
		.INIT('h1)
	) name16754 (
		_w27095_,
		_w27096_,
		_w27266_
	);
	LUT2 #(
		.INIT('h1)
	) name16755 (
		_w27097_,
		_w27098_,
		_w27267_
	);
	LUT2 #(
		.INIT('h1)
	) name16756 (
		_w27099_,
		_w27100_,
		_w27268_
	);
	LUT2 #(
		.INIT('h1)
	) name16757 (
		_w27101_,
		_w27102_,
		_w27269_
	);
	LUT2 #(
		.INIT('h1)
	) name16758 (
		_w27103_,
		_w27104_,
		_w27270_
	);
	LUT2 #(
		.INIT('h1)
	) name16759 (
		_w27105_,
		_w27106_,
		_w27271_
	);
	LUT2 #(
		.INIT('h1)
	) name16760 (
		_w27107_,
		_w27108_,
		_w27272_
	);
	LUT2 #(
		.INIT('h1)
	) name16761 (
		_w27109_,
		_w27110_,
		_w27273_
	);
	LUT2 #(
		.INIT('h1)
	) name16762 (
		_w27111_,
		_w27112_,
		_w27274_
	);
	LUT2 #(
		.INIT('h1)
	) name16763 (
		_w27113_,
		_w27114_,
		_w27275_
	);
	LUT2 #(
		.INIT('h1)
	) name16764 (
		_w27115_,
		_w27116_,
		_w27276_
	);
	LUT2 #(
		.INIT('h1)
	) name16765 (
		_w27117_,
		_w27118_,
		_w27277_
	);
	LUT2 #(
		.INIT('h1)
	) name16766 (
		_w27119_,
		_w27120_,
		_w27278_
	);
	LUT2 #(
		.INIT('h1)
	) name16767 (
		_w27121_,
		_w27122_,
		_w27279_
	);
	LUT2 #(
		.INIT('h1)
	) name16768 (
		_w27123_,
		_w27124_,
		_w27280_
	);
	LUT2 #(
		.INIT('h1)
	) name16769 (
		_w27125_,
		_w27126_,
		_w27281_
	);
	LUT2 #(
		.INIT('h1)
	) name16770 (
		_w27127_,
		_w27128_,
		_w27282_
	);
	LUT2 #(
		.INIT('h1)
	) name16771 (
		_w27129_,
		_w27130_,
		_w27283_
	);
	LUT2 #(
		.INIT('h1)
	) name16772 (
		_w27131_,
		_w27132_,
		_w27284_
	);
	LUT2 #(
		.INIT('h1)
	) name16773 (
		_w27133_,
		_w27134_,
		_w27285_
	);
	LUT2 #(
		.INIT('h1)
	) name16774 (
		_w27135_,
		_w27136_,
		_w27286_
	);
	LUT2 #(
		.INIT('h1)
	) name16775 (
		_w27137_,
		_w27138_,
		_w27287_
	);
	LUT2 #(
		.INIT('h1)
	) name16776 (
		_w27139_,
		_w27140_,
		_w27288_
	);
	LUT2 #(
		.INIT('h1)
	) name16777 (
		_w27141_,
		_w27142_,
		_w27289_
	);
	LUT2 #(
		.INIT('h1)
	) name16778 (
		_w27143_,
		_w27144_,
		_w27290_
	);
	LUT2 #(
		.INIT('h1)
	) name16779 (
		_w27145_,
		_w27146_,
		_w27291_
	);
	LUT2 #(
		.INIT('h1)
	) name16780 (
		_w27147_,
		_w27148_,
		_w27292_
	);
	LUT2 #(
		.INIT('h1)
	) name16781 (
		_w27149_,
		_w27150_,
		_w27293_
	);
	LUT2 #(
		.INIT('h1)
	) name16782 (
		_w27151_,
		_w27152_,
		_w27294_
	);
	LUT2 #(
		.INIT('h1)
	) name16783 (
		_w27153_,
		_w27154_,
		_w27295_
	);
	LUT2 #(
		.INIT('h1)
	) name16784 (
		_w27155_,
		_w27156_,
		_w27296_
	);
	LUT2 #(
		.INIT('h1)
	) name16785 (
		_w27157_,
		_w27158_,
		_w27297_
	);
	LUT2 #(
		.INIT('h1)
	) name16786 (
		_w27159_,
		_w27160_,
		_w27298_
	);
	LUT2 #(
		.INIT('h1)
	) name16787 (
		_w27161_,
		_w27162_,
		_w27299_
	);
	LUT2 #(
		.INIT('h1)
	) name16788 (
		_w27163_,
		_w27164_,
		_w27300_
	);
	LUT2 #(
		.INIT('h1)
	) name16789 (
		_w27165_,
		_w27166_,
		_w27301_
	);
	LUT2 #(
		.INIT('h1)
	) name16790 (
		_w27167_,
		_w27168_,
		_w27302_
	);
	LUT2 #(
		.INIT('h1)
	) name16791 (
		_w27169_,
		_w27170_,
		_w27303_
	);
	LUT2 #(
		.INIT('h1)
	) name16792 (
		_w27171_,
		_w27172_,
		_w27304_
	);
	LUT2 #(
		.INIT('h1)
	) name16793 (
		_w27173_,
		_w27174_,
		_w27305_
	);
	LUT2 #(
		.INIT('h1)
	) name16794 (
		_w27175_,
		_w27176_,
		_w27306_
	);
	LUT2 #(
		.INIT('h1)
	) name16795 (
		_w27177_,
		_w27178_,
		_w27307_
	);
	LUT2 #(
		.INIT('h1)
	) name16796 (
		_w27179_,
		_w27180_,
		_w27308_
	);
	LUT2 #(
		.INIT('h8)
	) name16797 (
		_w27307_,
		_w27308_,
		_w27309_
	);
	LUT2 #(
		.INIT('h8)
	) name16798 (
		_w27305_,
		_w27306_,
		_w27310_
	);
	LUT2 #(
		.INIT('h8)
	) name16799 (
		_w27303_,
		_w27304_,
		_w27311_
	);
	LUT2 #(
		.INIT('h8)
	) name16800 (
		_w27301_,
		_w27302_,
		_w27312_
	);
	LUT2 #(
		.INIT('h8)
	) name16801 (
		_w27299_,
		_w27300_,
		_w27313_
	);
	LUT2 #(
		.INIT('h8)
	) name16802 (
		_w27297_,
		_w27298_,
		_w27314_
	);
	LUT2 #(
		.INIT('h8)
	) name16803 (
		_w27295_,
		_w27296_,
		_w27315_
	);
	LUT2 #(
		.INIT('h8)
	) name16804 (
		_w27293_,
		_w27294_,
		_w27316_
	);
	LUT2 #(
		.INIT('h8)
	) name16805 (
		_w27291_,
		_w27292_,
		_w27317_
	);
	LUT2 #(
		.INIT('h8)
	) name16806 (
		_w27289_,
		_w27290_,
		_w27318_
	);
	LUT2 #(
		.INIT('h8)
	) name16807 (
		_w27287_,
		_w27288_,
		_w27319_
	);
	LUT2 #(
		.INIT('h8)
	) name16808 (
		_w27285_,
		_w27286_,
		_w27320_
	);
	LUT2 #(
		.INIT('h8)
	) name16809 (
		_w27283_,
		_w27284_,
		_w27321_
	);
	LUT2 #(
		.INIT('h8)
	) name16810 (
		_w27281_,
		_w27282_,
		_w27322_
	);
	LUT2 #(
		.INIT('h8)
	) name16811 (
		_w27279_,
		_w27280_,
		_w27323_
	);
	LUT2 #(
		.INIT('h8)
	) name16812 (
		_w27277_,
		_w27278_,
		_w27324_
	);
	LUT2 #(
		.INIT('h8)
	) name16813 (
		_w27275_,
		_w27276_,
		_w27325_
	);
	LUT2 #(
		.INIT('h8)
	) name16814 (
		_w27273_,
		_w27274_,
		_w27326_
	);
	LUT2 #(
		.INIT('h8)
	) name16815 (
		_w27271_,
		_w27272_,
		_w27327_
	);
	LUT2 #(
		.INIT('h8)
	) name16816 (
		_w27269_,
		_w27270_,
		_w27328_
	);
	LUT2 #(
		.INIT('h8)
	) name16817 (
		_w27267_,
		_w27268_,
		_w27329_
	);
	LUT2 #(
		.INIT('h8)
	) name16818 (
		_w27265_,
		_w27266_,
		_w27330_
	);
	LUT2 #(
		.INIT('h8)
	) name16819 (
		_w27263_,
		_w27264_,
		_w27331_
	);
	LUT2 #(
		.INIT('h8)
	) name16820 (
		_w27261_,
		_w27262_,
		_w27332_
	);
	LUT2 #(
		.INIT('h8)
	) name16821 (
		_w27259_,
		_w27260_,
		_w27333_
	);
	LUT2 #(
		.INIT('h8)
	) name16822 (
		_w27257_,
		_w27258_,
		_w27334_
	);
	LUT2 #(
		.INIT('h8)
	) name16823 (
		_w27255_,
		_w27256_,
		_w27335_
	);
	LUT2 #(
		.INIT('h8)
	) name16824 (
		_w27253_,
		_w27254_,
		_w27336_
	);
	LUT2 #(
		.INIT('h8)
	) name16825 (
		_w27251_,
		_w27252_,
		_w27337_
	);
	LUT2 #(
		.INIT('h8)
	) name16826 (
		_w27249_,
		_w27250_,
		_w27338_
	);
	LUT2 #(
		.INIT('h8)
	) name16827 (
		_w27247_,
		_w27248_,
		_w27339_
	);
	LUT2 #(
		.INIT('h8)
	) name16828 (
		_w27245_,
		_w27246_,
		_w27340_
	);
	LUT2 #(
		.INIT('h8)
	) name16829 (
		_w27243_,
		_w27244_,
		_w27341_
	);
	LUT2 #(
		.INIT('h8)
	) name16830 (
		_w27241_,
		_w27242_,
		_w27342_
	);
	LUT2 #(
		.INIT('h8)
	) name16831 (
		_w27239_,
		_w27240_,
		_w27343_
	);
	LUT2 #(
		.INIT('h8)
	) name16832 (
		_w27237_,
		_w27238_,
		_w27344_
	);
	LUT2 #(
		.INIT('h8)
	) name16833 (
		_w27235_,
		_w27236_,
		_w27345_
	);
	LUT2 #(
		.INIT('h8)
	) name16834 (
		_w27233_,
		_w27234_,
		_w27346_
	);
	LUT2 #(
		.INIT('h8)
	) name16835 (
		_w27231_,
		_w27232_,
		_w27347_
	);
	LUT2 #(
		.INIT('h8)
	) name16836 (
		_w27229_,
		_w27230_,
		_w27348_
	);
	LUT2 #(
		.INIT('h8)
	) name16837 (
		_w27227_,
		_w27228_,
		_w27349_
	);
	LUT2 #(
		.INIT('h8)
	) name16838 (
		_w27225_,
		_w27226_,
		_w27350_
	);
	LUT2 #(
		.INIT('h8)
	) name16839 (
		_w27223_,
		_w27224_,
		_w27351_
	);
	LUT2 #(
		.INIT('h8)
	) name16840 (
		_w27221_,
		_w27222_,
		_w27352_
	);
	LUT2 #(
		.INIT('h8)
	) name16841 (
		_w27219_,
		_w27220_,
		_w27353_
	);
	LUT2 #(
		.INIT('h8)
	) name16842 (
		_w27217_,
		_w27218_,
		_w27354_
	);
	LUT2 #(
		.INIT('h8)
	) name16843 (
		_w27215_,
		_w27216_,
		_w27355_
	);
	LUT2 #(
		.INIT('h8)
	) name16844 (
		_w27213_,
		_w27214_,
		_w27356_
	);
	LUT2 #(
		.INIT('h8)
	) name16845 (
		_w27211_,
		_w27212_,
		_w27357_
	);
	LUT2 #(
		.INIT('h8)
	) name16846 (
		_w27209_,
		_w27210_,
		_w27358_
	);
	LUT2 #(
		.INIT('h8)
	) name16847 (
		_w27207_,
		_w27208_,
		_w27359_
	);
	LUT2 #(
		.INIT('h8)
	) name16848 (
		_w27205_,
		_w27206_,
		_w27360_
	);
	LUT2 #(
		.INIT('h8)
	) name16849 (
		_w27203_,
		_w27204_,
		_w27361_
	);
	LUT2 #(
		.INIT('h8)
	) name16850 (
		_w27201_,
		_w27202_,
		_w27362_
	);
	LUT2 #(
		.INIT('h8)
	) name16851 (
		_w27199_,
		_w27200_,
		_w27363_
	);
	LUT2 #(
		.INIT('h8)
	) name16852 (
		_w27197_,
		_w27198_,
		_w27364_
	);
	LUT2 #(
		.INIT('h8)
	) name16853 (
		_w27195_,
		_w27196_,
		_w27365_
	);
	LUT2 #(
		.INIT('h8)
	) name16854 (
		_w27193_,
		_w27194_,
		_w27366_
	);
	LUT2 #(
		.INIT('h8)
	) name16855 (
		_w27191_,
		_w27192_,
		_w27367_
	);
	LUT2 #(
		.INIT('h8)
	) name16856 (
		_w27189_,
		_w27190_,
		_w27368_
	);
	LUT2 #(
		.INIT('h8)
	) name16857 (
		_w27187_,
		_w27188_,
		_w27369_
	);
	LUT2 #(
		.INIT('h8)
	) name16858 (
		_w27185_,
		_w27186_,
		_w27370_
	);
	LUT2 #(
		.INIT('h8)
	) name16859 (
		_w27183_,
		_w27184_,
		_w27371_
	);
	LUT2 #(
		.INIT('h8)
	) name16860 (
		_w27181_,
		_w27182_,
		_w27372_
	);
	LUT2 #(
		.INIT('h8)
	) name16861 (
		_w27371_,
		_w27372_,
		_w27373_
	);
	LUT2 #(
		.INIT('h8)
	) name16862 (
		_w27369_,
		_w27370_,
		_w27374_
	);
	LUT2 #(
		.INIT('h8)
	) name16863 (
		_w27367_,
		_w27368_,
		_w27375_
	);
	LUT2 #(
		.INIT('h8)
	) name16864 (
		_w27365_,
		_w27366_,
		_w27376_
	);
	LUT2 #(
		.INIT('h8)
	) name16865 (
		_w27363_,
		_w27364_,
		_w27377_
	);
	LUT2 #(
		.INIT('h8)
	) name16866 (
		_w27361_,
		_w27362_,
		_w27378_
	);
	LUT2 #(
		.INIT('h8)
	) name16867 (
		_w27359_,
		_w27360_,
		_w27379_
	);
	LUT2 #(
		.INIT('h8)
	) name16868 (
		_w27357_,
		_w27358_,
		_w27380_
	);
	LUT2 #(
		.INIT('h8)
	) name16869 (
		_w27355_,
		_w27356_,
		_w27381_
	);
	LUT2 #(
		.INIT('h8)
	) name16870 (
		_w27353_,
		_w27354_,
		_w27382_
	);
	LUT2 #(
		.INIT('h8)
	) name16871 (
		_w27351_,
		_w27352_,
		_w27383_
	);
	LUT2 #(
		.INIT('h8)
	) name16872 (
		_w27349_,
		_w27350_,
		_w27384_
	);
	LUT2 #(
		.INIT('h8)
	) name16873 (
		_w27347_,
		_w27348_,
		_w27385_
	);
	LUT2 #(
		.INIT('h8)
	) name16874 (
		_w27345_,
		_w27346_,
		_w27386_
	);
	LUT2 #(
		.INIT('h8)
	) name16875 (
		_w27343_,
		_w27344_,
		_w27387_
	);
	LUT2 #(
		.INIT('h8)
	) name16876 (
		_w27341_,
		_w27342_,
		_w27388_
	);
	LUT2 #(
		.INIT('h8)
	) name16877 (
		_w27339_,
		_w27340_,
		_w27389_
	);
	LUT2 #(
		.INIT('h8)
	) name16878 (
		_w27337_,
		_w27338_,
		_w27390_
	);
	LUT2 #(
		.INIT('h8)
	) name16879 (
		_w27335_,
		_w27336_,
		_w27391_
	);
	LUT2 #(
		.INIT('h8)
	) name16880 (
		_w27333_,
		_w27334_,
		_w27392_
	);
	LUT2 #(
		.INIT('h8)
	) name16881 (
		_w27331_,
		_w27332_,
		_w27393_
	);
	LUT2 #(
		.INIT('h8)
	) name16882 (
		_w27329_,
		_w27330_,
		_w27394_
	);
	LUT2 #(
		.INIT('h8)
	) name16883 (
		_w27327_,
		_w27328_,
		_w27395_
	);
	LUT2 #(
		.INIT('h8)
	) name16884 (
		_w27325_,
		_w27326_,
		_w27396_
	);
	LUT2 #(
		.INIT('h8)
	) name16885 (
		_w27323_,
		_w27324_,
		_w27397_
	);
	LUT2 #(
		.INIT('h8)
	) name16886 (
		_w27321_,
		_w27322_,
		_w27398_
	);
	LUT2 #(
		.INIT('h8)
	) name16887 (
		_w27319_,
		_w27320_,
		_w27399_
	);
	LUT2 #(
		.INIT('h8)
	) name16888 (
		_w27317_,
		_w27318_,
		_w27400_
	);
	LUT2 #(
		.INIT('h8)
	) name16889 (
		_w27315_,
		_w27316_,
		_w27401_
	);
	LUT2 #(
		.INIT('h8)
	) name16890 (
		_w27313_,
		_w27314_,
		_w27402_
	);
	LUT2 #(
		.INIT('h8)
	) name16891 (
		_w27311_,
		_w27312_,
		_w27403_
	);
	LUT2 #(
		.INIT('h8)
	) name16892 (
		_w27309_,
		_w27310_,
		_w27404_
	);
	LUT2 #(
		.INIT('h8)
	) name16893 (
		_w27403_,
		_w27404_,
		_w27405_
	);
	LUT2 #(
		.INIT('h8)
	) name16894 (
		_w27401_,
		_w27402_,
		_w27406_
	);
	LUT2 #(
		.INIT('h8)
	) name16895 (
		_w27399_,
		_w27400_,
		_w27407_
	);
	LUT2 #(
		.INIT('h8)
	) name16896 (
		_w27397_,
		_w27398_,
		_w27408_
	);
	LUT2 #(
		.INIT('h8)
	) name16897 (
		_w27395_,
		_w27396_,
		_w27409_
	);
	LUT2 #(
		.INIT('h8)
	) name16898 (
		_w27393_,
		_w27394_,
		_w27410_
	);
	LUT2 #(
		.INIT('h8)
	) name16899 (
		_w27391_,
		_w27392_,
		_w27411_
	);
	LUT2 #(
		.INIT('h8)
	) name16900 (
		_w27389_,
		_w27390_,
		_w27412_
	);
	LUT2 #(
		.INIT('h8)
	) name16901 (
		_w27387_,
		_w27388_,
		_w27413_
	);
	LUT2 #(
		.INIT('h8)
	) name16902 (
		_w27385_,
		_w27386_,
		_w27414_
	);
	LUT2 #(
		.INIT('h8)
	) name16903 (
		_w27383_,
		_w27384_,
		_w27415_
	);
	LUT2 #(
		.INIT('h8)
	) name16904 (
		_w27381_,
		_w27382_,
		_w27416_
	);
	LUT2 #(
		.INIT('h8)
	) name16905 (
		_w27379_,
		_w27380_,
		_w27417_
	);
	LUT2 #(
		.INIT('h8)
	) name16906 (
		_w27377_,
		_w27378_,
		_w27418_
	);
	LUT2 #(
		.INIT('h8)
	) name16907 (
		_w27375_,
		_w27376_,
		_w27419_
	);
	LUT2 #(
		.INIT('h8)
	) name16908 (
		_w27373_,
		_w27374_,
		_w27420_
	);
	LUT2 #(
		.INIT('h8)
	) name16909 (
		_w27419_,
		_w27420_,
		_w27421_
	);
	LUT2 #(
		.INIT('h8)
	) name16910 (
		_w27417_,
		_w27418_,
		_w27422_
	);
	LUT2 #(
		.INIT('h8)
	) name16911 (
		_w27415_,
		_w27416_,
		_w27423_
	);
	LUT2 #(
		.INIT('h8)
	) name16912 (
		_w27413_,
		_w27414_,
		_w27424_
	);
	LUT2 #(
		.INIT('h8)
	) name16913 (
		_w27411_,
		_w27412_,
		_w27425_
	);
	LUT2 #(
		.INIT('h8)
	) name16914 (
		_w27409_,
		_w27410_,
		_w27426_
	);
	LUT2 #(
		.INIT('h8)
	) name16915 (
		_w27407_,
		_w27408_,
		_w27427_
	);
	LUT2 #(
		.INIT('h8)
	) name16916 (
		_w27405_,
		_w27406_,
		_w27428_
	);
	LUT2 #(
		.INIT('h8)
	) name16917 (
		_w27427_,
		_w27428_,
		_w27429_
	);
	LUT2 #(
		.INIT('h8)
	) name16918 (
		_w27425_,
		_w27426_,
		_w27430_
	);
	LUT2 #(
		.INIT('h8)
	) name16919 (
		_w27423_,
		_w27424_,
		_w27431_
	);
	LUT2 #(
		.INIT('h8)
	) name16920 (
		_w27421_,
		_w27422_,
		_w27432_
	);
	LUT2 #(
		.INIT('h8)
	) name16921 (
		_w27431_,
		_w27432_,
		_w27433_
	);
	LUT2 #(
		.INIT('h8)
	) name16922 (
		_w27429_,
		_w27430_,
		_w27434_
	);
	LUT2 #(
		.INIT('h8)
	) name16923 (
		_w27433_,
		_w27434_,
		_w27435_
	);
	LUT2 #(
		.INIT('h1)
	) name16924 (
		wb_rst_i_pad,
		_w27435_,
		_w27436_
	);
	LUT2 #(
		.INIT('h1)
	) name16925 (
		_w22944_,
		_w27436_,
		_w27437_
	);
	LUT2 #(
		.INIT('h8)
	) name16926 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		_w22959_,
		_w27438_
	);
	LUT2 #(
		.INIT('h8)
	) name16927 (
		\ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 ,
		_w23499_,
		_w27439_
	);
	LUT2 #(
		.INIT('h8)
	) name16928 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		_w23501_,
		_w27440_
	);
	LUT2 #(
		.INIT('h8)
	) name16929 (
		\ethreg1_MIIRX_DATA_DataOut_reg[9]/NET0131 ,
		_w23507_,
		_w27441_
	);
	LUT2 #(
		.INIT('h8)
	) name16930 (
		\ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 ,
		_w22952_,
		_w27442_
	);
	LUT2 #(
		.INIT('h8)
	) name16931 (
		\ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 ,
		_w22956_,
		_w27443_
	);
	LUT2 #(
		.INIT('h8)
	) name16932 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w23513_,
		_w27444_
	);
	LUT2 #(
		.INIT('h8)
	) name16933 (
		\ethreg1_PACKETLEN_1_DataOut_reg[1]/NET0131 ,
		_w22966_,
		_w27445_
	);
	LUT2 #(
		.INIT('h8)
	) name16934 (
		\ethreg1_MODER_1_DataOut_reg[1]/NET0131 ,
		_w23519_,
		_w27446_
	);
	LUT2 #(
		.INIT('h8)
	) name16935 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 ,
		_w23522_,
		_w27447_
	);
	LUT2 #(
		.INIT('h1)
	) name16936 (
		_w27438_,
		_w27439_,
		_w27448_
	);
	LUT2 #(
		.INIT('h1)
	) name16937 (
		_w27440_,
		_w27441_,
		_w27449_
	);
	LUT2 #(
		.INIT('h1)
	) name16938 (
		_w27442_,
		_w27443_,
		_w27450_
	);
	LUT2 #(
		.INIT('h1)
	) name16939 (
		_w27444_,
		_w27446_,
		_w27451_
	);
	LUT2 #(
		.INIT('h4)
	) name16940 (
		_w27447_,
		_w27451_,
		_w27452_
	);
	LUT2 #(
		.INIT('h8)
	) name16941 (
		_w27449_,
		_w27450_,
		_w27453_
	);
	LUT2 #(
		.INIT('h8)
	) name16942 (
		_w22944_,
		_w27448_,
		_w27454_
	);
	LUT2 #(
		.INIT('h8)
	) name16943 (
		_w27453_,
		_w27454_,
		_w27455_
	);
	LUT2 #(
		.INIT('h4)
	) name16944 (
		_w27445_,
		_w27452_,
		_w27456_
	);
	LUT2 #(
		.INIT('h8)
	) name16945 (
		_w27455_,
		_w27456_,
		_w27457_
	);
	LUT2 #(
		.INIT('h1)
	) name16946 (
		_w27437_,
		_w27457_,
		_w27458_
	);
	LUT2 #(
		.INIT('h1)
	) name16947 (
		_w16743_,
		_w22944_,
		_w27459_
	);
	LUT2 #(
		.INIT('h8)
	) name16948 (
		\ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 ,
		_w22952_,
		_w27460_
	);
	LUT2 #(
		.INIT('h8)
	) name16949 (
		\ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 ,
		_w22956_,
		_w27461_
	);
	LUT2 #(
		.INIT('h8)
	) name16950 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		_w22959_,
		_w27462_
	);
	LUT2 #(
		.INIT('h8)
	) name16951 (
		\ethreg1_PACKETLEN_2_DataOut_reg[4]/NET0131 ,
		_w22966_,
		_w27463_
	);
	LUT2 #(
		.INIT('h1)
	) name16952 (
		_w27460_,
		_w27461_,
		_w27464_
	);
	LUT2 #(
		.INIT('h4)
	) name16953 (
		_w27462_,
		_w27464_,
		_w27465_
	);
	LUT2 #(
		.INIT('h8)
	) name16954 (
		_w22944_,
		_w27465_,
		_w27466_
	);
	LUT2 #(
		.INIT('h4)
	) name16955 (
		_w27463_,
		_w27466_,
		_w27467_
	);
	LUT2 #(
		.INIT('h1)
	) name16956 (
		_w27459_,
		_w27467_,
		_w27468_
	);
	LUT2 #(
		.INIT('h8)
	) name16957 (
		\wishbone_bd_ram_mem1_reg[69][11]/P0001 ,
		_w12738_,
		_w27469_
	);
	LUT2 #(
		.INIT('h8)
	) name16958 (
		\wishbone_bd_ram_mem1_reg[157][11]/P0001 ,
		_w12926_,
		_w27470_
	);
	LUT2 #(
		.INIT('h8)
	) name16959 (
		\wishbone_bd_ram_mem1_reg[106][11]/P0001 ,
		_w12713_,
		_w27471_
	);
	LUT2 #(
		.INIT('h8)
	) name16960 (
		\wishbone_bd_ram_mem1_reg[177][11]/P0001 ,
		_w12996_,
		_w27472_
	);
	LUT2 #(
		.INIT('h8)
	) name16961 (
		\wishbone_bd_ram_mem1_reg[64][11]/P0001 ,
		_w12976_,
		_w27473_
	);
	LUT2 #(
		.INIT('h8)
	) name16962 (
		\wishbone_bd_ram_mem1_reg[95][11]/P0001 ,
		_w12844_,
		_w27474_
	);
	LUT2 #(
		.INIT('h8)
	) name16963 (
		\wishbone_bd_ram_mem1_reg[68][11]/P0001 ,
		_w12946_,
		_w27475_
	);
	LUT2 #(
		.INIT('h8)
	) name16964 (
		\wishbone_bd_ram_mem1_reg[46][11]/P0001 ,
		_w12884_,
		_w27476_
	);
	LUT2 #(
		.INIT('h8)
	) name16965 (
		\wishbone_bd_ram_mem1_reg[118][11]/P0001 ,
		_w12830_,
		_w27477_
	);
	LUT2 #(
		.INIT('h8)
	) name16966 (
		\wishbone_bd_ram_mem1_reg[28][11]/P0001 ,
		_w13170_,
		_w27478_
	);
	LUT2 #(
		.INIT('h8)
	) name16967 (
		\wishbone_bd_ram_mem1_reg[171][11]/P0001 ,
		_w12910_,
		_w27479_
	);
	LUT2 #(
		.INIT('h8)
	) name16968 (
		\wishbone_bd_ram_mem1_reg[163][11]/P0001 ,
		_w12882_,
		_w27480_
	);
	LUT2 #(
		.INIT('h8)
	) name16969 (
		\wishbone_bd_ram_mem1_reg[27][11]/P0001 ,
		_w12880_,
		_w27481_
	);
	LUT2 #(
		.INIT('h8)
	) name16970 (
		\wishbone_bd_ram_mem1_reg[190][11]/P0001 ,
		_w12858_,
		_w27482_
	);
	LUT2 #(
		.INIT('h8)
	) name16971 (
		\wishbone_bd_ram_mem1_reg[107][11]/P0001 ,
		_w12749_,
		_w27483_
	);
	LUT2 #(
		.INIT('h8)
	) name16972 (
		\wishbone_bd_ram_mem1_reg[36][11]/P0001 ,
		_w12800_,
		_w27484_
	);
	LUT2 #(
		.INIT('h8)
	) name16973 (
		\wishbone_bd_ram_mem1_reg[182][11]/P0001 ,
		_w12820_,
		_w27485_
	);
	LUT2 #(
		.INIT('h8)
	) name16974 (
		\wishbone_bd_ram_mem1_reg[74][11]/P0001 ,
		_w12812_,
		_w27486_
	);
	LUT2 #(
		.INIT('h8)
	) name16975 (
		\wishbone_bd_ram_mem1_reg[131][11]/P0001 ,
		_w12852_,
		_w27487_
	);
	LUT2 #(
		.INIT('h8)
	) name16976 (
		\wishbone_bd_ram_mem1_reg[38][11]/P0001 ,
		_w13182_,
		_w27488_
	);
	LUT2 #(
		.INIT('h8)
	) name16977 (
		\wishbone_bd_ram_mem1_reg[121][11]/P0001 ,
		_w13078_,
		_w27489_
	);
	LUT2 #(
		.INIT('h8)
	) name16978 (
		\wishbone_bd_ram_mem1_reg[176][11]/P0001 ,
		_w12868_,
		_w27490_
	);
	LUT2 #(
		.INIT('h8)
	) name16979 (
		\wishbone_bd_ram_mem1_reg[242][11]/P0001 ,
		_w12932_,
		_w27491_
	);
	LUT2 #(
		.INIT('h8)
	) name16980 (
		\wishbone_bd_ram_mem1_reg[79][11]/P0001 ,
		_w13212_,
		_w27492_
	);
	LUT2 #(
		.INIT('h8)
	) name16981 (
		\wishbone_bd_ram_mem1_reg[245][11]/P0001 ,
		_w13022_,
		_w27493_
	);
	LUT2 #(
		.INIT('h8)
	) name16982 (
		\wishbone_bd_ram_mem1_reg[56][11]/P0001 ,
		_w12778_,
		_w27494_
	);
	LUT2 #(
		.INIT('h8)
	) name16983 (
		\wishbone_bd_ram_mem1_reg[183][11]/P0001 ,
		_w12787_,
		_w27495_
	);
	LUT2 #(
		.INIT('h8)
	) name16984 (
		\wishbone_bd_ram_mem1_reg[124][11]/P0001 ,
		_w13058_,
		_w27496_
	);
	LUT2 #(
		.INIT('h8)
	) name16985 (
		\wishbone_bd_ram_mem1_reg[221][11]/P0001 ,
		_w12802_,
		_w27497_
	);
	LUT2 #(
		.INIT('h8)
	) name16986 (
		\wishbone_bd_ram_mem1_reg[218][11]/P0001 ,
		_w13206_,
		_w27498_
	);
	LUT2 #(
		.INIT('h8)
	) name16987 (
		\wishbone_bd_ram_mem1_reg[162][11]/P0001 ,
		_w13098_,
		_w27499_
	);
	LUT2 #(
		.INIT('h8)
	) name16988 (
		\wishbone_bd_ram_mem1_reg[21][11]/P0001 ,
		_w12906_,
		_w27500_
	);
	LUT2 #(
		.INIT('h8)
	) name16989 (
		\wishbone_bd_ram_mem1_reg[123][11]/P0001 ,
		_w13114_,
		_w27501_
	);
	LUT2 #(
		.INIT('h8)
	) name16990 (
		\wishbone_bd_ram_mem1_reg[217][11]/P0001 ,
		_w13188_,
		_w27502_
	);
	LUT2 #(
		.INIT('h8)
	) name16991 (
		\wishbone_bd_ram_mem1_reg[250][11]/P0001 ,
		_w13128_,
		_w27503_
	);
	LUT2 #(
		.INIT('h8)
	) name16992 (
		\wishbone_bd_ram_mem1_reg[154][11]/P0001 ,
		_w12962_,
		_w27504_
	);
	LUT2 #(
		.INIT('h8)
	) name16993 (
		\wishbone_bd_ram_mem1_reg[62][11]/P0001 ,
		_w12673_,
		_w27505_
	);
	LUT2 #(
		.INIT('h8)
	) name16994 (
		\wishbone_bd_ram_mem1_reg[134][11]/P0001 ,
		_w12763_,
		_w27506_
	);
	LUT2 #(
		.INIT('h8)
	) name16995 (
		\wishbone_bd_ram_mem1_reg[184][11]/P0001 ,
		_w13062_,
		_w27507_
	);
	LUT2 #(
		.INIT('h8)
	) name16996 (
		\wishbone_bd_ram_mem1_reg[219][11]/P0001 ,
		_w12806_,
		_w27508_
	);
	LUT2 #(
		.INIT('h8)
	) name16997 (
		\wishbone_bd_ram_mem1_reg[33][11]/P0001 ,
		_w12980_,
		_w27509_
	);
	LUT2 #(
		.INIT('h8)
	) name16998 (
		\wishbone_bd_ram_mem1_reg[253][11]/P0001 ,
		_w13100_,
		_w27510_
	);
	LUT2 #(
		.INIT('h8)
	) name16999 (
		\wishbone_bd_ram_mem1_reg[113][11]/P0001 ,
		_w13026_,
		_w27511_
	);
	LUT2 #(
		.INIT('h8)
	) name17000 (
		\wishbone_bd_ram_mem1_reg[153][11]/P0001 ,
		_w12890_,
		_w27512_
	);
	LUT2 #(
		.INIT('h8)
	) name17001 (
		\wishbone_bd_ram_mem1_reg[185][11]/P0001 ,
		_w12940_,
		_w27513_
	);
	LUT2 #(
		.INIT('h8)
	) name17002 (
		\wishbone_bd_ram_mem1_reg[232][11]/P0001 ,
		_w12758_,
		_w27514_
	);
	LUT2 #(
		.INIT('h8)
	) name17003 (
		\wishbone_bd_ram_mem1_reg[55][11]/P0001 ,
		_w12785_,
		_w27515_
	);
	LUT2 #(
		.INIT('h8)
	) name17004 (
		\wishbone_bd_ram_mem1_reg[101][11]/P0001 ,
		_w13192_,
		_w27516_
	);
	LUT2 #(
		.INIT('h8)
	) name17005 (
		\wishbone_bd_ram_mem1_reg[8][11]/P0001 ,
		_w12920_,
		_w27517_
	);
	LUT2 #(
		.INIT('h8)
	) name17006 (
		\wishbone_bd_ram_mem1_reg[234][11]/P0001 ,
		_w13214_,
		_w27518_
	);
	LUT2 #(
		.INIT('h8)
	) name17007 (
		\wishbone_bd_ram_mem1_reg[148][11]/P0001 ,
		_w13000_,
		_w27519_
	);
	LUT2 #(
		.INIT('h8)
	) name17008 (
		\wishbone_bd_ram_mem1_reg[98][11]/P0001 ,
		_w12816_,
		_w27520_
	);
	LUT2 #(
		.INIT('h8)
	) name17009 (
		\wishbone_bd_ram_mem1_reg[246][11]/P0001 ,
		_w13076_,
		_w27521_
	);
	LUT2 #(
		.INIT('h8)
	) name17010 (
		\wishbone_bd_ram_mem1_reg[122][11]/P0001 ,
		_w13130_,
		_w27522_
	);
	LUT2 #(
		.INIT('h8)
	) name17011 (
		\wishbone_bd_ram_mem1_reg[174][11]/P0001 ,
		_w12972_,
		_w27523_
	);
	LUT2 #(
		.INIT('h8)
	) name17012 (
		\wishbone_bd_ram_mem1_reg[180][11]/P0001 ,
		_w12791_,
		_w27524_
	);
	LUT2 #(
		.INIT('h8)
	) name17013 (
		\wishbone_bd_ram_mem1_reg[90][11]/P0001 ,
		_w12978_,
		_w27525_
	);
	LUT2 #(
		.INIT('h8)
	) name17014 (
		\wishbone_bd_ram_mem1_reg[206][11]/P0001 ,
		_w12954_,
		_w27526_
	);
	LUT2 #(
		.INIT('h8)
	) name17015 (
		\wishbone_bd_ram_mem1_reg[82][11]/P0001 ,
		_w12942_,
		_w27527_
	);
	LUT2 #(
		.INIT('h8)
	) name17016 (
		\wishbone_bd_ram_mem1_reg[111][11]/P0001 ,
		_w12744_,
		_w27528_
	);
	LUT2 #(
		.INIT('h8)
	) name17017 (
		\wishbone_bd_ram_mem1_reg[222][11]/P0001 ,
		_w13094_,
		_w27529_
	);
	LUT2 #(
		.INIT('h8)
	) name17018 (
		\wishbone_bd_ram_mem1_reg[191][11]/P0001 ,
		_w13034_,
		_w27530_
	);
	LUT2 #(
		.INIT('h8)
	) name17019 (
		\wishbone_bd_ram_mem1_reg[99][11]/P0001 ,
		_w13038_,
		_w27531_
	);
	LUT2 #(
		.INIT('h8)
	) name17020 (
		\wishbone_bd_ram_mem1_reg[192][11]/P0001 ,
		_w12938_,
		_w27532_
	);
	LUT2 #(
		.INIT('h8)
	) name17021 (
		\wishbone_bd_ram_mem1_reg[48][11]/P0001 ,
		_w12970_,
		_w27533_
	);
	LUT2 #(
		.INIT('h8)
	) name17022 (
		\wishbone_bd_ram_mem1_reg[231][11]/P0001 ,
		_w12856_,
		_w27534_
	);
	LUT2 #(
		.INIT('h8)
	) name17023 (
		\wishbone_bd_ram_mem1_reg[136][11]/P0001 ,
		_w13064_,
		_w27535_
	);
	LUT2 #(
		.INIT('h8)
	) name17024 (
		\wishbone_bd_ram_mem1_reg[127][11]/P0001 ,
		_w13164_,
		_w27536_
	);
	LUT2 #(
		.INIT('h8)
	) name17025 (
		\wishbone_bd_ram_mem1_reg[161][11]/P0001 ,
		_w12754_,
		_w27537_
	);
	LUT2 #(
		.INIT('h8)
	) name17026 (
		\wishbone_bd_ram_mem1_reg[224][11]/P0001 ,
		_w12902_,
		_w27538_
	);
	LUT2 #(
		.INIT('h8)
	) name17027 (
		\wishbone_bd_ram_mem1_reg[146][11]/P0001 ,
		_w13060_,
		_w27539_
	);
	LUT2 #(
		.INIT('h8)
	) name17028 (
		\wishbone_bd_ram_mem1_reg[168][11]/P0001 ,
		_w13208_,
		_w27540_
	);
	LUT2 #(
		.INIT('h8)
	) name17029 (
		\wishbone_bd_ram_mem1_reg[65][11]/P0001 ,
		_w13176_,
		_w27541_
	);
	LUT2 #(
		.INIT('h8)
	) name17030 (
		\wishbone_bd_ram_mem1_reg[197][11]/P0001 ,
		_w12834_,
		_w27542_
	);
	LUT2 #(
		.INIT('h8)
	) name17031 (
		\wishbone_bd_ram_mem1_reg[125][11]/P0001 ,
		_w12956_,
		_w27543_
	);
	LUT2 #(
		.INIT('h8)
	) name17032 (
		\wishbone_bd_ram_mem1_reg[202][11]/P0001 ,
		_w12870_,
		_w27544_
	);
	LUT2 #(
		.INIT('h8)
	) name17033 (
		\wishbone_bd_ram_mem1_reg[189][11]/P0001 ,
		_w13042_,
		_w27545_
	);
	LUT2 #(
		.INIT('h8)
	) name17034 (
		\wishbone_bd_ram_mem1_reg[237][11]/P0001 ,
		_w12990_,
		_w27546_
	);
	LUT2 #(
		.INIT('h8)
	) name17035 (
		\wishbone_bd_ram_mem1_reg[213][11]/P0001 ,
		_w13002_,
		_w27547_
	);
	LUT2 #(
		.INIT('h8)
	) name17036 (
		\wishbone_bd_ram_mem1_reg[42][11]/P0001 ,
		_w12842_,
		_w27548_
	);
	LUT2 #(
		.INIT('h8)
	) name17037 (
		\wishbone_bd_ram_mem1_reg[31][11]/P0001 ,
		_w13198_,
		_w27549_
	);
	LUT2 #(
		.INIT('h8)
	) name17038 (
		\wishbone_bd_ram_mem1_reg[142][11]/P0001 ,
		_w12928_,
		_w27550_
	);
	LUT2 #(
		.INIT('h8)
	) name17039 (
		\wishbone_bd_ram_mem1_reg[58][11]/P0001 ,
		_w13070_,
		_w27551_
	);
	LUT2 #(
		.INIT('h8)
	) name17040 (
		\wishbone_bd_ram_mem1_reg[4][11]/P0001 ,
		_w12666_,
		_w27552_
	);
	LUT2 #(
		.INIT('h8)
	) name17041 (
		\wishbone_bd_ram_mem1_reg[16][11]/P0001 ,
		_w13140_,
		_w27553_
	);
	LUT2 #(
		.INIT('h8)
	) name17042 (
		\wishbone_bd_ram_mem1_reg[84][11]/P0001 ,
		_w12934_,
		_w27554_
	);
	LUT2 #(
		.INIT('h8)
	) name17043 (
		\wishbone_bd_ram_mem1_reg[18][11]/P0001 ,
		_w12679_,
		_w27555_
	);
	LUT2 #(
		.INIT('h8)
	) name17044 (
		\wishbone_bd_ram_mem1_reg[138][11]/P0001 ,
		_w12958_,
		_w27556_
	);
	LUT2 #(
		.INIT('h8)
	) name17045 (
		\wishbone_bd_ram_mem1_reg[110][11]/P0001 ,
		_w13046_,
		_w27557_
	);
	LUT2 #(
		.INIT('h8)
	) name17046 (
		\wishbone_bd_ram_mem1_reg[239][11]/P0001 ,
		_w12862_,
		_w27558_
	);
	LUT2 #(
		.INIT('h8)
	) name17047 (
		\wishbone_bd_ram_mem1_reg[178][11]/P0001 ,
		_w12886_,
		_w27559_
	);
	LUT2 #(
		.INIT('h8)
	) name17048 (
		\wishbone_bd_ram_mem1_reg[179][11]/P0001 ,
		_w13050_,
		_w27560_
	);
	LUT2 #(
		.INIT('h8)
	) name17049 (
		\wishbone_bd_ram_mem1_reg[210][11]/P0001 ,
		_w12924_,
		_w27561_
	);
	LUT2 #(
		.INIT('h8)
	) name17050 (
		\wishbone_bd_ram_mem1_reg[151][11]/P0001 ,
		_w13142_,
		_w27562_
	);
	LUT2 #(
		.INIT('h8)
	) name17051 (
		\wishbone_bd_ram_mem1_reg[80][11]/P0001 ,
		_w12689_,
		_w27563_
	);
	LUT2 #(
		.INIT('h8)
	) name17052 (
		\wishbone_bd_ram_mem1_reg[83][11]/P0001 ,
		_w12916_,
		_w27564_
	);
	LUT2 #(
		.INIT('h8)
	) name17053 (
		\wishbone_bd_ram_mem1_reg[214][11]/P0001 ,
		_w12984_,
		_w27565_
	);
	LUT2 #(
		.INIT('h8)
	) name17054 (
		\wishbone_bd_ram_mem1_reg[173][11]/P0001 ,
		_w12854_,
		_w27566_
	);
	LUT2 #(
		.INIT('h8)
	) name17055 (
		\wishbone_bd_ram_mem1_reg[20][11]/P0001 ,
		_w13174_,
		_w27567_
	);
	LUT2 #(
		.INIT('h8)
	) name17056 (
		\wishbone_bd_ram_mem1_reg[40][11]/P0001 ,
		_w13132_,
		_w27568_
	);
	LUT2 #(
		.INIT('h8)
	) name17057 (
		\wishbone_bd_ram_mem1_reg[91][11]/P0001 ,
		_w13074_,
		_w27569_
	);
	LUT2 #(
		.INIT('h8)
	) name17058 (
		\wishbone_bd_ram_mem1_reg[44][11]/P0001 ,
		_w12896_,
		_w27570_
	);
	LUT2 #(
		.INIT('h8)
	) name17059 (
		\wishbone_bd_ram_mem1_reg[30][11]/P0001 ,
		_w13104_,
		_w27571_
	);
	LUT2 #(
		.INIT('h8)
	) name17060 (
		\wishbone_bd_ram_mem1_reg[220][11]/P0001 ,
		_w13066_,
		_w27572_
	);
	LUT2 #(
		.INIT('h8)
	) name17061 (
		\wishbone_bd_ram_mem1_reg[75][11]/P0001 ,
		_w12826_,
		_w27573_
	);
	LUT2 #(
		.INIT('h8)
	) name17062 (
		\wishbone_bd_ram_mem1_reg[10][11]/P0001 ,
		_w13172_,
		_w27574_
	);
	LUT2 #(
		.INIT('h8)
	) name17063 (
		\wishbone_bd_ram_mem1_reg[12][11]/P0001 ,
		_w13118_,
		_w27575_
	);
	LUT2 #(
		.INIT('h8)
	) name17064 (
		\wishbone_bd_ram_mem1_reg[61][11]/P0001 ,
		_w12725_,
		_w27576_
	);
	LUT2 #(
		.INIT('h8)
	) name17065 (
		\wishbone_bd_ram_mem1_reg[181][11]/P0001 ,
		_w12828_,
		_w27577_
	);
	LUT2 #(
		.INIT('h8)
	) name17066 (
		\wishbone_bd_ram_mem1_reg[26][11]/P0001 ,
		_w12699_,
		_w27578_
	);
	LUT2 #(
		.INIT('h8)
	) name17067 (
		\wishbone_bd_ram_mem1_reg[147][11]/P0001 ,
		_w13146_,
		_w27579_
	);
	LUT2 #(
		.INIT('h8)
	) name17068 (
		\wishbone_bd_ram_mem1_reg[211][11]/P0001 ,
		_w13166_,
		_w27580_
	);
	LUT2 #(
		.INIT('h8)
	) name17069 (
		\wishbone_bd_ram_mem1_reg[164][11]/P0001 ,
		_w12876_,
		_w27581_
	);
	LUT2 #(
		.INIT('h8)
	) name17070 (
		\wishbone_bd_ram_mem1_reg[78][11]/P0001 ,
		_w12874_,
		_w27582_
	);
	LUT2 #(
		.INIT('h8)
	) name17071 (
		\wishbone_bd_ram_mem1_reg[35][11]/P0001 ,
		_w12703_,
		_w27583_
	);
	LUT2 #(
		.INIT('h8)
	) name17072 (
		\wishbone_bd_ram_mem1_reg[160][11]/P0001 ,
		_w12872_,
		_w27584_
	);
	LUT2 #(
		.INIT('h8)
	) name17073 (
		\wishbone_bd_ram_mem1_reg[175][11]/P0001 ,
		_w13126_,
		_w27585_
	);
	LUT2 #(
		.INIT('h8)
	) name17074 (
		\wishbone_bd_ram_mem1_reg[71][11]/P0001 ,
		_w12798_,
		_w27586_
	);
	LUT2 #(
		.INIT('h8)
	) name17075 (
		\wishbone_bd_ram_mem1_reg[196][11]/P0001 ,
		_w13090_,
		_w27587_
	);
	LUT2 #(
		.INIT('h8)
	) name17076 (
		\wishbone_bd_ram_mem1_reg[119][11]/P0001 ,
		_w13048_,
		_w27588_
	);
	LUT2 #(
		.INIT('h8)
	) name17077 (
		\wishbone_bd_ram_mem1_reg[207][11]/P0001 ,
		_w13180_,
		_w27589_
	);
	LUT2 #(
		.INIT('h8)
	) name17078 (
		\wishbone_bd_ram_mem1_reg[32][11]/P0001 ,
		_w13120_,
		_w27590_
	);
	LUT2 #(
		.INIT('h8)
	) name17079 (
		\wishbone_bd_ram_mem1_reg[203][11]/P0001 ,
		_w13158_,
		_w27591_
	);
	LUT2 #(
		.INIT('h8)
	) name17080 (
		\wishbone_bd_ram_mem1_reg[7][11]/P0001 ,
		_w12728_,
		_w27592_
	);
	LUT2 #(
		.INIT('h8)
	) name17081 (
		\wishbone_bd_ram_mem1_reg[96][11]/P0001 ,
		_w12912_,
		_w27593_
	);
	LUT2 #(
		.INIT('h8)
	) name17082 (
		\wishbone_bd_ram_mem1_reg[6][11]/P0001 ,
		_w12968_,
		_w27594_
	);
	LUT2 #(
		.INIT('h8)
	) name17083 (
		\wishbone_bd_ram_mem1_reg[54][11]/P0001 ,
		_w12770_,
		_w27595_
	);
	LUT2 #(
		.INIT('h8)
	) name17084 (
		\wishbone_bd_ram_mem1_reg[194][11]/P0001 ,
		_w12772_,
		_w27596_
	);
	LUT2 #(
		.INIT('h8)
	) name17085 (
		\wishbone_bd_ram_mem1_reg[39][11]/P0001 ,
		_w13018_,
		_w27597_
	);
	LUT2 #(
		.INIT('h8)
	) name17086 (
		\wishbone_bd_ram_mem1_reg[133][11]/P0001 ,
		_w12761_,
		_w27598_
	);
	LUT2 #(
		.INIT('h8)
	) name17087 (
		\wishbone_bd_ram_mem1_reg[159][11]/P0001 ,
		_w12774_,
		_w27599_
	);
	LUT2 #(
		.INIT('h8)
	) name17088 (
		\wishbone_bd_ram_mem1_reg[139][11]/P0001 ,
		_w12814_,
		_w27600_
	);
	LUT2 #(
		.INIT('h8)
	) name17089 (
		\wishbone_bd_ram_mem1_reg[24][11]/P0001 ,
		_w13084_,
		_w27601_
	);
	LUT2 #(
		.INIT('h8)
	) name17090 (
		\wishbone_bd_ram_mem1_reg[240][11]/P0001 ,
		_w12864_,
		_w27602_
	);
	LUT2 #(
		.INIT('h8)
	) name17091 (
		\wishbone_bd_ram_mem1_reg[230][11]/P0001 ,
		_w13036_,
		_w27603_
	);
	LUT2 #(
		.INIT('h8)
	) name17092 (
		\wishbone_bd_ram_mem1_reg[126][11]/P0001 ,
		_w13218_,
		_w27604_
	);
	LUT2 #(
		.INIT('h8)
	) name17093 (
		\wishbone_bd_ram_mem1_reg[5][11]/P0001 ,
		_w12878_,
		_w27605_
	);
	LUT2 #(
		.INIT('h8)
	) name17094 (
		\wishbone_bd_ram_mem1_reg[143][11]/P0001 ,
		_w12922_,
		_w27606_
	);
	LUT2 #(
		.INIT('h8)
	) name17095 (
		\wishbone_bd_ram_mem1_reg[226][11]/P0001 ,
		_w13138_,
		_w27607_
	);
	LUT2 #(
		.INIT('h8)
	) name17096 (
		\wishbone_bd_ram_mem1_reg[70][11]/P0001 ,
		_w12840_,
		_w27608_
	);
	LUT2 #(
		.INIT('h8)
	) name17097 (
		\wishbone_bd_ram_mem1_reg[60][11]/P0001 ,
		_w13204_,
		_w27609_
	);
	LUT2 #(
		.INIT('h8)
	) name17098 (
		\wishbone_bd_ram_mem1_reg[228][11]/P0001 ,
		_w12765_,
		_w27610_
	);
	LUT2 #(
		.INIT('h8)
	) name17099 (
		\wishbone_bd_ram_mem1_reg[92][11]/P0001 ,
		_w13010_,
		_w27611_
	);
	LUT2 #(
		.INIT('h8)
	) name17100 (
		\wishbone_bd_ram_mem1_reg[13][11]/P0001 ,
		_w13178_,
		_w27612_
	);
	LUT2 #(
		.INIT('h8)
	) name17101 (
		\wishbone_bd_ram_mem1_reg[50][11]/P0001 ,
		_w13150_,
		_w27613_
	);
	LUT2 #(
		.INIT('h8)
	) name17102 (
		\wishbone_bd_ram_mem1_reg[229][11]/P0001 ,
		_w12711_,
		_w27614_
	);
	LUT2 #(
		.INIT('h8)
	) name17103 (
		\wishbone_bd_ram_mem1_reg[130][11]/P0001 ,
		_w12914_,
		_w27615_
	);
	LUT2 #(
		.INIT('h8)
	) name17104 (
		\wishbone_bd_ram_mem1_reg[187][11]/P0001 ,
		_w13196_,
		_w27616_
	);
	LUT2 #(
		.INIT('h8)
	) name17105 (
		\wishbone_bd_ram_mem1_reg[37][11]/P0001 ,
		_w13102_,
		_w27617_
	);
	LUT2 #(
		.INIT('h8)
	) name17106 (
		\wishbone_bd_ram_mem1_reg[167][11]/P0001 ,
		_w12986_,
		_w27618_
	);
	LUT2 #(
		.INIT('h8)
	) name17107 (
		\wishbone_bd_ram_mem1_reg[254][11]/P0001 ,
		_w12892_,
		_w27619_
	);
	LUT2 #(
		.INIT('h8)
	) name17108 (
		\wishbone_bd_ram_mem1_reg[198][11]/P0001 ,
		_w12832_,
		_w27620_
	);
	LUT2 #(
		.INIT('h8)
	) name17109 (
		\wishbone_bd_ram_mem1_reg[105][11]/P0001 ,
		_w12751_,
		_w27621_
	);
	LUT2 #(
		.INIT('h8)
	) name17110 (
		\wishbone_bd_ram_mem1_reg[52][11]/P0001 ,
		_w13082_,
		_w27622_
	);
	LUT2 #(
		.INIT('h8)
	) name17111 (
		\wishbone_bd_ram_mem1_reg[155][11]/P0001 ,
		_w13122_,
		_w27623_
	);
	LUT2 #(
		.INIT('h8)
	) name17112 (
		\wishbone_bd_ram_mem1_reg[85][11]/P0001 ,
		_w13216_,
		_w27624_
	);
	LUT2 #(
		.INIT('h8)
	) name17113 (
		\wishbone_bd_ram_mem1_reg[22][11]/P0001 ,
		_w13110_,
		_w27625_
	);
	LUT2 #(
		.INIT('h8)
	) name17114 (
		\wishbone_bd_ram_mem1_reg[193][11]/P0001 ,
		_w13056_,
		_w27626_
	);
	LUT2 #(
		.INIT('h8)
	) name17115 (
		\wishbone_bd_ram_mem1_reg[11][11]/P0001 ,
		_w13194_,
		_w27627_
	);
	LUT2 #(
		.INIT('h8)
	) name17116 (
		\wishbone_bd_ram_mem1_reg[145][11]/P0001 ,
		_w13106_,
		_w27628_
	);
	LUT2 #(
		.INIT('h8)
	) name17117 (
		\wishbone_bd_ram_mem1_reg[116][11]/P0001 ,
		_w12998_,
		_w27629_
	);
	LUT2 #(
		.INIT('h8)
	) name17118 (
		\wishbone_bd_ram_mem1_reg[29][11]/P0001 ,
		_w12952_,
		_w27630_
	);
	LUT2 #(
		.INIT('h8)
	) name17119 (
		\wishbone_bd_ram_mem1_reg[59][11]/P0001 ,
		_w12780_,
		_w27631_
	);
	LUT2 #(
		.INIT('h8)
	) name17120 (
		\wishbone_bd_ram_mem1_reg[204][11]/P0001 ,
		_w13162_,
		_w27632_
	);
	LUT2 #(
		.INIT('h8)
	) name17121 (
		\wishbone_bd_ram_mem1_reg[102][11]/P0001 ,
		_w12685_,
		_w27633_
	);
	LUT2 #(
		.INIT('h8)
	) name17122 (
		\wishbone_bd_ram_mem1_reg[158][11]/P0001 ,
		_w12898_,
		_w27634_
	);
	LUT2 #(
		.INIT('h8)
	) name17123 (
		\wishbone_bd_ram_mem1_reg[140][11]/P0001 ,
		_w12894_,
		_w27635_
	);
	LUT2 #(
		.INIT('h8)
	) name17124 (
		\wishbone_bd_ram_mem1_reg[137][11]/P0001 ,
		_w13168_,
		_w27636_
	);
	LUT2 #(
		.INIT('h8)
	) name17125 (
		\wishbone_bd_ram_mem1_reg[23][11]/P0001 ,
		_w13008_,
		_w27637_
	);
	LUT2 #(
		.INIT('h8)
	) name17126 (
		\wishbone_bd_ram_mem1_reg[249][11]/P0001 ,
		_w12900_,
		_w27638_
	);
	LUT2 #(
		.INIT('h8)
	) name17127 (
		\wishbone_bd_ram_mem1_reg[1][11]/P0001 ,
		_w13014_,
		_w27639_
	);
	LUT2 #(
		.INIT('h8)
	) name17128 (
		\wishbone_bd_ram_mem1_reg[209][11]/P0001 ,
		_w13152_,
		_w27640_
	);
	LUT2 #(
		.INIT('h8)
	) name17129 (
		\wishbone_bd_ram_mem1_reg[15][11]/P0001 ,
		_w13210_,
		_w27641_
	);
	LUT2 #(
		.INIT('h8)
	) name17130 (
		\wishbone_bd_ram_mem1_reg[97][11]/P0001 ,
		_w13096_,
		_w27642_
	);
	LUT2 #(
		.INIT('h8)
	) name17131 (
		\wishbone_bd_ram_mem1_reg[94][11]/P0001 ,
		_w13186_,
		_w27643_
	);
	LUT2 #(
		.INIT('h8)
	) name17132 (
		\wishbone_bd_ram_mem1_reg[195][11]/P0001 ,
		_w13144_,
		_w27644_
	);
	LUT2 #(
		.INIT('h8)
	) name17133 (
		\wishbone_bd_ram_mem1_reg[156][11]/P0001 ,
		_w13190_,
		_w27645_
	);
	LUT2 #(
		.INIT('h8)
	) name17134 (
		\wishbone_bd_ram_mem1_reg[225][11]/P0001 ,
		_w13092_,
		_w27646_
	);
	LUT2 #(
		.INIT('h8)
	) name17135 (
		\wishbone_bd_ram_mem1_reg[238][11]/P0001 ,
		_w13160_,
		_w27647_
	);
	LUT2 #(
		.INIT('h8)
	) name17136 (
		\wishbone_bd_ram_mem1_reg[57][11]/P0001 ,
		_w13116_,
		_w27648_
	);
	LUT2 #(
		.INIT('h8)
	) name17137 (
		\wishbone_bd_ram_mem1_reg[235][11]/P0001 ,
		_w12696_,
		_w27649_
	);
	LUT2 #(
		.INIT('h8)
	) name17138 (
		\wishbone_bd_ram_mem1_reg[135][11]/P0001 ,
		_w13124_,
		_w27650_
	);
	LUT2 #(
		.INIT('h8)
	) name17139 (
		\wishbone_bd_ram_mem1_reg[149][11]/P0001 ,
		_w12741_,
		_w27651_
	);
	LUT2 #(
		.INIT('h8)
	) name17140 (
		\wishbone_bd_ram_mem1_reg[63][11]/P0001 ,
		_w12850_,
		_w27652_
	);
	LUT2 #(
		.INIT('h8)
	) name17141 (
		\wishbone_bd_ram_mem1_reg[251][11]/P0001 ,
		_w13054_,
		_w27653_
	);
	LUT2 #(
		.INIT('h8)
	) name17142 (
		\wishbone_bd_ram_mem1_reg[77][11]/P0001 ,
		_w12982_,
		_w27654_
	);
	LUT2 #(
		.INIT('h8)
	) name17143 (
		\wishbone_bd_ram_mem1_reg[165][11]/P0001 ,
		_w13044_,
		_w27655_
	);
	LUT2 #(
		.INIT('h8)
	) name17144 (
		\wishbone_bd_ram_mem1_reg[244][11]/P0001 ,
		_w12747_,
		_w27656_
	);
	LUT2 #(
		.INIT('h8)
	) name17145 (
		\wishbone_bd_ram_mem1_reg[86][11]/P0001 ,
		_w12735_,
		_w27657_
	);
	LUT2 #(
		.INIT('h8)
	) name17146 (
		\wishbone_bd_ram_mem1_reg[19][11]/P0001 ,
		_w13012_,
		_w27658_
	);
	LUT2 #(
		.INIT('h8)
	) name17147 (
		\wishbone_bd_ram_mem1_reg[166][11]/P0001 ,
		_w13040_,
		_w27659_
	);
	LUT2 #(
		.INIT('h8)
	) name17148 (
		\wishbone_bd_ram_mem1_reg[34][11]/P0001 ,
		_w12930_,
		_w27660_
	);
	LUT2 #(
		.INIT('h8)
	) name17149 (
		\wishbone_bd_ram_mem1_reg[150][11]/P0001 ,
		_w13136_,
		_w27661_
	);
	LUT2 #(
		.INIT('h8)
	) name17150 (
		\wishbone_bd_ram_mem1_reg[216][11]/P0001 ,
		_w13028_,
		_w27662_
	);
	LUT2 #(
		.INIT('h8)
	) name17151 (
		\wishbone_bd_ram_mem1_reg[208][11]/P0001 ,
		_w13032_,
		_w27663_
	);
	LUT2 #(
		.INIT('h8)
	) name17152 (
		\wishbone_bd_ram_mem1_reg[115][11]/P0001 ,
		_w13112_,
		_w27664_
	);
	LUT2 #(
		.INIT('h8)
	) name17153 (
		\wishbone_bd_ram_mem1_reg[14][11]/P0001 ,
		_w13086_,
		_w27665_
	);
	LUT2 #(
		.INIT('h8)
	) name17154 (
		\wishbone_bd_ram_mem1_reg[128][11]/P0001 ,
		_w12793_,
		_w27666_
	);
	LUT2 #(
		.INIT('h8)
	) name17155 (
		\wishbone_bd_ram_mem1_reg[144][11]/P0001 ,
		_w12756_,
		_w27667_
	);
	LUT2 #(
		.INIT('h8)
	) name17156 (
		\wishbone_bd_ram_mem1_reg[170][11]/P0001 ,
		_w13030_,
		_w27668_
	);
	LUT2 #(
		.INIT('h8)
	) name17157 (
		\wishbone_bd_ram_mem1_reg[186][11]/P0001 ,
		_w12783_,
		_w27669_
	);
	LUT2 #(
		.INIT('h8)
	) name17158 (
		\wishbone_bd_ram_mem1_reg[25][11]/P0001 ,
		_w13108_,
		_w27670_
	);
	LUT2 #(
		.INIT('h8)
	) name17159 (
		\wishbone_bd_ram_mem1_reg[188][11]/P0001 ,
		_w12948_,
		_w27671_
	);
	LUT2 #(
		.INIT('h8)
	) name17160 (
		\wishbone_bd_ram_mem1_reg[172][11]/P0001 ,
		_w12944_,
		_w27672_
	);
	LUT2 #(
		.INIT('h8)
	) name17161 (
		\wishbone_bd_ram_mem1_reg[49][11]/P0001 ,
		_w12994_,
		_w27673_
	);
	LUT2 #(
		.INIT('h8)
	) name17162 (
		\wishbone_bd_ram_mem1_reg[104][11]/P0001 ,
		_w13148_,
		_w27674_
	);
	LUT2 #(
		.INIT('h8)
	) name17163 (
		\wishbone_bd_ram_mem1_reg[76][11]/P0001 ,
		_w13184_,
		_w27675_
	);
	LUT2 #(
		.INIT('h8)
	) name17164 (
		\wishbone_bd_ram_mem1_reg[73][11]/P0001 ,
		_w12918_,
		_w27676_
	);
	LUT2 #(
		.INIT('h8)
	) name17165 (
		\wishbone_bd_ram_mem1_reg[200][11]/P0001 ,
		_w12988_,
		_w27677_
	);
	LUT2 #(
		.INIT('h8)
	) name17166 (
		\wishbone_bd_ram_mem1_reg[114][11]/P0001 ,
		_w13202_,
		_w27678_
	);
	LUT2 #(
		.INIT('h8)
	) name17167 (
		\wishbone_bd_ram_mem1_reg[252][11]/P0001 ,
		_w13080_,
		_w27679_
	);
	LUT2 #(
		.INIT('h8)
	) name17168 (
		\wishbone_bd_ram_mem1_reg[201][11]/P0001 ,
		_w12822_,
		_w27680_
	);
	LUT2 #(
		.INIT('h8)
	) name17169 (
		\wishbone_bd_ram_mem1_reg[103][11]/P0001 ,
		_w12846_,
		_w27681_
	);
	LUT2 #(
		.INIT('h8)
	) name17170 (
		\wishbone_bd_ram_mem1_reg[205][11]/P0001 ,
		_w13068_,
		_w27682_
	);
	LUT2 #(
		.INIT('h8)
	) name17171 (
		\wishbone_bd_ram_mem1_reg[132][11]/P0001 ,
		_w12992_,
		_w27683_
	);
	LUT2 #(
		.INIT('h8)
	) name17172 (
		\wishbone_bd_ram_mem1_reg[247][11]/P0001 ,
		_w12818_,
		_w27684_
	);
	LUT2 #(
		.INIT('h8)
	) name17173 (
		\wishbone_bd_ram_mem1_reg[241][11]/P0001 ,
		_w13006_,
		_w27685_
	);
	LUT2 #(
		.INIT('h8)
	) name17174 (
		\wishbone_bd_ram_mem1_reg[141][11]/P0001 ,
		_w13004_,
		_w27686_
	);
	LUT2 #(
		.INIT('h8)
	) name17175 (
		\wishbone_bd_ram_mem1_reg[51][11]/P0001 ,
		_w13024_,
		_w27687_
	);
	LUT2 #(
		.INIT('h8)
	) name17176 (
		\wishbone_bd_ram_mem1_reg[129][11]/P0001 ,
		_w12776_,
		_w27688_
	);
	LUT2 #(
		.INIT('h8)
	) name17177 (
		\wishbone_bd_ram_mem1_reg[236][11]/P0001 ,
		_w12731_,
		_w27689_
	);
	LUT2 #(
		.INIT('h8)
	) name17178 (
		\wishbone_bd_ram_mem1_reg[2][11]/P0001 ,
		_w13088_,
		_w27690_
	);
	LUT2 #(
		.INIT('h8)
	) name17179 (
		\wishbone_bd_ram_mem1_reg[199][11]/P0001 ,
		_w12768_,
		_w27691_
	);
	LUT2 #(
		.INIT('h8)
	) name17180 (
		\wishbone_bd_ram_mem1_reg[81][11]/P0001 ,
		_w12950_,
		_w27692_
	);
	LUT2 #(
		.INIT('h8)
	) name17181 (
		\wishbone_bd_ram_mem1_reg[67][11]/P0001 ,
		_w13134_,
		_w27693_
	);
	LUT2 #(
		.INIT('h8)
	) name17182 (
		\wishbone_bd_ram_mem1_reg[9][11]/P0001 ,
		_w12808_,
		_w27694_
	);
	LUT2 #(
		.INIT('h8)
	) name17183 (
		\wishbone_bd_ram_mem1_reg[100][11]/P0001 ,
		_w12960_,
		_w27695_
	);
	LUT2 #(
		.INIT('h8)
	) name17184 (
		\wishbone_bd_ram_mem1_reg[0][11]/P0001 ,
		_w12717_,
		_w27696_
	);
	LUT2 #(
		.INIT('h8)
	) name17185 (
		\wishbone_bd_ram_mem1_reg[223][11]/P0001 ,
		_w12838_,
		_w27697_
	);
	LUT2 #(
		.INIT('h8)
	) name17186 (
		\wishbone_bd_ram_mem1_reg[43][11]/P0001 ,
		_w13200_,
		_w27698_
	);
	LUT2 #(
		.INIT('h8)
	) name17187 (
		\wishbone_bd_ram_mem1_reg[233][11]/P0001 ,
		_w12836_,
		_w27699_
	);
	LUT2 #(
		.INIT('h8)
	) name17188 (
		\wishbone_bd_ram_mem1_reg[152][11]/P0001 ,
		_w12966_,
		_w27700_
	);
	LUT2 #(
		.INIT('h8)
	) name17189 (
		\wishbone_bd_ram_mem1_reg[109][11]/P0001 ,
		_w12888_,
		_w27701_
	);
	LUT2 #(
		.INIT('h8)
	) name17190 (
		\wishbone_bd_ram_mem1_reg[88][11]/P0001 ,
		_w12860_,
		_w27702_
	);
	LUT2 #(
		.INIT('h8)
	) name17191 (
		\wishbone_bd_ram_mem1_reg[3][11]/P0001 ,
		_w12866_,
		_w27703_
	);
	LUT2 #(
		.INIT('h8)
	) name17192 (
		\wishbone_bd_ram_mem1_reg[17][11]/P0001 ,
		_w12848_,
		_w27704_
	);
	LUT2 #(
		.INIT('h8)
	) name17193 (
		\wishbone_bd_ram_mem1_reg[41][11]/P0001 ,
		_w13052_,
		_w27705_
	);
	LUT2 #(
		.INIT('h8)
	) name17194 (
		\wishbone_bd_ram_mem1_reg[89][11]/P0001 ,
		_w12964_,
		_w27706_
	);
	LUT2 #(
		.INIT('h8)
	) name17195 (
		\wishbone_bd_ram_mem1_reg[45][11]/P0001 ,
		_w12908_,
		_w27707_
	);
	LUT2 #(
		.INIT('h8)
	) name17196 (
		\wishbone_bd_ram_mem1_reg[248][11]/P0001 ,
		_w12789_,
		_w27708_
	);
	LUT2 #(
		.INIT('h8)
	) name17197 (
		\wishbone_bd_ram_mem1_reg[227][11]/P0001 ,
		_w12936_,
		_w27709_
	);
	LUT2 #(
		.INIT('h8)
	) name17198 (
		\wishbone_bd_ram_mem1_reg[255][11]/P0001 ,
		_w13072_,
		_w27710_
	);
	LUT2 #(
		.INIT('h8)
	) name17199 (
		\wishbone_bd_ram_mem1_reg[53][11]/P0001 ,
		_w13020_,
		_w27711_
	);
	LUT2 #(
		.INIT('h8)
	) name17200 (
		\wishbone_bd_ram_mem1_reg[169][11]/P0001 ,
		_w12722_,
		_w27712_
	);
	LUT2 #(
		.INIT('h8)
	) name17201 (
		\wishbone_bd_ram_mem1_reg[215][11]/P0001 ,
		_w12974_,
		_w27713_
	);
	LUT2 #(
		.INIT('h8)
	) name17202 (
		\wishbone_bd_ram_mem1_reg[93][11]/P0001 ,
		_w13016_,
		_w27714_
	);
	LUT2 #(
		.INIT('h8)
	) name17203 (
		\wishbone_bd_ram_mem1_reg[120][11]/P0001 ,
		_w12707_,
		_w27715_
	);
	LUT2 #(
		.INIT('h8)
	) name17204 (
		\wishbone_bd_ram_mem1_reg[212][11]/P0001 ,
		_w12796_,
		_w27716_
	);
	LUT2 #(
		.INIT('h8)
	) name17205 (
		\wishbone_bd_ram_mem1_reg[47][11]/P0001 ,
		_w12904_,
		_w27717_
	);
	LUT2 #(
		.INIT('h8)
	) name17206 (
		\wishbone_bd_ram_mem1_reg[117][11]/P0001 ,
		_w12715_,
		_w27718_
	);
	LUT2 #(
		.INIT('h8)
	) name17207 (
		\wishbone_bd_ram_mem1_reg[112][11]/P0001 ,
		_w12733_,
		_w27719_
	);
	LUT2 #(
		.INIT('h8)
	) name17208 (
		\wishbone_bd_ram_mem1_reg[87][11]/P0001 ,
		_w13154_,
		_w27720_
	);
	LUT2 #(
		.INIT('h8)
	) name17209 (
		\wishbone_bd_ram_mem1_reg[72][11]/P0001 ,
		_w12810_,
		_w27721_
	);
	LUT2 #(
		.INIT('h8)
	) name17210 (
		\wishbone_bd_ram_mem1_reg[66][11]/P0001 ,
		_w12824_,
		_w27722_
	);
	LUT2 #(
		.INIT('h8)
	) name17211 (
		\wishbone_bd_ram_mem1_reg[108][11]/P0001 ,
		_w13156_,
		_w27723_
	);
	LUT2 #(
		.INIT('h8)
	) name17212 (
		\wishbone_bd_ram_mem1_reg[243][11]/P0001 ,
		_w12804_,
		_w27724_
	);
	LUT2 #(
		.INIT('h1)
	) name17213 (
		_w27469_,
		_w27470_,
		_w27725_
	);
	LUT2 #(
		.INIT('h1)
	) name17214 (
		_w27471_,
		_w27472_,
		_w27726_
	);
	LUT2 #(
		.INIT('h1)
	) name17215 (
		_w27473_,
		_w27474_,
		_w27727_
	);
	LUT2 #(
		.INIT('h1)
	) name17216 (
		_w27475_,
		_w27476_,
		_w27728_
	);
	LUT2 #(
		.INIT('h1)
	) name17217 (
		_w27477_,
		_w27478_,
		_w27729_
	);
	LUT2 #(
		.INIT('h1)
	) name17218 (
		_w27479_,
		_w27480_,
		_w27730_
	);
	LUT2 #(
		.INIT('h1)
	) name17219 (
		_w27481_,
		_w27482_,
		_w27731_
	);
	LUT2 #(
		.INIT('h1)
	) name17220 (
		_w27483_,
		_w27484_,
		_w27732_
	);
	LUT2 #(
		.INIT('h1)
	) name17221 (
		_w27485_,
		_w27486_,
		_w27733_
	);
	LUT2 #(
		.INIT('h1)
	) name17222 (
		_w27487_,
		_w27488_,
		_w27734_
	);
	LUT2 #(
		.INIT('h1)
	) name17223 (
		_w27489_,
		_w27490_,
		_w27735_
	);
	LUT2 #(
		.INIT('h1)
	) name17224 (
		_w27491_,
		_w27492_,
		_w27736_
	);
	LUT2 #(
		.INIT('h1)
	) name17225 (
		_w27493_,
		_w27494_,
		_w27737_
	);
	LUT2 #(
		.INIT('h1)
	) name17226 (
		_w27495_,
		_w27496_,
		_w27738_
	);
	LUT2 #(
		.INIT('h1)
	) name17227 (
		_w27497_,
		_w27498_,
		_w27739_
	);
	LUT2 #(
		.INIT('h1)
	) name17228 (
		_w27499_,
		_w27500_,
		_w27740_
	);
	LUT2 #(
		.INIT('h1)
	) name17229 (
		_w27501_,
		_w27502_,
		_w27741_
	);
	LUT2 #(
		.INIT('h1)
	) name17230 (
		_w27503_,
		_w27504_,
		_w27742_
	);
	LUT2 #(
		.INIT('h1)
	) name17231 (
		_w27505_,
		_w27506_,
		_w27743_
	);
	LUT2 #(
		.INIT('h1)
	) name17232 (
		_w27507_,
		_w27508_,
		_w27744_
	);
	LUT2 #(
		.INIT('h1)
	) name17233 (
		_w27509_,
		_w27510_,
		_w27745_
	);
	LUT2 #(
		.INIT('h1)
	) name17234 (
		_w27511_,
		_w27512_,
		_w27746_
	);
	LUT2 #(
		.INIT('h1)
	) name17235 (
		_w27513_,
		_w27514_,
		_w27747_
	);
	LUT2 #(
		.INIT('h1)
	) name17236 (
		_w27515_,
		_w27516_,
		_w27748_
	);
	LUT2 #(
		.INIT('h1)
	) name17237 (
		_w27517_,
		_w27518_,
		_w27749_
	);
	LUT2 #(
		.INIT('h1)
	) name17238 (
		_w27519_,
		_w27520_,
		_w27750_
	);
	LUT2 #(
		.INIT('h1)
	) name17239 (
		_w27521_,
		_w27522_,
		_w27751_
	);
	LUT2 #(
		.INIT('h1)
	) name17240 (
		_w27523_,
		_w27524_,
		_w27752_
	);
	LUT2 #(
		.INIT('h1)
	) name17241 (
		_w27525_,
		_w27526_,
		_w27753_
	);
	LUT2 #(
		.INIT('h1)
	) name17242 (
		_w27527_,
		_w27528_,
		_w27754_
	);
	LUT2 #(
		.INIT('h1)
	) name17243 (
		_w27529_,
		_w27530_,
		_w27755_
	);
	LUT2 #(
		.INIT('h1)
	) name17244 (
		_w27531_,
		_w27532_,
		_w27756_
	);
	LUT2 #(
		.INIT('h1)
	) name17245 (
		_w27533_,
		_w27534_,
		_w27757_
	);
	LUT2 #(
		.INIT('h1)
	) name17246 (
		_w27535_,
		_w27536_,
		_w27758_
	);
	LUT2 #(
		.INIT('h1)
	) name17247 (
		_w27537_,
		_w27538_,
		_w27759_
	);
	LUT2 #(
		.INIT('h1)
	) name17248 (
		_w27539_,
		_w27540_,
		_w27760_
	);
	LUT2 #(
		.INIT('h1)
	) name17249 (
		_w27541_,
		_w27542_,
		_w27761_
	);
	LUT2 #(
		.INIT('h1)
	) name17250 (
		_w27543_,
		_w27544_,
		_w27762_
	);
	LUT2 #(
		.INIT('h1)
	) name17251 (
		_w27545_,
		_w27546_,
		_w27763_
	);
	LUT2 #(
		.INIT('h1)
	) name17252 (
		_w27547_,
		_w27548_,
		_w27764_
	);
	LUT2 #(
		.INIT('h1)
	) name17253 (
		_w27549_,
		_w27550_,
		_w27765_
	);
	LUT2 #(
		.INIT('h1)
	) name17254 (
		_w27551_,
		_w27552_,
		_w27766_
	);
	LUT2 #(
		.INIT('h1)
	) name17255 (
		_w27553_,
		_w27554_,
		_w27767_
	);
	LUT2 #(
		.INIT('h1)
	) name17256 (
		_w27555_,
		_w27556_,
		_w27768_
	);
	LUT2 #(
		.INIT('h1)
	) name17257 (
		_w27557_,
		_w27558_,
		_w27769_
	);
	LUT2 #(
		.INIT('h1)
	) name17258 (
		_w27559_,
		_w27560_,
		_w27770_
	);
	LUT2 #(
		.INIT('h1)
	) name17259 (
		_w27561_,
		_w27562_,
		_w27771_
	);
	LUT2 #(
		.INIT('h1)
	) name17260 (
		_w27563_,
		_w27564_,
		_w27772_
	);
	LUT2 #(
		.INIT('h1)
	) name17261 (
		_w27565_,
		_w27566_,
		_w27773_
	);
	LUT2 #(
		.INIT('h1)
	) name17262 (
		_w27567_,
		_w27568_,
		_w27774_
	);
	LUT2 #(
		.INIT('h1)
	) name17263 (
		_w27569_,
		_w27570_,
		_w27775_
	);
	LUT2 #(
		.INIT('h1)
	) name17264 (
		_w27571_,
		_w27572_,
		_w27776_
	);
	LUT2 #(
		.INIT('h1)
	) name17265 (
		_w27573_,
		_w27574_,
		_w27777_
	);
	LUT2 #(
		.INIT('h1)
	) name17266 (
		_w27575_,
		_w27576_,
		_w27778_
	);
	LUT2 #(
		.INIT('h1)
	) name17267 (
		_w27577_,
		_w27578_,
		_w27779_
	);
	LUT2 #(
		.INIT('h1)
	) name17268 (
		_w27579_,
		_w27580_,
		_w27780_
	);
	LUT2 #(
		.INIT('h1)
	) name17269 (
		_w27581_,
		_w27582_,
		_w27781_
	);
	LUT2 #(
		.INIT('h1)
	) name17270 (
		_w27583_,
		_w27584_,
		_w27782_
	);
	LUT2 #(
		.INIT('h1)
	) name17271 (
		_w27585_,
		_w27586_,
		_w27783_
	);
	LUT2 #(
		.INIT('h1)
	) name17272 (
		_w27587_,
		_w27588_,
		_w27784_
	);
	LUT2 #(
		.INIT('h1)
	) name17273 (
		_w27589_,
		_w27590_,
		_w27785_
	);
	LUT2 #(
		.INIT('h1)
	) name17274 (
		_w27591_,
		_w27592_,
		_w27786_
	);
	LUT2 #(
		.INIT('h1)
	) name17275 (
		_w27593_,
		_w27594_,
		_w27787_
	);
	LUT2 #(
		.INIT('h1)
	) name17276 (
		_w27595_,
		_w27596_,
		_w27788_
	);
	LUT2 #(
		.INIT('h1)
	) name17277 (
		_w27597_,
		_w27598_,
		_w27789_
	);
	LUT2 #(
		.INIT('h1)
	) name17278 (
		_w27599_,
		_w27600_,
		_w27790_
	);
	LUT2 #(
		.INIT('h1)
	) name17279 (
		_w27601_,
		_w27602_,
		_w27791_
	);
	LUT2 #(
		.INIT('h1)
	) name17280 (
		_w27603_,
		_w27604_,
		_w27792_
	);
	LUT2 #(
		.INIT('h1)
	) name17281 (
		_w27605_,
		_w27606_,
		_w27793_
	);
	LUT2 #(
		.INIT('h1)
	) name17282 (
		_w27607_,
		_w27608_,
		_w27794_
	);
	LUT2 #(
		.INIT('h1)
	) name17283 (
		_w27609_,
		_w27610_,
		_w27795_
	);
	LUT2 #(
		.INIT('h1)
	) name17284 (
		_w27611_,
		_w27612_,
		_w27796_
	);
	LUT2 #(
		.INIT('h1)
	) name17285 (
		_w27613_,
		_w27614_,
		_w27797_
	);
	LUT2 #(
		.INIT('h1)
	) name17286 (
		_w27615_,
		_w27616_,
		_w27798_
	);
	LUT2 #(
		.INIT('h1)
	) name17287 (
		_w27617_,
		_w27618_,
		_w27799_
	);
	LUT2 #(
		.INIT('h1)
	) name17288 (
		_w27619_,
		_w27620_,
		_w27800_
	);
	LUT2 #(
		.INIT('h1)
	) name17289 (
		_w27621_,
		_w27622_,
		_w27801_
	);
	LUT2 #(
		.INIT('h1)
	) name17290 (
		_w27623_,
		_w27624_,
		_w27802_
	);
	LUT2 #(
		.INIT('h1)
	) name17291 (
		_w27625_,
		_w27626_,
		_w27803_
	);
	LUT2 #(
		.INIT('h1)
	) name17292 (
		_w27627_,
		_w27628_,
		_w27804_
	);
	LUT2 #(
		.INIT('h1)
	) name17293 (
		_w27629_,
		_w27630_,
		_w27805_
	);
	LUT2 #(
		.INIT('h1)
	) name17294 (
		_w27631_,
		_w27632_,
		_w27806_
	);
	LUT2 #(
		.INIT('h1)
	) name17295 (
		_w27633_,
		_w27634_,
		_w27807_
	);
	LUT2 #(
		.INIT('h1)
	) name17296 (
		_w27635_,
		_w27636_,
		_w27808_
	);
	LUT2 #(
		.INIT('h1)
	) name17297 (
		_w27637_,
		_w27638_,
		_w27809_
	);
	LUT2 #(
		.INIT('h1)
	) name17298 (
		_w27639_,
		_w27640_,
		_w27810_
	);
	LUT2 #(
		.INIT('h1)
	) name17299 (
		_w27641_,
		_w27642_,
		_w27811_
	);
	LUT2 #(
		.INIT('h1)
	) name17300 (
		_w27643_,
		_w27644_,
		_w27812_
	);
	LUT2 #(
		.INIT('h1)
	) name17301 (
		_w27645_,
		_w27646_,
		_w27813_
	);
	LUT2 #(
		.INIT('h1)
	) name17302 (
		_w27647_,
		_w27648_,
		_w27814_
	);
	LUT2 #(
		.INIT('h1)
	) name17303 (
		_w27649_,
		_w27650_,
		_w27815_
	);
	LUT2 #(
		.INIT('h1)
	) name17304 (
		_w27651_,
		_w27652_,
		_w27816_
	);
	LUT2 #(
		.INIT('h1)
	) name17305 (
		_w27653_,
		_w27654_,
		_w27817_
	);
	LUT2 #(
		.INIT('h1)
	) name17306 (
		_w27655_,
		_w27656_,
		_w27818_
	);
	LUT2 #(
		.INIT('h1)
	) name17307 (
		_w27657_,
		_w27658_,
		_w27819_
	);
	LUT2 #(
		.INIT('h1)
	) name17308 (
		_w27659_,
		_w27660_,
		_w27820_
	);
	LUT2 #(
		.INIT('h1)
	) name17309 (
		_w27661_,
		_w27662_,
		_w27821_
	);
	LUT2 #(
		.INIT('h1)
	) name17310 (
		_w27663_,
		_w27664_,
		_w27822_
	);
	LUT2 #(
		.INIT('h1)
	) name17311 (
		_w27665_,
		_w27666_,
		_w27823_
	);
	LUT2 #(
		.INIT('h1)
	) name17312 (
		_w27667_,
		_w27668_,
		_w27824_
	);
	LUT2 #(
		.INIT('h1)
	) name17313 (
		_w27669_,
		_w27670_,
		_w27825_
	);
	LUT2 #(
		.INIT('h1)
	) name17314 (
		_w27671_,
		_w27672_,
		_w27826_
	);
	LUT2 #(
		.INIT('h1)
	) name17315 (
		_w27673_,
		_w27674_,
		_w27827_
	);
	LUT2 #(
		.INIT('h1)
	) name17316 (
		_w27675_,
		_w27676_,
		_w27828_
	);
	LUT2 #(
		.INIT('h1)
	) name17317 (
		_w27677_,
		_w27678_,
		_w27829_
	);
	LUT2 #(
		.INIT('h1)
	) name17318 (
		_w27679_,
		_w27680_,
		_w27830_
	);
	LUT2 #(
		.INIT('h1)
	) name17319 (
		_w27681_,
		_w27682_,
		_w27831_
	);
	LUT2 #(
		.INIT('h1)
	) name17320 (
		_w27683_,
		_w27684_,
		_w27832_
	);
	LUT2 #(
		.INIT('h1)
	) name17321 (
		_w27685_,
		_w27686_,
		_w27833_
	);
	LUT2 #(
		.INIT('h1)
	) name17322 (
		_w27687_,
		_w27688_,
		_w27834_
	);
	LUT2 #(
		.INIT('h1)
	) name17323 (
		_w27689_,
		_w27690_,
		_w27835_
	);
	LUT2 #(
		.INIT('h1)
	) name17324 (
		_w27691_,
		_w27692_,
		_w27836_
	);
	LUT2 #(
		.INIT('h1)
	) name17325 (
		_w27693_,
		_w27694_,
		_w27837_
	);
	LUT2 #(
		.INIT('h1)
	) name17326 (
		_w27695_,
		_w27696_,
		_w27838_
	);
	LUT2 #(
		.INIT('h1)
	) name17327 (
		_w27697_,
		_w27698_,
		_w27839_
	);
	LUT2 #(
		.INIT('h1)
	) name17328 (
		_w27699_,
		_w27700_,
		_w27840_
	);
	LUT2 #(
		.INIT('h1)
	) name17329 (
		_w27701_,
		_w27702_,
		_w27841_
	);
	LUT2 #(
		.INIT('h1)
	) name17330 (
		_w27703_,
		_w27704_,
		_w27842_
	);
	LUT2 #(
		.INIT('h1)
	) name17331 (
		_w27705_,
		_w27706_,
		_w27843_
	);
	LUT2 #(
		.INIT('h1)
	) name17332 (
		_w27707_,
		_w27708_,
		_w27844_
	);
	LUT2 #(
		.INIT('h1)
	) name17333 (
		_w27709_,
		_w27710_,
		_w27845_
	);
	LUT2 #(
		.INIT('h1)
	) name17334 (
		_w27711_,
		_w27712_,
		_w27846_
	);
	LUT2 #(
		.INIT('h1)
	) name17335 (
		_w27713_,
		_w27714_,
		_w27847_
	);
	LUT2 #(
		.INIT('h1)
	) name17336 (
		_w27715_,
		_w27716_,
		_w27848_
	);
	LUT2 #(
		.INIT('h1)
	) name17337 (
		_w27717_,
		_w27718_,
		_w27849_
	);
	LUT2 #(
		.INIT('h1)
	) name17338 (
		_w27719_,
		_w27720_,
		_w27850_
	);
	LUT2 #(
		.INIT('h1)
	) name17339 (
		_w27721_,
		_w27722_,
		_w27851_
	);
	LUT2 #(
		.INIT('h1)
	) name17340 (
		_w27723_,
		_w27724_,
		_w27852_
	);
	LUT2 #(
		.INIT('h8)
	) name17341 (
		_w27851_,
		_w27852_,
		_w27853_
	);
	LUT2 #(
		.INIT('h8)
	) name17342 (
		_w27849_,
		_w27850_,
		_w27854_
	);
	LUT2 #(
		.INIT('h8)
	) name17343 (
		_w27847_,
		_w27848_,
		_w27855_
	);
	LUT2 #(
		.INIT('h8)
	) name17344 (
		_w27845_,
		_w27846_,
		_w27856_
	);
	LUT2 #(
		.INIT('h8)
	) name17345 (
		_w27843_,
		_w27844_,
		_w27857_
	);
	LUT2 #(
		.INIT('h8)
	) name17346 (
		_w27841_,
		_w27842_,
		_w27858_
	);
	LUT2 #(
		.INIT('h8)
	) name17347 (
		_w27839_,
		_w27840_,
		_w27859_
	);
	LUT2 #(
		.INIT('h8)
	) name17348 (
		_w27837_,
		_w27838_,
		_w27860_
	);
	LUT2 #(
		.INIT('h8)
	) name17349 (
		_w27835_,
		_w27836_,
		_w27861_
	);
	LUT2 #(
		.INIT('h8)
	) name17350 (
		_w27833_,
		_w27834_,
		_w27862_
	);
	LUT2 #(
		.INIT('h8)
	) name17351 (
		_w27831_,
		_w27832_,
		_w27863_
	);
	LUT2 #(
		.INIT('h8)
	) name17352 (
		_w27829_,
		_w27830_,
		_w27864_
	);
	LUT2 #(
		.INIT('h8)
	) name17353 (
		_w27827_,
		_w27828_,
		_w27865_
	);
	LUT2 #(
		.INIT('h8)
	) name17354 (
		_w27825_,
		_w27826_,
		_w27866_
	);
	LUT2 #(
		.INIT('h8)
	) name17355 (
		_w27823_,
		_w27824_,
		_w27867_
	);
	LUT2 #(
		.INIT('h8)
	) name17356 (
		_w27821_,
		_w27822_,
		_w27868_
	);
	LUT2 #(
		.INIT('h8)
	) name17357 (
		_w27819_,
		_w27820_,
		_w27869_
	);
	LUT2 #(
		.INIT('h8)
	) name17358 (
		_w27817_,
		_w27818_,
		_w27870_
	);
	LUT2 #(
		.INIT('h8)
	) name17359 (
		_w27815_,
		_w27816_,
		_w27871_
	);
	LUT2 #(
		.INIT('h8)
	) name17360 (
		_w27813_,
		_w27814_,
		_w27872_
	);
	LUT2 #(
		.INIT('h8)
	) name17361 (
		_w27811_,
		_w27812_,
		_w27873_
	);
	LUT2 #(
		.INIT('h8)
	) name17362 (
		_w27809_,
		_w27810_,
		_w27874_
	);
	LUT2 #(
		.INIT('h8)
	) name17363 (
		_w27807_,
		_w27808_,
		_w27875_
	);
	LUT2 #(
		.INIT('h8)
	) name17364 (
		_w27805_,
		_w27806_,
		_w27876_
	);
	LUT2 #(
		.INIT('h8)
	) name17365 (
		_w27803_,
		_w27804_,
		_w27877_
	);
	LUT2 #(
		.INIT('h8)
	) name17366 (
		_w27801_,
		_w27802_,
		_w27878_
	);
	LUT2 #(
		.INIT('h8)
	) name17367 (
		_w27799_,
		_w27800_,
		_w27879_
	);
	LUT2 #(
		.INIT('h8)
	) name17368 (
		_w27797_,
		_w27798_,
		_w27880_
	);
	LUT2 #(
		.INIT('h8)
	) name17369 (
		_w27795_,
		_w27796_,
		_w27881_
	);
	LUT2 #(
		.INIT('h8)
	) name17370 (
		_w27793_,
		_w27794_,
		_w27882_
	);
	LUT2 #(
		.INIT('h8)
	) name17371 (
		_w27791_,
		_w27792_,
		_w27883_
	);
	LUT2 #(
		.INIT('h8)
	) name17372 (
		_w27789_,
		_w27790_,
		_w27884_
	);
	LUT2 #(
		.INIT('h8)
	) name17373 (
		_w27787_,
		_w27788_,
		_w27885_
	);
	LUT2 #(
		.INIT('h8)
	) name17374 (
		_w27785_,
		_w27786_,
		_w27886_
	);
	LUT2 #(
		.INIT('h8)
	) name17375 (
		_w27783_,
		_w27784_,
		_w27887_
	);
	LUT2 #(
		.INIT('h8)
	) name17376 (
		_w27781_,
		_w27782_,
		_w27888_
	);
	LUT2 #(
		.INIT('h8)
	) name17377 (
		_w27779_,
		_w27780_,
		_w27889_
	);
	LUT2 #(
		.INIT('h8)
	) name17378 (
		_w27777_,
		_w27778_,
		_w27890_
	);
	LUT2 #(
		.INIT('h8)
	) name17379 (
		_w27775_,
		_w27776_,
		_w27891_
	);
	LUT2 #(
		.INIT('h8)
	) name17380 (
		_w27773_,
		_w27774_,
		_w27892_
	);
	LUT2 #(
		.INIT('h8)
	) name17381 (
		_w27771_,
		_w27772_,
		_w27893_
	);
	LUT2 #(
		.INIT('h8)
	) name17382 (
		_w27769_,
		_w27770_,
		_w27894_
	);
	LUT2 #(
		.INIT('h8)
	) name17383 (
		_w27767_,
		_w27768_,
		_w27895_
	);
	LUT2 #(
		.INIT('h8)
	) name17384 (
		_w27765_,
		_w27766_,
		_w27896_
	);
	LUT2 #(
		.INIT('h8)
	) name17385 (
		_w27763_,
		_w27764_,
		_w27897_
	);
	LUT2 #(
		.INIT('h8)
	) name17386 (
		_w27761_,
		_w27762_,
		_w27898_
	);
	LUT2 #(
		.INIT('h8)
	) name17387 (
		_w27759_,
		_w27760_,
		_w27899_
	);
	LUT2 #(
		.INIT('h8)
	) name17388 (
		_w27757_,
		_w27758_,
		_w27900_
	);
	LUT2 #(
		.INIT('h8)
	) name17389 (
		_w27755_,
		_w27756_,
		_w27901_
	);
	LUT2 #(
		.INIT('h8)
	) name17390 (
		_w27753_,
		_w27754_,
		_w27902_
	);
	LUT2 #(
		.INIT('h8)
	) name17391 (
		_w27751_,
		_w27752_,
		_w27903_
	);
	LUT2 #(
		.INIT('h8)
	) name17392 (
		_w27749_,
		_w27750_,
		_w27904_
	);
	LUT2 #(
		.INIT('h8)
	) name17393 (
		_w27747_,
		_w27748_,
		_w27905_
	);
	LUT2 #(
		.INIT('h8)
	) name17394 (
		_w27745_,
		_w27746_,
		_w27906_
	);
	LUT2 #(
		.INIT('h8)
	) name17395 (
		_w27743_,
		_w27744_,
		_w27907_
	);
	LUT2 #(
		.INIT('h8)
	) name17396 (
		_w27741_,
		_w27742_,
		_w27908_
	);
	LUT2 #(
		.INIT('h8)
	) name17397 (
		_w27739_,
		_w27740_,
		_w27909_
	);
	LUT2 #(
		.INIT('h8)
	) name17398 (
		_w27737_,
		_w27738_,
		_w27910_
	);
	LUT2 #(
		.INIT('h8)
	) name17399 (
		_w27735_,
		_w27736_,
		_w27911_
	);
	LUT2 #(
		.INIT('h8)
	) name17400 (
		_w27733_,
		_w27734_,
		_w27912_
	);
	LUT2 #(
		.INIT('h8)
	) name17401 (
		_w27731_,
		_w27732_,
		_w27913_
	);
	LUT2 #(
		.INIT('h8)
	) name17402 (
		_w27729_,
		_w27730_,
		_w27914_
	);
	LUT2 #(
		.INIT('h8)
	) name17403 (
		_w27727_,
		_w27728_,
		_w27915_
	);
	LUT2 #(
		.INIT('h8)
	) name17404 (
		_w27725_,
		_w27726_,
		_w27916_
	);
	LUT2 #(
		.INIT('h8)
	) name17405 (
		_w27915_,
		_w27916_,
		_w27917_
	);
	LUT2 #(
		.INIT('h8)
	) name17406 (
		_w27913_,
		_w27914_,
		_w27918_
	);
	LUT2 #(
		.INIT('h8)
	) name17407 (
		_w27911_,
		_w27912_,
		_w27919_
	);
	LUT2 #(
		.INIT('h8)
	) name17408 (
		_w27909_,
		_w27910_,
		_w27920_
	);
	LUT2 #(
		.INIT('h8)
	) name17409 (
		_w27907_,
		_w27908_,
		_w27921_
	);
	LUT2 #(
		.INIT('h8)
	) name17410 (
		_w27905_,
		_w27906_,
		_w27922_
	);
	LUT2 #(
		.INIT('h8)
	) name17411 (
		_w27903_,
		_w27904_,
		_w27923_
	);
	LUT2 #(
		.INIT('h8)
	) name17412 (
		_w27901_,
		_w27902_,
		_w27924_
	);
	LUT2 #(
		.INIT('h8)
	) name17413 (
		_w27899_,
		_w27900_,
		_w27925_
	);
	LUT2 #(
		.INIT('h8)
	) name17414 (
		_w27897_,
		_w27898_,
		_w27926_
	);
	LUT2 #(
		.INIT('h8)
	) name17415 (
		_w27895_,
		_w27896_,
		_w27927_
	);
	LUT2 #(
		.INIT('h8)
	) name17416 (
		_w27893_,
		_w27894_,
		_w27928_
	);
	LUT2 #(
		.INIT('h8)
	) name17417 (
		_w27891_,
		_w27892_,
		_w27929_
	);
	LUT2 #(
		.INIT('h8)
	) name17418 (
		_w27889_,
		_w27890_,
		_w27930_
	);
	LUT2 #(
		.INIT('h8)
	) name17419 (
		_w27887_,
		_w27888_,
		_w27931_
	);
	LUT2 #(
		.INIT('h8)
	) name17420 (
		_w27885_,
		_w27886_,
		_w27932_
	);
	LUT2 #(
		.INIT('h8)
	) name17421 (
		_w27883_,
		_w27884_,
		_w27933_
	);
	LUT2 #(
		.INIT('h8)
	) name17422 (
		_w27881_,
		_w27882_,
		_w27934_
	);
	LUT2 #(
		.INIT('h8)
	) name17423 (
		_w27879_,
		_w27880_,
		_w27935_
	);
	LUT2 #(
		.INIT('h8)
	) name17424 (
		_w27877_,
		_w27878_,
		_w27936_
	);
	LUT2 #(
		.INIT('h8)
	) name17425 (
		_w27875_,
		_w27876_,
		_w27937_
	);
	LUT2 #(
		.INIT('h8)
	) name17426 (
		_w27873_,
		_w27874_,
		_w27938_
	);
	LUT2 #(
		.INIT('h8)
	) name17427 (
		_w27871_,
		_w27872_,
		_w27939_
	);
	LUT2 #(
		.INIT('h8)
	) name17428 (
		_w27869_,
		_w27870_,
		_w27940_
	);
	LUT2 #(
		.INIT('h8)
	) name17429 (
		_w27867_,
		_w27868_,
		_w27941_
	);
	LUT2 #(
		.INIT('h8)
	) name17430 (
		_w27865_,
		_w27866_,
		_w27942_
	);
	LUT2 #(
		.INIT('h8)
	) name17431 (
		_w27863_,
		_w27864_,
		_w27943_
	);
	LUT2 #(
		.INIT('h8)
	) name17432 (
		_w27861_,
		_w27862_,
		_w27944_
	);
	LUT2 #(
		.INIT('h8)
	) name17433 (
		_w27859_,
		_w27860_,
		_w27945_
	);
	LUT2 #(
		.INIT('h8)
	) name17434 (
		_w27857_,
		_w27858_,
		_w27946_
	);
	LUT2 #(
		.INIT('h8)
	) name17435 (
		_w27855_,
		_w27856_,
		_w27947_
	);
	LUT2 #(
		.INIT('h8)
	) name17436 (
		_w27853_,
		_w27854_,
		_w27948_
	);
	LUT2 #(
		.INIT('h8)
	) name17437 (
		_w27947_,
		_w27948_,
		_w27949_
	);
	LUT2 #(
		.INIT('h8)
	) name17438 (
		_w27945_,
		_w27946_,
		_w27950_
	);
	LUT2 #(
		.INIT('h8)
	) name17439 (
		_w27943_,
		_w27944_,
		_w27951_
	);
	LUT2 #(
		.INIT('h8)
	) name17440 (
		_w27941_,
		_w27942_,
		_w27952_
	);
	LUT2 #(
		.INIT('h8)
	) name17441 (
		_w27939_,
		_w27940_,
		_w27953_
	);
	LUT2 #(
		.INIT('h8)
	) name17442 (
		_w27937_,
		_w27938_,
		_w27954_
	);
	LUT2 #(
		.INIT('h8)
	) name17443 (
		_w27935_,
		_w27936_,
		_w27955_
	);
	LUT2 #(
		.INIT('h8)
	) name17444 (
		_w27933_,
		_w27934_,
		_w27956_
	);
	LUT2 #(
		.INIT('h8)
	) name17445 (
		_w27931_,
		_w27932_,
		_w27957_
	);
	LUT2 #(
		.INIT('h8)
	) name17446 (
		_w27929_,
		_w27930_,
		_w27958_
	);
	LUT2 #(
		.INIT('h8)
	) name17447 (
		_w27927_,
		_w27928_,
		_w27959_
	);
	LUT2 #(
		.INIT('h8)
	) name17448 (
		_w27925_,
		_w27926_,
		_w27960_
	);
	LUT2 #(
		.INIT('h8)
	) name17449 (
		_w27923_,
		_w27924_,
		_w27961_
	);
	LUT2 #(
		.INIT('h8)
	) name17450 (
		_w27921_,
		_w27922_,
		_w27962_
	);
	LUT2 #(
		.INIT('h8)
	) name17451 (
		_w27919_,
		_w27920_,
		_w27963_
	);
	LUT2 #(
		.INIT('h8)
	) name17452 (
		_w27917_,
		_w27918_,
		_w27964_
	);
	LUT2 #(
		.INIT('h8)
	) name17453 (
		_w27963_,
		_w27964_,
		_w27965_
	);
	LUT2 #(
		.INIT('h8)
	) name17454 (
		_w27961_,
		_w27962_,
		_w27966_
	);
	LUT2 #(
		.INIT('h8)
	) name17455 (
		_w27959_,
		_w27960_,
		_w27967_
	);
	LUT2 #(
		.INIT('h8)
	) name17456 (
		_w27957_,
		_w27958_,
		_w27968_
	);
	LUT2 #(
		.INIT('h8)
	) name17457 (
		_w27955_,
		_w27956_,
		_w27969_
	);
	LUT2 #(
		.INIT('h8)
	) name17458 (
		_w27953_,
		_w27954_,
		_w27970_
	);
	LUT2 #(
		.INIT('h8)
	) name17459 (
		_w27951_,
		_w27952_,
		_w27971_
	);
	LUT2 #(
		.INIT('h8)
	) name17460 (
		_w27949_,
		_w27950_,
		_w27972_
	);
	LUT2 #(
		.INIT('h8)
	) name17461 (
		_w27971_,
		_w27972_,
		_w27973_
	);
	LUT2 #(
		.INIT('h8)
	) name17462 (
		_w27969_,
		_w27970_,
		_w27974_
	);
	LUT2 #(
		.INIT('h8)
	) name17463 (
		_w27967_,
		_w27968_,
		_w27975_
	);
	LUT2 #(
		.INIT('h8)
	) name17464 (
		_w27965_,
		_w27966_,
		_w27976_
	);
	LUT2 #(
		.INIT('h8)
	) name17465 (
		_w27975_,
		_w27976_,
		_w27977_
	);
	LUT2 #(
		.INIT('h8)
	) name17466 (
		_w27973_,
		_w27974_,
		_w27978_
	);
	LUT2 #(
		.INIT('h8)
	) name17467 (
		_w27977_,
		_w27978_,
		_w27979_
	);
	LUT2 #(
		.INIT('h1)
	) name17468 (
		wb_rst_i_pad,
		_w27979_,
		_w27980_
	);
	LUT2 #(
		.INIT('h1)
	) name17469 (
		_w22944_,
		_w27980_,
		_w27981_
	);
	LUT2 #(
		.INIT('h8)
	) name17470 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		_w22959_,
		_w27982_
	);
	LUT2 #(
		.INIT('h8)
	) name17471 (
		\ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 ,
		_w23499_,
		_w27983_
	);
	LUT2 #(
		.INIT('h8)
	) name17472 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		_w23501_,
		_w27984_
	);
	LUT2 #(
		.INIT('h8)
	) name17473 (
		\ethreg1_MIIRX_DATA_DataOut_reg[11]/NET0131 ,
		_w23507_,
		_w27985_
	);
	LUT2 #(
		.INIT('h8)
	) name17474 (
		\ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 ,
		_w22952_,
		_w27986_
	);
	LUT2 #(
		.INIT('h8)
	) name17475 (
		\ethreg1_PACKETLEN_1_DataOut_reg[3]/NET0131 ,
		_w22966_,
		_w27987_
	);
	LUT2 #(
		.INIT('h8)
	) name17476 (
		\ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 ,
		_w22956_,
		_w27988_
	);
	LUT2 #(
		.INIT('h8)
	) name17477 (
		\ethreg1_MODER_1_DataOut_reg[3]/NET0131 ,
		_w23519_,
		_w27989_
	);
	LUT2 #(
		.INIT('h8)
	) name17478 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		_w23513_,
		_w27990_
	);
	LUT2 #(
		.INIT('h8)
	) name17479 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 ,
		_w23522_,
		_w27991_
	);
	LUT2 #(
		.INIT('h1)
	) name17480 (
		_w27982_,
		_w27983_,
		_w27992_
	);
	LUT2 #(
		.INIT('h1)
	) name17481 (
		_w27984_,
		_w27985_,
		_w27993_
	);
	LUT2 #(
		.INIT('h1)
	) name17482 (
		_w27986_,
		_w27988_,
		_w27994_
	);
	LUT2 #(
		.INIT('h1)
	) name17483 (
		_w27989_,
		_w27990_,
		_w27995_
	);
	LUT2 #(
		.INIT('h4)
	) name17484 (
		_w27991_,
		_w27995_,
		_w27996_
	);
	LUT2 #(
		.INIT('h8)
	) name17485 (
		_w27993_,
		_w27994_,
		_w27997_
	);
	LUT2 #(
		.INIT('h8)
	) name17486 (
		_w22944_,
		_w27992_,
		_w27998_
	);
	LUT2 #(
		.INIT('h8)
	) name17487 (
		_w27997_,
		_w27998_,
		_w27999_
	);
	LUT2 #(
		.INIT('h4)
	) name17488 (
		_w27987_,
		_w27996_,
		_w28000_
	);
	LUT2 #(
		.INIT('h8)
	) name17489 (
		_w27999_,
		_w28000_,
		_w28001_
	);
	LUT2 #(
		.INIT('h1)
	) name17490 (
		_w27981_,
		_w28001_,
		_w28002_
	);
	LUT2 #(
		.INIT('h4)
	) name17491 (
		\wishbone_TxLength_reg[10]/NET0131 ,
		_w17290_,
		_w28003_
	);
	LUT2 #(
		.INIT('h1)
	) name17492 (
		\wishbone_TxLength_reg[11]/NET0131 ,
		_w28003_,
		_w28004_
	);
	LUT2 #(
		.INIT('h8)
	) name17493 (
		\wishbone_TxLength_reg[11]/NET0131 ,
		_w28003_,
		_w28005_
	);
	LUT2 #(
		.INIT('h2)
	) name17494 (
		_w18569_,
		_w28004_,
		_w28006_
	);
	LUT2 #(
		.INIT('h4)
	) name17495 (
		_w28005_,
		_w28006_,
		_w28007_
	);
	LUT2 #(
		.INIT('h1)
	) name17496 (
		_w20857_,
		_w28007_,
		_w28008_
	);
	LUT2 #(
		.INIT('h8)
	) name17497 (
		\wishbone_bd_ram_mem0_reg[8][2]/P0001 ,
		_w12920_,
		_w28009_
	);
	LUT2 #(
		.INIT('h8)
	) name17498 (
		\wishbone_bd_ram_mem0_reg[60][2]/P0001 ,
		_w13204_,
		_w28010_
	);
	LUT2 #(
		.INIT('h8)
	) name17499 (
		\wishbone_bd_ram_mem0_reg[42][2]/P0001 ,
		_w12842_,
		_w28011_
	);
	LUT2 #(
		.INIT('h8)
	) name17500 (
		\wishbone_bd_ram_mem0_reg[95][2]/P0001 ,
		_w12844_,
		_w28012_
	);
	LUT2 #(
		.INIT('h8)
	) name17501 (
		\wishbone_bd_ram_mem0_reg[80][2]/P0001 ,
		_w12689_,
		_w28013_
	);
	LUT2 #(
		.INIT('h8)
	) name17502 (
		\wishbone_bd_ram_mem0_reg[235][2]/P0001 ,
		_w12696_,
		_w28014_
	);
	LUT2 #(
		.INIT('h8)
	) name17503 (
		\wishbone_bd_ram_mem0_reg[135][2]/P0001 ,
		_w13124_,
		_w28015_
	);
	LUT2 #(
		.INIT('h8)
	) name17504 (
		\wishbone_bd_ram_mem0_reg[31][2]/P0001 ,
		_w13198_,
		_w28016_
	);
	LUT2 #(
		.INIT('h8)
	) name17505 (
		\wishbone_bd_ram_mem0_reg[121][2]/P0001 ,
		_w13078_,
		_w28017_
	);
	LUT2 #(
		.INIT('h8)
	) name17506 (
		\wishbone_bd_ram_mem0_reg[246][2]/P0001 ,
		_w13076_,
		_w28018_
	);
	LUT2 #(
		.INIT('h8)
	) name17507 (
		\wishbone_bd_ram_mem0_reg[200][2]/P0001 ,
		_w12988_,
		_w28019_
	);
	LUT2 #(
		.INIT('h8)
	) name17508 (
		\wishbone_bd_ram_mem0_reg[136][2]/P0001 ,
		_w13064_,
		_w28020_
	);
	LUT2 #(
		.INIT('h8)
	) name17509 (
		\wishbone_bd_ram_mem0_reg[16][2]/P0001 ,
		_w13140_,
		_w28021_
	);
	LUT2 #(
		.INIT('h8)
	) name17510 (
		\wishbone_bd_ram_mem0_reg[219][2]/P0001 ,
		_w12806_,
		_w28022_
	);
	LUT2 #(
		.INIT('h8)
	) name17511 (
		\wishbone_bd_ram_mem0_reg[38][2]/P0001 ,
		_w13182_,
		_w28023_
	);
	LUT2 #(
		.INIT('h8)
	) name17512 (
		\wishbone_bd_ram_mem0_reg[23][2]/P0001 ,
		_w13008_,
		_w28024_
	);
	LUT2 #(
		.INIT('h8)
	) name17513 (
		\wishbone_bd_ram_mem0_reg[212][2]/P0001 ,
		_w12796_,
		_w28025_
	);
	LUT2 #(
		.INIT('h8)
	) name17514 (
		\wishbone_bd_ram_mem0_reg[25][2]/P0001 ,
		_w13108_,
		_w28026_
	);
	LUT2 #(
		.INIT('h8)
	) name17515 (
		\wishbone_bd_ram_mem0_reg[85][2]/P0001 ,
		_w13216_,
		_w28027_
	);
	LUT2 #(
		.INIT('h8)
	) name17516 (
		\wishbone_bd_ram_mem0_reg[72][2]/P0001 ,
		_w12810_,
		_w28028_
	);
	LUT2 #(
		.INIT('h8)
	) name17517 (
		\wishbone_bd_ram_mem0_reg[157][2]/P0001 ,
		_w12926_,
		_w28029_
	);
	LUT2 #(
		.INIT('h8)
	) name17518 (
		\wishbone_bd_ram_mem0_reg[124][2]/P0001 ,
		_w13058_,
		_w28030_
	);
	LUT2 #(
		.INIT('h8)
	) name17519 (
		\wishbone_bd_ram_mem0_reg[113][2]/P0001 ,
		_w13026_,
		_w28031_
	);
	LUT2 #(
		.INIT('h8)
	) name17520 (
		\wishbone_bd_ram_mem0_reg[146][2]/P0001 ,
		_w13060_,
		_w28032_
	);
	LUT2 #(
		.INIT('h8)
	) name17521 (
		\wishbone_bd_ram_mem0_reg[188][2]/P0001 ,
		_w12948_,
		_w28033_
	);
	LUT2 #(
		.INIT('h8)
	) name17522 (
		\wishbone_bd_ram_mem0_reg[26][2]/P0001 ,
		_w12699_,
		_w28034_
	);
	LUT2 #(
		.INIT('h8)
	) name17523 (
		\wishbone_bd_ram_mem0_reg[108][2]/P0001 ,
		_w13156_,
		_w28035_
	);
	LUT2 #(
		.INIT('h8)
	) name17524 (
		\wishbone_bd_ram_mem0_reg[228][2]/P0001 ,
		_w12765_,
		_w28036_
	);
	LUT2 #(
		.INIT('h8)
	) name17525 (
		\wishbone_bd_ram_mem0_reg[196][2]/P0001 ,
		_w13090_,
		_w28037_
	);
	LUT2 #(
		.INIT('h8)
	) name17526 (
		\wishbone_bd_ram_mem0_reg[100][2]/P0001 ,
		_w12960_,
		_w28038_
	);
	LUT2 #(
		.INIT('h8)
	) name17527 (
		\wishbone_bd_ram_mem0_reg[198][2]/P0001 ,
		_w12832_,
		_w28039_
	);
	LUT2 #(
		.INIT('h8)
	) name17528 (
		\wishbone_bd_ram_mem0_reg[224][2]/P0001 ,
		_w12902_,
		_w28040_
	);
	LUT2 #(
		.INIT('h8)
	) name17529 (
		\wishbone_bd_ram_mem0_reg[150][2]/P0001 ,
		_w13136_,
		_w28041_
	);
	LUT2 #(
		.INIT('h8)
	) name17530 (
		\wishbone_bd_ram_mem0_reg[253][2]/P0001 ,
		_w13100_,
		_w28042_
	);
	LUT2 #(
		.INIT('h8)
	) name17531 (
		\wishbone_bd_ram_mem0_reg[159][2]/P0001 ,
		_w12774_,
		_w28043_
	);
	LUT2 #(
		.INIT('h8)
	) name17532 (
		\wishbone_bd_ram_mem0_reg[138][2]/P0001 ,
		_w12958_,
		_w28044_
	);
	LUT2 #(
		.INIT('h8)
	) name17533 (
		\wishbone_bd_ram_mem0_reg[3][2]/P0001 ,
		_w12866_,
		_w28045_
	);
	LUT2 #(
		.INIT('h8)
	) name17534 (
		\wishbone_bd_ram_mem0_reg[10][2]/P0001 ,
		_w13172_,
		_w28046_
	);
	LUT2 #(
		.INIT('h8)
	) name17535 (
		\wishbone_bd_ram_mem0_reg[12][2]/P0001 ,
		_w13118_,
		_w28047_
	);
	LUT2 #(
		.INIT('h8)
	) name17536 (
		\wishbone_bd_ram_mem0_reg[109][2]/P0001 ,
		_w12888_,
		_w28048_
	);
	LUT2 #(
		.INIT('h8)
	) name17537 (
		\wishbone_bd_ram_mem0_reg[191][2]/P0001 ,
		_w13034_,
		_w28049_
	);
	LUT2 #(
		.INIT('h8)
	) name17538 (
		\wishbone_bd_ram_mem0_reg[202][2]/P0001 ,
		_w12870_,
		_w28050_
	);
	LUT2 #(
		.INIT('h8)
	) name17539 (
		\wishbone_bd_ram_mem0_reg[180][2]/P0001 ,
		_w12791_,
		_w28051_
	);
	LUT2 #(
		.INIT('h8)
	) name17540 (
		\wishbone_bd_ram_mem0_reg[119][2]/P0001 ,
		_w13048_,
		_w28052_
	);
	LUT2 #(
		.INIT('h8)
	) name17541 (
		\wishbone_bd_ram_mem0_reg[175][2]/P0001 ,
		_w13126_,
		_w28053_
	);
	LUT2 #(
		.INIT('h8)
	) name17542 (
		\wishbone_bd_ram_mem0_reg[229][2]/P0001 ,
		_w12711_,
		_w28054_
	);
	LUT2 #(
		.INIT('h8)
	) name17543 (
		\wishbone_bd_ram_mem0_reg[51][2]/P0001 ,
		_w13024_,
		_w28055_
	);
	LUT2 #(
		.INIT('h8)
	) name17544 (
		\wishbone_bd_ram_mem0_reg[250][2]/P0001 ,
		_w13128_,
		_w28056_
	);
	LUT2 #(
		.INIT('h8)
	) name17545 (
		\wishbone_bd_ram_mem0_reg[242][2]/P0001 ,
		_w12932_,
		_w28057_
	);
	LUT2 #(
		.INIT('h8)
	) name17546 (
		\wishbone_bd_ram_mem0_reg[238][2]/P0001 ,
		_w13160_,
		_w28058_
	);
	LUT2 #(
		.INIT('h8)
	) name17547 (
		\wishbone_bd_ram_mem0_reg[223][2]/P0001 ,
		_w12838_,
		_w28059_
	);
	LUT2 #(
		.INIT('h8)
	) name17548 (
		\wishbone_bd_ram_mem0_reg[86][2]/P0001 ,
		_w12735_,
		_w28060_
	);
	LUT2 #(
		.INIT('h8)
	) name17549 (
		\wishbone_bd_ram_mem0_reg[76][2]/P0001 ,
		_w13184_,
		_w28061_
	);
	LUT2 #(
		.INIT('h8)
	) name17550 (
		\wishbone_bd_ram_mem0_reg[132][2]/P0001 ,
		_w12992_,
		_w28062_
	);
	LUT2 #(
		.INIT('h8)
	) name17551 (
		\wishbone_bd_ram_mem0_reg[102][2]/P0001 ,
		_w12685_,
		_w28063_
	);
	LUT2 #(
		.INIT('h8)
	) name17552 (
		\wishbone_bd_ram_mem0_reg[114][2]/P0001 ,
		_w13202_,
		_w28064_
	);
	LUT2 #(
		.INIT('h8)
	) name17553 (
		\wishbone_bd_ram_mem0_reg[192][2]/P0001 ,
		_w12938_,
		_w28065_
	);
	LUT2 #(
		.INIT('h8)
	) name17554 (
		\wishbone_bd_ram_mem0_reg[62][2]/P0001 ,
		_w12673_,
		_w28066_
	);
	LUT2 #(
		.INIT('h8)
	) name17555 (
		\wishbone_bd_ram_mem0_reg[137][2]/P0001 ,
		_w13168_,
		_w28067_
	);
	LUT2 #(
		.INIT('h8)
	) name17556 (
		\wishbone_bd_ram_mem0_reg[93][2]/P0001 ,
		_w13016_,
		_w28068_
	);
	LUT2 #(
		.INIT('h8)
	) name17557 (
		\wishbone_bd_ram_mem0_reg[221][2]/P0001 ,
		_w12802_,
		_w28069_
	);
	LUT2 #(
		.INIT('h8)
	) name17558 (
		\wishbone_bd_ram_mem0_reg[131][2]/P0001 ,
		_w12852_,
		_w28070_
	);
	LUT2 #(
		.INIT('h8)
	) name17559 (
		\wishbone_bd_ram_mem0_reg[222][2]/P0001 ,
		_w13094_,
		_w28071_
	);
	LUT2 #(
		.INIT('h8)
	) name17560 (
		\wishbone_bd_ram_mem0_reg[255][2]/P0001 ,
		_w13072_,
		_w28072_
	);
	LUT2 #(
		.INIT('h8)
	) name17561 (
		\wishbone_bd_ram_mem0_reg[233][2]/P0001 ,
		_w12836_,
		_w28073_
	);
	LUT2 #(
		.INIT('h8)
	) name17562 (
		\wishbone_bd_ram_mem0_reg[183][2]/P0001 ,
		_w12787_,
		_w28074_
	);
	LUT2 #(
		.INIT('h8)
	) name17563 (
		\wishbone_bd_ram_mem0_reg[70][2]/P0001 ,
		_w12840_,
		_w28075_
	);
	LUT2 #(
		.INIT('h8)
	) name17564 (
		\wishbone_bd_ram_mem0_reg[2][2]/P0001 ,
		_w13088_,
		_w28076_
	);
	LUT2 #(
		.INIT('h8)
	) name17565 (
		\wishbone_bd_ram_mem0_reg[104][2]/P0001 ,
		_w13148_,
		_w28077_
	);
	LUT2 #(
		.INIT('h8)
	) name17566 (
		\wishbone_bd_ram_mem0_reg[153][2]/P0001 ,
		_w12890_,
		_w28078_
	);
	LUT2 #(
		.INIT('h8)
	) name17567 (
		\wishbone_bd_ram_mem0_reg[44][2]/P0001 ,
		_w12896_,
		_w28079_
	);
	LUT2 #(
		.INIT('h8)
	) name17568 (
		\wishbone_bd_ram_mem0_reg[59][2]/P0001 ,
		_w12780_,
		_w28080_
	);
	LUT2 #(
		.INIT('h8)
	) name17569 (
		\wishbone_bd_ram_mem0_reg[1][2]/P0001 ,
		_w13014_,
		_w28081_
	);
	LUT2 #(
		.INIT('h8)
	) name17570 (
		\wishbone_bd_ram_mem0_reg[170][2]/P0001 ,
		_w13030_,
		_w28082_
	);
	LUT2 #(
		.INIT('h8)
	) name17571 (
		\wishbone_bd_ram_mem0_reg[103][2]/P0001 ,
		_w12846_,
		_w28083_
	);
	LUT2 #(
		.INIT('h8)
	) name17572 (
		\wishbone_bd_ram_mem0_reg[194][2]/P0001 ,
		_w12772_,
		_w28084_
	);
	LUT2 #(
		.INIT('h8)
	) name17573 (
		\wishbone_bd_ram_mem0_reg[166][2]/P0001 ,
		_w13040_,
		_w28085_
	);
	LUT2 #(
		.INIT('h8)
	) name17574 (
		\wishbone_bd_ram_mem0_reg[207][2]/P0001 ,
		_w13180_,
		_w28086_
	);
	LUT2 #(
		.INIT('h8)
	) name17575 (
		\wishbone_bd_ram_mem0_reg[178][2]/P0001 ,
		_w12886_,
		_w28087_
	);
	LUT2 #(
		.INIT('h8)
	) name17576 (
		\wishbone_bd_ram_mem0_reg[118][2]/P0001 ,
		_w12830_,
		_w28088_
	);
	LUT2 #(
		.INIT('h8)
	) name17577 (
		\wishbone_bd_ram_mem0_reg[91][2]/P0001 ,
		_w13074_,
		_w28089_
	);
	LUT2 #(
		.INIT('h8)
	) name17578 (
		\wishbone_bd_ram_mem0_reg[193][2]/P0001 ,
		_w13056_,
		_w28090_
	);
	LUT2 #(
		.INIT('h8)
	) name17579 (
		\wishbone_bd_ram_mem0_reg[160][2]/P0001 ,
		_w12872_,
		_w28091_
	);
	LUT2 #(
		.INIT('h8)
	) name17580 (
		\wishbone_bd_ram_mem0_reg[236][2]/P0001 ,
		_w12731_,
		_w28092_
	);
	LUT2 #(
		.INIT('h8)
	) name17581 (
		\wishbone_bd_ram_mem0_reg[43][2]/P0001 ,
		_w13200_,
		_w28093_
	);
	LUT2 #(
		.INIT('h8)
	) name17582 (
		\wishbone_bd_ram_mem0_reg[13][2]/P0001 ,
		_w13178_,
		_w28094_
	);
	LUT2 #(
		.INIT('h8)
	) name17583 (
		\wishbone_bd_ram_mem0_reg[50][2]/P0001 ,
		_w13150_,
		_w28095_
	);
	LUT2 #(
		.INIT('h8)
	) name17584 (
		\wishbone_bd_ram_mem0_reg[87][2]/P0001 ,
		_w13154_,
		_w28096_
	);
	LUT2 #(
		.INIT('h8)
	) name17585 (
		\wishbone_bd_ram_mem0_reg[28][2]/P0001 ,
		_w13170_,
		_w28097_
	);
	LUT2 #(
		.INIT('h8)
	) name17586 (
		\wishbone_bd_ram_mem0_reg[248][2]/P0001 ,
		_w12789_,
		_w28098_
	);
	LUT2 #(
		.INIT('h8)
	) name17587 (
		\wishbone_bd_ram_mem0_reg[11][2]/P0001 ,
		_w13194_,
		_w28099_
	);
	LUT2 #(
		.INIT('h8)
	) name17588 (
		\wishbone_bd_ram_mem0_reg[231][2]/P0001 ,
		_w12856_,
		_w28100_
	);
	LUT2 #(
		.INIT('h8)
	) name17589 (
		\wishbone_bd_ram_mem0_reg[240][2]/P0001 ,
		_w12864_,
		_w28101_
	);
	LUT2 #(
		.INIT('h8)
	) name17590 (
		\wishbone_bd_ram_mem0_reg[179][2]/P0001 ,
		_w13050_,
		_w28102_
	);
	LUT2 #(
		.INIT('h8)
	) name17591 (
		\wishbone_bd_ram_mem0_reg[34][2]/P0001 ,
		_w12930_,
		_w28103_
	);
	LUT2 #(
		.INIT('h8)
	) name17592 (
		\wishbone_bd_ram_mem0_reg[186][2]/P0001 ,
		_w12783_,
		_w28104_
	);
	LUT2 #(
		.INIT('h8)
	) name17593 (
		\wishbone_bd_ram_mem0_reg[190][2]/P0001 ,
		_w12858_,
		_w28105_
	);
	LUT2 #(
		.INIT('h8)
	) name17594 (
		\wishbone_bd_ram_mem0_reg[140][2]/P0001 ,
		_w12894_,
		_w28106_
	);
	LUT2 #(
		.INIT('h8)
	) name17595 (
		\wishbone_bd_ram_mem0_reg[149][2]/P0001 ,
		_w12741_,
		_w28107_
	);
	LUT2 #(
		.INIT('h8)
	) name17596 (
		\wishbone_bd_ram_mem0_reg[24][2]/P0001 ,
		_w13084_,
		_w28108_
	);
	LUT2 #(
		.INIT('h8)
	) name17597 (
		\wishbone_bd_ram_mem0_reg[214][2]/P0001 ,
		_w12984_,
		_w28109_
	);
	LUT2 #(
		.INIT('h8)
	) name17598 (
		\wishbone_bd_ram_mem0_reg[174][2]/P0001 ,
		_w12972_,
		_w28110_
	);
	LUT2 #(
		.INIT('h8)
	) name17599 (
		\wishbone_bd_ram_mem0_reg[96][2]/P0001 ,
		_w12912_,
		_w28111_
	);
	LUT2 #(
		.INIT('h8)
	) name17600 (
		\wishbone_bd_ram_mem0_reg[189][2]/P0001 ,
		_w13042_,
		_w28112_
	);
	LUT2 #(
		.INIT('h8)
	) name17601 (
		\wishbone_bd_ram_mem0_reg[163][2]/P0001 ,
		_w12882_,
		_w28113_
	);
	LUT2 #(
		.INIT('h8)
	) name17602 (
		\wishbone_bd_ram_mem0_reg[73][2]/P0001 ,
		_w12918_,
		_w28114_
	);
	LUT2 #(
		.INIT('h8)
	) name17603 (
		\wishbone_bd_ram_mem0_reg[64][2]/P0001 ,
		_w12976_,
		_w28115_
	);
	LUT2 #(
		.INIT('h8)
	) name17604 (
		\wishbone_bd_ram_mem0_reg[145][2]/P0001 ,
		_w13106_,
		_w28116_
	);
	LUT2 #(
		.INIT('h8)
	) name17605 (
		\wishbone_bd_ram_mem0_reg[210][2]/P0001 ,
		_w12924_,
		_w28117_
	);
	LUT2 #(
		.INIT('h8)
	) name17606 (
		\wishbone_bd_ram_mem0_reg[47][2]/P0001 ,
		_w12904_,
		_w28118_
	);
	LUT2 #(
		.INIT('h8)
	) name17607 (
		\wishbone_bd_ram_mem0_reg[195][2]/P0001 ,
		_w13144_,
		_w28119_
	);
	LUT2 #(
		.INIT('h8)
	) name17608 (
		\wishbone_bd_ram_mem0_reg[39][2]/P0001 ,
		_w13018_,
		_w28120_
	);
	LUT2 #(
		.INIT('h8)
	) name17609 (
		\wishbone_bd_ram_mem0_reg[199][2]/P0001 ,
		_w12768_,
		_w28121_
	);
	LUT2 #(
		.INIT('h8)
	) name17610 (
		\wishbone_bd_ram_mem0_reg[164][2]/P0001 ,
		_w12876_,
		_w28122_
	);
	LUT2 #(
		.INIT('h8)
	) name17611 (
		\wishbone_bd_ram_mem0_reg[249][2]/P0001 ,
		_w12900_,
		_w28123_
	);
	LUT2 #(
		.INIT('h8)
	) name17612 (
		\wishbone_bd_ram_mem0_reg[98][2]/P0001 ,
		_w12816_,
		_w28124_
	);
	LUT2 #(
		.INIT('h8)
	) name17613 (
		\wishbone_bd_ram_mem0_reg[88][2]/P0001 ,
		_w12860_,
		_w28125_
	);
	LUT2 #(
		.INIT('h8)
	) name17614 (
		\wishbone_bd_ram_mem0_reg[82][2]/P0001 ,
		_w12942_,
		_w28126_
	);
	LUT2 #(
		.INIT('h8)
	) name17615 (
		\wishbone_bd_ram_mem0_reg[169][2]/P0001 ,
		_w12722_,
		_w28127_
	);
	LUT2 #(
		.INIT('h8)
	) name17616 (
		\wishbone_bd_ram_mem0_reg[84][2]/P0001 ,
		_w12934_,
		_w28128_
	);
	LUT2 #(
		.INIT('h8)
	) name17617 (
		\wishbone_bd_ram_mem0_reg[112][2]/P0001 ,
		_w12733_,
		_w28129_
	);
	LUT2 #(
		.INIT('h8)
	) name17618 (
		\wishbone_bd_ram_mem0_reg[245][2]/P0001 ,
		_w13022_,
		_w28130_
	);
	LUT2 #(
		.INIT('h8)
	) name17619 (
		\wishbone_bd_ram_mem0_reg[57][2]/P0001 ,
		_w13116_,
		_w28131_
	);
	LUT2 #(
		.INIT('h8)
	) name17620 (
		\wishbone_bd_ram_mem0_reg[206][2]/P0001 ,
		_w12954_,
		_w28132_
	);
	LUT2 #(
		.INIT('h8)
	) name17621 (
		\wishbone_bd_ram_mem0_reg[143][2]/P0001 ,
		_w12922_,
		_w28133_
	);
	LUT2 #(
		.INIT('h8)
	) name17622 (
		\wishbone_bd_ram_mem0_reg[7][2]/P0001 ,
		_w12728_,
		_w28134_
	);
	LUT2 #(
		.INIT('h8)
	) name17623 (
		\wishbone_bd_ram_mem0_reg[142][2]/P0001 ,
		_w12928_,
		_w28135_
	);
	LUT2 #(
		.INIT('h8)
	) name17624 (
		\wishbone_bd_ram_mem0_reg[237][2]/P0001 ,
		_w12990_,
		_w28136_
	);
	LUT2 #(
		.INIT('h8)
	) name17625 (
		\wishbone_bd_ram_mem0_reg[171][2]/P0001 ,
		_w12910_,
		_w28137_
	);
	LUT2 #(
		.INIT('h8)
	) name17626 (
		\wishbone_bd_ram_mem0_reg[156][2]/P0001 ,
		_w13190_,
		_w28138_
	);
	LUT2 #(
		.INIT('h8)
	) name17627 (
		\wishbone_bd_ram_mem0_reg[32][2]/P0001 ,
		_w13120_,
		_w28139_
	);
	LUT2 #(
		.INIT('h8)
	) name17628 (
		\wishbone_bd_ram_mem0_reg[35][2]/P0001 ,
		_w12703_,
		_w28140_
	);
	LUT2 #(
		.INIT('h8)
	) name17629 (
		\wishbone_bd_ram_mem0_reg[89][2]/P0001 ,
		_w12964_,
		_w28141_
	);
	LUT2 #(
		.INIT('h8)
	) name17630 (
		\wishbone_bd_ram_mem0_reg[74][2]/P0001 ,
		_w12812_,
		_w28142_
	);
	LUT2 #(
		.INIT('h8)
	) name17631 (
		\wishbone_bd_ram_mem0_reg[203][2]/P0001 ,
		_w13158_,
		_w28143_
	);
	LUT2 #(
		.INIT('h8)
	) name17632 (
		\wishbone_bd_ram_mem0_reg[90][2]/P0001 ,
		_w12978_,
		_w28144_
	);
	LUT2 #(
		.INIT('h8)
	) name17633 (
		\wishbone_bd_ram_mem0_reg[27][2]/P0001 ,
		_w12880_,
		_w28145_
	);
	LUT2 #(
		.INIT('h8)
	) name17634 (
		\wishbone_bd_ram_mem0_reg[77][2]/P0001 ,
		_w12982_,
		_w28146_
	);
	LUT2 #(
		.INIT('h8)
	) name17635 (
		\wishbone_bd_ram_mem0_reg[216][2]/P0001 ,
		_w13028_,
		_w28147_
	);
	LUT2 #(
		.INIT('h8)
	) name17636 (
		\wishbone_bd_ram_mem0_reg[167][2]/P0001 ,
		_w12986_,
		_w28148_
	);
	LUT2 #(
		.INIT('h8)
	) name17637 (
		\wishbone_bd_ram_mem0_reg[185][2]/P0001 ,
		_w12940_,
		_w28149_
	);
	LUT2 #(
		.INIT('h8)
	) name17638 (
		\wishbone_bd_ram_mem0_reg[110][2]/P0001 ,
		_w13046_,
		_w28150_
	);
	LUT2 #(
		.INIT('h8)
	) name17639 (
		\wishbone_bd_ram_mem0_reg[232][2]/P0001 ,
		_w12758_,
		_w28151_
	);
	LUT2 #(
		.INIT('h8)
	) name17640 (
		\wishbone_bd_ram_mem0_reg[61][2]/P0001 ,
		_w12725_,
		_w28152_
	);
	LUT2 #(
		.INIT('h8)
	) name17641 (
		\wishbone_bd_ram_mem0_reg[107][2]/P0001 ,
		_w12749_,
		_w28153_
	);
	LUT2 #(
		.INIT('h8)
	) name17642 (
		\wishbone_bd_ram_mem0_reg[101][2]/P0001 ,
		_w13192_,
		_w28154_
	);
	LUT2 #(
		.INIT('h8)
	) name17643 (
		\wishbone_bd_ram_mem0_reg[184][2]/P0001 ,
		_w13062_,
		_w28155_
	);
	LUT2 #(
		.INIT('h8)
	) name17644 (
		\wishbone_bd_ram_mem0_reg[215][2]/P0001 ,
		_w12974_,
		_w28156_
	);
	LUT2 #(
		.INIT('h8)
	) name17645 (
		\wishbone_bd_ram_mem0_reg[134][2]/P0001 ,
		_w12763_,
		_w28157_
	);
	LUT2 #(
		.INIT('h8)
	) name17646 (
		\wishbone_bd_ram_mem0_reg[111][2]/P0001 ,
		_w12744_,
		_w28158_
	);
	LUT2 #(
		.INIT('h8)
	) name17647 (
		\wishbone_bd_ram_mem0_reg[129][2]/P0001 ,
		_w12776_,
		_w28159_
	);
	LUT2 #(
		.INIT('h8)
	) name17648 (
		\wishbone_bd_ram_mem0_reg[92][2]/P0001 ,
		_w13010_,
		_w28160_
	);
	LUT2 #(
		.INIT('h8)
	) name17649 (
		\wishbone_bd_ram_mem0_reg[46][2]/P0001 ,
		_w12884_,
		_w28161_
	);
	LUT2 #(
		.INIT('h8)
	) name17650 (
		\wishbone_bd_ram_mem0_reg[4][2]/P0001 ,
		_w12666_,
		_w28162_
	);
	LUT2 #(
		.INIT('h8)
	) name17651 (
		\wishbone_bd_ram_mem0_reg[168][2]/P0001 ,
		_w13208_,
		_w28163_
	);
	LUT2 #(
		.INIT('h8)
	) name17652 (
		\wishbone_bd_ram_mem0_reg[56][2]/P0001 ,
		_w12778_,
		_w28164_
	);
	LUT2 #(
		.INIT('h8)
	) name17653 (
		\wishbone_bd_ram_mem0_reg[99][2]/P0001 ,
		_w13038_,
		_w28165_
	);
	LUT2 #(
		.INIT('h8)
	) name17654 (
		\wishbone_bd_ram_mem0_reg[213][2]/P0001 ,
		_w13002_,
		_w28166_
	);
	LUT2 #(
		.INIT('h8)
	) name17655 (
		\wishbone_bd_ram_mem0_reg[41][2]/P0001 ,
		_w13052_,
		_w28167_
	);
	LUT2 #(
		.INIT('h8)
	) name17656 (
		\wishbone_bd_ram_mem0_reg[220][2]/P0001 ,
		_w13066_,
		_w28168_
	);
	LUT2 #(
		.INIT('h8)
	) name17657 (
		\wishbone_bd_ram_mem0_reg[53][2]/P0001 ,
		_w13020_,
		_w28169_
	);
	LUT2 #(
		.INIT('h8)
	) name17658 (
		\wishbone_bd_ram_mem0_reg[49][2]/P0001 ,
		_w12994_,
		_w28170_
	);
	LUT2 #(
		.INIT('h8)
	) name17659 (
		\wishbone_bd_ram_mem0_reg[117][2]/P0001 ,
		_w12715_,
		_w28171_
	);
	LUT2 #(
		.INIT('h8)
	) name17660 (
		\wishbone_bd_ram_mem0_reg[177][2]/P0001 ,
		_w12996_,
		_w28172_
	);
	LUT2 #(
		.INIT('h8)
	) name17661 (
		\wishbone_bd_ram_mem0_reg[125][2]/P0001 ,
		_w12956_,
		_w28173_
	);
	LUT2 #(
		.INIT('h8)
	) name17662 (
		\wishbone_bd_ram_mem0_reg[45][2]/P0001 ,
		_w12908_,
		_w28174_
	);
	LUT2 #(
		.INIT('h8)
	) name17663 (
		\wishbone_bd_ram_mem0_reg[106][2]/P0001 ,
		_w12713_,
		_w28175_
	);
	LUT2 #(
		.INIT('h8)
	) name17664 (
		\wishbone_bd_ram_mem0_reg[130][2]/P0001 ,
		_w12914_,
		_w28176_
	);
	LUT2 #(
		.INIT('h8)
	) name17665 (
		\wishbone_bd_ram_mem0_reg[48][2]/P0001 ,
		_w12970_,
		_w28177_
	);
	LUT2 #(
		.INIT('h8)
	) name17666 (
		\wishbone_bd_ram_mem0_reg[154][2]/P0001 ,
		_w12962_,
		_w28178_
	);
	LUT2 #(
		.INIT('h8)
	) name17667 (
		\wishbone_bd_ram_mem0_reg[0][2]/P0001 ,
		_w12717_,
		_w28179_
	);
	LUT2 #(
		.INIT('h8)
	) name17668 (
		\wishbone_bd_ram_mem0_reg[243][2]/P0001 ,
		_w12804_,
		_w28180_
	);
	LUT2 #(
		.INIT('h8)
	) name17669 (
		\wishbone_bd_ram_mem0_reg[36][2]/P0001 ,
		_w12800_,
		_w28181_
	);
	LUT2 #(
		.INIT('h8)
	) name17670 (
		\wishbone_bd_ram_mem0_reg[251][2]/P0001 ,
		_w13054_,
		_w28182_
	);
	LUT2 #(
		.INIT('h8)
	) name17671 (
		\wishbone_bd_ram_mem0_reg[241][2]/P0001 ,
		_w13006_,
		_w28183_
	);
	LUT2 #(
		.INIT('h8)
	) name17672 (
		\wishbone_bd_ram_mem0_reg[97][2]/P0001 ,
		_w13096_,
		_w28184_
	);
	LUT2 #(
		.INIT('h8)
	) name17673 (
		\wishbone_bd_ram_mem0_reg[19][2]/P0001 ,
		_w13012_,
		_w28185_
	);
	LUT2 #(
		.INIT('h8)
	) name17674 (
		\wishbone_bd_ram_mem0_reg[37][2]/P0001 ,
		_w13102_,
		_w28186_
	);
	LUT2 #(
		.INIT('h8)
	) name17675 (
		\wishbone_bd_ram_mem0_reg[123][2]/P0001 ,
		_w13114_,
		_w28187_
	);
	LUT2 #(
		.INIT('h8)
	) name17676 (
		\wishbone_bd_ram_mem0_reg[244][2]/P0001 ,
		_w12747_,
		_w28188_
	);
	LUT2 #(
		.INIT('h8)
	) name17677 (
		\wishbone_bd_ram_mem0_reg[247][2]/P0001 ,
		_w12818_,
		_w28189_
	);
	LUT2 #(
		.INIT('h8)
	) name17678 (
		\wishbone_bd_ram_mem0_reg[58][2]/P0001 ,
		_w13070_,
		_w28190_
	);
	LUT2 #(
		.INIT('h8)
	) name17679 (
		\wishbone_bd_ram_mem0_reg[197][2]/P0001 ,
		_w12834_,
		_w28191_
	);
	LUT2 #(
		.INIT('h8)
	) name17680 (
		\wishbone_bd_ram_mem0_reg[234][2]/P0001 ,
		_w13214_,
		_w28192_
	);
	LUT2 #(
		.INIT('h8)
	) name17681 (
		\wishbone_bd_ram_mem0_reg[254][2]/P0001 ,
		_w12892_,
		_w28193_
	);
	LUT2 #(
		.INIT('h8)
	) name17682 (
		\wishbone_bd_ram_mem0_reg[230][2]/P0001 ,
		_w13036_,
		_w28194_
	);
	LUT2 #(
		.INIT('h8)
	) name17683 (
		\wishbone_bd_ram_mem0_reg[227][2]/P0001 ,
		_w12936_,
		_w28195_
	);
	LUT2 #(
		.INIT('h8)
	) name17684 (
		\wishbone_bd_ram_mem0_reg[52][2]/P0001 ,
		_w13082_,
		_w28196_
	);
	LUT2 #(
		.INIT('h8)
	) name17685 (
		\wishbone_bd_ram_mem0_reg[79][2]/P0001 ,
		_w13212_,
		_w28197_
	);
	LUT2 #(
		.INIT('h8)
	) name17686 (
		\wishbone_bd_ram_mem0_reg[71][2]/P0001 ,
		_w12798_,
		_w28198_
	);
	LUT2 #(
		.INIT('h8)
	) name17687 (
		\wishbone_bd_ram_mem0_reg[30][2]/P0001 ,
		_w13104_,
		_w28199_
	);
	LUT2 #(
		.INIT('h8)
	) name17688 (
		\wishbone_bd_ram_mem0_reg[133][2]/P0001 ,
		_w12761_,
		_w28200_
	);
	LUT2 #(
		.INIT('h8)
	) name17689 (
		\wishbone_bd_ram_mem0_reg[226][2]/P0001 ,
		_w13138_,
		_w28201_
	);
	LUT2 #(
		.INIT('h8)
	) name17690 (
		\wishbone_bd_ram_mem0_reg[139][2]/P0001 ,
		_w12814_,
		_w28202_
	);
	LUT2 #(
		.INIT('h8)
	) name17691 (
		\wishbone_bd_ram_mem0_reg[105][2]/P0001 ,
		_w12751_,
		_w28203_
	);
	LUT2 #(
		.INIT('h8)
	) name17692 (
		\wishbone_bd_ram_mem0_reg[162][2]/P0001 ,
		_w13098_,
		_w28204_
	);
	LUT2 #(
		.INIT('h8)
	) name17693 (
		\wishbone_bd_ram_mem0_reg[252][2]/P0001 ,
		_w13080_,
		_w28205_
	);
	LUT2 #(
		.INIT('h8)
	) name17694 (
		\wishbone_bd_ram_mem0_reg[152][2]/P0001 ,
		_w12966_,
		_w28206_
	);
	LUT2 #(
		.INIT('h8)
	) name17695 (
		\wishbone_bd_ram_mem0_reg[5][2]/P0001 ,
		_w12878_,
		_w28207_
	);
	LUT2 #(
		.INIT('h8)
	) name17696 (
		\wishbone_bd_ram_mem0_reg[120][2]/P0001 ,
		_w12707_,
		_w28208_
	);
	LUT2 #(
		.INIT('h8)
	) name17697 (
		\wishbone_bd_ram_mem0_reg[66][2]/P0001 ,
		_w12824_,
		_w28209_
	);
	LUT2 #(
		.INIT('h8)
	) name17698 (
		\wishbone_bd_ram_mem0_reg[55][2]/P0001 ,
		_w12785_,
		_w28210_
	);
	LUT2 #(
		.INIT('h8)
	) name17699 (
		\wishbone_bd_ram_mem0_reg[15][2]/P0001 ,
		_w13210_,
		_w28211_
	);
	LUT2 #(
		.INIT('h8)
	) name17700 (
		\wishbone_bd_ram_mem0_reg[116][2]/P0001 ,
		_w12998_,
		_w28212_
	);
	LUT2 #(
		.INIT('h8)
	) name17701 (
		\wishbone_bd_ram_mem0_reg[161][2]/P0001 ,
		_w12754_,
		_w28213_
	);
	LUT2 #(
		.INIT('h8)
	) name17702 (
		\wishbone_bd_ram_mem0_reg[40][2]/P0001 ,
		_w13132_,
		_w28214_
	);
	LUT2 #(
		.INIT('h8)
	) name17703 (
		\wishbone_bd_ram_mem0_reg[14][2]/P0001 ,
		_w13086_,
		_w28215_
	);
	LUT2 #(
		.INIT('h8)
	) name17704 (
		\wishbone_bd_ram_mem0_reg[6][2]/P0001 ,
		_w12968_,
		_w28216_
	);
	LUT2 #(
		.INIT('h8)
	) name17705 (
		\wishbone_bd_ram_mem0_reg[20][2]/P0001 ,
		_w13174_,
		_w28217_
	);
	LUT2 #(
		.INIT('h8)
	) name17706 (
		\wishbone_bd_ram_mem0_reg[67][2]/P0001 ,
		_w13134_,
		_w28218_
	);
	LUT2 #(
		.INIT('h8)
	) name17707 (
		\wishbone_bd_ram_mem0_reg[181][2]/P0001 ,
		_w12828_,
		_w28219_
	);
	LUT2 #(
		.INIT('h8)
	) name17708 (
		\wishbone_bd_ram_mem0_reg[155][2]/P0001 ,
		_w13122_,
		_w28220_
	);
	LUT2 #(
		.INIT('h8)
	) name17709 (
		\wishbone_bd_ram_mem0_reg[9][2]/P0001 ,
		_w12808_,
		_w28221_
	);
	LUT2 #(
		.INIT('h8)
	) name17710 (
		\wishbone_bd_ram_mem0_reg[69][2]/P0001 ,
		_w12738_,
		_w28222_
	);
	LUT2 #(
		.INIT('h8)
	) name17711 (
		\wishbone_bd_ram_mem0_reg[218][2]/P0001 ,
		_w13206_,
		_w28223_
	);
	LUT2 #(
		.INIT('h8)
	) name17712 (
		\wishbone_bd_ram_mem0_reg[225][2]/P0001 ,
		_w13092_,
		_w28224_
	);
	LUT2 #(
		.INIT('h8)
	) name17713 (
		\wishbone_bd_ram_mem0_reg[128][2]/P0001 ,
		_w12793_,
		_w28225_
	);
	LUT2 #(
		.INIT('h8)
	) name17714 (
		\wishbone_bd_ram_mem0_reg[182][2]/P0001 ,
		_w12820_,
		_w28226_
	);
	LUT2 #(
		.INIT('h8)
	) name17715 (
		\wishbone_bd_ram_mem0_reg[158][2]/P0001 ,
		_w12898_,
		_w28227_
	);
	LUT2 #(
		.INIT('h8)
	) name17716 (
		\wishbone_bd_ram_mem0_reg[148][2]/P0001 ,
		_w13000_,
		_w28228_
	);
	LUT2 #(
		.INIT('h8)
	) name17717 (
		\wishbone_bd_ram_mem0_reg[144][2]/P0001 ,
		_w12756_,
		_w28229_
	);
	LUT2 #(
		.INIT('h8)
	) name17718 (
		\wishbone_bd_ram_mem0_reg[33][2]/P0001 ,
		_w12980_,
		_w28230_
	);
	LUT2 #(
		.INIT('h8)
	) name17719 (
		\wishbone_bd_ram_mem0_reg[209][2]/P0001 ,
		_w13152_,
		_w28231_
	);
	LUT2 #(
		.INIT('h8)
	) name17720 (
		\wishbone_bd_ram_mem0_reg[165][2]/P0001 ,
		_w13044_,
		_w28232_
	);
	LUT2 #(
		.INIT('h8)
	) name17721 (
		\wishbone_bd_ram_mem0_reg[17][2]/P0001 ,
		_w12848_,
		_w28233_
	);
	LUT2 #(
		.INIT('h8)
	) name17722 (
		\wishbone_bd_ram_mem0_reg[205][2]/P0001 ,
		_w13068_,
		_w28234_
	);
	LUT2 #(
		.INIT('h8)
	) name17723 (
		\wishbone_bd_ram_mem0_reg[187][2]/P0001 ,
		_w13196_,
		_w28235_
	);
	LUT2 #(
		.INIT('h8)
	) name17724 (
		\wishbone_bd_ram_mem0_reg[204][2]/P0001 ,
		_w13162_,
		_w28236_
	);
	LUT2 #(
		.INIT('h8)
	) name17725 (
		\wishbone_bd_ram_mem0_reg[126][2]/P0001 ,
		_w13218_,
		_w28237_
	);
	LUT2 #(
		.INIT('h8)
	) name17726 (
		\wishbone_bd_ram_mem0_reg[211][2]/P0001 ,
		_w13166_,
		_w28238_
	);
	LUT2 #(
		.INIT('h8)
	) name17727 (
		\wishbone_bd_ram_mem0_reg[63][2]/P0001 ,
		_w12850_,
		_w28239_
	);
	LUT2 #(
		.INIT('h8)
	) name17728 (
		\wishbone_bd_ram_mem0_reg[239][2]/P0001 ,
		_w12862_,
		_w28240_
	);
	LUT2 #(
		.INIT('h8)
	) name17729 (
		\wishbone_bd_ram_mem0_reg[122][2]/P0001 ,
		_w13130_,
		_w28241_
	);
	LUT2 #(
		.INIT('h8)
	) name17730 (
		\wishbone_bd_ram_mem0_reg[29][2]/P0001 ,
		_w12952_,
		_w28242_
	);
	LUT2 #(
		.INIT('h8)
	) name17731 (
		\wishbone_bd_ram_mem0_reg[65][2]/P0001 ,
		_w13176_,
		_w28243_
	);
	LUT2 #(
		.INIT('h8)
	) name17732 (
		\wishbone_bd_ram_mem0_reg[18][2]/P0001 ,
		_w12679_,
		_w28244_
	);
	LUT2 #(
		.INIT('h8)
	) name17733 (
		\wishbone_bd_ram_mem0_reg[201][2]/P0001 ,
		_w12822_,
		_w28245_
	);
	LUT2 #(
		.INIT('h8)
	) name17734 (
		\wishbone_bd_ram_mem0_reg[173][2]/P0001 ,
		_w12854_,
		_w28246_
	);
	LUT2 #(
		.INIT('h8)
	) name17735 (
		\wishbone_bd_ram_mem0_reg[75][2]/P0001 ,
		_w12826_,
		_w28247_
	);
	LUT2 #(
		.INIT('h8)
	) name17736 (
		\wishbone_bd_ram_mem0_reg[94][2]/P0001 ,
		_w13186_,
		_w28248_
	);
	LUT2 #(
		.INIT('h8)
	) name17737 (
		\wishbone_bd_ram_mem0_reg[217][2]/P0001 ,
		_w13188_,
		_w28249_
	);
	LUT2 #(
		.INIT('h8)
	) name17738 (
		\wishbone_bd_ram_mem0_reg[147][2]/P0001 ,
		_w13146_,
		_w28250_
	);
	LUT2 #(
		.INIT('h8)
	) name17739 (
		\wishbone_bd_ram_mem0_reg[208][2]/P0001 ,
		_w13032_,
		_w28251_
	);
	LUT2 #(
		.INIT('h8)
	) name17740 (
		\wishbone_bd_ram_mem0_reg[115][2]/P0001 ,
		_w13112_,
		_w28252_
	);
	LUT2 #(
		.INIT('h8)
	) name17741 (
		\wishbone_bd_ram_mem0_reg[172][2]/P0001 ,
		_w12944_,
		_w28253_
	);
	LUT2 #(
		.INIT('h8)
	) name17742 (
		\wishbone_bd_ram_mem0_reg[83][2]/P0001 ,
		_w12916_,
		_w28254_
	);
	LUT2 #(
		.INIT('h8)
	) name17743 (
		\wishbone_bd_ram_mem0_reg[21][2]/P0001 ,
		_w12906_,
		_w28255_
	);
	LUT2 #(
		.INIT('h8)
	) name17744 (
		\wishbone_bd_ram_mem0_reg[127][2]/P0001 ,
		_w13164_,
		_w28256_
	);
	LUT2 #(
		.INIT('h8)
	) name17745 (
		\wishbone_bd_ram_mem0_reg[141][2]/P0001 ,
		_w13004_,
		_w28257_
	);
	LUT2 #(
		.INIT('h8)
	) name17746 (
		\wishbone_bd_ram_mem0_reg[54][2]/P0001 ,
		_w12770_,
		_w28258_
	);
	LUT2 #(
		.INIT('h8)
	) name17747 (
		\wishbone_bd_ram_mem0_reg[81][2]/P0001 ,
		_w12950_,
		_w28259_
	);
	LUT2 #(
		.INIT('h8)
	) name17748 (
		\wishbone_bd_ram_mem0_reg[22][2]/P0001 ,
		_w13110_,
		_w28260_
	);
	LUT2 #(
		.INIT('h8)
	) name17749 (
		\wishbone_bd_ram_mem0_reg[68][2]/P0001 ,
		_w12946_,
		_w28261_
	);
	LUT2 #(
		.INIT('h8)
	) name17750 (
		\wishbone_bd_ram_mem0_reg[176][2]/P0001 ,
		_w12868_,
		_w28262_
	);
	LUT2 #(
		.INIT('h8)
	) name17751 (
		\wishbone_bd_ram_mem0_reg[78][2]/P0001 ,
		_w12874_,
		_w28263_
	);
	LUT2 #(
		.INIT('h8)
	) name17752 (
		\wishbone_bd_ram_mem0_reg[151][2]/P0001 ,
		_w13142_,
		_w28264_
	);
	LUT2 #(
		.INIT('h1)
	) name17753 (
		_w28009_,
		_w28010_,
		_w28265_
	);
	LUT2 #(
		.INIT('h1)
	) name17754 (
		_w28011_,
		_w28012_,
		_w28266_
	);
	LUT2 #(
		.INIT('h1)
	) name17755 (
		_w28013_,
		_w28014_,
		_w28267_
	);
	LUT2 #(
		.INIT('h1)
	) name17756 (
		_w28015_,
		_w28016_,
		_w28268_
	);
	LUT2 #(
		.INIT('h1)
	) name17757 (
		_w28017_,
		_w28018_,
		_w28269_
	);
	LUT2 #(
		.INIT('h1)
	) name17758 (
		_w28019_,
		_w28020_,
		_w28270_
	);
	LUT2 #(
		.INIT('h1)
	) name17759 (
		_w28021_,
		_w28022_,
		_w28271_
	);
	LUT2 #(
		.INIT('h1)
	) name17760 (
		_w28023_,
		_w28024_,
		_w28272_
	);
	LUT2 #(
		.INIT('h1)
	) name17761 (
		_w28025_,
		_w28026_,
		_w28273_
	);
	LUT2 #(
		.INIT('h1)
	) name17762 (
		_w28027_,
		_w28028_,
		_w28274_
	);
	LUT2 #(
		.INIT('h1)
	) name17763 (
		_w28029_,
		_w28030_,
		_w28275_
	);
	LUT2 #(
		.INIT('h1)
	) name17764 (
		_w28031_,
		_w28032_,
		_w28276_
	);
	LUT2 #(
		.INIT('h1)
	) name17765 (
		_w28033_,
		_w28034_,
		_w28277_
	);
	LUT2 #(
		.INIT('h1)
	) name17766 (
		_w28035_,
		_w28036_,
		_w28278_
	);
	LUT2 #(
		.INIT('h1)
	) name17767 (
		_w28037_,
		_w28038_,
		_w28279_
	);
	LUT2 #(
		.INIT('h1)
	) name17768 (
		_w28039_,
		_w28040_,
		_w28280_
	);
	LUT2 #(
		.INIT('h1)
	) name17769 (
		_w28041_,
		_w28042_,
		_w28281_
	);
	LUT2 #(
		.INIT('h1)
	) name17770 (
		_w28043_,
		_w28044_,
		_w28282_
	);
	LUT2 #(
		.INIT('h1)
	) name17771 (
		_w28045_,
		_w28046_,
		_w28283_
	);
	LUT2 #(
		.INIT('h1)
	) name17772 (
		_w28047_,
		_w28048_,
		_w28284_
	);
	LUT2 #(
		.INIT('h1)
	) name17773 (
		_w28049_,
		_w28050_,
		_w28285_
	);
	LUT2 #(
		.INIT('h1)
	) name17774 (
		_w28051_,
		_w28052_,
		_w28286_
	);
	LUT2 #(
		.INIT('h1)
	) name17775 (
		_w28053_,
		_w28054_,
		_w28287_
	);
	LUT2 #(
		.INIT('h1)
	) name17776 (
		_w28055_,
		_w28056_,
		_w28288_
	);
	LUT2 #(
		.INIT('h1)
	) name17777 (
		_w28057_,
		_w28058_,
		_w28289_
	);
	LUT2 #(
		.INIT('h1)
	) name17778 (
		_w28059_,
		_w28060_,
		_w28290_
	);
	LUT2 #(
		.INIT('h1)
	) name17779 (
		_w28061_,
		_w28062_,
		_w28291_
	);
	LUT2 #(
		.INIT('h1)
	) name17780 (
		_w28063_,
		_w28064_,
		_w28292_
	);
	LUT2 #(
		.INIT('h1)
	) name17781 (
		_w28065_,
		_w28066_,
		_w28293_
	);
	LUT2 #(
		.INIT('h1)
	) name17782 (
		_w28067_,
		_w28068_,
		_w28294_
	);
	LUT2 #(
		.INIT('h1)
	) name17783 (
		_w28069_,
		_w28070_,
		_w28295_
	);
	LUT2 #(
		.INIT('h1)
	) name17784 (
		_w28071_,
		_w28072_,
		_w28296_
	);
	LUT2 #(
		.INIT('h1)
	) name17785 (
		_w28073_,
		_w28074_,
		_w28297_
	);
	LUT2 #(
		.INIT('h1)
	) name17786 (
		_w28075_,
		_w28076_,
		_w28298_
	);
	LUT2 #(
		.INIT('h1)
	) name17787 (
		_w28077_,
		_w28078_,
		_w28299_
	);
	LUT2 #(
		.INIT('h1)
	) name17788 (
		_w28079_,
		_w28080_,
		_w28300_
	);
	LUT2 #(
		.INIT('h1)
	) name17789 (
		_w28081_,
		_w28082_,
		_w28301_
	);
	LUT2 #(
		.INIT('h1)
	) name17790 (
		_w28083_,
		_w28084_,
		_w28302_
	);
	LUT2 #(
		.INIT('h1)
	) name17791 (
		_w28085_,
		_w28086_,
		_w28303_
	);
	LUT2 #(
		.INIT('h1)
	) name17792 (
		_w28087_,
		_w28088_,
		_w28304_
	);
	LUT2 #(
		.INIT('h1)
	) name17793 (
		_w28089_,
		_w28090_,
		_w28305_
	);
	LUT2 #(
		.INIT('h1)
	) name17794 (
		_w28091_,
		_w28092_,
		_w28306_
	);
	LUT2 #(
		.INIT('h1)
	) name17795 (
		_w28093_,
		_w28094_,
		_w28307_
	);
	LUT2 #(
		.INIT('h1)
	) name17796 (
		_w28095_,
		_w28096_,
		_w28308_
	);
	LUT2 #(
		.INIT('h1)
	) name17797 (
		_w28097_,
		_w28098_,
		_w28309_
	);
	LUT2 #(
		.INIT('h1)
	) name17798 (
		_w28099_,
		_w28100_,
		_w28310_
	);
	LUT2 #(
		.INIT('h1)
	) name17799 (
		_w28101_,
		_w28102_,
		_w28311_
	);
	LUT2 #(
		.INIT('h1)
	) name17800 (
		_w28103_,
		_w28104_,
		_w28312_
	);
	LUT2 #(
		.INIT('h1)
	) name17801 (
		_w28105_,
		_w28106_,
		_w28313_
	);
	LUT2 #(
		.INIT('h1)
	) name17802 (
		_w28107_,
		_w28108_,
		_w28314_
	);
	LUT2 #(
		.INIT('h1)
	) name17803 (
		_w28109_,
		_w28110_,
		_w28315_
	);
	LUT2 #(
		.INIT('h1)
	) name17804 (
		_w28111_,
		_w28112_,
		_w28316_
	);
	LUT2 #(
		.INIT('h1)
	) name17805 (
		_w28113_,
		_w28114_,
		_w28317_
	);
	LUT2 #(
		.INIT('h1)
	) name17806 (
		_w28115_,
		_w28116_,
		_w28318_
	);
	LUT2 #(
		.INIT('h1)
	) name17807 (
		_w28117_,
		_w28118_,
		_w28319_
	);
	LUT2 #(
		.INIT('h1)
	) name17808 (
		_w28119_,
		_w28120_,
		_w28320_
	);
	LUT2 #(
		.INIT('h1)
	) name17809 (
		_w28121_,
		_w28122_,
		_w28321_
	);
	LUT2 #(
		.INIT('h1)
	) name17810 (
		_w28123_,
		_w28124_,
		_w28322_
	);
	LUT2 #(
		.INIT('h1)
	) name17811 (
		_w28125_,
		_w28126_,
		_w28323_
	);
	LUT2 #(
		.INIT('h1)
	) name17812 (
		_w28127_,
		_w28128_,
		_w28324_
	);
	LUT2 #(
		.INIT('h1)
	) name17813 (
		_w28129_,
		_w28130_,
		_w28325_
	);
	LUT2 #(
		.INIT('h1)
	) name17814 (
		_w28131_,
		_w28132_,
		_w28326_
	);
	LUT2 #(
		.INIT('h1)
	) name17815 (
		_w28133_,
		_w28134_,
		_w28327_
	);
	LUT2 #(
		.INIT('h1)
	) name17816 (
		_w28135_,
		_w28136_,
		_w28328_
	);
	LUT2 #(
		.INIT('h1)
	) name17817 (
		_w28137_,
		_w28138_,
		_w28329_
	);
	LUT2 #(
		.INIT('h1)
	) name17818 (
		_w28139_,
		_w28140_,
		_w28330_
	);
	LUT2 #(
		.INIT('h1)
	) name17819 (
		_w28141_,
		_w28142_,
		_w28331_
	);
	LUT2 #(
		.INIT('h1)
	) name17820 (
		_w28143_,
		_w28144_,
		_w28332_
	);
	LUT2 #(
		.INIT('h1)
	) name17821 (
		_w28145_,
		_w28146_,
		_w28333_
	);
	LUT2 #(
		.INIT('h1)
	) name17822 (
		_w28147_,
		_w28148_,
		_w28334_
	);
	LUT2 #(
		.INIT('h1)
	) name17823 (
		_w28149_,
		_w28150_,
		_w28335_
	);
	LUT2 #(
		.INIT('h1)
	) name17824 (
		_w28151_,
		_w28152_,
		_w28336_
	);
	LUT2 #(
		.INIT('h1)
	) name17825 (
		_w28153_,
		_w28154_,
		_w28337_
	);
	LUT2 #(
		.INIT('h1)
	) name17826 (
		_w28155_,
		_w28156_,
		_w28338_
	);
	LUT2 #(
		.INIT('h1)
	) name17827 (
		_w28157_,
		_w28158_,
		_w28339_
	);
	LUT2 #(
		.INIT('h1)
	) name17828 (
		_w28159_,
		_w28160_,
		_w28340_
	);
	LUT2 #(
		.INIT('h1)
	) name17829 (
		_w28161_,
		_w28162_,
		_w28341_
	);
	LUT2 #(
		.INIT('h1)
	) name17830 (
		_w28163_,
		_w28164_,
		_w28342_
	);
	LUT2 #(
		.INIT('h1)
	) name17831 (
		_w28165_,
		_w28166_,
		_w28343_
	);
	LUT2 #(
		.INIT('h1)
	) name17832 (
		_w28167_,
		_w28168_,
		_w28344_
	);
	LUT2 #(
		.INIT('h1)
	) name17833 (
		_w28169_,
		_w28170_,
		_w28345_
	);
	LUT2 #(
		.INIT('h1)
	) name17834 (
		_w28171_,
		_w28172_,
		_w28346_
	);
	LUT2 #(
		.INIT('h1)
	) name17835 (
		_w28173_,
		_w28174_,
		_w28347_
	);
	LUT2 #(
		.INIT('h1)
	) name17836 (
		_w28175_,
		_w28176_,
		_w28348_
	);
	LUT2 #(
		.INIT('h1)
	) name17837 (
		_w28177_,
		_w28178_,
		_w28349_
	);
	LUT2 #(
		.INIT('h1)
	) name17838 (
		_w28179_,
		_w28180_,
		_w28350_
	);
	LUT2 #(
		.INIT('h1)
	) name17839 (
		_w28181_,
		_w28182_,
		_w28351_
	);
	LUT2 #(
		.INIT('h1)
	) name17840 (
		_w28183_,
		_w28184_,
		_w28352_
	);
	LUT2 #(
		.INIT('h1)
	) name17841 (
		_w28185_,
		_w28186_,
		_w28353_
	);
	LUT2 #(
		.INIT('h1)
	) name17842 (
		_w28187_,
		_w28188_,
		_w28354_
	);
	LUT2 #(
		.INIT('h1)
	) name17843 (
		_w28189_,
		_w28190_,
		_w28355_
	);
	LUT2 #(
		.INIT('h1)
	) name17844 (
		_w28191_,
		_w28192_,
		_w28356_
	);
	LUT2 #(
		.INIT('h1)
	) name17845 (
		_w28193_,
		_w28194_,
		_w28357_
	);
	LUT2 #(
		.INIT('h1)
	) name17846 (
		_w28195_,
		_w28196_,
		_w28358_
	);
	LUT2 #(
		.INIT('h1)
	) name17847 (
		_w28197_,
		_w28198_,
		_w28359_
	);
	LUT2 #(
		.INIT('h1)
	) name17848 (
		_w28199_,
		_w28200_,
		_w28360_
	);
	LUT2 #(
		.INIT('h1)
	) name17849 (
		_w28201_,
		_w28202_,
		_w28361_
	);
	LUT2 #(
		.INIT('h1)
	) name17850 (
		_w28203_,
		_w28204_,
		_w28362_
	);
	LUT2 #(
		.INIT('h1)
	) name17851 (
		_w28205_,
		_w28206_,
		_w28363_
	);
	LUT2 #(
		.INIT('h1)
	) name17852 (
		_w28207_,
		_w28208_,
		_w28364_
	);
	LUT2 #(
		.INIT('h1)
	) name17853 (
		_w28209_,
		_w28210_,
		_w28365_
	);
	LUT2 #(
		.INIT('h1)
	) name17854 (
		_w28211_,
		_w28212_,
		_w28366_
	);
	LUT2 #(
		.INIT('h1)
	) name17855 (
		_w28213_,
		_w28214_,
		_w28367_
	);
	LUT2 #(
		.INIT('h1)
	) name17856 (
		_w28215_,
		_w28216_,
		_w28368_
	);
	LUT2 #(
		.INIT('h1)
	) name17857 (
		_w28217_,
		_w28218_,
		_w28369_
	);
	LUT2 #(
		.INIT('h1)
	) name17858 (
		_w28219_,
		_w28220_,
		_w28370_
	);
	LUT2 #(
		.INIT('h1)
	) name17859 (
		_w28221_,
		_w28222_,
		_w28371_
	);
	LUT2 #(
		.INIT('h1)
	) name17860 (
		_w28223_,
		_w28224_,
		_w28372_
	);
	LUT2 #(
		.INIT('h1)
	) name17861 (
		_w28225_,
		_w28226_,
		_w28373_
	);
	LUT2 #(
		.INIT('h1)
	) name17862 (
		_w28227_,
		_w28228_,
		_w28374_
	);
	LUT2 #(
		.INIT('h1)
	) name17863 (
		_w28229_,
		_w28230_,
		_w28375_
	);
	LUT2 #(
		.INIT('h1)
	) name17864 (
		_w28231_,
		_w28232_,
		_w28376_
	);
	LUT2 #(
		.INIT('h1)
	) name17865 (
		_w28233_,
		_w28234_,
		_w28377_
	);
	LUT2 #(
		.INIT('h1)
	) name17866 (
		_w28235_,
		_w28236_,
		_w28378_
	);
	LUT2 #(
		.INIT('h1)
	) name17867 (
		_w28237_,
		_w28238_,
		_w28379_
	);
	LUT2 #(
		.INIT('h1)
	) name17868 (
		_w28239_,
		_w28240_,
		_w28380_
	);
	LUT2 #(
		.INIT('h1)
	) name17869 (
		_w28241_,
		_w28242_,
		_w28381_
	);
	LUT2 #(
		.INIT('h1)
	) name17870 (
		_w28243_,
		_w28244_,
		_w28382_
	);
	LUT2 #(
		.INIT('h1)
	) name17871 (
		_w28245_,
		_w28246_,
		_w28383_
	);
	LUT2 #(
		.INIT('h1)
	) name17872 (
		_w28247_,
		_w28248_,
		_w28384_
	);
	LUT2 #(
		.INIT('h1)
	) name17873 (
		_w28249_,
		_w28250_,
		_w28385_
	);
	LUT2 #(
		.INIT('h1)
	) name17874 (
		_w28251_,
		_w28252_,
		_w28386_
	);
	LUT2 #(
		.INIT('h1)
	) name17875 (
		_w28253_,
		_w28254_,
		_w28387_
	);
	LUT2 #(
		.INIT('h1)
	) name17876 (
		_w28255_,
		_w28256_,
		_w28388_
	);
	LUT2 #(
		.INIT('h1)
	) name17877 (
		_w28257_,
		_w28258_,
		_w28389_
	);
	LUT2 #(
		.INIT('h1)
	) name17878 (
		_w28259_,
		_w28260_,
		_w28390_
	);
	LUT2 #(
		.INIT('h1)
	) name17879 (
		_w28261_,
		_w28262_,
		_w28391_
	);
	LUT2 #(
		.INIT('h1)
	) name17880 (
		_w28263_,
		_w28264_,
		_w28392_
	);
	LUT2 #(
		.INIT('h8)
	) name17881 (
		_w28391_,
		_w28392_,
		_w28393_
	);
	LUT2 #(
		.INIT('h8)
	) name17882 (
		_w28389_,
		_w28390_,
		_w28394_
	);
	LUT2 #(
		.INIT('h8)
	) name17883 (
		_w28387_,
		_w28388_,
		_w28395_
	);
	LUT2 #(
		.INIT('h8)
	) name17884 (
		_w28385_,
		_w28386_,
		_w28396_
	);
	LUT2 #(
		.INIT('h8)
	) name17885 (
		_w28383_,
		_w28384_,
		_w28397_
	);
	LUT2 #(
		.INIT('h8)
	) name17886 (
		_w28381_,
		_w28382_,
		_w28398_
	);
	LUT2 #(
		.INIT('h8)
	) name17887 (
		_w28379_,
		_w28380_,
		_w28399_
	);
	LUT2 #(
		.INIT('h8)
	) name17888 (
		_w28377_,
		_w28378_,
		_w28400_
	);
	LUT2 #(
		.INIT('h8)
	) name17889 (
		_w28375_,
		_w28376_,
		_w28401_
	);
	LUT2 #(
		.INIT('h8)
	) name17890 (
		_w28373_,
		_w28374_,
		_w28402_
	);
	LUT2 #(
		.INIT('h8)
	) name17891 (
		_w28371_,
		_w28372_,
		_w28403_
	);
	LUT2 #(
		.INIT('h8)
	) name17892 (
		_w28369_,
		_w28370_,
		_w28404_
	);
	LUT2 #(
		.INIT('h8)
	) name17893 (
		_w28367_,
		_w28368_,
		_w28405_
	);
	LUT2 #(
		.INIT('h8)
	) name17894 (
		_w28365_,
		_w28366_,
		_w28406_
	);
	LUT2 #(
		.INIT('h8)
	) name17895 (
		_w28363_,
		_w28364_,
		_w28407_
	);
	LUT2 #(
		.INIT('h8)
	) name17896 (
		_w28361_,
		_w28362_,
		_w28408_
	);
	LUT2 #(
		.INIT('h8)
	) name17897 (
		_w28359_,
		_w28360_,
		_w28409_
	);
	LUT2 #(
		.INIT('h8)
	) name17898 (
		_w28357_,
		_w28358_,
		_w28410_
	);
	LUT2 #(
		.INIT('h8)
	) name17899 (
		_w28355_,
		_w28356_,
		_w28411_
	);
	LUT2 #(
		.INIT('h8)
	) name17900 (
		_w28353_,
		_w28354_,
		_w28412_
	);
	LUT2 #(
		.INIT('h8)
	) name17901 (
		_w28351_,
		_w28352_,
		_w28413_
	);
	LUT2 #(
		.INIT('h8)
	) name17902 (
		_w28349_,
		_w28350_,
		_w28414_
	);
	LUT2 #(
		.INIT('h8)
	) name17903 (
		_w28347_,
		_w28348_,
		_w28415_
	);
	LUT2 #(
		.INIT('h8)
	) name17904 (
		_w28345_,
		_w28346_,
		_w28416_
	);
	LUT2 #(
		.INIT('h8)
	) name17905 (
		_w28343_,
		_w28344_,
		_w28417_
	);
	LUT2 #(
		.INIT('h8)
	) name17906 (
		_w28341_,
		_w28342_,
		_w28418_
	);
	LUT2 #(
		.INIT('h8)
	) name17907 (
		_w28339_,
		_w28340_,
		_w28419_
	);
	LUT2 #(
		.INIT('h8)
	) name17908 (
		_w28337_,
		_w28338_,
		_w28420_
	);
	LUT2 #(
		.INIT('h8)
	) name17909 (
		_w28335_,
		_w28336_,
		_w28421_
	);
	LUT2 #(
		.INIT('h8)
	) name17910 (
		_w28333_,
		_w28334_,
		_w28422_
	);
	LUT2 #(
		.INIT('h8)
	) name17911 (
		_w28331_,
		_w28332_,
		_w28423_
	);
	LUT2 #(
		.INIT('h8)
	) name17912 (
		_w28329_,
		_w28330_,
		_w28424_
	);
	LUT2 #(
		.INIT('h8)
	) name17913 (
		_w28327_,
		_w28328_,
		_w28425_
	);
	LUT2 #(
		.INIT('h8)
	) name17914 (
		_w28325_,
		_w28326_,
		_w28426_
	);
	LUT2 #(
		.INIT('h8)
	) name17915 (
		_w28323_,
		_w28324_,
		_w28427_
	);
	LUT2 #(
		.INIT('h8)
	) name17916 (
		_w28321_,
		_w28322_,
		_w28428_
	);
	LUT2 #(
		.INIT('h8)
	) name17917 (
		_w28319_,
		_w28320_,
		_w28429_
	);
	LUT2 #(
		.INIT('h8)
	) name17918 (
		_w28317_,
		_w28318_,
		_w28430_
	);
	LUT2 #(
		.INIT('h8)
	) name17919 (
		_w28315_,
		_w28316_,
		_w28431_
	);
	LUT2 #(
		.INIT('h8)
	) name17920 (
		_w28313_,
		_w28314_,
		_w28432_
	);
	LUT2 #(
		.INIT('h8)
	) name17921 (
		_w28311_,
		_w28312_,
		_w28433_
	);
	LUT2 #(
		.INIT('h8)
	) name17922 (
		_w28309_,
		_w28310_,
		_w28434_
	);
	LUT2 #(
		.INIT('h8)
	) name17923 (
		_w28307_,
		_w28308_,
		_w28435_
	);
	LUT2 #(
		.INIT('h8)
	) name17924 (
		_w28305_,
		_w28306_,
		_w28436_
	);
	LUT2 #(
		.INIT('h8)
	) name17925 (
		_w28303_,
		_w28304_,
		_w28437_
	);
	LUT2 #(
		.INIT('h8)
	) name17926 (
		_w28301_,
		_w28302_,
		_w28438_
	);
	LUT2 #(
		.INIT('h8)
	) name17927 (
		_w28299_,
		_w28300_,
		_w28439_
	);
	LUT2 #(
		.INIT('h8)
	) name17928 (
		_w28297_,
		_w28298_,
		_w28440_
	);
	LUT2 #(
		.INIT('h8)
	) name17929 (
		_w28295_,
		_w28296_,
		_w28441_
	);
	LUT2 #(
		.INIT('h8)
	) name17930 (
		_w28293_,
		_w28294_,
		_w28442_
	);
	LUT2 #(
		.INIT('h8)
	) name17931 (
		_w28291_,
		_w28292_,
		_w28443_
	);
	LUT2 #(
		.INIT('h8)
	) name17932 (
		_w28289_,
		_w28290_,
		_w28444_
	);
	LUT2 #(
		.INIT('h8)
	) name17933 (
		_w28287_,
		_w28288_,
		_w28445_
	);
	LUT2 #(
		.INIT('h8)
	) name17934 (
		_w28285_,
		_w28286_,
		_w28446_
	);
	LUT2 #(
		.INIT('h8)
	) name17935 (
		_w28283_,
		_w28284_,
		_w28447_
	);
	LUT2 #(
		.INIT('h8)
	) name17936 (
		_w28281_,
		_w28282_,
		_w28448_
	);
	LUT2 #(
		.INIT('h8)
	) name17937 (
		_w28279_,
		_w28280_,
		_w28449_
	);
	LUT2 #(
		.INIT('h8)
	) name17938 (
		_w28277_,
		_w28278_,
		_w28450_
	);
	LUT2 #(
		.INIT('h8)
	) name17939 (
		_w28275_,
		_w28276_,
		_w28451_
	);
	LUT2 #(
		.INIT('h8)
	) name17940 (
		_w28273_,
		_w28274_,
		_w28452_
	);
	LUT2 #(
		.INIT('h8)
	) name17941 (
		_w28271_,
		_w28272_,
		_w28453_
	);
	LUT2 #(
		.INIT('h8)
	) name17942 (
		_w28269_,
		_w28270_,
		_w28454_
	);
	LUT2 #(
		.INIT('h8)
	) name17943 (
		_w28267_,
		_w28268_,
		_w28455_
	);
	LUT2 #(
		.INIT('h8)
	) name17944 (
		_w28265_,
		_w28266_,
		_w28456_
	);
	LUT2 #(
		.INIT('h8)
	) name17945 (
		_w28455_,
		_w28456_,
		_w28457_
	);
	LUT2 #(
		.INIT('h8)
	) name17946 (
		_w28453_,
		_w28454_,
		_w28458_
	);
	LUT2 #(
		.INIT('h8)
	) name17947 (
		_w28451_,
		_w28452_,
		_w28459_
	);
	LUT2 #(
		.INIT('h8)
	) name17948 (
		_w28449_,
		_w28450_,
		_w28460_
	);
	LUT2 #(
		.INIT('h8)
	) name17949 (
		_w28447_,
		_w28448_,
		_w28461_
	);
	LUT2 #(
		.INIT('h8)
	) name17950 (
		_w28445_,
		_w28446_,
		_w28462_
	);
	LUT2 #(
		.INIT('h8)
	) name17951 (
		_w28443_,
		_w28444_,
		_w28463_
	);
	LUT2 #(
		.INIT('h8)
	) name17952 (
		_w28441_,
		_w28442_,
		_w28464_
	);
	LUT2 #(
		.INIT('h8)
	) name17953 (
		_w28439_,
		_w28440_,
		_w28465_
	);
	LUT2 #(
		.INIT('h8)
	) name17954 (
		_w28437_,
		_w28438_,
		_w28466_
	);
	LUT2 #(
		.INIT('h8)
	) name17955 (
		_w28435_,
		_w28436_,
		_w28467_
	);
	LUT2 #(
		.INIT('h8)
	) name17956 (
		_w28433_,
		_w28434_,
		_w28468_
	);
	LUT2 #(
		.INIT('h8)
	) name17957 (
		_w28431_,
		_w28432_,
		_w28469_
	);
	LUT2 #(
		.INIT('h8)
	) name17958 (
		_w28429_,
		_w28430_,
		_w28470_
	);
	LUT2 #(
		.INIT('h8)
	) name17959 (
		_w28427_,
		_w28428_,
		_w28471_
	);
	LUT2 #(
		.INIT('h8)
	) name17960 (
		_w28425_,
		_w28426_,
		_w28472_
	);
	LUT2 #(
		.INIT('h8)
	) name17961 (
		_w28423_,
		_w28424_,
		_w28473_
	);
	LUT2 #(
		.INIT('h8)
	) name17962 (
		_w28421_,
		_w28422_,
		_w28474_
	);
	LUT2 #(
		.INIT('h8)
	) name17963 (
		_w28419_,
		_w28420_,
		_w28475_
	);
	LUT2 #(
		.INIT('h8)
	) name17964 (
		_w28417_,
		_w28418_,
		_w28476_
	);
	LUT2 #(
		.INIT('h8)
	) name17965 (
		_w28415_,
		_w28416_,
		_w28477_
	);
	LUT2 #(
		.INIT('h8)
	) name17966 (
		_w28413_,
		_w28414_,
		_w28478_
	);
	LUT2 #(
		.INIT('h8)
	) name17967 (
		_w28411_,
		_w28412_,
		_w28479_
	);
	LUT2 #(
		.INIT('h8)
	) name17968 (
		_w28409_,
		_w28410_,
		_w28480_
	);
	LUT2 #(
		.INIT('h8)
	) name17969 (
		_w28407_,
		_w28408_,
		_w28481_
	);
	LUT2 #(
		.INIT('h8)
	) name17970 (
		_w28405_,
		_w28406_,
		_w28482_
	);
	LUT2 #(
		.INIT('h8)
	) name17971 (
		_w28403_,
		_w28404_,
		_w28483_
	);
	LUT2 #(
		.INIT('h8)
	) name17972 (
		_w28401_,
		_w28402_,
		_w28484_
	);
	LUT2 #(
		.INIT('h8)
	) name17973 (
		_w28399_,
		_w28400_,
		_w28485_
	);
	LUT2 #(
		.INIT('h8)
	) name17974 (
		_w28397_,
		_w28398_,
		_w28486_
	);
	LUT2 #(
		.INIT('h8)
	) name17975 (
		_w28395_,
		_w28396_,
		_w28487_
	);
	LUT2 #(
		.INIT('h8)
	) name17976 (
		_w28393_,
		_w28394_,
		_w28488_
	);
	LUT2 #(
		.INIT('h8)
	) name17977 (
		_w28487_,
		_w28488_,
		_w28489_
	);
	LUT2 #(
		.INIT('h8)
	) name17978 (
		_w28485_,
		_w28486_,
		_w28490_
	);
	LUT2 #(
		.INIT('h8)
	) name17979 (
		_w28483_,
		_w28484_,
		_w28491_
	);
	LUT2 #(
		.INIT('h8)
	) name17980 (
		_w28481_,
		_w28482_,
		_w28492_
	);
	LUT2 #(
		.INIT('h8)
	) name17981 (
		_w28479_,
		_w28480_,
		_w28493_
	);
	LUT2 #(
		.INIT('h8)
	) name17982 (
		_w28477_,
		_w28478_,
		_w28494_
	);
	LUT2 #(
		.INIT('h8)
	) name17983 (
		_w28475_,
		_w28476_,
		_w28495_
	);
	LUT2 #(
		.INIT('h8)
	) name17984 (
		_w28473_,
		_w28474_,
		_w28496_
	);
	LUT2 #(
		.INIT('h8)
	) name17985 (
		_w28471_,
		_w28472_,
		_w28497_
	);
	LUT2 #(
		.INIT('h8)
	) name17986 (
		_w28469_,
		_w28470_,
		_w28498_
	);
	LUT2 #(
		.INIT('h8)
	) name17987 (
		_w28467_,
		_w28468_,
		_w28499_
	);
	LUT2 #(
		.INIT('h8)
	) name17988 (
		_w28465_,
		_w28466_,
		_w28500_
	);
	LUT2 #(
		.INIT('h8)
	) name17989 (
		_w28463_,
		_w28464_,
		_w28501_
	);
	LUT2 #(
		.INIT('h8)
	) name17990 (
		_w28461_,
		_w28462_,
		_w28502_
	);
	LUT2 #(
		.INIT('h8)
	) name17991 (
		_w28459_,
		_w28460_,
		_w28503_
	);
	LUT2 #(
		.INIT('h8)
	) name17992 (
		_w28457_,
		_w28458_,
		_w28504_
	);
	LUT2 #(
		.INIT('h8)
	) name17993 (
		_w28503_,
		_w28504_,
		_w28505_
	);
	LUT2 #(
		.INIT('h8)
	) name17994 (
		_w28501_,
		_w28502_,
		_w28506_
	);
	LUT2 #(
		.INIT('h8)
	) name17995 (
		_w28499_,
		_w28500_,
		_w28507_
	);
	LUT2 #(
		.INIT('h8)
	) name17996 (
		_w28497_,
		_w28498_,
		_w28508_
	);
	LUT2 #(
		.INIT('h8)
	) name17997 (
		_w28495_,
		_w28496_,
		_w28509_
	);
	LUT2 #(
		.INIT('h8)
	) name17998 (
		_w28493_,
		_w28494_,
		_w28510_
	);
	LUT2 #(
		.INIT('h8)
	) name17999 (
		_w28491_,
		_w28492_,
		_w28511_
	);
	LUT2 #(
		.INIT('h8)
	) name18000 (
		_w28489_,
		_w28490_,
		_w28512_
	);
	LUT2 #(
		.INIT('h8)
	) name18001 (
		_w28511_,
		_w28512_,
		_w28513_
	);
	LUT2 #(
		.INIT('h8)
	) name18002 (
		_w28509_,
		_w28510_,
		_w28514_
	);
	LUT2 #(
		.INIT('h8)
	) name18003 (
		_w28507_,
		_w28508_,
		_w28515_
	);
	LUT2 #(
		.INIT('h8)
	) name18004 (
		_w28505_,
		_w28506_,
		_w28516_
	);
	LUT2 #(
		.INIT('h8)
	) name18005 (
		_w28515_,
		_w28516_,
		_w28517_
	);
	LUT2 #(
		.INIT('h8)
	) name18006 (
		_w28513_,
		_w28514_,
		_w28518_
	);
	LUT2 #(
		.INIT('h8)
	) name18007 (
		_w28517_,
		_w28518_,
		_w28519_
	);
	LUT2 #(
		.INIT('h1)
	) name18008 (
		wb_rst_i_pad,
		_w28519_,
		_w28520_
	);
	LUT2 #(
		.INIT('h1)
	) name18009 (
		_w22944_,
		_w28520_,
		_w28521_
	);
	LUT2 #(
		.INIT('h8)
	) name18010 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		_w22959_,
		_w28522_
	);
	LUT2 #(
		.INIT('h8)
	) name18011 (
		\ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 ,
		_w23499_,
		_w28523_
	);
	LUT2 #(
		.INIT('h8)
	) name18012 (
		\ethreg1_IPGR1_0_DataOut_reg[2]/NET0131 ,
		_w24710_,
		_w28524_
	);
	LUT2 #(
		.INIT('h8)
	) name18013 (
		_w23512_,
		_w24706_,
		_w28525_
	);
	LUT2 #(
		.INIT('h8)
	) name18014 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		_w28525_,
		_w28526_
	);
	LUT2 #(
		.INIT('h8)
	) name18015 (
		\ethreg1_PACKETLEN_0_DataOut_reg[2]/NET0131 ,
		_w22966_,
		_w28527_
	);
	LUT2 #(
		.INIT('h8)
	) name18016 (
		\ethreg1_MODER_0_DataOut_reg[2]/NET0131 ,
		_w23519_,
		_w28528_
	);
	LUT2 #(
		.INIT('h8)
	) name18017 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 ,
		_w23522_,
		_w28529_
	);
	LUT2 #(
		.INIT('h8)
	) name18018 (
		_w23521_,
		_w24716_,
		_w28530_
	);
	LUT2 #(
		.INIT('h8)
	) name18019 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		_w28530_,
		_w28531_
	);
	LUT2 #(
		.INIT('h8)
	) name18020 (
		\ethreg1_IPGR2_0_DataOut_reg[2]/NET0131 ,
		_w24724_,
		_w28532_
	);
	LUT2 #(
		.INIT('h8)
	) name18021 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 ,
		_w23513_,
		_w28533_
	);
	LUT2 #(
		.INIT('h8)
	) name18022 (
		_w23506_,
		_w23521_,
		_w28534_
	);
	LUT2 #(
		.INIT('h8)
	) name18023 (
		\miim1_Nvalid_reg/NET0131 ,
		_w28534_,
		_w28535_
	);
	LUT2 #(
		.INIT('h8)
	) name18024 (
		_w23506_,
		_w24706_,
		_w28536_
	);
	LUT2 #(
		.INIT('h8)
	) name18025 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		_w28536_,
		_w28537_
	);
	LUT2 #(
		.INIT('h8)
	) name18026 (
		\ethreg1_irq_rxb_reg/NET0131 ,
		_w24707_,
		_w28538_
	);
	LUT2 #(
		.INIT('h8)
	) name18027 (
		\ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 ,
		_w24722_,
		_w28539_
	);
	LUT2 #(
		.INIT('h8)
	) name18028 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		_w23501_,
		_w28540_
	);
	LUT2 #(
		.INIT('h8)
	) name18029 (
		\ethreg1_MIIRX_DATA_DataOut_reg[2]/NET0131 ,
		_w23507_,
		_w28541_
	);
	LUT2 #(
		.INIT('h8)
	) name18030 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		_w24713_,
		_w28542_
	);
	LUT2 #(
		.INIT('h8)
	) name18031 (
		\ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 ,
		_w22956_,
		_w28543_
	);
	LUT2 #(
		.INIT('h8)
	) name18032 (
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		_w24726_,
		_w28544_
	);
	LUT2 #(
		.INIT('h8)
	) name18033 (
		\ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 ,
		_w22952_,
		_w28545_
	);
	LUT2 #(
		.INIT('h8)
	) name18034 (
		\ethreg1_IPGT_0_DataOut_reg[2]/NET0131 ,
		_w24717_,
		_w28546_
	);
	LUT2 #(
		.INIT('h1)
	) name18035 (
		_w28522_,
		_w28523_,
		_w28547_
	);
	LUT2 #(
		.INIT('h1)
	) name18036 (
		_w28524_,
		_w28526_,
		_w28548_
	);
	LUT2 #(
		.INIT('h1)
	) name18037 (
		_w28528_,
		_w28529_,
		_w28549_
	);
	LUT2 #(
		.INIT('h1)
	) name18038 (
		_w28531_,
		_w28532_,
		_w28550_
	);
	LUT2 #(
		.INIT('h1)
	) name18039 (
		_w28533_,
		_w28535_,
		_w28551_
	);
	LUT2 #(
		.INIT('h1)
	) name18040 (
		_w28537_,
		_w28538_,
		_w28552_
	);
	LUT2 #(
		.INIT('h1)
	) name18041 (
		_w28539_,
		_w28540_,
		_w28553_
	);
	LUT2 #(
		.INIT('h1)
	) name18042 (
		_w28541_,
		_w28542_,
		_w28554_
	);
	LUT2 #(
		.INIT('h1)
	) name18043 (
		_w28543_,
		_w28544_,
		_w28555_
	);
	LUT2 #(
		.INIT('h1)
	) name18044 (
		_w28545_,
		_w28546_,
		_w28556_
	);
	LUT2 #(
		.INIT('h8)
	) name18045 (
		_w28555_,
		_w28556_,
		_w28557_
	);
	LUT2 #(
		.INIT('h8)
	) name18046 (
		_w28553_,
		_w28554_,
		_w28558_
	);
	LUT2 #(
		.INIT('h8)
	) name18047 (
		_w28551_,
		_w28552_,
		_w28559_
	);
	LUT2 #(
		.INIT('h8)
	) name18048 (
		_w28549_,
		_w28550_,
		_w28560_
	);
	LUT2 #(
		.INIT('h8)
	) name18049 (
		_w28547_,
		_w28548_,
		_w28561_
	);
	LUT2 #(
		.INIT('h8)
	) name18050 (
		_w22944_,
		_w28561_,
		_w28562_
	);
	LUT2 #(
		.INIT('h8)
	) name18051 (
		_w28559_,
		_w28560_,
		_w28563_
	);
	LUT2 #(
		.INIT('h8)
	) name18052 (
		_w28557_,
		_w28558_,
		_w28564_
	);
	LUT2 #(
		.INIT('h4)
	) name18053 (
		_w28527_,
		_w28564_,
		_w28565_
	);
	LUT2 #(
		.INIT('h8)
	) name18054 (
		_w28562_,
		_w28563_,
		_w28566_
	);
	LUT2 #(
		.INIT('h8)
	) name18055 (
		_w28565_,
		_w28566_,
		_w28567_
	);
	LUT2 #(
		.INIT('h1)
	) name18056 (
		_w28521_,
		_w28567_,
		_w28568_
	);
	LUT2 #(
		.INIT('h1)
	) name18057 (
		_w22944_,
		_w24094_,
		_w28569_
	);
	LUT2 #(
		.INIT('h8)
	) name18058 (
		\ethreg1_IPGT_0_DataOut_reg[0]/NET0131 ,
		_w24717_,
		_w28570_
	);
	LUT2 #(
		.INIT('h8)
	) name18059 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		_w22959_,
		_w28571_
	);
	LUT2 #(
		.INIT('h8)
	) name18060 (
		\ethreg1_IPGR1_0_DataOut_reg[0]/NET0131 ,
		_w24710_,
		_w28572_
	);
	LUT2 #(
		.INIT('h8)
	) name18061 (
		\ethreg1_MIIRX_DATA_DataOut_reg[0]/NET0131 ,
		_w23507_,
		_w28573_
	);
	LUT2 #(
		.INIT('h8)
	) name18062 (
		\ethreg1_PACKETLEN_0_DataOut_reg[0]/NET0131 ,
		_w22966_,
		_w28574_
	);
	LUT2 #(
		.INIT('h8)
	) name18063 (
		\ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 ,
		_w23499_,
		_w28575_
	);
	LUT2 #(
		.INIT('h8)
	) name18064 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		_w28525_,
		_w28576_
	);
	LUT2 #(
		.INIT('h8)
	) name18065 (
		\ethreg1_irq_txb_reg/NET0131 ,
		_w24707_,
		_w28577_
	);
	LUT2 #(
		.INIT('h8)
	) name18066 (
		\ethreg1_MIICOMMAND0_DataOut_reg[0]/NET0131 ,
		_w28536_,
		_w28578_
	);
	LUT2 #(
		.INIT('h8)
	) name18067 (
		\ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 ,
		_w22956_,
		_w28579_
	);
	LUT2 #(
		.INIT('h8)
	) name18068 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		_w23519_,
		_w28580_
	);
	LUT2 #(
		.INIT('h8)
	) name18069 (
		\ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 ,
		_w22952_,
		_w28581_
	);
	LUT2 #(
		.INIT('h8)
	) name18070 (
		\ethreg1_IPGR2_0_DataOut_reg[0]/NET0131 ,
		_w24724_,
		_w28582_
	);
	LUT2 #(
		.INIT('h8)
	) name18071 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 ,
		_w23513_,
		_w28583_
	);
	LUT2 #(
		.INIT('h8)
	) name18072 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		_w23501_,
		_w28584_
	);
	LUT2 #(
		.INIT('h8)
	) name18073 (
		\miim1_shftrg_LinkFail_reg/NET0131 ,
		_w28534_,
		_w28585_
	);
	LUT2 #(
		.INIT('h8)
	) name18074 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 ,
		_w23522_,
		_w28586_
	);
	LUT2 #(
		.INIT('h8)
	) name18075 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		_w28530_,
		_w28587_
	);
	LUT2 #(
		.INIT('h8)
	) name18076 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		_w24713_,
		_w28588_
	);
	LUT2 #(
		.INIT('h8)
	) name18077 (
		\ethreg1_MIIMODER_0_DataOut_reg[0]/NET0131 ,
		_w24726_,
		_w28589_
	);
	LUT2 #(
		.INIT('h8)
	) name18078 (
		\ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 ,
		_w24722_,
		_w28590_
	);
	LUT2 #(
		.INIT('h1)
	) name18079 (
		_w28570_,
		_w28571_,
		_w28591_
	);
	LUT2 #(
		.INIT('h1)
	) name18080 (
		_w28572_,
		_w28573_,
		_w28592_
	);
	LUT2 #(
		.INIT('h1)
	) name18081 (
		_w28575_,
		_w28576_,
		_w28593_
	);
	LUT2 #(
		.INIT('h1)
	) name18082 (
		_w28577_,
		_w28578_,
		_w28594_
	);
	LUT2 #(
		.INIT('h1)
	) name18083 (
		_w28579_,
		_w28580_,
		_w28595_
	);
	LUT2 #(
		.INIT('h1)
	) name18084 (
		_w28581_,
		_w28582_,
		_w28596_
	);
	LUT2 #(
		.INIT('h1)
	) name18085 (
		_w28583_,
		_w28584_,
		_w28597_
	);
	LUT2 #(
		.INIT('h1)
	) name18086 (
		_w28585_,
		_w28586_,
		_w28598_
	);
	LUT2 #(
		.INIT('h1)
	) name18087 (
		_w28587_,
		_w28588_,
		_w28599_
	);
	LUT2 #(
		.INIT('h1)
	) name18088 (
		_w28589_,
		_w28590_,
		_w28600_
	);
	LUT2 #(
		.INIT('h8)
	) name18089 (
		_w28599_,
		_w28600_,
		_w28601_
	);
	LUT2 #(
		.INIT('h8)
	) name18090 (
		_w28597_,
		_w28598_,
		_w28602_
	);
	LUT2 #(
		.INIT('h8)
	) name18091 (
		_w28595_,
		_w28596_,
		_w28603_
	);
	LUT2 #(
		.INIT('h8)
	) name18092 (
		_w28593_,
		_w28594_,
		_w28604_
	);
	LUT2 #(
		.INIT('h8)
	) name18093 (
		_w28591_,
		_w28592_,
		_w28605_
	);
	LUT2 #(
		.INIT('h8)
	) name18094 (
		_w22944_,
		_w28605_,
		_w28606_
	);
	LUT2 #(
		.INIT('h8)
	) name18095 (
		_w28603_,
		_w28604_,
		_w28607_
	);
	LUT2 #(
		.INIT('h8)
	) name18096 (
		_w28601_,
		_w28602_,
		_w28608_
	);
	LUT2 #(
		.INIT('h4)
	) name18097 (
		_w28574_,
		_w28608_,
		_w28609_
	);
	LUT2 #(
		.INIT('h8)
	) name18098 (
		_w28606_,
		_w28607_,
		_w28610_
	);
	LUT2 #(
		.INIT('h8)
	) name18099 (
		_w28609_,
		_w28610_,
		_w28611_
	);
	LUT2 #(
		.INIT('h1)
	) name18100 (
		_w28569_,
		_w28611_,
		_w28612_
	);
	LUT2 #(
		.INIT('h1)
	) name18101 (
		_w16210_,
		_w22944_,
		_w28613_
	);
	LUT2 #(
		.INIT('h8)
	) name18102 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		_w24713_,
		_w28614_
	);
	LUT2 #(
		.INIT('h8)
	) name18103 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		_w22959_,
		_w28615_
	);
	LUT2 #(
		.INIT('h8)
	) name18104 (
		\ethreg1_IPGR2_0_DataOut_reg[1]/NET0131 ,
		_w24724_,
		_w28616_
	);
	LUT2 #(
		.INIT('h8)
	) name18105 (
		\ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 ,
		_w22952_,
		_w28617_
	);
	LUT2 #(
		.INIT('h8)
	) name18106 (
		\ethreg1_PACKETLEN_0_DataOut_reg[1]/NET0131 ,
		_w22966_,
		_w28618_
	);
	LUT2 #(
		.INIT('h8)
	) name18107 (
		\ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 ,
		_w22956_,
		_w28619_
	);
	LUT2 #(
		.INIT('h8)
	) name18108 (
		\ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 ,
		_w23499_,
		_w28620_
	);
	LUT2 #(
		.INIT('h8)
	) name18109 (
		\ethreg1_MIIRX_DATA_DataOut_reg[1]/NET0131 ,
		_w23507_,
		_w28621_
	);
	LUT2 #(
		.INIT('h1)
	) name18110 (
		_w28534_,
		_w28536_,
		_w28622_
	);
	LUT2 #(
		.INIT('h2)
	) name18111 (
		\ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 ,
		_w28622_,
		_w28623_
	);
	LUT2 #(
		.INIT('h8)
	) name18112 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		_w24726_,
		_w28624_
	);
	LUT2 #(
		.INIT('h8)
	) name18113 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 ,
		_w23513_,
		_w28625_
	);
	LUT2 #(
		.INIT('h8)
	) name18114 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		_w23501_,
		_w28626_
	);
	LUT2 #(
		.INIT('h8)
	) name18115 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 ,
		_w23522_,
		_w28627_
	);
	LUT2 #(
		.INIT('h8)
	) name18116 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		_w28530_,
		_w28628_
	);
	LUT2 #(
		.INIT('h8)
	) name18117 (
		\ethreg1_irq_txe_reg/NET0131 ,
		_w24707_,
		_w28629_
	);
	LUT2 #(
		.INIT('h8)
	) name18118 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		_w28525_,
		_w28630_
	);
	LUT2 #(
		.INIT('h1)
	) name18119 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w28631_
	);
	LUT2 #(
		.INIT('h1)
	) name18120 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		\miim1_InProgress_q3_reg/NET0131 ,
		_w28632_
	);
	LUT2 #(
		.INIT('h1)
	) name18121 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_Nvalid_reg/NET0131 ,
		_w28633_
	);
	LUT2 #(
		.INIT('h1)
	) name18122 (
		\miim1_RStatStart_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w28634_
	);
	LUT2 #(
		.INIT('h8)
	) name18123 (
		_w28633_,
		_w28634_,
		_w28635_
	);
	LUT2 #(
		.INIT('h8)
	) name18124 (
		_w28631_,
		_w28632_,
		_w28636_
	);
	LUT2 #(
		.INIT('h8)
	) name18125 (
		_w28635_,
		_w28636_,
		_w28637_
	);
	LUT2 #(
		.INIT('h2)
	) name18126 (
		_w28534_,
		_w28637_,
		_w28638_
	);
	LUT2 #(
		.INIT('h8)
	) name18127 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		_w23519_,
		_w28639_
	);
	LUT2 #(
		.INIT('h8)
	) name18128 (
		\ethreg1_IPGR1_0_DataOut_reg[1]/NET0131 ,
		_w24710_,
		_w28640_
	);
	LUT2 #(
		.INIT('h8)
	) name18129 (
		\ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 ,
		_w24722_,
		_w28641_
	);
	LUT2 #(
		.INIT('h8)
	) name18130 (
		\ethreg1_IPGT_0_DataOut_reg[1]/NET0131 ,
		_w24717_,
		_w28642_
	);
	LUT2 #(
		.INIT('h1)
	) name18131 (
		_w28614_,
		_w28615_,
		_w28643_
	);
	LUT2 #(
		.INIT('h1)
	) name18132 (
		_w28616_,
		_w28617_,
		_w28644_
	);
	LUT2 #(
		.INIT('h1)
	) name18133 (
		_w28619_,
		_w28620_,
		_w28645_
	);
	LUT2 #(
		.INIT('h1)
	) name18134 (
		_w28621_,
		_w28624_,
		_w28646_
	);
	LUT2 #(
		.INIT('h1)
	) name18135 (
		_w28625_,
		_w28626_,
		_w28647_
	);
	LUT2 #(
		.INIT('h1)
	) name18136 (
		_w28627_,
		_w28628_,
		_w28648_
	);
	LUT2 #(
		.INIT('h1)
	) name18137 (
		_w28629_,
		_w28630_,
		_w28649_
	);
	LUT2 #(
		.INIT('h1)
	) name18138 (
		_w28638_,
		_w28639_,
		_w28650_
	);
	LUT2 #(
		.INIT('h1)
	) name18139 (
		_w28640_,
		_w28641_,
		_w28651_
	);
	LUT2 #(
		.INIT('h4)
	) name18140 (
		_w28642_,
		_w28651_,
		_w28652_
	);
	LUT2 #(
		.INIT('h8)
	) name18141 (
		_w28649_,
		_w28650_,
		_w28653_
	);
	LUT2 #(
		.INIT('h8)
	) name18142 (
		_w28647_,
		_w28648_,
		_w28654_
	);
	LUT2 #(
		.INIT('h8)
	) name18143 (
		_w28645_,
		_w28646_,
		_w28655_
	);
	LUT2 #(
		.INIT('h8)
	) name18144 (
		_w28643_,
		_w28644_,
		_w28656_
	);
	LUT2 #(
		.INIT('h2)
	) name18145 (
		_w22944_,
		_w28623_,
		_w28657_
	);
	LUT2 #(
		.INIT('h8)
	) name18146 (
		_w28656_,
		_w28657_,
		_w28658_
	);
	LUT2 #(
		.INIT('h8)
	) name18147 (
		_w28654_,
		_w28655_,
		_w28659_
	);
	LUT2 #(
		.INIT('h8)
	) name18148 (
		_w28652_,
		_w28653_,
		_w28660_
	);
	LUT2 #(
		.INIT('h4)
	) name18149 (
		_w28618_,
		_w28660_,
		_w28661_
	);
	LUT2 #(
		.INIT('h8)
	) name18150 (
		_w28658_,
		_w28659_,
		_w28662_
	);
	LUT2 #(
		.INIT('h8)
	) name18151 (
		_w28661_,
		_w28662_,
		_w28663_
	);
	LUT2 #(
		.INIT('h1)
	) name18152 (
		_w28613_,
		_w28663_,
		_w28664_
	);
	LUT2 #(
		.INIT('h2)
	) name18153 (
		\wishbone_TxLength_reg[7]/NET0131 ,
		_w17812_,
		_w28665_
	);
	LUT2 #(
		.INIT('h8)
	) name18154 (
		_w12657_,
		_w15113_,
		_w28666_
	);
	LUT2 #(
		.INIT('h1)
	) name18155 (
		_w28665_,
		_w28666_,
		_w28667_
	);
	LUT2 #(
		.INIT('h2)
	) name18156 (
		_w18569_,
		_w28667_,
		_w28668_
	);
	LUT2 #(
		.INIT('h1)
	) name18157 (
		_w22416_,
		_w28668_,
		_w28669_
	);
	LUT2 #(
		.INIT('h2)
	) name18158 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w12657_,
		_w28670_
	);
	LUT2 #(
		.INIT('h2)
	) name18159 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w16766_,
		_w28671_
	);
	LUT2 #(
		.INIT('h1)
	) name18160 (
		_w23564_,
		_w28671_,
		_w28672_
	);
	LUT2 #(
		.INIT('h2)
	) name18161 (
		_w16762_,
		_w28672_,
		_w28673_
	);
	LUT2 #(
		.INIT('h2)
	) name18162 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w13481_,
		_w28674_
	);
	LUT2 #(
		.INIT('h1)
	) name18163 (
		_w23553_,
		_w28674_,
		_w28675_
	);
	LUT2 #(
		.INIT('h4)
	) name18164 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w16757_,
		_w28676_
	);
	LUT2 #(
		.INIT('h2)
	) name18165 (
		_w16756_,
		_w28676_,
		_w28677_
	);
	LUT2 #(
		.INIT('h1)
	) name18166 (
		_w16748_,
		_w28677_,
		_w28678_
	);
	LUT2 #(
		.INIT('h1)
	) name18167 (
		_w28675_,
		_w28678_,
		_w28679_
	);
	LUT2 #(
		.INIT('h8)
	) name18168 (
		_w16757_,
		_w28677_,
		_w28680_
	);
	LUT2 #(
		.INIT('h2)
	) name18169 (
		\wishbone_TxLength_reg[5]/NET0131 ,
		_w16753_,
		_w28681_
	);
	LUT2 #(
		.INIT('h1)
	) name18170 (
		_w23561_,
		_w28681_,
		_w28682_
	);
	LUT2 #(
		.INIT('h2)
	) name18171 (
		_w16750_,
		_w28682_,
		_w28683_
	);
	LUT2 #(
		.INIT('h1)
	) name18172 (
		_w28679_,
		_w28680_,
		_w28684_
	);
	LUT2 #(
		.INIT('h4)
	) name18173 (
		_w28673_,
		_w28684_,
		_w28685_
	);
	LUT2 #(
		.INIT('h4)
	) name18174 (
		_w28683_,
		_w28685_,
		_w28686_
	);
	LUT2 #(
		.INIT('h2)
	) name18175 (
		_w13500_,
		_w28686_,
		_w28687_
	);
	LUT2 #(
		.INIT('h1)
	) name18176 (
		_w28670_,
		_w28687_,
		_w28688_
	);
	LUT2 #(
		.INIT('h1)
	) name18177 (
		_w12656_,
		_w28688_,
		_w28689_
	);
	LUT2 #(
		.INIT('h1)
	) name18178 (
		_w21901_,
		_w28689_,
		_w28690_
	);
	LUT2 #(
		.INIT('h8)
	) name18179 (
		\ethreg1_COLLCONF_2_DataOut_reg[0]/NET0131 ,
		_w24730_,
		_w28691_
	);
	LUT2 #(
		.INIT('h8)
	) name18180 (
		\ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 ,
		_w22956_,
		_w28692_
	);
	LUT2 #(
		.INIT('h8)
	) name18181 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		_w22959_,
		_w28693_
	);
	LUT2 #(
		.INIT('h8)
	) name18182 (
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		_w23519_,
		_w28694_
	);
	LUT2 #(
		.INIT('h8)
	) name18183 (
		\ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 ,
		_w22952_,
		_w28695_
	);
	LUT2 #(
		.INIT('h8)
	) name18184 (
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		_w23499_,
		_w28696_
	);
	LUT2 #(
		.INIT('h8)
	) name18185 (
		\ethreg1_PACKETLEN_2_DataOut_reg[0]/NET0131 ,
		_w22966_,
		_w28697_
	);
	LUT2 #(
		.INIT('h1)
	) name18186 (
		_w28692_,
		_w28693_,
		_w28698_
	);
	LUT2 #(
		.INIT('h1)
	) name18187 (
		_w28694_,
		_w28695_,
		_w28699_
	);
	LUT2 #(
		.INIT('h4)
	) name18188 (
		_w28696_,
		_w28699_,
		_w28700_
	);
	LUT2 #(
		.INIT('h8)
	) name18189 (
		_w28698_,
		_w28700_,
		_w28701_
	);
	LUT2 #(
		.INIT('h1)
	) name18190 (
		_w28691_,
		_w28697_,
		_w28702_
	);
	LUT2 #(
		.INIT('h8)
	) name18191 (
		_w28701_,
		_w28702_,
		_w28703_
	);
	LUT2 #(
		.INIT('h2)
	) name18192 (
		_w22944_,
		_w28703_,
		_w28704_
	);
	LUT2 #(
		.INIT('h2)
	) name18193 (
		_w19088_,
		_w22944_,
		_w28705_
	);
	LUT2 #(
		.INIT('h1)
	) name18194 (
		_w28704_,
		_w28705_,
		_w28706_
	);
	LUT2 #(
		.INIT('h8)
	) name18195 (
		\wishbone_bd_ram_mem0_reg[58][6]/P0001 ,
		_w13070_,
		_w28707_
	);
	LUT2 #(
		.INIT('h8)
	) name18196 (
		\wishbone_bd_ram_mem0_reg[56][6]/P0001 ,
		_w12778_,
		_w28708_
	);
	LUT2 #(
		.INIT('h8)
	) name18197 (
		\wishbone_bd_ram_mem0_reg[126][6]/P0001 ,
		_w13218_,
		_w28709_
	);
	LUT2 #(
		.INIT('h8)
	) name18198 (
		\wishbone_bd_ram_mem0_reg[125][6]/P0001 ,
		_w12956_,
		_w28710_
	);
	LUT2 #(
		.INIT('h8)
	) name18199 (
		\wishbone_bd_ram_mem0_reg[161][6]/P0001 ,
		_w12754_,
		_w28711_
	);
	LUT2 #(
		.INIT('h8)
	) name18200 (
		\wishbone_bd_ram_mem0_reg[243][6]/P0001 ,
		_w12804_,
		_w28712_
	);
	LUT2 #(
		.INIT('h8)
	) name18201 (
		\wishbone_bd_ram_mem0_reg[38][6]/P0001 ,
		_w13182_,
		_w28713_
	);
	LUT2 #(
		.INIT('h8)
	) name18202 (
		\wishbone_bd_ram_mem0_reg[22][6]/P0001 ,
		_w13110_,
		_w28714_
	);
	LUT2 #(
		.INIT('h8)
	) name18203 (
		\wishbone_bd_ram_mem0_reg[130][6]/P0001 ,
		_w12914_,
		_w28715_
	);
	LUT2 #(
		.INIT('h8)
	) name18204 (
		\wishbone_bd_ram_mem0_reg[18][6]/P0001 ,
		_w12679_,
		_w28716_
	);
	LUT2 #(
		.INIT('h8)
	) name18205 (
		\wishbone_bd_ram_mem0_reg[199][6]/P0001 ,
		_w12768_,
		_w28717_
	);
	LUT2 #(
		.INIT('h8)
	) name18206 (
		\wishbone_bd_ram_mem0_reg[45][6]/P0001 ,
		_w12908_,
		_w28718_
	);
	LUT2 #(
		.INIT('h8)
	) name18207 (
		\wishbone_bd_ram_mem0_reg[44][6]/P0001 ,
		_w12896_,
		_w28719_
	);
	LUT2 #(
		.INIT('h8)
	) name18208 (
		\wishbone_bd_ram_mem0_reg[94][6]/P0001 ,
		_w13186_,
		_w28720_
	);
	LUT2 #(
		.INIT('h8)
	) name18209 (
		\wishbone_bd_ram_mem0_reg[29][6]/P0001 ,
		_w12952_,
		_w28721_
	);
	LUT2 #(
		.INIT('h8)
	) name18210 (
		\wishbone_bd_ram_mem0_reg[66][6]/P0001 ,
		_w12824_,
		_w28722_
	);
	LUT2 #(
		.INIT('h8)
	) name18211 (
		\wishbone_bd_ram_mem0_reg[223][6]/P0001 ,
		_w12838_,
		_w28723_
	);
	LUT2 #(
		.INIT('h8)
	) name18212 (
		\wishbone_bd_ram_mem0_reg[196][6]/P0001 ,
		_w13090_,
		_w28724_
	);
	LUT2 #(
		.INIT('h8)
	) name18213 (
		\wishbone_bd_ram_mem0_reg[62][6]/P0001 ,
		_w12673_,
		_w28725_
	);
	LUT2 #(
		.INIT('h8)
	) name18214 (
		\wishbone_bd_ram_mem0_reg[52][6]/P0001 ,
		_w13082_,
		_w28726_
	);
	LUT2 #(
		.INIT('h8)
	) name18215 (
		\wishbone_bd_ram_mem0_reg[61][6]/P0001 ,
		_w12725_,
		_w28727_
	);
	LUT2 #(
		.INIT('h8)
	) name18216 (
		\wishbone_bd_ram_mem0_reg[162][6]/P0001 ,
		_w13098_,
		_w28728_
	);
	LUT2 #(
		.INIT('h8)
	) name18217 (
		\wishbone_bd_ram_mem0_reg[203][6]/P0001 ,
		_w13158_,
		_w28729_
	);
	LUT2 #(
		.INIT('h8)
	) name18218 (
		\wishbone_bd_ram_mem0_reg[231][6]/P0001 ,
		_w12856_,
		_w28730_
	);
	LUT2 #(
		.INIT('h8)
	) name18219 (
		\wishbone_bd_ram_mem0_reg[198][6]/P0001 ,
		_w12832_,
		_w28731_
	);
	LUT2 #(
		.INIT('h8)
	) name18220 (
		\wishbone_bd_ram_mem0_reg[98][6]/P0001 ,
		_w12816_,
		_w28732_
	);
	LUT2 #(
		.INIT('h8)
	) name18221 (
		\wishbone_bd_ram_mem0_reg[120][6]/P0001 ,
		_w12707_,
		_w28733_
	);
	LUT2 #(
		.INIT('h8)
	) name18222 (
		\wishbone_bd_ram_mem0_reg[63][6]/P0001 ,
		_w12850_,
		_w28734_
	);
	LUT2 #(
		.INIT('h8)
	) name18223 (
		\wishbone_bd_ram_mem0_reg[193][6]/P0001 ,
		_w13056_,
		_w28735_
	);
	LUT2 #(
		.INIT('h8)
	) name18224 (
		\wishbone_bd_ram_mem0_reg[59][6]/P0001 ,
		_w12780_,
		_w28736_
	);
	LUT2 #(
		.INIT('h8)
	) name18225 (
		\wishbone_bd_ram_mem0_reg[71][6]/P0001 ,
		_w12798_,
		_w28737_
	);
	LUT2 #(
		.INIT('h8)
	) name18226 (
		\wishbone_bd_ram_mem0_reg[191][6]/P0001 ,
		_w13034_,
		_w28738_
	);
	LUT2 #(
		.INIT('h8)
	) name18227 (
		\wishbone_bd_ram_mem0_reg[53][6]/P0001 ,
		_w13020_,
		_w28739_
	);
	LUT2 #(
		.INIT('h8)
	) name18228 (
		\wishbone_bd_ram_mem0_reg[187][6]/P0001 ,
		_w13196_,
		_w28740_
	);
	LUT2 #(
		.INIT('h8)
	) name18229 (
		\wishbone_bd_ram_mem0_reg[36][6]/P0001 ,
		_w12800_,
		_w28741_
	);
	LUT2 #(
		.INIT('h8)
	) name18230 (
		\wishbone_bd_ram_mem0_reg[155][6]/P0001 ,
		_w13122_,
		_w28742_
	);
	LUT2 #(
		.INIT('h8)
	) name18231 (
		\wishbone_bd_ram_mem0_reg[26][6]/P0001 ,
		_w12699_,
		_w28743_
	);
	LUT2 #(
		.INIT('h8)
	) name18232 (
		\wishbone_bd_ram_mem0_reg[117][6]/P0001 ,
		_w12715_,
		_w28744_
	);
	LUT2 #(
		.INIT('h8)
	) name18233 (
		\wishbone_bd_ram_mem0_reg[241][6]/P0001 ,
		_w13006_,
		_w28745_
	);
	LUT2 #(
		.INIT('h8)
	) name18234 (
		\wishbone_bd_ram_mem0_reg[248][6]/P0001 ,
		_w12789_,
		_w28746_
	);
	LUT2 #(
		.INIT('h8)
	) name18235 (
		\wishbone_bd_ram_mem0_reg[244][6]/P0001 ,
		_w12747_,
		_w28747_
	);
	LUT2 #(
		.INIT('h8)
	) name18236 (
		\wishbone_bd_ram_mem0_reg[215][6]/P0001 ,
		_w12974_,
		_w28748_
	);
	LUT2 #(
		.INIT('h8)
	) name18237 (
		\wishbone_bd_ram_mem0_reg[153][6]/P0001 ,
		_w12890_,
		_w28749_
	);
	LUT2 #(
		.INIT('h8)
	) name18238 (
		\wishbone_bd_ram_mem0_reg[131][6]/P0001 ,
		_w12852_,
		_w28750_
	);
	LUT2 #(
		.INIT('h8)
	) name18239 (
		\wishbone_bd_ram_mem0_reg[211][6]/P0001 ,
		_w13166_,
		_w28751_
	);
	LUT2 #(
		.INIT('h8)
	) name18240 (
		\wishbone_bd_ram_mem0_reg[81][6]/P0001 ,
		_w12950_,
		_w28752_
	);
	LUT2 #(
		.INIT('h8)
	) name18241 (
		\wishbone_bd_ram_mem0_reg[35][6]/P0001 ,
		_w12703_,
		_w28753_
	);
	LUT2 #(
		.INIT('h8)
	) name18242 (
		\wishbone_bd_ram_mem0_reg[238][6]/P0001 ,
		_w13160_,
		_w28754_
	);
	LUT2 #(
		.INIT('h8)
	) name18243 (
		\wishbone_bd_ram_mem0_reg[114][6]/P0001 ,
		_w13202_,
		_w28755_
	);
	LUT2 #(
		.INIT('h8)
	) name18244 (
		\wishbone_bd_ram_mem0_reg[227][6]/P0001 ,
		_w12936_,
		_w28756_
	);
	LUT2 #(
		.INIT('h8)
	) name18245 (
		\wishbone_bd_ram_mem0_reg[1][6]/P0001 ,
		_w13014_,
		_w28757_
	);
	LUT2 #(
		.INIT('h8)
	) name18246 (
		\wishbone_bd_ram_mem0_reg[60][6]/P0001 ,
		_w13204_,
		_w28758_
	);
	LUT2 #(
		.INIT('h8)
	) name18247 (
		\wishbone_bd_ram_mem0_reg[19][6]/P0001 ,
		_w13012_,
		_w28759_
	);
	LUT2 #(
		.INIT('h8)
	) name18248 (
		\wishbone_bd_ram_mem0_reg[133][6]/P0001 ,
		_w12761_,
		_w28760_
	);
	LUT2 #(
		.INIT('h8)
	) name18249 (
		\wishbone_bd_ram_mem0_reg[96][6]/P0001 ,
		_w12912_,
		_w28761_
	);
	LUT2 #(
		.INIT('h8)
	) name18250 (
		\wishbone_bd_ram_mem0_reg[224][6]/P0001 ,
		_w12902_,
		_w28762_
	);
	LUT2 #(
		.INIT('h8)
	) name18251 (
		\wishbone_bd_ram_mem0_reg[88][6]/P0001 ,
		_w12860_,
		_w28763_
	);
	LUT2 #(
		.INIT('h8)
	) name18252 (
		\wishbone_bd_ram_mem0_reg[254][6]/P0001 ,
		_w12892_,
		_w28764_
	);
	LUT2 #(
		.INIT('h8)
	) name18253 (
		\wishbone_bd_ram_mem0_reg[87][6]/P0001 ,
		_w13154_,
		_w28765_
	);
	LUT2 #(
		.INIT('h8)
	) name18254 (
		\wishbone_bd_ram_mem0_reg[100][6]/P0001 ,
		_w12960_,
		_w28766_
	);
	LUT2 #(
		.INIT('h8)
	) name18255 (
		\wishbone_bd_ram_mem0_reg[219][6]/P0001 ,
		_w12806_,
		_w28767_
	);
	LUT2 #(
		.INIT('h8)
	) name18256 (
		\wishbone_bd_ram_mem0_reg[179][6]/P0001 ,
		_w13050_,
		_w28768_
	);
	LUT2 #(
		.INIT('h8)
	) name18257 (
		\wishbone_bd_ram_mem0_reg[146][6]/P0001 ,
		_w13060_,
		_w28769_
	);
	LUT2 #(
		.INIT('h8)
	) name18258 (
		\wishbone_bd_ram_mem0_reg[204][6]/P0001 ,
		_w13162_,
		_w28770_
	);
	LUT2 #(
		.INIT('h8)
	) name18259 (
		\wishbone_bd_ram_mem0_reg[221][6]/P0001 ,
		_w12802_,
		_w28771_
	);
	LUT2 #(
		.INIT('h8)
	) name18260 (
		\wishbone_bd_ram_mem0_reg[127][6]/P0001 ,
		_w13164_,
		_w28772_
	);
	LUT2 #(
		.INIT('h8)
	) name18261 (
		\wishbone_bd_ram_mem0_reg[74][6]/P0001 ,
		_w12812_,
		_w28773_
	);
	LUT2 #(
		.INIT('h8)
	) name18262 (
		\wishbone_bd_ram_mem0_reg[4][6]/P0001 ,
		_w12666_,
		_w28774_
	);
	LUT2 #(
		.INIT('h8)
	) name18263 (
		\wishbone_bd_ram_mem0_reg[89][6]/P0001 ,
		_w12964_,
		_w28775_
	);
	LUT2 #(
		.INIT('h8)
	) name18264 (
		\wishbone_bd_ram_mem0_reg[104][6]/P0001 ,
		_w13148_,
		_w28776_
	);
	LUT2 #(
		.INIT('h8)
	) name18265 (
		\wishbone_bd_ram_mem0_reg[194][6]/P0001 ,
		_w12772_,
		_w28777_
	);
	LUT2 #(
		.INIT('h8)
	) name18266 (
		\wishbone_bd_ram_mem0_reg[92][6]/P0001 ,
		_w13010_,
		_w28778_
	);
	LUT2 #(
		.INIT('h8)
	) name18267 (
		\wishbone_bd_ram_mem0_reg[79][6]/P0001 ,
		_w13212_,
		_w28779_
	);
	LUT2 #(
		.INIT('h8)
	) name18268 (
		\wishbone_bd_ram_mem0_reg[212][6]/P0001 ,
		_w12796_,
		_w28780_
	);
	LUT2 #(
		.INIT('h8)
	) name18269 (
		\wishbone_bd_ram_mem0_reg[151][6]/P0001 ,
		_w13142_,
		_w28781_
	);
	LUT2 #(
		.INIT('h8)
	) name18270 (
		\wishbone_bd_ram_mem0_reg[225][6]/P0001 ,
		_w13092_,
		_w28782_
	);
	LUT2 #(
		.INIT('h8)
	) name18271 (
		\wishbone_bd_ram_mem0_reg[174][6]/P0001 ,
		_w12972_,
		_w28783_
	);
	LUT2 #(
		.INIT('h8)
	) name18272 (
		\wishbone_bd_ram_mem0_reg[178][6]/P0001 ,
		_w12886_,
		_w28784_
	);
	LUT2 #(
		.INIT('h8)
	) name18273 (
		\wishbone_bd_ram_mem0_reg[217][6]/P0001 ,
		_w13188_,
		_w28785_
	);
	LUT2 #(
		.INIT('h8)
	) name18274 (
		\wishbone_bd_ram_mem0_reg[72][6]/P0001 ,
		_w12810_,
		_w28786_
	);
	LUT2 #(
		.INIT('h8)
	) name18275 (
		\wishbone_bd_ram_mem0_reg[210][6]/P0001 ,
		_w12924_,
		_w28787_
	);
	LUT2 #(
		.INIT('h8)
	) name18276 (
		\wishbone_bd_ram_mem0_reg[121][6]/P0001 ,
		_w13078_,
		_w28788_
	);
	LUT2 #(
		.INIT('h8)
	) name18277 (
		\wishbone_bd_ram_mem0_reg[149][6]/P0001 ,
		_w12741_,
		_w28789_
	);
	LUT2 #(
		.INIT('h8)
	) name18278 (
		\wishbone_bd_ram_mem0_reg[183][6]/P0001 ,
		_w12787_,
		_w28790_
	);
	LUT2 #(
		.INIT('h8)
	) name18279 (
		\wishbone_bd_ram_mem0_reg[80][6]/P0001 ,
		_w12689_,
		_w28791_
	);
	LUT2 #(
		.INIT('h8)
	) name18280 (
		\wishbone_bd_ram_mem0_reg[33][6]/P0001 ,
		_w12980_,
		_w28792_
	);
	LUT2 #(
		.INIT('h8)
	) name18281 (
		\wishbone_bd_ram_mem0_reg[21][6]/P0001 ,
		_w12906_,
		_w28793_
	);
	LUT2 #(
		.INIT('h8)
	) name18282 (
		\wishbone_bd_ram_mem0_reg[73][6]/P0001 ,
		_w12918_,
		_w28794_
	);
	LUT2 #(
		.INIT('h8)
	) name18283 (
		\wishbone_bd_ram_mem0_reg[51][6]/P0001 ,
		_w13024_,
		_w28795_
	);
	LUT2 #(
		.INIT('h8)
	) name18284 (
		\wishbone_bd_ram_mem0_reg[252][6]/P0001 ,
		_w13080_,
		_w28796_
	);
	LUT2 #(
		.INIT('h8)
	) name18285 (
		\wishbone_bd_ram_mem0_reg[32][6]/P0001 ,
		_w13120_,
		_w28797_
	);
	LUT2 #(
		.INIT('h8)
	) name18286 (
		\wishbone_bd_ram_mem0_reg[144][6]/P0001 ,
		_w12756_,
		_w28798_
	);
	LUT2 #(
		.INIT('h8)
	) name18287 (
		\wishbone_bd_ram_mem0_reg[249][6]/P0001 ,
		_w12900_,
		_w28799_
	);
	LUT2 #(
		.INIT('h8)
	) name18288 (
		\wishbone_bd_ram_mem0_reg[255][6]/P0001 ,
		_w13072_,
		_w28800_
	);
	LUT2 #(
		.INIT('h8)
	) name18289 (
		\wishbone_bd_ram_mem0_reg[84][6]/P0001 ,
		_w12934_,
		_w28801_
	);
	LUT2 #(
		.INIT('h8)
	) name18290 (
		\wishbone_bd_ram_mem0_reg[237][6]/P0001 ,
		_w12990_,
		_w28802_
	);
	LUT2 #(
		.INIT('h8)
	) name18291 (
		\wishbone_bd_ram_mem0_reg[181][6]/P0001 ,
		_w12828_,
		_w28803_
	);
	LUT2 #(
		.INIT('h8)
	) name18292 (
		\wishbone_bd_ram_mem0_reg[113][6]/P0001 ,
		_w13026_,
		_w28804_
	);
	LUT2 #(
		.INIT('h8)
	) name18293 (
		\wishbone_bd_ram_mem0_reg[49][6]/P0001 ,
		_w12994_,
		_w28805_
	);
	LUT2 #(
		.INIT('h8)
	) name18294 (
		\wishbone_bd_ram_mem0_reg[13][6]/P0001 ,
		_w13178_,
		_w28806_
	);
	LUT2 #(
		.INIT('h8)
	) name18295 (
		\wishbone_bd_ram_mem0_reg[138][6]/P0001 ,
		_w12958_,
		_w28807_
	);
	LUT2 #(
		.INIT('h8)
	) name18296 (
		\wishbone_bd_ram_mem0_reg[177][6]/P0001 ,
		_w12996_,
		_w28808_
	);
	LUT2 #(
		.INIT('h8)
	) name18297 (
		\wishbone_bd_ram_mem0_reg[171][6]/P0001 ,
		_w12910_,
		_w28809_
	);
	LUT2 #(
		.INIT('h8)
	) name18298 (
		\wishbone_bd_ram_mem0_reg[182][6]/P0001 ,
		_w12820_,
		_w28810_
	);
	LUT2 #(
		.INIT('h8)
	) name18299 (
		\wishbone_bd_ram_mem0_reg[76][6]/P0001 ,
		_w13184_,
		_w28811_
	);
	LUT2 #(
		.INIT('h8)
	) name18300 (
		\wishbone_bd_ram_mem0_reg[109][6]/P0001 ,
		_w12888_,
		_w28812_
	);
	LUT2 #(
		.INIT('h8)
	) name18301 (
		\wishbone_bd_ram_mem0_reg[2][6]/P0001 ,
		_w13088_,
		_w28813_
	);
	LUT2 #(
		.INIT('h8)
	) name18302 (
		\wishbone_bd_ram_mem0_reg[186][6]/P0001 ,
		_w12783_,
		_w28814_
	);
	LUT2 #(
		.INIT('h8)
	) name18303 (
		\wishbone_bd_ram_mem0_reg[154][6]/P0001 ,
		_w12962_,
		_w28815_
	);
	LUT2 #(
		.INIT('h8)
	) name18304 (
		\wishbone_bd_ram_mem0_reg[118][6]/P0001 ,
		_w12830_,
		_w28816_
	);
	LUT2 #(
		.INIT('h8)
	) name18305 (
		\wishbone_bd_ram_mem0_reg[137][6]/P0001 ,
		_w13168_,
		_w28817_
	);
	LUT2 #(
		.INIT('h8)
	) name18306 (
		\wishbone_bd_ram_mem0_reg[20][6]/P0001 ,
		_w13174_,
		_w28818_
	);
	LUT2 #(
		.INIT('h8)
	) name18307 (
		\wishbone_bd_ram_mem0_reg[3][6]/P0001 ,
		_w12866_,
		_w28819_
	);
	LUT2 #(
		.INIT('h8)
	) name18308 (
		\wishbone_bd_ram_mem0_reg[85][6]/P0001 ,
		_w13216_,
		_w28820_
	);
	LUT2 #(
		.INIT('h8)
	) name18309 (
		\wishbone_bd_ram_mem0_reg[9][6]/P0001 ,
		_w12808_,
		_w28821_
	);
	LUT2 #(
		.INIT('h8)
	) name18310 (
		\wishbone_bd_ram_mem0_reg[145][6]/P0001 ,
		_w13106_,
		_w28822_
	);
	LUT2 #(
		.INIT('h8)
	) name18311 (
		\wishbone_bd_ram_mem0_reg[197][6]/P0001 ,
		_w12834_,
		_w28823_
	);
	LUT2 #(
		.INIT('h8)
	) name18312 (
		\wishbone_bd_ram_mem0_reg[208][6]/P0001 ,
		_w13032_,
		_w28824_
	);
	LUT2 #(
		.INIT('h8)
	) name18313 (
		\wishbone_bd_ram_mem0_reg[176][6]/P0001 ,
		_w12868_,
		_w28825_
	);
	LUT2 #(
		.INIT('h8)
	) name18314 (
		\wishbone_bd_ram_mem0_reg[65][6]/P0001 ,
		_w13176_,
		_w28826_
	);
	LUT2 #(
		.INIT('h8)
	) name18315 (
		\wishbone_bd_ram_mem0_reg[139][6]/P0001 ,
		_w12814_,
		_w28827_
	);
	LUT2 #(
		.INIT('h8)
	) name18316 (
		\wishbone_bd_ram_mem0_reg[207][6]/P0001 ,
		_w13180_,
		_w28828_
	);
	LUT2 #(
		.INIT('h8)
	) name18317 (
		\wishbone_bd_ram_mem0_reg[128][6]/P0001 ,
		_w12793_,
		_w28829_
	);
	LUT2 #(
		.INIT('h8)
	) name18318 (
		\wishbone_bd_ram_mem0_reg[216][6]/P0001 ,
		_w13028_,
		_w28830_
	);
	LUT2 #(
		.INIT('h8)
	) name18319 (
		\wishbone_bd_ram_mem0_reg[64][6]/P0001 ,
		_w12976_,
		_w28831_
	);
	LUT2 #(
		.INIT('h8)
	) name18320 (
		\wishbone_bd_ram_mem0_reg[147][6]/P0001 ,
		_w13146_,
		_w28832_
	);
	LUT2 #(
		.INIT('h8)
	) name18321 (
		\wishbone_bd_ram_mem0_reg[218][6]/P0001 ,
		_w13206_,
		_w28833_
	);
	LUT2 #(
		.INIT('h8)
	) name18322 (
		\wishbone_bd_ram_mem0_reg[188][6]/P0001 ,
		_w12948_,
		_w28834_
	);
	LUT2 #(
		.INIT('h8)
	) name18323 (
		\wishbone_bd_ram_mem0_reg[107][6]/P0001 ,
		_w12749_,
		_w28835_
	);
	LUT2 #(
		.INIT('h8)
	) name18324 (
		\wishbone_bd_ram_mem0_reg[165][6]/P0001 ,
		_w13044_,
		_w28836_
	);
	LUT2 #(
		.INIT('h8)
	) name18325 (
		\wishbone_bd_ram_mem0_reg[15][6]/P0001 ,
		_w13210_,
		_w28837_
	);
	LUT2 #(
		.INIT('h8)
	) name18326 (
		\wishbone_bd_ram_mem0_reg[115][6]/P0001 ,
		_w13112_,
		_w28838_
	);
	LUT2 #(
		.INIT('h8)
	) name18327 (
		\wishbone_bd_ram_mem0_reg[180][6]/P0001 ,
		_w12791_,
		_w28839_
	);
	LUT2 #(
		.INIT('h8)
	) name18328 (
		\wishbone_bd_ram_mem0_reg[46][6]/P0001 ,
		_w12884_,
		_w28840_
	);
	LUT2 #(
		.INIT('h8)
	) name18329 (
		\wishbone_bd_ram_mem0_reg[78][6]/P0001 ,
		_w12874_,
		_w28841_
	);
	LUT2 #(
		.INIT('h8)
	) name18330 (
		\wishbone_bd_ram_mem0_reg[230][6]/P0001 ,
		_w13036_,
		_w28842_
	);
	LUT2 #(
		.INIT('h8)
	) name18331 (
		\wishbone_bd_ram_mem0_reg[43][6]/P0001 ,
		_w13200_,
		_w28843_
	);
	LUT2 #(
		.INIT('h8)
	) name18332 (
		\wishbone_bd_ram_mem0_reg[86][6]/P0001 ,
		_w12735_,
		_w28844_
	);
	LUT2 #(
		.INIT('h8)
	) name18333 (
		\wishbone_bd_ram_mem0_reg[213][6]/P0001 ,
		_w13002_,
		_w28845_
	);
	LUT2 #(
		.INIT('h8)
	) name18334 (
		\wishbone_bd_ram_mem0_reg[150][6]/P0001 ,
		_w13136_,
		_w28846_
	);
	LUT2 #(
		.INIT('h8)
	) name18335 (
		\wishbone_bd_ram_mem0_reg[140][6]/P0001 ,
		_w12894_,
		_w28847_
	);
	LUT2 #(
		.INIT('h8)
	) name18336 (
		\wishbone_bd_ram_mem0_reg[202][6]/P0001 ,
		_w12870_,
		_w28848_
	);
	LUT2 #(
		.INIT('h8)
	) name18337 (
		\wishbone_bd_ram_mem0_reg[112][6]/P0001 ,
		_w12733_,
		_w28849_
	);
	LUT2 #(
		.INIT('h8)
	) name18338 (
		\wishbone_bd_ram_mem0_reg[135][6]/P0001 ,
		_w13124_,
		_w28850_
	);
	LUT2 #(
		.INIT('h8)
	) name18339 (
		\wishbone_bd_ram_mem0_reg[102][6]/P0001 ,
		_w12685_,
		_w28851_
	);
	LUT2 #(
		.INIT('h8)
	) name18340 (
		\wishbone_bd_ram_mem0_reg[129][6]/P0001 ,
		_w12776_,
		_w28852_
	);
	LUT2 #(
		.INIT('h8)
	) name18341 (
		\wishbone_bd_ram_mem0_reg[164][6]/P0001 ,
		_w12876_,
		_w28853_
	);
	LUT2 #(
		.INIT('h8)
	) name18342 (
		\wishbone_bd_ram_mem0_reg[233][6]/P0001 ,
		_w12836_,
		_w28854_
	);
	LUT2 #(
		.INIT('h8)
	) name18343 (
		\wishbone_bd_ram_mem0_reg[34][6]/P0001 ,
		_w12930_,
		_w28855_
	);
	LUT2 #(
		.INIT('h8)
	) name18344 (
		\wishbone_bd_ram_mem0_reg[222][6]/P0001 ,
		_w13094_,
		_w28856_
	);
	LUT2 #(
		.INIT('h8)
	) name18345 (
		\wishbone_bd_ram_mem0_reg[152][6]/P0001 ,
		_w12966_,
		_w28857_
	);
	LUT2 #(
		.INIT('h8)
	) name18346 (
		\wishbone_bd_ram_mem0_reg[93][6]/P0001 ,
		_w13016_,
		_w28858_
	);
	LUT2 #(
		.INIT('h8)
	) name18347 (
		\wishbone_bd_ram_mem0_reg[14][6]/P0001 ,
		_w13086_,
		_w28859_
	);
	LUT2 #(
		.INIT('h8)
	) name18348 (
		\wishbone_bd_ram_mem0_reg[5][6]/P0001 ,
		_w12878_,
		_w28860_
	);
	LUT2 #(
		.INIT('h8)
	) name18349 (
		\wishbone_bd_ram_mem0_reg[134][6]/P0001 ,
		_w12763_,
		_w28861_
	);
	LUT2 #(
		.INIT('h8)
	) name18350 (
		\wishbone_bd_ram_mem0_reg[77][6]/P0001 ,
		_w12982_,
		_w28862_
	);
	LUT2 #(
		.INIT('h8)
	) name18351 (
		\wishbone_bd_ram_mem0_reg[136][6]/P0001 ,
		_w13064_,
		_w28863_
	);
	LUT2 #(
		.INIT('h8)
	) name18352 (
		\wishbone_bd_ram_mem0_reg[239][6]/P0001 ,
		_w12862_,
		_w28864_
	);
	LUT2 #(
		.INIT('h8)
	) name18353 (
		\wishbone_bd_ram_mem0_reg[25][6]/P0001 ,
		_w13108_,
		_w28865_
	);
	LUT2 #(
		.INIT('h8)
	) name18354 (
		\wishbone_bd_ram_mem0_reg[106][6]/P0001 ,
		_w12713_,
		_w28866_
	);
	LUT2 #(
		.INIT('h8)
	) name18355 (
		\wishbone_bd_ram_mem0_reg[251][6]/P0001 ,
		_w13054_,
		_w28867_
	);
	LUT2 #(
		.INIT('h8)
	) name18356 (
		\wishbone_bd_ram_mem0_reg[235][6]/P0001 ,
		_w12696_,
		_w28868_
	);
	LUT2 #(
		.INIT('h8)
	) name18357 (
		\wishbone_bd_ram_mem0_reg[111][6]/P0001 ,
		_w12744_,
		_w28869_
	);
	LUT2 #(
		.INIT('h8)
	) name18358 (
		\wishbone_bd_ram_mem0_reg[247][6]/P0001 ,
		_w12818_,
		_w28870_
	);
	LUT2 #(
		.INIT('h8)
	) name18359 (
		\wishbone_bd_ram_mem0_reg[39][6]/P0001 ,
		_w13018_,
		_w28871_
	);
	LUT2 #(
		.INIT('h8)
	) name18360 (
		\wishbone_bd_ram_mem0_reg[116][6]/P0001 ,
		_w12998_,
		_w28872_
	);
	LUT2 #(
		.INIT('h8)
	) name18361 (
		\wishbone_bd_ram_mem0_reg[90][6]/P0001 ,
		_w12978_,
		_w28873_
	);
	LUT2 #(
		.INIT('h8)
	) name18362 (
		\wishbone_bd_ram_mem0_reg[156][6]/P0001 ,
		_w13190_,
		_w28874_
	);
	LUT2 #(
		.INIT('h8)
	) name18363 (
		\wishbone_bd_ram_mem0_reg[82][6]/P0001 ,
		_w12942_,
		_w28875_
	);
	LUT2 #(
		.INIT('h8)
	) name18364 (
		\wishbone_bd_ram_mem0_reg[105][6]/P0001 ,
		_w12751_,
		_w28876_
	);
	LUT2 #(
		.INIT('h8)
	) name18365 (
		\wishbone_bd_ram_mem0_reg[37][6]/P0001 ,
		_w13102_,
		_w28877_
	);
	LUT2 #(
		.INIT('h8)
	) name18366 (
		\wishbone_bd_ram_mem0_reg[185][6]/P0001 ,
		_w12940_,
		_w28878_
	);
	LUT2 #(
		.INIT('h8)
	) name18367 (
		\wishbone_bd_ram_mem0_reg[48][6]/P0001 ,
		_w12970_,
		_w28879_
	);
	LUT2 #(
		.INIT('h8)
	) name18368 (
		\wishbone_bd_ram_mem0_reg[253][6]/P0001 ,
		_w13100_,
		_w28880_
	);
	LUT2 #(
		.INIT('h8)
	) name18369 (
		\wishbone_bd_ram_mem0_reg[172][6]/P0001 ,
		_w12944_,
		_w28881_
	);
	LUT2 #(
		.INIT('h8)
	) name18370 (
		\wishbone_bd_ram_mem0_reg[228][6]/P0001 ,
		_w12765_,
		_w28882_
	);
	LUT2 #(
		.INIT('h8)
	) name18371 (
		\wishbone_bd_ram_mem0_reg[192][6]/P0001 ,
		_w12938_,
		_w28883_
	);
	LUT2 #(
		.INIT('h8)
	) name18372 (
		\wishbone_bd_ram_mem0_reg[169][6]/P0001 ,
		_w12722_,
		_w28884_
	);
	LUT2 #(
		.INIT('h8)
	) name18373 (
		\wishbone_bd_ram_mem0_reg[201][6]/P0001 ,
		_w12822_,
		_w28885_
	);
	LUT2 #(
		.INIT('h8)
	) name18374 (
		\wishbone_bd_ram_mem0_reg[200][6]/P0001 ,
		_w12988_,
		_w28886_
	);
	LUT2 #(
		.INIT('h8)
	) name18375 (
		\wishbone_bd_ram_mem0_reg[173][6]/P0001 ,
		_w12854_,
		_w28887_
	);
	LUT2 #(
		.INIT('h8)
	) name18376 (
		\wishbone_bd_ram_mem0_reg[67][6]/P0001 ,
		_w13134_,
		_w28888_
	);
	LUT2 #(
		.INIT('h8)
	) name18377 (
		\wishbone_bd_ram_mem0_reg[205][6]/P0001 ,
		_w13068_,
		_w28889_
	);
	LUT2 #(
		.INIT('h8)
	) name18378 (
		\wishbone_bd_ram_mem0_reg[158][6]/P0001 ,
		_w12898_,
		_w28890_
	);
	LUT2 #(
		.INIT('h8)
	) name18379 (
		\wishbone_bd_ram_mem0_reg[214][6]/P0001 ,
		_w12984_,
		_w28891_
	);
	LUT2 #(
		.INIT('h8)
	) name18380 (
		\wishbone_bd_ram_mem0_reg[108][6]/P0001 ,
		_w13156_,
		_w28892_
	);
	LUT2 #(
		.INIT('h8)
	) name18381 (
		\wishbone_bd_ram_mem0_reg[10][6]/P0001 ,
		_w13172_,
		_w28893_
	);
	LUT2 #(
		.INIT('h8)
	) name18382 (
		\wishbone_bd_ram_mem0_reg[27][6]/P0001 ,
		_w12880_,
		_w28894_
	);
	LUT2 #(
		.INIT('h8)
	) name18383 (
		\wishbone_bd_ram_mem0_reg[16][6]/P0001 ,
		_w13140_,
		_w28895_
	);
	LUT2 #(
		.INIT('h8)
	) name18384 (
		\wishbone_bd_ram_mem0_reg[11][6]/P0001 ,
		_w13194_,
		_w28896_
	);
	LUT2 #(
		.INIT('h8)
	) name18385 (
		\wishbone_bd_ram_mem0_reg[24][6]/P0001 ,
		_w13084_,
		_w28897_
	);
	LUT2 #(
		.INIT('h8)
	) name18386 (
		\wishbone_bd_ram_mem0_reg[184][6]/P0001 ,
		_w13062_,
		_w28898_
	);
	LUT2 #(
		.INIT('h8)
	) name18387 (
		\wishbone_bd_ram_mem0_reg[246][6]/P0001 ,
		_w13076_,
		_w28899_
	);
	LUT2 #(
		.INIT('h8)
	) name18388 (
		\wishbone_bd_ram_mem0_reg[110][6]/P0001 ,
		_w13046_,
		_w28900_
	);
	LUT2 #(
		.INIT('h8)
	) name18389 (
		\wishbone_bd_ram_mem0_reg[91][6]/P0001 ,
		_w13074_,
		_w28901_
	);
	LUT2 #(
		.INIT('h8)
	) name18390 (
		\wishbone_bd_ram_mem0_reg[234][6]/P0001 ,
		_w13214_,
		_w28902_
	);
	LUT2 #(
		.INIT('h8)
	) name18391 (
		\wishbone_bd_ram_mem0_reg[240][6]/P0001 ,
		_w12864_,
		_w28903_
	);
	LUT2 #(
		.INIT('h8)
	) name18392 (
		\wishbone_bd_ram_mem0_reg[68][6]/P0001 ,
		_w12946_,
		_w28904_
	);
	LUT2 #(
		.INIT('h8)
	) name18393 (
		\wishbone_bd_ram_mem0_reg[28][6]/P0001 ,
		_w13170_,
		_w28905_
	);
	LUT2 #(
		.INIT('h8)
	) name18394 (
		\wishbone_bd_ram_mem0_reg[103][6]/P0001 ,
		_w12846_,
		_w28906_
	);
	LUT2 #(
		.INIT('h8)
	) name18395 (
		\wishbone_bd_ram_mem0_reg[101][6]/P0001 ,
		_w13192_,
		_w28907_
	);
	LUT2 #(
		.INIT('h8)
	) name18396 (
		\wishbone_bd_ram_mem0_reg[7][6]/P0001 ,
		_w12728_,
		_w28908_
	);
	LUT2 #(
		.INIT('h8)
	) name18397 (
		\wishbone_bd_ram_mem0_reg[142][6]/P0001 ,
		_w12928_,
		_w28909_
	);
	LUT2 #(
		.INIT('h8)
	) name18398 (
		\wishbone_bd_ram_mem0_reg[54][6]/P0001 ,
		_w12770_,
		_w28910_
	);
	LUT2 #(
		.INIT('h8)
	) name18399 (
		\wishbone_bd_ram_mem0_reg[95][6]/P0001 ,
		_w12844_,
		_w28911_
	);
	LUT2 #(
		.INIT('h8)
	) name18400 (
		\wishbone_bd_ram_mem0_reg[8][6]/P0001 ,
		_w12920_,
		_w28912_
	);
	LUT2 #(
		.INIT('h8)
	) name18401 (
		\wishbone_bd_ram_mem0_reg[70][6]/P0001 ,
		_w12840_,
		_w28913_
	);
	LUT2 #(
		.INIT('h8)
	) name18402 (
		\wishbone_bd_ram_mem0_reg[83][6]/P0001 ,
		_w12916_,
		_w28914_
	);
	LUT2 #(
		.INIT('h8)
	) name18403 (
		\wishbone_bd_ram_mem0_reg[141][6]/P0001 ,
		_w13004_,
		_w28915_
	);
	LUT2 #(
		.INIT('h8)
	) name18404 (
		\wishbone_bd_ram_mem0_reg[40][6]/P0001 ,
		_w13132_,
		_w28916_
	);
	LUT2 #(
		.INIT('h8)
	) name18405 (
		\wishbone_bd_ram_mem0_reg[229][6]/P0001 ,
		_w12711_,
		_w28917_
	);
	LUT2 #(
		.INIT('h8)
	) name18406 (
		\wishbone_bd_ram_mem0_reg[57][6]/P0001 ,
		_w13116_,
		_w28918_
	);
	LUT2 #(
		.INIT('h8)
	) name18407 (
		\wishbone_bd_ram_mem0_reg[50][6]/P0001 ,
		_w13150_,
		_w28919_
	);
	LUT2 #(
		.INIT('h8)
	) name18408 (
		\wishbone_bd_ram_mem0_reg[12][6]/P0001 ,
		_w13118_,
		_w28920_
	);
	LUT2 #(
		.INIT('h8)
	) name18409 (
		\wishbone_bd_ram_mem0_reg[99][6]/P0001 ,
		_w13038_,
		_w28921_
	);
	LUT2 #(
		.INIT('h8)
	) name18410 (
		\wishbone_bd_ram_mem0_reg[206][6]/P0001 ,
		_w12954_,
		_w28922_
	);
	LUT2 #(
		.INIT('h8)
	) name18411 (
		\wishbone_bd_ram_mem0_reg[148][6]/P0001 ,
		_w13000_,
		_w28923_
	);
	LUT2 #(
		.INIT('h8)
	) name18412 (
		\wishbone_bd_ram_mem0_reg[132][6]/P0001 ,
		_w12992_,
		_w28924_
	);
	LUT2 #(
		.INIT('h8)
	) name18413 (
		\wishbone_bd_ram_mem0_reg[124][6]/P0001 ,
		_w13058_,
		_w28925_
	);
	LUT2 #(
		.INIT('h8)
	) name18414 (
		\wishbone_bd_ram_mem0_reg[163][6]/P0001 ,
		_w12882_,
		_w28926_
	);
	LUT2 #(
		.INIT('h8)
	) name18415 (
		\wishbone_bd_ram_mem0_reg[143][6]/P0001 ,
		_w12922_,
		_w28927_
	);
	LUT2 #(
		.INIT('h8)
	) name18416 (
		\wishbone_bd_ram_mem0_reg[17][6]/P0001 ,
		_w12848_,
		_w28928_
	);
	LUT2 #(
		.INIT('h8)
	) name18417 (
		\wishbone_bd_ram_mem0_reg[236][6]/P0001 ,
		_w12731_,
		_w28929_
	);
	LUT2 #(
		.INIT('h8)
	) name18418 (
		\wishbone_bd_ram_mem0_reg[168][6]/P0001 ,
		_w13208_,
		_w28930_
	);
	LUT2 #(
		.INIT('h8)
	) name18419 (
		\wishbone_bd_ram_mem0_reg[189][6]/P0001 ,
		_w13042_,
		_w28931_
	);
	LUT2 #(
		.INIT('h8)
	) name18420 (
		\wishbone_bd_ram_mem0_reg[55][6]/P0001 ,
		_w12785_,
		_w28932_
	);
	LUT2 #(
		.INIT('h8)
	) name18421 (
		\wishbone_bd_ram_mem0_reg[190][6]/P0001 ,
		_w12858_,
		_w28933_
	);
	LUT2 #(
		.INIT('h8)
	) name18422 (
		\wishbone_bd_ram_mem0_reg[170][6]/P0001 ,
		_w13030_,
		_w28934_
	);
	LUT2 #(
		.INIT('h8)
	) name18423 (
		\wishbone_bd_ram_mem0_reg[242][6]/P0001 ,
		_w12932_,
		_w28935_
	);
	LUT2 #(
		.INIT('h8)
	) name18424 (
		\wishbone_bd_ram_mem0_reg[220][6]/P0001 ,
		_w13066_,
		_w28936_
	);
	LUT2 #(
		.INIT('h8)
	) name18425 (
		\wishbone_bd_ram_mem0_reg[123][6]/P0001 ,
		_w13114_,
		_w28937_
	);
	LUT2 #(
		.INIT('h8)
	) name18426 (
		\wishbone_bd_ram_mem0_reg[6][6]/P0001 ,
		_w12968_,
		_w28938_
	);
	LUT2 #(
		.INIT('h8)
	) name18427 (
		\wishbone_bd_ram_mem0_reg[75][6]/P0001 ,
		_w12826_,
		_w28939_
	);
	LUT2 #(
		.INIT('h8)
	) name18428 (
		\wishbone_bd_ram_mem0_reg[47][6]/P0001 ,
		_w12904_,
		_w28940_
	);
	LUT2 #(
		.INIT('h8)
	) name18429 (
		\wishbone_bd_ram_mem0_reg[42][6]/P0001 ,
		_w12842_,
		_w28941_
	);
	LUT2 #(
		.INIT('h8)
	) name18430 (
		\wishbone_bd_ram_mem0_reg[0][6]/P0001 ,
		_w12717_,
		_w28942_
	);
	LUT2 #(
		.INIT('h8)
	) name18431 (
		\wishbone_bd_ram_mem0_reg[250][6]/P0001 ,
		_w13128_,
		_w28943_
	);
	LUT2 #(
		.INIT('h8)
	) name18432 (
		\wishbone_bd_ram_mem0_reg[119][6]/P0001 ,
		_w13048_,
		_w28944_
	);
	LUT2 #(
		.INIT('h8)
	) name18433 (
		\wishbone_bd_ram_mem0_reg[159][6]/P0001 ,
		_w12774_,
		_w28945_
	);
	LUT2 #(
		.INIT('h8)
	) name18434 (
		\wishbone_bd_ram_mem0_reg[232][6]/P0001 ,
		_w12758_,
		_w28946_
	);
	LUT2 #(
		.INIT('h8)
	) name18435 (
		\wishbone_bd_ram_mem0_reg[245][6]/P0001 ,
		_w13022_,
		_w28947_
	);
	LUT2 #(
		.INIT('h8)
	) name18436 (
		\wishbone_bd_ram_mem0_reg[166][6]/P0001 ,
		_w13040_,
		_w28948_
	);
	LUT2 #(
		.INIT('h8)
	) name18437 (
		\wishbone_bd_ram_mem0_reg[97][6]/P0001 ,
		_w13096_,
		_w28949_
	);
	LUT2 #(
		.INIT('h8)
	) name18438 (
		\wishbone_bd_ram_mem0_reg[31][6]/P0001 ,
		_w13198_,
		_w28950_
	);
	LUT2 #(
		.INIT('h8)
	) name18439 (
		\wishbone_bd_ram_mem0_reg[226][6]/P0001 ,
		_w13138_,
		_w28951_
	);
	LUT2 #(
		.INIT('h8)
	) name18440 (
		\wishbone_bd_ram_mem0_reg[23][6]/P0001 ,
		_w13008_,
		_w28952_
	);
	LUT2 #(
		.INIT('h8)
	) name18441 (
		\wishbone_bd_ram_mem0_reg[30][6]/P0001 ,
		_w13104_,
		_w28953_
	);
	LUT2 #(
		.INIT('h8)
	) name18442 (
		\wishbone_bd_ram_mem0_reg[209][6]/P0001 ,
		_w13152_,
		_w28954_
	);
	LUT2 #(
		.INIT('h8)
	) name18443 (
		\wishbone_bd_ram_mem0_reg[157][6]/P0001 ,
		_w12926_,
		_w28955_
	);
	LUT2 #(
		.INIT('h8)
	) name18444 (
		\wishbone_bd_ram_mem0_reg[122][6]/P0001 ,
		_w13130_,
		_w28956_
	);
	LUT2 #(
		.INIT('h8)
	) name18445 (
		\wishbone_bd_ram_mem0_reg[167][6]/P0001 ,
		_w12986_,
		_w28957_
	);
	LUT2 #(
		.INIT('h8)
	) name18446 (
		\wishbone_bd_ram_mem0_reg[41][6]/P0001 ,
		_w13052_,
		_w28958_
	);
	LUT2 #(
		.INIT('h8)
	) name18447 (
		\wishbone_bd_ram_mem0_reg[69][6]/P0001 ,
		_w12738_,
		_w28959_
	);
	LUT2 #(
		.INIT('h8)
	) name18448 (
		\wishbone_bd_ram_mem0_reg[195][6]/P0001 ,
		_w13144_,
		_w28960_
	);
	LUT2 #(
		.INIT('h8)
	) name18449 (
		\wishbone_bd_ram_mem0_reg[160][6]/P0001 ,
		_w12872_,
		_w28961_
	);
	LUT2 #(
		.INIT('h8)
	) name18450 (
		\wishbone_bd_ram_mem0_reg[175][6]/P0001 ,
		_w13126_,
		_w28962_
	);
	LUT2 #(
		.INIT('h1)
	) name18451 (
		_w28707_,
		_w28708_,
		_w28963_
	);
	LUT2 #(
		.INIT('h1)
	) name18452 (
		_w28709_,
		_w28710_,
		_w28964_
	);
	LUT2 #(
		.INIT('h1)
	) name18453 (
		_w28711_,
		_w28712_,
		_w28965_
	);
	LUT2 #(
		.INIT('h1)
	) name18454 (
		_w28713_,
		_w28714_,
		_w28966_
	);
	LUT2 #(
		.INIT('h1)
	) name18455 (
		_w28715_,
		_w28716_,
		_w28967_
	);
	LUT2 #(
		.INIT('h1)
	) name18456 (
		_w28717_,
		_w28718_,
		_w28968_
	);
	LUT2 #(
		.INIT('h1)
	) name18457 (
		_w28719_,
		_w28720_,
		_w28969_
	);
	LUT2 #(
		.INIT('h1)
	) name18458 (
		_w28721_,
		_w28722_,
		_w28970_
	);
	LUT2 #(
		.INIT('h1)
	) name18459 (
		_w28723_,
		_w28724_,
		_w28971_
	);
	LUT2 #(
		.INIT('h1)
	) name18460 (
		_w28725_,
		_w28726_,
		_w28972_
	);
	LUT2 #(
		.INIT('h1)
	) name18461 (
		_w28727_,
		_w28728_,
		_w28973_
	);
	LUT2 #(
		.INIT('h1)
	) name18462 (
		_w28729_,
		_w28730_,
		_w28974_
	);
	LUT2 #(
		.INIT('h1)
	) name18463 (
		_w28731_,
		_w28732_,
		_w28975_
	);
	LUT2 #(
		.INIT('h1)
	) name18464 (
		_w28733_,
		_w28734_,
		_w28976_
	);
	LUT2 #(
		.INIT('h1)
	) name18465 (
		_w28735_,
		_w28736_,
		_w28977_
	);
	LUT2 #(
		.INIT('h1)
	) name18466 (
		_w28737_,
		_w28738_,
		_w28978_
	);
	LUT2 #(
		.INIT('h1)
	) name18467 (
		_w28739_,
		_w28740_,
		_w28979_
	);
	LUT2 #(
		.INIT('h1)
	) name18468 (
		_w28741_,
		_w28742_,
		_w28980_
	);
	LUT2 #(
		.INIT('h1)
	) name18469 (
		_w28743_,
		_w28744_,
		_w28981_
	);
	LUT2 #(
		.INIT('h1)
	) name18470 (
		_w28745_,
		_w28746_,
		_w28982_
	);
	LUT2 #(
		.INIT('h1)
	) name18471 (
		_w28747_,
		_w28748_,
		_w28983_
	);
	LUT2 #(
		.INIT('h1)
	) name18472 (
		_w28749_,
		_w28750_,
		_w28984_
	);
	LUT2 #(
		.INIT('h1)
	) name18473 (
		_w28751_,
		_w28752_,
		_w28985_
	);
	LUT2 #(
		.INIT('h1)
	) name18474 (
		_w28753_,
		_w28754_,
		_w28986_
	);
	LUT2 #(
		.INIT('h1)
	) name18475 (
		_w28755_,
		_w28756_,
		_w28987_
	);
	LUT2 #(
		.INIT('h1)
	) name18476 (
		_w28757_,
		_w28758_,
		_w28988_
	);
	LUT2 #(
		.INIT('h1)
	) name18477 (
		_w28759_,
		_w28760_,
		_w28989_
	);
	LUT2 #(
		.INIT('h1)
	) name18478 (
		_w28761_,
		_w28762_,
		_w28990_
	);
	LUT2 #(
		.INIT('h1)
	) name18479 (
		_w28763_,
		_w28764_,
		_w28991_
	);
	LUT2 #(
		.INIT('h1)
	) name18480 (
		_w28765_,
		_w28766_,
		_w28992_
	);
	LUT2 #(
		.INIT('h1)
	) name18481 (
		_w28767_,
		_w28768_,
		_w28993_
	);
	LUT2 #(
		.INIT('h1)
	) name18482 (
		_w28769_,
		_w28770_,
		_w28994_
	);
	LUT2 #(
		.INIT('h1)
	) name18483 (
		_w28771_,
		_w28772_,
		_w28995_
	);
	LUT2 #(
		.INIT('h1)
	) name18484 (
		_w28773_,
		_w28774_,
		_w28996_
	);
	LUT2 #(
		.INIT('h1)
	) name18485 (
		_w28775_,
		_w28776_,
		_w28997_
	);
	LUT2 #(
		.INIT('h1)
	) name18486 (
		_w28777_,
		_w28778_,
		_w28998_
	);
	LUT2 #(
		.INIT('h1)
	) name18487 (
		_w28779_,
		_w28780_,
		_w28999_
	);
	LUT2 #(
		.INIT('h1)
	) name18488 (
		_w28781_,
		_w28782_,
		_w29000_
	);
	LUT2 #(
		.INIT('h1)
	) name18489 (
		_w28783_,
		_w28784_,
		_w29001_
	);
	LUT2 #(
		.INIT('h1)
	) name18490 (
		_w28785_,
		_w28786_,
		_w29002_
	);
	LUT2 #(
		.INIT('h1)
	) name18491 (
		_w28787_,
		_w28788_,
		_w29003_
	);
	LUT2 #(
		.INIT('h1)
	) name18492 (
		_w28789_,
		_w28790_,
		_w29004_
	);
	LUT2 #(
		.INIT('h1)
	) name18493 (
		_w28791_,
		_w28792_,
		_w29005_
	);
	LUT2 #(
		.INIT('h1)
	) name18494 (
		_w28793_,
		_w28794_,
		_w29006_
	);
	LUT2 #(
		.INIT('h1)
	) name18495 (
		_w28795_,
		_w28796_,
		_w29007_
	);
	LUT2 #(
		.INIT('h1)
	) name18496 (
		_w28797_,
		_w28798_,
		_w29008_
	);
	LUT2 #(
		.INIT('h1)
	) name18497 (
		_w28799_,
		_w28800_,
		_w29009_
	);
	LUT2 #(
		.INIT('h1)
	) name18498 (
		_w28801_,
		_w28802_,
		_w29010_
	);
	LUT2 #(
		.INIT('h1)
	) name18499 (
		_w28803_,
		_w28804_,
		_w29011_
	);
	LUT2 #(
		.INIT('h1)
	) name18500 (
		_w28805_,
		_w28806_,
		_w29012_
	);
	LUT2 #(
		.INIT('h1)
	) name18501 (
		_w28807_,
		_w28808_,
		_w29013_
	);
	LUT2 #(
		.INIT('h1)
	) name18502 (
		_w28809_,
		_w28810_,
		_w29014_
	);
	LUT2 #(
		.INIT('h1)
	) name18503 (
		_w28811_,
		_w28812_,
		_w29015_
	);
	LUT2 #(
		.INIT('h1)
	) name18504 (
		_w28813_,
		_w28814_,
		_w29016_
	);
	LUT2 #(
		.INIT('h1)
	) name18505 (
		_w28815_,
		_w28816_,
		_w29017_
	);
	LUT2 #(
		.INIT('h1)
	) name18506 (
		_w28817_,
		_w28818_,
		_w29018_
	);
	LUT2 #(
		.INIT('h1)
	) name18507 (
		_w28819_,
		_w28820_,
		_w29019_
	);
	LUT2 #(
		.INIT('h1)
	) name18508 (
		_w28821_,
		_w28822_,
		_w29020_
	);
	LUT2 #(
		.INIT('h1)
	) name18509 (
		_w28823_,
		_w28824_,
		_w29021_
	);
	LUT2 #(
		.INIT('h1)
	) name18510 (
		_w28825_,
		_w28826_,
		_w29022_
	);
	LUT2 #(
		.INIT('h1)
	) name18511 (
		_w28827_,
		_w28828_,
		_w29023_
	);
	LUT2 #(
		.INIT('h1)
	) name18512 (
		_w28829_,
		_w28830_,
		_w29024_
	);
	LUT2 #(
		.INIT('h1)
	) name18513 (
		_w28831_,
		_w28832_,
		_w29025_
	);
	LUT2 #(
		.INIT('h1)
	) name18514 (
		_w28833_,
		_w28834_,
		_w29026_
	);
	LUT2 #(
		.INIT('h1)
	) name18515 (
		_w28835_,
		_w28836_,
		_w29027_
	);
	LUT2 #(
		.INIT('h1)
	) name18516 (
		_w28837_,
		_w28838_,
		_w29028_
	);
	LUT2 #(
		.INIT('h1)
	) name18517 (
		_w28839_,
		_w28840_,
		_w29029_
	);
	LUT2 #(
		.INIT('h1)
	) name18518 (
		_w28841_,
		_w28842_,
		_w29030_
	);
	LUT2 #(
		.INIT('h1)
	) name18519 (
		_w28843_,
		_w28844_,
		_w29031_
	);
	LUT2 #(
		.INIT('h1)
	) name18520 (
		_w28845_,
		_w28846_,
		_w29032_
	);
	LUT2 #(
		.INIT('h1)
	) name18521 (
		_w28847_,
		_w28848_,
		_w29033_
	);
	LUT2 #(
		.INIT('h1)
	) name18522 (
		_w28849_,
		_w28850_,
		_w29034_
	);
	LUT2 #(
		.INIT('h1)
	) name18523 (
		_w28851_,
		_w28852_,
		_w29035_
	);
	LUT2 #(
		.INIT('h1)
	) name18524 (
		_w28853_,
		_w28854_,
		_w29036_
	);
	LUT2 #(
		.INIT('h1)
	) name18525 (
		_w28855_,
		_w28856_,
		_w29037_
	);
	LUT2 #(
		.INIT('h1)
	) name18526 (
		_w28857_,
		_w28858_,
		_w29038_
	);
	LUT2 #(
		.INIT('h1)
	) name18527 (
		_w28859_,
		_w28860_,
		_w29039_
	);
	LUT2 #(
		.INIT('h1)
	) name18528 (
		_w28861_,
		_w28862_,
		_w29040_
	);
	LUT2 #(
		.INIT('h1)
	) name18529 (
		_w28863_,
		_w28864_,
		_w29041_
	);
	LUT2 #(
		.INIT('h1)
	) name18530 (
		_w28865_,
		_w28866_,
		_w29042_
	);
	LUT2 #(
		.INIT('h1)
	) name18531 (
		_w28867_,
		_w28868_,
		_w29043_
	);
	LUT2 #(
		.INIT('h1)
	) name18532 (
		_w28869_,
		_w28870_,
		_w29044_
	);
	LUT2 #(
		.INIT('h1)
	) name18533 (
		_w28871_,
		_w28872_,
		_w29045_
	);
	LUT2 #(
		.INIT('h1)
	) name18534 (
		_w28873_,
		_w28874_,
		_w29046_
	);
	LUT2 #(
		.INIT('h1)
	) name18535 (
		_w28875_,
		_w28876_,
		_w29047_
	);
	LUT2 #(
		.INIT('h1)
	) name18536 (
		_w28877_,
		_w28878_,
		_w29048_
	);
	LUT2 #(
		.INIT('h1)
	) name18537 (
		_w28879_,
		_w28880_,
		_w29049_
	);
	LUT2 #(
		.INIT('h1)
	) name18538 (
		_w28881_,
		_w28882_,
		_w29050_
	);
	LUT2 #(
		.INIT('h1)
	) name18539 (
		_w28883_,
		_w28884_,
		_w29051_
	);
	LUT2 #(
		.INIT('h1)
	) name18540 (
		_w28885_,
		_w28886_,
		_w29052_
	);
	LUT2 #(
		.INIT('h1)
	) name18541 (
		_w28887_,
		_w28888_,
		_w29053_
	);
	LUT2 #(
		.INIT('h1)
	) name18542 (
		_w28889_,
		_w28890_,
		_w29054_
	);
	LUT2 #(
		.INIT('h1)
	) name18543 (
		_w28891_,
		_w28892_,
		_w29055_
	);
	LUT2 #(
		.INIT('h1)
	) name18544 (
		_w28893_,
		_w28894_,
		_w29056_
	);
	LUT2 #(
		.INIT('h1)
	) name18545 (
		_w28895_,
		_w28896_,
		_w29057_
	);
	LUT2 #(
		.INIT('h1)
	) name18546 (
		_w28897_,
		_w28898_,
		_w29058_
	);
	LUT2 #(
		.INIT('h1)
	) name18547 (
		_w28899_,
		_w28900_,
		_w29059_
	);
	LUT2 #(
		.INIT('h1)
	) name18548 (
		_w28901_,
		_w28902_,
		_w29060_
	);
	LUT2 #(
		.INIT('h1)
	) name18549 (
		_w28903_,
		_w28904_,
		_w29061_
	);
	LUT2 #(
		.INIT('h1)
	) name18550 (
		_w28905_,
		_w28906_,
		_w29062_
	);
	LUT2 #(
		.INIT('h1)
	) name18551 (
		_w28907_,
		_w28908_,
		_w29063_
	);
	LUT2 #(
		.INIT('h1)
	) name18552 (
		_w28909_,
		_w28910_,
		_w29064_
	);
	LUT2 #(
		.INIT('h1)
	) name18553 (
		_w28911_,
		_w28912_,
		_w29065_
	);
	LUT2 #(
		.INIT('h1)
	) name18554 (
		_w28913_,
		_w28914_,
		_w29066_
	);
	LUT2 #(
		.INIT('h1)
	) name18555 (
		_w28915_,
		_w28916_,
		_w29067_
	);
	LUT2 #(
		.INIT('h1)
	) name18556 (
		_w28917_,
		_w28918_,
		_w29068_
	);
	LUT2 #(
		.INIT('h1)
	) name18557 (
		_w28919_,
		_w28920_,
		_w29069_
	);
	LUT2 #(
		.INIT('h1)
	) name18558 (
		_w28921_,
		_w28922_,
		_w29070_
	);
	LUT2 #(
		.INIT('h1)
	) name18559 (
		_w28923_,
		_w28924_,
		_w29071_
	);
	LUT2 #(
		.INIT('h1)
	) name18560 (
		_w28925_,
		_w28926_,
		_w29072_
	);
	LUT2 #(
		.INIT('h1)
	) name18561 (
		_w28927_,
		_w28928_,
		_w29073_
	);
	LUT2 #(
		.INIT('h1)
	) name18562 (
		_w28929_,
		_w28930_,
		_w29074_
	);
	LUT2 #(
		.INIT('h1)
	) name18563 (
		_w28931_,
		_w28932_,
		_w29075_
	);
	LUT2 #(
		.INIT('h1)
	) name18564 (
		_w28933_,
		_w28934_,
		_w29076_
	);
	LUT2 #(
		.INIT('h1)
	) name18565 (
		_w28935_,
		_w28936_,
		_w29077_
	);
	LUT2 #(
		.INIT('h1)
	) name18566 (
		_w28937_,
		_w28938_,
		_w29078_
	);
	LUT2 #(
		.INIT('h1)
	) name18567 (
		_w28939_,
		_w28940_,
		_w29079_
	);
	LUT2 #(
		.INIT('h1)
	) name18568 (
		_w28941_,
		_w28942_,
		_w29080_
	);
	LUT2 #(
		.INIT('h1)
	) name18569 (
		_w28943_,
		_w28944_,
		_w29081_
	);
	LUT2 #(
		.INIT('h1)
	) name18570 (
		_w28945_,
		_w28946_,
		_w29082_
	);
	LUT2 #(
		.INIT('h1)
	) name18571 (
		_w28947_,
		_w28948_,
		_w29083_
	);
	LUT2 #(
		.INIT('h1)
	) name18572 (
		_w28949_,
		_w28950_,
		_w29084_
	);
	LUT2 #(
		.INIT('h1)
	) name18573 (
		_w28951_,
		_w28952_,
		_w29085_
	);
	LUT2 #(
		.INIT('h1)
	) name18574 (
		_w28953_,
		_w28954_,
		_w29086_
	);
	LUT2 #(
		.INIT('h1)
	) name18575 (
		_w28955_,
		_w28956_,
		_w29087_
	);
	LUT2 #(
		.INIT('h1)
	) name18576 (
		_w28957_,
		_w28958_,
		_w29088_
	);
	LUT2 #(
		.INIT('h1)
	) name18577 (
		_w28959_,
		_w28960_,
		_w29089_
	);
	LUT2 #(
		.INIT('h1)
	) name18578 (
		_w28961_,
		_w28962_,
		_w29090_
	);
	LUT2 #(
		.INIT('h8)
	) name18579 (
		_w29089_,
		_w29090_,
		_w29091_
	);
	LUT2 #(
		.INIT('h8)
	) name18580 (
		_w29087_,
		_w29088_,
		_w29092_
	);
	LUT2 #(
		.INIT('h8)
	) name18581 (
		_w29085_,
		_w29086_,
		_w29093_
	);
	LUT2 #(
		.INIT('h8)
	) name18582 (
		_w29083_,
		_w29084_,
		_w29094_
	);
	LUT2 #(
		.INIT('h8)
	) name18583 (
		_w29081_,
		_w29082_,
		_w29095_
	);
	LUT2 #(
		.INIT('h8)
	) name18584 (
		_w29079_,
		_w29080_,
		_w29096_
	);
	LUT2 #(
		.INIT('h8)
	) name18585 (
		_w29077_,
		_w29078_,
		_w29097_
	);
	LUT2 #(
		.INIT('h8)
	) name18586 (
		_w29075_,
		_w29076_,
		_w29098_
	);
	LUT2 #(
		.INIT('h8)
	) name18587 (
		_w29073_,
		_w29074_,
		_w29099_
	);
	LUT2 #(
		.INIT('h8)
	) name18588 (
		_w29071_,
		_w29072_,
		_w29100_
	);
	LUT2 #(
		.INIT('h8)
	) name18589 (
		_w29069_,
		_w29070_,
		_w29101_
	);
	LUT2 #(
		.INIT('h8)
	) name18590 (
		_w29067_,
		_w29068_,
		_w29102_
	);
	LUT2 #(
		.INIT('h8)
	) name18591 (
		_w29065_,
		_w29066_,
		_w29103_
	);
	LUT2 #(
		.INIT('h8)
	) name18592 (
		_w29063_,
		_w29064_,
		_w29104_
	);
	LUT2 #(
		.INIT('h8)
	) name18593 (
		_w29061_,
		_w29062_,
		_w29105_
	);
	LUT2 #(
		.INIT('h8)
	) name18594 (
		_w29059_,
		_w29060_,
		_w29106_
	);
	LUT2 #(
		.INIT('h8)
	) name18595 (
		_w29057_,
		_w29058_,
		_w29107_
	);
	LUT2 #(
		.INIT('h8)
	) name18596 (
		_w29055_,
		_w29056_,
		_w29108_
	);
	LUT2 #(
		.INIT('h8)
	) name18597 (
		_w29053_,
		_w29054_,
		_w29109_
	);
	LUT2 #(
		.INIT('h8)
	) name18598 (
		_w29051_,
		_w29052_,
		_w29110_
	);
	LUT2 #(
		.INIT('h8)
	) name18599 (
		_w29049_,
		_w29050_,
		_w29111_
	);
	LUT2 #(
		.INIT('h8)
	) name18600 (
		_w29047_,
		_w29048_,
		_w29112_
	);
	LUT2 #(
		.INIT('h8)
	) name18601 (
		_w29045_,
		_w29046_,
		_w29113_
	);
	LUT2 #(
		.INIT('h8)
	) name18602 (
		_w29043_,
		_w29044_,
		_w29114_
	);
	LUT2 #(
		.INIT('h8)
	) name18603 (
		_w29041_,
		_w29042_,
		_w29115_
	);
	LUT2 #(
		.INIT('h8)
	) name18604 (
		_w29039_,
		_w29040_,
		_w29116_
	);
	LUT2 #(
		.INIT('h8)
	) name18605 (
		_w29037_,
		_w29038_,
		_w29117_
	);
	LUT2 #(
		.INIT('h8)
	) name18606 (
		_w29035_,
		_w29036_,
		_w29118_
	);
	LUT2 #(
		.INIT('h8)
	) name18607 (
		_w29033_,
		_w29034_,
		_w29119_
	);
	LUT2 #(
		.INIT('h8)
	) name18608 (
		_w29031_,
		_w29032_,
		_w29120_
	);
	LUT2 #(
		.INIT('h8)
	) name18609 (
		_w29029_,
		_w29030_,
		_w29121_
	);
	LUT2 #(
		.INIT('h8)
	) name18610 (
		_w29027_,
		_w29028_,
		_w29122_
	);
	LUT2 #(
		.INIT('h8)
	) name18611 (
		_w29025_,
		_w29026_,
		_w29123_
	);
	LUT2 #(
		.INIT('h8)
	) name18612 (
		_w29023_,
		_w29024_,
		_w29124_
	);
	LUT2 #(
		.INIT('h8)
	) name18613 (
		_w29021_,
		_w29022_,
		_w29125_
	);
	LUT2 #(
		.INIT('h8)
	) name18614 (
		_w29019_,
		_w29020_,
		_w29126_
	);
	LUT2 #(
		.INIT('h8)
	) name18615 (
		_w29017_,
		_w29018_,
		_w29127_
	);
	LUT2 #(
		.INIT('h8)
	) name18616 (
		_w29015_,
		_w29016_,
		_w29128_
	);
	LUT2 #(
		.INIT('h8)
	) name18617 (
		_w29013_,
		_w29014_,
		_w29129_
	);
	LUT2 #(
		.INIT('h8)
	) name18618 (
		_w29011_,
		_w29012_,
		_w29130_
	);
	LUT2 #(
		.INIT('h8)
	) name18619 (
		_w29009_,
		_w29010_,
		_w29131_
	);
	LUT2 #(
		.INIT('h8)
	) name18620 (
		_w29007_,
		_w29008_,
		_w29132_
	);
	LUT2 #(
		.INIT('h8)
	) name18621 (
		_w29005_,
		_w29006_,
		_w29133_
	);
	LUT2 #(
		.INIT('h8)
	) name18622 (
		_w29003_,
		_w29004_,
		_w29134_
	);
	LUT2 #(
		.INIT('h8)
	) name18623 (
		_w29001_,
		_w29002_,
		_w29135_
	);
	LUT2 #(
		.INIT('h8)
	) name18624 (
		_w28999_,
		_w29000_,
		_w29136_
	);
	LUT2 #(
		.INIT('h8)
	) name18625 (
		_w28997_,
		_w28998_,
		_w29137_
	);
	LUT2 #(
		.INIT('h8)
	) name18626 (
		_w28995_,
		_w28996_,
		_w29138_
	);
	LUT2 #(
		.INIT('h8)
	) name18627 (
		_w28993_,
		_w28994_,
		_w29139_
	);
	LUT2 #(
		.INIT('h8)
	) name18628 (
		_w28991_,
		_w28992_,
		_w29140_
	);
	LUT2 #(
		.INIT('h8)
	) name18629 (
		_w28989_,
		_w28990_,
		_w29141_
	);
	LUT2 #(
		.INIT('h8)
	) name18630 (
		_w28987_,
		_w28988_,
		_w29142_
	);
	LUT2 #(
		.INIT('h8)
	) name18631 (
		_w28985_,
		_w28986_,
		_w29143_
	);
	LUT2 #(
		.INIT('h8)
	) name18632 (
		_w28983_,
		_w28984_,
		_w29144_
	);
	LUT2 #(
		.INIT('h8)
	) name18633 (
		_w28981_,
		_w28982_,
		_w29145_
	);
	LUT2 #(
		.INIT('h8)
	) name18634 (
		_w28979_,
		_w28980_,
		_w29146_
	);
	LUT2 #(
		.INIT('h8)
	) name18635 (
		_w28977_,
		_w28978_,
		_w29147_
	);
	LUT2 #(
		.INIT('h8)
	) name18636 (
		_w28975_,
		_w28976_,
		_w29148_
	);
	LUT2 #(
		.INIT('h8)
	) name18637 (
		_w28973_,
		_w28974_,
		_w29149_
	);
	LUT2 #(
		.INIT('h8)
	) name18638 (
		_w28971_,
		_w28972_,
		_w29150_
	);
	LUT2 #(
		.INIT('h8)
	) name18639 (
		_w28969_,
		_w28970_,
		_w29151_
	);
	LUT2 #(
		.INIT('h8)
	) name18640 (
		_w28967_,
		_w28968_,
		_w29152_
	);
	LUT2 #(
		.INIT('h8)
	) name18641 (
		_w28965_,
		_w28966_,
		_w29153_
	);
	LUT2 #(
		.INIT('h8)
	) name18642 (
		_w28963_,
		_w28964_,
		_w29154_
	);
	LUT2 #(
		.INIT('h8)
	) name18643 (
		_w29153_,
		_w29154_,
		_w29155_
	);
	LUT2 #(
		.INIT('h8)
	) name18644 (
		_w29151_,
		_w29152_,
		_w29156_
	);
	LUT2 #(
		.INIT('h8)
	) name18645 (
		_w29149_,
		_w29150_,
		_w29157_
	);
	LUT2 #(
		.INIT('h8)
	) name18646 (
		_w29147_,
		_w29148_,
		_w29158_
	);
	LUT2 #(
		.INIT('h8)
	) name18647 (
		_w29145_,
		_w29146_,
		_w29159_
	);
	LUT2 #(
		.INIT('h8)
	) name18648 (
		_w29143_,
		_w29144_,
		_w29160_
	);
	LUT2 #(
		.INIT('h8)
	) name18649 (
		_w29141_,
		_w29142_,
		_w29161_
	);
	LUT2 #(
		.INIT('h8)
	) name18650 (
		_w29139_,
		_w29140_,
		_w29162_
	);
	LUT2 #(
		.INIT('h8)
	) name18651 (
		_w29137_,
		_w29138_,
		_w29163_
	);
	LUT2 #(
		.INIT('h8)
	) name18652 (
		_w29135_,
		_w29136_,
		_w29164_
	);
	LUT2 #(
		.INIT('h8)
	) name18653 (
		_w29133_,
		_w29134_,
		_w29165_
	);
	LUT2 #(
		.INIT('h8)
	) name18654 (
		_w29131_,
		_w29132_,
		_w29166_
	);
	LUT2 #(
		.INIT('h8)
	) name18655 (
		_w29129_,
		_w29130_,
		_w29167_
	);
	LUT2 #(
		.INIT('h8)
	) name18656 (
		_w29127_,
		_w29128_,
		_w29168_
	);
	LUT2 #(
		.INIT('h8)
	) name18657 (
		_w29125_,
		_w29126_,
		_w29169_
	);
	LUT2 #(
		.INIT('h8)
	) name18658 (
		_w29123_,
		_w29124_,
		_w29170_
	);
	LUT2 #(
		.INIT('h8)
	) name18659 (
		_w29121_,
		_w29122_,
		_w29171_
	);
	LUT2 #(
		.INIT('h8)
	) name18660 (
		_w29119_,
		_w29120_,
		_w29172_
	);
	LUT2 #(
		.INIT('h8)
	) name18661 (
		_w29117_,
		_w29118_,
		_w29173_
	);
	LUT2 #(
		.INIT('h8)
	) name18662 (
		_w29115_,
		_w29116_,
		_w29174_
	);
	LUT2 #(
		.INIT('h8)
	) name18663 (
		_w29113_,
		_w29114_,
		_w29175_
	);
	LUT2 #(
		.INIT('h8)
	) name18664 (
		_w29111_,
		_w29112_,
		_w29176_
	);
	LUT2 #(
		.INIT('h8)
	) name18665 (
		_w29109_,
		_w29110_,
		_w29177_
	);
	LUT2 #(
		.INIT('h8)
	) name18666 (
		_w29107_,
		_w29108_,
		_w29178_
	);
	LUT2 #(
		.INIT('h8)
	) name18667 (
		_w29105_,
		_w29106_,
		_w29179_
	);
	LUT2 #(
		.INIT('h8)
	) name18668 (
		_w29103_,
		_w29104_,
		_w29180_
	);
	LUT2 #(
		.INIT('h8)
	) name18669 (
		_w29101_,
		_w29102_,
		_w29181_
	);
	LUT2 #(
		.INIT('h8)
	) name18670 (
		_w29099_,
		_w29100_,
		_w29182_
	);
	LUT2 #(
		.INIT('h8)
	) name18671 (
		_w29097_,
		_w29098_,
		_w29183_
	);
	LUT2 #(
		.INIT('h8)
	) name18672 (
		_w29095_,
		_w29096_,
		_w29184_
	);
	LUT2 #(
		.INIT('h8)
	) name18673 (
		_w29093_,
		_w29094_,
		_w29185_
	);
	LUT2 #(
		.INIT('h8)
	) name18674 (
		_w29091_,
		_w29092_,
		_w29186_
	);
	LUT2 #(
		.INIT('h8)
	) name18675 (
		_w29185_,
		_w29186_,
		_w29187_
	);
	LUT2 #(
		.INIT('h8)
	) name18676 (
		_w29183_,
		_w29184_,
		_w29188_
	);
	LUT2 #(
		.INIT('h8)
	) name18677 (
		_w29181_,
		_w29182_,
		_w29189_
	);
	LUT2 #(
		.INIT('h8)
	) name18678 (
		_w29179_,
		_w29180_,
		_w29190_
	);
	LUT2 #(
		.INIT('h8)
	) name18679 (
		_w29177_,
		_w29178_,
		_w29191_
	);
	LUT2 #(
		.INIT('h8)
	) name18680 (
		_w29175_,
		_w29176_,
		_w29192_
	);
	LUT2 #(
		.INIT('h8)
	) name18681 (
		_w29173_,
		_w29174_,
		_w29193_
	);
	LUT2 #(
		.INIT('h8)
	) name18682 (
		_w29171_,
		_w29172_,
		_w29194_
	);
	LUT2 #(
		.INIT('h8)
	) name18683 (
		_w29169_,
		_w29170_,
		_w29195_
	);
	LUT2 #(
		.INIT('h8)
	) name18684 (
		_w29167_,
		_w29168_,
		_w29196_
	);
	LUT2 #(
		.INIT('h8)
	) name18685 (
		_w29165_,
		_w29166_,
		_w29197_
	);
	LUT2 #(
		.INIT('h8)
	) name18686 (
		_w29163_,
		_w29164_,
		_w29198_
	);
	LUT2 #(
		.INIT('h8)
	) name18687 (
		_w29161_,
		_w29162_,
		_w29199_
	);
	LUT2 #(
		.INIT('h8)
	) name18688 (
		_w29159_,
		_w29160_,
		_w29200_
	);
	LUT2 #(
		.INIT('h8)
	) name18689 (
		_w29157_,
		_w29158_,
		_w29201_
	);
	LUT2 #(
		.INIT('h8)
	) name18690 (
		_w29155_,
		_w29156_,
		_w29202_
	);
	LUT2 #(
		.INIT('h8)
	) name18691 (
		_w29201_,
		_w29202_,
		_w29203_
	);
	LUT2 #(
		.INIT('h8)
	) name18692 (
		_w29199_,
		_w29200_,
		_w29204_
	);
	LUT2 #(
		.INIT('h8)
	) name18693 (
		_w29197_,
		_w29198_,
		_w29205_
	);
	LUT2 #(
		.INIT('h8)
	) name18694 (
		_w29195_,
		_w29196_,
		_w29206_
	);
	LUT2 #(
		.INIT('h8)
	) name18695 (
		_w29193_,
		_w29194_,
		_w29207_
	);
	LUT2 #(
		.INIT('h8)
	) name18696 (
		_w29191_,
		_w29192_,
		_w29208_
	);
	LUT2 #(
		.INIT('h8)
	) name18697 (
		_w29189_,
		_w29190_,
		_w29209_
	);
	LUT2 #(
		.INIT('h8)
	) name18698 (
		_w29187_,
		_w29188_,
		_w29210_
	);
	LUT2 #(
		.INIT('h8)
	) name18699 (
		_w29209_,
		_w29210_,
		_w29211_
	);
	LUT2 #(
		.INIT('h8)
	) name18700 (
		_w29207_,
		_w29208_,
		_w29212_
	);
	LUT2 #(
		.INIT('h8)
	) name18701 (
		_w29205_,
		_w29206_,
		_w29213_
	);
	LUT2 #(
		.INIT('h8)
	) name18702 (
		_w29203_,
		_w29204_,
		_w29214_
	);
	LUT2 #(
		.INIT('h8)
	) name18703 (
		_w29213_,
		_w29214_,
		_w29215_
	);
	LUT2 #(
		.INIT('h8)
	) name18704 (
		_w29211_,
		_w29212_,
		_w29216_
	);
	LUT2 #(
		.INIT('h8)
	) name18705 (
		_w29215_,
		_w29216_,
		_w29217_
	);
	LUT2 #(
		.INIT('h1)
	) name18706 (
		wb_rst_i_pad,
		_w29217_,
		_w29218_
	);
	LUT2 #(
		.INIT('h1)
	) name18707 (
		_w22944_,
		_w29218_,
		_w29219_
	);
	LUT2 #(
		.INIT('h8)
	) name18708 (
		\ethreg1_IPGT_0_DataOut_reg[6]/NET0131 ,
		_w24717_,
		_w29220_
	);
	LUT2 #(
		.INIT('h8)
	) name18709 (
		\ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 ,
		_w22956_,
		_w29221_
	);
	LUT2 #(
		.INIT('h8)
	) name18710 (
		\ethreg1_IPGR2_0_DataOut_reg[6]/NET0131 ,
		_w24724_,
		_w29222_
	);
	LUT2 #(
		.INIT('h8)
	) name18711 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		_w24726_,
		_w29223_
	);
	LUT2 #(
		.INIT('h8)
	) name18712 (
		\ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 ,
		_w22952_,
		_w29224_
	);
	LUT2 #(
		.INIT('h8)
	) name18713 (
		\ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 ,
		_w24722_,
		_w29225_
	);
	LUT2 #(
		.INIT('h8)
	) name18714 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		_w22959_,
		_w29226_
	);
	LUT2 #(
		.INIT('h8)
	) name18715 (
		\ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 ,
		_w23499_,
		_w29227_
	);
	LUT2 #(
		.INIT('h8)
	) name18716 (
		\ethreg1_IPGR1_0_DataOut_reg[6]/NET0131 ,
		_w24710_,
		_w29228_
	);
	LUT2 #(
		.INIT('h8)
	) name18717 (
		\ethreg1_PACKETLEN_0_DataOut_reg[6]/NET0131 ,
		_w22966_,
		_w29229_
	);
	LUT2 #(
		.INIT('h8)
	) name18718 (
		\ethreg1_MODER_0_DataOut_reg[6]/NET0131 ,
		_w23519_,
		_w29230_
	);
	LUT2 #(
		.INIT('h8)
	) name18719 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		_w24713_,
		_w29231_
	);
	LUT2 #(
		.INIT('h8)
	) name18720 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		_w23501_,
		_w29232_
	);
	LUT2 #(
		.INIT('h8)
	) name18721 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 ,
		_w23522_,
		_w29233_
	);
	LUT2 #(
		.INIT('h8)
	) name18722 (
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w24707_,
		_w29234_
	);
	LUT2 #(
		.INIT('h8)
	) name18723 (
		\ethreg1_MIIRX_DATA_DataOut_reg[6]/NET0131 ,
		_w23507_,
		_w29235_
	);
	LUT2 #(
		.INIT('h1)
	) name18724 (
		_w29220_,
		_w29221_,
		_w29236_
	);
	LUT2 #(
		.INIT('h1)
	) name18725 (
		_w29222_,
		_w29223_,
		_w29237_
	);
	LUT2 #(
		.INIT('h1)
	) name18726 (
		_w29224_,
		_w29225_,
		_w29238_
	);
	LUT2 #(
		.INIT('h1)
	) name18727 (
		_w29226_,
		_w29227_,
		_w29239_
	);
	LUT2 #(
		.INIT('h1)
	) name18728 (
		_w29228_,
		_w29230_,
		_w29240_
	);
	LUT2 #(
		.INIT('h1)
	) name18729 (
		_w29231_,
		_w29232_,
		_w29241_
	);
	LUT2 #(
		.INIT('h1)
	) name18730 (
		_w29233_,
		_w29234_,
		_w29242_
	);
	LUT2 #(
		.INIT('h4)
	) name18731 (
		_w29235_,
		_w29242_,
		_w29243_
	);
	LUT2 #(
		.INIT('h8)
	) name18732 (
		_w29240_,
		_w29241_,
		_w29244_
	);
	LUT2 #(
		.INIT('h8)
	) name18733 (
		_w29238_,
		_w29239_,
		_w29245_
	);
	LUT2 #(
		.INIT('h8)
	) name18734 (
		_w29236_,
		_w29237_,
		_w29246_
	);
	LUT2 #(
		.INIT('h8)
	) name18735 (
		_w22944_,
		_w29246_,
		_w29247_
	);
	LUT2 #(
		.INIT('h8)
	) name18736 (
		_w29244_,
		_w29245_,
		_w29248_
	);
	LUT2 #(
		.INIT('h4)
	) name18737 (
		_w29229_,
		_w29243_,
		_w29249_
	);
	LUT2 #(
		.INIT('h8)
	) name18738 (
		_w29248_,
		_w29249_,
		_w29250_
	);
	LUT2 #(
		.INIT('h8)
	) name18739 (
		_w29247_,
		_w29250_,
		_w29251_
	);
	LUT2 #(
		.INIT('h1)
	) name18740 (
		_w29219_,
		_w29251_,
		_w29252_
	);
	LUT2 #(
		.INIT('h1)
	) name18741 (
		_w20126_,
		_w22944_,
		_w29253_
	);
	LUT2 #(
		.INIT('h8)
	) name18742 (
		\ethreg1_COLLCONF_2_DataOut_reg[1]/NET0131 ,
		_w24730_,
		_w29254_
	);
	LUT2 #(
		.INIT('h8)
	) name18743 (
		\ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 ,
		_w22956_,
		_w29255_
	);
	LUT2 #(
		.INIT('h8)
	) name18744 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		_w22959_,
		_w29256_
	);
	LUT2 #(
		.INIT('h8)
	) name18745 (
		\ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 ,
		_w22952_,
		_w29257_
	);
	LUT2 #(
		.INIT('h8)
	) name18746 (
		\ethreg1_PACKETLEN_2_DataOut_reg[1]/NET0131 ,
		_w22966_,
		_w29258_
	);
	LUT2 #(
		.INIT('h1)
	) name18747 (
		_w29255_,
		_w29256_,
		_w29259_
	);
	LUT2 #(
		.INIT('h4)
	) name18748 (
		_w29257_,
		_w29259_,
		_w29260_
	);
	LUT2 #(
		.INIT('h8)
	) name18749 (
		_w22944_,
		_w29260_,
		_w29261_
	);
	LUT2 #(
		.INIT('h1)
	) name18750 (
		_w29254_,
		_w29258_,
		_w29262_
	);
	LUT2 #(
		.INIT('h8)
	) name18751 (
		_w29261_,
		_w29262_,
		_w29263_
	);
	LUT2 #(
		.INIT('h1)
	) name18752 (
		_w29253_,
		_w29263_,
		_w29264_
	);
	LUT2 #(
		.INIT('h1)
	) name18753 (
		_w18564_,
		_w22944_,
		_w29265_
	);
	LUT2 #(
		.INIT('h8)
	) name18754 (
		\ethreg1_COLLCONF_2_DataOut_reg[2]/NET0131 ,
		_w24730_,
		_w29266_
	);
	LUT2 #(
		.INIT('h8)
	) name18755 (
		\ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 ,
		_w22956_,
		_w29267_
	);
	LUT2 #(
		.INIT('h8)
	) name18756 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		_w22959_,
		_w29268_
	);
	LUT2 #(
		.INIT('h8)
	) name18757 (
		\ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 ,
		_w22952_,
		_w29269_
	);
	LUT2 #(
		.INIT('h8)
	) name18758 (
		\ethreg1_PACKETLEN_2_DataOut_reg[2]/NET0131 ,
		_w22966_,
		_w29270_
	);
	LUT2 #(
		.INIT('h1)
	) name18759 (
		_w29267_,
		_w29268_,
		_w29271_
	);
	LUT2 #(
		.INIT('h4)
	) name18760 (
		_w29269_,
		_w29271_,
		_w29272_
	);
	LUT2 #(
		.INIT('h8)
	) name18761 (
		_w22944_,
		_w29272_,
		_w29273_
	);
	LUT2 #(
		.INIT('h1)
	) name18762 (
		_w29266_,
		_w29270_,
		_w29274_
	);
	LUT2 #(
		.INIT('h8)
	) name18763 (
		_w29273_,
		_w29274_,
		_w29275_
	);
	LUT2 #(
		.INIT('h1)
	) name18764 (
		_w29265_,
		_w29275_,
		_w29276_
	);
	LUT2 #(
		.INIT('h1)
	) name18765 (
		_w21383_,
		_w22944_,
		_w29277_
	);
	LUT2 #(
		.INIT('h8)
	) name18766 (
		\ethreg1_COLLCONF_2_DataOut_reg[3]/NET0131 ,
		_w24730_,
		_w29278_
	);
	LUT2 #(
		.INIT('h8)
	) name18767 (
		\ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 ,
		_w22956_,
		_w29279_
	);
	LUT2 #(
		.INIT('h8)
	) name18768 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		_w22959_,
		_w29280_
	);
	LUT2 #(
		.INIT('h8)
	) name18769 (
		\ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 ,
		_w22952_,
		_w29281_
	);
	LUT2 #(
		.INIT('h8)
	) name18770 (
		\ethreg1_PACKETLEN_2_DataOut_reg[3]/NET0131 ,
		_w22966_,
		_w29282_
	);
	LUT2 #(
		.INIT('h1)
	) name18771 (
		_w29279_,
		_w29280_,
		_w29283_
	);
	LUT2 #(
		.INIT('h4)
	) name18772 (
		_w29281_,
		_w29283_,
		_w29284_
	);
	LUT2 #(
		.INIT('h8)
	) name18773 (
		_w22944_,
		_w29284_,
		_w29285_
	);
	LUT2 #(
		.INIT('h1)
	) name18774 (
		_w29278_,
		_w29282_,
		_w29286_
	);
	LUT2 #(
		.INIT('h8)
	) name18775 (
		_w29285_,
		_w29286_,
		_w29287_
	);
	LUT2 #(
		.INIT('h1)
	) name18776 (
		_w29277_,
		_w29287_,
		_w29288_
	);
	LUT2 #(
		.INIT('h8)
	) name18777 (
		_w15696_,
		_w21383_,
		_w29289_
	);
	LUT2 #(
		.INIT('h8)
	) name18778 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w17862_,
		_w29290_
	);
	LUT2 #(
		.INIT('h8)
	) name18779 (
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w29290_,
		_w29291_
	);
	LUT2 #(
		.INIT('h8)
	) name18780 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		_w29291_,
		_w29292_
	);
	LUT2 #(
		.INIT('h1)
	) name18781 (
		\wishbone_RxPointerMSB_reg[19]/NET0131 ,
		_w29292_,
		_w29293_
	);
	LUT2 #(
		.INIT('h1)
	) name18782 (
		_w15696_,
		_w17866_,
		_w29294_
	);
	LUT2 #(
		.INIT('h4)
	) name18783 (
		_w29293_,
		_w29294_,
		_w29295_
	);
	LUT2 #(
		.INIT('h1)
	) name18784 (
		_w29289_,
		_w29295_,
		_w29296_
	);
	LUT2 #(
		.INIT('h1)
	) name18785 (
		\wishbone_RxPointerMSB_reg[20]/NET0131 ,
		_w17866_,
		_w29297_
	);
	LUT2 #(
		.INIT('h1)
	) name18786 (
		_w15696_,
		_w17867_,
		_w29298_
	);
	LUT2 #(
		.INIT('h4)
	) name18787 (
		_w29297_,
		_w29298_,
		_w29299_
	);
	LUT2 #(
		.INIT('h8)
	) name18788 (
		_w15696_,
		_w16743_,
		_w29300_
	);
	LUT2 #(
		.INIT('h1)
	) name18789 (
		_w29299_,
		_w29300_,
		_w29301_
	);
	LUT2 #(
		.INIT('h8)
	) name18790 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		_w17867_,
		_w29302_
	);
	LUT2 #(
		.INIT('h1)
	) name18791 (
		\wishbone_RxPointerMSB_reg[21]/NET0131 ,
		_w17867_,
		_w29303_
	);
	LUT2 #(
		.INIT('h1)
	) name18792 (
		_w15696_,
		_w29302_,
		_w29304_
	);
	LUT2 #(
		.INIT('h4)
	) name18793 (
		_w29303_,
		_w29304_,
		_w29305_
	);
	LUT2 #(
		.INIT('h8)
	) name18794 (
		_w15696_,
		_w21900_,
		_w29306_
	);
	LUT2 #(
		.INIT('h1)
	) name18795 (
		_w29305_,
		_w29306_,
		_w29307_
	);
	LUT2 #(
		.INIT('h8)
	) name18796 (
		_w15696_,
		_w22932_,
		_w29308_
	);
	LUT2 #(
		.INIT('h1)
	) name18797 (
		\wishbone_RxPointerMSB_reg[22]/NET0131 ,
		_w29302_,
		_w29309_
	);
	LUT2 #(
		.INIT('h1)
	) name18798 (
		_w15696_,
		_w17869_,
		_w29310_
	);
	LUT2 #(
		.INIT('h4)
	) name18799 (
		_w29309_,
		_w29310_,
		_w29311_
	);
	LUT2 #(
		.INIT('h1)
	) name18800 (
		_w29308_,
		_w29311_,
		_w29312_
	);
	LUT2 #(
		.INIT('h1)
	) name18801 (
		\wishbone_RxPointerMSB_reg[23]/NET0131 ,
		_w17869_,
		_w29313_
	);
	LUT2 #(
		.INIT('h1)
	) name18802 (
		_w15696_,
		_w17870_,
		_w29314_
	);
	LUT2 #(
		.INIT('h4)
	) name18803 (
		_w29313_,
		_w29314_,
		_w29315_
	);
	LUT2 #(
		.INIT('h8)
	) name18804 (
		_w15696_,
		_w22415_,
		_w29316_
	);
	LUT2 #(
		.INIT('h1)
	) name18805 (
		_w29315_,
		_w29316_,
		_w29317_
	);
	LUT2 #(
		.INIT('h1)
	) name18806 (
		\wishbone_RxPointerMSB_reg[24]/NET0131 ,
		_w17870_,
		_w29318_
	);
	LUT2 #(
		.INIT('h1)
	) name18807 (
		_w15696_,
		_w17871_,
		_w29319_
	);
	LUT2 #(
		.INIT('h4)
	) name18808 (
		_w29318_,
		_w29319_,
		_w29320_
	);
	LUT2 #(
		.INIT('h8)
	) name18809 (
		_w15110_,
		_w15696_,
		_w29321_
	);
	LUT2 #(
		.INIT('h1)
	) name18810 (
		_w29320_,
		_w29321_,
		_w29322_
	);
	LUT2 #(
		.INIT('h1)
	) name18811 (
		\wishbone_RxPointerMSB_reg[25]/NET0131 ,
		_w17871_,
		_w29323_
	);
	LUT2 #(
		.INIT('h1)
	) name18812 (
		_w15696_,
		_w17872_,
		_w29324_
	);
	LUT2 #(
		.INIT('h4)
	) name18813 (
		_w29323_,
		_w29324_,
		_w29325_
	);
	LUT2 #(
		.INIT('h8)
	) name18814 (
		_w15696_,
		_w17810_,
		_w29326_
	);
	LUT2 #(
		.INIT('h1)
	) name18815 (
		_w29325_,
		_w29326_,
		_w29327_
	);
	LUT2 #(
		.INIT('h1)
	) name18816 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		_w17872_,
		_w29328_
	);
	LUT2 #(
		.INIT('h8)
	) name18817 (
		\wishbone_RxPointerMSB_reg[26]/NET0131 ,
		_w17872_,
		_w29329_
	);
	LUT2 #(
		.INIT('h1)
	) name18818 (
		_w15696_,
		_w29328_,
		_w29330_
	);
	LUT2 #(
		.INIT('h4)
	) name18819 (
		_w29329_,
		_w29330_,
		_w29331_
	);
	LUT2 #(
		.INIT('h8)
	) name18820 (
		_w15696_,
		_w17287_,
		_w29332_
	);
	LUT2 #(
		.INIT('h1)
	) name18821 (
		_w29331_,
		_w29332_,
		_w29333_
	);
	LUT2 #(
		.INIT('h1)
	) name18822 (
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w29329_,
		_w29334_
	);
	LUT2 #(
		.INIT('h8)
	) name18823 (
		\wishbone_RxPointerMSB_reg[27]/NET0131 ,
		_w29329_,
		_w29335_
	);
	LUT2 #(
		.INIT('h1)
	) name18824 (
		_w15696_,
		_w29334_,
		_w29336_
	);
	LUT2 #(
		.INIT('h4)
	) name18825 (
		_w29335_,
		_w29336_,
		_w29337_
	);
	LUT2 #(
		.INIT('h8)
	) name18826 (
		_w15696_,
		_w20856_,
		_w29338_
	);
	LUT2 #(
		.INIT('h1)
	) name18827 (
		_w29337_,
		_w29338_,
		_w29339_
	);
	LUT2 #(
		.INIT('h8)
	) name18828 (
		_w13475_,
		_w15696_,
		_w29340_
	);
	LUT2 #(
		.INIT('h1)
	) name18829 (
		\wishbone_RxPointerMSB_reg[28]/NET0131 ,
		_w29335_,
		_w29341_
	);
	LUT2 #(
		.INIT('h1)
	) name18830 (
		_w15696_,
		_w17875_,
		_w29342_
	);
	LUT2 #(
		.INIT('h4)
	) name18831 (
		_w29341_,
		_w29342_,
		_w29343_
	);
	LUT2 #(
		.INIT('h1)
	) name18832 (
		_w29340_,
		_w29343_,
		_w29344_
	);
	LUT2 #(
		.INIT('h1)
	) name18833 (
		\wishbone_RxPointerMSB_reg[29]/NET0131 ,
		_w17875_,
		_w29345_
	);
	LUT2 #(
		.INIT('h1)
	) name18834 (
		_w15696_,
		_w17876_,
		_w29346_
	);
	LUT2 #(
		.INIT('h4)
	) name18835 (
		_w29345_,
		_w29346_,
		_w29347_
	);
	LUT2 #(
		.INIT('h8)
	) name18836 (
		_w14019_,
		_w15696_,
		_w29348_
	);
	LUT2 #(
		.INIT('h1)
	) name18837 (
		_w29347_,
		_w29348_,
		_w29349_
	);
	LUT2 #(
		.INIT('h1)
	) name18838 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w17879_,
		_w29350_
	);
	LUT2 #(
		.INIT('h8)
	) name18839 (
		\wishbone_RxPointerMSB_reg[31]/NET0131 ,
		_w17879_,
		_w29351_
	);
	LUT2 #(
		.INIT('h1)
	) name18840 (
		_w29350_,
		_w29351_,
		_w29352_
	);
	LUT2 #(
		.INIT('h1)
	) name18841 (
		_w15696_,
		_w29352_,
		_w29353_
	);
	LUT2 #(
		.INIT('h2)
	) name18842 (
		_w15696_,
		_w19604_,
		_w29354_
	);
	LUT2 #(
		.INIT('h1)
	) name18843 (
		_w29353_,
		_w29354_,
		_w29355_
	);
	LUT2 #(
		.INIT('h8)
	) name18844 (
		_w15696_,
		_w27436_,
		_w29356_
	);
	LUT2 #(
		.INIT('h8)
	) name18845 (
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w17854_,
		_w29357_
	);
	LUT2 #(
		.INIT('h1)
	) name18846 (
		\wishbone_RxPointerMSB_reg[9]/NET0131 ,
		_w29357_,
		_w29358_
	);
	LUT2 #(
		.INIT('h1)
	) name18847 (
		_w15696_,
		_w17856_,
		_w29359_
	);
	LUT2 #(
		.INIT('h4)
	) name18848 (
		_w29358_,
		_w29359_,
		_w29360_
	);
	LUT2 #(
		.INIT('h1)
	) name18849 (
		_w29356_,
		_w29360_,
		_w29361_
	);
	LUT2 #(
		.INIT('h1)
	) name18850 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w17902_,
		_w29362_
	);
	LUT2 #(
		.INIT('h8)
	) name18851 (
		\wishbone_TxPointerMSB_reg[19]/NET0131 ,
		_w17902_,
		_w29363_
	);
	LUT2 #(
		.INIT('h1)
	) name18852 (
		_w17883_,
		_w29362_,
		_w29364_
	);
	LUT2 #(
		.INIT('h4)
	) name18853 (
		_w29363_,
		_w29364_,
		_w29365_
	);
	LUT2 #(
		.INIT('h8)
	) name18854 (
		_w17883_,
		_w21383_,
		_w29366_
	);
	LUT2 #(
		.INIT('h1)
	) name18855 (
		_w29365_,
		_w29366_,
		_w29367_
	);
	LUT2 #(
		.INIT('h8)
	) name18856 (
		_w16743_,
		_w17883_,
		_w29368_
	);
	LUT2 #(
		.INIT('h1)
	) name18857 (
		\wishbone_TxPointerMSB_reg[20]/NET0131 ,
		_w29363_,
		_w29369_
	);
	LUT2 #(
		.INIT('h1)
	) name18858 (
		_w17883_,
		_w17904_,
		_w29370_
	);
	LUT2 #(
		.INIT('h4)
	) name18859 (
		_w29369_,
		_w29370_,
		_w29371_
	);
	LUT2 #(
		.INIT('h1)
	) name18860 (
		_w29368_,
		_w29371_,
		_w29372_
	);
	LUT2 #(
		.INIT('h1)
	) name18861 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w17904_,
		_w29373_
	);
	LUT2 #(
		.INIT('h8)
	) name18862 (
		\wishbone_TxPointerMSB_reg[21]/NET0131 ,
		_w17904_,
		_w29374_
	);
	LUT2 #(
		.INIT('h1)
	) name18863 (
		_w17883_,
		_w29373_,
		_w29375_
	);
	LUT2 #(
		.INIT('h4)
	) name18864 (
		_w29374_,
		_w29375_,
		_w29376_
	);
	LUT2 #(
		.INIT('h8)
	) name18865 (
		_w17883_,
		_w21900_,
		_w29377_
	);
	LUT2 #(
		.INIT('h1)
	) name18866 (
		_w29376_,
		_w29377_,
		_w29378_
	);
	LUT2 #(
		.INIT('h8)
	) name18867 (
		_w17883_,
		_w22932_,
		_w29379_
	);
	LUT2 #(
		.INIT('h1)
	) name18868 (
		\wishbone_TxPointerMSB_reg[22]/NET0131 ,
		_w29374_,
		_w29380_
	);
	LUT2 #(
		.INIT('h1)
	) name18869 (
		_w17883_,
		_w17906_,
		_w29381_
	);
	LUT2 #(
		.INIT('h4)
	) name18870 (
		_w29380_,
		_w29381_,
		_w29382_
	);
	LUT2 #(
		.INIT('h1)
	) name18871 (
		_w29379_,
		_w29382_,
		_w29383_
	);
	LUT2 #(
		.INIT('h1)
	) name18872 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		_w17906_,
		_w29384_
	);
	LUT2 #(
		.INIT('h8)
	) name18873 (
		\wishbone_TxPointerMSB_reg[23]/NET0131 ,
		_w17906_,
		_w29385_
	);
	LUT2 #(
		.INIT('h1)
	) name18874 (
		_w17883_,
		_w29384_,
		_w29386_
	);
	LUT2 #(
		.INIT('h4)
	) name18875 (
		_w29385_,
		_w29386_,
		_w29387_
	);
	LUT2 #(
		.INIT('h8)
	) name18876 (
		_w17883_,
		_w22415_,
		_w29388_
	);
	LUT2 #(
		.INIT('h1)
	) name18877 (
		_w29387_,
		_w29388_,
		_w29389_
	);
	LUT2 #(
		.INIT('h8)
	) name18878 (
		_w15110_,
		_w17883_,
		_w29390_
	);
	LUT2 #(
		.INIT('h1)
	) name18879 (
		\wishbone_TxPointerMSB_reg[24]/NET0131 ,
		_w29385_,
		_w29391_
	);
	LUT2 #(
		.INIT('h1)
	) name18880 (
		_w17883_,
		_w17908_,
		_w29392_
	);
	LUT2 #(
		.INIT('h4)
	) name18881 (
		_w29391_,
		_w29392_,
		_w29393_
	);
	LUT2 #(
		.INIT('h1)
	) name18882 (
		_w29390_,
		_w29393_,
		_w29394_
	);
	LUT2 #(
		.INIT('h1)
	) name18883 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w17908_,
		_w29395_
	);
	LUT2 #(
		.INIT('h8)
	) name18884 (
		\wishbone_TxPointerMSB_reg[25]/NET0131 ,
		_w17908_,
		_w29396_
	);
	LUT2 #(
		.INIT('h1)
	) name18885 (
		_w17883_,
		_w29395_,
		_w29397_
	);
	LUT2 #(
		.INIT('h4)
	) name18886 (
		_w29396_,
		_w29397_,
		_w29398_
	);
	LUT2 #(
		.INIT('h8)
	) name18887 (
		_w17810_,
		_w17883_,
		_w29399_
	);
	LUT2 #(
		.INIT('h1)
	) name18888 (
		_w29398_,
		_w29399_,
		_w29400_
	);
	LUT2 #(
		.INIT('h8)
	) name18889 (
		_w17287_,
		_w17883_,
		_w29401_
	);
	LUT2 #(
		.INIT('h1)
	) name18890 (
		\wishbone_TxPointerMSB_reg[26]/NET0131 ,
		_w29396_,
		_w29402_
	);
	LUT2 #(
		.INIT('h1)
	) name18891 (
		_w17883_,
		_w17910_,
		_w29403_
	);
	LUT2 #(
		.INIT('h4)
	) name18892 (
		_w29402_,
		_w29403_,
		_w29404_
	);
	LUT2 #(
		.INIT('h1)
	) name18893 (
		_w29401_,
		_w29404_,
		_w29405_
	);
	LUT2 #(
		.INIT('h8)
	) name18894 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w17910_,
		_w29406_
	);
	LUT2 #(
		.INIT('h1)
	) name18895 (
		\wishbone_TxPointerMSB_reg[27]/NET0131 ,
		_w17910_,
		_w29407_
	);
	LUT2 #(
		.INIT('h1)
	) name18896 (
		_w17883_,
		_w29406_,
		_w29408_
	);
	LUT2 #(
		.INIT('h4)
	) name18897 (
		_w29407_,
		_w29408_,
		_w29409_
	);
	LUT2 #(
		.INIT('h8)
	) name18898 (
		_w17883_,
		_w20856_,
		_w29410_
	);
	LUT2 #(
		.INIT('h1)
	) name18899 (
		_w29409_,
		_w29410_,
		_w29411_
	);
	LUT2 #(
		.INIT('h2)
	) name18900 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		_w17911_,
		_w29412_
	);
	LUT2 #(
		.INIT('h4)
	) name18901 (
		\wishbone_TxPointerMSB_reg[29]/NET0131 ,
		_w17911_,
		_w29413_
	);
	LUT2 #(
		.INIT('h1)
	) name18902 (
		_w29412_,
		_w29413_,
		_w29414_
	);
	LUT2 #(
		.INIT('h1)
	) name18903 (
		_w17883_,
		_w29414_,
		_w29415_
	);
	LUT2 #(
		.INIT('h8)
	) name18904 (
		_w14019_,
		_w17883_,
		_w29416_
	);
	LUT2 #(
		.INIT('h1)
	) name18905 (
		_w29415_,
		_w29416_,
		_w29417_
	);
	LUT2 #(
		.INIT('h8)
	) name18906 (
		_w13475_,
		_w17883_,
		_w29418_
	);
	LUT2 #(
		.INIT('h1)
	) name18907 (
		\wishbone_TxPointerMSB_reg[28]/NET0131 ,
		_w29406_,
		_w29419_
	);
	LUT2 #(
		.INIT('h1)
	) name18908 (
		_w17883_,
		_w17911_,
		_w29420_
	);
	LUT2 #(
		.INIT('h4)
	) name18909 (
		_w29419_,
		_w29420_,
		_w29421_
	);
	LUT2 #(
		.INIT('h1)
	) name18910 (
		_w29418_,
		_w29421_,
		_w29422_
	);
	LUT2 #(
		.INIT('h8)
	) name18911 (
		_w17884_,
		_w17912_,
		_w29423_
	);
	LUT2 #(
		.INIT('h8)
	) name18912 (
		_w17910_,
		_w29423_,
		_w29424_
	);
	LUT2 #(
		.INIT('h2)
	) name18913 (
		\wishbone_TxPointerMSB_reg[31]/NET0131 ,
		_w29424_,
		_w29425_
	);
	LUT2 #(
		.INIT('h4)
	) name18914 (
		\wishbone_TxPointerMSB_reg[31]/NET0131 ,
		_w29424_,
		_w29426_
	);
	LUT2 #(
		.INIT('h1)
	) name18915 (
		_w29425_,
		_w29426_,
		_w29427_
	);
	LUT2 #(
		.INIT('h1)
	) name18916 (
		_w17883_,
		_w29427_,
		_w29428_
	);
	LUT2 #(
		.INIT('h8)
	) name18917 (
		_w17883_,
		_w19604_,
		_w29429_
	);
	LUT2 #(
		.INIT('h1)
	) name18918 (
		_w29428_,
		_w29429_,
		_w29430_
	);
	LUT2 #(
		.INIT('h1)
	) name18919 (
		\wishbone_TxPointerMSB_reg[9]/NET0131 ,
		_w17892_,
		_w29431_
	);
	LUT2 #(
		.INIT('h1)
	) name18920 (
		_w17883_,
		_w17893_,
		_w29432_
	);
	LUT2 #(
		.INIT('h4)
	) name18921 (
		_w29431_,
		_w29432_,
		_w29433_
	);
	LUT2 #(
		.INIT('h8)
	) name18922 (
		_w17883_,
		_w27436_,
		_w29434_
	);
	LUT2 #(
		.INIT('h1)
	) name18923 (
		_w29433_,
		_w29434_,
		_w29435_
	);
	LUT2 #(
		.INIT('h8)
	) name18924 (
		\wishbone_bd_ram_mem1_reg[85][13]/P0001 ,
		_w13216_,
		_w29436_
	);
	LUT2 #(
		.INIT('h8)
	) name18925 (
		\wishbone_bd_ram_mem1_reg[103][13]/P0001 ,
		_w12846_,
		_w29437_
	);
	LUT2 #(
		.INIT('h8)
	) name18926 (
		\wishbone_bd_ram_mem1_reg[114][13]/P0001 ,
		_w13202_,
		_w29438_
	);
	LUT2 #(
		.INIT('h8)
	) name18927 (
		\wishbone_bd_ram_mem1_reg[52][13]/P0001 ,
		_w13082_,
		_w29439_
	);
	LUT2 #(
		.INIT('h8)
	) name18928 (
		\wishbone_bd_ram_mem1_reg[34][13]/P0001 ,
		_w12930_,
		_w29440_
	);
	LUT2 #(
		.INIT('h8)
	) name18929 (
		\wishbone_bd_ram_mem1_reg[247][13]/P0001 ,
		_w12818_,
		_w29441_
	);
	LUT2 #(
		.INIT('h8)
	) name18930 (
		\wishbone_bd_ram_mem1_reg[131][13]/P0001 ,
		_w12852_,
		_w29442_
	);
	LUT2 #(
		.INIT('h8)
	) name18931 (
		\wishbone_bd_ram_mem1_reg[158][13]/P0001 ,
		_w12898_,
		_w29443_
	);
	LUT2 #(
		.INIT('h8)
	) name18932 (
		\wishbone_bd_ram_mem1_reg[77][13]/P0001 ,
		_w12982_,
		_w29444_
	);
	LUT2 #(
		.INIT('h8)
	) name18933 (
		\wishbone_bd_ram_mem1_reg[239][13]/P0001 ,
		_w12862_,
		_w29445_
	);
	LUT2 #(
		.INIT('h8)
	) name18934 (
		\wishbone_bd_ram_mem1_reg[42][13]/P0001 ,
		_w12842_,
		_w29446_
	);
	LUT2 #(
		.INIT('h8)
	) name18935 (
		\wishbone_bd_ram_mem1_reg[155][13]/P0001 ,
		_w13122_,
		_w29447_
	);
	LUT2 #(
		.INIT('h8)
	) name18936 (
		\wishbone_bd_ram_mem1_reg[24][13]/P0001 ,
		_w13084_,
		_w29448_
	);
	LUT2 #(
		.INIT('h8)
	) name18937 (
		\wishbone_bd_ram_mem1_reg[138][13]/P0001 ,
		_w12958_,
		_w29449_
	);
	LUT2 #(
		.INIT('h8)
	) name18938 (
		\wishbone_bd_ram_mem1_reg[40][13]/P0001 ,
		_w13132_,
		_w29450_
	);
	LUT2 #(
		.INIT('h8)
	) name18939 (
		\wishbone_bd_ram_mem1_reg[31][13]/P0001 ,
		_w13198_,
		_w29451_
	);
	LUT2 #(
		.INIT('h8)
	) name18940 (
		\wishbone_bd_ram_mem1_reg[102][13]/P0001 ,
		_w12685_,
		_w29452_
	);
	LUT2 #(
		.INIT('h8)
	) name18941 (
		\wishbone_bd_ram_mem1_reg[75][13]/P0001 ,
		_w12826_,
		_w29453_
	);
	LUT2 #(
		.INIT('h8)
	) name18942 (
		\wishbone_bd_ram_mem1_reg[8][13]/P0001 ,
		_w12920_,
		_w29454_
	);
	LUT2 #(
		.INIT('h8)
	) name18943 (
		\wishbone_bd_ram_mem1_reg[21][13]/P0001 ,
		_w12906_,
		_w29455_
	);
	LUT2 #(
		.INIT('h8)
	) name18944 (
		\wishbone_bd_ram_mem1_reg[18][13]/P0001 ,
		_w12679_,
		_w29456_
	);
	LUT2 #(
		.INIT('h8)
	) name18945 (
		\wishbone_bd_ram_mem1_reg[76][13]/P0001 ,
		_w13184_,
		_w29457_
	);
	LUT2 #(
		.INIT('h8)
	) name18946 (
		\wishbone_bd_ram_mem1_reg[224][13]/P0001 ,
		_w12902_,
		_w29458_
	);
	LUT2 #(
		.INIT('h8)
	) name18947 (
		\wishbone_bd_ram_mem1_reg[27][13]/P0001 ,
		_w12880_,
		_w29459_
	);
	LUT2 #(
		.INIT('h8)
	) name18948 (
		\wishbone_bd_ram_mem1_reg[208][13]/P0001 ,
		_w13032_,
		_w29460_
	);
	LUT2 #(
		.INIT('h8)
	) name18949 (
		\wishbone_bd_ram_mem1_reg[79][13]/P0001 ,
		_w13212_,
		_w29461_
	);
	LUT2 #(
		.INIT('h8)
	) name18950 (
		\wishbone_bd_ram_mem1_reg[60][13]/P0001 ,
		_w13204_,
		_w29462_
	);
	LUT2 #(
		.INIT('h8)
	) name18951 (
		\wishbone_bd_ram_mem1_reg[214][13]/P0001 ,
		_w12984_,
		_w29463_
	);
	LUT2 #(
		.INIT('h8)
	) name18952 (
		\wishbone_bd_ram_mem1_reg[45][13]/P0001 ,
		_w12908_,
		_w29464_
	);
	LUT2 #(
		.INIT('h8)
	) name18953 (
		\wishbone_bd_ram_mem1_reg[110][13]/P0001 ,
		_w13046_,
		_w29465_
	);
	LUT2 #(
		.INIT('h8)
	) name18954 (
		\wishbone_bd_ram_mem1_reg[66][13]/P0001 ,
		_w12824_,
		_w29466_
	);
	LUT2 #(
		.INIT('h8)
	) name18955 (
		\wishbone_bd_ram_mem1_reg[170][13]/P0001 ,
		_w13030_,
		_w29467_
	);
	LUT2 #(
		.INIT('h8)
	) name18956 (
		\wishbone_bd_ram_mem1_reg[133][13]/P0001 ,
		_w12761_,
		_w29468_
	);
	LUT2 #(
		.INIT('h8)
	) name18957 (
		\wishbone_bd_ram_mem1_reg[111][13]/P0001 ,
		_w12744_,
		_w29469_
	);
	LUT2 #(
		.INIT('h8)
	) name18958 (
		\wishbone_bd_ram_mem1_reg[206][13]/P0001 ,
		_w12954_,
		_w29470_
	);
	LUT2 #(
		.INIT('h8)
	) name18959 (
		\wishbone_bd_ram_mem1_reg[112][13]/P0001 ,
		_w12733_,
		_w29471_
	);
	LUT2 #(
		.INIT('h8)
	) name18960 (
		\wishbone_bd_ram_mem1_reg[160][13]/P0001 ,
		_w12872_,
		_w29472_
	);
	LUT2 #(
		.INIT('h8)
	) name18961 (
		\wishbone_bd_ram_mem1_reg[167][13]/P0001 ,
		_w12986_,
		_w29473_
	);
	LUT2 #(
		.INIT('h8)
	) name18962 (
		\wishbone_bd_ram_mem1_reg[250][13]/P0001 ,
		_w13128_,
		_w29474_
	);
	LUT2 #(
		.INIT('h8)
	) name18963 (
		\wishbone_bd_ram_mem1_reg[240][13]/P0001 ,
		_w12864_,
		_w29475_
	);
	LUT2 #(
		.INIT('h8)
	) name18964 (
		\wishbone_bd_ram_mem1_reg[220][13]/P0001 ,
		_w13066_,
		_w29476_
	);
	LUT2 #(
		.INIT('h8)
	) name18965 (
		\wishbone_bd_ram_mem1_reg[251][13]/P0001 ,
		_w13054_,
		_w29477_
	);
	LUT2 #(
		.INIT('h8)
	) name18966 (
		\wishbone_bd_ram_mem1_reg[148][13]/P0001 ,
		_w13000_,
		_w29478_
	);
	LUT2 #(
		.INIT('h8)
	) name18967 (
		\wishbone_bd_ram_mem1_reg[108][13]/P0001 ,
		_w13156_,
		_w29479_
	);
	LUT2 #(
		.INIT('h8)
	) name18968 (
		\wishbone_bd_ram_mem1_reg[200][13]/P0001 ,
		_w12988_,
		_w29480_
	);
	LUT2 #(
		.INIT('h8)
	) name18969 (
		\wishbone_bd_ram_mem1_reg[91][13]/P0001 ,
		_w13074_,
		_w29481_
	);
	LUT2 #(
		.INIT('h8)
	) name18970 (
		\wishbone_bd_ram_mem1_reg[101][13]/P0001 ,
		_w13192_,
		_w29482_
	);
	LUT2 #(
		.INIT('h8)
	) name18971 (
		\wishbone_bd_ram_mem1_reg[132][13]/P0001 ,
		_w12992_,
		_w29483_
	);
	LUT2 #(
		.INIT('h8)
	) name18972 (
		\wishbone_bd_ram_mem1_reg[88][13]/P0001 ,
		_w12860_,
		_w29484_
	);
	LUT2 #(
		.INIT('h8)
	) name18973 (
		\wishbone_bd_ram_mem1_reg[109][13]/P0001 ,
		_w12888_,
		_w29485_
	);
	LUT2 #(
		.INIT('h8)
	) name18974 (
		\wishbone_bd_ram_mem1_reg[50][13]/P0001 ,
		_w13150_,
		_w29486_
	);
	LUT2 #(
		.INIT('h8)
	) name18975 (
		\wishbone_bd_ram_mem1_reg[118][13]/P0001 ,
		_w12830_,
		_w29487_
	);
	LUT2 #(
		.INIT('h8)
	) name18976 (
		\wishbone_bd_ram_mem1_reg[178][13]/P0001 ,
		_w12886_,
		_w29488_
	);
	LUT2 #(
		.INIT('h8)
	) name18977 (
		\wishbone_bd_ram_mem1_reg[92][13]/P0001 ,
		_w13010_,
		_w29489_
	);
	LUT2 #(
		.INIT('h8)
	) name18978 (
		\wishbone_bd_ram_mem1_reg[69][13]/P0001 ,
		_w12738_,
		_w29490_
	);
	LUT2 #(
		.INIT('h8)
	) name18979 (
		\wishbone_bd_ram_mem1_reg[191][13]/P0001 ,
		_w13034_,
		_w29491_
	);
	LUT2 #(
		.INIT('h8)
	) name18980 (
		\wishbone_bd_ram_mem1_reg[120][13]/P0001 ,
		_w12707_,
		_w29492_
	);
	LUT2 #(
		.INIT('h8)
	) name18981 (
		\wishbone_bd_ram_mem1_reg[237][13]/P0001 ,
		_w12990_,
		_w29493_
	);
	LUT2 #(
		.INIT('h8)
	) name18982 (
		\wishbone_bd_ram_mem1_reg[116][13]/P0001 ,
		_w12998_,
		_w29494_
	);
	LUT2 #(
		.INIT('h8)
	) name18983 (
		\wishbone_bd_ram_mem1_reg[122][13]/P0001 ,
		_w13130_,
		_w29495_
	);
	LUT2 #(
		.INIT('h8)
	) name18984 (
		\wishbone_bd_ram_mem1_reg[7][13]/P0001 ,
		_w12728_,
		_w29496_
	);
	LUT2 #(
		.INIT('h8)
	) name18985 (
		\wishbone_bd_ram_mem1_reg[12][13]/P0001 ,
		_w13118_,
		_w29497_
	);
	LUT2 #(
		.INIT('h8)
	) name18986 (
		\wishbone_bd_ram_mem1_reg[169][13]/P0001 ,
		_w12722_,
		_w29498_
	);
	LUT2 #(
		.INIT('h8)
	) name18987 (
		\wishbone_bd_ram_mem1_reg[49][13]/P0001 ,
		_w12994_,
		_w29499_
	);
	LUT2 #(
		.INIT('h8)
	) name18988 (
		\wishbone_bd_ram_mem1_reg[184][13]/P0001 ,
		_w13062_,
		_w29500_
	);
	LUT2 #(
		.INIT('h8)
	) name18989 (
		\wishbone_bd_ram_mem1_reg[47][13]/P0001 ,
		_w12904_,
		_w29501_
	);
	LUT2 #(
		.INIT('h8)
	) name18990 (
		\wishbone_bd_ram_mem1_reg[74][13]/P0001 ,
		_w12812_,
		_w29502_
	);
	LUT2 #(
		.INIT('h8)
	) name18991 (
		\wishbone_bd_ram_mem1_reg[84][13]/P0001 ,
		_w12934_,
		_w29503_
	);
	LUT2 #(
		.INIT('h8)
	) name18992 (
		\wishbone_bd_ram_mem1_reg[90][13]/P0001 ,
		_w12978_,
		_w29504_
	);
	LUT2 #(
		.INIT('h8)
	) name18993 (
		\wishbone_bd_ram_mem1_reg[255][13]/P0001 ,
		_w13072_,
		_w29505_
	);
	LUT2 #(
		.INIT('h8)
	) name18994 (
		\wishbone_bd_ram_mem1_reg[177][13]/P0001 ,
		_w12996_,
		_w29506_
	);
	LUT2 #(
		.INIT('h8)
	) name18995 (
		\wishbone_bd_ram_mem1_reg[213][13]/P0001 ,
		_w13002_,
		_w29507_
	);
	LUT2 #(
		.INIT('h8)
	) name18996 (
		\wishbone_bd_ram_mem1_reg[13][13]/P0001 ,
		_w13178_,
		_w29508_
	);
	LUT2 #(
		.INIT('h8)
	) name18997 (
		\wishbone_bd_ram_mem1_reg[143][13]/P0001 ,
		_w12922_,
		_w29509_
	);
	LUT2 #(
		.INIT('h8)
	) name18998 (
		\wishbone_bd_ram_mem1_reg[5][13]/P0001 ,
		_w12878_,
		_w29510_
	);
	LUT2 #(
		.INIT('h8)
	) name18999 (
		\wishbone_bd_ram_mem1_reg[217][13]/P0001 ,
		_w13188_,
		_w29511_
	);
	LUT2 #(
		.INIT('h8)
	) name19000 (
		\wishbone_bd_ram_mem1_reg[30][13]/P0001 ,
		_w13104_,
		_w29512_
	);
	LUT2 #(
		.INIT('h8)
	) name19001 (
		\wishbone_bd_ram_mem1_reg[54][13]/P0001 ,
		_w12770_,
		_w29513_
	);
	LUT2 #(
		.INIT('h8)
	) name19002 (
		\wishbone_bd_ram_mem1_reg[176][13]/P0001 ,
		_w12868_,
		_w29514_
	);
	LUT2 #(
		.INIT('h8)
	) name19003 (
		\wishbone_bd_ram_mem1_reg[175][13]/P0001 ,
		_w13126_,
		_w29515_
	);
	LUT2 #(
		.INIT('h8)
	) name19004 (
		\wishbone_bd_ram_mem1_reg[188][13]/P0001 ,
		_w12948_,
		_w29516_
	);
	LUT2 #(
		.INIT('h8)
	) name19005 (
		\wishbone_bd_ram_mem1_reg[134][13]/P0001 ,
		_w12763_,
		_w29517_
	);
	LUT2 #(
		.INIT('h8)
	) name19006 (
		\wishbone_bd_ram_mem1_reg[37][13]/P0001 ,
		_w13102_,
		_w29518_
	);
	LUT2 #(
		.INIT('h8)
	) name19007 (
		\wishbone_bd_ram_mem1_reg[203][13]/P0001 ,
		_w13158_,
		_w29519_
	);
	LUT2 #(
		.INIT('h8)
	) name19008 (
		\wishbone_bd_ram_mem1_reg[65][13]/P0001 ,
		_w13176_,
		_w29520_
	);
	LUT2 #(
		.INIT('h8)
	) name19009 (
		\wishbone_bd_ram_mem1_reg[126][13]/P0001 ,
		_w13218_,
		_w29521_
	);
	LUT2 #(
		.INIT('h8)
	) name19010 (
		\wishbone_bd_ram_mem1_reg[57][13]/P0001 ,
		_w13116_,
		_w29522_
	);
	LUT2 #(
		.INIT('h8)
	) name19011 (
		\wishbone_bd_ram_mem1_reg[82][13]/P0001 ,
		_w12942_,
		_w29523_
	);
	LUT2 #(
		.INIT('h8)
	) name19012 (
		\wishbone_bd_ram_mem1_reg[154][13]/P0001 ,
		_w12962_,
		_w29524_
	);
	LUT2 #(
		.INIT('h8)
	) name19013 (
		\wishbone_bd_ram_mem1_reg[233][13]/P0001 ,
		_w12836_,
		_w29525_
	);
	LUT2 #(
		.INIT('h8)
	) name19014 (
		\wishbone_bd_ram_mem1_reg[87][13]/P0001 ,
		_w13154_,
		_w29526_
	);
	LUT2 #(
		.INIT('h8)
	) name19015 (
		\wishbone_bd_ram_mem1_reg[179][13]/P0001 ,
		_w13050_,
		_w29527_
	);
	LUT2 #(
		.INIT('h8)
	) name19016 (
		\wishbone_bd_ram_mem1_reg[201][13]/P0001 ,
		_w12822_,
		_w29528_
	);
	LUT2 #(
		.INIT('h8)
	) name19017 (
		\wishbone_bd_ram_mem1_reg[209][13]/P0001 ,
		_w13152_,
		_w29529_
	);
	LUT2 #(
		.INIT('h8)
	) name19018 (
		\wishbone_bd_ram_mem1_reg[29][13]/P0001 ,
		_w12952_,
		_w29530_
	);
	LUT2 #(
		.INIT('h8)
	) name19019 (
		\wishbone_bd_ram_mem1_reg[36][13]/P0001 ,
		_w12800_,
		_w29531_
	);
	LUT2 #(
		.INIT('h8)
	) name19020 (
		\wishbone_bd_ram_mem1_reg[97][13]/P0001 ,
		_w13096_,
		_w29532_
	);
	LUT2 #(
		.INIT('h8)
	) name19021 (
		\wishbone_bd_ram_mem1_reg[95][13]/P0001 ,
		_w12844_,
		_w29533_
	);
	LUT2 #(
		.INIT('h8)
	) name19022 (
		\wishbone_bd_ram_mem1_reg[130][13]/P0001 ,
		_w12914_,
		_w29534_
	);
	LUT2 #(
		.INIT('h8)
	) name19023 (
		\wishbone_bd_ram_mem1_reg[107][13]/P0001 ,
		_w12749_,
		_w29535_
	);
	LUT2 #(
		.INIT('h8)
	) name19024 (
		\wishbone_bd_ram_mem1_reg[232][13]/P0001 ,
		_w12758_,
		_w29536_
	);
	LUT2 #(
		.INIT('h8)
	) name19025 (
		\wishbone_bd_ram_mem1_reg[56][13]/P0001 ,
		_w12778_,
		_w29537_
	);
	LUT2 #(
		.INIT('h8)
	) name19026 (
		\wishbone_bd_ram_mem1_reg[171][13]/P0001 ,
		_w12910_,
		_w29538_
	);
	LUT2 #(
		.INIT('h8)
	) name19027 (
		\wishbone_bd_ram_mem1_reg[38][13]/P0001 ,
		_w13182_,
		_w29539_
	);
	LUT2 #(
		.INIT('h8)
	) name19028 (
		\wishbone_bd_ram_mem1_reg[136][13]/P0001 ,
		_w13064_,
		_w29540_
	);
	LUT2 #(
		.INIT('h8)
	) name19029 (
		\wishbone_bd_ram_mem1_reg[6][13]/P0001 ,
		_w12968_,
		_w29541_
	);
	LUT2 #(
		.INIT('h8)
	) name19030 (
		\wishbone_bd_ram_mem1_reg[180][13]/P0001 ,
		_w12791_,
		_w29542_
	);
	LUT2 #(
		.INIT('h8)
	) name19031 (
		\wishbone_bd_ram_mem1_reg[166][13]/P0001 ,
		_w13040_,
		_w29543_
	);
	LUT2 #(
		.INIT('h8)
	) name19032 (
		\wishbone_bd_ram_mem1_reg[152][13]/P0001 ,
		_w12966_,
		_w29544_
	);
	LUT2 #(
		.INIT('h8)
	) name19033 (
		\wishbone_bd_ram_mem1_reg[145][13]/P0001 ,
		_w13106_,
		_w29545_
	);
	LUT2 #(
		.INIT('h8)
	) name19034 (
		\wishbone_bd_ram_mem1_reg[218][13]/P0001 ,
		_w13206_,
		_w29546_
	);
	LUT2 #(
		.INIT('h8)
	) name19035 (
		\wishbone_bd_ram_mem1_reg[141][13]/P0001 ,
		_w13004_,
		_w29547_
	);
	LUT2 #(
		.INIT('h8)
	) name19036 (
		\wishbone_bd_ram_mem1_reg[182][13]/P0001 ,
		_w12820_,
		_w29548_
	);
	LUT2 #(
		.INIT('h8)
	) name19037 (
		\wishbone_bd_ram_mem1_reg[199][13]/P0001 ,
		_w12768_,
		_w29549_
	);
	LUT2 #(
		.INIT('h8)
	) name19038 (
		\wishbone_bd_ram_mem1_reg[216][13]/P0001 ,
		_w13028_,
		_w29550_
	);
	LUT2 #(
		.INIT('h8)
	) name19039 (
		\wishbone_bd_ram_mem1_reg[146][13]/P0001 ,
		_w13060_,
		_w29551_
	);
	LUT2 #(
		.INIT('h8)
	) name19040 (
		\wishbone_bd_ram_mem1_reg[78][13]/P0001 ,
		_w12874_,
		_w29552_
	);
	LUT2 #(
		.INIT('h8)
	) name19041 (
		\wishbone_bd_ram_mem1_reg[137][13]/P0001 ,
		_w13168_,
		_w29553_
	);
	LUT2 #(
		.INIT('h8)
	) name19042 (
		\wishbone_bd_ram_mem1_reg[115][13]/P0001 ,
		_w13112_,
		_w29554_
	);
	LUT2 #(
		.INIT('h8)
	) name19043 (
		\wishbone_bd_ram_mem1_reg[80][13]/P0001 ,
		_w12689_,
		_w29555_
	);
	LUT2 #(
		.INIT('h8)
	) name19044 (
		\wishbone_bd_ram_mem1_reg[100][13]/P0001 ,
		_w12960_,
		_w29556_
	);
	LUT2 #(
		.INIT('h8)
	) name19045 (
		\wishbone_bd_ram_mem1_reg[229][13]/P0001 ,
		_w12711_,
		_w29557_
	);
	LUT2 #(
		.INIT('h8)
	) name19046 (
		\wishbone_bd_ram_mem1_reg[96][13]/P0001 ,
		_w12912_,
		_w29558_
	);
	LUT2 #(
		.INIT('h8)
	) name19047 (
		\wishbone_bd_ram_mem1_reg[252][13]/P0001 ,
		_w13080_,
		_w29559_
	);
	LUT2 #(
		.INIT('h8)
	) name19048 (
		\wishbone_bd_ram_mem1_reg[44][13]/P0001 ,
		_w12896_,
		_w29560_
	);
	LUT2 #(
		.INIT('h8)
	) name19049 (
		\wishbone_bd_ram_mem1_reg[219][13]/P0001 ,
		_w12806_,
		_w29561_
	);
	LUT2 #(
		.INIT('h8)
	) name19050 (
		\wishbone_bd_ram_mem1_reg[150][13]/P0001 ,
		_w13136_,
		_w29562_
	);
	LUT2 #(
		.INIT('h8)
	) name19051 (
		\wishbone_bd_ram_mem1_reg[194][13]/P0001 ,
		_w12772_,
		_w29563_
	);
	LUT2 #(
		.INIT('h8)
	) name19052 (
		\wishbone_bd_ram_mem1_reg[151][13]/P0001 ,
		_w13142_,
		_w29564_
	);
	LUT2 #(
		.INIT('h8)
	) name19053 (
		\wishbone_bd_ram_mem1_reg[11][13]/P0001 ,
		_w13194_,
		_w29565_
	);
	LUT2 #(
		.INIT('h8)
	) name19054 (
		\wishbone_bd_ram_mem1_reg[28][13]/P0001 ,
		_w13170_,
		_w29566_
	);
	LUT2 #(
		.INIT('h8)
	) name19055 (
		\wishbone_bd_ram_mem1_reg[226][13]/P0001 ,
		_w13138_,
		_w29567_
	);
	LUT2 #(
		.INIT('h8)
	) name19056 (
		\wishbone_bd_ram_mem1_reg[144][13]/P0001 ,
		_w12756_,
		_w29568_
	);
	LUT2 #(
		.INIT('h8)
	) name19057 (
		\wishbone_bd_ram_mem1_reg[25][13]/P0001 ,
		_w13108_,
		_w29569_
	);
	LUT2 #(
		.INIT('h8)
	) name19058 (
		\wishbone_bd_ram_mem1_reg[89][13]/P0001 ,
		_w12964_,
		_w29570_
	);
	LUT2 #(
		.INIT('h8)
	) name19059 (
		\wishbone_bd_ram_mem1_reg[192][13]/P0001 ,
		_w12938_,
		_w29571_
	);
	LUT2 #(
		.INIT('h8)
	) name19060 (
		\wishbone_bd_ram_mem1_reg[128][13]/P0001 ,
		_w12793_,
		_w29572_
	);
	LUT2 #(
		.INIT('h8)
	) name19061 (
		\wishbone_bd_ram_mem1_reg[236][13]/P0001 ,
		_w12731_,
		_w29573_
	);
	LUT2 #(
		.INIT('h8)
	) name19062 (
		\wishbone_bd_ram_mem1_reg[198][13]/P0001 ,
		_w12832_,
		_w29574_
	);
	LUT2 #(
		.INIT('h8)
	) name19063 (
		\wishbone_bd_ram_mem1_reg[147][13]/P0001 ,
		_w13146_,
		_w29575_
	);
	LUT2 #(
		.INIT('h8)
	) name19064 (
		\wishbone_bd_ram_mem1_reg[183][13]/P0001 ,
		_w12787_,
		_w29576_
	);
	LUT2 #(
		.INIT('h8)
	) name19065 (
		\wishbone_bd_ram_mem1_reg[15][13]/P0001 ,
		_w13210_,
		_w29577_
	);
	LUT2 #(
		.INIT('h8)
	) name19066 (
		\wishbone_bd_ram_mem1_reg[32][13]/P0001 ,
		_w13120_,
		_w29578_
	);
	LUT2 #(
		.INIT('h8)
	) name19067 (
		\wishbone_bd_ram_mem1_reg[16][13]/P0001 ,
		_w13140_,
		_w29579_
	);
	LUT2 #(
		.INIT('h8)
	) name19068 (
		\wishbone_bd_ram_mem1_reg[33][13]/P0001 ,
		_w12980_,
		_w29580_
	);
	LUT2 #(
		.INIT('h8)
	) name19069 (
		\wishbone_bd_ram_mem1_reg[162][13]/P0001 ,
		_w13098_,
		_w29581_
	);
	LUT2 #(
		.INIT('h8)
	) name19070 (
		\wishbone_bd_ram_mem1_reg[2][13]/P0001 ,
		_w13088_,
		_w29582_
	);
	LUT2 #(
		.INIT('h8)
	) name19071 (
		\wishbone_bd_ram_mem1_reg[238][13]/P0001 ,
		_w13160_,
		_w29583_
	);
	LUT2 #(
		.INIT('h8)
	) name19072 (
		\wishbone_bd_ram_mem1_reg[157][13]/P0001 ,
		_w12926_,
		_w29584_
	);
	LUT2 #(
		.INIT('h8)
	) name19073 (
		\wishbone_bd_ram_mem1_reg[186][13]/P0001 ,
		_w12783_,
		_w29585_
	);
	LUT2 #(
		.INIT('h8)
	) name19074 (
		\wishbone_bd_ram_mem1_reg[105][13]/P0001 ,
		_w12751_,
		_w29586_
	);
	LUT2 #(
		.INIT('h8)
	) name19075 (
		\wishbone_bd_ram_mem1_reg[245][13]/P0001 ,
		_w13022_,
		_w29587_
	);
	LUT2 #(
		.INIT('h8)
	) name19076 (
		\wishbone_bd_ram_mem1_reg[181][13]/P0001 ,
		_w12828_,
		_w29588_
	);
	LUT2 #(
		.INIT('h8)
	) name19077 (
		\wishbone_bd_ram_mem1_reg[9][13]/P0001 ,
		_w12808_,
		_w29589_
	);
	LUT2 #(
		.INIT('h8)
	) name19078 (
		\wishbone_bd_ram_mem1_reg[14][13]/P0001 ,
		_w13086_,
		_w29590_
	);
	LUT2 #(
		.INIT('h8)
	) name19079 (
		\wishbone_bd_ram_mem1_reg[212][13]/P0001 ,
		_w12796_,
		_w29591_
	);
	LUT2 #(
		.INIT('h8)
	) name19080 (
		\wishbone_bd_ram_mem1_reg[23][13]/P0001 ,
		_w13008_,
		_w29592_
	);
	LUT2 #(
		.INIT('h8)
	) name19081 (
		\wishbone_bd_ram_mem1_reg[124][13]/P0001 ,
		_w13058_,
		_w29593_
	);
	LUT2 #(
		.INIT('h8)
	) name19082 (
		\wishbone_bd_ram_mem1_reg[123][13]/P0001 ,
		_w13114_,
		_w29594_
	);
	LUT2 #(
		.INIT('h8)
	) name19083 (
		\wishbone_bd_ram_mem1_reg[0][13]/P0001 ,
		_w12717_,
		_w29595_
	);
	LUT2 #(
		.INIT('h8)
	) name19084 (
		\wishbone_bd_ram_mem1_reg[196][13]/P0001 ,
		_w13090_,
		_w29596_
	);
	LUT2 #(
		.INIT('h8)
	) name19085 (
		\wishbone_bd_ram_mem1_reg[189][13]/P0001 ,
		_w13042_,
		_w29597_
	);
	LUT2 #(
		.INIT('h8)
	) name19086 (
		\wishbone_bd_ram_mem1_reg[83][13]/P0001 ,
		_w12916_,
		_w29598_
	);
	LUT2 #(
		.INIT('h8)
	) name19087 (
		\wishbone_bd_ram_mem1_reg[231][13]/P0001 ,
		_w12856_,
		_w29599_
	);
	LUT2 #(
		.INIT('h8)
	) name19088 (
		\wishbone_bd_ram_mem1_reg[173][13]/P0001 ,
		_w12854_,
		_w29600_
	);
	LUT2 #(
		.INIT('h8)
	) name19089 (
		\wishbone_bd_ram_mem1_reg[46][13]/P0001 ,
		_w12884_,
		_w29601_
	);
	LUT2 #(
		.INIT('h8)
	) name19090 (
		\wishbone_bd_ram_mem1_reg[119][13]/P0001 ,
		_w13048_,
		_w29602_
	);
	LUT2 #(
		.INIT('h8)
	) name19091 (
		\wishbone_bd_ram_mem1_reg[43][13]/P0001 ,
		_w13200_,
		_w29603_
	);
	LUT2 #(
		.INIT('h8)
	) name19092 (
		\wishbone_bd_ram_mem1_reg[73][13]/P0001 ,
		_w12918_,
		_w29604_
	);
	LUT2 #(
		.INIT('h8)
	) name19093 (
		\wishbone_bd_ram_mem1_reg[225][13]/P0001 ,
		_w13092_,
		_w29605_
	);
	LUT2 #(
		.INIT('h8)
	) name19094 (
		\wishbone_bd_ram_mem1_reg[106][13]/P0001 ,
		_w12713_,
		_w29606_
	);
	LUT2 #(
		.INIT('h8)
	) name19095 (
		\wishbone_bd_ram_mem1_reg[98][13]/P0001 ,
		_w12816_,
		_w29607_
	);
	LUT2 #(
		.INIT('h8)
	) name19096 (
		\wishbone_bd_ram_mem1_reg[129][13]/P0001 ,
		_w12776_,
		_w29608_
	);
	LUT2 #(
		.INIT('h8)
	) name19097 (
		\wishbone_bd_ram_mem1_reg[254][13]/P0001 ,
		_w12892_,
		_w29609_
	);
	LUT2 #(
		.INIT('h8)
	) name19098 (
		\wishbone_bd_ram_mem1_reg[139][13]/P0001 ,
		_w12814_,
		_w29610_
	);
	LUT2 #(
		.INIT('h8)
	) name19099 (
		\wishbone_bd_ram_mem1_reg[159][13]/P0001 ,
		_w12774_,
		_w29611_
	);
	LUT2 #(
		.INIT('h8)
	) name19100 (
		\wishbone_bd_ram_mem1_reg[244][13]/P0001 ,
		_w12747_,
		_w29612_
	);
	LUT2 #(
		.INIT('h8)
	) name19101 (
		\wishbone_bd_ram_mem1_reg[228][13]/P0001 ,
		_w12765_,
		_w29613_
	);
	LUT2 #(
		.INIT('h8)
	) name19102 (
		\wishbone_bd_ram_mem1_reg[163][13]/P0001 ,
		_w12882_,
		_w29614_
	);
	LUT2 #(
		.INIT('h8)
	) name19103 (
		\wishbone_bd_ram_mem1_reg[121][13]/P0001 ,
		_w13078_,
		_w29615_
	);
	LUT2 #(
		.INIT('h8)
	) name19104 (
		\wishbone_bd_ram_mem1_reg[140][13]/P0001 ,
		_w12894_,
		_w29616_
	);
	LUT2 #(
		.INIT('h8)
	) name19105 (
		\wishbone_bd_ram_mem1_reg[67][13]/P0001 ,
		_w13134_,
		_w29617_
	);
	LUT2 #(
		.INIT('h8)
	) name19106 (
		\wishbone_bd_ram_mem1_reg[185][13]/P0001 ,
		_w12940_,
		_w29618_
	);
	LUT2 #(
		.INIT('h8)
	) name19107 (
		\wishbone_bd_ram_mem1_reg[202][13]/P0001 ,
		_w12870_,
		_w29619_
	);
	LUT2 #(
		.INIT('h8)
	) name19108 (
		\wishbone_bd_ram_mem1_reg[190][13]/P0001 ,
		_w12858_,
		_w29620_
	);
	LUT2 #(
		.INIT('h8)
	) name19109 (
		\wishbone_bd_ram_mem1_reg[4][13]/P0001 ,
		_w12666_,
		_w29621_
	);
	LUT2 #(
		.INIT('h8)
	) name19110 (
		\wishbone_bd_ram_mem1_reg[193][13]/P0001 ,
		_w13056_,
		_w29622_
	);
	LUT2 #(
		.INIT('h8)
	) name19111 (
		\wishbone_bd_ram_mem1_reg[204][13]/P0001 ,
		_w13162_,
		_w29623_
	);
	LUT2 #(
		.INIT('h8)
	) name19112 (
		\wishbone_bd_ram_mem1_reg[243][13]/P0001 ,
		_w12804_,
		_w29624_
	);
	LUT2 #(
		.INIT('h8)
	) name19113 (
		\wishbone_bd_ram_mem1_reg[210][13]/P0001 ,
		_w12924_,
		_w29625_
	);
	LUT2 #(
		.INIT('h8)
	) name19114 (
		\wishbone_bd_ram_mem1_reg[205][13]/P0001 ,
		_w13068_,
		_w29626_
	);
	LUT2 #(
		.INIT('h8)
	) name19115 (
		\wishbone_bd_ram_mem1_reg[48][13]/P0001 ,
		_w12970_,
		_w29627_
	);
	LUT2 #(
		.INIT('h8)
	) name19116 (
		\wishbone_bd_ram_mem1_reg[187][13]/P0001 ,
		_w13196_,
		_w29628_
	);
	LUT2 #(
		.INIT('h8)
	) name19117 (
		\wishbone_bd_ram_mem1_reg[10][13]/P0001 ,
		_w13172_,
		_w29629_
	);
	LUT2 #(
		.INIT('h8)
	) name19118 (
		\wishbone_bd_ram_mem1_reg[94][13]/P0001 ,
		_w13186_,
		_w29630_
	);
	LUT2 #(
		.INIT('h8)
	) name19119 (
		\wishbone_bd_ram_mem1_reg[234][13]/P0001 ,
		_w13214_,
		_w29631_
	);
	LUT2 #(
		.INIT('h8)
	) name19120 (
		\wishbone_bd_ram_mem1_reg[172][13]/P0001 ,
		_w12944_,
		_w29632_
	);
	LUT2 #(
		.INIT('h8)
	) name19121 (
		\wishbone_bd_ram_mem1_reg[26][13]/P0001 ,
		_w12699_,
		_w29633_
	);
	LUT2 #(
		.INIT('h8)
	) name19122 (
		\wishbone_bd_ram_mem1_reg[164][13]/P0001 ,
		_w12876_,
		_w29634_
	);
	LUT2 #(
		.INIT('h8)
	) name19123 (
		\wishbone_bd_ram_mem1_reg[3][13]/P0001 ,
		_w12866_,
		_w29635_
	);
	LUT2 #(
		.INIT('h8)
	) name19124 (
		\wishbone_bd_ram_mem1_reg[195][13]/P0001 ,
		_w13144_,
		_w29636_
	);
	LUT2 #(
		.INIT('h8)
	) name19125 (
		\wishbone_bd_ram_mem1_reg[70][13]/P0001 ,
		_w12840_,
		_w29637_
	);
	LUT2 #(
		.INIT('h8)
	) name19126 (
		\wishbone_bd_ram_mem1_reg[165][13]/P0001 ,
		_w13044_,
		_w29638_
	);
	LUT2 #(
		.INIT('h8)
	) name19127 (
		\wishbone_bd_ram_mem1_reg[71][13]/P0001 ,
		_w12798_,
		_w29639_
	);
	LUT2 #(
		.INIT('h8)
	) name19128 (
		\wishbone_bd_ram_mem1_reg[39][13]/P0001 ,
		_w13018_,
		_w29640_
	);
	LUT2 #(
		.INIT('h8)
	) name19129 (
		\wishbone_bd_ram_mem1_reg[113][13]/P0001 ,
		_w13026_,
		_w29641_
	);
	LUT2 #(
		.INIT('h8)
	) name19130 (
		\wishbone_bd_ram_mem1_reg[168][13]/P0001 ,
		_w13208_,
		_w29642_
	);
	LUT2 #(
		.INIT('h8)
	) name19131 (
		\wishbone_bd_ram_mem1_reg[22][13]/P0001 ,
		_w13110_,
		_w29643_
	);
	LUT2 #(
		.INIT('h8)
	) name19132 (
		\wishbone_bd_ram_mem1_reg[68][13]/P0001 ,
		_w12946_,
		_w29644_
	);
	LUT2 #(
		.INIT('h8)
	) name19133 (
		\wishbone_bd_ram_mem1_reg[17][13]/P0001 ,
		_w12848_,
		_w29645_
	);
	LUT2 #(
		.INIT('h8)
	) name19134 (
		\wishbone_bd_ram_mem1_reg[249][13]/P0001 ,
		_w12900_,
		_w29646_
	);
	LUT2 #(
		.INIT('h8)
	) name19135 (
		\wishbone_bd_ram_mem1_reg[19][13]/P0001 ,
		_w13012_,
		_w29647_
	);
	LUT2 #(
		.INIT('h8)
	) name19136 (
		\wishbone_bd_ram_mem1_reg[153][13]/P0001 ,
		_w12890_,
		_w29648_
	);
	LUT2 #(
		.INIT('h8)
	) name19137 (
		\wishbone_bd_ram_mem1_reg[127][13]/P0001 ,
		_w13164_,
		_w29649_
	);
	LUT2 #(
		.INIT('h8)
	) name19138 (
		\wishbone_bd_ram_mem1_reg[55][13]/P0001 ,
		_w12785_,
		_w29650_
	);
	LUT2 #(
		.INIT('h8)
	) name19139 (
		\wishbone_bd_ram_mem1_reg[53][13]/P0001 ,
		_w13020_,
		_w29651_
	);
	LUT2 #(
		.INIT('h8)
	) name19140 (
		\wishbone_bd_ram_mem1_reg[104][13]/P0001 ,
		_w13148_,
		_w29652_
	);
	LUT2 #(
		.INIT('h8)
	) name19141 (
		\wishbone_bd_ram_mem1_reg[62][13]/P0001 ,
		_w12673_,
		_w29653_
	);
	LUT2 #(
		.INIT('h8)
	) name19142 (
		\wishbone_bd_ram_mem1_reg[41][13]/P0001 ,
		_w13052_,
		_w29654_
	);
	LUT2 #(
		.INIT('h8)
	) name19143 (
		\wishbone_bd_ram_mem1_reg[117][13]/P0001 ,
		_w12715_,
		_w29655_
	);
	LUT2 #(
		.INIT('h8)
	) name19144 (
		\wishbone_bd_ram_mem1_reg[161][13]/P0001 ,
		_w12754_,
		_w29656_
	);
	LUT2 #(
		.INIT('h8)
	) name19145 (
		\wishbone_bd_ram_mem1_reg[20][13]/P0001 ,
		_w13174_,
		_w29657_
	);
	LUT2 #(
		.INIT('h8)
	) name19146 (
		\wishbone_bd_ram_mem1_reg[86][13]/P0001 ,
		_w12735_,
		_w29658_
	);
	LUT2 #(
		.INIT('h8)
	) name19147 (
		\wishbone_bd_ram_mem1_reg[227][13]/P0001 ,
		_w12936_,
		_w29659_
	);
	LUT2 #(
		.INIT('h8)
	) name19148 (
		\wishbone_bd_ram_mem1_reg[72][13]/P0001 ,
		_w12810_,
		_w29660_
	);
	LUT2 #(
		.INIT('h8)
	) name19149 (
		\wishbone_bd_ram_mem1_reg[223][13]/P0001 ,
		_w12838_,
		_w29661_
	);
	LUT2 #(
		.INIT('h8)
	) name19150 (
		\wishbone_bd_ram_mem1_reg[207][13]/P0001 ,
		_w13180_,
		_w29662_
	);
	LUT2 #(
		.INIT('h8)
	) name19151 (
		\wishbone_bd_ram_mem1_reg[242][13]/P0001 ,
		_w12932_,
		_w29663_
	);
	LUT2 #(
		.INIT('h8)
	) name19152 (
		\wishbone_bd_ram_mem1_reg[211][13]/P0001 ,
		_w13166_,
		_w29664_
	);
	LUT2 #(
		.INIT('h8)
	) name19153 (
		\wishbone_bd_ram_mem1_reg[156][13]/P0001 ,
		_w13190_,
		_w29665_
	);
	LUT2 #(
		.INIT('h8)
	) name19154 (
		\wishbone_bd_ram_mem1_reg[142][13]/P0001 ,
		_w12928_,
		_w29666_
	);
	LUT2 #(
		.INIT('h8)
	) name19155 (
		\wishbone_bd_ram_mem1_reg[51][13]/P0001 ,
		_w13024_,
		_w29667_
	);
	LUT2 #(
		.INIT('h8)
	) name19156 (
		\wishbone_bd_ram_mem1_reg[215][13]/P0001 ,
		_w12974_,
		_w29668_
	);
	LUT2 #(
		.INIT('h8)
	) name19157 (
		\wishbone_bd_ram_mem1_reg[64][13]/P0001 ,
		_w12976_,
		_w29669_
	);
	LUT2 #(
		.INIT('h8)
	) name19158 (
		\wishbone_bd_ram_mem1_reg[1][13]/P0001 ,
		_w13014_,
		_w29670_
	);
	LUT2 #(
		.INIT('h8)
	) name19159 (
		\wishbone_bd_ram_mem1_reg[58][13]/P0001 ,
		_w13070_,
		_w29671_
	);
	LUT2 #(
		.INIT('h8)
	) name19160 (
		\wishbone_bd_ram_mem1_reg[221][13]/P0001 ,
		_w12802_,
		_w29672_
	);
	LUT2 #(
		.INIT('h8)
	) name19161 (
		\wishbone_bd_ram_mem1_reg[230][13]/P0001 ,
		_w13036_,
		_w29673_
	);
	LUT2 #(
		.INIT('h8)
	) name19162 (
		\wishbone_bd_ram_mem1_reg[35][13]/P0001 ,
		_w12703_,
		_w29674_
	);
	LUT2 #(
		.INIT('h8)
	) name19163 (
		\wishbone_bd_ram_mem1_reg[241][13]/P0001 ,
		_w13006_,
		_w29675_
	);
	LUT2 #(
		.INIT('h8)
	) name19164 (
		\wishbone_bd_ram_mem1_reg[93][13]/P0001 ,
		_w13016_,
		_w29676_
	);
	LUT2 #(
		.INIT('h8)
	) name19165 (
		\wishbone_bd_ram_mem1_reg[125][13]/P0001 ,
		_w12956_,
		_w29677_
	);
	LUT2 #(
		.INIT('h8)
	) name19166 (
		\wishbone_bd_ram_mem1_reg[63][13]/P0001 ,
		_w12850_,
		_w29678_
	);
	LUT2 #(
		.INIT('h8)
	) name19167 (
		\wishbone_bd_ram_mem1_reg[246][13]/P0001 ,
		_w13076_,
		_w29679_
	);
	LUT2 #(
		.INIT('h8)
	) name19168 (
		\wishbone_bd_ram_mem1_reg[81][13]/P0001 ,
		_w12950_,
		_w29680_
	);
	LUT2 #(
		.INIT('h8)
	) name19169 (
		\wishbone_bd_ram_mem1_reg[253][13]/P0001 ,
		_w13100_,
		_w29681_
	);
	LUT2 #(
		.INIT('h8)
	) name19170 (
		\wishbone_bd_ram_mem1_reg[197][13]/P0001 ,
		_w12834_,
		_w29682_
	);
	LUT2 #(
		.INIT('h8)
	) name19171 (
		\wishbone_bd_ram_mem1_reg[174][13]/P0001 ,
		_w12972_,
		_w29683_
	);
	LUT2 #(
		.INIT('h8)
	) name19172 (
		\wishbone_bd_ram_mem1_reg[149][13]/P0001 ,
		_w12741_,
		_w29684_
	);
	LUT2 #(
		.INIT('h8)
	) name19173 (
		\wishbone_bd_ram_mem1_reg[222][13]/P0001 ,
		_w13094_,
		_w29685_
	);
	LUT2 #(
		.INIT('h8)
	) name19174 (
		\wishbone_bd_ram_mem1_reg[99][13]/P0001 ,
		_w13038_,
		_w29686_
	);
	LUT2 #(
		.INIT('h8)
	) name19175 (
		\wishbone_bd_ram_mem1_reg[248][13]/P0001 ,
		_w12789_,
		_w29687_
	);
	LUT2 #(
		.INIT('h8)
	) name19176 (
		\wishbone_bd_ram_mem1_reg[135][13]/P0001 ,
		_w13124_,
		_w29688_
	);
	LUT2 #(
		.INIT('h8)
	) name19177 (
		\wishbone_bd_ram_mem1_reg[59][13]/P0001 ,
		_w12780_,
		_w29689_
	);
	LUT2 #(
		.INIT('h8)
	) name19178 (
		\wishbone_bd_ram_mem1_reg[61][13]/P0001 ,
		_w12725_,
		_w29690_
	);
	LUT2 #(
		.INIT('h8)
	) name19179 (
		\wishbone_bd_ram_mem1_reg[235][13]/P0001 ,
		_w12696_,
		_w29691_
	);
	LUT2 #(
		.INIT('h1)
	) name19180 (
		_w29436_,
		_w29437_,
		_w29692_
	);
	LUT2 #(
		.INIT('h1)
	) name19181 (
		_w29438_,
		_w29439_,
		_w29693_
	);
	LUT2 #(
		.INIT('h1)
	) name19182 (
		_w29440_,
		_w29441_,
		_w29694_
	);
	LUT2 #(
		.INIT('h1)
	) name19183 (
		_w29442_,
		_w29443_,
		_w29695_
	);
	LUT2 #(
		.INIT('h1)
	) name19184 (
		_w29444_,
		_w29445_,
		_w29696_
	);
	LUT2 #(
		.INIT('h1)
	) name19185 (
		_w29446_,
		_w29447_,
		_w29697_
	);
	LUT2 #(
		.INIT('h1)
	) name19186 (
		_w29448_,
		_w29449_,
		_w29698_
	);
	LUT2 #(
		.INIT('h1)
	) name19187 (
		_w29450_,
		_w29451_,
		_w29699_
	);
	LUT2 #(
		.INIT('h1)
	) name19188 (
		_w29452_,
		_w29453_,
		_w29700_
	);
	LUT2 #(
		.INIT('h1)
	) name19189 (
		_w29454_,
		_w29455_,
		_w29701_
	);
	LUT2 #(
		.INIT('h1)
	) name19190 (
		_w29456_,
		_w29457_,
		_w29702_
	);
	LUT2 #(
		.INIT('h1)
	) name19191 (
		_w29458_,
		_w29459_,
		_w29703_
	);
	LUT2 #(
		.INIT('h1)
	) name19192 (
		_w29460_,
		_w29461_,
		_w29704_
	);
	LUT2 #(
		.INIT('h1)
	) name19193 (
		_w29462_,
		_w29463_,
		_w29705_
	);
	LUT2 #(
		.INIT('h1)
	) name19194 (
		_w29464_,
		_w29465_,
		_w29706_
	);
	LUT2 #(
		.INIT('h1)
	) name19195 (
		_w29466_,
		_w29467_,
		_w29707_
	);
	LUT2 #(
		.INIT('h1)
	) name19196 (
		_w29468_,
		_w29469_,
		_w29708_
	);
	LUT2 #(
		.INIT('h1)
	) name19197 (
		_w29470_,
		_w29471_,
		_w29709_
	);
	LUT2 #(
		.INIT('h1)
	) name19198 (
		_w29472_,
		_w29473_,
		_w29710_
	);
	LUT2 #(
		.INIT('h1)
	) name19199 (
		_w29474_,
		_w29475_,
		_w29711_
	);
	LUT2 #(
		.INIT('h1)
	) name19200 (
		_w29476_,
		_w29477_,
		_w29712_
	);
	LUT2 #(
		.INIT('h1)
	) name19201 (
		_w29478_,
		_w29479_,
		_w29713_
	);
	LUT2 #(
		.INIT('h1)
	) name19202 (
		_w29480_,
		_w29481_,
		_w29714_
	);
	LUT2 #(
		.INIT('h1)
	) name19203 (
		_w29482_,
		_w29483_,
		_w29715_
	);
	LUT2 #(
		.INIT('h1)
	) name19204 (
		_w29484_,
		_w29485_,
		_w29716_
	);
	LUT2 #(
		.INIT('h1)
	) name19205 (
		_w29486_,
		_w29487_,
		_w29717_
	);
	LUT2 #(
		.INIT('h1)
	) name19206 (
		_w29488_,
		_w29489_,
		_w29718_
	);
	LUT2 #(
		.INIT('h1)
	) name19207 (
		_w29490_,
		_w29491_,
		_w29719_
	);
	LUT2 #(
		.INIT('h1)
	) name19208 (
		_w29492_,
		_w29493_,
		_w29720_
	);
	LUT2 #(
		.INIT('h1)
	) name19209 (
		_w29494_,
		_w29495_,
		_w29721_
	);
	LUT2 #(
		.INIT('h1)
	) name19210 (
		_w29496_,
		_w29497_,
		_w29722_
	);
	LUT2 #(
		.INIT('h1)
	) name19211 (
		_w29498_,
		_w29499_,
		_w29723_
	);
	LUT2 #(
		.INIT('h1)
	) name19212 (
		_w29500_,
		_w29501_,
		_w29724_
	);
	LUT2 #(
		.INIT('h1)
	) name19213 (
		_w29502_,
		_w29503_,
		_w29725_
	);
	LUT2 #(
		.INIT('h1)
	) name19214 (
		_w29504_,
		_w29505_,
		_w29726_
	);
	LUT2 #(
		.INIT('h1)
	) name19215 (
		_w29506_,
		_w29507_,
		_w29727_
	);
	LUT2 #(
		.INIT('h1)
	) name19216 (
		_w29508_,
		_w29509_,
		_w29728_
	);
	LUT2 #(
		.INIT('h1)
	) name19217 (
		_w29510_,
		_w29511_,
		_w29729_
	);
	LUT2 #(
		.INIT('h1)
	) name19218 (
		_w29512_,
		_w29513_,
		_w29730_
	);
	LUT2 #(
		.INIT('h1)
	) name19219 (
		_w29514_,
		_w29515_,
		_w29731_
	);
	LUT2 #(
		.INIT('h1)
	) name19220 (
		_w29516_,
		_w29517_,
		_w29732_
	);
	LUT2 #(
		.INIT('h1)
	) name19221 (
		_w29518_,
		_w29519_,
		_w29733_
	);
	LUT2 #(
		.INIT('h1)
	) name19222 (
		_w29520_,
		_w29521_,
		_w29734_
	);
	LUT2 #(
		.INIT('h1)
	) name19223 (
		_w29522_,
		_w29523_,
		_w29735_
	);
	LUT2 #(
		.INIT('h1)
	) name19224 (
		_w29524_,
		_w29525_,
		_w29736_
	);
	LUT2 #(
		.INIT('h1)
	) name19225 (
		_w29526_,
		_w29527_,
		_w29737_
	);
	LUT2 #(
		.INIT('h1)
	) name19226 (
		_w29528_,
		_w29529_,
		_w29738_
	);
	LUT2 #(
		.INIT('h1)
	) name19227 (
		_w29530_,
		_w29531_,
		_w29739_
	);
	LUT2 #(
		.INIT('h1)
	) name19228 (
		_w29532_,
		_w29533_,
		_w29740_
	);
	LUT2 #(
		.INIT('h1)
	) name19229 (
		_w29534_,
		_w29535_,
		_w29741_
	);
	LUT2 #(
		.INIT('h1)
	) name19230 (
		_w29536_,
		_w29537_,
		_w29742_
	);
	LUT2 #(
		.INIT('h1)
	) name19231 (
		_w29538_,
		_w29539_,
		_w29743_
	);
	LUT2 #(
		.INIT('h1)
	) name19232 (
		_w29540_,
		_w29541_,
		_w29744_
	);
	LUT2 #(
		.INIT('h1)
	) name19233 (
		_w29542_,
		_w29543_,
		_w29745_
	);
	LUT2 #(
		.INIT('h1)
	) name19234 (
		_w29544_,
		_w29545_,
		_w29746_
	);
	LUT2 #(
		.INIT('h1)
	) name19235 (
		_w29546_,
		_w29547_,
		_w29747_
	);
	LUT2 #(
		.INIT('h1)
	) name19236 (
		_w29548_,
		_w29549_,
		_w29748_
	);
	LUT2 #(
		.INIT('h1)
	) name19237 (
		_w29550_,
		_w29551_,
		_w29749_
	);
	LUT2 #(
		.INIT('h1)
	) name19238 (
		_w29552_,
		_w29553_,
		_w29750_
	);
	LUT2 #(
		.INIT('h1)
	) name19239 (
		_w29554_,
		_w29555_,
		_w29751_
	);
	LUT2 #(
		.INIT('h1)
	) name19240 (
		_w29556_,
		_w29557_,
		_w29752_
	);
	LUT2 #(
		.INIT('h1)
	) name19241 (
		_w29558_,
		_w29559_,
		_w29753_
	);
	LUT2 #(
		.INIT('h1)
	) name19242 (
		_w29560_,
		_w29561_,
		_w29754_
	);
	LUT2 #(
		.INIT('h1)
	) name19243 (
		_w29562_,
		_w29563_,
		_w29755_
	);
	LUT2 #(
		.INIT('h1)
	) name19244 (
		_w29564_,
		_w29565_,
		_w29756_
	);
	LUT2 #(
		.INIT('h1)
	) name19245 (
		_w29566_,
		_w29567_,
		_w29757_
	);
	LUT2 #(
		.INIT('h1)
	) name19246 (
		_w29568_,
		_w29569_,
		_w29758_
	);
	LUT2 #(
		.INIT('h1)
	) name19247 (
		_w29570_,
		_w29571_,
		_w29759_
	);
	LUT2 #(
		.INIT('h1)
	) name19248 (
		_w29572_,
		_w29573_,
		_w29760_
	);
	LUT2 #(
		.INIT('h1)
	) name19249 (
		_w29574_,
		_w29575_,
		_w29761_
	);
	LUT2 #(
		.INIT('h1)
	) name19250 (
		_w29576_,
		_w29577_,
		_w29762_
	);
	LUT2 #(
		.INIT('h1)
	) name19251 (
		_w29578_,
		_w29579_,
		_w29763_
	);
	LUT2 #(
		.INIT('h1)
	) name19252 (
		_w29580_,
		_w29581_,
		_w29764_
	);
	LUT2 #(
		.INIT('h1)
	) name19253 (
		_w29582_,
		_w29583_,
		_w29765_
	);
	LUT2 #(
		.INIT('h1)
	) name19254 (
		_w29584_,
		_w29585_,
		_w29766_
	);
	LUT2 #(
		.INIT('h1)
	) name19255 (
		_w29586_,
		_w29587_,
		_w29767_
	);
	LUT2 #(
		.INIT('h1)
	) name19256 (
		_w29588_,
		_w29589_,
		_w29768_
	);
	LUT2 #(
		.INIT('h1)
	) name19257 (
		_w29590_,
		_w29591_,
		_w29769_
	);
	LUT2 #(
		.INIT('h1)
	) name19258 (
		_w29592_,
		_w29593_,
		_w29770_
	);
	LUT2 #(
		.INIT('h1)
	) name19259 (
		_w29594_,
		_w29595_,
		_w29771_
	);
	LUT2 #(
		.INIT('h1)
	) name19260 (
		_w29596_,
		_w29597_,
		_w29772_
	);
	LUT2 #(
		.INIT('h1)
	) name19261 (
		_w29598_,
		_w29599_,
		_w29773_
	);
	LUT2 #(
		.INIT('h1)
	) name19262 (
		_w29600_,
		_w29601_,
		_w29774_
	);
	LUT2 #(
		.INIT('h1)
	) name19263 (
		_w29602_,
		_w29603_,
		_w29775_
	);
	LUT2 #(
		.INIT('h1)
	) name19264 (
		_w29604_,
		_w29605_,
		_w29776_
	);
	LUT2 #(
		.INIT('h1)
	) name19265 (
		_w29606_,
		_w29607_,
		_w29777_
	);
	LUT2 #(
		.INIT('h1)
	) name19266 (
		_w29608_,
		_w29609_,
		_w29778_
	);
	LUT2 #(
		.INIT('h1)
	) name19267 (
		_w29610_,
		_w29611_,
		_w29779_
	);
	LUT2 #(
		.INIT('h1)
	) name19268 (
		_w29612_,
		_w29613_,
		_w29780_
	);
	LUT2 #(
		.INIT('h1)
	) name19269 (
		_w29614_,
		_w29615_,
		_w29781_
	);
	LUT2 #(
		.INIT('h1)
	) name19270 (
		_w29616_,
		_w29617_,
		_w29782_
	);
	LUT2 #(
		.INIT('h1)
	) name19271 (
		_w29618_,
		_w29619_,
		_w29783_
	);
	LUT2 #(
		.INIT('h1)
	) name19272 (
		_w29620_,
		_w29621_,
		_w29784_
	);
	LUT2 #(
		.INIT('h1)
	) name19273 (
		_w29622_,
		_w29623_,
		_w29785_
	);
	LUT2 #(
		.INIT('h1)
	) name19274 (
		_w29624_,
		_w29625_,
		_w29786_
	);
	LUT2 #(
		.INIT('h1)
	) name19275 (
		_w29626_,
		_w29627_,
		_w29787_
	);
	LUT2 #(
		.INIT('h1)
	) name19276 (
		_w29628_,
		_w29629_,
		_w29788_
	);
	LUT2 #(
		.INIT('h1)
	) name19277 (
		_w29630_,
		_w29631_,
		_w29789_
	);
	LUT2 #(
		.INIT('h1)
	) name19278 (
		_w29632_,
		_w29633_,
		_w29790_
	);
	LUT2 #(
		.INIT('h1)
	) name19279 (
		_w29634_,
		_w29635_,
		_w29791_
	);
	LUT2 #(
		.INIT('h1)
	) name19280 (
		_w29636_,
		_w29637_,
		_w29792_
	);
	LUT2 #(
		.INIT('h1)
	) name19281 (
		_w29638_,
		_w29639_,
		_w29793_
	);
	LUT2 #(
		.INIT('h1)
	) name19282 (
		_w29640_,
		_w29641_,
		_w29794_
	);
	LUT2 #(
		.INIT('h1)
	) name19283 (
		_w29642_,
		_w29643_,
		_w29795_
	);
	LUT2 #(
		.INIT('h1)
	) name19284 (
		_w29644_,
		_w29645_,
		_w29796_
	);
	LUT2 #(
		.INIT('h1)
	) name19285 (
		_w29646_,
		_w29647_,
		_w29797_
	);
	LUT2 #(
		.INIT('h1)
	) name19286 (
		_w29648_,
		_w29649_,
		_w29798_
	);
	LUT2 #(
		.INIT('h1)
	) name19287 (
		_w29650_,
		_w29651_,
		_w29799_
	);
	LUT2 #(
		.INIT('h1)
	) name19288 (
		_w29652_,
		_w29653_,
		_w29800_
	);
	LUT2 #(
		.INIT('h1)
	) name19289 (
		_w29654_,
		_w29655_,
		_w29801_
	);
	LUT2 #(
		.INIT('h1)
	) name19290 (
		_w29656_,
		_w29657_,
		_w29802_
	);
	LUT2 #(
		.INIT('h1)
	) name19291 (
		_w29658_,
		_w29659_,
		_w29803_
	);
	LUT2 #(
		.INIT('h1)
	) name19292 (
		_w29660_,
		_w29661_,
		_w29804_
	);
	LUT2 #(
		.INIT('h1)
	) name19293 (
		_w29662_,
		_w29663_,
		_w29805_
	);
	LUT2 #(
		.INIT('h1)
	) name19294 (
		_w29664_,
		_w29665_,
		_w29806_
	);
	LUT2 #(
		.INIT('h1)
	) name19295 (
		_w29666_,
		_w29667_,
		_w29807_
	);
	LUT2 #(
		.INIT('h1)
	) name19296 (
		_w29668_,
		_w29669_,
		_w29808_
	);
	LUT2 #(
		.INIT('h1)
	) name19297 (
		_w29670_,
		_w29671_,
		_w29809_
	);
	LUT2 #(
		.INIT('h1)
	) name19298 (
		_w29672_,
		_w29673_,
		_w29810_
	);
	LUT2 #(
		.INIT('h1)
	) name19299 (
		_w29674_,
		_w29675_,
		_w29811_
	);
	LUT2 #(
		.INIT('h1)
	) name19300 (
		_w29676_,
		_w29677_,
		_w29812_
	);
	LUT2 #(
		.INIT('h1)
	) name19301 (
		_w29678_,
		_w29679_,
		_w29813_
	);
	LUT2 #(
		.INIT('h1)
	) name19302 (
		_w29680_,
		_w29681_,
		_w29814_
	);
	LUT2 #(
		.INIT('h1)
	) name19303 (
		_w29682_,
		_w29683_,
		_w29815_
	);
	LUT2 #(
		.INIT('h1)
	) name19304 (
		_w29684_,
		_w29685_,
		_w29816_
	);
	LUT2 #(
		.INIT('h1)
	) name19305 (
		_w29686_,
		_w29687_,
		_w29817_
	);
	LUT2 #(
		.INIT('h1)
	) name19306 (
		_w29688_,
		_w29689_,
		_w29818_
	);
	LUT2 #(
		.INIT('h1)
	) name19307 (
		_w29690_,
		_w29691_,
		_w29819_
	);
	LUT2 #(
		.INIT('h8)
	) name19308 (
		_w29818_,
		_w29819_,
		_w29820_
	);
	LUT2 #(
		.INIT('h8)
	) name19309 (
		_w29816_,
		_w29817_,
		_w29821_
	);
	LUT2 #(
		.INIT('h8)
	) name19310 (
		_w29814_,
		_w29815_,
		_w29822_
	);
	LUT2 #(
		.INIT('h8)
	) name19311 (
		_w29812_,
		_w29813_,
		_w29823_
	);
	LUT2 #(
		.INIT('h8)
	) name19312 (
		_w29810_,
		_w29811_,
		_w29824_
	);
	LUT2 #(
		.INIT('h8)
	) name19313 (
		_w29808_,
		_w29809_,
		_w29825_
	);
	LUT2 #(
		.INIT('h8)
	) name19314 (
		_w29806_,
		_w29807_,
		_w29826_
	);
	LUT2 #(
		.INIT('h8)
	) name19315 (
		_w29804_,
		_w29805_,
		_w29827_
	);
	LUT2 #(
		.INIT('h8)
	) name19316 (
		_w29802_,
		_w29803_,
		_w29828_
	);
	LUT2 #(
		.INIT('h8)
	) name19317 (
		_w29800_,
		_w29801_,
		_w29829_
	);
	LUT2 #(
		.INIT('h8)
	) name19318 (
		_w29798_,
		_w29799_,
		_w29830_
	);
	LUT2 #(
		.INIT('h8)
	) name19319 (
		_w29796_,
		_w29797_,
		_w29831_
	);
	LUT2 #(
		.INIT('h8)
	) name19320 (
		_w29794_,
		_w29795_,
		_w29832_
	);
	LUT2 #(
		.INIT('h8)
	) name19321 (
		_w29792_,
		_w29793_,
		_w29833_
	);
	LUT2 #(
		.INIT('h8)
	) name19322 (
		_w29790_,
		_w29791_,
		_w29834_
	);
	LUT2 #(
		.INIT('h8)
	) name19323 (
		_w29788_,
		_w29789_,
		_w29835_
	);
	LUT2 #(
		.INIT('h8)
	) name19324 (
		_w29786_,
		_w29787_,
		_w29836_
	);
	LUT2 #(
		.INIT('h8)
	) name19325 (
		_w29784_,
		_w29785_,
		_w29837_
	);
	LUT2 #(
		.INIT('h8)
	) name19326 (
		_w29782_,
		_w29783_,
		_w29838_
	);
	LUT2 #(
		.INIT('h8)
	) name19327 (
		_w29780_,
		_w29781_,
		_w29839_
	);
	LUT2 #(
		.INIT('h8)
	) name19328 (
		_w29778_,
		_w29779_,
		_w29840_
	);
	LUT2 #(
		.INIT('h8)
	) name19329 (
		_w29776_,
		_w29777_,
		_w29841_
	);
	LUT2 #(
		.INIT('h8)
	) name19330 (
		_w29774_,
		_w29775_,
		_w29842_
	);
	LUT2 #(
		.INIT('h8)
	) name19331 (
		_w29772_,
		_w29773_,
		_w29843_
	);
	LUT2 #(
		.INIT('h8)
	) name19332 (
		_w29770_,
		_w29771_,
		_w29844_
	);
	LUT2 #(
		.INIT('h8)
	) name19333 (
		_w29768_,
		_w29769_,
		_w29845_
	);
	LUT2 #(
		.INIT('h8)
	) name19334 (
		_w29766_,
		_w29767_,
		_w29846_
	);
	LUT2 #(
		.INIT('h8)
	) name19335 (
		_w29764_,
		_w29765_,
		_w29847_
	);
	LUT2 #(
		.INIT('h8)
	) name19336 (
		_w29762_,
		_w29763_,
		_w29848_
	);
	LUT2 #(
		.INIT('h8)
	) name19337 (
		_w29760_,
		_w29761_,
		_w29849_
	);
	LUT2 #(
		.INIT('h8)
	) name19338 (
		_w29758_,
		_w29759_,
		_w29850_
	);
	LUT2 #(
		.INIT('h8)
	) name19339 (
		_w29756_,
		_w29757_,
		_w29851_
	);
	LUT2 #(
		.INIT('h8)
	) name19340 (
		_w29754_,
		_w29755_,
		_w29852_
	);
	LUT2 #(
		.INIT('h8)
	) name19341 (
		_w29752_,
		_w29753_,
		_w29853_
	);
	LUT2 #(
		.INIT('h8)
	) name19342 (
		_w29750_,
		_w29751_,
		_w29854_
	);
	LUT2 #(
		.INIT('h8)
	) name19343 (
		_w29748_,
		_w29749_,
		_w29855_
	);
	LUT2 #(
		.INIT('h8)
	) name19344 (
		_w29746_,
		_w29747_,
		_w29856_
	);
	LUT2 #(
		.INIT('h8)
	) name19345 (
		_w29744_,
		_w29745_,
		_w29857_
	);
	LUT2 #(
		.INIT('h8)
	) name19346 (
		_w29742_,
		_w29743_,
		_w29858_
	);
	LUT2 #(
		.INIT('h8)
	) name19347 (
		_w29740_,
		_w29741_,
		_w29859_
	);
	LUT2 #(
		.INIT('h8)
	) name19348 (
		_w29738_,
		_w29739_,
		_w29860_
	);
	LUT2 #(
		.INIT('h8)
	) name19349 (
		_w29736_,
		_w29737_,
		_w29861_
	);
	LUT2 #(
		.INIT('h8)
	) name19350 (
		_w29734_,
		_w29735_,
		_w29862_
	);
	LUT2 #(
		.INIT('h8)
	) name19351 (
		_w29732_,
		_w29733_,
		_w29863_
	);
	LUT2 #(
		.INIT('h8)
	) name19352 (
		_w29730_,
		_w29731_,
		_w29864_
	);
	LUT2 #(
		.INIT('h8)
	) name19353 (
		_w29728_,
		_w29729_,
		_w29865_
	);
	LUT2 #(
		.INIT('h8)
	) name19354 (
		_w29726_,
		_w29727_,
		_w29866_
	);
	LUT2 #(
		.INIT('h8)
	) name19355 (
		_w29724_,
		_w29725_,
		_w29867_
	);
	LUT2 #(
		.INIT('h8)
	) name19356 (
		_w29722_,
		_w29723_,
		_w29868_
	);
	LUT2 #(
		.INIT('h8)
	) name19357 (
		_w29720_,
		_w29721_,
		_w29869_
	);
	LUT2 #(
		.INIT('h8)
	) name19358 (
		_w29718_,
		_w29719_,
		_w29870_
	);
	LUT2 #(
		.INIT('h8)
	) name19359 (
		_w29716_,
		_w29717_,
		_w29871_
	);
	LUT2 #(
		.INIT('h8)
	) name19360 (
		_w29714_,
		_w29715_,
		_w29872_
	);
	LUT2 #(
		.INIT('h8)
	) name19361 (
		_w29712_,
		_w29713_,
		_w29873_
	);
	LUT2 #(
		.INIT('h8)
	) name19362 (
		_w29710_,
		_w29711_,
		_w29874_
	);
	LUT2 #(
		.INIT('h8)
	) name19363 (
		_w29708_,
		_w29709_,
		_w29875_
	);
	LUT2 #(
		.INIT('h8)
	) name19364 (
		_w29706_,
		_w29707_,
		_w29876_
	);
	LUT2 #(
		.INIT('h8)
	) name19365 (
		_w29704_,
		_w29705_,
		_w29877_
	);
	LUT2 #(
		.INIT('h8)
	) name19366 (
		_w29702_,
		_w29703_,
		_w29878_
	);
	LUT2 #(
		.INIT('h8)
	) name19367 (
		_w29700_,
		_w29701_,
		_w29879_
	);
	LUT2 #(
		.INIT('h8)
	) name19368 (
		_w29698_,
		_w29699_,
		_w29880_
	);
	LUT2 #(
		.INIT('h8)
	) name19369 (
		_w29696_,
		_w29697_,
		_w29881_
	);
	LUT2 #(
		.INIT('h8)
	) name19370 (
		_w29694_,
		_w29695_,
		_w29882_
	);
	LUT2 #(
		.INIT('h8)
	) name19371 (
		_w29692_,
		_w29693_,
		_w29883_
	);
	LUT2 #(
		.INIT('h8)
	) name19372 (
		_w29882_,
		_w29883_,
		_w29884_
	);
	LUT2 #(
		.INIT('h8)
	) name19373 (
		_w29880_,
		_w29881_,
		_w29885_
	);
	LUT2 #(
		.INIT('h8)
	) name19374 (
		_w29878_,
		_w29879_,
		_w29886_
	);
	LUT2 #(
		.INIT('h8)
	) name19375 (
		_w29876_,
		_w29877_,
		_w29887_
	);
	LUT2 #(
		.INIT('h8)
	) name19376 (
		_w29874_,
		_w29875_,
		_w29888_
	);
	LUT2 #(
		.INIT('h8)
	) name19377 (
		_w29872_,
		_w29873_,
		_w29889_
	);
	LUT2 #(
		.INIT('h8)
	) name19378 (
		_w29870_,
		_w29871_,
		_w29890_
	);
	LUT2 #(
		.INIT('h8)
	) name19379 (
		_w29868_,
		_w29869_,
		_w29891_
	);
	LUT2 #(
		.INIT('h8)
	) name19380 (
		_w29866_,
		_w29867_,
		_w29892_
	);
	LUT2 #(
		.INIT('h8)
	) name19381 (
		_w29864_,
		_w29865_,
		_w29893_
	);
	LUT2 #(
		.INIT('h8)
	) name19382 (
		_w29862_,
		_w29863_,
		_w29894_
	);
	LUT2 #(
		.INIT('h8)
	) name19383 (
		_w29860_,
		_w29861_,
		_w29895_
	);
	LUT2 #(
		.INIT('h8)
	) name19384 (
		_w29858_,
		_w29859_,
		_w29896_
	);
	LUT2 #(
		.INIT('h8)
	) name19385 (
		_w29856_,
		_w29857_,
		_w29897_
	);
	LUT2 #(
		.INIT('h8)
	) name19386 (
		_w29854_,
		_w29855_,
		_w29898_
	);
	LUT2 #(
		.INIT('h8)
	) name19387 (
		_w29852_,
		_w29853_,
		_w29899_
	);
	LUT2 #(
		.INIT('h8)
	) name19388 (
		_w29850_,
		_w29851_,
		_w29900_
	);
	LUT2 #(
		.INIT('h8)
	) name19389 (
		_w29848_,
		_w29849_,
		_w29901_
	);
	LUT2 #(
		.INIT('h8)
	) name19390 (
		_w29846_,
		_w29847_,
		_w29902_
	);
	LUT2 #(
		.INIT('h8)
	) name19391 (
		_w29844_,
		_w29845_,
		_w29903_
	);
	LUT2 #(
		.INIT('h8)
	) name19392 (
		_w29842_,
		_w29843_,
		_w29904_
	);
	LUT2 #(
		.INIT('h8)
	) name19393 (
		_w29840_,
		_w29841_,
		_w29905_
	);
	LUT2 #(
		.INIT('h8)
	) name19394 (
		_w29838_,
		_w29839_,
		_w29906_
	);
	LUT2 #(
		.INIT('h8)
	) name19395 (
		_w29836_,
		_w29837_,
		_w29907_
	);
	LUT2 #(
		.INIT('h8)
	) name19396 (
		_w29834_,
		_w29835_,
		_w29908_
	);
	LUT2 #(
		.INIT('h8)
	) name19397 (
		_w29832_,
		_w29833_,
		_w29909_
	);
	LUT2 #(
		.INIT('h8)
	) name19398 (
		_w29830_,
		_w29831_,
		_w29910_
	);
	LUT2 #(
		.INIT('h8)
	) name19399 (
		_w29828_,
		_w29829_,
		_w29911_
	);
	LUT2 #(
		.INIT('h8)
	) name19400 (
		_w29826_,
		_w29827_,
		_w29912_
	);
	LUT2 #(
		.INIT('h8)
	) name19401 (
		_w29824_,
		_w29825_,
		_w29913_
	);
	LUT2 #(
		.INIT('h8)
	) name19402 (
		_w29822_,
		_w29823_,
		_w29914_
	);
	LUT2 #(
		.INIT('h8)
	) name19403 (
		_w29820_,
		_w29821_,
		_w29915_
	);
	LUT2 #(
		.INIT('h8)
	) name19404 (
		_w29914_,
		_w29915_,
		_w29916_
	);
	LUT2 #(
		.INIT('h8)
	) name19405 (
		_w29912_,
		_w29913_,
		_w29917_
	);
	LUT2 #(
		.INIT('h8)
	) name19406 (
		_w29910_,
		_w29911_,
		_w29918_
	);
	LUT2 #(
		.INIT('h8)
	) name19407 (
		_w29908_,
		_w29909_,
		_w29919_
	);
	LUT2 #(
		.INIT('h8)
	) name19408 (
		_w29906_,
		_w29907_,
		_w29920_
	);
	LUT2 #(
		.INIT('h8)
	) name19409 (
		_w29904_,
		_w29905_,
		_w29921_
	);
	LUT2 #(
		.INIT('h8)
	) name19410 (
		_w29902_,
		_w29903_,
		_w29922_
	);
	LUT2 #(
		.INIT('h8)
	) name19411 (
		_w29900_,
		_w29901_,
		_w29923_
	);
	LUT2 #(
		.INIT('h8)
	) name19412 (
		_w29898_,
		_w29899_,
		_w29924_
	);
	LUT2 #(
		.INIT('h8)
	) name19413 (
		_w29896_,
		_w29897_,
		_w29925_
	);
	LUT2 #(
		.INIT('h8)
	) name19414 (
		_w29894_,
		_w29895_,
		_w29926_
	);
	LUT2 #(
		.INIT('h8)
	) name19415 (
		_w29892_,
		_w29893_,
		_w29927_
	);
	LUT2 #(
		.INIT('h8)
	) name19416 (
		_w29890_,
		_w29891_,
		_w29928_
	);
	LUT2 #(
		.INIT('h8)
	) name19417 (
		_w29888_,
		_w29889_,
		_w29929_
	);
	LUT2 #(
		.INIT('h8)
	) name19418 (
		_w29886_,
		_w29887_,
		_w29930_
	);
	LUT2 #(
		.INIT('h8)
	) name19419 (
		_w29884_,
		_w29885_,
		_w29931_
	);
	LUT2 #(
		.INIT('h8)
	) name19420 (
		_w29930_,
		_w29931_,
		_w29932_
	);
	LUT2 #(
		.INIT('h8)
	) name19421 (
		_w29928_,
		_w29929_,
		_w29933_
	);
	LUT2 #(
		.INIT('h8)
	) name19422 (
		_w29926_,
		_w29927_,
		_w29934_
	);
	LUT2 #(
		.INIT('h8)
	) name19423 (
		_w29924_,
		_w29925_,
		_w29935_
	);
	LUT2 #(
		.INIT('h8)
	) name19424 (
		_w29922_,
		_w29923_,
		_w29936_
	);
	LUT2 #(
		.INIT('h8)
	) name19425 (
		_w29920_,
		_w29921_,
		_w29937_
	);
	LUT2 #(
		.INIT('h8)
	) name19426 (
		_w29918_,
		_w29919_,
		_w29938_
	);
	LUT2 #(
		.INIT('h8)
	) name19427 (
		_w29916_,
		_w29917_,
		_w29939_
	);
	LUT2 #(
		.INIT('h8)
	) name19428 (
		_w29938_,
		_w29939_,
		_w29940_
	);
	LUT2 #(
		.INIT('h8)
	) name19429 (
		_w29936_,
		_w29937_,
		_w29941_
	);
	LUT2 #(
		.INIT('h8)
	) name19430 (
		_w29934_,
		_w29935_,
		_w29942_
	);
	LUT2 #(
		.INIT('h8)
	) name19431 (
		_w29932_,
		_w29933_,
		_w29943_
	);
	LUT2 #(
		.INIT('h8)
	) name19432 (
		_w29942_,
		_w29943_,
		_w29944_
	);
	LUT2 #(
		.INIT('h8)
	) name19433 (
		_w29940_,
		_w29941_,
		_w29945_
	);
	LUT2 #(
		.INIT('h8)
	) name19434 (
		_w29944_,
		_w29945_,
		_w29946_
	);
	LUT2 #(
		.INIT('h1)
	) name19435 (
		wb_rst_i_pad,
		_w29946_,
		_w29947_
	);
	LUT2 #(
		.INIT('h1)
	) name19436 (
		_w22944_,
		_w29947_,
		_w29948_
	);
	LUT2 #(
		.INIT('h8)
	) name19437 (
		\ethreg1_MODER_1_DataOut_reg[5]/NET0131 ,
		_w23519_,
		_w29949_
	);
	LUT2 #(
		.INIT('h8)
	) name19438 (
		\ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 ,
		_w23499_,
		_w29950_
	);
	LUT2 #(
		.INIT('h8)
	) name19439 (
		\ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 ,
		_w22952_,
		_w29951_
	);
	LUT2 #(
		.INIT('h8)
	) name19440 (
		\ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 ,
		_w22956_,
		_w29952_
	);
	LUT2 #(
		.INIT('h8)
	) name19441 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 ,
		_w23522_,
		_w29953_
	);
	LUT2 #(
		.INIT('h8)
	) name19442 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		_w22959_,
		_w29954_
	);
	LUT2 #(
		.INIT('h8)
	) name19443 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		_w23501_,
		_w29955_
	);
	LUT2 #(
		.INIT('h8)
	) name19444 (
		\ethreg1_MIIRX_DATA_DataOut_reg[13]/NET0131 ,
		_w23507_,
		_w29956_
	);
	LUT2 #(
		.INIT('h8)
	) name19445 (
		\ethreg1_PACKETLEN_1_DataOut_reg[5]/NET0131 ,
		_w22966_,
		_w29957_
	);
	LUT2 #(
		.INIT('h1)
	) name19446 (
		_w29949_,
		_w29950_,
		_w29958_
	);
	LUT2 #(
		.INIT('h1)
	) name19447 (
		_w29951_,
		_w29952_,
		_w29959_
	);
	LUT2 #(
		.INIT('h1)
	) name19448 (
		_w29953_,
		_w29954_,
		_w29960_
	);
	LUT2 #(
		.INIT('h1)
	) name19449 (
		_w29955_,
		_w29956_,
		_w29961_
	);
	LUT2 #(
		.INIT('h8)
	) name19450 (
		_w29960_,
		_w29961_,
		_w29962_
	);
	LUT2 #(
		.INIT('h8)
	) name19451 (
		_w29958_,
		_w29959_,
		_w29963_
	);
	LUT2 #(
		.INIT('h8)
	) name19452 (
		_w22944_,
		_w29963_,
		_w29964_
	);
	LUT2 #(
		.INIT('h4)
	) name19453 (
		_w29957_,
		_w29962_,
		_w29965_
	);
	LUT2 #(
		.INIT('h8)
	) name19454 (
		_w29964_,
		_w29965_,
		_w29966_
	);
	LUT2 #(
		.INIT('h1)
	) name19455 (
		_w29948_,
		_w29966_,
		_w29967_
	);
	LUT2 #(
		.INIT('h8)
	) name19456 (
		\wishbone_bd_ram_mem1_reg[18][14]/P0001 ,
		_w12679_,
		_w29968_
	);
	LUT2 #(
		.INIT('h8)
	) name19457 (
		\wishbone_bd_ram_mem1_reg[58][14]/P0001 ,
		_w13070_,
		_w29969_
	);
	LUT2 #(
		.INIT('h8)
	) name19458 (
		\wishbone_bd_ram_mem1_reg[171][14]/P0001 ,
		_w12910_,
		_w29970_
	);
	LUT2 #(
		.INIT('h8)
	) name19459 (
		\wishbone_bd_ram_mem1_reg[118][14]/P0001 ,
		_w12830_,
		_w29971_
	);
	LUT2 #(
		.INIT('h8)
	) name19460 (
		\wishbone_bd_ram_mem1_reg[33][14]/P0001 ,
		_w12980_,
		_w29972_
	);
	LUT2 #(
		.INIT('h8)
	) name19461 (
		\wishbone_bd_ram_mem1_reg[113][14]/P0001 ,
		_w13026_,
		_w29973_
	);
	LUT2 #(
		.INIT('h8)
	) name19462 (
		\wishbone_bd_ram_mem1_reg[44][14]/P0001 ,
		_w12896_,
		_w29974_
	);
	LUT2 #(
		.INIT('h8)
	) name19463 (
		\wishbone_bd_ram_mem1_reg[237][14]/P0001 ,
		_w12990_,
		_w29975_
	);
	LUT2 #(
		.INIT('h8)
	) name19464 (
		\wishbone_bd_ram_mem1_reg[29][14]/P0001 ,
		_w12952_,
		_w29976_
	);
	LUT2 #(
		.INIT('h8)
	) name19465 (
		\wishbone_bd_ram_mem1_reg[241][14]/P0001 ,
		_w13006_,
		_w29977_
	);
	LUT2 #(
		.INIT('h8)
	) name19466 (
		\wishbone_bd_ram_mem1_reg[211][14]/P0001 ,
		_w13166_,
		_w29978_
	);
	LUT2 #(
		.INIT('h8)
	) name19467 (
		\wishbone_bd_ram_mem1_reg[66][14]/P0001 ,
		_w12824_,
		_w29979_
	);
	LUT2 #(
		.INIT('h8)
	) name19468 (
		\wishbone_bd_ram_mem1_reg[78][14]/P0001 ,
		_w12874_,
		_w29980_
	);
	LUT2 #(
		.INIT('h8)
	) name19469 (
		\wishbone_bd_ram_mem1_reg[46][14]/P0001 ,
		_w12884_,
		_w29981_
	);
	LUT2 #(
		.INIT('h8)
	) name19470 (
		\wishbone_bd_ram_mem1_reg[157][14]/P0001 ,
		_w12926_,
		_w29982_
	);
	LUT2 #(
		.INIT('h8)
	) name19471 (
		\wishbone_bd_ram_mem1_reg[81][14]/P0001 ,
		_w12950_,
		_w29983_
	);
	LUT2 #(
		.INIT('h8)
	) name19472 (
		\wishbone_bd_ram_mem1_reg[197][14]/P0001 ,
		_w12834_,
		_w29984_
	);
	LUT2 #(
		.INIT('h8)
	) name19473 (
		\wishbone_bd_ram_mem1_reg[222][14]/P0001 ,
		_w13094_,
		_w29985_
	);
	LUT2 #(
		.INIT('h8)
	) name19474 (
		\wishbone_bd_ram_mem1_reg[16][14]/P0001 ,
		_w13140_,
		_w29986_
	);
	LUT2 #(
		.INIT('h8)
	) name19475 (
		\wishbone_bd_ram_mem1_reg[135][14]/P0001 ,
		_w13124_,
		_w29987_
	);
	LUT2 #(
		.INIT('h8)
	) name19476 (
		\wishbone_bd_ram_mem1_reg[68][14]/P0001 ,
		_w12946_,
		_w29988_
	);
	LUT2 #(
		.INIT('h8)
	) name19477 (
		\wishbone_bd_ram_mem1_reg[132][14]/P0001 ,
		_w12992_,
		_w29989_
	);
	LUT2 #(
		.INIT('h8)
	) name19478 (
		\wishbone_bd_ram_mem1_reg[87][14]/P0001 ,
		_w13154_,
		_w29990_
	);
	LUT2 #(
		.INIT('h8)
	) name19479 (
		\wishbone_bd_ram_mem1_reg[108][14]/P0001 ,
		_w13156_,
		_w29991_
	);
	LUT2 #(
		.INIT('h8)
	) name19480 (
		\wishbone_bd_ram_mem1_reg[210][14]/P0001 ,
		_w12924_,
		_w29992_
	);
	LUT2 #(
		.INIT('h8)
	) name19481 (
		\wishbone_bd_ram_mem1_reg[85][14]/P0001 ,
		_w13216_,
		_w29993_
	);
	LUT2 #(
		.INIT('h8)
	) name19482 (
		\wishbone_bd_ram_mem1_reg[50][14]/P0001 ,
		_w13150_,
		_w29994_
	);
	LUT2 #(
		.INIT('h8)
	) name19483 (
		\wishbone_bd_ram_mem1_reg[176][14]/P0001 ,
		_w12868_,
		_w29995_
	);
	LUT2 #(
		.INIT('h8)
	) name19484 (
		\wishbone_bd_ram_mem1_reg[75][14]/P0001 ,
		_w12826_,
		_w29996_
	);
	LUT2 #(
		.INIT('h8)
	) name19485 (
		\wishbone_bd_ram_mem1_reg[70][14]/P0001 ,
		_w12840_,
		_w29997_
	);
	LUT2 #(
		.INIT('h8)
	) name19486 (
		\wishbone_bd_ram_mem1_reg[155][14]/P0001 ,
		_w13122_,
		_w29998_
	);
	LUT2 #(
		.INIT('h8)
	) name19487 (
		\wishbone_bd_ram_mem1_reg[243][14]/P0001 ,
		_w12804_,
		_w29999_
	);
	LUT2 #(
		.INIT('h8)
	) name19488 (
		\wishbone_bd_ram_mem1_reg[14][14]/P0001 ,
		_w13086_,
		_w30000_
	);
	LUT2 #(
		.INIT('h8)
	) name19489 (
		\wishbone_bd_ram_mem1_reg[93][14]/P0001 ,
		_w13016_,
		_w30001_
	);
	LUT2 #(
		.INIT('h8)
	) name19490 (
		\wishbone_bd_ram_mem1_reg[32][14]/P0001 ,
		_w13120_,
		_w30002_
	);
	LUT2 #(
		.INIT('h8)
	) name19491 (
		\wishbone_bd_ram_mem1_reg[215][14]/P0001 ,
		_w12974_,
		_w30003_
	);
	LUT2 #(
		.INIT('h8)
	) name19492 (
		\wishbone_bd_ram_mem1_reg[17][14]/P0001 ,
		_w12848_,
		_w30004_
	);
	LUT2 #(
		.INIT('h8)
	) name19493 (
		\wishbone_bd_ram_mem1_reg[25][14]/P0001 ,
		_w13108_,
		_w30005_
	);
	LUT2 #(
		.INIT('h8)
	) name19494 (
		\wishbone_bd_ram_mem1_reg[105][14]/P0001 ,
		_w12751_,
		_w30006_
	);
	LUT2 #(
		.INIT('h8)
	) name19495 (
		\wishbone_bd_ram_mem1_reg[234][14]/P0001 ,
		_w13214_,
		_w30007_
	);
	LUT2 #(
		.INIT('h8)
	) name19496 (
		\wishbone_bd_ram_mem1_reg[185][14]/P0001 ,
		_w12940_,
		_w30008_
	);
	LUT2 #(
		.INIT('h8)
	) name19497 (
		\wishbone_bd_ram_mem1_reg[129][14]/P0001 ,
		_w12776_,
		_w30009_
	);
	LUT2 #(
		.INIT('h8)
	) name19498 (
		\wishbone_bd_ram_mem1_reg[240][14]/P0001 ,
		_w12864_,
		_w30010_
	);
	LUT2 #(
		.INIT('h8)
	) name19499 (
		\wishbone_bd_ram_mem1_reg[175][14]/P0001 ,
		_w13126_,
		_w30011_
	);
	LUT2 #(
		.INIT('h8)
	) name19500 (
		\wishbone_bd_ram_mem1_reg[199][14]/P0001 ,
		_w12768_,
		_w30012_
	);
	LUT2 #(
		.INIT('h8)
	) name19501 (
		\wishbone_bd_ram_mem1_reg[133][14]/P0001 ,
		_w12761_,
		_w30013_
	);
	LUT2 #(
		.INIT('h8)
	) name19502 (
		\wishbone_bd_ram_mem1_reg[165][14]/P0001 ,
		_w13044_,
		_w30014_
	);
	LUT2 #(
		.INIT('h8)
	) name19503 (
		\wishbone_bd_ram_mem1_reg[169][14]/P0001 ,
		_w12722_,
		_w30015_
	);
	LUT2 #(
		.INIT('h8)
	) name19504 (
		\wishbone_bd_ram_mem1_reg[212][14]/P0001 ,
		_w12796_,
		_w30016_
	);
	LUT2 #(
		.INIT('h8)
	) name19505 (
		\wishbone_bd_ram_mem1_reg[233][14]/P0001 ,
		_w12836_,
		_w30017_
	);
	LUT2 #(
		.INIT('h8)
	) name19506 (
		\wishbone_bd_ram_mem1_reg[43][14]/P0001 ,
		_w13200_,
		_w30018_
	);
	LUT2 #(
		.INIT('h8)
	) name19507 (
		\wishbone_bd_ram_mem1_reg[27][14]/P0001 ,
		_w12880_,
		_w30019_
	);
	LUT2 #(
		.INIT('h8)
	) name19508 (
		\wishbone_bd_ram_mem1_reg[138][14]/P0001 ,
		_w12958_,
		_w30020_
	);
	LUT2 #(
		.INIT('h8)
	) name19509 (
		\wishbone_bd_ram_mem1_reg[116][14]/P0001 ,
		_w12998_,
		_w30021_
	);
	LUT2 #(
		.INIT('h8)
	) name19510 (
		\wishbone_bd_ram_mem1_reg[121][14]/P0001 ,
		_w13078_,
		_w30022_
	);
	LUT2 #(
		.INIT('h8)
	) name19511 (
		\wishbone_bd_ram_mem1_reg[204][14]/P0001 ,
		_w13162_,
		_w30023_
	);
	LUT2 #(
		.INIT('h8)
	) name19512 (
		\wishbone_bd_ram_mem1_reg[125][14]/P0001 ,
		_w12956_,
		_w30024_
	);
	LUT2 #(
		.INIT('h8)
	) name19513 (
		\wishbone_bd_ram_mem1_reg[219][14]/P0001 ,
		_w12806_,
		_w30025_
	);
	LUT2 #(
		.INIT('h8)
	) name19514 (
		\wishbone_bd_ram_mem1_reg[11][14]/P0001 ,
		_w13194_,
		_w30026_
	);
	LUT2 #(
		.INIT('h8)
	) name19515 (
		\wishbone_bd_ram_mem1_reg[36][14]/P0001 ,
		_w12800_,
		_w30027_
	);
	LUT2 #(
		.INIT('h8)
	) name19516 (
		\wishbone_bd_ram_mem1_reg[178][14]/P0001 ,
		_w12886_,
		_w30028_
	);
	LUT2 #(
		.INIT('h8)
	) name19517 (
		\wishbone_bd_ram_mem1_reg[1][14]/P0001 ,
		_w13014_,
		_w30029_
	);
	LUT2 #(
		.INIT('h8)
	) name19518 (
		\wishbone_bd_ram_mem1_reg[232][14]/P0001 ,
		_w12758_,
		_w30030_
	);
	LUT2 #(
		.INIT('h8)
	) name19519 (
		\wishbone_bd_ram_mem1_reg[235][14]/P0001 ,
		_w12696_,
		_w30031_
	);
	LUT2 #(
		.INIT('h8)
	) name19520 (
		\wishbone_bd_ram_mem1_reg[114][14]/P0001 ,
		_w13202_,
		_w30032_
	);
	LUT2 #(
		.INIT('h8)
	) name19521 (
		\wishbone_bd_ram_mem1_reg[209][14]/P0001 ,
		_w13152_,
		_w30033_
	);
	LUT2 #(
		.INIT('h8)
	) name19522 (
		\wishbone_bd_ram_mem1_reg[28][14]/P0001 ,
		_w13170_,
		_w30034_
	);
	LUT2 #(
		.INIT('h8)
	) name19523 (
		\wishbone_bd_ram_mem1_reg[69][14]/P0001 ,
		_w12738_,
		_w30035_
	);
	LUT2 #(
		.INIT('h8)
	) name19524 (
		\wishbone_bd_ram_mem1_reg[0][14]/P0001 ,
		_w12717_,
		_w30036_
	);
	LUT2 #(
		.INIT('h8)
	) name19525 (
		\wishbone_bd_ram_mem1_reg[56][14]/P0001 ,
		_w12778_,
		_w30037_
	);
	LUT2 #(
		.INIT('h8)
	) name19526 (
		\wishbone_bd_ram_mem1_reg[247][14]/P0001 ,
		_w12818_,
		_w30038_
	);
	LUT2 #(
		.INIT('h8)
	) name19527 (
		\wishbone_bd_ram_mem1_reg[101][14]/P0001 ,
		_w13192_,
		_w30039_
	);
	LUT2 #(
		.INIT('h8)
	) name19528 (
		\wishbone_bd_ram_mem1_reg[242][14]/P0001 ,
		_w12932_,
		_w30040_
	);
	LUT2 #(
		.INIT('h8)
	) name19529 (
		\wishbone_bd_ram_mem1_reg[223][14]/P0001 ,
		_w12838_,
		_w30041_
	);
	LUT2 #(
		.INIT('h8)
	) name19530 (
		\wishbone_bd_ram_mem1_reg[214][14]/P0001 ,
		_w12984_,
		_w30042_
	);
	LUT2 #(
		.INIT('h8)
	) name19531 (
		\wishbone_bd_ram_mem1_reg[190][14]/P0001 ,
		_w12858_,
		_w30043_
	);
	LUT2 #(
		.INIT('h8)
	) name19532 (
		\wishbone_bd_ram_mem1_reg[177][14]/P0001 ,
		_w12996_,
		_w30044_
	);
	LUT2 #(
		.INIT('h8)
	) name19533 (
		\wishbone_bd_ram_mem1_reg[217][14]/P0001 ,
		_w13188_,
		_w30045_
	);
	LUT2 #(
		.INIT('h8)
	) name19534 (
		\wishbone_bd_ram_mem1_reg[194][14]/P0001 ,
		_w12772_,
		_w30046_
	);
	LUT2 #(
		.INIT('h8)
	) name19535 (
		\wishbone_bd_ram_mem1_reg[255][14]/P0001 ,
		_w13072_,
		_w30047_
	);
	LUT2 #(
		.INIT('h8)
	) name19536 (
		\wishbone_bd_ram_mem1_reg[198][14]/P0001 ,
		_w12832_,
		_w30048_
	);
	LUT2 #(
		.INIT('h8)
	) name19537 (
		\wishbone_bd_ram_mem1_reg[137][14]/P0001 ,
		_w13168_,
		_w30049_
	);
	LUT2 #(
		.INIT('h8)
	) name19538 (
		\wishbone_bd_ram_mem1_reg[4][14]/P0001 ,
		_w12666_,
		_w30050_
	);
	LUT2 #(
		.INIT('h8)
	) name19539 (
		\wishbone_bd_ram_mem1_reg[220][14]/P0001 ,
		_w13066_,
		_w30051_
	);
	LUT2 #(
		.INIT('h8)
	) name19540 (
		\wishbone_bd_ram_mem1_reg[107][14]/P0001 ,
		_w12749_,
		_w30052_
	);
	LUT2 #(
		.INIT('h8)
	) name19541 (
		\wishbone_bd_ram_mem1_reg[95][14]/P0001 ,
		_w12844_,
		_w30053_
	);
	LUT2 #(
		.INIT('h8)
	) name19542 (
		\wishbone_bd_ram_mem1_reg[164][14]/P0001 ,
		_w12876_,
		_w30054_
	);
	LUT2 #(
		.INIT('h8)
	) name19543 (
		\wishbone_bd_ram_mem1_reg[207][14]/P0001 ,
		_w13180_,
		_w30055_
	);
	LUT2 #(
		.INIT('h8)
	) name19544 (
		\wishbone_bd_ram_mem1_reg[45][14]/P0001 ,
		_w12908_,
		_w30056_
	);
	LUT2 #(
		.INIT('h8)
	) name19545 (
		\wishbone_bd_ram_mem1_reg[202][14]/P0001 ,
		_w12870_,
		_w30057_
	);
	LUT2 #(
		.INIT('h8)
	) name19546 (
		\wishbone_bd_ram_mem1_reg[76][14]/P0001 ,
		_w13184_,
		_w30058_
	);
	LUT2 #(
		.INIT('h8)
	) name19547 (
		\wishbone_bd_ram_mem1_reg[170][14]/P0001 ,
		_w13030_,
		_w30059_
	);
	LUT2 #(
		.INIT('h8)
	) name19548 (
		\wishbone_bd_ram_mem1_reg[206][14]/P0001 ,
		_w12954_,
		_w30060_
	);
	LUT2 #(
		.INIT('h8)
	) name19549 (
		\wishbone_bd_ram_mem1_reg[140][14]/P0001 ,
		_w12894_,
		_w30061_
	);
	LUT2 #(
		.INIT('h8)
	) name19550 (
		\wishbone_bd_ram_mem1_reg[2][14]/P0001 ,
		_w13088_,
		_w30062_
	);
	LUT2 #(
		.INIT('h8)
	) name19551 (
		\wishbone_bd_ram_mem1_reg[112][14]/P0001 ,
		_w12733_,
		_w30063_
	);
	LUT2 #(
		.INIT('h8)
	) name19552 (
		\wishbone_bd_ram_mem1_reg[248][14]/P0001 ,
		_w12789_,
		_w30064_
	);
	LUT2 #(
		.INIT('h8)
	) name19553 (
		\wishbone_bd_ram_mem1_reg[126][14]/P0001 ,
		_w13218_,
		_w30065_
	);
	LUT2 #(
		.INIT('h8)
	) name19554 (
		\wishbone_bd_ram_mem1_reg[8][14]/P0001 ,
		_w12920_,
		_w30066_
	);
	LUT2 #(
		.INIT('h8)
	) name19555 (
		\wishbone_bd_ram_mem1_reg[218][14]/P0001 ,
		_w13206_,
		_w30067_
	);
	LUT2 #(
		.INIT('h8)
	) name19556 (
		\wishbone_bd_ram_mem1_reg[123][14]/P0001 ,
		_w13114_,
		_w30068_
	);
	LUT2 #(
		.INIT('h8)
	) name19557 (
		\wishbone_bd_ram_mem1_reg[189][14]/P0001 ,
		_w13042_,
		_w30069_
	);
	LUT2 #(
		.INIT('h8)
	) name19558 (
		\wishbone_bd_ram_mem1_reg[146][14]/P0001 ,
		_w13060_,
		_w30070_
	);
	LUT2 #(
		.INIT('h8)
	) name19559 (
		\wishbone_bd_ram_mem1_reg[72][14]/P0001 ,
		_w12810_,
		_w30071_
	);
	LUT2 #(
		.INIT('h8)
	) name19560 (
		\wishbone_bd_ram_mem1_reg[134][14]/P0001 ,
		_w12763_,
		_w30072_
	);
	LUT2 #(
		.INIT('h8)
	) name19561 (
		\wishbone_bd_ram_mem1_reg[54][14]/P0001 ,
		_w12770_,
		_w30073_
	);
	LUT2 #(
		.INIT('h8)
	) name19562 (
		\wishbone_bd_ram_mem1_reg[203][14]/P0001 ,
		_w13158_,
		_w30074_
	);
	LUT2 #(
		.INIT('h8)
	) name19563 (
		\wishbone_bd_ram_mem1_reg[230][14]/P0001 ,
		_w13036_,
		_w30075_
	);
	LUT2 #(
		.INIT('h8)
	) name19564 (
		\wishbone_bd_ram_mem1_reg[98][14]/P0001 ,
		_w12816_,
		_w30076_
	);
	LUT2 #(
		.INIT('h8)
	) name19565 (
		\wishbone_bd_ram_mem1_reg[172][14]/P0001 ,
		_w12944_,
		_w30077_
	);
	LUT2 #(
		.INIT('h8)
	) name19566 (
		\wishbone_bd_ram_mem1_reg[53][14]/P0001 ,
		_w13020_,
		_w30078_
	);
	LUT2 #(
		.INIT('h8)
	) name19567 (
		\wishbone_bd_ram_mem1_reg[148][14]/P0001 ,
		_w13000_,
		_w30079_
	);
	LUT2 #(
		.INIT('h8)
	) name19568 (
		\wishbone_bd_ram_mem1_reg[205][14]/P0001 ,
		_w13068_,
		_w30080_
	);
	LUT2 #(
		.INIT('h8)
	) name19569 (
		\wishbone_bd_ram_mem1_reg[12][14]/P0001 ,
		_w13118_,
		_w30081_
	);
	LUT2 #(
		.INIT('h8)
	) name19570 (
		\wishbone_bd_ram_mem1_reg[253][14]/P0001 ,
		_w13100_,
		_w30082_
	);
	LUT2 #(
		.INIT('h8)
	) name19571 (
		\wishbone_bd_ram_mem1_reg[156][14]/P0001 ,
		_w13190_,
		_w30083_
	);
	LUT2 #(
		.INIT('h8)
	) name19572 (
		\wishbone_bd_ram_mem1_reg[224][14]/P0001 ,
		_w12902_,
		_w30084_
	);
	LUT2 #(
		.INIT('h8)
	) name19573 (
		\wishbone_bd_ram_mem1_reg[41][14]/P0001 ,
		_w13052_,
		_w30085_
	);
	LUT2 #(
		.INIT('h8)
	) name19574 (
		\wishbone_bd_ram_mem1_reg[195][14]/P0001 ,
		_w13144_,
		_w30086_
	);
	LUT2 #(
		.INIT('h8)
	) name19575 (
		\wishbone_bd_ram_mem1_reg[183][14]/P0001 ,
		_w12787_,
		_w30087_
	);
	LUT2 #(
		.INIT('h8)
	) name19576 (
		\wishbone_bd_ram_mem1_reg[231][14]/P0001 ,
		_w12856_,
		_w30088_
	);
	LUT2 #(
		.INIT('h8)
	) name19577 (
		\wishbone_bd_ram_mem1_reg[221][14]/P0001 ,
		_w12802_,
		_w30089_
	);
	LUT2 #(
		.INIT('h8)
	) name19578 (
		\wishbone_bd_ram_mem1_reg[13][14]/P0001 ,
		_w13178_,
		_w30090_
	);
	LUT2 #(
		.INIT('h8)
	) name19579 (
		\wishbone_bd_ram_mem1_reg[238][14]/P0001 ,
		_w13160_,
		_w30091_
	);
	LUT2 #(
		.INIT('h8)
	) name19580 (
		\wishbone_bd_ram_mem1_reg[131][14]/P0001 ,
		_w12852_,
		_w30092_
	);
	LUT2 #(
		.INIT('h8)
	) name19581 (
		\wishbone_bd_ram_mem1_reg[73][14]/P0001 ,
		_w12918_,
		_w30093_
	);
	LUT2 #(
		.INIT('h8)
	) name19582 (
		\wishbone_bd_ram_mem1_reg[31][14]/P0001 ,
		_w13198_,
		_w30094_
	);
	LUT2 #(
		.INIT('h8)
	) name19583 (
		\wishbone_bd_ram_mem1_reg[216][14]/P0001 ,
		_w13028_,
		_w30095_
	);
	LUT2 #(
		.INIT('h8)
	) name19584 (
		\wishbone_bd_ram_mem1_reg[149][14]/P0001 ,
		_w12741_,
		_w30096_
	);
	LUT2 #(
		.INIT('h8)
	) name19585 (
		\wishbone_bd_ram_mem1_reg[35][14]/P0001 ,
		_w12703_,
		_w30097_
	);
	LUT2 #(
		.INIT('h8)
	) name19586 (
		\wishbone_bd_ram_mem1_reg[147][14]/P0001 ,
		_w13146_,
		_w30098_
	);
	LUT2 #(
		.INIT('h8)
	) name19587 (
		\wishbone_bd_ram_mem1_reg[159][14]/P0001 ,
		_w12774_,
		_w30099_
	);
	LUT2 #(
		.INIT('h8)
	) name19588 (
		\wishbone_bd_ram_mem1_reg[143][14]/P0001 ,
		_w12922_,
		_w30100_
	);
	LUT2 #(
		.INIT('h8)
	) name19589 (
		\wishbone_bd_ram_mem1_reg[154][14]/P0001 ,
		_w12962_,
		_w30101_
	);
	LUT2 #(
		.INIT('h8)
	) name19590 (
		\wishbone_bd_ram_mem1_reg[130][14]/P0001 ,
		_w12914_,
		_w30102_
	);
	LUT2 #(
		.INIT('h8)
	) name19591 (
		\wishbone_bd_ram_mem1_reg[103][14]/P0001 ,
		_w12846_,
		_w30103_
	);
	LUT2 #(
		.INIT('h8)
	) name19592 (
		\wishbone_bd_ram_mem1_reg[102][14]/P0001 ,
		_w12685_,
		_w30104_
	);
	LUT2 #(
		.INIT('h8)
	) name19593 (
		\wishbone_bd_ram_mem1_reg[141][14]/P0001 ,
		_w13004_,
		_w30105_
	);
	LUT2 #(
		.INIT('h8)
	) name19594 (
		\wishbone_bd_ram_mem1_reg[239][14]/P0001 ,
		_w12862_,
		_w30106_
	);
	LUT2 #(
		.INIT('h8)
	) name19595 (
		\wishbone_bd_ram_mem1_reg[63][14]/P0001 ,
		_w12850_,
		_w30107_
	);
	LUT2 #(
		.INIT('h8)
	) name19596 (
		\wishbone_bd_ram_mem1_reg[250][14]/P0001 ,
		_w13128_,
		_w30108_
	);
	LUT2 #(
		.INIT('h8)
	) name19597 (
		\wishbone_bd_ram_mem1_reg[79][14]/P0001 ,
		_w13212_,
		_w30109_
	);
	LUT2 #(
		.INIT('h8)
	) name19598 (
		\wishbone_bd_ram_mem1_reg[74][14]/P0001 ,
		_w12812_,
		_w30110_
	);
	LUT2 #(
		.INIT('h8)
	) name19599 (
		\wishbone_bd_ram_mem1_reg[160][14]/P0001 ,
		_w12872_,
		_w30111_
	);
	LUT2 #(
		.INIT('h8)
	) name19600 (
		\wishbone_bd_ram_mem1_reg[77][14]/P0001 ,
		_w12982_,
		_w30112_
	);
	LUT2 #(
		.INIT('h8)
	) name19601 (
		\wishbone_bd_ram_mem1_reg[22][14]/P0001 ,
		_w13110_,
		_w30113_
	);
	LUT2 #(
		.INIT('h8)
	) name19602 (
		\wishbone_bd_ram_mem1_reg[21][14]/P0001 ,
		_w12906_,
		_w30114_
	);
	LUT2 #(
		.INIT('h8)
	) name19603 (
		\wishbone_bd_ram_mem1_reg[227][14]/P0001 ,
		_w12936_,
		_w30115_
	);
	LUT2 #(
		.INIT('h8)
	) name19604 (
		\wishbone_bd_ram_mem1_reg[49][14]/P0001 ,
		_w12994_,
		_w30116_
	);
	LUT2 #(
		.INIT('h8)
	) name19605 (
		\wishbone_bd_ram_mem1_reg[184][14]/P0001 ,
		_w13062_,
		_w30117_
	);
	LUT2 #(
		.INIT('h8)
	) name19606 (
		\wishbone_bd_ram_mem1_reg[82][14]/P0001 ,
		_w12942_,
		_w30118_
	);
	LUT2 #(
		.INIT('h8)
	) name19607 (
		\wishbone_bd_ram_mem1_reg[142][14]/P0001 ,
		_w12928_,
		_w30119_
	);
	LUT2 #(
		.INIT('h8)
	) name19608 (
		\wishbone_bd_ram_mem1_reg[162][14]/P0001 ,
		_w13098_,
		_w30120_
	);
	LUT2 #(
		.INIT('h8)
	) name19609 (
		\wishbone_bd_ram_mem1_reg[37][14]/P0001 ,
		_w13102_,
		_w30121_
	);
	LUT2 #(
		.INIT('h8)
	) name19610 (
		\wishbone_bd_ram_mem1_reg[23][14]/P0001 ,
		_w13008_,
		_w30122_
	);
	LUT2 #(
		.INIT('h8)
	) name19611 (
		\wishbone_bd_ram_mem1_reg[57][14]/P0001 ,
		_w13116_,
		_w30123_
	);
	LUT2 #(
		.INIT('h8)
	) name19612 (
		\wishbone_bd_ram_mem1_reg[167][14]/P0001 ,
		_w12986_,
		_w30124_
	);
	LUT2 #(
		.INIT('h8)
	) name19613 (
		\wishbone_bd_ram_mem1_reg[226][14]/P0001 ,
		_w13138_,
		_w30125_
	);
	LUT2 #(
		.INIT('h8)
	) name19614 (
		\wishbone_bd_ram_mem1_reg[83][14]/P0001 ,
		_w12916_,
		_w30126_
	);
	LUT2 #(
		.INIT('h8)
	) name19615 (
		\wishbone_bd_ram_mem1_reg[127][14]/P0001 ,
		_w13164_,
		_w30127_
	);
	LUT2 #(
		.INIT('h8)
	) name19616 (
		\wishbone_bd_ram_mem1_reg[100][14]/P0001 ,
		_w12960_,
		_w30128_
	);
	LUT2 #(
		.INIT('h8)
	) name19617 (
		\wishbone_bd_ram_mem1_reg[60][14]/P0001 ,
		_w13204_,
		_w30129_
	);
	LUT2 #(
		.INIT('h8)
	) name19618 (
		\wishbone_bd_ram_mem1_reg[168][14]/P0001 ,
		_w13208_,
		_w30130_
	);
	LUT2 #(
		.INIT('h8)
	) name19619 (
		\wishbone_bd_ram_mem1_reg[106][14]/P0001 ,
		_w12713_,
		_w30131_
	);
	LUT2 #(
		.INIT('h8)
	) name19620 (
		\wishbone_bd_ram_mem1_reg[174][14]/P0001 ,
		_w12972_,
		_w30132_
	);
	LUT2 #(
		.INIT('h8)
	) name19621 (
		\wishbone_bd_ram_mem1_reg[244][14]/P0001 ,
		_w12747_,
		_w30133_
	);
	LUT2 #(
		.INIT('h8)
	) name19622 (
		\wishbone_bd_ram_mem1_reg[40][14]/P0001 ,
		_w13132_,
		_w30134_
	);
	LUT2 #(
		.INIT('h8)
	) name19623 (
		\wishbone_bd_ram_mem1_reg[90][14]/P0001 ,
		_w12978_,
		_w30135_
	);
	LUT2 #(
		.INIT('h8)
	) name19624 (
		\wishbone_bd_ram_mem1_reg[158][14]/P0001 ,
		_w12898_,
		_w30136_
	);
	LUT2 #(
		.INIT('h8)
	) name19625 (
		\wishbone_bd_ram_mem1_reg[59][14]/P0001 ,
		_w12780_,
		_w30137_
	);
	LUT2 #(
		.INIT('h8)
	) name19626 (
		\wishbone_bd_ram_mem1_reg[65][14]/P0001 ,
		_w13176_,
		_w30138_
	);
	LUT2 #(
		.INIT('h8)
	) name19627 (
		\wishbone_bd_ram_mem1_reg[86][14]/P0001 ,
		_w12735_,
		_w30139_
	);
	LUT2 #(
		.INIT('h8)
	) name19628 (
		\wishbone_bd_ram_mem1_reg[124][14]/P0001 ,
		_w13058_,
		_w30140_
	);
	LUT2 #(
		.INIT('h8)
	) name19629 (
		\wishbone_bd_ram_mem1_reg[181][14]/P0001 ,
		_w12828_,
		_w30141_
	);
	LUT2 #(
		.INIT('h8)
	) name19630 (
		\wishbone_bd_ram_mem1_reg[228][14]/P0001 ,
		_w12765_,
		_w30142_
	);
	LUT2 #(
		.INIT('h8)
	) name19631 (
		\wishbone_bd_ram_mem1_reg[122][14]/P0001 ,
		_w13130_,
		_w30143_
	);
	LUT2 #(
		.INIT('h8)
	) name19632 (
		\wishbone_bd_ram_mem1_reg[104][14]/P0001 ,
		_w13148_,
		_w30144_
	);
	LUT2 #(
		.INIT('h8)
	) name19633 (
		\wishbone_bd_ram_mem1_reg[99][14]/P0001 ,
		_w13038_,
		_w30145_
	);
	LUT2 #(
		.INIT('h8)
	) name19634 (
		\wishbone_bd_ram_mem1_reg[208][14]/P0001 ,
		_w13032_,
		_w30146_
	);
	LUT2 #(
		.INIT('h8)
	) name19635 (
		\wishbone_bd_ram_mem1_reg[166][14]/P0001 ,
		_w13040_,
		_w30147_
	);
	LUT2 #(
		.INIT('h8)
	) name19636 (
		\wishbone_bd_ram_mem1_reg[26][14]/P0001 ,
		_w12699_,
		_w30148_
	);
	LUT2 #(
		.INIT('h8)
	) name19637 (
		\wishbone_bd_ram_mem1_reg[9][14]/P0001 ,
		_w12808_,
		_w30149_
	);
	LUT2 #(
		.INIT('h8)
	) name19638 (
		\wishbone_bd_ram_mem1_reg[89][14]/P0001 ,
		_w12964_,
		_w30150_
	);
	LUT2 #(
		.INIT('h8)
	) name19639 (
		\wishbone_bd_ram_mem1_reg[150][14]/P0001 ,
		_w13136_,
		_w30151_
	);
	LUT2 #(
		.INIT('h8)
	) name19640 (
		\wishbone_bd_ram_mem1_reg[117][14]/P0001 ,
		_w12715_,
		_w30152_
	);
	LUT2 #(
		.INIT('h8)
	) name19641 (
		\wishbone_bd_ram_mem1_reg[67][14]/P0001 ,
		_w13134_,
		_w30153_
	);
	LUT2 #(
		.INIT('h8)
	) name19642 (
		\wishbone_bd_ram_mem1_reg[246][14]/P0001 ,
		_w13076_,
		_w30154_
	);
	LUT2 #(
		.INIT('h8)
	) name19643 (
		\wishbone_bd_ram_mem1_reg[111][14]/P0001 ,
		_w12744_,
		_w30155_
	);
	LUT2 #(
		.INIT('h8)
	) name19644 (
		\wishbone_bd_ram_mem1_reg[5][14]/P0001 ,
		_w12878_,
		_w30156_
	);
	LUT2 #(
		.INIT('h8)
	) name19645 (
		\wishbone_bd_ram_mem1_reg[229][14]/P0001 ,
		_w12711_,
		_w30157_
	);
	LUT2 #(
		.INIT('h8)
	) name19646 (
		\wishbone_bd_ram_mem1_reg[182][14]/P0001 ,
		_w12820_,
		_w30158_
	);
	LUT2 #(
		.INIT('h8)
	) name19647 (
		\wishbone_bd_ram_mem1_reg[94][14]/P0001 ,
		_w13186_,
		_w30159_
	);
	LUT2 #(
		.INIT('h8)
	) name19648 (
		\wishbone_bd_ram_mem1_reg[91][14]/P0001 ,
		_w13074_,
		_w30160_
	);
	LUT2 #(
		.INIT('h8)
	) name19649 (
		\wishbone_bd_ram_mem1_reg[71][14]/P0001 ,
		_w12798_,
		_w30161_
	);
	LUT2 #(
		.INIT('h8)
	) name19650 (
		\wishbone_bd_ram_mem1_reg[7][14]/P0001 ,
		_w12728_,
		_w30162_
	);
	LUT2 #(
		.INIT('h8)
	) name19651 (
		\wishbone_bd_ram_mem1_reg[186][14]/P0001 ,
		_w12783_,
		_w30163_
	);
	LUT2 #(
		.INIT('h8)
	) name19652 (
		\wishbone_bd_ram_mem1_reg[213][14]/P0001 ,
		_w13002_,
		_w30164_
	);
	LUT2 #(
		.INIT('h8)
	) name19653 (
		\wishbone_bd_ram_mem1_reg[144][14]/P0001 ,
		_w12756_,
		_w30165_
	);
	LUT2 #(
		.INIT('h8)
	) name19654 (
		\wishbone_bd_ram_mem1_reg[42][14]/P0001 ,
		_w12842_,
		_w30166_
	);
	LUT2 #(
		.INIT('h8)
	) name19655 (
		\wishbone_bd_ram_mem1_reg[64][14]/P0001 ,
		_w12976_,
		_w30167_
	);
	LUT2 #(
		.INIT('h8)
	) name19656 (
		\wishbone_bd_ram_mem1_reg[254][14]/P0001 ,
		_w12892_,
		_w30168_
	);
	LUT2 #(
		.INIT('h8)
	) name19657 (
		\wishbone_bd_ram_mem1_reg[139][14]/P0001 ,
		_w12814_,
		_w30169_
	);
	LUT2 #(
		.INIT('h8)
	) name19658 (
		\wishbone_bd_ram_mem1_reg[109][14]/P0001 ,
		_w12888_,
		_w30170_
	);
	LUT2 #(
		.INIT('h8)
	) name19659 (
		\wishbone_bd_ram_mem1_reg[10][14]/P0001 ,
		_w13172_,
		_w30171_
	);
	LUT2 #(
		.INIT('h8)
	) name19660 (
		\wishbone_bd_ram_mem1_reg[236][14]/P0001 ,
		_w12731_,
		_w30172_
	);
	LUT2 #(
		.INIT('h8)
	) name19661 (
		\wishbone_bd_ram_mem1_reg[96][14]/P0001 ,
		_w12912_,
		_w30173_
	);
	LUT2 #(
		.INIT('h8)
	) name19662 (
		\wishbone_bd_ram_mem1_reg[55][14]/P0001 ,
		_w12785_,
		_w30174_
	);
	LUT2 #(
		.INIT('h8)
	) name19663 (
		\wishbone_bd_ram_mem1_reg[252][14]/P0001 ,
		_w13080_,
		_w30175_
	);
	LUT2 #(
		.INIT('h8)
	) name19664 (
		\wishbone_bd_ram_mem1_reg[161][14]/P0001 ,
		_w12754_,
		_w30176_
	);
	LUT2 #(
		.INIT('h8)
	) name19665 (
		\wishbone_bd_ram_mem1_reg[153][14]/P0001 ,
		_w12890_,
		_w30177_
	);
	LUT2 #(
		.INIT('h8)
	) name19666 (
		\wishbone_bd_ram_mem1_reg[84][14]/P0001 ,
		_w12934_,
		_w30178_
	);
	LUT2 #(
		.INIT('h8)
	) name19667 (
		\wishbone_bd_ram_mem1_reg[6][14]/P0001 ,
		_w12968_,
		_w30179_
	);
	LUT2 #(
		.INIT('h8)
	) name19668 (
		\wishbone_bd_ram_mem1_reg[38][14]/P0001 ,
		_w13182_,
		_w30180_
	);
	LUT2 #(
		.INIT('h8)
	) name19669 (
		\wishbone_bd_ram_mem1_reg[119][14]/P0001 ,
		_w13048_,
		_w30181_
	);
	LUT2 #(
		.INIT('h8)
	) name19670 (
		\wishbone_bd_ram_mem1_reg[163][14]/P0001 ,
		_w12882_,
		_w30182_
	);
	LUT2 #(
		.INIT('h8)
	) name19671 (
		\wishbone_bd_ram_mem1_reg[251][14]/P0001 ,
		_w13054_,
		_w30183_
	);
	LUT2 #(
		.INIT('h8)
	) name19672 (
		\wishbone_bd_ram_mem1_reg[80][14]/P0001 ,
		_w12689_,
		_w30184_
	);
	LUT2 #(
		.INIT('h8)
	) name19673 (
		\wishbone_bd_ram_mem1_reg[34][14]/P0001 ,
		_w12930_,
		_w30185_
	);
	LUT2 #(
		.INIT('h8)
	) name19674 (
		\wishbone_bd_ram_mem1_reg[92][14]/P0001 ,
		_w13010_,
		_w30186_
	);
	LUT2 #(
		.INIT('h8)
	) name19675 (
		\wishbone_bd_ram_mem1_reg[188][14]/P0001 ,
		_w12948_,
		_w30187_
	);
	LUT2 #(
		.INIT('h8)
	) name19676 (
		\wishbone_bd_ram_mem1_reg[180][14]/P0001 ,
		_w12791_,
		_w30188_
	);
	LUT2 #(
		.INIT('h8)
	) name19677 (
		\wishbone_bd_ram_mem1_reg[173][14]/P0001 ,
		_w12854_,
		_w30189_
	);
	LUT2 #(
		.INIT('h8)
	) name19678 (
		\wishbone_bd_ram_mem1_reg[191][14]/P0001 ,
		_w13034_,
		_w30190_
	);
	LUT2 #(
		.INIT('h8)
	) name19679 (
		\wishbone_bd_ram_mem1_reg[19][14]/P0001 ,
		_w13012_,
		_w30191_
	);
	LUT2 #(
		.INIT('h8)
	) name19680 (
		\wishbone_bd_ram_mem1_reg[145][14]/P0001 ,
		_w13106_,
		_w30192_
	);
	LUT2 #(
		.INIT('h8)
	) name19681 (
		\wishbone_bd_ram_mem1_reg[192][14]/P0001 ,
		_w12938_,
		_w30193_
	);
	LUT2 #(
		.INIT('h8)
	) name19682 (
		\wishbone_bd_ram_mem1_reg[51][14]/P0001 ,
		_w13024_,
		_w30194_
	);
	LUT2 #(
		.INIT('h8)
	) name19683 (
		\wishbone_bd_ram_mem1_reg[200][14]/P0001 ,
		_w12988_,
		_w30195_
	);
	LUT2 #(
		.INIT('h8)
	) name19684 (
		\wishbone_bd_ram_mem1_reg[151][14]/P0001 ,
		_w13142_,
		_w30196_
	);
	LUT2 #(
		.INIT('h8)
	) name19685 (
		\wishbone_bd_ram_mem1_reg[39][14]/P0001 ,
		_w13018_,
		_w30197_
	);
	LUT2 #(
		.INIT('h8)
	) name19686 (
		\wishbone_bd_ram_mem1_reg[152][14]/P0001 ,
		_w12966_,
		_w30198_
	);
	LUT2 #(
		.INIT('h8)
	) name19687 (
		\wishbone_bd_ram_mem1_reg[48][14]/P0001 ,
		_w12970_,
		_w30199_
	);
	LUT2 #(
		.INIT('h8)
	) name19688 (
		\wishbone_bd_ram_mem1_reg[225][14]/P0001 ,
		_w13092_,
		_w30200_
	);
	LUT2 #(
		.INIT('h8)
	) name19689 (
		\wishbone_bd_ram_mem1_reg[3][14]/P0001 ,
		_w12866_,
		_w30201_
	);
	LUT2 #(
		.INIT('h8)
	) name19690 (
		\wishbone_bd_ram_mem1_reg[47][14]/P0001 ,
		_w12904_,
		_w30202_
	);
	LUT2 #(
		.INIT('h8)
	) name19691 (
		\wishbone_bd_ram_mem1_reg[120][14]/P0001 ,
		_w12707_,
		_w30203_
	);
	LUT2 #(
		.INIT('h8)
	) name19692 (
		\wishbone_bd_ram_mem1_reg[187][14]/P0001 ,
		_w13196_,
		_w30204_
	);
	LUT2 #(
		.INIT('h8)
	) name19693 (
		\wishbone_bd_ram_mem1_reg[20][14]/P0001 ,
		_w13174_,
		_w30205_
	);
	LUT2 #(
		.INIT('h8)
	) name19694 (
		\wishbone_bd_ram_mem1_reg[136][14]/P0001 ,
		_w13064_,
		_w30206_
	);
	LUT2 #(
		.INIT('h8)
	) name19695 (
		\wishbone_bd_ram_mem1_reg[110][14]/P0001 ,
		_w13046_,
		_w30207_
	);
	LUT2 #(
		.INIT('h8)
	) name19696 (
		\wishbone_bd_ram_mem1_reg[201][14]/P0001 ,
		_w12822_,
		_w30208_
	);
	LUT2 #(
		.INIT('h8)
	) name19697 (
		\wishbone_bd_ram_mem1_reg[61][14]/P0001 ,
		_w12725_,
		_w30209_
	);
	LUT2 #(
		.INIT('h8)
	) name19698 (
		\wishbone_bd_ram_mem1_reg[245][14]/P0001 ,
		_w13022_,
		_w30210_
	);
	LUT2 #(
		.INIT('h8)
	) name19699 (
		\wishbone_bd_ram_mem1_reg[193][14]/P0001 ,
		_w13056_,
		_w30211_
	);
	LUT2 #(
		.INIT('h8)
	) name19700 (
		\wishbone_bd_ram_mem1_reg[249][14]/P0001 ,
		_w12900_,
		_w30212_
	);
	LUT2 #(
		.INIT('h8)
	) name19701 (
		\wishbone_bd_ram_mem1_reg[15][14]/P0001 ,
		_w13210_,
		_w30213_
	);
	LUT2 #(
		.INIT('h8)
	) name19702 (
		\wishbone_bd_ram_mem1_reg[52][14]/P0001 ,
		_w13082_,
		_w30214_
	);
	LUT2 #(
		.INIT('h8)
	) name19703 (
		\wishbone_bd_ram_mem1_reg[179][14]/P0001 ,
		_w13050_,
		_w30215_
	);
	LUT2 #(
		.INIT('h8)
	) name19704 (
		\wishbone_bd_ram_mem1_reg[24][14]/P0001 ,
		_w13084_,
		_w30216_
	);
	LUT2 #(
		.INIT('h8)
	) name19705 (
		\wishbone_bd_ram_mem1_reg[88][14]/P0001 ,
		_w12860_,
		_w30217_
	);
	LUT2 #(
		.INIT('h8)
	) name19706 (
		\wishbone_bd_ram_mem1_reg[115][14]/P0001 ,
		_w13112_,
		_w30218_
	);
	LUT2 #(
		.INIT('h8)
	) name19707 (
		\wishbone_bd_ram_mem1_reg[97][14]/P0001 ,
		_w13096_,
		_w30219_
	);
	LUT2 #(
		.INIT('h8)
	) name19708 (
		\wishbone_bd_ram_mem1_reg[62][14]/P0001 ,
		_w12673_,
		_w30220_
	);
	LUT2 #(
		.INIT('h8)
	) name19709 (
		\wishbone_bd_ram_mem1_reg[196][14]/P0001 ,
		_w13090_,
		_w30221_
	);
	LUT2 #(
		.INIT('h8)
	) name19710 (
		\wishbone_bd_ram_mem1_reg[30][14]/P0001 ,
		_w13104_,
		_w30222_
	);
	LUT2 #(
		.INIT('h8)
	) name19711 (
		\wishbone_bd_ram_mem1_reg[128][14]/P0001 ,
		_w12793_,
		_w30223_
	);
	LUT2 #(
		.INIT('h1)
	) name19712 (
		_w29968_,
		_w29969_,
		_w30224_
	);
	LUT2 #(
		.INIT('h1)
	) name19713 (
		_w29970_,
		_w29971_,
		_w30225_
	);
	LUT2 #(
		.INIT('h1)
	) name19714 (
		_w29972_,
		_w29973_,
		_w30226_
	);
	LUT2 #(
		.INIT('h1)
	) name19715 (
		_w29974_,
		_w29975_,
		_w30227_
	);
	LUT2 #(
		.INIT('h1)
	) name19716 (
		_w29976_,
		_w29977_,
		_w30228_
	);
	LUT2 #(
		.INIT('h1)
	) name19717 (
		_w29978_,
		_w29979_,
		_w30229_
	);
	LUT2 #(
		.INIT('h1)
	) name19718 (
		_w29980_,
		_w29981_,
		_w30230_
	);
	LUT2 #(
		.INIT('h1)
	) name19719 (
		_w29982_,
		_w29983_,
		_w30231_
	);
	LUT2 #(
		.INIT('h1)
	) name19720 (
		_w29984_,
		_w29985_,
		_w30232_
	);
	LUT2 #(
		.INIT('h1)
	) name19721 (
		_w29986_,
		_w29987_,
		_w30233_
	);
	LUT2 #(
		.INIT('h1)
	) name19722 (
		_w29988_,
		_w29989_,
		_w30234_
	);
	LUT2 #(
		.INIT('h1)
	) name19723 (
		_w29990_,
		_w29991_,
		_w30235_
	);
	LUT2 #(
		.INIT('h1)
	) name19724 (
		_w29992_,
		_w29993_,
		_w30236_
	);
	LUT2 #(
		.INIT('h1)
	) name19725 (
		_w29994_,
		_w29995_,
		_w30237_
	);
	LUT2 #(
		.INIT('h1)
	) name19726 (
		_w29996_,
		_w29997_,
		_w30238_
	);
	LUT2 #(
		.INIT('h1)
	) name19727 (
		_w29998_,
		_w29999_,
		_w30239_
	);
	LUT2 #(
		.INIT('h1)
	) name19728 (
		_w30000_,
		_w30001_,
		_w30240_
	);
	LUT2 #(
		.INIT('h1)
	) name19729 (
		_w30002_,
		_w30003_,
		_w30241_
	);
	LUT2 #(
		.INIT('h1)
	) name19730 (
		_w30004_,
		_w30005_,
		_w30242_
	);
	LUT2 #(
		.INIT('h1)
	) name19731 (
		_w30006_,
		_w30007_,
		_w30243_
	);
	LUT2 #(
		.INIT('h1)
	) name19732 (
		_w30008_,
		_w30009_,
		_w30244_
	);
	LUT2 #(
		.INIT('h1)
	) name19733 (
		_w30010_,
		_w30011_,
		_w30245_
	);
	LUT2 #(
		.INIT('h1)
	) name19734 (
		_w30012_,
		_w30013_,
		_w30246_
	);
	LUT2 #(
		.INIT('h1)
	) name19735 (
		_w30014_,
		_w30015_,
		_w30247_
	);
	LUT2 #(
		.INIT('h1)
	) name19736 (
		_w30016_,
		_w30017_,
		_w30248_
	);
	LUT2 #(
		.INIT('h1)
	) name19737 (
		_w30018_,
		_w30019_,
		_w30249_
	);
	LUT2 #(
		.INIT('h1)
	) name19738 (
		_w30020_,
		_w30021_,
		_w30250_
	);
	LUT2 #(
		.INIT('h1)
	) name19739 (
		_w30022_,
		_w30023_,
		_w30251_
	);
	LUT2 #(
		.INIT('h1)
	) name19740 (
		_w30024_,
		_w30025_,
		_w30252_
	);
	LUT2 #(
		.INIT('h1)
	) name19741 (
		_w30026_,
		_w30027_,
		_w30253_
	);
	LUT2 #(
		.INIT('h1)
	) name19742 (
		_w30028_,
		_w30029_,
		_w30254_
	);
	LUT2 #(
		.INIT('h1)
	) name19743 (
		_w30030_,
		_w30031_,
		_w30255_
	);
	LUT2 #(
		.INIT('h1)
	) name19744 (
		_w30032_,
		_w30033_,
		_w30256_
	);
	LUT2 #(
		.INIT('h1)
	) name19745 (
		_w30034_,
		_w30035_,
		_w30257_
	);
	LUT2 #(
		.INIT('h1)
	) name19746 (
		_w30036_,
		_w30037_,
		_w30258_
	);
	LUT2 #(
		.INIT('h1)
	) name19747 (
		_w30038_,
		_w30039_,
		_w30259_
	);
	LUT2 #(
		.INIT('h1)
	) name19748 (
		_w30040_,
		_w30041_,
		_w30260_
	);
	LUT2 #(
		.INIT('h1)
	) name19749 (
		_w30042_,
		_w30043_,
		_w30261_
	);
	LUT2 #(
		.INIT('h1)
	) name19750 (
		_w30044_,
		_w30045_,
		_w30262_
	);
	LUT2 #(
		.INIT('h1)
	) name19751 (
		_w30046_,
		_w30047_,
		_w30263_
	);
	LUT2 #(
		.INIT('h1)
	) name19752 (
		_w30048_,
		_w30049_,
		_w30264_
	);
	LUT2 #(
		.INIT('h1)
	) name19753 (
		_w30050_,
		_w30051_,
		_w30265_
	);
	LUT2 #(
		.INIT('h1)
	) name19754 (
		_w30052_,
		_w30053_,
		_w30266_
	);
	LUT2 #(
		.INIT('h1)
	) name19755 (
		_w30054_,
		_w30055_,
		_w30267_
	);
	LUT2 #(
		.INIT('h1)
	) name19756 (
		_w30056_,
		_w30057_,
		_w30268_
	);
	LUT2 #(
		.INIT('h1)
	) name19757 (
		_w30058_,
		_w30059_,
		_w30269_
	);
	LUT2 #(
		.INIT('h1)
	) name19758 (
		_w30060_,
		_w30061_,
		_w30270_
	);
	LUT2 #(
		.INIT('h1)
	) name19759 (
		_w30062_,
		_w30063_,
		_w30271_
	);
	LUT2 #(
		.INIT('h1)
	) name19760 (
		_w30064_,
		_w30065_,
		_w30272_
	);
	LUT2 #(
		.INIT('h1)
	) name19761 (
		_w30066_,
		_w30067_,
		_w30273_
	);
	LUT2 #(
		.INIT('h1)
	) name19762 (
		_w30068_,
		_w30069_,
		_w30274_
	);
	LUT2 #(
		.INIT('h1)
	) name19763 (
		_w30070_,
		_w30071_,
		_w30275_
	);
	LUT2 #(
		.INIT('h1)
	) name19764 (
		_w30072_,
		_w30073_,
		_w30276_
	);
	LUT2 #(
		.INIT('h1)
	) name19765 (
		_w30074_,
		_w30075_,
		_w30277_
	);
	LUT2 #(
		.INIT('h1)
	) name19766 (
		_w30076_,
		_w30077_,
		_w30278_
	);
	LUT2 #(
		.INIT('h1)
	) name19767 (
		_w30078_,
		_w30079_,
		_w30279_
	);
	LUT2 #(
		.INIT('h1)
	) name19768 (
		_w30080_,
		_w30081_,
		_w30280_
	);
	LUT2 #(
		.INIT('h1)
	) name19769 (
		_w30082_,
		_w30083_,
		_w30281_
	);
	LUT2 #(
		.INIT('h1)
	) name19770 (
		_w30084_,
		_w30085_,
		_w30282_
	);
	LUT2 #(
		.INIT('h1)
	) name19771 (
		_w30086_,
		_w30087_,
		_w30283_
	);
	LUT2 #(
		.INIT('h1)
	) name19772 (
		_w30088_,
		_w30089_,
		_w30284_
	);
	LUT2 #(
		.INIT('h1)
	) name19773 (
		_w30090_,
		_w30091_,
		_w30285_
	);
	LUT2 #(
		.INIT('h1)
	) name19774 (
		_w30092_,
		_w30093_,
		_w30286_
	);
	LUT2 #(
		.INIT('h1)
	) name19775 (
		_w30094_,
		_w30095_,
		_w30287_
	);
	LUT2 #(
		.INIT('h1)
	) name19776 (
		_w30096_,
		_w30097_,
		_w30288_
	);
	LUT2 #(
		.INIT('h1)
	) name19777 (
		_w30098_,
		_w30099_,
		_w30289_
	);
	LUT2 #(
		.INIT('h1)
	) name19778 (
		_w30100_,
		_w30101_,
		_w30290_
	);
	LUT2 #(
		.INIT('h1)
	) name19779 (
		_w30102_,
		_w30103_,
		_w30291_
	);
	LUT2 #(
		.INIT('h1)
	) name19780 (
		_w30104_,
		_w30105_,
		_w30292_
	);
	LUT2 #(
		.INIT('h1)
	) name19781 (
		_w30106_,
		_w30107_,
		_w30293_
	);
	LUT2 #(
		.INIT('h1)
	) name19782 (
		_w30108_,
		_w30109_,
		_w30294_
	);
	LUT2 #(
		.INIT('h1)
	) name19783 (
		_w30110_,
		_w30111_,
		_w30295_
	);
	LUT2 #(
		.INIT('h1)
	) name19784 (
		_w30112_,
		_w30113_,
		_w30296_
	);
	LUT2 #(
		.INIT('h1)
	) name19785 (
		_w30114_,
		_w30115_,
		_w30297_
	);
	LUT2 #(
		.INIT('h1)
	) name19786 (
		_w30116_,
		_w30117_,
		_w30298_
	);
	LUT2 #(
		.INIT('h1)
	) name19787 (
		_w30118_,
		_w30119_,
		_w30299_
	);
	LUT2 #(
		.INIT('h1)
	) name19788 (
		_w30120_,
		_w30121_,
		_w30300_
	);
	LUT2 #(
		.INIT('h1)
	) name19789 (
		_w30122_,
		_w30123_,
		_w30301_
	);
	LUT2 #(
		.INIT('h1)
	) name19790 (
		_w30124_,
		_w30125_,
		_w30302_
	);
	LUT2 #(
		.INIT('h1)
	) name19791 (
		_w30126_,
		_w30127_,
		_w30303_
	);
	LUT2 #(
		.INIT('h1)
	) name19792 (
		_w30128_,
		_w30129_,
		_w30304_
	);
	LUT2 #(
		.INIT('h1)
	) name19793 (
		_w30130_,
		_w30131_,
		_w30305_
	);
	LUT2 #(
		.INIT('h1)
	) name19794 (
		_w30132_,
		_w30133_,
		_w30306_
	);
	LUT2 #(
		.INIT('h1)
	) name19795 (
		_w30134_,
		_w30135_,
		_w30307_
	);
	LUT2 #(
		.INIT('h1)
	) name19796 (
		_w30136_,
		_w30137_,
		_w30308_
	);
	LUT2 #(
		.INIT('h1)
	) name19797 (
		_w30138_,
		_w30139_,
		_w30309_
	);
	LUT2 #(
		.INIT('h1)
	) name19798 (
		_w30140_,
		_w30141_,
		_w30310_
	);
	LUT2 #(
		.INIT('h1)
	) name19799 (
		_w30142_,
		_w30143_,
		_w30311_
	);
	LUT2 #(
		.INIT('h1)
	) name19800 (
		_w30144_,
		_w30145_,
		_w30312_
	);
	LUT2 #(
		.INIT('h1)
	) name19801 (
		_w30146_,
		_w30147_,
		_w30313_
	);
	LUT2 #(
		.INIT('h1)
	) name19802 (
		_w30148_,
		_w30149_,
		_w30314_
	);
	LUT2 #(
		.INIT('h1)
	) name19803 (
		_w30150_,
		_w30151_,
		_w30315_
	);
	LUT2 #(
		.INIT('h1)
	) name19804 (
		_w30152_,
		_w30153_,
		_w30316_
	);
	LUT2 #(
		.INIT('h1)
	) name19805 (
		_w30154_,
		_w30155_,
		_w30317_
	);
	LUT2 #(
		.INIT('h1)
	) name19806 (
		_w30156_,
		_w30157_,
		_w30318_
	);
	LUT2 #(
		.INIT('h1)
	) name19807 (
		_w30158_,
		_w30159_,
		_w30319_
	);
	LUT2 #(
		.INIT('h1)
	) name19808 (
		_w30160_,
		_w30161_,
		_w30320_
	);
	LUT2 #(
		.INIT('h1)
	) name19809 (
		_w30162_,
		_w30163_,
		_w30321_
	);
	LUT2 #(
		.INIT('h1)
	) name19810 (
		_w30164_,
		_w30165_,
		_w30322_
	);
	LUT2 #(
		.INIT('h1)
	) name19811 (
		_w30166_,
		_w30167_,
		_w30323_
	);
	LUT2 #(
		.INIT('h1)
	) name19812 (
		_w30168_,
		_w30169_,
		_w30324_
	);
	LUT2 #(
		.INIT('h1)
	) name19813 (
		_w30170_,
		_w30171_,
		_w30325_
	);
	LUT2 #(
		.INIT('h1)
	) name19814 (
		_w30172_,
		_w30173_,
		_w30326_
	);
	LUT2 #(
		.INIT('h1)
	) name19815 (
		_w30174_,
		_w30175_,
		_w30327_
	);
	LUT2 #(
		.INIT('h1)
	) name19816 (
		_w30176_,
		_w30177_,
		_w30328_
	);
	LUT2 #(
		.INIT('h1)
	) name19817 (
		_w30178_,
		_w30179_,
		_w30329_
	);
	LUT2 #(
		.INIT('h1)
	) name19818 (
		_w30180_,
		_w30181_,
		_w30330_
	);
	LUT2 #(
		.INIT('h1)
	) name19819 (
		_w30182_,
		_w30183_,
		_w30331_
	);
	LUT2 #(
		.INIT('h1)
	) name19820 (
		_w30184_,
		_w30185_,
		_w30332_
	);
	LUT2 #(
		.INIT('h1)
	) name19821 (
		_w30186_,
		_w30187_,
		_w30333_
	);
	LUT2 #(
		.INIT('h1)
	) name19822 (
		_w30188_,
		_w30189_,
		_w30334_
	);
	LUT2 #(
		.INIT('h1)
	) name19823 (
		_w30190_,
		_w30191_,
		_w30335_
	);
	LUT2 #(
		.INIT('h1)
	) name19824 (
		_w30192_,
		_w30193_,
		_w30336_
	);
	LUT2 #(
		.INIT('h1)
	) name19825 (
		_w30194_,
		_w30195_,
		_w30337_
	);
	LUT2 #(
		.INIT('h1)
	) name19826 (
		_w30196_,
		_w30197_,
		_w30338_
	);
	LUT2 #(
		.INIT('h1)
	) name19827 (
		_w30198_,
		_w30199_,
		_w30339_
	);
	LUT2 #(
		.INIT('h1)
	) name19828 (
		_w30200_,
		_w30201_,
		_w30340_
	);
	LUT2 #(
		.INIT('h1)
	) name19829 (
		_w30202_,
		_w30203_,
		_w30341_
	);
	LUT2 #(
		.INIT('h1)
	) name19830 (
		_w30204_,
		_w30205_,
		_w30342_
	);
	LUT2 #(
		.INIT('h1)
	) name19831 (
		_w30206_,
		_w30207_,
		_w30343_
	);
	LUT2 #(
		.INIT('h1)
	) name19832 (
		_w30208_,
		_w30209_,
		_w30344_
	);
	LUT2 #(
		.INIT('h1)
	) name19833 (
		_w30210_,
		_w30211_,
		_w30345_
	);
	LUT2 #(
		.INIT('h1)
	) name19834 (
		_w30212_,
		_w30213_,
		_w30346_
	);
	LUT2 #(
		.INIT('h1)
	) name19835 (
		_w30214_,
		_w30215_,
		_w30347_
	);
	LUT2 #(
		.INIT('h1)
	) name19836 (
		_w30216_,
		_w30217_,
		_w30348_
	);
	LUT2 #(
		.INIT('h1)
	) name19837 (
		_w30218_,
		_w30219_,
		_w30349_
	);
	LUT2 #(
		.INIT('h1)
	) name19838 (
		_w30220_,
		_w30221_,
		_w30350_
	);
	LUT2 #(
		.INIT('h1)
	) name19839 (
		_w30222_,
		_w30223_,
		_w30351_
	);
	LUT2 #(
		.INIT('h8)
	) name19840 (
		_w30350_,
		_w30351_,
		_w30352_
	);
	LUT2 #(
		.INIT('h8)
	) name19841 (
		_w30348_,
		_w30349_,
		_w30353_
	);
	LUT2 #(
		.INIT('h8)
	) name19842 (
		_w30346_,
		_w30347_,
		_w30354_
	);
	LUT2 #(
		.INIT('h8)
	) name19843 (
		_w30344_,
		_w30345_,
		_w30355_
	);
	LUT2 #(
		.INIT('h8)
	) name19844 (
		_w30342_,
		_w30343_,
		_w30356_
	);
	LUT2 #(
		.INIT('h8)
	) name19845 (
		_w30340_,
		_w30341_,
		_w30357_
	);
	LUT2 #(
		.INIT('h8)
	) name19846 (
		_w30338_,
		_w30339_,
		_w30358_
	);
	LUT2 #(
		.INIT('h8)
	) name19847 (
		_w30336_,
		_w30337_,
		_w30359_
	);
	LUT2 #(
		.INIT('h8)
	) name19848 (
		_w30334_,
		_w30335_,
		_w30360_
	);
	LUT2 #(
		.INIT('h8)
	) name19849 (
		_w30332_,
		_w30333_,
		_w30361_
	);
	LUT2 #(
		.INIT('h8)
	) name19850 (
		_w30330_,
		_w30331_,
		_w30362_
	);
	LUT2 #(
		.INIT('h8)
	) name19851 (
		_w30328_,
		_w30329_,
		_w30363_
	);
	LUT2 #(
		.INIT('h8)
	) name19852 (
		_w30326_,
		_w30327_,
		_w30364_
	);
	LUT2 #(
		.INIT('h8)
	) name19853 (
		_w30324_,
		_w30325_,
		_w30365_
	);
	LUT2 #(
		.INIT('h8)
	) name19854 (
		_w30322_,
		_w30323_,
		_w30366_
	);
	LUT2 #(
		.INIT('h8)
	) name19855 (
		_w30320_,
		_w30321_,
		_w30367_
	);
	LUT2 #(
		.INIT('h8)
	) name19856 (
		_w30318_,
		_w30319_,
		_w30368_
	);
	LUT2 #(
		.INIT('h8)
	) name19857 (
		_w30316_,
		_w30317_,
		_w30369_
	);
	LUT2 #(
		.INIT('h8)
	) name19858 (
		_w30314_,
		_w30315_,
		_w30370_
	);
	LUT2 #(
		.INIT('h8)
	) name19859 (
		_w30312_,
		_w30313_,
		_w30371_
	);
	LUT2 #(
		.INIT('h8)
	) name19860 (
		_w30310_,
		_w30311_,
		_w30372_
	);
	LUT2 #(
		.INIT('h8)
	) name19861 (
		_w30308_,
		_w30309_,
		_w30373_
	);
	LUT2 #(
		.INIT('h8)
	) name19862 (
		_w30306_,
		_w30307_,
		_w30374_
	);
	LUT2 #(
		.INIT('h8)
	) name19863 (
		_w30304_,
		_w30305_,
		_w30375_
	);
	LUT2 #(
		.INIT('h8)
	) name19864 (
		_w30302_,
		_w30303_,
		_w30376_
	);
	LUT2 #(
		.INIT('h8)
	) name19865 (
		_w30300_,
		_w30301_,
		_w30377_
	);
	LUT2 #(
		.INIT('h8)
	) name19866 (
		_w30298_,
		_w30299_,
		_w30378_
	);
	LUT2 #(
		.INIT('h8)
	) name19867 (
		_w30296_,
		_w30297_,
		_w30379_
	);
	LUT2 #(
		.INIT('h8)
	) name19868 (
		_w30294_,
		_w30295_,
		_w30380_
	);
	LUT2 #(
		.INIT('h8)
	) name19869 (
		_w30292_,
		_w30293_,
		_w30381_
	);
	LUT2 #(
		.INIT('h8)
	) name19870 (
		_w30290_,
		_w30291_,
		_w30382_
	);
	LUT2 #(
		.INIT('h8)
	) name19871 (
		_w30288_,
		_w30289_,
		_w30383_
	);
	LUT2 #(
		.INIT('h8)
	) name19872 (
		_w30286_,
		_w30287_,
		_w30384_
	);
	LUT2 #(
		.INIT('h8)
	) name19873 (
		_w30284_,
		_w30285_,
		_w30385_
	);
	LUT2 #(
		.INIT('h8)
	) name19874 (
		_w30282_,
		_w30283_,
		_w30386_
	);
	LUT2 #(
		.INIT('h8)
	) name19875 (
		_w30280_,
		_w30281_,
		_w30387_
	);
	LUT2 #(
		.INIT('h8)
	) name19876 (
		_w30278_,
		_w30279_,
		_w30388_
	);
	LUT2 #(
		.INIT('h8)
	) name19877 (
		_w30276_,
		_w30277_,
		_w30389_
	);
	LUT2 #(
		.INIT('h8)
	) name19878 (
		_w30274_,
		_w30275_,
		_w30390_
	);
	LUT2 #(
		.INIT('h8)
	) name19879 (
		_w30272_,
		_w30273_,
		_w30391_
	);
	LUT2 #(
		.INIT('h8)
	) name19880 (
		_w30270_,
		_w30271_,
		_w30392_
	);
	LUT2 #(
		.INIT('h8)
	) name19881 (
		_w30268_,
		_w30269_,
		_w30393_
	);
	LUT2 #(
		.INIT('h8)
	) name19882 (
		_w30266_,
		_w30267_,
		_w30394_
	);
	LUT2 #(
		.INIT('h8)
	) name19883 (
		_w30264_,
		_w30265_,
		_w30395_
	);
	LUT2 #(
		.INIT('h8)
	) name19884 (
		_w30262_,
		_w30263_,
		_w30396_
	);
	LUT2 #(
		.INIT('h8)
	) name19885 (
		_w30260_,
		_w30261_,
		_w30397_
	);
	LUT2 #(
		.INIT('h8)
	) name19886 (
		_w30258_,
		_w30259_,
		_w30398_
	);
	LUT2 #(
		.INIT('h8)
	) name19887 (
		_w30256_,
		_w30257_,
		_w30399_
	);
	LUT2 #(
		.INIT('h8)
	) name19888 (
		_w30254_,
		_w30255_,
		_w30400_
	);
	LUT2 #(
		.INIT('h8)
	) name19889 (
		_w30252_,
		_w30253_,
		_w30401_
	);
	LUT2 #(
		.INIT('h8)
	) name19890 (
		_w30250_,
		_w30251_,
		_w30402_
	);
	LUT2 #(
		.INIT('h8)
	) name19891 (
		_w30248_,
		_w30249_,
		_w30403_
	);
	LUT2 #(
		.INIT('h8)
	) name19892 (
		_w30246_,
		_w30247_,
		_w30404_
	);
	LUT2 #(
		.INIT('h8)
	) name19893 (
		_w30244_,
		_w30245_,
		_w30405_
	);
	LUT2 #(
		.INIT('h8)
	) name19894 (
		_w30242_,
		_w30243_,
		_w30406_
	);
	LUT2 #(
		.INIT('h8)
	) name19895 (
		_w30240_,
		_w30241_,
		_w30407_
	);
	LUT2 #(
		.INIT('h8)
	) name19896 (
		_w30238_,
		_w30239_,
		_w30408_
	);
	LUT2 #(
		.INIT('h8)
	) name19897 (
		_w30236_,
		_w30237_,
		_w30409_
	);
	LUT2 #(
		.INIT('h8)
	) name19898 (
		_w30234_,
		_w30235_,
		_w30410_
	);
	LUT2 #(
		.INIT('h8)
	) name19899 (
		_w30232_,
		_w30233_,
		_w30411_
	);
	LUT2 #(
		.INIT('h8)
	) name19900 (
		_w30230_,
		_w30231_,
		_w30412_
	);
	LUT2 #(
		.INIT('h8)
	) name19901 (
		_w30228_,
		_w30229_,
		_w30413_
	);
	LUT2 #(
		.INIT('h8)
	) name19902 (
		_w30226_,
		_w30227_,
		_w30414_
	);
	LUT2 #(
		.INIT('h8)
	) name19903 (
		_w30224_,
		_w30225_,
		_w30415_
	);
	LUT2 #(
		.INIT('h8)
	) name19904 (
		_w30414_,
		_w30415_,
		_w30416_
	);
	LUT2 #(
		.INIT('h8)
	) name19905 (
		_w30412_,
		_w30413_,
		_w30417_
	);
	LUT2 #(
		.INIT('h8)
	) name19906 (
		_w30410_,
		_w30411_,
		_w30418_
	);
	LUT2 #(
		.INIT('h8)
	) name19907 (
		_w30408_,
		_w30409_,
		_w30419_
	);
	LUT2 #(
		.INIT('h8)
	) name19908 (
		_w30406_,
		_w30407_,
		_w30420_
	);
	LUT2 #(
		.INIT('h8)
	) name19909 (
		_w30404_,
		_w30405_,
		_w30421_
	);
	LUT2 #(
		.INIT('h8)
	) name19910 (
		_w30402_,
		_w30403_,
		_w30422_
	);
	LUT2 #(
		.INIT('h8)
	) name19911 (
		_w30400_,
		_w30401_,
		_w30423_
	);
	LUT2 #(
		.INIT('h8)
	) name19912 (
		_w30398_,
		_w30399_,
		_w30424_
	);
	LUT2 #(
		.INIT('h8)
	) name19913 (
		_w30396_,
		_w30397_,
		_w30425_
	);
	LUT2 #(
		.INIT('h8)
	) name19914 (
		_w30394_,
		_w30395_,
		_w30426_
	);
	LUT2 #(
		.INIT('h8)
	) name19915 (
		_w30392_,
		_w30393_,
		_w30427_
	);
	LUT2 #(
		.INIT('h8)
	) name19916 (
		_w30390_,
		_w30391_,
		_w30428_
	);
	LUT2 #(
		.INIT('h8)
	) name19917 (
		_w30388_,
		_w30389_,
		_w30429_
	);
	LUT2 #(
		.INIT('h8)
	) name19918 (
		_w30386_,
		_w30387_,
		_w30430_
	);
	LUT2 #(
		.INIT('h8)
	) name19919 (
		_w30384_,
		_w30385_,
		_w30431_
	);
	LUT2 #(
		.INIT('h8)
	) name19920 (
		_w30382_,
		_w30383_,
		_w30432_
	);
	LUT2 #(
		.INIT('h8)
	) name19921 (
		_w30380_,
		_w30381_,
		_w30433_
	);
	LUT2 #(
		.INIT('h8)
	) name19922 (
		_w30378_,
		_w30379_,
		_w30434_
	);
	LUT2 #(
		.INIT('h8)
	) name19923 (
		_w30376_,
		_w30377_,
		_w30435_
	);
	LUT2 #(
		.INIT('h8)
	) name19924 (
		_w30374_,
		_w30375_,
		_w30436_
	);
	LUT2 #(
		.INIT('h8)
	) name19925 (
		_w30372_,
		_w30373_,
		_w30437_
	);
	LUT2 #(
		.INIT('h8)
	) name19926 (
		_w30370_,
		_w30371_,
		_w30438_
	);
	LUT2 #(
		.INIT('h8)
	) name19927 (
		_w30368_,
		_w30369_,
		_w30439_
	);
	LUT2 #(
		.INIT('h8)
	) name19928 (
		_w30366_,
		_w30367_,
		_w30440_
	);
	LUT2 #(
		.INIT('h8)
	) name19929 (
		_w30364_,
		_w30365_,
		_w30441_
	);
	LUT2 #(
		.INIT('h8)
	) name19930 (
		_w30362_,
		_w30363_,
		_w30442_
	);
	LUT2 #(
		.INIT('h8)
	) name19931 (
		_w30360_,
		_w30361_,
		_w30443_
	);
	LUT2 #(
		.INIT('h8)
	) name19932 (
		_w30358_,
		_w30359_,
		_w30444_
	);
	LUT2 #(
		.INIT('h8)
	) name19933 (
		_w30356_,
		_w30357_,
		_w30445_
	);
	LUT2 #(
		.INIT('h8)
	) name19934 (
		_w30354_,
		_w30355_,
		_w30446_
	);
	LUT2 #(
		.INIT('h8)
	) name19935 (
		_w30352_,
		_w30353_,
		_w30447_
	);
	LUT2 #(
		.INIT('h8)
	) name19936 (
		_w30446_,
		_w30447_,
		_w30448_
	);
	LUT2 #(
		.INIT('h8)
	) name19937 (
		_w30444_,
		_w30445_,
		_w30449_
	);
	LUT2 #(
		.INIT('h8)
	) name19938 (
		_w30442_,
		_w30443_,
		_w30450_
	);
	LUT2 #(
		.INIT('h8)
	) name19939 (
		_w30440_,
		_w30441_,
		_w30451_
	);
	LUT2 #(
		.INIT('h8)
	) name19940 (
		_w30438_,
		_w30439_,
		_w30452_
	);
	LUT2 #(
		.INIT('h8)
	) name19941 (
		_w30436_,
		_w30437_,
		_w30453_
	);
	LUT2 #(
		.INIT('h8)
	) name19942 (
		_w30434_,
		_w30435_,
		_w30454_
	);
	LUT2 #(
		.INIT('h8)
	) name19943 (
		_w30432_,
		_w30433_,
		_w30455_
	);
	LUT2 #(
		.INIT('h8)
	) name19944 (
		_w30430_,
		_w30431_,
		_w30456_
	);
	LUT2 #(
		.INIT('h8)
	) name19945 (
		_w30428_,
		_w30429_,
		_w30457_
	);
	LUT2 #(
		.INIT('h8)
	) name19946 (
		_w30426_,
		_w30427_,
		_w30458_
	);
	LUT2 #(
		.INIT('h8)
	) name19947 (
		_w30424_,
		_w30425_,
		_w30459_
	);
	LUT2 #(
		.INIT('h8)
	) name19948 (
		_w30422_,
		_w30423_,
		_w30460_
	);
	LUT2 #(
		.INIT('h8)
	) name19949 (
		_w30420_,
		_w30421_,
		_w30461_
	);
	LUT2 #(
		.INIT('h8)
	) name19950 (
		_w30418_,
		_w30419_,
		_w30462_
	);
	LUT2 #(
		.INIT('h8)
	) name19951 (
		_w30416_,
		_w30417_,
		_w30463_
	);
	LUT2 #(
		.INIT('h8)
	) name19952 (
		_w30462_,
		_w30463_,
		_w30464_
	);
	LUT2 #(
		.INIT('h8)
	) name19953 (
		_w30460_,
		_w30461_,
		_w30465_
	);
	LUT2 #(
		.INIT('h8)
	) name19954 (
		_w30458_,
		_w30459_,
		_w30466_
	);
	LUT2 #(
		.INIT('h8)
	) name19955 (
		_w30456_,
		_w30457_,
		_w30467_
	);
	LUT2 #(
		.INIT('h8)
	) name19956 (
		_w30454_,
		_w30455_,
		_w30468_
	);
	LUT2 #(
		.INIT('h8)
	) name19957 (
		_w30452_,
		_w30453_,
		_w30469_
	);
	LUT2 #(
		.INIT('h8)
	) name19958 (
		_w30450_,
		_w30451_,
		_w30470_
	);
	LUT2 #(
		.INIT('h8)
	) name19959 (
		_w30448_,
		_w30449_,
		_w30471_
	);
	LUT2 #(
		.INIT('h8)
	) name19960 (
		_w30470_,
		_w30471_,
		_w30472_
	);
	LUT2 #(
		.INIT('h8)
	) name19961 (
		_w30468_,
		_w30469_,
		_w30473_
	);
	LUT2 #(
		.INIT('h8)
	) name19962 (
		_w30466_,
		_w30467_,
		_w30474_
	);
	LUT2 #(
		.INIT('h8)
	) name19963 (
		_w30464_,
		_w30465_,
		_w30475_
	);
	LUT2 #(
		.INIT('h8)
	) name19964 (
		_w30474_,
		_w30475_,
		_w30476_
	);
	LUT2 #(
		.INIT('h8)
	) name19965 (
		_w30472_,
		_w30473_,
		_w30477_
	);
	LUT2 #(
		.INIT('h8)
	) name19966 (
		_w30476_,
		_w30477_,
		_w30478_
	);
	LUT2 #(
		.INIT('h1)
	) name19967 (
		wb_rst_i_pad,
		_w30478_,
		_w30479_
	);
	LUT2 #(
		.INIT('h1)
	) name19968 (
		_w22944_,
		_w30479_,
		_w30480_
	);
	LUT2 #(
		.INIT('h8)
	) name19969 (
		\ethreg1_MODER_1_DataOut_reg[6]/NET0131 ,
		_w23519_,
		_w30481_
	);
	LUT2 #(
		.INIT('h8)
	) name19970 (
		\ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 ,
		_w23499_,
		_w30482_
	);
	LUT2 #(
		.INIT('h8)
	) name19971 (
		\ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 ,
		_w22952_,
		_w30483_
	);
	LUT2 #(
		.INIT('h8)
	) name19972 (
		\ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 ,
		_w22956_,
		_w30484_
	);
	LUT2 #(
		.INIT('h8)
	) name19973 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 ,
		_w23522_,
		_w30485_
	);
	LUT2 #(
		.INIT('h8)
	) name19974 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		_w22959_,
		_w30486_
	);
	LUT2 #(
		.INIT('h8)
	) name19975 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		_w23501_,
		_w30487_
	);
	LUT2 #(
		.INIT('h8)
	) name19976 (
		\ethreg1_MIIRX_DATA_DataOut_reg[14]/NET0131 ,
		_w23507_,
		_w30488_
	);
	LUT2 #(
		.INIT('h8)
	) name19977 (
		\ethreg1_PACKETLEN_1_DataOut_reg[6]/NET0131 ,
		_w22966_,
		_w30489_
	);
	LUT2 #(
		.INIT('h1)
	) name19978 (
		_w30481_,
		_w30482_,
		_w30490_
	);
	LUT2 #(
		.INIT('h1)
	) name19979 (
		_w30483_,
		_w30484_,
		_w30491_
	);
	LUT2 #(
		.INIT('h1)
	) name19980 (
		_w30485_,
		_w30486_,
		_w30492_
	);
	LUT2 #(
		.INIT('h1)
	) name19981 (
		_w30487_,
		_w30488_,
		_w30493_
	);
	LUT2 #(
		.INIT('h8)
	) name19982 (
		_w30492_,
		_w30493_,
		_w30494_
	);
	LUT2 #(
		.INIT('h8)
	) name19983 (
		_w30490_,
		_w30491_,
		_w30495_
	);
	LUT2 #(
		.INIT('h8)
	) name19984 (
		_w22944_,
		_w30495_,
		_w30496_
	);
	LUT2 #(
		.INIT('h4)
	) name19985 (
		_w30489_,
		_w30494_,
		_w30497_
	);
	LUT2 #(
		.INIT('h8)
	) name19986 (
		_w30496_,
		_w30497_,
		_w30498_
	);
	LUT2 #(
		.INIT('h1)
	) name19987 (
		_w30480_,
		_w30498_,
		_w30499_
	);
	LUT2 #(
		.INIT('h1)
	) name19988 (
		_w15689_,
		_w22944_,
		_w30500_
	);
	LUT2 #(
		.INIT('h8)
	) name19989 (
		\ethreg1_MODER_1_DataOut_reg[7]/NET0131 ,
		_w23519_,
		_w30501_
	);
	LUT2 #(
		.INIT('h8)
	) name19990 (
		\ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 ,
		_w23499_,
		_w30502_
	);
	LUT2 #(
		.INIT('h8)
	) name19991 (
		\ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 ,
		_w22952_,
		_w30503_
	);
	LUT2 #(
		.INIT('h8)
	) name19992 (
		\ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 ,
		_w22956_,
		_w30504_
	);
	LUT2 #(
		.INIT('h8)
	) name19993 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 ,
		_w23522_,
		_w30505_
	);
	LUT2 #(
		.INIT('h8)
	) name19994 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		_w22959_,
		_w30506_
	);
	LUT2 #(
		.INIT('h8)
	) name19995 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		_w23501_,
		_w30507_
	);
	LUT2 #(
		.INIT('h8)
	) name19996 (
		\ethreg1_MIIRX_DATA_DataOut_reg[15]/NET0131 ,
		_w23507_,
		_w30508_
	);
	LUT2 #(
		.INIT('h8)
	) name19997 (
		\ethreg1_PACKETLEN_1_DataOut_reg[7]/NET0131 ,
		_w22966_,
		_w30509_
	);
	LUT2 #(
		.INIT('h1)
	) name19998 (
		_w30501_,
		_w30502_,
		_w30510_
	);
	LUT2 #(
		.INIT('h1)
	) name19999 (
		_w30503_,
		_w30504_,
		_w30511_
	);
	LUT2 #(
		.INIT('h1)
	) name20000 (
		_w30505_,
		_w30506_,
		_w30512_
	);
	LUT2 #(
		.INIT('h1)
	) name20001 (
		_w30507_,
		_w30508_,
		_w30513_
	);
	LUT2 #(
		.INIT('h8)
	) name20002 (
		_w30512_,
		_w30513_,
		_w30514_
	);
	LUT2 #(
		.INIT('h8)
	) name20003 (
		_w30510_,
		_w30511_,
		_w30515_
	);
	LUT2 #(
		.INIT('h8)
	) name20004 (
		_w22944_,
		_w30515_,
		_w30516_
	);
	LUT2 #(
		.INIT('h4)
	) name20005 (
		_w30509_,
		_w30514_,
		_w30517_
	);
	LUT2 #(
		.INIT('h8)
	) name20006 (
		_w30516_,
		_w30517_,
		_w30518_
	);
	LUT2 #(
		.INIT('h1)
	) name20007 (
		_w30500_,
		_w30518_,
		_w30519_
	);
	LUT2 #(
		.INIT('h8)
	) name20008 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w17858_,
		_w30520_
	);
	LUT2 #(
		.INIT('h1)
	) name20009 (
		\wishbone_RxPointerMSB_reg[12]/NET0131 ,
		_w17858_,
		_w30521_
	);
	LUT2 #(
		.INIT('h1)
	) name20010 (
		_w15696_,
		_w30520_,
		_w30522_
	);
	LUT2 #(
		.INIT('h4)
	) name20011 (
		_w30521_,
		_w30522_,
		_w30523_
	);
	LUT2 #(
		.INIT('h8)
	) name20012 (
		_w15696_,
		_w23494_,
		_w30524_
	);
	LUT2 #(
		.INIT('h1)
	) name20013 (
		_w30523_,
		_w30524_,
		_w30525_
	);
	LUT2 #(
		.INIT('h1)
	) name20014 (
		\wishbone_RxPointerMSB_reg[14]/NET0131 ,
		_w17860_,
		_w30526_
	);
	LUT2 #(
		.INIT('h1)
	) name20015 (
		_w15696_,
		_w17861_,
		_w30527_
	);
	LUT2 #(
		.INIT('h4)
	) name20016 (
		_w30526_,
		_w30527_,
		_w30528_
	);
	LUT2 #(
		.INIT('h8)
	) name20017 (
		_w15696_,
		_w30479_,
		_w30529_
	);
	LUT2 #(
		.INIT('h1)
	) name20018 (
		_w30528_,
		_w30529_,
		_w30530_
	);
	LUT2 #(
		.INIT('h1)
	) name20019 (
		\wishbone_RxPointerMSB_reg[4]/NET0131 ,
		_w17850_,
		_w30531_
	);
	LUT2 #(
		.INIT('h1)
	) name20020 (
		_w15696_,
		_w17851_,
		_w30532_
	);
	LUT2 #(
		.INIT('h4)
	) name20021 (
		_w30531_,
		_w30532_,
		_w30533_
	);
	LUT2 #(
		.INIT('h8)
	) name20022 (
		_w15696_,
		_w25266_,
		_w30534_
	);
	LUT2 #(
		.INIT('h1)
	) name20023 (
		_w30533_,
		_w30534_,
		_w30535_
	);
	LUT2 #(
		.INIT('h1)
	) name20024 (
		\wishbone_RxPointerMSB_reg[5]/NET0131 ,
		_w17851_,
		_w30536_
	);
	LUT2 #(
		.INIT('h1)
	) name20025 (
		_w15696_,
		_w17852_,
		_w30537_
	);
	LUT2 #(
		.INIT('h4)
	) name20026 (
		_w30536_,
		_w30537_,
		_w30538_
	);
	LUT2 #(
		.INIT('h8)
	) name20027 (
		_w15696_,
		_w25816_,
		_w30539_
	);
	LUT2 #(
		.INIT('h1)
	) name20028 (
		_w30538_,
		_w30539_,
		_w30540_
	);
	LUT2 #(
		.INIT('h1)
	) name20029 (
		\wishbone_RxPointerMSB_reg[7]/NET0131 ,
		_w17853_,
		_w30541_
	);
	LUT2 #(
		.INIT('h1)
	) name20030 (
		_w15696_,
		_w17854_,
		_w30542_
	);
	LUT2 #(
		.INIT('h4)
	) name20031 (
		_w30541_,
		_w30542_,
		_w30543_
	);
	LUT2 #(
		.INIT('h8)
	) name20032 (
		_w15696_,
		_w26364_,
		_w30544_
	);
	LUT2 #(
		.INIT('h1)
	) name20033 (
		_w30543_,
		_w30544_,
		_w30545_
	);
	LUT2 #(
		.INIT('h1)
	) name20034 (
		\wishbone_RxPointerMSB_reg[6]/NET0131 ,
		_w17852_,
		_w30546_
	);
	LUT2 #(
		.INIT('h1)
	) name20035 (
		_w15696_,
		_w17853_,
		_w30547_
	);
	LUT2 #(
		.INIT('h4)
	) name20036 (
		_w30546_,
		_w30547_,
		_w30548_
	);
	LUT2 #(
		.INIT('h8)
	) name20037 (
		_w15696_,
		_w29218_,
		_w30549_
	);
	LUT2 #(
		.INIT('h1)
	) name20038 (
		_w30548_,
		_w30549_,
		_w30550_
	);
	LUT2 #(
		.INIT('h1)
	) name20039 (
		\wishbone_TxPointerMSB_reg[12]/NET0131 ,
		_w17895_,
		_w30551_
	);
	LUT2 #(
		.INIT('h1)
	) name20040 (
		_w17883_,
		_w17896_,
		_w30552_
	);
	LUT2 #(
		.INIT('h4)
	) name20041 (
		_w30551_,
		_w30552_,
		_w30553_
	);
	LUT2 #(
		.INIT('h8)
	) name20042 (
		_w17883_,
		_w23494_,
		_w30554_
	);
	LUT2 #(
		.INIT('h1)
	) name20043 (
		_w30553_,
		_w30554_,
		_w30555_
	);
	LUT2 #(
		.INIT('h8)
	) name20044 (
		_w17883_,
		_w30479_,
		_w30556_
	);
	LUT2 #(
		.INIT('h8)
	) name20045 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		_w17896_,
		_w30557_
	);
	LUT2 #(
		.INIT('h1)
	) name20046 (
		\wishbone_TxPointerMSB_reg[14]/NET0131 ,
		_w30557_,
		_w30558_
	);
	LUT2 #(
		.INIT('h1)
	) name20047 (
		_w17883_,
		_w17898_,
		_w30559_
	);
	LUT2 #(
		.INIT('h4)
	) name20048 (
		_w30558_,
		_w30559_,
		_w30560_
	);
	LUT2 #(
		.INIT('h1)
	) name20049 (
		_w30556_,
		_w30560_,
		_w30561_
	);
	LUT2 #(
		.INIT('h1)
	) name20050 (
		\wishbone_TxPointerMSB_reg[4]/NET0131 ,
		_w17887_,
		_w30562_
	);
	LUT2 #(
		.INIT('h1)
	) name20051 (
		_w17883_,
		_w17888_,
		_w30563_
	);
	LUT2 #(
		.INIT('h4)
	) name20052 (
		_w30562_,
		_w30563_,
		_w30564_
	);
	LUT2 #(
		.INIT('h8)
	) name20053 (
		_w17883_,
		_w25266_,
		_w30565_
	);
	LUT2 #(
		.INIT('h1)
	) name20054 (
		_w30564_,
		_w30565_,
		_w30566_
	);
	LUT2 #(
		.INIT('h1)
	) name20055 (
		\wishbone_TxPointerMSB_reg[5]/NET0131 ,
		_w17888_,
		_w30567_
	);
	LUT2 #(
		.INIT('h1)
	) name20056 (
		_w17883_,
		_w17889_,
		_w30568_
	);
	LUT2 #(
		.INIT('h4)
	) name20057 (
		_w30567_,
		_w30568_,
		_w30569_
	);
	LUT2 #(
		.INIT('h8)
	) name20058 (
		_w17883_,
		_w25816_,
		_w30570_
	);
	LUT2 #(
		.INIT('h1)
	) name20059 (
		_w30569_,
		_w30570_,
		_w30571_
	);
	LUT2 #(
		.INIT('h1)
	) name20060 (
		\wishbone_TxPointerMSB_reg[6]/NET0131 ,
		_w17889_,
		_w30572_
	);
	LUT2 #(
		.INIT('h1)
	) name20061 (
		_w17883_,
		_w17890_,
		_w30573_
	);
	LUT2 #(
		.INIT('h4)
	) name20062 (
		_w30572_,
		_w30573_,
		_w30574_
	);
	LUT2 #(
		.INIT('h8)
	) name20063 (
		_w17883_,
		_w29218_,
		_w30575_
	);
	LUT2 #(
		.INIT('h1)
	) name20064 (
		_w30574_,
		_w30575_,
		_w30576_
	);
	LUT2 #(
		.INIT('h1)
	) name20065 (
		\wishbone_TxPointerMSB_reg[7]/NET0131 ,
		_w17890_,
		_w30577_
	);
	LUT2 #(
		.INIT('h1)
	) name20066 (
		_w17883_,
		_w17891_,
		_w30578_
	);
	LUT2 #(
		.INIT('h4)
	) name20067 (
		_w30577_,
		_w30578_,
		_w30579_
	);
	LUT2 #(
		.INIT('h8)
	) name20068 (
		_w17883_,
		_w26364_,
		_w30580_
	);
	LUT2 #(
		.INIT('h1)
	) name20069 (
		_w30579_,
		_w30580_,
		_w30581_
	);
	LUT2 #(
		.INIT('h1)
	) name20070 (
		\wishbone_RxPointerMSB_reg[11]/NET0131 ,
		_w17857_,
		_w30582_
	);
	LUT2 #(
		.INIT('h1)
	) name20071 (
		_w15696_,
		_w17858_,
		_w30583_
	);
	LUT2 #(
		.INIT('h4)
	) name20072 (
		_w30582_,
		_w30583_,
		_w30584_
	);
	LUT2 #(
		.INIT('h8)
	) name20073 (
		_w15696_,
		_w27980_,
		_w30585_
	);
	LUT2 #(
		.INIT('h1)
	) name20074 (
		_w30584_,
		_w30585_,
		_w30586_
	);
	LUT2 #(
		.INIT('h8)
	) name20075 (
		_w15696_,
		_w29947_,
		_w30587_
	);
	LUT2 #(
		.INIT('h1)
	) name20076 (
		\wishbone_RxPointerMSB_reg[13]/NET0131 ,
		_w30520_,
		_w30588_
	);
	LUT2 #(
		.INIT('h1)
	) name20077 (
		_w15696_,
		_w17860_,
		_w30589_
	);
	LUT2 #(
		.INIT('h4)
	) name20078 (
		_w30588_,
		_w30589_,
		_w30590_
	);
	LUT2 #(
		.INIT('h1)
	) name20079 (
		_w30587_,
		_w30590_,
		_w30591_
	);
	LUT2 #(
		.INIT('h1)
	) name20080 (
		\wishbone_RxPointerMSB_reg[15]/NET0131 ,
		_w17861_,
		_w30592_
	);
	LUT2 #(
		.INIT('h1)
	) name20081 (
		_w15696_,
		_w17862_,
		_w30593_
	);
	LUT2 #(
		.INIT('h4)
	) name20082 (
		_w30592_,
		_w30593_,
		_w30594_
	);
	LUT2 #(
		.INIT('h8)
	) name20083 (
		_w15689_,
		_w15696_,
		_w30595_
	);
	LUT2 #(
		.INIT('h1)
	) name20084 (
		_w30594_,
		_w30595_,
		_w30596_
	);
	LUT2 #(
		.INIT('h1)
	) name20085 (
		\wishbone_RxPointerMSB_reg[16]/NET0131 ,
		_w17862_,
		_w30597_
	);
	LUT2 #(
		.INIT('h1)
	) name20086 (
		_w15696_,
		_w29290_,
		_w30598_
	);
	LUT2 #(
		.INIT('h4)
	) name20087 (
		_w30597_,
		_w30598_,
		_w30599_
	);
	LUT2 #(
		.INIT('h8)
	) name20088 (
		_w15696_,
		_w19088_,
		_w30600_
	);
	LUT2 #(
		.INIT('h1)
	) name20089 (
		_w30599_,
		_w30600_,
		_w30601_
	);
	LUT2 #(
		.INIT('h1)
	) name20090 (
		\wishbone_RxPointerMSB_reg[17]/NET0131 ,
		_w29290_,
		_w30602_
	);
	LUT2 #(
		.INIT('h1)
	) name20091 (
		_w15696_,
		_w29291_,
		_w30603_
	);
	LUT2 #(
		.INIT('h4)
	) name20092 (
		_w30602_,
		_w30603_,
		_w30604_
	);
	LUT2 #(
		.INIT('h8)
	) name20093 (
		_w15696_,
		_w20126_,
		_w30605_
	);
	LUT2 #(
		.INIT('h1)
	) name20094 (
		_w30604_,
		_w30605_,
		_w30606_
	);
	LUT2 #(
		.INIT('h1)
	) name20095 (
		\wishbone_RxPointerMSB_reg[18]/NET0131 ,
		_w29291_,
		_w30607_
	);
	LUT2 #(
		.INIT('h1)
	) name20096 (
		_w15696_,
		_w29292_,
		_w30608_
	);
	LUT2 #(
		.INIT('h4)
	) name20097 (
		_w30607_,
		_w30608_,
		_w30609_
	);
	LUT2 #(
		.INIT('h8)
	) name20098 (
		_w15696_,
		_w18564_,
		_w30610_
	);
	LUT2 #(
		.INIT('h1)
	) name20099 (
		_w30609_,
		_w30610_,
		_w30611_
	);
	LUT2 #(
		.INIT('h1)
	) name20100 (
		\wishbone_RxPointerMSB_reg[2]/NET0131 ,
		_w15698_,
		_w30612_
	);
	LUT2 #(
		.INIT('h1)
	) name20101 (
		_w15696_,
		_w17849_,
		_w30613_
	);
	LUT2 #(
		.INIT('h4)
	) name20102 (
		_w30612_,
		_w30613_,
		_w30614_
	);
	LUT2 #(
		.INIT('h8)
	) name20103 (
		_w15696_,
		_w28520_,
		_w30615_
	);
	LUT2 #(
		.INIT('h1)
	) name20104 (
		_w30614_,
		_w30615_,
		_w30616_
	);
	LUT2 #(
		.INIT('h1)
	) name20105 (
		\wishbone_RxPointerMSB_reg[3]/NET0131 ,
		_w17849_,
		_w30617_
	);
	LUT2 #(
		.INIT('h1)
	) name20106 (
		_w15696_,
		_w17850_,
		_w30618_
	);
	LUT2 #(
		.INIT('h4)
	) name20107 (
		_w30617_,
		_w30618_,
		_w30619_
	);
	LUT2 #(
		.INIT('h8)
	) name20108 (
		_w15696_,
		_w24704_,
		_w30620_
	);
	LUT2 #(
		.INIT('h1)
	) name20109 (
		_w30619_,
		_w30620_,
		_w30621_
	);
	LUT2 #(
		.INIT('h1)
	) name20110 (
		\wishbone_RxPointerMSB_reg[8]/NET0131 ,
		_w17854_,
		_w30622_
	);
	LUT2 #(
		.INIT('h1)
	) name20111 (
		_w15696_,
		_w29357_,
		_w30623_
	);
	LUT2 #(
		.INIT('h4)
	) name20112 (
		_w30622_,
		_w30623_,
		_w30624_
	);
	LUT2 #(
		.INIT('h8)
	) name20113 (
		_w15696_,
		_w26900_,
		_w30625_
	);
	LUT2 #(
		.INIT('h1)
	) name20114 (
		_w30624_,
		_w30625_,
		_w30626_
	);
	LUT2 #(
		.INIT('h1)
	) name20115 (
		\wishbone_TxPointerMSB_reg[10]/NET0131 ,
		_w17893_,
		_w30627_
	);
	LUT2 #(
		.INIT('h1)
	) name20116 (
		_w17883_,
		_w17894_,
		_w30628_
	);
	LUT2 #(
		.INIT('h4)
	) name20117 (
		_w30627_,
		_w30628_,
		_w30629_
	);
	LUT2 #(
		.INIT('h8)
	) name20118 (
		\wishbone_bd_ram_mem1_reg[124][10]/P0001 ,
		_w13058_,
		_w30630_
	);
	LUT2 #(
		.INIT('h8)
	) name20119 (
		\wishbone_bd_ram_mem1_reg[3][10]/P0001 ,
		_w12866_,
		_w30631_
	);
	LUT2 #(
		.INIT('h8)
	) name20120 (
		\wishbone_bd_ram_mem1_reg[164][10]/P0001 ,
		_w12876_,
		_w30632_
	);
	LUT2 #(
		.INIT('h8)
	) name20121 (
		\wishbone_bd_ram_mem1_reg[29][10]/P0001 ,
		_w12952_,
		_w30633_
	);
	LUT2 #(
		.INIT('h8)
	) name20122 (
		\wishbone_bd_ram_mem1_reg[210][10]/P0001 ,
		_w12924_,
		_w30634_
	);
	LUT2 #(
		.INIT('h8)
	) name20123 (
		\wishbone_bd_ram_mem1_reg[159][10]/P0001 ,
		_w12774_,
		_w30635_
	);
	LUT2 #(
		.INIT('h8)
	) name20124 (
		\wishbone_bd_ram_mem1_reg[43][10]/P0001 ,
		_w13200_,
		_w30636_
	);
	LUT2 #(
		.INIT('h8)
	) name20125 (
		\wishbone_bd_ram_mem1_reg[253][10]/P0001 ,
		_w13100_,
		_w30637_
	);
	LUT2 #(
		.INIT('h8)
	) name20126 (
		\wishbone_bd_ram_mem1_reg[60][10]/P0001 ,
		_w13204_,
		_w30638_
	);
	LUT2 #(
		.INIT('h8)
	) name20127 (
		\wishbone_bd_ram_mem1_reg[30][10]/P0001 ,
		_w13104_,
		_w30639_
	);
	LUT2 #(
		.INIT('h8)
	) name20128 (
		\wishbone_bd_ram_mem1_reg[242][10]/P0001 ,
		_w12932_,
		_w30640_
	);
	LUT2 #(
		.INIT('h8)
	) name20129 (
		\wishbone_bd_ram_mem1_reg[48][10]/P0001 ,
		_w12970_,
		_w30641_
	);
	LUT2 #(
		.INIT('h8)
	) name20130 (
		\wishbone_bd_ram_mem1_reg[77][10]/P0001 ,
		_w12982_,
		_w30642_
	);
	LUT2 #(
		.INIT('h8)
	) name20131 (
		\wishbone_bd_ram_mem1_reg[249][10]/P0001 ,
		_w12900_,
		_w30643_
	);
	LUT2 #(
		.INIT('h8)
	) name20132 (
		\wishbone_bd_ram_mem1_reg[119][10]/P0001 ,
		_w13048_,
		_w30644_
	);
	LUT2 #(
		.INIT('h8)
	) name20133 (
		\wishbone_bd_ram_mem1_reg[92][10]/P0001 ,
		_w13010_,
		_w30645_
	);
	LUT2 #(
		.INIT('h8)
	) name20134 (
		\wishbone_bd_ram_mem1_reg[141][10]/P0001 ,
		_w13004_,
		_w30646_
	);
	LUT2 #(
		.INIT('h8)
	) name20135 (
		\wishbone_bd_ram_mem1_reg[137][10]/P0001 ,
		_w13168_,
		_w30647_
	);
	LUT2 #(
		.INIT('h8)
	) name20136 (
		\wishbone_bd_ram_mem1_reg[191][10]/P0001 ,
		_w13034_,
		_w30648_
	);
	LUT2 #(
		.INIT('h8)
	) name20137 (
		\wishbone_bd_ram_mem1_reg[177][10]/P0001 ,
		_w12996_,
		_w30649_
	);
	LUT2 #(
		.INIT('h8)
	) name20138 (
		\wishbone_bd_ram_mem1_reg[103][10]/P0001 ,
		_w12846_,
		_w30650_
	);
	LUT2 #(
		.INIT('h8)
	) name20139 (
		\wishbone_bd_ram_mem1_reg[56][10]/P0001 ,
		_w12778_,
		_w30651_
	);
	LUT2 #(
		.INIT('h8)
	) name20140 (
		\wishbone_bd_ram_mem1_reg[220][10]/P0001 ,
		_w13066_,
		_w30652_
	);
	LUT2 #(
		.INIT('h8)
	) name20141 (
		\wishbone_bd_ram_mem1_reg[131][10]/P0001 ,
		_w12852_,
		_w30653_
	);
	LUT2 #(
		.INIT('h8)
	) name20142 (
		\wishbone_bd_ram_mem1_reg[228][10]/P0001 ,
		_w12765_,
		_w30654_
	);
	LUT2 #(
		.INIT('h8)
	) name20143 (
		\wishbone_bd_ram_mem1_reg[65][10]/P0001 ,
		_w13176_,
		_w30655_
	);
	LUT2 #(
		.INIT('h8)
	) name20144 (
		\wishbone_bd_ram_mem1_reg[189][10]/P0001 ,
		_w13042_,
		_w30656_
	);
	LUT2 #(
		.INIT('h8)
	) name20145 (
		\wishbone_bd_ram_mem1_reg[82][10]/P0001 ,
		_w12942_,
		_w30657_
	);
	LUT2 #(
		.INIT('h8)
	) name20146 (
		\wishbone_bd_ram_mem1_reg[70][10]/P0001 ,
		_w12840_,
		_w30658_
	);
	LUT2 #(
		.INIT('h8)
	) name20147 (
		\wishbone_bd_ram_mem1_reg[10][10]/P0001 ,
		_w13172_,
		_w30659_
	);
	LUT2 #(
		.INIT('h8)
	) name20148 (
		\wishbone_bd_ram_mem1_reg[219][10]/P0001 ,
		_w12806_,
		_w30660_
	);
	LUT2 #(
		.INIT('h8)
	) name20149 (
		\wishbone_bd_ram_mem1_reg[236][10]/P0001 ,
		_w12731_,
		_w30661_
	);
	LUT2 #(
		.INIT('h8)
	) name20150 (
		\wishbone_bd_ram_mem1_reg[206][10]/P0001 ,
		_w12954_,
		_w30662_
	);
	LUT2 #(
		.INIT('h8)
	) name20151 (
		\wishbone_bd_ram_mem1_reg[163][10]/P0001 ,
		_w12882_,
		_w30663_
	);
	LUT2 #(
		.INIT('h8)
	) name20152 (
		\wishbone_bd_ram_mem1_reg[187][10]/P0001 ,
		_w13196_,
		_w30664_
	);
	LUT2 #(
		.INIT('h8)
	) name20153 (
		\wishbone_bd_ram_mem1_reg[162][10]/P0001 ,
		_w13098_,
		_w30665_
	);
	LUT2 #(
		.INIT('h8)
	) name20154 (
		\wishbone_bd_ram_mem1_reg[22][10]/P0001 ,
		_w13110_,
		_w30666_
	);
	LUT2 #(
		.INIT('h8)
	) name20155 (
		\wishbone_bd_ram_mem1_reg[140][10]/P0001 ,
		_w12894_,
		_w30667_
	);
	LUT2 #(
		.INIT('h8)
	) name20156 (
		\wishbone_bd_ram_mem1_reg[111][10]/P0001 ,
		_w12744_,
		_w30668_
	);
	LUT2 #(
		.INIT('h8)
	) name20157 (
		\wishbone_bd_ram_mem1_reg[165][10]/P0001 ,
		_w13044_,
		_w30669_
	);
	LUT2 #(
		.INIT('h8)
	) name20158 (
		\wishbone_bd_ram_mem1_reg[44][10]/P0001 ,
		_w12896_,
		_w30670_
	);
	LUT2 #(
		.INIT('h8)
	) name20159 (
		\wishbone_bd_ram_mem1_reg[188][10]/P0001 ,
		_w12948_,
		_w30671_
	);
	LUT2 #(
		.INIT('h8)
	) name20160 (
		\wishbone_bd_ram_mem1_reg[31][10]/P0001 ,
		_w13198_,
		_w30672_
	);
	LUT2 #(
		.INIT('h8)
	) name20161 (
		\wishbone_bd_ram_mem1_reg[96][10]/P0001 ,
		_w12912_,
		_w30673_
	);
	LUT2 #(
		.INIT('h8)
	) name20162 (
		\wishbone_bd_ram_mem1_reg[12][10]/P0001 ,
		_w13118_,
		_w30674_
	);
	LUT2 #(
		.INIT('h8)
	) name20163 (
		\wishbone_bd_ram_mem1_reg[99][10]/P0001 ,
		_w13038_,
		_w30675_
	);
	LUT2 #(
		.INIT('h8)
	) name20164 (
		\wishbone_bd_ram_mem1_reg[41][10]/P0001 ,
		_w13052_,
		_w30676_
	);
	LUT2 #(
		.INIT('h8)
	) name20165 (
		\wishbone_bd_ram_mem1_reg[54][10]/P0001 ,
		_w12770_,
		_w30677_
	);
	LUT2 #(
		.INIT('h8)
	) name20166 (
		\wishbone_bd_ram_mem1_reg[90][10]/P0001 ,
		_w12978_,
		_w30678_
	);
	LUT2 #(
		.INIT('h8)
	) name20167 (
		\wishbone_bd_ram_mem1_reg[252][10]/P0001 ,
		_w13080_,
		_w30679_
	);
	LUT2 #(
		.INIT('h8)
	) name20168 (
		\wishbone_bd_ram_mem1_reg[39][10]/P0001 ,
		_w13018_,
		_w30680_
	);
	LUT2 #(
		.INIT('h8)
	) name20169 (
		\wishbone_bd_ram_mem1_reg[175][10]/P0001 ,
		_w13126_,
		_w30681_
	);
	LUT2 #(
		.INIT('h8)
	) name20170 (
		\wishbone_bd_ram_mem1_reg[28][10]/P0001 ,
		_w13170_,
		_w30682_
	);
	LUT2 #(
		.INIT('h8)
	) name20171 (
		\wishbone_bd_ram_mem1_reg[100][10]/P0001 ,
		_w12960_,
		_w30683_
	);
	LUT2 #(
		.INIT('h8)
	) name20172 (
		\wishbone_bd_ram_mem1_reg[102][10]/P0001 ,
		_w12685_,
		_w30684_
	);
	LUT2 #(
		.INIT('h8)
	) name20173 (
		\wishbone_bd_ram_mem1_reg[161][10]/P0001 ,
		_w12754_,
		_w30685_
	);
	LUT2 #(
		.INIT('h8)
	) name20174 (
		\wishbone_bd_ram_mem1_reg[151][10]/P0001 ,
		_w13142_,
		_w30686_
	);
	LUT2 #(
		.INIT('h8)
	) name20175 (
		\wishbone_bd_ram_mem1_reg[240][10]/P0001 ,
		_w12864_,
		_w30687_
	);
	LUT2 #(
		.INIT('h8)
	) name20176 (
		\wishbone_bd_ram_mem1_reg[122][10]/P0001 ,
		_w13130_,
		_w30688_
	);
	LUT2 #(
		.INIT('h8)
	) name20177 (
		\wishbone_bd_ram_mem1_reg[215][10]/P0001 ,
		_w12974_,
		_w30689_
	);
	LUT2 #(
		.INIT('h8)
	) name20178 (
		\wishbone_bd_ram_mem1_reg[184][10]/P0001 ,
		_w13062_,
		_w30690_
	);
	LUT2 #(
		.INIT('h8)
	) name20179 (
		\wishbone_bd_ram_mem1_reg[139][10]/P0001 ,
		_w12814_,
		_w30691_
	);
	LUT2 #(
		.INIT('h8)
	) name20180 (
		\wishbone_bd_ram_mem1_reg[93][10]/P0001 ,
		_w13016_,
		_w30692_
	);
	LUT2 #(
		.INIT('h8)
	) name20181 (
		\wishbone_bd_ram_mem1_reg[76][10]/P0001 ,
		_w13184_,
		_w30693_
	);
	LUT2 #(
		.INIT('h8)
	) name20182 (
		\wishbone_bd_ram_mem1_reg[38][10]/P0001 ,
		_w13182_,
		_w30694_
	);
	LUT2 #(
		.INIT('h8)
	) name20183 (
		\wishbone_bd_ram_mem1_reg[64][10]/P0001 ,
		_w12976_,
		_w30695_
	);
	LUT2 #(
		.INIT('h8)
	) name20184 (
		\wishbone_bd_ram_mem1_reg[132][10]/P0001 ,
		_w12992_,
		_w30696_
	);
	LUT2 #(
		.INIT('h8)
	) name20185 (
		\wishbone_bd_ram_mem1_reg[235][10]/P0001 ,
		_w12696_,
		_w30697_
	);
	LUT2 #(
		.INIT('h8)
	) name20186 (
		\wishbone_bd_ram_mem1_reg[200][10]/P0001 ,
		_w12988_,
		_w30698_
	);
	LUT2 #(
		.INIT('h8)
	) name20187 (
		\wishbone_bd_ram_mem1_reg[148][10]/P0001 ,
		_w13000_,
		_w30699_
	);
	LUT2 #(
		.INIT('h8)
	) name20188 (
		\wishbone_bd_ram_mem1_reg[230][10]/P0001 ,
		_w13036_,
		_w30700_
	);
	LUT2 #(
		.INIT('h8)
	) name20189 (
		\wishbone_bd_ram_mem1_reg[14][10]/P0001 ,
		_w13086_,
		_w30701_
	);
	LUT2 #(
		.INIT('h8)
	) name20190 (
		\wishbone_bd_ram_mem1_reg[17][10]/P0001 ,
		_w12848_,
		_w30702_
	);
	LUT2 #(
		.INIT('h8)
	) name20191 (
		\wishbone_bd_ram_mem1_reg[0][10]/P0001 ,
		_w12717_,
		_w30703_
	);
	LUT2 #(
		.INIT('h8)
	) name20192 (
		\wishbone_bd_ram_mem1_reg[27][10]/P0001 ,
		_w12880_,
		_w30704_
	);
	LUT2 #(
		.INIT('h8)
	) name20193 (
		\wishbone_bd_ram_mem1_reg[158][10]/P0001 ,
		_w12898_,
		_w30705_
	);
	LUT2 #(
		.INIT('h8)
	) name20194 (
		\wishbone_bd_ram_mem1_reg[255][10]/P0001 ,
		_w13072_,
		_w30706_
	);
	LUT2 #(
		.INIT('h8)
	) name20195 (
		\wishbone_bd_ram_mem1_reg[71][10]/P0001 ,
		_w12798_,
		_w30707_
	);
	LUT2 #(
		.INIT('h8)
	) name20196 (
		\wishbone_bd_ram_mem1_reg[127][10]/P0001 ,
		_w13164_,
		_w30708_
	);
	LUT2 #(
		.INIT('h8)
	) name20197 (
		\wishbone_bd_ram_mem1_reg[21][10]/P0001 ,
		_w12906_,
		_w30709_
	);
	LUT2 #(
		.INIT('h8)
	) name20198 (
		\wishbone_bd_ram_mem1_reg[134][10]/P0001 ,
		_w12763_,
		_w30710_
	);
	LUT2 #(
		.INIT('h8)
	) name20199 (
		\wishbone_bd_ram_mem1_reg[199][10]/P0001 ,
		_w12768_,
		_w30711_
	);
	LUT2 #(
		.INIT('h8)
	) name20200 (
		\wishbone_bd_ram_mem1_reg[112][10]/P0001 ,
		_w12733_,
		_w30712_
	);
	LUT2 #(
		.INIT('h8)
	) name20201 (
		\wishbone_bd_ram_mem1_reg[78][10]/P0001 ,
		_w12874_,
		_w30713_
	);
	LUT2 #(
		.INIT('h8)
	) name20202 (
		\wishbone_bd_ram_mem1_reg[20][10]/P0001 ,
		_w13174_,
		_w30714_
	);
	LUT2 #(
		.INIT('h8)
	) name20203 (
		\wishbone_bd_ram_mem1_reg[88][10]/P0001 ,
		_w12860_,
		_w30715_
	);
	LUT2 #(
		.INIT('h8)
	) name20204 (
		\wishbone_bd_ram_mem1_reg[33][10]/P0001 ,
		_w12980_,
		_w30716_
	);
	LUT2 #(
		.INIT('h8)
	) name20205 (
		\wishbone_bd_ram_mem1_reg[222][10]/P0001 ,
		_w13094_,
		_w30717_
	);
	LUT2 #(
		.INIT('h8)
	) name20206 (
		\wishbone_bd_ram_mem1_reg[193][10]/P0001 ,
		_w13056_,
		_w30718_
	);
	LUT2 #(
		.INIT('h8)
	) name20207 (
		\wishbone_bd_ram_mem1_reg[116][10]/P0001 ,
		_w12998_,
		_w30719_
	);
	LUT2 #(
		.INIT('h8)
	) name20208 (
		\wishbone_bd_ram_mem1_reg[251][10]/P0001 ,
		_w13054_,
		_w30720_
	);
	LUT2 #(
		.INIT('h8)
	) name20209 (
		\wishbone_bd_ram_mem1_reg[113][10]/P0001 ,
		_w13026_,
		_w30721_
	);
	LUT2 #(
		.INIT('h8)
	) name20210 (
		\wishbone_bd_ram_mem1_reg[208][10]/P0001 ,
		_w13032_,
		_w30722_
	);
	LUT2 #(
		.INIT('h8)
	) name20211 (
		\wishbone_bd_ram_mem1_reg[107][10]/P0001 ,
		_w12749_,
		_w30723_
	);
	LUT2 #(
		.INIT('h8)
	) name20212 (
		\wishbone_bd_ram_mem1_reg[118][10]/P0001 ,
		_w12830_,
		_w30724_
	);
	LUT2 #(
		.INIT('h8)
	) name20213 (
		\wishbone_bd_ram_mem1_reg[155][10]/P0001 ,
		_w13122_,
		_w30725_
	);
	LUT2 #(
		.INIT('h8)
	) name20214 (
		\wishbone_bd_ram_mem1_reg[83][10]/P0001 ,
		_w12916_,
		_w30726_
	);
	LUT2 #(
		.INIT('h8)
	) name20215 (
		\wishbone_bd_ram_mem1_reg[79][10]/P0001 ,
		_w13212_,
		_w30727_
	);
	LUT2 #(
		.INIT('h8)
	) name20216 (
		\wishbone_bd_ram_mem1_reg[204][10]/P0001 ,
		_w13162_,
		_w30728_
	);
	LUT2 #(
		.INIT('h8)
	) name20217 (
		\wishbone_bd_ram_mem1_reg[243][10]/P0001 ,
		_w12804_,
		_w30729_
	);
	LUT2 #(
		.INIT('h8)
	) name20218 (
		\wishbone_bd_ram_mem1_reg[241][10]/P0001 ,
		_w13006_,
		_w30730_
	);
	LUT2 #(
		.INIT('h8)
	) name20219 (
		\wishbone_bd_ram_mem1_reg[146][10]/P0001 ,
		_w13060_,
		_w30731_
	);
	LUT2 #(
		.INIT('h8)
	) name20220 (
		\wishbone_bd_ram_mem1_reg[18][10]/P0001 ,
		_w12679_,
		_w30732_
	);
	LUT2 #(
		.INIT('h8)
	) name20221 (
		\wishbone_bd_ram_mem1_reg[58][10]/P0001 ,
		_w13070_,
		_w30733_
	);
	LUT2 #(
		.INIT('h8)
	) name20222 (
		\wishbone_bd_ram_mem1_reg[133][10]/P0001 ,
		_w12761_,
		_w30734_
	);
	LUT2 #(
		.INIT('h8)
	) name20223 (
		\wishbone_bd_ram_mem1_reg[52][10]/P0001 ,
		_w13082_,
		_w30735_
	);
	LUT2 #(
		.INIT('h8)
	) name20224 (
		\wishbone_bd_ram_mem1_reg[136][10]/P0001 ,
		_w13064_,
		_w30736_
	);
	LUT2 #(
		.INIT('h8)
	) name20225 (
		\wishbone_bd_ram_mem1_reg[86][10]/P0001 ,
		_w12735_,
		_w30737_
	);
	LUT2 #(
		.INIT('h8)
	) name20226 (
		\wishbone_bd_ram_mem1_reg[24][10]/P0001 ,
		_w13084_,
		_w30738_
	);
	LUT2 #(
		.INIT('h8)
	) name20227 (
		\wishbone_bd_ram_mem1_reg[149][10]/P0001 ,
		_w12741_,
		_w30739_
	);
	LUT2 #(
		.INIT('h8)
	) name20228 (
		\wishbone_bd_ram_mem1_reg[32][10]/P0001 ,
		_w13120_,
		_w30740_
	);
	LUT2 #(
		.INIT('h8)
	) name20229 (
		\wishbone_bd_ram_mem1_reg[42][10]/P0001 ,
		_w12842_,
		_w30741_
	);
	LUT2 #(
		.INIT('h8)
	) name20230 (
		\wishbone_bd_ram_mem1_reg[49][10]/P0001 ,
		_w12994_,
		_w30742_
	);
	LUT2 #(
		.INIT('h8)
	) name20231 (
		\wishbone_bd_ram_mem1_reg[128][10]/P0001 ,
		_w12793_,
		_w30743_
	);
	LUT2 #(
		.INIT('h8)
	) name20232 (
		\wishbone_bd_ram_mem1_reg[245][10]/P0001 ,
		_w13022_,
		_w30744_
	);
	LUT2 #(
		.INIT('h8)
	) name20233 (
		\wishbone_bd_ram_mem1_reg[120][10]/P0001 ,
		_w12707_,
		_w30745_
	);
	LUT2 #(
		.INIT('h8)
	) name20234 (
		\wishbone_bd_ram_mem1_reg[247][10]/P0001 ,
		_w12818_,
		_w30746_
	);
	LUT2 #(
		.INIT('h8)
	) name20235 (
		\wishbone_bd_ram_mem1_reg[180][10]/P0001 ,
		_w12791_,
		_w30747_
	);
	LUT2 #(
		.INIT('h8)
	) name20236 (
		\wishbone_bd_ram_mem1_reg[225][10]/P0001 ,
		_w13092_,
		_w30748_
	);
	LUT2 #(
		.INIT('h8)
	) name20237 (
		\wishbone_bd_ram_mem1_reg[145][10]/P0001 ,
		_w13106_,
		_w30749_
	);
	LUT2 #(
		.INIT('h8)
	) name20238 (
		\wishbone_bd_ram_mem1_reg[196][10]/P0001 ,
		_w13090_,
		_w30750_
	);
	LUT2 #(
		.INIT('h8)
	) name20239 (
		\wishbone_bd_ram_mem1_reg[81][10]/P0001 ,
		_w12950_,
		_w30751_
	);
	LUT2 #(
		.INIT('h8)
	) name20240 (
		\wishbone_bd_ram_mem1_reg[183][10]/P0001 ,
		_w12787_,
		_w30752_
	);
	LUT2 #(
		.INIT('h8)
	) name20241 (
		\wishbone_bd_ram_mem1_reg[250][10]/P0001 ,
		_w13128_,
		_w30753_
	);
	LUT2 #(
		.INIT('h8)
	) name20242 (
		\wishbone_bd_ram_mem1_reg[106][10]/P0001 ,
		_w12713_,
		_w30754_
	);
	LUT2 #(
		.INIT('h8)
	) name20243 (
		\wishbone_bd_ram_mem1_reg[212][10]/P0001 ,
		_w12796_,
		_w30755_
	);
	LUT2 #(
		.INIT('h8)
	) name20244 (
		\wishbone_bd_ram_mem1_reg[246][10]/P0001 ,
		_w13076_,
		_w30756_
	);
	LUT2 #(
		.INIT('h8)
	) name20245 (
		\wishbone_bd_ram_mem1_reg[181][10]/P0001 ,
		_w12828_,
		_w30757_
	);
	LUT2 #(
		.INIT('h8)
	) name20246 (
		\wishbone_bd_ram_mem1_reg[89][10]/P0001 ,
		_w12964_,
		_w30758_
	);
	LUT2 #(
		.INIT('h8)
	) name20247 (
		\wishbone_bd_ram_mem1_reg[218][10]/P0001 ,
		_w13206_,
		_w30759_
	);
	LUT2 #(
		.INIT('h8)
	) name20248 (
		\wishbone_bd_ram_mem1_reg[23][10]/P0001 ,
		_w13008_,
		_w30760_
	);
	LUT2 #(
		.INIT('h8)
	) name20249 (
		\wishbone_bd_ram_mem1_reg[11][10]/P0001 ,
		_w13194_,
		_w30761_
	);
	LUT2 #(
		.INIT('h8)
	) name20250 (
		\wishbone_bd_ram_mem1_reg[62][10]/P0001 ,
		_w12673_,
		_w30762_
	);
	LUT2 #(
		.INIT('h8)
	) name20251 (
		\wishbone_bd_ram_mem1_reg[75][10]/P0001 ,
		_w12826_,
		_w30763_
	);
	LUT2 #(
		.INIT('h8)
	) name20252 (
		\wishbone_bd_ram_mem1_reg[61][10]/P0001 ,
		_w12725_,
		_w30764_
	);
	LUT2 #(
		.INIT('h8)
	) name20253 (
		\wishbone_bd_ram_mem1_reg[211][10]/P0001 ,
		_w13166_,
		_w30765_
	);
	LUT2 #(
		.INIT('h8)
	) name20254 (
		\wishbone_bd_ram_mem1_reg[37][10]/P0001 ,
		_w13102_,
		_w30766_
	);
	LUT2 #(
		.INIT('h8)
	) name20255 (
		\wishbone_bd_ram_mem1_reg[57][10]/P0001 ,
		_w13116_,
		_w30767_
	);
	LUT2 #(
		.INIT('h8)
	) name20256 (
		\wishbone_bd_ram_mem1_reg[7][10]/P0001 ,
		_w12728_,
		_w30768_
	);
	LUT2 #(
		.INIT('h8)
	) name20257 (
		\wishbone_bd_ram_mem1_reg[108][10]/P0001 ,
		_w13156_,
		_w30769_
	);
	LUT2 #(
		.INIT('h8)
	) name20258 (
		\wishbone_bd_ram_mem1_reg[197][10]/P0001 ,
		_w12834_,
		_w30770_
	);
	LUT2 #(
		.INIT('h8)
	) name20259 (
		\wishbone_bd_ram_mem1_reg[36][10]/P0001 ,
		_w12800_,
		_w30771_
	);
	LUT2 #(
		.INIT('h8)
	) name20260 (
		\wishbone_bd_ram_mem1_reg[216][10]/P0001 ,
		_w13028_,
		_w30772_
	);
	LUT2 #(
		.INIT('h8)
	) name20261 (
		\wishbone_bd_ram_mem1_reg[26][10]/P0001 ,
		_w12699_,
		_w30773_
	);
	LUT2 #(
		.INIT('h8)
	) name20262 (
		\wishbone_bd_ram_mem1_reg[126][10]/P0001 ,
		_w13218_,
		_w30774_
	);
	LUT2 #(
		.INIT('h8)
	) name20263 (
		\wishbone_bd_ram_mem1_reg[207][10]/P0001 ,
		_w13180_,
		_w30775_
	);
	LUT2 #(
		.INIT('h8)
	) name20264 (
		\wishbone_bd_ram_mem1_reg[157][10]/P0001 ,
		_w12926_,
		_w30776_
	);
	LUT2 #(
		.INIT('h8)
	) name20265 (
		\wishbone_bd_ram_mem1_reg[19][10]/P0001 ,
		_w13012_,
		_w30777_
	);
	LUT2 #(
		.INIT('h8)
	) name20266 (
		\wishbone_bd_ram_mem1_reg[4][10]/P0001 ,
		_w12666_,
		_w30778_
	);
	LUT2 #(
		.INIT('h8)
	) name20267 (
		\wishbone_bd_ram_mem1_reg[190][10]/P0001 ,
		_w12858_,
		_w30779_
	);
	LUT2 #(
		.INIT('h8)
	) name20268 (
		\wishbone_bd_ram_mem1_reg[213][10]/P0001 ,
		_w13002_,
		_w30780_
	);
	LUT2 #(
		.INIT('h8)
	) name20269 (
		\wishbone_bd_ram_mem1_reg[101][10]/P0001 ,
		_w13192_,
		_w30781_
	);
	LUT2 #(
		.INIT('h8)
	) name20270 (
		\wishbone_bd_ram_mem1_reg[97][10]/P0001 ,
		_w13096_,
		_w30782_
	);
	LUT2 #(
		.INIT('h8)
	) name20271 (
		\wishbone_bd_ram_mem1_reg[16][10]/P0001 ,
		_w13140_,
		_w30783_
	);
	LUT2 #(
		.INIT('h8)
	) name20272 (
		\wishbone_bd_ram_mem1_reg[201][10]/P0001 ,
		_w12822_,
		_w30784_
	);
	LUT2 #(
		.INIT('h8)
	) name20273 (
		\wishbone_bd_ram_mem1_reg[59][10]/P0001 ,
		_w12780_,
		_w30785_
	);
	LUT2 #(
		.INIT('h8)
	) name20274 (
		\wishbone_bd_ram_mem1_reg[117][10]/P0001 ,
		_w12715_,
		_w30786_
	);
	LUT2 #(
		.INIT('h8)
	) name20275 (
		\wishbone_bd_ram_mem1_reg[142][10]/P0001 ,
		_w12928_,
		_w30787_
	);
	LUT2 #(
		.INIT('h8)
	) name20276 (
		\wishbone_bd_ram_mem1_reg[154][10]/P0001 ,
		_w12962_,
		_w30788_
	);
	LUT2 #(
		.INIT('h8)
	) name20277 (
		\wishbone_bd_ram_mem1_reg[156][10]/P0001 ,
		_w13190_,
		_w30789_
	);
	LUT2 #(
		.INIT('h8)
	) name20278 (
		\wishbone_bd_ram_mem1_reg[15][10]/P0001 ,
		_w13210_,
		_w30790_
	);
	LUT2 #(
		.INIT('h8)
	) name20279 (
		\wishbone_bd_ram_mem1_reg[5][10]/P0001 ,
		_w12878_,
		_w30791_
	);
	LUT2 #(
		.INIT('h8)
	) name20280 (
		\wishbone_bd_ram_mem1_reg[73][10]/P0001 ,
		_w12918_,
		_w30792_
	);
	LUT2 #(
		.INIT('h8)
	) name20281 (
		\wishbone_bd_ram_mem1_reg[114][10]/P0001 ,
		_w13202_,
		_w30793_
	);
	LUT2 #(
		.INIT('h8)
	) name20282 (
		\wishbone_bd_ram_mem1_reg[80][10]/P0001 ,
		_w12689_,
		_w30794_
	);
	LUT2 #(
		.INIT('h8)
	) name20283 (
		\wishbone_bd_ram_mem1_reg[138][10]/P0001 ,
		_w12958_,
		_w30795_
	);
	LUT2 #(
		.INIT('h8)
	) name20284 (
		\wishbone_bd_ram_mem1_reg[224][10]/P0001 ,
		_w12902_,
		_w30796_
	);
	LUT2 #(
		.INIT('h8)
	) name20285 (
		\wishbone_bd_ram_mem1_reg[174][10]/P0001 ,
		_w12972_,
		_w30797_
	);
	LUT2 #(
		.INIT('h8)
	) name20286 (
		\wishbone_bd_ram_mem1_reg[123][10]/P0001 ,
		_w13114_,
		_w30798_
	);
	LUT2 #(
		.INIT('h8)
	) name20287 (
		\wishbone_bd_ram_mem1_reg[152][10]/P0001 ,
		_w12966_,
		_w30799_
	);
	LUT2 #(
		.INIT('h8)
	) name20288 (
		\wishbone_bd_ram_mem1_reg[69][10]/P0001 ,
		_w12738_,
		_w30800_
	);
	LUT2 #(
		.INIT('h8)
	) name20289 (
		\wishbone_bd_ram_mem1_reg[68][10]/P0001 ,
		_w12946_,
		_w30801_
	);
	LUT2 #(
		.INIT('h8)
	) name20290 (
		\wishbone_bd_ram_mem1_reg[147][10]/P0001 ,
		_w13146_,
		_w30802_
	);
	LUT2 #(
		.INIT('h8)
	) name20291 (
		\wishbone_bd_ram_mem1_reg[167][10]/P0001 ,
		_w12986_,
		_w30803_
	);
	LUT2 #(
		.INIT('h8)
	) name20292 (
		\wishbone_bd_ram_mem1_reg[202][10]/P0001 ,
		_w12870_,
		_w30804_
	);
	LUT2 #(
		.INIT('h8)
	) name20293 (
		\wishbone_bd_ram_mem1_reg[115][10]/P0001 ,
		_w13112_,
		_w30805_
	);
	LUT2 #(
		.INIT('h8)
	) name20294 (
		\wishbone_bd_ram_mem1_reg[98][10]/P0001 ,
		_w12816_,
		_w30806_
	);
	LUT2 #(
		.INIT('h8)
	) name20295 (
		\wishbone_bd_ram_mem1_reg[237][10]/P0001 ,
		_w12990_,
		_w30807_
	);
	LUT2 #(
		.INIT('h8)
	) name20296 (
		\wishbone_bd_ram_mem1_reg[234][10]/P0001 ,
		_w13214_,
		_w30808_
	);
	LUT2 #(
		.INIT('h8)
	) name20297 (
		\wishbone_bd_ram_mem1_reg[47][10]/P0001 ,
		_w12904_,
		_w30809_
	);
	LUT2 #(
		.INIT('h8)
	) name20298 (
		\wishbone_bd_ram_mem1_reg[203][10]/P0001 ,
		_w13158_,
		_w30810_
	);
	LUT2 #(
		.INIT('h8)
	) name20299 (
		\wishbone_bd_ram_mem1_reg[121][10]/P0001 ,
		_w13078_,
		_w30811_
	);
	LUT2 #(
		.INIT('h8)
	) name20300 (
		\wishbone_bd_ram_mem1_reg[209][10]/P0001 ,
		_w13152_,
		_w30812_
	);
	LUT2 #(
		.INIT('h8)
	) name20301 (
		\wishbone_bd_ram_mem1_reg[91][10]/P0001 ,
		_w13074_,
		_w30813_
	);
	LUT2 #(
		.INIT('h8)
	) name20302 (
		\wishbone_bd_ram_mem1_reg[229][10]/P0001 ,
		_w12711_,
		_w30814_
	);
	LUT2 #(
		.INIT('h8)
	) name20303 (
		\wishbone_bd_ram_mem1_reg[170][10]/P0001 ,
		_w13030_,
		_w30815_
	);
	LUT2 #(
		.INIT('h8)
	) name20304 (
		\wishbone_bd_ram_mem1_reg[53][10]/P0001 ,
		_w13020_,
		_w30816_
	);
	LUT2 #(
		.INIT('h8)
	) name20305 (
		\wishbone_bd_ram_mem1_reg[185][10]/P0001 ,
		_w12940_,
		_w30817_
	);
	LUT2 #(
		.INIT('h8)
	) name20306 (
		\wishbone_bd_ram_mem1_reg[1][10]/P0001 ,
		_w13014_,
		_w30818_
	);
	LUT2 #(
		.INIT('h8)
	) name20307 (
		\wishbone_bd_ram_mem1_reg[135][10]/P0001 ,
		_w13124_,
		_w30819_
	);
	LUT2 #(
		.INIT('h8)
	) name20308 (
		\wishbone_bd_ram_mem1_reg[104][10]/P0001 ,
		_w13148_,
		_w30820_
	);
	LUT2 #(
		.INIT('h8)
	) name20309 (
		\wishbone_bd_ram_mem1_reg[176][10]/P0001 ,
		_w12868_,
		_w30821_
	);
	LUT2 #(
		.INIT('h8)
	) name20310 (
		\wishbone_bd_ram_mem1_reg[217][10]/P0001 ,
		_w13188_,
		_w30822_
	);
	LUT2 #(
		.INIT('h8)
	) name20311 (
		\wishbone_bd_ram_mem1_reg[87][10]/P0001 ,
		_w13154_,
		_w30823_
	);
	LUT2 #(
		.INIT('h8)
	) name20312 (
		\wishbone_bd_ram_mem1_reg[238][10]/P0001 ,
		_w13160_,
		_w30824_
	);
	LUT2 #(
		.INIT('h8)
	) name20313 (
		\wishbone_bd_ram_mem1_reg[55][10]/P0001 ,
		_w12785_,
		_w30825_
	);
	LUT2 #(
		.INIT('h8)
	) name20314 (
		\wishbone_bd_ram_mem1_reg[94][10]/P0001 ,
		_w13186_,
		_w30826_
	);
	LUT2 #(
		.INIT('h8)
	) name20315 (
		\wishbone_bd_ram_mem1_reg[50][10]/P0001 ,
		_w13150_,
		_w30827_
	);
	LUT2 #(
		.INIT('h8)
	) name20316 (
		\wishbone_bd_ram_mem1_reg[67][10]/P0001 ,
		_w13134_,
		_w30828_
	);
	LUT2 #(
		.INIT('h8)
	) name20317 (
		\wishbone_bd_ram_mem1_reg[84][10]/P0001 ,
		_w12934_,
		_w30829_
	);
	LUT2 #(
		.INIT('h8)
	) name20318 (
		\wishbone_bd_ram_mem1_reg[232][10]/P0001 ,
		_w12758_,
		_w30830_
	);
	LUT2 #(
		.INIT('h8)
	) name20319 (
		\wishbone_bd_ram_mem1_reg[46][10]/P0001 ,
		_w12884_,
		_w30831_
	);
	LUT2 #(
		.INIT('h8)
	) name20320 (
		\wishbone_bd_ram_mem1_reg[74][10]/P0001 ,
		_w12812_,
		_w30832_
	);
	LUT2 #(
		.INIT('h8)
	) name20321 (
		\wishbone_bd_ram_mem1_reg[214][10]/P0001 ,
		_w12984_,
		_w30833_
	);
	LUT2 #(
		.INIT('h8)
	) name20322 (
		\wishbone_bd_ram_mem1_reg[166][10]/P0001 ,
		_w13040_,
		_w30834_
	);
	LUT2 #(
		.INIT('h8)
	) name20323 (
		\wishbone_bd_ram_mem1_reg[95][10]/P0001 ,
		_w12844_,
		_w30835_
	);
	LUT2 #(
		.INIT('h8)
	) name20324 (
		\wishbone_bd_ram_mem1_reg[178][10]/P0001 ,
		_w12886_,
		_w30836_
	);
	LUT2 #(
		.INIT('h8)
	) name20325 (
		\wishbone_bd_ram_mem1_reg[25][10]/P0001 ,
		_w13108_,
		_w30837_
	);
	LUT2 #(
		.INIT('h8)
	) name20326 (
		\wishbone_bd_ram_mem1_reg[171][10]/P0001 ,
		_w12910_,
		_w30838_
	);
	LUT2 #(
		.INIT('h8)
	) name20327 (
		\wishbone_bd_ram_mem1_reg[72][10]/P0001 ,
		_w12810_,
		_w30839_
	);
	LUT2 #(
		.INIT('h8)
	) name20328 (
		\wishbone_bd_ram_mem1_reg[221][10]/P0001 ,
		_w12802_,
		_w30840_
	);
	LUT2 #(
		.INIT('h8)
	) name20329 (
		\wishbone_bd_ram_mem1_reg[227][10]/P0001 ,
		_w12936_,
		_w30841_
	);
	LUT2 #(
		.INIT('h8)
	) name20330 (
		\wishbone_bd_ram_mem1_reg[182][10]/P0001 ,
		_w12820_,
		_w30842_
	);
	LUT2 #(
		.INIT('h8)
	) name20331 (
		\wishbone_bd_ram_mem1_reg[9][10]/P0001 ,
		_w12808_,
		_w30843_
	);
	LUT2 #(
		.INIT('h8)
	) name20332 (
		\wishbone_bd_ram_mem1_reg[110][10]/P0001 ,
		_w13046_,
		_w30844_
	);
	LUT2 #(
		.INIT('h8)
	) name20333 (
		\wishbone_bd_ram_mem1_reg[85][10]/P0001 ,
		_w13216_,
		_w30845_
	);
	LUT2 #(
		.INIT('h8)
	) name20334 (
		\wishbone_bd_ram_mem1_reg[168][10]/P0001 ,
		_w13208_,
		_w30846_
	);
	LUT2 #(
		.INIT('h8)
	) name20335 (
		\wishbone_bd_ram_mem1_reg[143][10]/P0001 ,
		_w12922_,
		_w30847_
	);
	LUT2 #(
		.INIT('h8)
	) name20336 (
		\wishbone_bd_ram_mem1_reg[248][10]/P0001 ,
		_w12789_,
		_w30848_
	);
	LUT2 #(
		.INIT('h8)
	) name20337 (
		\wishbone_bd_ram_mem1_reg[51][10]/P0001 ,
		_w13024_,
		_w30849_
	);
	LUT2 #(
		.INIT('h8)
	) name20338 (
		\wishbone_bd_ram_mem1_reg[125][10]/P0001 ,
		_w12956_,
		_w30850_
	);
	LUT2 #(
		.INIT('h8)
	) name20339 (
		\wishbone_bd_ram_mem1_reg[153][10]/P0001 ,
		_w12890_,
		_w30851_
	);
	LUT2 #(
		.INIT('h8)
	) name20340 (
		\wishbone_bd_ram_mem1_reg[179][10]/P0001 ,
		_w13050_,
		_w30852_
	);
	LUT2 #(
		.INIT('h8)
	) name20341 (
		\wishbone_bd_ram_mem1_reg[129][10]/P0001 ,
		_w12776_,
		_w30853_
	);
	LUT2 #(
		.INIT('h8)
	) name20342 (
		\wishbone_bd_ram_mem1_reg[34][10]/P0001 ,
		_w12930_,
		_w30854_
	);
	LUT2 #(
		.INIT('h8)
	) name20343 (
		\wishbone_bd_ram_mem1_reg[198][10]/P0001 ,
		_w12832_,
		_w30855_
	);
	LUT2 #(
		.INIT('h8)
	) name20344 (
		\wishbone_bd_ram_mem1_reg[226][10]/P0001 ,
		_w13138_,
		_w30856_
	);
	LUT2 #(
		.INIT('h8)
	) name20345 (
		\wishbone_bd_ram_mem1_reg[244][10]/P0001 ,
		_w12747_,
		_w30857_
	);
	LUT2 #(
		.INIT('h8)
	) name20346 (
		\wishbone_bd_ram_mem1_reg[13][10]/P0001 ,
		_w13178_,
		_w30858_
	);
	LUT2 #(
		.INIT('h8)
	) name20347 (
		\wishbone_bd_ram_mem1_reg[45][10]/P0001 ,
		_w12908_,
		_w30859_
	);
	LUT2 #(
		.INIT('h8)
	) name20348 (
		\wishbone_bd_ram_mem1_reg[109][10]/P0001 ,
		_w12888_,
		_w30860_
	);
	LUT2 #(
		.INIT('h8)
	) name20349 (
		\wishbone_bd_ram_mem1_reg[63][10]/P0001 ,
		_w12850_,
		_w30861_
	);
	LUT2 #(
		.INIT('h8)
	) name20350 (
		\wishbone_bd_ram_mem1_reg[35][10]/P0001 ,
		_w12703_,
		_w30862_
	);
	LUT2 #(
		.INIT('h8)
	) name20351 (
		\wishbone_bd_ram_mem1_reg[173][10]/P0001 ,
		_w12854_,
		_w30863_
	);
	LUT2 #(
		.INIT('h8)
	) name20352 (
		\wishbone_bd_ram_mem1_reg[233][10]/P0001 ,
		_w12836_,
		_w30864_
	);
	LUT2 #(
		.INIT('h8)
	) name20353 (
		\wishbone_bd_ram_mem1_reg[40][10]/P0001 ,
		_w13132_,
		_w30865_
	);
	LUT2 #(
		.INIT('h8)
	) name20354 (
		\wishbone_bd_ram_mem1_reg[66][10]/P0001 ,
		_w12824_,
		_w30866_
	);
	LUT2 #(
		.INIT('h8)
	) name20355 (
		\wishbone_bd_ram_mem1_reg[192][10]/P0001 ,
		_w12938_,
		_w30867_
	);
	LUT2 #(
		.INIT('h8)
	) name20356 (
		\wishbone_bd_ram_mem1_reg[195][10]/P0001 ,
		_w13144_,
		_w30868_
	);
	LUT2 #(
		.INIT('h8)
	) name20357 (
		\wishbone_bd_ram_mem1_reg[160][10]/P0001 ,
		_w12872_,
		_w30869_
	);
	LUT2 #(
		.INIT('h8)
	) name20358 (
		\wishbone_bd_ram_mem1_reg[194][10]/P0001 ,
		_w12772_,
		_w30870_
	);
	LUT2 #(
		.INIT('h8)
	) name20359 (
		\wishbone_bd_ram_mem1_reg[231][10]/P0001 ,
		_w12856_,
		_w30871_
	);
	LUT2 #(
		.INIT('h8)
	) name20360 (
		\wishbone_bd_ram_mem1_reg[169][10]/P0001 ,
		_w12722_,
		_w30872_
	);
	LUT2 #(
		.INIT('h8)
	) name20361 (
		\wishbone_bd_ram_mem1_reg[105][10]/P0001 ,
		_w12751_,
		_w30873_
	);
	LUT2 #(
		.INIT('h8)
	) name20362 (
		\wishbone_bd_ram_mem1_reg[254][10]/P0001 ,
		_w12892_,
		_w30874_
	);
	LUT2 #(
		.INIT('h8)
	) name20363 (
		\wishbone_bd_ram_mem1_reg[6][10]/P0001 ,
		_w12968_,
		_w30875_
	);
	LUT2 #(
		.INIT('h8)
	) name20364 (
		\wishbone_bd_ram_mem1_reg[2][10]/P0001 ,
		_w13088_,
		_w30876_
	);
	LUT2 #(
		.INIT('h8)
	) name20365 (
		\wishbone_bd_ram_mem1_reg[8][10]/P0001 ,
		_w12920_,
		_w30877_
	);
	LUT2 #(
		.INIT('h8)
	) name20366 (
		\wishbone_bd_ram_mem1_reg[205][10]/P0001 ,
		_w13068_,
		_w30878_
	);
	LUT2 #(
		.INIT('h8)
	) name20367 (
		\wishbone_bd_ram_mem1_reg[150][10]/P0001 ,
		_w13136_,
		_w30879_
	);
	LUT2 #(
		.INIT('h8)
	) name20368 (
		\wishbone_bd_ram_mem1_reg[239][10]/P0001 ,
		_w12862_,
		_w30880_
	);
	LUT2 #(
		.INIT('h8)
	) name20369 (
		\wishbone_bd_ram_mem1_reg[172][10]/P0001 ,
		_w12944_,
		_w30881_
	);
	LUT2 #(
		.INIT('h8)
	) name20370 (
		\wishbone_bd_ram_mem1_reg[130][10]/P0001 ,
		_w12914_,
		_w30882_
	);
	LUT2 #(
		.INIT('h8)
	) name20371 (
		\wishbone_bd_ram_mem1_reg[186][10]/P0001 ,
		_w12783_,
		_w30883_
	);
	LUT2 #(
		.INIT('h8)
	) name20372 (
		\wishbone_bd_ram_mem1_reg[223][10]/P0001 ,
		_w12838_,
		_w30884_
	);
	LUT2 #(
		.INIT('h8)
	) name20373 (
		\wishbone_bd_ram_mem1_reg[144][10]/P0001 ,
		_w12756_,
		_w30885_
	);
	LUT2 #(
		.INIT('h1)
	) name20374 (
		_w30630_,
		_w30631_,
		_w30886_
	);
	LUT2 #(
		.INIT('h1)
	) name20375 (
		_w30632_,
		_w30633_,
		_w30887_
	);
	LUT2 #(
		.INIT('h1)
	) name20376 (
		_w30634_,
		_w30635_,
		_w30888_
	);
	LUT2 #(
		.INIT('h1)
	) name20377 (
		_w30636_,
		_w30637_,
		_w30889_
	);
	LUT2 #(
		.INIT('h1)
	) name20378 (
		_w30638_,
		_w30639_,
		_w30890_
	);
	LUT2 #(
		.INIT('h1)
	) name20379 (
		_w30640_,
		_w30641_,
		_w30891_
	);
	LUT2 #(
		.INIT('h1)
	) name20380 (
		_w30642_,
		_w30643_,
		_w30892_
	);
	LUT2 #(
		.INIT('h1)
	) name20381 (
		_w30644_,
		_w30645_,
		_w30893_
	);
	LUT2 #(
		.INIT('h1)
	) name20382 (
		_w30646_,
		_w30647_,
		_w30894_
	);
	LUT2 #(
		.INIT('h1)
	) name20383 (
		_w30648_,
		_w30649_,
		_w30895_
	);
	LUT2 #(
		.INIT('h1)
	) name20384 (
		_w30650_,
		_w30651_,
		_w30896_
	);
	LUT2 #(
		.INIT('h1)
	) name20385 (
		_w30652_,
		_w30653_,
		_w30897_
	);
	LUT2 #(
		.INIT('h1)
	) name20386 (
		_w30654_,
		_w30655_,
		_w30898_
	);
	LUT2 #(
		.INIT('h1)
	) name20387 (
		_w30656_,
		_w30657_,
		_w30899_
	);
	LUT2 #(
		.INIT('h1)
	) name20388 (
		_w30658_,
		_w30659_,
		_w30900_
	);
	LUT2 #(
		.INIT('h1)
	) name20389 (
		_w30660_,
		_w30661_,
		_w30901_
	);
	LUT2 #(
		.INIT('h1)
	) name20390 (
		_w30662_,
		_w30663_,
		_w30902_
	);
	LUT2 #(
		.INIT('h1)
	) name20391 (
		_w30664_,
		_w30665_,
		_w30903_
	);
	LUT2 #(
		.INIT('h1)
	) name20392 (
		_w30666_,
		_w30667_,
		_w30904_
	);
	LUT2 #(
		.INIT('h1)
	) name20393 (
		_w30668_,
		_w30669_,
		_w30905_
	);
	LUT2 #(
		.INIT('h1)
	) name20394 (
		_w30670_,
		_w30671_,
		_w30906_
	);
	LUT2 #(
		.INIT('h1)
	) name20395 (
		_w30672_,
		_w30673_,
		_w30907_
	);
	LUT2 #(
		.INIT('h1)
	) name20396 (
		_w30674_,
		_w30675_,
		_w30908_
	);
	LUT2 #(
		.INIT('h1)
	) name20397 (
		_w30676_,
		_w30677_,
		_w30909_
	);
	LUT2 #(
		.INIT('h1)
	) name20398 (
		_w30678_,
		_w30679_,
		_w30910_
	);
	LUT2 #(
		.INIT('h1)
	) name20399 (
		_w30680_,
		_w30681_,
		_w30911_
	);
	LUT2 #(
		.INIT('h1)
	) name20400 (
		_w30682_,
		_w30683_,
		_w30912_
	);
	LUT2 #(
		.INIT('h1)
	) name20401 (
		_w30684_,
		_w30685_,
		_w30913_
	);
	LUT2 #(
		.INIT('h1)
	) name20402 (
		_w30686_,
		_w30687_,
		_w30914_
	);
	LUT2 #(
		.INIT('h1)
	) name20403 (
		_w30688_,
		_w30689_,
		_w30915_
	);
	LUT2 #(
		.INIT('h1)
	) name20404 (
		_w30690_,
		_w30691_,
		_w30916_
	);
	LUT2 #(
		.INIT('h1)
	) name20405 (
		_w30692_,
		_w30693_,
		_w30917_
	);
	LUT2 #(
		.INIT('h1)
	) name20406 (
		_w30694_,
		_w30695_,
		_w30918_
	);
	LUT2 #(
		.INIT('h1)
	) name20407 (
		_w30696_,
		_w30697_,
		_w30919_
	);
	LUT2 #(
		.INIT('h1)
	) name20408 (
		_w30698_,
		_w30699_,
		_w30920_
	);
	LUT2 #(
		.INIT('h1)
	) name20409 (
		_w30700_,
		_w30701_,
		_w30921_
	);
	LUT2 #(
		.INIT('h1)
	) name20410 (
		_w30702_,
		_w30703_,
		_w30922_
	);
	LUT2 #(
		.INIT('h1)
	) name20411 (
		_w30704_,
		_w30705_,
		_w30923_
	);
	LUT2 #(
		.INIT('h1)
	) name20412 (
		_w30706_,
		_w30707_,
		_w30924_
	);
	LUT2 #(
		.INIT('h1)
	) name20413 (
		_w30708_,
		_w30709_,
		_w30925_
	);
	LUT2 #(
		.INIT('h1)
	) name20414 (
		_w30710_,
		_w30711_,
		_w30926_
	);
	LUT2 #(
		.INIT('h1)
	) name20415 (
		_w30712_,
		_w30713_,
		_w30927_
	);
	LUT2 #(
		.INIT('h1)
	) name20416 (
		_w30714_,
		_w30715_,
		_w30928_
	);
	LUT2 #(
		.INIT('h1)
	) name20417 (
		_w30716_,
		_w30717_,
		_w30929_
	);
	LUT2 #(
		.INIT('h1)
	) name20418 (
		_w30718_,
		_w30719_,
		_w30930_
	);
	LUT2 #(
		.INIT('h1)
	) name20419 (
		_w30720_,
		_w30721_,
		_w30931_
	);
	LUT2 #(
		.INIT('h1)
	) name20420 (
		_w30722_,
		_w30723_,
		_w30932_
	);
	LUT2 #(
		.INIT('h1)
	) name20421 (
		_w30724_,
		_w30725_,
		_w30933_
	);
	LUT2 #(
		.INIT('h1)
	) name20422 (
		_w30726_,
		_w30727_,
		_w30934_
	);
	LUT2 #(
		.INIT('h1)
	) name20423 (
		_w30728_,
		_w30729_,
		_w30935_
	);
	LUT2 #(
		.INIT('h1)
	) name20424 (
		_w30730_,
		_w30731_,
		_w30936_
	);
	LUT2 #(
		.INIT('h1)
	) name20425 (
		_w30732_,
		_w30733_,
		_w30937_
	);
	LUT2 #(
		.INIT('h1)
	) name20426 (
		_w30734_,
		_w30735_,
		_w30938_
	);
	LUT2 #(
		.INIT('h1)
	) name20427 (
		_w30736_,
		_w30737_,
		_w30939_
	);
	LUT2 #(
		.INIT('h1)
	) name20428 (
		_w30738_,
		_w30739_,
		_w30940_
	);
	LUT2 #(
		.INIT('h1)
	) name20429 (
		_w30740_,
		_w30741_,
		_w30941_
	);
	LUT2 #(
		.INIT('h1)
	) name20430 (
		_w30742_,
		_w30743_,
		_w30942_
	);
	LUT2 #(
		.INIT('h1)
	) name20431 (
		_w30744_,
		_w30745_,
		_w30943_
	);
	LUT2 #(
		.INIT('h1)
	) name20432 (
		_w30746_,
		_w30747_,
		_w30944_
	);
	LUT2 #(
		.INIT('h1)
	) name20433 (
		_w30748_,
		_w30749_,
		_w30945_
	);
	LUT2 #(
		.INIT('h1)
	) name20434 (
		_w30750_,
		_w30751_,
		_w30946_
	);
	LUT2 #(
		.INIT('h1)
	) name20435 (
		_w30752_,
		_w30753_,
		_w30947_
	);
	LUT2 #(
		.INIT('h1)
	) name20436 (
		_w30754_,
		_w30755_,
		_w30948_
	);
	LUT2 #(
		.INIT('h1)
	) name20437 (
		_w30756_,
		_w30757_,
		_w30949_
	);
	LUT2 #(
		.INIT('h1)
	) name20438 (
		_w30758_,
		_w30759_,
		_w30950_
	);
	LUT2 #(
		.INIT('h1)
	) name20439 (
		_w30760_,
		_w30761_,
		_w30951_
	);
	LUT2 #(
		.INIT('h1)
	) name20440 (
		_w30762_,
		_w30763_,
		_w30952_
	);
	LUT2 #(
		.INIT('h1)
	) name20441 (
		_w30764_,
		_w30765_,
		_w30953_
	);
	LUT2 #(
		.INIT('h1)
	) name20442 (
		_w30766_,
		_w30767_,
		_w30954_
	);
	LUT2 #(
		.INIT('h1)
	) name20443 (
		_w30768_,
		_w30769_,
		_w30955_
	);
	LUT2 #(
		.INIT('h1)
	) name20444 (
		_w30770_,
		_w30771_,
		_w30956_
	);
	LUT2 #(
		.INIT('h1)
	) name20445 (
		_w30772_,
		_w30773_,
		_w30957_
	);
	LUT2 #(
		.INIT('h1)
	) name20446 (
		_w30774_,
		_w30775_,
		_w30958_
	);
	LUT2 #(
		.INIT('h1)
	) name20447 (
		_w30776_,
		_w30777_,
		_w30959_
	);
	LUT2 #(
		.INIT('h1)
	) name20448 (
		_w30778_,
		_w30779_,
		_w30960_
	);
	LUT2 #(
		.INIT('h1)
	) name20449 (
		_w30780_,
		_w30781_,
		_w30961_
	);
	LUT2 #(
		.INIT('h1)
	) name20450 (
		_w30782_,
		_w30783_,
		_w30962_
	);
	LUT2 #(
		.INIT('h1)
	) name20451 (
		_w30784_,
		_w30785_,
		_w30963_
	);
	LUT2 #(
		.INIT('h1)
	) name20452 (
		_w30786_,
		_w30787_,
		_w30964_
	);
	LUT2 #(
		.INIT('h1)
	) name20453 (
		_w30788_,
		_w30789_,
		_w30965_
	);
	LUT2 #(
		.INIT('h1)
	) name20454 (
		_w30790_,
		_w30791_,
		_w30966_
	);
	LUT2 #(
		.INIT('h1)
	) name20455 (
		_w30792_,
		_w30793_,
		_w30967_
	);
	LUT2 #(
		.INIT('h1)
	) name20456 (
		_w30794_,
		_w30795_,
		_w30968_
	);
	LUT2 #(
		.INIT('h1)
	) name20457 (
		_w30796_,
		_w30797_,
		_w30969_
	);
	LUT2 #(
		.INIT('h1)
	) name20458 (
		_w30798_,
		_w30799_,
		_w30970_
	);
	LUT2 #(
		.INIT('h1)
	) name20459 (
		_w30800_,
		_w30801_,
		_w30971_
	);
	LUT2 #(
		.INIT('h1)
	) name20460 (
		_w30802_,
		_w30803_,
		_w30972_
	);
	LUT2 #(
		.INIT('h1)
	) name20461 (
		_w30804_,
		_w30805_,
		_w30973_
	);
	LUT2 #(
		.INIT('h1)
	) name20462 (
		_w30806_,
		_w30807_,
		_w30974_
	);
	LUT2 #(
		.INIT('h1)
	) name20463 (
		_w30808_,
		_w30809_,
		_w30975_
	);
	LUT2 #(
		.INIT('h1)
	) name20464 (
		_w30810_,
		_w30811_,
		_w30976_
	);
	LUT2 #(
		.INIT('h1)
	) name20465 (
		_w30812_,
		_w30813_,
		_w30977_
	);
	LUT2 #(
		.INIT('h1)
	) name20466 (
		_w30814_,
		_w30815_,
		_w30978_
	);
	LUT2 #(
		.INIT('h1)
	) name20467 (
		_w30816_,
		_w30817_,
		_w30979_
	);
	LUT2 #(
		.INIT('h1)
	) name20468 (
		_w30818_,
		_w30819_,
		_w30980_
	);
	LUT2 #(
		.INIT('h1)
	) name20469 (
		_w30820_,
		_w30821_,
		_w30981_
	);
	LUT2 #(
		.INIT('h1)
	) name20470 (
		_w30822_,
		_w30823_,
		_w30982_
	);
	LUT2 #(
		.INIT('h1)
	) name20471 (
		_w30824_,
		_w30825_,
		_w30983_
	);
	LUT2 #(
		.INIT('h1)
	) name20472 (
		_w30826_,
		_w30827_,
		_w30984_
	);
	LUT2 #(
		.INIT('h1)
	) name20473 (
		_w30828_,
		_w30829_,
		_w30985_
	);
	LUT2 #(
		.INIT('h1)
	) name20474 (
		_w30830_,
		_w30831_,
		_w30986_
	);
	LUT2 #(
		.INIT('h1)
	) name20475 (
		_w30832_,
		_w30833_,
		_w30987_
	);
	LUT2 #(
		.INIT('h1)
	) name20476 (
		_w30834_,
		_w30835_,
		_w30988_
	);
	LUT2 #(
		.INIT('h1)
	) name20477 (
		_w30836_,
		_w30837_,
		_w30989_
	);
	LUT2 #(
		.INIT('h1)
	) name20478 (
		_w30838_,
		_w30839_,
		_w30990_
	);
	LUT2 #(
		.INIT('h1)
	) name20479 (
		_w30840_,
		_w30841_,
		_w30991_
	);
	LUT2 #(
		.INIT('h1)
	) name20480 (
		_w30842_,
		_w30843_,
		_w30992_
	);
	LUT2 #(
		.INIT('h1)
	) name20481 (
		_w30844_,
		_w30845_,
		_w30993_
	);
	LUT2 #(
		.INIT('h1)
	) name20482 (
		_w30846_,
		_w30847_,
		_w30994_
	);
	LUT2 #(
		.INIT('h1)
	) name20483 (
		_w30848_,
		_w30849_,
		_w30995_
	);
	LUT2 #(
		.INIT('h1)
	) name20484 (
		_w30850_,
		_w30851_,
		_w30996_
	);
	LUT2 #(
		.INIT('h1)
	) name20485 (
		_w30852_,
		_w30853_,
		_w30997_
	);
	LUT2 #(
		.INIT('h1)
	) name20486 (
		_w30854_,
		_w30855_,
		_w30998_
	);
	LUT2 #(
		.INIT('h1)
	) name20487 (
		_w30856_,
		_w30857_,
		_w30999_
	);
	LUT2 #(
		.INIT('h1)
	) name20488 (
		_w30858_,
		_w30859_,
		_w31000_
	);
	LUT2 #(
		.INIT('h1)
	) name20489 (
		_w30860_,
		_w30861_,
		_w31001_
	);
	LUT2 #(
		.INIT('h1)
	) name20490 (
		_w30862_,
		_w30863_,
		_w31002_
	);
	LUT2 #(
		.INIT('h1)
	) name20491 (
		_w30864_,
		_w30865_,
		_w31003_
	);
	LUT2 #(
		.INIT('h1)
	) name20492 (
		_w30866_,
		_w30867_,
		_w31004_
	);
	LUT2 #(
		.INIT('h1)
	) name20493 (
		_w30868_,
		_w30869_,
		_w31005_
	);
	LUT2 #(
		.INIT('h1)
	) name20494 (
		_w30870_,
		_w30871_,
		_w31006_
	);
	LUT2 #(
		.INIT('h1)
	) name20495 (
		_w30872_,
		_w30873_,
		_w31007_
	);
	LUT2 #(
		.INIT('h1)
	) name20496 (
		_w30874_,
		_w30875_,
		_w31008_
	);
	LUT2 #(
		.INIT('h1)
	) name20497 (
		_w30876_,
		_w30877_,
		_w31009_
	);
	LUT2 #(
		.INIT('h1)
	) name20498 (
		_w30878_,
		_w30879_,
		_w31010_
	);
	LUT2 #(
		.INIT('h1)
	) name20499 (
		_w30880_,
		_w30881_,
		_w31011_
	);
	LUT2 #(
		.INIT('h1)
	) name20500 (
		_w30882_,
		_w30883_,
		_w31012_
	);
	LUT2 #(
		.INIT('h1)
	) name20501 (
		_w30884_,
		_w30885_,
		_w31013_
	);
	LUT2 #(
		.INIT('h8)
	) name20502 (
		_w31012_,
		_w31013_,
		_w31014_
	);
	LUT2 #(
		.INIT('h8)
	) name20503 (
		_w31010_,
		_w31011_,
		_w31015_
	);
	LUT2 #(
		.INIT('h8)
	) name20504 (
		_w31008_,
		_w31009_,
		_w31016_
	);
	LUT2 #(
		.INIT('h8)
	) name20505 (
		_w31006_,
		_w31007_,
		_w31017_
	);
	LUT2 #(
		.INIT('h8)
	) name20506 (
		_w31004_,
		_w31005_,
		_w31018_
	);
	LUT2 #(
		.INIT('h8)
	) name20507 (
		_w31002_,
		_w31003_,
		_w31019_
	);
	LUT2 #(
		.INIT('h8)
	) name20508 (
		_w31000_,
		_w31001_,
		_w31020_
	);
	LUT2 #(
		.INIT('h8)
	) name20509 (
		_w30998_,
		_w30999_,
		_w31021_
	);
	LUT2 #(
		.INIT('h8)
	) name20510 (
		_w30996_,
		_w30997_,
		_w31022_
	);
	LUT2 #(
		.INIT('h8)
	) name20511 (
		_w30994_,
		_w30995_,
		_w31023_
	);
	LUT2 #(
		.INIT('h8)
	) name20512 (
		_w30992_,
		_w30993_,
		_w31024_
	);
	LUT2 #(
		.INIT('h8)
	) name20513 (
		_w30990_,
		_w30991_,
		_w31025_
	);
	LUT2 #(
		.INIT('h8)
	) name20514 (
		_w30988_,
		_w30989_,
		_w31026_
	);
	LUT2 #(
		.INIT('h8)
	) name20515 (
		_w30986_,
		_w30987_,
		_w31027_
	);
	LUT2 #(
		.INIT('h8)
	) name20516 (
		_w30984_,
		_w30985_,
		_w31028_
	);
	LUT2 #(
		.INIT('h8)
	) name20517 (
		_w30982_,
		_w30983_,
		_w31029_
	);
	LUT2 #(
		.INIT('h8)
	) name20518 (
		_w30980_,
		_w30981_,
		_w31030_
	);
	LUT2 #(
		.INIT('h8)
	) name20519 (
		_w30978_,
		_w30979_,
		_w31031_
	);
	LUT2 #(
		.INIT('h8)
	) name20520 (
		_w30976_,
		_w30977_,
		_w31032_
	);
	LUT2 #(
		.INIT('h8)
	) name20521 (
		_w30974_,
		_w30975_,
		_w31033_
	);
	LUT2 #(
		.INIT('h8)
	) name20522 (
		_w30972_,
		_w30973_,
		_w31034_
	);
	LUT2 #(
		.INIT('h8)
	) name20523 (
		_w30970_,
		_w30971_,
		_w31035_
	);
	LUT2 #(
		.INIT('h8)
	) name20524 (
		_w30968_,
		_w30969_,
		_w31036_
	);
	LUT2 #(
		.INIT('h8)
	) name20525 (
		_w30966_,
		_w30967_,
		_w31037_
	);
	LUT2 #(
		.INIT('h8)
	) name20526 (
		_w30964_,
		_w30965_,
		_w31038_
	);
	LUT2 #(
		.INIT('h8)
	) name20527 (
		_w30962_,
		_w30963_,
		_w31039_
	);
	LUT2 #(
		.INIT('h8)
	) name20528 (
		_w30960_,
		_w30961_,
		_w31040_
	);
	LUT2 #(
		.INIT('h8)
	) name20529 (
		_w30958_,
		_w30959_,
		_w31041_
	);
	LUT2 #(
		.INIT('h8)
	) name20530 (
		_w30956_,
		_w30957_,
		_w31042_
	);
	LUT2 #(
		.INIT('h8)
	) name20531 (
		_w30954_,
		_w30955_,
		_w31043_
	);
	LUT2 #(
		.INIT('h8)
	) name20532 (
		_w30952_,
		_w30953_,
		_w31044_
	);
	LUT2 #(
		.INIT('h8)
	) name20533 (
		_w30950_,
		_w30951_,
		_w31045_
	);
	LUT2 #(
		.INIT('h8)
	) name20534 (
		_w30948_,
		_w30949_,
		_w31046_
	);
	LUT2 #(
		.INIT('h8)
	) name20535 (
		_w30946_,
		_w30947_,
		_w31047_
	);
	LUT2 #(
		.INIT('h8)
	) name20536 (
		_w30944_,
		_w30945_,
		_w31048_
	);
	LUT2 #(
		.INIT('h8)
	) name20537 (
		_w30942_,
		_w30943_,
		_w31049_
	);
	LUT2 #(
		.INIT('h8)
	) name20538 (
		_w30940_,
		_w30941_,
		_w31050_
	);
	LUT2 #(
		.INIT('h8)
	) name20539 (
		_w30938_,
		_w30939_,
		_w31051_
	);
	LUT2 #(
		.INIT('h8)
	) name20540 (
		_w30936_,
		_w30937_,
		_w31052_
	);
	LUT2 #(
		.INIT('h8)
	) name20541 (
		_w30934_,
		_w30935_,
		_w31053_
	);
	LUT2 #(
		.INIT('h8)
	) name20542 (
		_w30932_,
		_w30933_,
		_w31054_
	);
	LUT2 #(
		.INIT('h8)
	) name20543 (
		_w30930_,
		_w30931_,
		_w31055_
	);
	LUT2 #(
		.INIT('h8)
	) name20544 (
		_w30928_,
		_w30929_,
		_w31056_
	);
	LUT2 #(
		.INIT('h8)
	) name20545 (
		_w30926_,
		_w30927_,
		_w31057_
	);
	LUT2 #(
		.INIT('h8)
	) name20546 (
		_w30924_,
		_w30925_,
		_w31058_
	);
	LUT2 #(
		.INIT('h8)
	) name20547 (
		_w30922_,
		_w30923_,
		_w31059_
	);
	LUT2 #(
		.INIT('h8)
	) name20548 (
		_w30920_,
		_w30921_,
		_w31060_
	);
	LUT2 #(
		.INIT('h8)
	) name20549 (
		_w30918_,
		_w30919_,
		_w31061_
	);
	LUT2 #(
		.INIT('h8)
	) name20550 (
		_w30916_,
		_w30917_,
		_w31062_
	);
	LUT2 #(
		.INIT('h8)
	) name20551 (
		_w30914_,
		_w30915_,
		_w31063_
	);
	LUT2 #(
		.INIT('h8)
	) name20552 (
		_w30912_,
		_w30913_,
		_w31064_
	);
	LUT2 #(
		.INIT('h8)
	) name20553 (
		_w30910_,
		_w30911_,
		_w31065_
	);
	LUT2 #(
		.INIT('h8)
	) name20554 (
		_w30908_,
		_w30909_,
		_w31066_
	);
	LUT2 #(
		.INIT('h8)
	) name20555 (
		_w30906_,
		_w30907_,
		_w31067_
	);
	LUT2 #(
		.INIT('h8)
	) name20556 (
		_w30904_,
		_w30905_,
		_w31068_
	);
	LUT2 #(
		.INIT('h8)
	) name20557 (
		_w30902_,
		_w30903_,
		_w31069_
	);
	LUT2 #(
		.INIT('h8)
	) name20558 (
		_w30900_,
		_w30901_,
		_w31070_
	);
	LUT2 #(
		.INIT('h8)
	) name20559 (
		_w30898_,
		_w30899_,
		_w31071_
	);
	LUT2 #(
		.INIT('h8)
	) name20560 (
		_w30896_,
		_w30897_,
		_w31072_
	);
	LUT2 #(
		.INIT('h8)
	) name20561 (
		_w30894_,
		_w30895_,
		_w31073_
	);
	LUT2 #(
		.INIT('h8)
	) name20562 (
		_w30892_,
		_w30893_,
		_w31074_
	);
	LUT2 #(
		.INIT('h8)
	) name20563 (
		_w30890_,
		_w30891_,
		_w31075_
	);
	LUT2 #(
		.INIT('h8)
	) name20564 (
		_w30888_,
		_w30889_,
		_w31076_
	);
	LUT2 #(
		.INIT('h8)
	) name20565 (
		_w30886_,
		_w30887_,
		_w31077_
	);
	LUT2 #(
		.INIT('h8)
	) name20566 (
		_w31076_,
		_w31077_,
		_w31078_
	);
	LUT2 #(
		.INIT('h8)
	) name20567 (
		_w31074_,
		_w31075_,
		_w31079_
	);
	LUT2 #(
		.INIT('h8)
	) name20568 (
		_w31072_,
		_w31073_,
		_w31080_
	);
	LUT2 #(
		.INIT('h8)
	) name20569 (
		_w31070_,
		_w31071_,
		_w31081_
	);
	LUT2 #(
		.INIT('h8)
	) name20570 (
		_w31068_,
		_w31069_,
		_w31082_
	);
	LUT2 #(
		.INIT('h8)
	) name20571 (
		_w31066_,
		_w31067_,
		_w31083_
	);
	LUT2 #(
		.INIT('h8)
	) name20572 (
		_w31064_,
		_w31065_,
		_w31084_
	);
	LUT2 #(
		.INIT('h8)
	) name20573 (
		_w31062_,
		_w31063_,
		_w31085_
	);
	LUT2 #(
		.INIT('h8)
	) name20574 (
		_w31060_,
		_w31061_,
		_w31086_
	);
	LUT2 #(
		.INIT('h8)
	) name20575 (
		_w31058_,
		_w31059_,
		_w31087_
	);
	LUT2 #(
		.INIT('h8)
	) name20576 (
		_w31056_,
		_w31057_,
		_w31088_
	);
	LUT2 #(
		.INIT('h8)
	) name20577 (
		_w31054_,
		_w31055_,
		_w31089_
	);
	LUT2 #(
		.INIT('h8)
	) name20578 (
		_w31052_,
		_w31053_,
		_w31090_
	);
	LUT2 #(
		.INIT('h8)
	) name20579 (
		_w31050_,
		_w31051_,
		_w31091_
	);
	LUT2 #(
		.INIT('h8)
	) name20580 (
		_w31048_,
		_w31049_,
		_w31092_
	);
	LUT2 #(
		.INIT('h8)
	) name20581 (
		_w31046_,
		_w31047_,
		_w31093_
	);
	LUT2 #(
		.INIT('h8)
	) name20582 (
		_w31044_,
		_w31045_,
		_w31094_
	);
	LUT2 #(
		.INIT('h8)
	) name20583 (
		_w31042_,
		_w31043_,
		_w31095_
	);
	LUT2 #(
		.INIT('h8)
	) name20584 (
		_w31040_,
		_w31041_,
		_w31096_
	);
	LUT2 #(
		.INIT('h8)
	) name20585 (
		_w31038_,
		_w31039_,
		_w31097_
	);
	LUT2 #(
		.INIT('h8)
	) name20586 (
		_w31036_,
		_w31037_,
		_w31098_
	);
	LUT2 #(
		.INIT('h8)
	) name20587 (
		_w31034_,
		_w31035_,
		_w31099_
	);
	LUT2 #(
		.INIT('h8)
	) name20588 (
		_w31032_,
		_w31033_,
		_w31100_
	);
	LUT2 #(
		.INIT('h8)
	) name20589 (
		_w31030_,
		_w31031_,
		_w31101_
	);
	LUT2 #(
		.INIT('h8)
	) name20590 (
		_w31028_,
		_w31029_,
		_w31102_
	);
	LUT2 #(
		.INIT('h8)
	) name20591 (
		_w31026_,
		_w31027_,
		_w31103_
	);
	LUT2 #(
		.INIT('h8)
	) name20592 (
		_w31024_,
		_w31025_,
		_w31104_
	);
	LUT2 #(
		.INIT('h8)
	) name20593 (
		_w31022_,
		_w31023_,
		_w31105_
	);
	LUT2 #(
		.INIT('h8)
	) name20594 (
		_w31020_,
		_w31021_,
		_w31106_
	);
	LUT2 #(
		.INIT('h8)
	) name20595 (
		_w31018_,
		_w31019_,
		_w31107_
	);
	LUT2 #(
		.INIT('h8)
	) name20596 (
		_w31016_,
		_w31017_,
		_w31108_
	);
	LUT2 #(
		.INIT('h8)
	) name20597 (
		_w31014_,
		_w31015_,
		_w31109_
	);
	LUT2 #(
		.INIT('h8)
	) name20598 (
		_w31108_,
		_w31109_,
		_w31110_
	);
	LUT2 #(
		.INIT('h8)
	) name20599 (
		_w31106_,
		_w31107_,
		_w31111_
	);
	LUT2 #(
		.INIT('h8)
	) name20600 (
		_w31104_,
		_w31105_,
		_w31112_
	);
	LUT2 #(
		.INIT('h8)
	) name20601 (
		_w31102_,
		_w31103_,
		_w31113_
	);
	LUT2 #(
		.INIT('h8)
	) name20602 (
		_w31100_,
		_w31101_,
		_w31114_
	);
	LUT2 #(
		.INIT('h8)
	) name20603 (
		_w31098_,
		_w31099_,
		_w31115_
	);
	LUT2 #(
		.INIT('h8)
	) name20604 (
		_w31096_,
		_w31097_,
		_w31116_
	);
	LUT2 #(
		.INIT('h8)
	) name20605 (
		_w31094_,
		_w31095_,
		_w31117_
	);
	LUT2 #(
		.INIT('h8)
	) name20606 (
		_w31092_,
		_w31093_,
		_w31118_
	);
	LUT2 #(
		.INIT('h8)
	) name20607 (
		_w31090_,
		_w31091_,
		_w31119_
	);
	LUT2 #(
		.INIT('h8)
	) name20608 (
		_w31088_,
		_w31089_,
		_w31120_
	);
	LUT2 #(
		.INIT('h8)
	) name20609 (
		_w31086_,
		_w31087_,
		_w31121_
	);
	LUT2 #(
		.INIT('h8)
	) name20610 (
		_w31084_,
		_w31085_,
		_w31122_
	);
	LUT2 #(
		.INIT('h8)
	) name20611 (
		_w31082_,
		_w31083_,
		_w31123_
	);
	LUT2 #(
		.INIT('h8)
	) name20612 (
		_w31080_,
		_w31081_,
		_w31124_
	);
	LUT2 #(
		.INIT('h8)
	) name20613 (
		_w31078_,
		_w31079_,
		_w31125_
	);
	LUT2 #(
		.INIT('h8)
	) name20614 (
		_w31124_,
		_w31125_,
		_w31126_
	);
	LUT2 #(
		.INIT('h8)
	) name20615 (
		_w31122_,
		_w31123_,
		_w31127_
	);
	LUT2 #(
		.INIT('h8)
	) name20616 (
		_w31120_,
		_w31121_,
		_w31128_
	);
	LUT2 #(
		.INIT('h8)
	) name20617 (
		_w31118_,
		_w31119_,
		_w31129_
	);
	LUT2 #(
		.INIT('h8)
	) name20618 (
		_w31116_,
		_w31117_,
		_w31130_
	);
	LUT2 #(
		.INIT('h8)
	) name20619 (
		_w31114_,
		_w31115_,
		_w31131_
	);
	LUT2 #(
		.INIT('h8)
	) name20620 (
		_w31112_,
		_w31113_,
		_w31132_
	);
	LUT2 #(
		.INIT('h8)
	) name20621 (
		_w31110_,
		_w31111_,
		_w31133_
	);
	LUT2 #(
		.INIT('h8)
	) name20622 (
		_w31132_,
		_w31133_,
		_w31134_
	);
	LUT2 #(
		.INIT('h8)
	) name20623 (
		_w31130_,
		_w31131_,
		_w31135_
	);
	LUT2 #(
		.INIT('h8)
	) name20624 (
		_w31128_,
		_w31129_,
		_w31136_
	);
	LUT2 #(
		.INIT('h8)
	) name20625 (
		_w31126_,
		_w31127_,
		_w31137_
	);
	LUT2 #(
		.INIT('h8)
	) name20626 (
		_w31136_,
		_w31137_,
		_w31138_
	);
	LUT2 #(
		.INIT('h8)
	) name20627 (
		_w31134_,
		_w31135_,
		_w31139_
	);
	LUT2 #(
		.INIT('h8)
	) name20628 (
		_w31138_,
		_w31139_,
		_w31140_
	);
	LUT2 #(
		.INIT('h1)
	) name20629 (
		wb_rst_i_pad,
		_w31140_,
		_w31141_
	);
	LUT2 #(
		.INIT('h8)
	) name20630 (
		_w17883_,
		_w31141_,
		_w31142_
	);
	LUT2 #(
		.INIT('h1)
	) name20631 (
		_w30629_,
		_w31142_,
		_w31143_
	);
	LUT2 #(
		.INIT('h1)
	) name20632 (
		\wishbone_TxPointerMSB_reg[11]/NET0131 ,
		_w17894_,
		_w31144_
	);
	LUT2 #(
		.INIT('h1)
	) name20633 (
		_w17883_,
		_w17895_,
		_w31145_
	);
	LUT2 #(
		.INIT('h4)
	) name20634 (
		_w31144_,
		_w31145_,
		_w31146_
	);
	LUT2 #(
		.INIT('h8)
	) name20635 (
		_w17883_,
		_w27980_,
		_w31147_
	);
	LUT2 #(
		.INIT('h1)
	) name20636 (
		_w31146_,
		_w31147_,
		_w31148_
	);
	LUT2 #(
		.INIT('h1)
	) name20637 (
		\wishbone_TxPointerMSB_reg[13]/NET0131 ,
		_w17896_,
		_w31149_
	);
	LUT2 #(
		.INIT('h1)
	) name20638 (
		_w17883_,
		_w30557_,
		_w31150_
	);
	LUT2 #(
		.INIT('h4)
	) name20639 (
		_w31149_,
		_w31150_,
		_w31151_
	);
	LUT2 #(
		.INIT('h8)
	) name20640 (
		_w17883_,
		_w29947_,
		_w31152_
	);
	LUT2 #(
		.INIT('h1)
	) name20641 (
		_w31151_,
		_w31152_,
		_w31153_
	);
	LUT2 #(
		.INIT('h8)
	) name20642 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w17898_,
		_w31154_
	);
	LUT2 #(
		.INIT('h1)
	) name20643 (
		\wishbone_TxPointerMSB_reg[15]/NET0131 ,
		_w17898_,
		_w31155_
	);
	LUT2 #(
		.INIT('h1)
	) name20644 (
		_w17883_,
		_w31154_,
		_w31156_
	);
	LUT2 #(
		.INIT('h4)
	) name20645 (
		_w31155_,
		_w31156_,
		_w31157_
	);
	LUT2 #(
		.INIT('h8)
	) name20646 (
		_w15689_,
		_w17883_,
		_w31158_
	);
	LUT2 #(
		.INIT('h1)
	) name20647 (
		_w31157_,
		_w31158_,
		_w31159_
	);
	LUT2 #(
		.INIT('h8)
	) name20648 (
		_w17883_,
		_w19088_,
		_w31160_
	);
	LUT2 #(
		.INIT('h1)
	) name20649 (
		\wishbone_TxPointerMSB_reg[16]/NET0131 ,
		_w31154_,
		_w31161_
	);
	LUT2 #(
		.INIT('h1)
	) name20650 (
		_w17883_,
		_w17900_,
		_w31162_
	);
	LUT2 #(
		.INIT('h4)
	) name20651 (
		_w31161_,
		_w31162_,
		_w31163_
	);
	LUT2 #(
		.INIT('h1)
	) name20652 (
		_w31160_,
		_w31163_,
		_w31164_
	);
	LUT2 #(
		.INIT('h1)
	) name20653 (
		\wishbone_TxPointerMSB_reg[17]/NET0131 ,
		_w17900_,
		_w31165_
	);
	LUT2 #(
		.INIT('h1)
	) name20654 (
		_w17883_,
		_w17901_,
		_w31166_
	);
	LUT2 #(
		.INIT('h4)
	) name20655 (
		_w31165_,
		_w31166_,
		_w31167_
	);
	LUT2 #(
		.INIT('h8)
	) name20656 (
		_w17883_,
		_w20126_,
		_w31168_
	);
	LUT2 #(
		.INIT('h1)
	) name20657 (
		_w31167_,
		_w31168_,
		_w31169_
	);
	LUT2 #(
		.INIT('h1)
	) name20658 (
		\wishbone_TxPointerMSB_reg[18]/NET0131 ,
		_w17901_,
		_w31170_
	);
	LUT2 #(
		.INIT('h1)
	) name20659 (
		_w17883_,
		_w17902_,
		_w31171_
	);
	LUT2 #(
		.INIT('h4)
	) name20660 (
		_w31170_,
		_w31171_,
		_w31172_
	);
	LUT2 #(
		.INIT('h8)
	) name20661 (
		_w17883_,
		_w18564_,
		_w31173_
	);
	LUT2 #(
		.INIT('h1)
	) name20662 (
		_w31172_,
		_w31173_,
		_w31174_
	);
	LUT2 #(
		.INIT('h1)
	) name20663 (
		\wishbone_TxPointerMSB_reg[2]/NET0131 ,
		_w17885_,
		_w31175_
	);
	LUT2 #(
		.INIT('h1)
	) name20664 (
		_w17883_,
		_w17886_,
		_w31176_
	);
	LUT2 #(
		.INIT('h4)
	) name20665 (
		_w31175_,
		_w31176_,
		_w31177_
	);
	LUT2 #(
		.INIT('h8)
	) name20666 (
		_w17883_,
		_w28520_,
		_w31178_
	);
	LUT2 #(
		.INIT('h1)
	) name20667 (
		_w31177_,
		_w31178_,
		_w31179_
	);
	LUT2 #(
		.INIT('h1)
	) name20668 (
		\wishbone_TxPointerMSB_reg[3]/NET0131 ,
		_w17886_,
		_w31180_
	);
	LUT2 #(
		.INIT('h1)
	) name20669 (
		_w17883_,
		_w17887_,
		_w31181_
	);
	LUT2 #(
		.INIT('h4)
	) name20670 (
		_w31180_,
		_w31181_,
		_w31182_
	);
	LUT2 #(
		.INIT('h8)
	) name20671 (
		_w17883_,
		_w24704_,
		_w31183_
	);
	LUT2 #(
		.INIT('h1)
	) name20672 (
		_w31182_,
		_w31183_,
		_w31184_
	);
	LUT2 #(
		.INIT('h1)
	) name20673 (
		\wishbone_TxPointerMSB_reg[8]/NET0131 ,
		_w17891_,
		_w31185_
	);
	LUT2 #(
		.INIT('h1)
	) name20674 (
		_w17883_,
		_w17892_,
		_w31186_
	);
	LUT2 #(
		.INIT('h4)
	) name20675 (
		_w31185_,
		_w31186_,
		_w31187_
	);
	LUT2 #(
		.INIT('h8)
	) name20676 (
		_w17883_,
		_w26900_,
		_w31188_
	);
	LUT2 #(
		.INIT('h1)
	) name20677 (
		_w31187_,
		_w31188_,
		_w31189_
	);
	LUT2 #(
		.INIT('h1)
	) name20678 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		_w31190_
	);
	LUT2 #(
		.INIT('h4)
	) name20679 (
		\miim1_clkgen_Counter_reg[2]/NET0131 ,
		_w31190_,
		_w31191_
	);
	LUT2 #(
		.INIT('h4)
	) name20680 (
		\miim1_clkgen_Counter_reg[3]/NET0131 ,
		_w31191_,
		_w31192_
	);
	LUT2 #(
		.INIT('h4)
	) name20681 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		_w31192_,
		_w31193_
	);
	LUT2 #(
		.INIT('h2)
	) name20682 (
		\miim1_clkgen_Counter_reg[4]/NET0131 ,
		_w31192_,
		_w31194_
	);
	LUT2 #(
		.INIT('h1)
	) name20683 (
		_w31193_,
		_w31194_,
		_w31195_
	);
	LUT2 #(
		.INIT('h1)
	) name20684 (
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w31196_
	);
	LUT2 #(
		.INIT('h1)
	) name20685 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w31197_
	);
	LUT2 #(
		.INIT('h1)
	) name20686 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w31198_
	);
	LUT2 #(
		.INIT('h8)
	) name20687 (
		_w31197_,
		_w31198_,
		_w31199_
	);
	LUT2 #(
		.INIT('h8)
	) name20688 (
		_w31196_,
		_w31199_,
		_w31200_
	);
	LUT2 #(
		.INIT('h1)
	) name20689 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		_w31200_,
		_w31201_
	);
	LUT2 #(
		.INIT('h4)
	) name20690 (
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		_w31201_,
		_w31202_
	);
	LUT2 #(
		.INIT('h4)
	) name20691 (
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w31202_,
		_w31203_
	);
	LUT2 #(
		.INIT('h4)
	) name20692 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		_w31203_,
		_w31204_
	);
	LUT2 #(
		.INIT('h2)
	) name20693 (
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w31204_,
		_w31205_
	);
	LUT2 #(
		.INIT('h4)
	) name20694 (
		\ethreg1_MIIMODER_0_DataOut_reg[5]/NET0131 ,
		_w31204_,
		_w31206_
	);
	LUT2 #(
		.INIT('h4)
	) name20695 (
		\miim1_clkgen_Counter_reg[5]/NET0131 ,
		_w31193_,
		_w31207_
	);
	LUT2 #(
		.INIT('h4)
	) name20696 (
		\miim1_clkgen_Counter_reg[6]/NET0131 ,
		_w31207_,
		_w31208_
	);
	LUT2 #(
		.INIT('h4)
	) name20697 (
		_w31205_,
		_w31208_,
		_w31209_
	);
	LUT2 #(
		.INIT('h4)
	) name20698 (
		_w31206_,
		_w31209_,
		_w31210_
	);
	LUT2 #(
		.INIT('h1)
	) name20699 (
		_w31195_,
		_w31210_,
		_w31211_
	);
	LUT2 #(
		.INIT('h1)
	) name20700 (
		\RxAbort_wb_reg/NET0131 ,
		\wishbone_ShiftEnded_rck_reg/NET0131 ,
		_w31212_
	);
	LUT2 #(
		.INIT('h8)
	) name20701 (
		\rxethmac1_RxValid_reg/NET0131 ,
		\wishbone_RxReady_reg/NET0131 ,
		_w31213_
	);
	LUT2 #(
		.INIT('h8)
	) name20702 (
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w31213_,
		_w31214_
	);
	LUT2 #(
		.INIT('h1)
	) name20703 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w31214_,
		_w31215_
	);
	LUT2 #(
		.INIT('h2)
	) name20704 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w31215_,
		_w31216_
	);
	LUT2 #(
		.INIT('h4)
	) name20705 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w31215_,
		_w31217_
	);
	LUT2 #(
		.INIT('h1)
	) name20706 (
		_w31216_,
		_w31217_,
		_w31218_
	);
	LUT2 #(
		.INIT('h1)
	) name20707 (
		_w15139_,
		_w31218_,
		_w31219_
	);
	LUT2 #(
		.INIT('h4)
	) name20708 (
		_w15140_,
		_w31212_,
		_w31220_
	);
	LUT2 #(
		.INIT('h4)
	) name20709 (
		_w31219_,
		_w31220_,
		_w31221_
	);
	LUT2 #(
		.INIT('h4)
	) name20710 (
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w14570_,
		_w31222_
	);
	LUT2 #(
		.INIT('h4)
	) name20711 (
		_w14571_,
		_w14582_,
		_w31223_
	);
	LUT2 #(
		.INIT('h4)
	) name20712 (
		_w31222_,
		_w31223_,
		_w31224_
	);
	LUT2 #(
		.INIT('h2)
	) name20713 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		_w31225_
	);
	LUT2 #(
		.INIT('h8)
	) name20714 (
		_w11828_,
		_w12645_,
		_w31226_
	);
	LUT2 #(
		.INIT('h8)
	) name20715 (
		_w12651_,
		_w31226_,
		_w31227_
	);
	LUT2 #(
		.INIT('h2)
	) name20716 (
		_w11828_,
		_w31225_,
		_w31228_
	);
	LUT2 #(
		.INIT('h4)
	) name20717 (
		_w31227_,
		_w31228_,
		_w31229_
	);
	LUT2 #(
		.INIT('h8)
	) name20718 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w31229_,
		_w31230_
	);
	LUT2 #(
		.INIT('h8)
	) name20719 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w31230_,
		_w31231_
	);
	LUT2 #(
		.INIT('h8)
	) name20720 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		_w31231_,
		_w31232_
	);
	LUT2 #(
		.INIT('h8)
	) name20721 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w31232_,
		_w31233_
	);
	LUT2 #(
		.INIT('h1)
	) name20722 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w31233_,
		_w31234_
	);
	LUT2 #(
		.INIT('h8)
	) name20723 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[4]/NET0131 ,
		_w31233_,
		_w31235_
	);
	LUT2 #(
		.INIT('h1)
	) name20724 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w31234_,
		_w31236_
	);
	LUT2 #(
		.INIT('h4)
	) name20725 (
		_w31235_,
		_w31236_,
		_w31237_
	);
	LUT2 #(
		.INIT('h2)
	) name20726 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w31238_
	);
	LUT2 #(
		.INIT('h4)
	) name20727 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w31239_
	);
	LUT2 #(
		.INIT('h1)
	) name20728 (
		_w31238_,
		_w31239_,
		_w31240_
	);
	LUT2 #(
		.INIT('h8)
	) name20729 (
		_w15139_,
		_w31240_,
		_w31241_
	);
	LUT2 #(
		.INIT('h1)
	) name20730 (
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		_w31216_,
		_w31242_
	);
	LUT2 #(
		.INIT('h8)
	) name20731 (
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		_w31216_,
		_w31243_
	);
	LUT2 #(
		.INIT('h1)
	) name20732 (
		_w31242_,
		_w31243_,
		_w31244_
	);
	LUT2 #(
		.INIT('h1)
	) name20733 (
		_w15139_,
		_w31244_,
		_w31245_
	);
	LUT2 #(
		.INIT('h2)
	) name20734 (
		_w31212_,
		_w31241_,
		_w31246_
	);
	LUT2 #(
		.INIT('h4)
	) name20735 (
		_w31245_,
		_w31246_,
		_w31247_
	);
	LUT2 #(
		.INIT('h1)
	) name20736 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[0]/NET0131 ,
		_w31229_,
		_w31248_
	);
	LUT2 #(
		.INIT('h1)
	) name20737 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w31230_,
		_w31249_
	);
	LUT2 #(
		.INIT('h4)
	) name20738 (
		_w31248_,
		_w31249_,
		_w31250_
	);
	LUT2 #(
		.INIT('h1)
	) name20739 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[2]/NET0131 ,
		_w31231_,
		_w31251_
	);
	LUT2 #(
		.INIT('h1)
	) name20740 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w31232_,
		_w31252_
	);
	LUT2 #(
		.INIT('h4)
	) name20741 (
		_w31251_,
		_w31252_,
		_w31253_
	);
	LUT2 #(
		.INIT('h1)
	) name20742 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[3]/NET0131 ,
		_w31232_,
		_w31254_
	);
	LUT2 #(
		.INIT('h1)
	) name20743 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w31233_,
		_w31255_
	);
	LUT2 #(
		.INIT('h4)
	) name20744 (
		_w31254_,
		_w31255_,
		_w31256_
	);
	LUT2 #(
		.INIT('h1)
	) name20745 (
		\txethmac1_txcounters1_ByteCnt_reg[10]/NET0131 ,
		_w14576_,
		_w31257_
	);
	LUT2 #(
		.INIT('h4)
	) name20746 (
		_w14577_,
		_w14582_,
		_w31258_
	);
	LUT2 #(
		.INIT('h4)
	) name20747 (
		_w31257_,
		_w31258_,
		_w31259_
	);
	LUT2 #(
		.INIT('h1)
	) name20748 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w14578_,
		_w31260_
	);
	LUT2 #(
		.INIT('h8)
	) name20749 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w14578_,
		_w31261_
	);
	LUT2 #(
		.INIT('h2)
	) name20750 (
		_w14582_,
		_w31260_,
		_w31262_
	);
	LUT2 #(
		.INIT('h4)
	) name20751 (
		_w31261_,
		_w31262_,
		_w31263_
	);
	LUT2 #(
		.INIT('h8)
	) name20752 (
		\txethmac1_txcounters1_ByteCnt_reg[12]/NET0131 ,
		_w14566_,
		_w31264_
	);
	LUT2 #(
		.INIT('h4)
	) name20753 (
		_w14570_,
		_w31264_,
		_w31265_
	);
	LUT2 #(
		.INIT('h1)
	) name20754 (
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w31265_,
		_w31266_
	);
	LUT2 #(
		.INIT('h8)
	) name20755 (
		\txethmac1_txcounters1_ByteCnt_reg[13]/NET0131 ,
		_w31265_,
		_w31267_
	);
	LUT2 #(
		.INIT('h2)
	) name20756 (
		_w14582_,
		_w31266_,
		_w31268_
	);
	LUT2 #(
		.INIT('h4)
	) name20757 (
		_w31267_,
		_w31268_,
		_w31269_
	);
	LUT2 #(
		.INIT('h1)
	) name20758 (
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w31267_,
		_w31270_
	);
	LUT2 #(
		.INIT('h8)
	) name20759 (
		\txethmac1_txcounters1_ByteCnt_reg[14]/NET0131 ,
		_w31267_,
		_w31271_
	);
	LUT2 #(
		.INIT('h2)
	) name20760 (
		_w14582_,
		_w31270_,
		_w31272_
	);
	LUT2 #(
		.INIT('h4)
	) name20761 (
		_w31271_,
		_w31272_,
		_w31273_
	);
	LUT2 #(
		.INIT('h1)
	) name20762 (
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w14571_,
		_w31274_
	);
	LUT2 #(
		.INIT('h4)
	) name20763 (
		_w14572_,
		_w14582_,
		_w31275_
	);
	LUT2 #(
		.INIT('h4)
	) name20764 (
		_w31274_,
		_w31275_,
		_w31276_
	);
	LUT2 #(
		.INIT('h1)
	) name20765 (
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w14572_,
		_w31277_
	);
	LUT2 #(
		.INIT('h4)
	) name20766 (
		_w14573_,
		_w14582_,
		_w31278_
	);
	LUT2 #(
		.INIT('h4)
	) name20767 (
		_w31277_,
		_w31278_,
		_w31279_
	);
	LUT2 #(
		.INIT('h1)
	) name20768 (
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w14573_,
		_w31280_
	);
	LUT2 #(
		.INIT('h4)
	) name20769 (
		_w14574_,
		_w14582_,
		_w31281_
	);
	LUT2 #(
		.INIT('h4)
	) name20770 (
		_w31280_,
		_w31281_,
		_w31282_
	);
	LUT2 #(
		.INIT('h8)
	) name20771 (
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w14574_,
		_w31283_
	);
	LUT2 #(
		.INIT('h1)
	) name20772 (
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w14574_,
		_w31284_
	);
	LUT2 #(
		.INIT('h2)
	) name20773 (
		_w14582_,
		_w31283_,
		_w31285_
	);
	LUT2 #(
		.INIT('h4)
	) name20774 (
		_w31284_,
		_w31285_,
		_w31286_
	);
	LUT2 #(
		.INIT('h8)
	) name20775 (
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w31283_,
		_w31287_
	);
	LUT2 #(
		.INIT('h1)
	) name20776 (
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w31283_,
		_w31288_
	);
	LUT2 #(
		.INIT('h2)
	) name20777 (
		_w14582_,
		_w31287_,
		_w31289_
	);
	LUT2 #(
		.INIT('h4)
	) name20778 (
		_w31288_,
		_w31289_,
		_w31290_
	);
	LUT2 #(
		.INIT('h8)
	) name20779 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w31287_,
		_w31291_
	);
	LUT2 #(
		.INIT('h1)
	) name20780 (
		\txethmac1_txcounters1_ByteCnt_reg[6]/NET0131 ,
		_w31287_,
		_w31292_
	);
	LUT2 #(
		.INIT('h2)
	) name20781 (
		_w14582_,
		_w31291_,
		_w31293_
	);
	LUT2 #(
		.INIT('h4)
	) name20782 (
		_w31292_,
		_w31293_,
		_w31294_
	);
	LUT2 #(
		.INIT('h8)
	) name20783 (
		_w14554_,
		_w31287_,
		_w31295_
	);
	LUT2 #(
		.INIT('h1)
	) name20784 (
		\txethmac1_txcounters1_ByteCnt_reg[7]/NET0131 ,
		_w31291_,
		_w31296_
	);
	LUT2 #(
		.INIT('h2)
	) name20785 (
		_w14582_,
		_w31295_,
		_w31297_
	);
	LUT2 #(
		.INIT('h4)
	) name20786 (
		_w31296_,
		_w31297_,
		_w31298_
	);
	LUT2 #(
		.INIT('h1)
	) name20787 (
		\txethmac1_txcounters1_ByteCnt_reg[8]/NET0131 ,
		_w31295_,
		_w31299_
	);
	LUT2 #(
		.INIT('h4)
	) name20788 (
		_w14575_,
		_w14582_,
		_w31300_
	);
	LUT2 #(
		.INIT('h4)
	) name20789 (
		_w31299_,
		_w31300_,
		_w31301_
	);
	LUT2 #(
		.INIT('h2)
	) name20790 (
		_w14564_,
		_w14570_,
		_w31302_
	);
	LUT2 #(
		.INIT('h2)
	) name20791 (
		_w14563_,
		_w14570_,
		_w31303_
	);
	LUT2 #(
		.INIT('h1)
	) name20792 (
		\txethmac1_txcounters1_ByteCnt_reg[9]/NET0131 ,
		_w31303_,
		_w31304_
	);
	LUT2 #(
		.INIT('h2)
	) name20793 (
		_w14582_,
		_w31302_,
		_w31305_
	);
	LUT2 #(
		.INIT('h4)
	) name20794 (
		_w31304_,
		_w31305_,
		_w31306_
	);
	LUT2 #(
		.INIT('h2)
	) name20795 (
		\txethmac1_txcrc_Crc_reg[3]/NET0131 ,
		_w12458_,
		_w31307_
	);
	LUT2 #(
		.INIT('h4)
	) name20796 (
		\txethmac1_txcrc_Crc_reg[3]/NET0131 ,
		_w12458_,
		_w31308_
	);
	LUT2 #(
		.INIT('h2)
	) name20797 (
		_w11181_,
		_w31307_,
		_w31309_
	);
	LUT2 #(
		.INIT('h4)
	) name20798 (
		_w31308_,
		_w31309_,
		_w31310_
	);
	LUT2 #(
		.INIT('h2)
	) name20799 (
		\txethmac1_txcrc_Crc_reg[2]/NET0131 ,
		_w11422_,
		_w31311_
	);
	LUT2 #(
		.INIT('h4)
	) name20800 (
		\txethmac1_txcrc_Crc_reg[2]/NET0131 ,
		_w11422_,
		_w31312_
	);
	LUT2 #(
		.INIT('h2)
	) name20801 (
		_w11181_,
		_w31311_,
		_w31313_
	);
	LUT2 #(
		.INIT('h4)
	) name20802 (
		_w31312_,
		_w31313_,
		_w31314_
	);
	LUT2 #(
		.INIT('h4)
	) name20803 (
		_w12557_,
		_w12566_,
		_w31315_
	);
	LUT2 #(
		.INIT('h2)
	) name20804 (
		_w12543_,
		_w12563_,
		_w31316_
	);
	LUT2 #(
		.INIT('h2)
	) name20805 (
		_w12554_,
		_w12557_,
		_w31317_
	);
	LUT2 #(
		.INIT('h4)
	) name20806 (
		_w12543_,
		_w31317_,
		_w31318_
	);
	LUT2 #(
		.INIT('h1)
	) name20807 (
		_w12564_,
		_w12568_,
		_w31319_
	);
	LUT2 #(
		.INIT('h4)
	) name20808 (
		_w31318_,
		_w31319_,
		_w31320_
	);
	LUT2 #(
		.INIT('h1)
	) name20809 (
		_w31316_,
		_w31320_,
		_w31321_
	);
	LUT2 #(
		.INIT('h4)
	) name20810 (
		_w31315_,
		_w31321_,
		_w31322_
	);
	LUT2 #(
		.INIT('h8)
	) name20811 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12611_,
		_w31323_
	);
	LUT2 #(
		.INIT('h4)
	) name20812 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12558_,
		_w31324_
	);
	LUT2 #(
		.INIT('h8)
	) name20813 (
		_w12542_,
		_w12568_,
		_w31325_
	);
	LUT2 #(
		.INIT('h4)
	) name20814 (
		_w31324_,
		_w31325_,
		_w31326_
	);
	LUT2 #(
		.INIT('h4)
	) name20815 (
		_w31317_,
		_w31326_,
		_w31327_
	);
	LUT2 #(
		.INIT('h4)
	) name20816 (
		_w31323_,
		_w31327_,
		_w31328_
	);
	LUT2 #(
		.INIT('h1)
	) name20817 (
		_w31318_,
		_w31328_,
		_w31329_
	);
	LUT2 #(
		.INIT('h8)
	) name20818 (
		_w31322_,
		_w31329_,
		_w31330_
	);
	LUT2 #(
		.INIT('h2)
	) name20819 (
		\m_wb_sel_o[0]_pad ,
		_w31330_,
		_w31331_
	);
	LUT2 #(
		.INIT('h2)
	) name20820 (
		_w12636_,
		_w31331_,
		_w31332_
	);
	LUT2 #(
		.INIT('h2)
	) name20821 (
		\macstatus1_InvalidSymbol_reg/NET0131 ,
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w31333_
	);
	LUT2 #(
		.INIT('h8)
	) name20822 (
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		mtxerr_pad_o_pad,
		_w31334_
	);
	LUT2 #(
		.INIT('h2)
	) name20823 (
		\RxEnSync_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		_w31335_
	);
	LUT2 #(
		.INIT('h8)
	) name20824 (
		mrxerr_pad_i_pad,
		_w31335_,
		_w31336_
	);
	LUT2 #(
		.INIT('h1)
	) name20825 (
		_w31334_,
		_w31336_,
		_w31337_
	);
	LUT2 #(
		.INIT('h1)
	) name20826 (
		_w10586_,
		_w31337_,
		_w31338_
	);
	LUT2 #(
		.INIT('h1)
	) name20827 (
		_w10666_,
		_w11229_,
		_w31339_
	);
	LUT2 #(
		.INIT('h8)
	) name20828 (
		_w11786_,
		_w31339_,
		_w31340_
	);
	LUT2 #(
		.INIT('h8)
	) name20829 (
		_w31338_,
		_w31340_,
		_w31341_
	);
	LUT2 #(
		.INIT('h1)
	) name20830 (
		_w31333_,
		_w31341_,
		_w31342_
	);
	LUT2 #(
		.INIT('h8)
	) name20831 (
		\wishbone_ShiftEndedSync_c1_reg/NET0131 ,
		\wishbone_ShiftEndedSync_c2_reg/NET0131 ,
		_w31343_
	);
	LUT2 #(
		.INIT('h2)
	) name20832 (
		\wishbone_ShiftEnded_rck_reg/NET0131 ,
		_w31343_,
		_w31344_
	);
	LUT2 #(
		.INIT('h8)
	) name20833 (
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w31345_
	);
	LUT2 #(
		.INIT('h8)
	) name20834 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		\rxethmac1_RxValid_reg/NET0131 ,
		_w31346_
	);
	LUT2 #(
		.INIT('h8)
	) name20835 (
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w31345_,
		_w31347_
	);
	LUT2 #(
		.INIT('h8)
	) name20836 (
		_w31346_,
		_w31347_,
		_w31348_
	);
	LUT2 #(
		.INIT('h1)
	) name20837 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w31348_,
		_w31349_
	);
	LUT2 #(
		.INIT('h1)
	) name20838 (
		_w15147_,
		_w31349_,
		_w31350_
	);
	LUT2 #(
		.INIT('h1)
	) name20839 (
		_w31344_,
		_w31350_,
		_w31351_
	);
	LUT2 #(
		.INIT('h1)
	) name20840 (
		\RxAbort_wb_reg/NET0131 ,
		_w31351_,
		_w31352_
	);
	LUT2 #(
		.INIT('h1)
	) name20841 (
		\maccontrol1_receivecontrol1_ByteCnt_reg[1]/NET0131 ,
		_w31230_,
		_w31353_
	);
	LUT2 #(
		.INIT('h1)
	) name20842 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w31231_,
		_w31354_
	);
	LUT2 #(
		.INIT('h4)
	) name20843 (
		_w31353_,
		_w31354_,
		_w31355_
	);
	LUT2 #(
		.INIT('h2)
	) name20844 (
		m_wb_stb_o_pad,
		_w31322_,
		_w31356_
	);
	LUT2 #(
		.INIT('h2)
	) name20845 (
		_w12636_,
		_w31356_,
		_w31357_
	);
	LUT2 #(
		.INIT('h1)
	) name20846 (
		_w31315_,
		_w31328_,
		_w31358_
	);
	LUT2 #(
		.INIT('h4)
	) name20847 (
		_w12561_,
		_w31358_,
		_w31359_
	);
	LUT2 #(
		.INIT('h8)
	) name20848 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		_w31360_
	);
	LUT2 #(
		.INIT('h4)
	) name20849 (
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w31360_,
		_w31361_
	);
	LUT2 #(
		.INIT('h2)
	) name20850 (
		_w12561_,
		_w31361_,
		_w31362_
	);
	LUT2 #(
		.INIT('h1)
	) name20851 (
		_w31359_,
		_w31362_,
		_w31363_
	);
	LUT2 #(
		.INIT('h2)
	) name20852 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w31363_,
		_w31364_
	);
	LUT2 #(
		.INIT('h8)
	) name20853 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w31365_
	);
	LUT2 #(
		.INIT('h2)
	) name20854 (
		\wishbone_TxLength_reg[2]/NET0131 ,
		_w16763_,
		_w31366_
	);
	LUT2 #(
		.INIT('h1)
	) name20855 (
		\wishbone_TxLength_reg[3]/NET0131 ,
		_w31366_,
		_w31367_
	);
	LUT2 #(
		.INIT('h2)
	) name20856 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w31367_,
		_w31368_
	);
	LUT2 #(
		.INIT('h8)
	) name20857 (
		_w13479_,
		_w13482_,
		_w31369_
	);
	LUT2 #(
		.INIT('h8)
	) name20858 (
		_w13498_,
		_w31369_,
		_w31370_
	);
	LUT2 #(
		.INIT('h4)
	) name20859 (
		_w31368_,
		_w31370_,
		_w31371_
	);
	LUT2 #(
		.INIT('h1)
	) name20860 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w31365_,
		_w31372_
	);
	LUT2 #(
		.INIT('h4)
	) name20861 (
		_w31371_,
		_w31372_,
		_w31373_
	);
	LUT2 #(
		.INIT('h4)
	) name20862 (
		_w31358_,
		_w31373_,
		_w31374_
	);
	LUT2 #(
		.INIT('h1)
	) name20863 (
		_w31364_,
		_w31374_,
		_w31375_
	);
	LUT2 #(
		.INIT('h2)
	) name20864 (
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w31322_,
		_w31376_
	);
	LUT2 #(
		.INIT('h2)
	) name20865 (
		_w12573_,
		_w31376_,
		_w31377_
	);
	LUT2 #(
		.INIT('h8)
	) name20866 (
		_w12628_,
		_w12629_,
		_w31378_
	);
	LUT2 #(
		.INIT('h8)
	) name20867 (
		_w12562_,
		_w12570_,
		_w31379_
	);
	LUT2 #(
		.INIT('h2)
	) name20868 (
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w31318_,
		_w31380_
	);
	LUT2 #(
		.INIT('h4)
	) name20869 (
		_w31378_,
		_w31380_,
		_w31381_
	);
	LUT2 #(
		.INIT('h1)
	) name20870 (
		_w12621_,
		_w31379_,
		_w31382_
	);
	LUT2 #(
		.INIT('h8)
	) name20871 (
		_w31381_,
		_w31382_,
		_w31383_
	);
	LUT2 #(
		.INIT('h4)
	) name20872 (
		_w12561_,
		_w31383_,
		_w31384_
	);
	LUT2 #(
		.INIT('h1)
	) name20873 (
		_w31328_,
		_w31384_,
		_w31385_
	);
	LUT2 #(
		.INIT('h1)
	) name20874 (
		\txethmac1_StatusLatch_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w31386_
	);
	LUT2 #(
		.INIT('h4)
	) name20875 (
		_w11266_,
		_w31386_,
		_w31387_
	);
	LUT2 #(
		.INIT('h1)
	) name20876 (
		_w11099_,
		_w31387_,
		_w31388_
	);
	LUT2 #(
		.INIT('h8)
	) name20877 (
		_w10582_,
		_w12122_,
		_w31389_
	);
	LUT2 #(
		.INIT('h2)
	) name20878 (
		_w31338_,
		_w31389_,
		_w31390_
	);
	LUT2 #(
		.INIT('h4)
	) name20879 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifo_reg/NET0131 ,
		_w31391_
	);
	LUT2 #(
		.INIT('h2)
	) name20880 (
		_w15147_,
		_w31391_,
		_w31392_
	);
	LUT2 #(
		.INIT('h1)
	) name20881 (
		\RxAbort_wb_reg/NET0131 ,
		_w31392_,
		_w31393_
	);
	LUT2 #(
		.INIT('h2)
	) name20882 (
		\ethreg1_MIIMODER_0_DataOut_reg[4]/NET0131 ,
		_w31203_,
		_w31394_
	);
	LUT2 #(
		.INIT('h4)
	) name20883 (
		_w31204_,
		_w31208_,
		_w31395_
	);
	LUT2 #(
		.INIT('h4)
	) name20884 (
		_w31394_,
		_w31395_,
		_w31396_
	);
	LUT2 #(
		.INIT('h2)
	) name20885 (
		\miim1_clkgen_Counter_reg[3]/NET0131 ,
		_w31191_,
		_w31397_
	);
	LUT2 #(
		.INIT('h1)
	) name20886 (
		_w31192_,
		_w31397_,
		_w31398_
	);
	LUT2 #(
		.INIT('h4)
	) name20887 (
		_w31208_,
		_w31398_,
		_w31399_
	);
	LUT2 #(
		.INIT('h1)
	) name20888 (
		_w31396_,
		_w31399_,
		_w31400_
	);
	LUT2 #(
		.INIT('h8)
	) name20889 (
		mdc_pad_o_pad,
		_w31208_,
		_w31401_
	);
	LUT2 #(
		.INIT('h2)
	) name20890 (
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w31401_,
		_w31402_
	);
	LUT2 #(
		.INIT('h1)
	) name20891 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		_w31403_
	);
	LUT2 #(
		.INIT('h1)
	) name20892 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w31404_
	);
	LUT2 #(
		.INIT('h2)
	) name20893 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w31405_
	);
	LUT2 #(
		.INIT('h1)
	) name20894 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w31406_
	);
	LUT2 #(
		.INIT('h8)
	) name20895 (
		_w31405_,
		_w31406_,
		_w31407_
	);
	LUT2 #(
		.INIT('h8)
	) name20896 (
		_w31403_,
		_w31404_,
		_w31408_
	);
	LUT2 #(
		.INIT('h8)
	) name20897 (
		_w31407_,
		_w31408_,
		_w31409_
	);
	LUT2 #(
		.INIT('h8)
	) name20898 (
		\miim1_InProgress_reg/NET0131 ,
		_w31409_,
		_w31410_
	);
	LUT2 #(
		.INIT('h4)
	) name20899 (
		\miim1_BitCounter_reg[6]/NET0131 ,
		\miim1_InProgress_reg/NET0131 ,
		_w31411_
	);
	LUT2 #(
		.INIT('h4)
	) name20900 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w31411_,
		_w31412_
	);
	LUT2 #(
		.INIT('h4)
	) name20901 (
		\miim1_BitCounter_reg[2]/NET0131 ,
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w31413_
	);
	LUT2 #(
		.INIT('h8)
	) name20902 (
		_w31403_,
		_w31413_,
		_w31414_
	);
	LUT2 #(
		.INIT('h1)
	) name20903 (
		\ethreg1_MIIMODER_1_DataOut_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w31415_
	);
	LUT2 #(
		.INIT('h8)
	) name20904 (
		_w31412_,
		_w31415_,
		_w31416_
	);
	LUT2 #(
		.INIT('h8)
	) name20905 (
		_w31414_,
		_w31416_,
		_w31417_
	);
	LUT2 #(
		.INIT('h1)
	) name20906 (
		_w31410_,
		_w31417_,
		_w31418_
	);
	LUT2 #(
		.INIT('h2)
	) name20907 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[2]/NET0131 ,
		_w31418_,
		_w31419_
	);
	LUT2 #(
		.INIT('h8)
	) name20908 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w31411_,
		_w31420_
	);
	LUT2 #(
		.INIT('h8)
	) name20909 (
		\miim1_WriteOp_reg/NET0131 ,
		_w31414_,
		_w31421_
	);
	LUT2 #(
		.INIT('h8)
	) name20910 (
		_w31420_,
		_w31421_,
		_w31422_
	);
	LUT2 #(
		.INIT('h8)
	) name20911 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w31412_,
		_w31423_
	);
	LUT2 #(
		.INIT('h8)
	) name20912 (
		_w31414_,
		_w31423_,
		_w31424_
	);
	LUT2 #(
		.INIT('h1)
	) name20913 (
		_w31422_,
		_w31424_,
		_w31425_
	);
	LUT2 #(
		.INIT('h8)
	) name20914 (
		_w31418_,
		_w31425_,
		_w31426_
	);
	LUT2 #(
		.INIT('h8)
	) name20915 (
		\miim1_shftrg_ShiftReg_reg[0]/NET0131 ,
		_w31426_,
		_w31427_
	);
	LUT2 #(
		.INIT('h4)
	) name20916 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w31422_,
		_w31428_
	);
	LUT2 #(
		.INIT('h8)
	) name20917 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[1]/NET0131 ,
		_w31428_,
		_w31429_
	);
	LUT2 #(
		.INIT('h8)
	) name20918 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w31422_,
		_w31430_
	);
	LUT2 #(
		.INIT('h8)
	) name20919 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[1]/NET0131 ,
		_w31430_,
		_w31431_
	);
	LUT2 #(
		.INIT('h1)
	) name20920 (
		_w31419_,
		_w31424_,
		_w31432_
	);
	LUT2 #(
		.INIT('h1)
	) name20921 (
		_w31429_,
		_w31431_,
		_w31433_
	);
	LUT2 #(
		.INIT('h8)
	) name20922 (
		_w31432_,
		_w31433_,
		_w31434_
	);
	LUT2 #(
		.INIT('h4)
	) name20923 (
		_w31427_,
		_w31434_,
		_w31435_
	);
	LUT2 #(
		.INIT('h2)
	) name20924 (
		_w31401_,
		_w31435_,
		_w31436_
	);
	LUT2 #(
		.INIT('h1)
	) name20925 (
		_w31402_,
		_w31436_,
		_w31437_
	);
	LUT2 #(
		.INIT('h2)
	) name20926 (
		\miim1_shftrg_ShiftReg_reg[2]/NET0131 ,
		_w31401_,
		_w31438_
	);
	LUT2 #(
		.INIT('h8)
	) name20927 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[2]/NET0131 ,
		_w31430_,
		_w31439_
	);
	LUT2 #(
		.INIT('h8)
	) name20928 (
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w31426_,
		_w31440_
	);
	LUT2 #(
		.INIT('h8)
	) name20929 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 ,
		_w31428_,
		_w31441_
	);
	LUT2 #(
		.INIT('h2)
	) name20930 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[3]/NET0131 ,
		_w31418_,
		_w31442_
	);
	LUT2 #(
		.INIT('h8)
	) name20931 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		_w31424_,
		_w31443_
	);
	LUT2 #(
		.INIT('h1)
	) name20932 (
		_w31439_,
		_w31443_,
		_w31444_
	);
	LUT2 #(
		.INIT('h1)
	) name20933 (
		_w31441_,
		_w31442_,
		_w31445_
	);
	LUT2 #(
		.INIT('h8)
	) name20934 (
		_w31444_,
		_w31445_,
		_w31446_
	);
	LUT2 #(
		.INIT('h4)
	) name20935 (
		_w31440_,
		_w31446_,
		_w31447_
	);
	LUT2 #(
		.INIT('h2)
	) name20936 (
		_w31401_,
		_w31447_,
		_w31448_
	);
	LUT2 #(
		.INIT('h1)
	) name20937 (
		_w31438_,
		_w31448_,
		_w31449_
	);
	LUT2 #(
		.INIT('h2)
	) name20938 (
		\miim1_shftrg_ShiftReg_reg[3]/NET0131 ,
		_w31401_,
		_w31450_
	);
	LUT2 #(
		.INIT('h8)
	) name20939 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[3]/NET0131 ,
		_w31430_,
		_w31451_
	);
	LUT2 #(
		.INIT('h8)
	) name20940 (
		\miim1_shftrg_ShiftReg_reg[2]/NET0131 ,
		_w31426_,
		_w31452_
	);
	LUT2 #(
		.INIT('h8)
	) name20941 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[3]/NET0131 ,
		_w31428_,
		_w31453_
	);
	LUT2 #(
		.INIT('h2)
	) name20942 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[4]/NET0131 ,
		_w31418_,
		_w31454_
	);
	LUT2 #(
		.INIT('h8)
	) name20943 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w31424_,
		_w31455_
	);
	LUT2 #(
		.INIT('h1)
	) name20944 (
		_w31451_,
		_w31455_,
		_w31456_
	);
	LUT2 #(
		.INIT('h1)
	) name20945 (
		_w31453_,
		_w31454_,
		_w31457_
	);
	LUT2 #(
		.INIT('h8)
	) name20946 (
		_w31456_,
		_w31457_,
		_w31458_
	);
	LUT2 #(
		.INIT('h4)
	) name20947 (
		_w31452_,
		_w31458_,
		_w31459_
	);
	LUT2 #(
		.INIT('h2)
	) name20948 (
		_w31401_,
		_w31459_,
		_w31460_
	);
	LUT2 #(
		.INIT('h1)
	) name20949 (
		_w31450_,
		_w31460_,
		_w31461_
	);
	LUT2 #(
		.INIT('h2)
	) name20950 (
		\miim1_shftrg_ShiftReg_reg[4]/NET0131 ,
		_w31401_,
		_w31462_
	);
	LUT2 #(
		.INIT('h8)
	) name20951 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[4]/NET0131 ,
		_w31430_,
		_w31463_
	);
	LUT2 #(
		.INIT('h8)
	) name20952 (
		\miim1_shftrg_ShiftReg_reg[3]/NET0131 ,
		_w31426_,
		_w31464_
	);
	LUT2 #(
		.INIT('h8)
	) name20953 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[4]/NET0131 ,
		_w31428_,
		_w31465_
	);
	LUT2 #(
		.INIT('h2)
	) name20954 (
		\miim1_WriteOp_reg/NET0131 ,
		_w31418_,
		_w31466_
	);
	LUT2 #(
		.INIT('h8)
	) name20955 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		_w31424_,
		_w31467_
	);
	LUT2 #(
		.INIT('h1)
	) name20956 (
		_w31463_,
		_w31467_,
		_w31468_
	);
	LUT2 #(
		.INIT('h1)
	) name20957 (
		_w31465_,
		_w31466_,
		_w31469_
	);
	LUT2 #(
		.INIT('h8)
	) name20958 (
		_w31468_,
		_w31469_,
		_w31470_
	);
	LUT2 #(
		.INIT('h4)
	) name20959 (
		_w31464_,
		_w31470_,
		_w31471_
	);
	LUT2 #(
		.INIT('h2)
	) name20960 (
		_w31401_,
		_w31471_,
		_w31472_
	);
	LUT2 #(
		.INIT('h1)
	) name20961 (
		_w31462_,
		_w31472_,
		_w31473_
	);
	LUT2 #(
		.INIT('h2)
	) name20962 (
		\miim1_shftrg_ShiftReg_reg[5]/NET0131 ,
		_w31401_,
		_w31474_
	);
	LUT2 #(
		.INIT('h8)
	) name20963 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[5]/NET0131 ,
		_w31430_,
		_w31475_
	);
	LUT2 #(
		.INIT('h8)
	) name20964 (
		\miim1_shftrg_ShiftReg_reg[4]/NET0131 ,
		_w31426_,
		_w31476_
	);
	LUT2 #(
		.INIT('h8)
	) name20965 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[5]/NET0131 ,
		_w31428_,
		_w31477_
	);
	LUT2 #(
		.INIT('h1)
	) name20966 (
		\miim1_WriteOp_reg/NET0131 ,
		_w31418_,
		_w31478_
	);
	LUT2 #(
		.INIT('h8)
	) name20967 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		_w31424_,
		_w31479_
	);
	LUT2 #(
		.INIT('h1)
	) name20968 (
		_w31475_,
		_w31479_,
		_w31480_
	);
	LUT2 #(
		.INIT('h1)
	) name20969 (
		_w31477_,
		_w31478_,
		_w31481_
	);
	LUT2 #(
		.INIT('h8)
	) name20970 (
		_w31480_,
		_w31481_,
		_w31482_
	);
	LUT2 #(
		.INIT('h4)
	) name20971 (
		_w31476_,
		_w31482_,
		_w31483_
	);
	LUT2 #(
		.INIT('h2)
	) name20972 (
		_w31401_,
		_w31483_,
		_w31484_
	);
	LUT2 #(
		.INIT('h1)
	) name20973 (
		_w31474_,
		_w31484_,
		_w31485_
	);
	LUT2 #(
		.INIT('h2)
	) name20974 (
		\miim1_shftrg_ShiftReg_reg[6]/NET0131 ,
		_w31401_,
		_w31486_
	);
	LUT2 #(
		.INIT('h8)
	) name20975 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w31424_,
		_w31487_
	);
	LUT2 #(
		.INIT('h8)
	) name20976 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[6]/NET0131 ,
		_w31428_,
		_w31488_
	);
	LUT2 #(
		.INIT('h8)
	) name20977 (
		\miim1_shftrg_ShiftReg_reg[5]/NET0131 ,
		_w31425_,
		_w31489_
	);
	LUT2 #(
		.INIT('h8)
	) name20978 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[6]/NET0131 ,
		_w31430_,
		_w31490_
	);
	LUT2 #(
		.INIT('h2)
	) name20979 (
		_w31418_,
		_w31487_,
		_w31491_
	);
	LUT2 #(
		.INIT('h4)
	) name20980 (
		_w31488_,
		_w31491_,
		_w31492_
	);
	LUT2 #(
		.INIT('h1)
	) name20981 (
		_w31489_,
		_w31490_,
		_w31493_
	);
	LUT2 #(
		.INIT('h8)
	) name20982 (
		_w31492_,
		_w31493_,
		_w31494_
	);
	LUT2 #(
		.INIT('h2)
	) name20983 (
		_w31401_,
		_w31494_,
		_w31495_
	);
	LUT2 #(
		.INIT('h1)
	) name20984 (
		_w31486_,
		_w31495_,
		_w31496_
	);
	LUT2 #(
		.INIT('h4)
	) name20985 (
		\txethmac1_TxAbort_reg/NET0131 ,
		_w11385_,
		_w31497_
	);
	LUT2 #(
		.INIT('h4)
	) name20986 (
		_w11266_,
		_w11388_,
		_w31498_
	);
	LUT2 #(
		.INIT('h1)
	) name20987 (
		_w31497_,
		_w31498_,
		_w31499_
	);
	LUT2 #(
		.INIT('h8)
	) name20988 (
		\rxethmac1_CrcHashGood_reg/P0001 ,
		\rxethmac1_Multicast_reg/NET0131 ,
		_w31500_
	);
	LUT2 #(
		.INIT('h1)
	) name20989 (
		\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 ,
		_w31500_,
		_w31501_
	);
	LUT2 #(
		.INIT('h8)
	) name20990 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		_w31502_
	);
	LUT2 #(
		.INIT('h1)
	) name20991 (
		\ethreg1_RXHASH0_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31503_
	);
	LUT2 #(
		.INIT('h4)
	) name20992 (
		\ethreg1_RXHASH1_3_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31504_
	);
	LUT2 #(
		.INIT('h2)
	) name20993 (
		_w31502_,
		_w31503_,
		_w31505_
	);
	LUT2 #(
		.INIT('h4)
	) name20994 (
		_w31504_,
		_w31505_,
		_w31506_
	);
	LUT2 #(
		.INIT('h4)
	) name20995 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		_w31507_
	);
	LUT2 #(
		.INIT('h1)
	) name20996 (
		\ethreg1_RXHASH0_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31508_
	);
	LUT2 #(
		.INIT('h4)
	) name20997 (
		\ethreg1_RXHASH1_2_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31509_
	);
	LUT2 #(
		.INIT('h2)
	) name20998 (
		_w31507_,
		_w31508_,
		_w31510_
	);
	LUT2 #(
		.INIT('h4)
	) name20999 (
		_w31509_,
		_w31510_,
		_w31511_
	);
	LUT2 #(
		.INIT('h1)
	) name21000 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		_w31512_
	);
	LUT2 #(
		.INIT('h1)
	) name21001 (
		\ethreg1_RXHASH0_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31513_
	);
	LUT2 #(
		.INIT('h4)
	) name21002 (
		\ethreg1_RXHASH1_0_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31514_
	);
	LUT2 #(
		.INIT('h2)
	) name21003 (
		_w31512_,
		_w31513_,
		_w31515_
	);
	LUT2 #(
		.INIT('h4)
	) name21004 (
		_w31514_,
		_w31515_,
		_w31516_
	);
	LUT2 #(
		.INIT('h2)
	) name21005 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		_w31517_
	);
	LUT2 #(
		.INIT('h1)
	) name21006 (
		\ethreg1_RXHASH0_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31518_
	);
	LUT2 #(
		.INIT('h4)
	) name21007 (
		\ethreg1_RXHASH1_1_DataOut_reg[5]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31519_
	);
	LUT2 #(
		.INIT('h2)
	) name21008 (
		_w31517_,
		_w31518_,
		_w31520_
	);
	LUT2 #(
		.INIT('h4)
	) name21009 (
		_w31519_,
		_w31520_,
		_w31521_
	);
	LUT2 #(
		.INIT('h2)
	) name21010 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31506_,
		_w31522_
	);
	LUT2 #(
		.INIT('h1)
	) name21011 (
		_w31511_,
		_w31516_,
		_w31523_
	);
	LUT2 #(
		.INIT('h4)
	) name21012 (
		_w31521_,
		_w31523_,
		_w31524_
	);
	LUT2 #(
		.INIT('h8)
	) name21013 (
		_w31522_,
		_w31524_,
		_w31525_
	);
	LUT2 #(
		.INIT('h1)
	) name21014 (
		\ethreg1_RXHASH0_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31526_
	);
	LUT2 #(
		.INIT('h4)
	) name21015 (
		\ethreg1_RXHASH1_0_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31527_
	);
	LUT2 #(
		.INIT('h2)
	) name21016 (
		_w31512_,
		_w31526_,
		_w31528_
	);
	LUT2 #(
		.INIT('h4)
	) name21017 (
		_w31527_,
		_w31528_,
		_w31529_
	);
	LUT2 #(
		.INIT('h1)
	) name21018 (
		\ethreg1_RXHASH0_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31530_
	);
	LUT2 #(
		.INIT('h4)
	) name21019 (
		\ethreg1_RXHASH1_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31531_
	);
	LUT2 #(
		.INIT('h2)
	) name21020 (
		_w31517_,
		_w31530_,
		_w31532_
	);
	LUT2 #(
		.INIT('h4)
	) name21021 (
		_w31531_,
		_w31532_,
		_w31533_
	);
	LUT2 #(
		.INIT('h1)
	) name21022 (
		\ethreg1_RXHASH0_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31534_
	);
	LUT2 #(
		.INIT('h4)
	) name21023 (
		\ethreg1_RXHASH1_2_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31535_
	);
	LUT2 #(
		.INIT('h2)
	) name21024 (
		_w31507_,
		_w31534_,
		_w31536_
	);
	LUT2 #(
		.INIT('h4)
	) name21025 (
		_w31535_,
		_w31536_,
		_w31537_
	);
	LUT2 #(
		.INIT('h1)
	) name21026 (
		\ethreg1_RXHASH0_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31538_
	);
	LUT2 #(
		.INIT('h4)
	) name21027 (
		\ethreg1_RXHASH1_3_DataOut_reg[4]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31539_
	);
	LUT2 #(
		.INIT('h2)
	) name21028 (
		_w31502_,
		_w31538_,
		_w31540_
	);
	LUT2 #(
		.INIT('h4)
	) name21029 (
		_w31539_,
		_w31540_,
		_w31541_
	);
	LUT2 #(
		.INIT('h1)
	) name21030 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31529_,
		_w31542_
	);
	LUT2 #(
		.INIT('h1)
	) name21031 (
		_w31533_,
		_w31537_,
		_w31543_
	);
	LUT2 #(
		.INIT('h4)
	) name21032 (
		_w31541_,
		_w31543_,
		_w31544_
	);
	LUT2 #(
		.INIT('h8)
	) name21033 (
		_w31542_,
		_w31544_,
		_w31545_
	);
	LUT2 #(
		.INIT('h1)
	) name21034 (
		_w31525_,
		_w31545_,
		_w31546_
	);
	LUT2 #(
		.INIT('h1)
	) name21035 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		_w31546_,
		_w31547_
	);
	LUT2 #(
		.INIT('h1)
	) name21036 (
		\ethreg1_RXHASH0_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31548_
	);
	LUT2 #(
		.INIT('h4)
	) name21037 (
		\ethreg1_RXHASH1_0_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31549_
	);
	LUT2 #(
		.INIT('h2)
	) name21038 (
		_w31512_,
		_w31548_,
		_w31550_
	);
	LUT2 #(
		.INIT('h4)
	) name21039 (
		_w31549_,
		_w31550_,
		_w31551_
	);
	LUT2 #(
		.INIT('h1)
	) name21040 (
		\ethreg1_RXHASH0_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31552_
	);
	LUT2 #(
		.INIT('h4)
	) name21041 (
		\ethreg1_RXHASH1_1_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31553_
	);
	LUT2 #(
		.INIT('h2)
	) name21042 (
		_w31517_,
		_w31552_,
		_w31554_
	);
	LUT2 #(
		.INIT('h4)
	) name21043 (
		_w31553_,
		_w31554_,
		_w31555_
	);
	LUT2 #(
		.INIT('h1)
	) name21044 (
		\ethreg1_RXHASH0_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31556_
	);
	LUT2 #(
		.INIT('h4)
	) name21045 (
		\ethreg1_RXHASH1_2_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31557_
	);
	LUT2 #(
		.INIT('h2)
	) name21046 (
		_w31507_,
		_w31556_,
		_w31558_
	);
	LUT2 #(
		.INIT('h4)
	) name21047 (
		_w31557_,
		_w31558_,
		_w31559_
	);
	LUT2 #(
		.INIT('h1)
	) name21048 (
		\ethreg1_RXHASH0_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31560_
	);
	LUT2 #(
		.INIT('h4)
	) name21049 (
		\ethreg1_RXHASH1_3_DataOut_reg[6]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31561_
	);
	LUT2 #(
		.INIT('h2)
	) name21050 (
		_w31502_,
		_w31560_,
		_w31562_
	);
	LUT2 #(
		.INIT('h4)
	) name21051 (
		_w31561_,
		_w31562_,
		_w31563_
	);
	LUT2 #(
		.INIT('h1)
	) name21052 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31551_,
		_w31564_
	);
	LUT2 #(
		.INIT('h1)
	) name21053 (
		_w31555_,
		_w31559_,
		_w31565_
	);
	LUT2 #(
		.INIT('h4)
	) name21054 (
		_w31563_,
		_w31565_,
		_w31566_
	);
	LUT2 #(
		.INIT('h8)
	) name21055 (
		_w31564_,
		_w31566_,
		_w31567_
	);
	LUT2 #(
		.INIT('h1)
	) name21056 (
		\ethreg1_RXHASH0_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31568_
	);
	LUT2 #(
		.INIT('h4)
	) name21057 (
		\ethreg1_RXHASH1_0_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31569_
	);
	LUT2 #(
		.INIT('h2)
	) name21058 (
		_w31512_,
		_w31568_,
		_w31570_
	);
	LUT2 #(
		.INIT('h4)
	) name21059 (
		_w31569_,
		_w31570_,
		_w31571_
	);
	LUT2 #(
		.INIT('h1)
	) name21060 (
		\ethreg1_RXHASH0_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31572_
	);
	LUT2 #(
		.INIT('h4)
	) name21061 (
		\ethreg1_RXHASH1_2_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31573_
	);
	LUT2 #(
		.INIT('h2)
	) name21062 (
		_w31507_,
		_w31572_,
		_w31574_
	);
	LUT2 #(
		.INIT('h4)
	) name21063 (
		_w31573_,
		_w31574_,
		_w31575_
	);
	LUT2 #(
		.INIT('h1)
	) name21064 (
		\ethreg1_RXHASH0_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31576_
	);
	LUT2 #(
		.INIT('h4)
	) name21065 (
		\ethreg1_RXHASH1_3_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31577_
	);
	LUT2 #(
		.INIT('h2)
	) name21066 (
		_w31502_,
		_w31576_,
		_w31578_
	);
	LUT2 #(
		.INIT('h4)
	) name21067 (
		_w31577_,
		_w31578_,
		_w31579_
	);
	LUT2 #(
		.INIT('h1)
	) name21068 (
		\ethreg1_RXHASH0_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31580_
	);
	LUT2 #(
		.INIT('h4)
	) name21069 (
		\ethreg1_RXHASH1_1_DataOut_reg[7]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31581_
	);
	LUT2 #(
		.INIT('h2)
	) name21070 (
		_w31517_,
		_w31580_,
		_w31582_
	);
	LUT2 #(
		.INIT('h4)
	) name21071 (
		_w31581_,
		_w31582_,
		_w31583_
	);
	LUT2 #(
		.INIT('h2)
	) name21072 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31571_,
		_w31584_
	);
	LUT2 #(
		.INIT('h1)
	) name21073 (
		_w31575_,
		_w31579_,
		_w31585_
	);
	LUT2 #(
		.INIT('h4)
	) name21074 (
		_w31583_,
		_w31585_,
		_w31586_
	);
	LUT2 #(
		.INIT('h8)
	) name21075 (
		_w31584_,
		_w31586_,
		_w31587_
	);
	LUT2 #(
		.INIT('h1)
	) name21076 (
		_w31567_,
		_w31587_,
		_w31588_
	);
	LUT2 #(
		.INIT('h2)
	) name21077 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		_w31588_,
		_w31589_
	);
	LUT2 #(
		.INIT('h2)
	) name21078 (
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w31547_,
		_w31590_
	);
	LUT2 #(
		.INIT('h4)
	) name21079 (
		_w31589_,
		_w31590_,
		_w31591_
	);
	LUT2 #(
		.INIT('h1)
	) name21080 (
		\ethreg1_RXHASH0_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31592_
	);
	LUT2 #(
		.INIT('h4)
	) name21081 (
		\ethreg1_RXHASH1_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31593_
	);
	LUT2 #(
		.INIT('h2)
	) name21082 (
		_w31512_,
		_w31592_,
		_w31594_
	);
	LUT2 #(
		.INIT('h4)
	) name21083 (
		_w31593_,
		_w31594_,
		_w31595_
	);
	LUT2 #(
		.INIT('h1)
	) name21084 (
		\ethreg1_RXHASH0_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31596_
	);
	LUT2 #(
		.INIT('h4)
	) name21085 (
		\ethreg1_RXHASH1_1_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31597_
	);
	LUT2 #(
		.INIT('h2)
	) name21086 (
		_w31517_,
		_w31596_,
		_w31598_
	);
	LUT2 #(
		.INIT('h4)
	) name21087 (
		_w31597_,
		_w31598_,
		_w31599_
	);
	LUT2 #(
		.INIT('h1)
	) name21088 (
		\ethreg1_RXHASH0_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31600_
	);
	LUT2 #(
		.INIT('h4)
	) name21089 (
		\ethreg1_RXHASH1_3_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31601_
	);
	LUT2 #(
		.INIT('h2)
	) name21090 (
		_w31502_,
		_w31600_,
		_w31602_
	);
	LUT2 #(
		.INIT('h4)
	) name21091 (
		_w31601_,
		_w31602_,
		_w31603_
	);
	LUT2 #(
		.INIT('h1)
	) name21092 (
		\ethreg1_RXHASH0_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31604_
	);
	LUT2 #(
		.INIT('h4)
	) name21093 (
		\ethreg1_RXHASH1_2_DataOut_reg[1]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31605_
	);
	LUT2 #(
		.INIT('h2)
	) name21094 (
		_w31507_,
		_w31604_,
		_w31606_
	);
	LUT2 #(
		.INIT('h4)
	) name21095 (
		_w31605_,
		_w31606_,
		_w31607_
	);
	LUT2 #(
		.INIT('h2)
	) name21096 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31595_,
		_w31608_
	);
	LUT2 #(
		.INIT('h1)
	) name21097 (
		_w31599_,
		_w31603_,
		_w31609_
	);
	LUT2 #(
		.INIT('h4)
	) name21098 (
		_w31607_,
		_w31609_,
		_w31610_
	);
	LUT2 #(
		.INIT('h8)
	) name21099 (
		_w31608_,
		_w31610_,
		_w31611_
	);
	LUT2 #(
		.INIT('h1)
	) name21100 (
		\ethreg1_RXHASH0_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31612_
	);
	LUT2 #(
		.INIT('h4)
	) name21101 (
		\ethreg1_RXHASH1_3_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31613_
	);
	LUT2 #(
		.INIT('h2)
	) name21102 (
		_w31502_,
		_w31612_,
		_w31614_
	);
	LUT2 #(
		.INIT('h4)
	) name21103 (
		_w31613_,
		_w31614_,
		_w31615_
	);
	LUT2 #(
		.INIT('h1)
	) name21104 (
		\ethreg1_RXHASH0_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31616_
	);
	LUT2 #(
		.INIT('h4)
	) name21105 (
		\ethreg1_RXHASH1_2_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31617_
	);
	LUT2 #(
		.INIT('h2)
	) name21106 (
		_w31507_,
		_w31616_,
		_w31618_
	);
	LUT2 #(
		.INIT('h4)
	) name21107 (
		_w31617_,
		_w31618_,
		_w31619_
	);
	LUT2 #(
		.INIT('h1)
	) name21108 (
		\ethreg1_RXHASH0_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31620_
	);
	LUT2 #(
		.INIT('h4)
	) name21109 (
		\ethreg1_RXHASH1_1_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31621_
	);
	LUT2 #(
		.INIT('h2)
	) name21110 (
		_w31517_,
		_w31620_,
		_w31622_
	);
	LUT2 #(
		.INIT('h4)
	) name21111 (
		_w31621_,
		_w31622_,
		_w31623_
	);
	LUT2 #(
		.INIT('h1)
	) name21112 (
		\ethreg1_RXHASH0_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31624_
	);
	LUT2 #(
		.INIT('h4)
	) name21113 (
		\ethreg1_RXHASH1_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31625_
	);
	LUT2 #(
		.INIT('h2)
	) name21114 (
		_w31512_,
		_w31624_,
		_w31626_
	);
	LUT2 #(
		.INIT('h4)
	) name21115 (
		_w31625_,
		_w31626_,
		_w31627_
	);
	LUT2 #(
		.INIT('h1)
	) name21116 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31615_,
		_w31628_
	);
	LUT2 #(
		.INIT('h1)
	) name21117 (
		_w31619_,
		_w31623_,
		_w31629_
	);
	LUT2 #(
		.INIT('h4)
	) name21118 (
		_w31627_,
		_w31629_,
		_w31630_
	);
	LUT2 #(
		.INIT('h8)
	) name21119 (
		_w31628_,
		_w31630_,
		_w31631_
	);
	LUT2 #(
		.INIT('h1)
	) name21120 (
		_w31611_,
		_w31631_,
		_w31632_
	);
	LUT2 #(
		.INIT('h1)
	) name21121 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		_w31632_,
		_w31633_
	);
	LUT2 #(
		.INIT('h1)
	) name21122 (
		\ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31634_
	);
	LUT2 #(
		.INIT('h4)
	) name21123 (
		\ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31635_
	);
	LUT2 #(
		.INIT('h2)
	) name21124 (
		_w31517_,
		_w31634_,
		_w31636_
	);
	LUT2 #(
		.INIT('h4)
	) name21125 (
		_w31635_,
		_w31636_,
		_w31637_
	);
	LUT2 #(
		.INIT('h1)
	) name21126 (
		\ethreg1_RXHASH0_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31638_
	);
	LUT2 #(
		.INIT('h4)
	) name21127 (
		\ethreg1_RXHASH1_3_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31639_
	);
	LUT2 #(
		.INIT('h2)
	) name21128 (
		_w31502_,
		_w31638_,
		_w31640_
	);
	LUT2 #(
		.INIT('h4)
	) name21129 (
		_w31639_,
		_w31640_,
		_w31641_
	);
	LUT2 #(
		.INIT('h1)
	) name21130 (
		\ethreg1_RXHASH0_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31642_
	);
	LUT2 #(
		.INIT('h4)
	) name21131 (
		\ethreg1_RXHASH1_2_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31643_
	);
	LUT2 #(
		.INIT('h2)
	) name21132 (
		_w31507_,
		_w31642_,
		_w31644_
	);
	LUT2 #(
		.INIT('h4)
	) name21133 (
		_w31643_,
		_w31644_,
		_w31645_
	);
	LUT2 #(
		.INIT('h1)
	) name21134 (
		\ethreg1_RXHASH0_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31646_
	);
	LUT2 #(
		.INIT('h4)
	) name21135 (
		\ethreg1_RXHASH1_0_DataOut_reg[2]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31647_
	);
	LUT2 #(
		.INIT('h2)
	) name21136 (
		_w31512_,
		_w31646_,
		_w31648_
	);
	LUT2 #(
		.INIT('h4)
	) name21137 (
		_w31647_,
		_w31648_,
		_w31649_
	);
	LUT2 #(
		.INIT('h1)
	) name21138 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31637_,
		_w31650_
	);
	LUT2 #(
		.INIT('h1)
	) name21139 (
		_w31641_,
		_w31645_,
		_w31651_
	);
	LUT2 #(
		.INIT('h4)
	) name21140 (
		_w31649_,
		_w31651_,
		_w31652_
	);
	LUT2 #(
		.INIT('h8)
	) name21141 (
		_w31650_,
		_w31652_,
		_w31653_
	);
	LUT2 #(
		.INIT('h1)
	) name21142 (
		\ethreg1_RXHASH0_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31654_
	);
	LUT2 #(
		.INIT('h4)
	) name21143 (
		\ethreg1_RXHASH1_1_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31655_
	);
	LUT2 #(
		.INIT('h2)
	) name21144 (
		_w31517_,
		_w31654_,
		_w31656_
	);
	LUT2 #(
		.INIT('h4)
	) name21145 (
		_w31655_,
		_w31656_,
		_w31657_
	);
	LUT2 #(
		.INIT('h1)
	) name21146 (
		\ethreg1_RXHASH0_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31658_
	);
	LUT2 #(
		.INIT('h4)
	) name21147 (
		\ethreg1_RXHASH1_2_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31659_
	);
	LUT2 #(
		.INIT('h2)
	) name21148 (
		_w31507_,
		_w31658_,
		_w31660_
	);
	LUT2 #(
		.INIT('h4)
	) name21149 (
		_w31659_,
		_w31660_,
		_w31661_
	);
	LUT2 #(
		.INIT('h1)
	) name21150 (
		\ethreg1_RXHASH0_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31662_
	);
	LUT2 #(
		.INIT('h4)
	) name21151 (
		\ethreg1_RXHASH1_3_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31663_
	);
	LUT2 #(
		.INIT('h2)
	) name21152 (
		_w31502_,
		_w31662_,
		_w31664_
	);
	LUT2 #(
		.INIT('h4)
	) name21153 (
		_w31663_,
		_w31664_,
		_w31665_
	);
	LUT2 #(
		.INIT('h1)
	) name21154 (
		\ethreg1_RXHASH0_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31666_
	);
	LUT2 #(
		.INIT('h4)
	) name21155 (
		\ethreg1_RXHASH1_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w31667_
	);
	LUT2 #(
		.INIT('h2)
	) name21156 (
		_w31512_,
		_w31666_,
		_w31668_
	);
	LUT2 #(
		.INIT('h4)
	) name21157 (
		_w31667_,
		_w31668_,
		_w31669_
	);
	LUT2 #(
		.INIT('h2)
	) name21158 (
		\rxethmac1_CrcHash_reg[0]/P0001 ,
		_w31657_,
		_w31670_
	);
	LUT2 #(
		.INIT('h1)
	) name21159 (
		_w31661_,
		_w31665_,
		_w31671_
	);
	LUT2 #(
		.INIT('h4)
	) name21160 (
		_w31669_,
		_w31671_,
		_w31672_
	);
	LUT2 #(
		.INIT('h8)
	) name21161 (
		_w31670_,
		_w31672_,
		_w31673_
	);
	LUT2 #(
		.INIT('h1)
	) name21162 (
		_w31653_,
		_w31673_,
		_w31674_
	);
	LUT2 #(
		.INIT('h2)
	) name21163 (
		\rxethmac1_CrcHash_reg[1]/P0001 ,
		_w31674_,
		_w31675_
	);
	LUT2 #(
		.INIT('h1)
	) name21164 (
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w31633_,
		_w31676_
	);
	LUT2 #(
		.INIT('h4)
	) name21165 (
		_w31675_,
		_w31676_,
		_w31677_
	);
	LUT2 #(
		.INIT('h2)
	) name21166 (
		_w31500_,
		_w31591_,
		_w31678_
	);
	LUT2 #(
		.INIT('h4)
	) name21167 (
		_w31677_,
		_w31678_,
		_w31679_
	);
	LUT2 #(
		.INIT('h2)
	) name21168 (
		_w12477_,
		_w31501_,
		_w31680_
	);
	LUT2 #(
		.INIT('h4)
	) name21169 (
		_w31679_,
		_w31680_,
		_w31681_
	);
	LUT2 #(
		.INIT('h8)
	) name21170 (
		\wb_sel_i[0]_pad ,
		_w22942_,
		_w31682_
	);
	LUT2 #(
		.INIT('h4)
	) name21171 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w31683_
	);
	LUT2 #(
		.INIT('h8)
	) name21172 (
		_w31682_,
		_w31683_,
		_w31684_
	);
	LUT2 #(
		.INIT('h1)
	) name21173 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w31685_
	);
	LUT2 #(
		.INIT('h4)
	) name21174 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w31686_
	);
	LUT2 #(
		.INIT('h1)
	) name21175 (
		\wb_dat_i[0]_pad ,
		\wb_dat_i[1]_pad ,
		_w31687_
	);
	LUT2 #(
		.INIT('h1)
	) name21176 (
		\wb_dat_i[2]_pad ,
		\wb_dat_i[3]_pad ,
		_w31688_
	);
	LUT2 #(
		.INIT('h1)
	) name21177 (
		\wb_dat_i[4]_pad ,
		\wb_dat_i[5]_pad ,
		_w31689_
	);
	LUT2 #(
		.INIT('h4)
	) name21178 (
		\wb_dat_i[6]_pad ,
		_w31689_,
		_w31690_
	);
	LUT2 #(
		.INIT('h8)
	) name21179 (
		_w31687_,
		_w31688_,
		_w31691_
	);
	LUT2 #(
		.INIT('h8)
	) name21180 (
		_w31690_,
		_w31691_,
		_w31692_
	);
	LUT2 #(
		.INIT('h2)
	) name21181 (
		\wb_dat_i[7]_pad ,
		_w31692_,
		_w31693_
	);
	LUT2 #(
		.INIT('h1)
	) name21182 (
		\wb_adr_i[6]_pad ,
		\wb_dat_i[10]_pad ,
		_w31694_
	);
	LUT2 #(
		.INIT('h1)
	) name21183 (
		\wb_dat_i[11]_pad ,
		\wb_dat_i[12]_pad ,
		_w31695_
	);
	LUT2 #(
		.INIT('h1)
	) name21184 (
		\wb_dat_i[13]_pad ,
		\wb_dat_i[14]_pad ,
		_w31696_
	);
	LUT2 #(
		.INIT('h1)
	) name21185 (
		\wb_dat_i[15]_pad ,
		\wb_dat_i[16]_pad ,
		_w31697_
	);
	LUT2 #(
		.INIT('h1)
	) name21186 (
		\wb_dat_i[17]_pad ,
		\wb_dat_i[18]_pad ,
		_w31698_
	);
	LUT2 #(
		.INIT('h1)
	) name21187 (
		\wb_dat_i[19]_pad ,
		\wb_dat_i[20]_pad ,
		_w31699_
	);
	LUT2 #(
		.INIT('h1)
	) name21188 (
		\wb_dat_i[21]_pad ,
		\wb_dat_i[22]_pad ,
		_w31700_
	);
	LUT2 #(
		.INIT('h1)
	) name21189 (
		\wb_dat_i[23]_pad ,
		\wb_dat_i[24]_pad ,
		_w31701_
	);
	LUT2 #(
		.INIT('h1)
	) name21190 (
		\wb_dat_i[25]_pad ,
		\wb_dat_i[26]_pad ,
		_w31702_
	);
	LUT2 #(
		.INIT('h1)
	) name21191 (
		\wb_dat_i[27]_pad ,
		\wb_dat_i[28]_pad ,
		_w31703_
	);
	LUT2 #(
		.INIT('h1)
	) name21192 (
		\wb_dat_i[29]_pad ,
		\wb_dat_i[30]_pad ,
		_w31704_
	);
	LUT2 #(
		.INIT('h1)
	) name21193 (
		\wb_dat_i[31]_pad ,
		\wb_dat_i[8]_pad ,
		_w31705_
	);
	LUT2 #(
		.INIT('h4)
	) name21194 (
		\wb_dat_i[9]_pad ,
		_w31705_,
		_w31706_
	);
	LUT2 #(
		.INIT('h8)
	) name21195 (
		_w31703_,
		_w31704_,
		_w31707_
	);
	LUT2 #(
		.INIT('h8)
	) name21196 (
		_w31701_,
		_w31702_,
		_w31708_
	);
	LUT2 #(
		.INIT('h8)
	) name21197 (
		_w31699_,
		_w31700_,
		_w31709_
	);
	LUT2 #(
		.INIT('h8)
	) name21198 (
		_w31697_,
		_w31698_,
		_w31710_
	);
	LUT2 #(
		.INIT('h8)
	) name21199 (
		_w31695_,
		_w31696_,
		_w31711_
	);
	LUT2 #(
		.INIT('h8)
	) name21200 (
		_w31685_,
		_w31694_,
		_w31712_
	);
	LUT2 #(
		.INIT('h8)
	) name21201 (
		_w31686_,
		_w31712_,
		_w31713_
	);
	LUT2 #(
		.INIT('h8)
	) name21202 (
		_w31710_,
		_w31711_,
		_w31714_
	);
	LUT2 #(
		.INIT('h8)
	) name21203 (
		_w31708_,
		_w31709_,
		_w31715_
	);
	LUT2 #(
		.INIT('h8)
	) name21204 (
		_w31706_,
		_w31707_,
		_w31716_
	);
	LUT2 #(
		.INIT('h8)
	) name21205 (
		_w22962_,
		_w31716_,
		_w31717_
	);
	LUT2 #(
		.INIT('h8)
	) name21206 (
		_w31714_,
		_w31715_,
		_w31718_
	);
	LUT2 #(
		.INIT('h8)
	) name21207 (
		_w31713_,
		_w31718_,
		_w31719_
	);
	LUT2 #(
		.INIT('h4)
	) name21208 (
		_w31693_,
		_w31717_,
		_w31720_
	);
	LUT2 #(
		.INIT('h8)
	) name21209 (
		_w31719_,
		_w31720_,
		_w31721_
	);
	LUT2 #(
		.INIT('h8)
	) name21210 (
		_w31684_,
		_w31721_,
		_w31722_
	);
	LUT2 #(
		.INIT('h4)
	) name21211 (
		\rxethmac1_crcrx_Crc_reg[17]/NET0131 ,
		_w10580_,
		_w31723_
	);
	LUT2 #(
		.INIT('h2)
	) name21212 (
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w11244_,
		_w31724_
	);
	LUT2 #(
		.INIT('h4)
	) name21213 (
		\rxethmac1_crcrx_Crc_reg[2]/NET0131 ,
		_w11244_,
		_w31725_
	);
	LUT2 #(
		.INIT('h2)
	) name21214 (
		_w10580_,
		_w31724_,
		_w31726_
	);
	LUT2 #(
		.INIT('h4)
	) name21215 (
		_w31725_,
		_w31726_,
		_w31727_
	);
	LUT2 #(
		.INIT('h8)
	) name21216 (
		\maccontrol1_receivecontrol1_OpCodeOK_reg/NET0131 ,
		\maccontrol1_receivecontrol1_TypeLengthOK_reg/NET0131 ,
		_w31728_
	);
	LUT2 #(
		.INIT('h8)
	) name21217 (
		_w11831_,
		_w31728_,
		_w31729_
	);
	LUT2 #(
		.INIT('h8)
	) name21218 (
		_w12646_,
		_w31729_,
		_w31730_
	);
	LUT2 #(
		.INIT('h8)
	) name21219 (
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w31730_,
		_w31731_
	);
	LUT2 #(
		.INIT('h1)
	) name21220 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w31731_,
		_w31732_
	);
	LUT2 #(
		.INIT('h1)
	) name21221 (
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w31732_,
		_w31733_
	);
	LUT2 #(
		.INIT('h2)
	) name21222 (
		\txethmac1_txcrc_Crc_reg[0]/NET0131 ,
		_w12458_,
		_w31734_
	);
	LUT2 #(
		.INIT('h4)
	) name21223 (
		\txethmac1_txcrc_Crc_reg[0]/NET0131 ,
		_w12458_,
		_w31735_
	);
	LUT2 #(
		.INIT('h2)
	) name21224 (
		_w11181_,
		_w31734_,
		_w31736_
	);
	LUT2 #(
		.INIT('h4)
	) name21225 (
		_w31735_,
		_w31736_,
		_w31737_
	);
	LUT2 #(
		.INIT('h8)
	) name21226 (
		_w11908_,
		_w31226_,
		_w31738_
	);
	LUT2 #(
		.INIT('h1)
	) name21227 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 ,
		_w31738_,
		_w31739_
	);
	LUT2 #(
		.INIT('h4)
	) name21228 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w31738_,
		_w31740_
	);
	LUT2 #(
		.INIT('h1)
	) name21229 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31739_,
		_w31741_
	);
	LUT2 #(
		.INIT('h4)
	) name21230 (
		_w31740_,
		_w31741_,
		_w31742_
	);
	LUT2 #(
		.INIT('h8)
	) name21231 (
		_w11831_,
		_w31226_,
		_w31743_
	);
	LUT2 #(
		.INIT('h1)
	) name21232 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 ,
		_w31743_,
		_w31744_
	);
	LUT2 #(
		.INIT('h4)
	) name21233 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w31743_,
		_w31745_
	);
	LUT2 #(
		.INIT('h1)
	) name21234 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31744_,
		_w31746_
	);
	LUT2 #(
		.INIT('h4)
	) name21235 (
		_w31745_,
		_w31746_,
		_w31747_
	);
	LUT2 #(
		.INIT('h1)
	) name21236 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 ,
		_w31743_,
		_w31748_
	);
	LUT2 #(
		.INIT('h4)
	) name21237 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w31743_,
		_w31749_
	);
	LUT2 #(
		.INIT('h1)
	) name21238 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31748_,
		_w31750_
	);
	LUT2 #(
		.INIT('h4)
	) name21239 (
		_w31749_,
		_w31750_,
		_w31751_
	);
	LUT2 #(
		.INIT('h1)
	) name21240 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 ,
		_w31743_,
		_w31752_
	);
	LUT2 #(
		.INIT('h4)
	) name21241 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w31743_,
		_w31753_
	);
	LUT2 #(
		.INIT('h1)
	) name21242 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31752_,
		_w31754_
	);
	LUT2 #(
		.INIT('h4)
	) name21243 (
		_w31753_,
		_w31754_,
		_w31755_
	);
	LUT2 #(
		.INIT('h1)
	) name21244 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 ,
		_w31743_,
		_w31756_
	);
	LUT2 #(
		.INIT('h4)
	) name21245 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w31743_,
		_w31757_
	);
	LUT2 #(
		.INIT('h1)
	) name21246 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31756_,
		_w31758_
	);
	LUT2 #(
		.INIT('h4)
	) name21247 (
		_w31757_,
		_w31758_,
		_w31759_
	);
	LUT2 #(
		.INIT('h1)
	) name21248 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 ,
		_w31743_,
		_w31760_
	);
	LUT2 #(
		.INIT('h4)
	) name21249 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w31743_,
		_w31761_
	);
	LUT2 #(
		.INIT('h1)
	) name21250 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31760_,
		_w31762_
	);
	LUT2 #(
		.INIT('h4)
	) name21251 (
		_w31761_,
		_w31762_,
		_w31763_
	);
	LUT2 #(
		.INIT('h1)
	) name21252 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 ,
		_w31743_,
		_w31764_
	);
	LUT2 #(
		.INIT('h4)
	) name21253 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w31743_,
		_w31765_
	);
	LUT2 #(
		.INIT('h1)
	) name21254 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31764_,
		_w31766_
	);
	LUT2 #(
		.INIT('h4)
	) name21255 (
		_w31765_,
		_w31766_,
		_w31767_
	);
	LUT2 #(
		.INIT('h1)
	) name21256 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 ,
		_w31738_,
		_w31768_
	);
	LUT2 #(
		.INIT('h4)
	) name21257 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w31738_,
		_w31769_
	);
	LUT2 #(
		.INIT('h1)
	) name21258 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31768_,
		_w31770_
	);
	LUT2 #(
		.INIT('h4)
	) name21259 (
		_w31769_,
		_w31770_,
		_w31771_
	);
	LUT2 #(
		.INIT('h1)
	) name21260 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 ,
		_w31738_,
		_w31772_
	);
	LUT2 #(
		.INIT('h4)
	) name21261 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w31738_,
		_w31773_
	);
	LUT2 #(
		.INIT('h1)
	) name21262 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31772_,
		_w31774_
	);
	LUT2 #(
		.INIT('h4)
	) name21263 (
		_w31773_,
		_w31774_,
		_w31775_
	);
	LUT2 #(
		.INIT('h1)
	) name21264 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 ,
		_w31738_,
		_w31776_
	);
	LUT2 #(
		.INIT('h4)
	) name21265 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w31738_,
		_w31777_
	);
	LUT2 #(
		.INIT('h1)
	) name21266 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31776_,
		_w31778_
	);
	LUT2 #(
		.INIT('h4)
	) name21267 (
		_w31777_,
		_w31778_,
		_w31779_
	);
	LUT2 #(
		.INIT('h1)
	) name21268 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 ,
		_w31738_,
		_w31780_
	);
	LUT2 #(
		.INIT('h4)
	) name21269 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w31738_,
		_w31781_
	);
	LUT2 #(
		.INIT('h1)
	) name21270 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31780_,
		_w31782_
	);
	LUT2 #(
		.INIT('h4)
	) name21271 (
		_w31781_,
		_w31782_,
		_w31783_
	);
	LUT2 #(
		.INIT('h1)
	) name21272 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 ,
		_w31738_,
		_w31784_
	);
	LUT2 #(
		.INIT('h4)
	) name21273 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w31738_,
		_w31785_
	);
	LUT2 #(
		.INIT('h1)
	) name21274 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31784_,
		_w31786_
	);
	LUT2 #(
		.INIT('h4)
	) name21275 (
		_w31785_,
		_w31786_,
		_w31787_
	);
	LUT2 #(
		.INIT('h1)
	) name21276 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 ,
		_w31738_,
		_w31788_
	);
	LUT2 #(
		.INIT('h4)
	) name21277 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w31738_,
		_w31789_
	);
	LUT2 #(
		.INIT('h1)
	) name21278 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31788_,
		_w31790_
	);
	LUT2 #(
		.INIT('h4)
	) name21279 (
		_w31789_,
		_w31790_,
		_w31791_
	);
	LUT2 #(
		.INIT('h1)
	) name21280 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 ,
		_w31738_,
		_w31792_
	);
	LUT2 #(
		.INIT('h4)
	) name21281 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w31738_,
		_w31793_
	);
	LUT2 #(
		.INIT('h1)
	) name21282 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31792_,
		_w31794_
	);
	LUT2 #(
		.INIT('h4)
	) name21283 (
		_w31793_,
		_w31794_,
		_w31795_
	);
	LUT2 #(
		.INIT('h1)
	) name21284 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 ,
		_w31743_,
		_w31796_
	);
	LUT2 #(
		.INIT('h4)
	) name21285 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w31743_,
		_w31797_
	);
	LUT2 #(
		.INIT('h1)
	) name21286 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31796_,
		_w31798_
	);
	LUT2 #(
		.INIT('h4)
	) name21287 (
		_w31797_,
		_w31798_,
		_w31799_
	);
	LUT2 #(
		.INIT('h1)
	) name21288 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 ,
		_w31743_,
		_w31800_
	);
	LUT2 #(
		.INIT('h4)
	) name21289 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w31743_,
		_w31801_
	);
	LUT2 #(
		.INIT('h1)
	) name21290 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31800_,
		_w31802_
	);
	LUT2 #(
		.INIT('h4)
	) name21291 (
		_w31801_,
		_w31802_,
		_w31803_
	);
	LUT2 #(
		.INIT('h1)
	) name21292 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		_w12632_,
		_w31804_
	);
	LUT2 #(
		.INIT('h2)
	) name21293 (
		\m_wb_sel_o[1]_pad ,
		_w31330_,
		_w31805_
	);
	LUT2 #(
		.INIT('h1)
	) name21294 (
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w12632_,
		_w31806_
	);
	LUT2 #(
		.INIT('h2)
	) name21295 (
		_w12573_,
		_w31806_,
		_w31807_
	);
	LUT2 #(
		.INIT('h4)
	) name21296 (
		_w31804_,
		_w31807_,
		_w31808_
	);
	LUT2 #(
		.INIT('h4)
	) name21297 (
		_w31805_,
		_w31808_,
		_w31809_
	);
	LUT2 #(
		.INIT('h2)
	) name21298 (
		\m_wb_sel_o[2]_pad ,
		_w31330_,
		_w31810_
	);
	LUT2 #(
		.INIT('h2)
	) name21299 (
		_w31807_,
		_w31810_,
		_w31811_
	);
	LUT2 #(
		.INIT('h2)
	) name21300 (
		\m_wb_sel_o[3]_pad ,
		_w31330_,
		_w31812_
	);
	LUT2 #(
		.INIT('h1)
	) name21301 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		\wishbone_RxPointerLSB_rst_reg[1]/NET0131 ,
		_w31813_
	);
	LUT2 #(
		.INIT('h4)
	) name21302 (
		_w12632_,
		_w31813_,
		_w31814_
	);
	LUT2 #(
		.INIT('h2)
	) name21303 (
		_w12573_,
		_w31814_,
		_w31815_
	);
	LUT2 #(
		.INIT('h4)
	) name21304 (
		_w31812_,
		_w31815_,
		_w31816_
	);
	LUT2 #(
		.INIT('h2)
	) name21305 (
		_w31321_,
		_w31328_,
		_w31817_
	);
	LUT2 #(
		.INIT('h2)
	) name21306 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w31817_,
		_w31818_
	);
	LUT2 #(
		.INIT('h2)
	) name21307 (
		_w12632_,
		_w31818_,
		_w31819_
	);
	LUT2 #(
		.INIT('h2)
	) name21308 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w31817_,
		_w31820_
	);
	LUT2 #(
		.INIT('h2)
	) name21309 (
		_w12573_,
		_w31820_,
		_w31821_
	);
	LUT2 #(
		.INIT('h1)
	) name21310 (
		\macstatus1_RxColWindow_reg/NET0131 ,
		\rxethmac1_rxstatem1_StateIdle_reg/NET0131 ,
		_w31822_
	);
	LUT2 #(
		.INIT('h2)
	) name21311 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w31823_
	);
	LUT2 #(
		.INIT('h4)
	) name21312 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[1]/NET0131 ,
		_w31824_
	);
	LUT2 #(
		.INIT('h1)
	) name21313 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w31825_
	);
	LUT2 #(
		.INIT('h8)
	) name21314 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_ByteCnt_reg[0]/NET0131 ,
		_w31826_
	);
	LUT2 #(
		.INIT('h1)
	) name21315 (
		_w31825_,
		_w31826_,
		_w31827_
	);
	LUT2 #(
		.INIT('h1)
	) name21316 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w31828_
	);
	LUT2 #(
		.INIT('h8)
	) name21317 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		_w11492_,
		_w31829_
	);
	LUT2 #(
		.INIT('h1)
	) name21318 (
		_w31828_,
		_w31829_,
		_w31830_
	);
	LUT2 #(
		.INIT('h1)
	) name21319 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		_w11495_,
		_w31831_
	);
	LUT2 #(
		.INIT('h8)
	) name21320 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		_w11495_,
		_w31832_
	);
	LUT2 #(
		.INIT('h1)
	) name21321 (
		_w31831_,
		_w31832_,
		_w31833_
	);
	LUT2 #(
		.INIT('h1)
	) name21322 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w31834_
	);
	LUT2 #(
		.INIT('h8)
	) name21323 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		_w11506_,
		_w31835_
	);
	LUT2 #(
		.INIT('h1)
	) name21324 (
		_w31834_,
		_w31835_,
		_w31836_
	);
	LUT2 #(
		.INIT('h2)
	) name21325 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w31837_
	);
	LUT2 #(
		.INIT('h4)
	) name21326 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		_w11488_,
		_w31838_
	);
	LUT2 #(
		.INIT('h4)
	) name21327 (
		mcoll_pad_i_pad,
		\rxethmac1_rxstatem1_StateData1_reg/NET0131 ,
		_w31839_
	);
	LUT2 #(
		.INIT('h4)
	) name21328 (
		_w31823_,
		_w31839_,
		_w31840_
	);
	LUT2 #(
		.INIT('h4)
	) name21329 (
		_w31824_,
		_w31840_,
		_w31841_
	);
	LUT2 #(
		.INIT('h4)
	) name21330 (
		_w31827_,
		_w31841_,
		_w31842_
	);
	LUT2 #(
		.INIT('h4)
	) name21331 (
		_w31833_,
		_w31842_,
		_w31843_
	);
	LUT2 #(
		.INIT('h4)
	) name21332 (
		_w31830_,
		_w31843_,
		_w31844_
	);
	LUT2 #(
		.INIT('h1)
	) name21333 (
		_w31837_,
		_w31838_,
		_w31845_
	);
	LUT2 #(
		.INIT('h8)
	) name21334 (
		_w31844_,
		_w31845_,
		_w31846_
	);
	LUT2 #(
		.INIT('h4)
	) name21335 (
		_w31836_,
		_w31846_,
		_w31847_
	);
	LUT2 #(
		.INIT('h1)
	) name21336 (
		_w31822_,
		_w31847_,
		_w31848_
	);
	LUT2 #(
		.INIT('h8)
	) name21337 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w31849_
	);
	LUT2 #(
		.INIT('h2)
	) name21338 (
		_w10576_,
		_w31849_,
		_w31850_
	);
	LUT2 #(
		.INIT('h8)
	) name21339 (
		_w10527_,
		_w31850_,
		_w31851_
	);
	LUT2 #(
		.INIT('h2)
	) name21340 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w31851_,
		_w31852_
	);
	LUT2 #(
		.INIT('h2)
	) name21341 (
		\rxethmac1_DelayData_reg/NET0131 ,
		_w31852_,
		_w31853_
	);
	LUT2 #(
		.INIT('h8)
	) name21342 (
		\rxethmac1_RxData_d_reg[0]/NET0131 ,
		_w31853_,
		_w31854_
	);
	LUT2 #(
		.INIT('h8)
	) name21343 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		_w31852_,
		_w31855_
	);
	LUT2 #(
		.INIT('h1)
	) name21344 (
		_w31854_,
		_w31855_,
		_w31856_
	);
	LUT2 #(
		.INIT('h1)
	) name21345 (
		\txethmac1_StopExcessiveDeferOccured_reg/NET0131 ,
		_w11095_,
		_w31857_
	);
	LUT2 #(
		.INIT('h1)
	) name21346 (
		_w11099_,
		_w31857_,
		_w31858_
	);
	LUT2 #(
		.INIT('h8)
	) name21347 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrmWAddr_reg/NET0131 ,
		_w31227_,
		_w31859_
	);
	LUT2 #(
		.INIT('h8)
	) name21348 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[0]/NET0131 ,
		_w31859_,
		_w31860_
	);
	LUT2 #(
		.INIT('h1)
	) name21349 (
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w31859_,
		_w31861_
	);
	LUT2 #(
		.INIT('h8)
	) name21350 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[0]/NET0131 ,
		_w31861_,
		_w31862_
	);
	LUT2 #(
		.INIT('h1)
	) name21351 (
		_w31860_,
		_w31862_,
		_w31863_
	);
	LUT2 #(
		.INIT('h8)
	) name21352 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[10]/NET0131 ,
		_w31859_,
		_w31864_
	);
	LUT2 #(
		.INIT('h8)
	) name21353 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[10]/NET0131 ,
		_w31861_,
		_w31865_
	);
	LUT2 #(
		.INIT('h1)
	) name21354 (
		_w31864_,
		_w31865_,
		_w31866_
	);
	LUT2 #(
		.INIT('h8)
	) name21355 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[11]/NET0131 ,
		_w31859_,
		_w31867_
	);
	LUT2 #(
		.INIT('h8)
	) name21356 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[11]/NET0131 ,
		_w31861_,
		_w31868_
	);
	LUT2 #(
		.INIT('h1)
	) name21357 (
		_w31867_,
		_w31868_,
		_w31869_
	);
	LUT2 #(
		.INIT('h8)
	) name21358 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[12]/NET0131 ,
		_w31859_,
		_w31870_
	);
	LUT2 #(
		.INIT('h8)
	) name21359 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[12]/NET0131 ,
		_w31861_,
		_w31871_
	);
	LUT2 #(
		.INIT('h1)
	) name21360 (
		_w31870_,
		_w31871_,
		_w31872_
	);
	LUT2 #(
		.INIT('h8)
	) name21361 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[13]/NET0131 ,
		_w31859_,
		_w31873_
	);
	LUT2 #(
		.INIT('h8)
	) name21362 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[13]/NET0131 ,
		_w31861_,
		_w31874_
	);
	LUT2 #(
		.INIT('h1)
	) name21363 (
		_w31873_,
		_w31874_,
		_w31875_
	);
	LUT2 #(
		.INIT('h8)
	) name21364 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[15]/NET0131 ,
		_w31859_,
		_w31876_
	);
	LUT2 #(
		.INIT('h8)
	) name21365 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[15]/NET0131 ,
		_w31861_,
		_w31877_
	);
	LUT2 #(
		.INIT('h1)
	) name21366 (
		_w31876_,
		_w31877_,
		_w31878_
	);
	LUT2 #(
		.INIT('h8)
	) name21367 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[14]/NET0131 ,
		_w31859_,
		_w31879_
	);
	LUT2 #(
		.INIT('h8)
	) name21368 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[14]/NET0131 ,
		_w31861_,
		_w31880_
	);
	LUT2 #(
		.INIT('h1)
	) name21369 (
		_w31879_,
		_w31880_,
		_w31881_
	);
	LUT2 #(
		.INIT('h8)
	) name21370 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[1]/NET0131 ,
		_w31859_,
		_w31882_
	);
	LUT2 #(
		.INIT('h8)
	) name21371 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[1]/NET0131 ,
		_w31861_,
		_w31883_
	);
	LUT2 #(
		.INIT('h1)
	) name21372 (
		_w31882_,
		_w31883_,
		_w31884_
	);
	LUT2 #(
		.INIT('h8)
	) name21373 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[2]/NET0131 ,
		_w31859_,
		_w31885_
	);
	LUT2 #(
		.INIT('h8)
	) name21374 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[2]/NET0131 ,
		_w31861_,
		_w31886_
	);
	LUT2 #(
		.INIT('h1)
	) name21375 (
		_w31885_,
		_w31886_,
		_w31887_
	);
	LUT2 #(
		.INIT('h8)
	) name21376 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[3]/NET0131 ,
		_w31859_,
		_w31888_
	);
	LUT2 #(
		.INIT('h8)
	) name21377 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[3]/NET0131 ,
		_w31861_,
		_w31889_
	);
	LUT2 #(
		.INIT('h1)
	) name21378 (
		_w31888_,
		_w31889_,
		_w31890_
	);
	LUT2 #(
		.INIT('h8)
	) name21379 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[4]/NET0131 ,
		_w31859_,
		_w31891_
	);
	LUT2 #(
		.INIT('h8)
	) name21380 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[4]/NET0131 ,
		_w31861_,
		_w31892_
	);
	LUT2 #(
		.INIT('h1)
	) name21381 (
		_w31891_,
		_w31892_,
		_w31893_
	);
	LUT2 #(
		.INIT('h8)
	) name21382 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[5]/NET0131 ,
		_w31859_,
		_w31894_
	);
	LUT2 #(
		.INIT('h8)
	) name21383 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[5]/NET0131 ,
		_w31861_,
		_w31895_
	);
	LUT2 #(
		.INIT('h1)
	) name21384 (
		_w31894_,
		_w31895_,
		_w31896_
	);
	LUT2 #(
		.INIT('h8)
	) name21385 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[6]/NET0131 ,
		_w31859_,
		_w31897_
	);
	LUT2 #(
		.INIT('h8)
	) name21386 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[6]/NET0131 ,
		_w31861_,
		_w31898_
	);
	LUT2 #(
		.INIT('h1)
	) name21387 (
		_w31897_,
		_w31898_,
		_w31899_
	);
	LUT2 #(
		.INIT('h8)
	) name21388 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[7]/NET0131 ,
		_w31859_,
		_w31900_
	);
	LUT2 #(
		.INIT('h8)
	) name21389 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[7]/NET0131 ,
		_w31861_,
		_w31901_
	);
	LUT2 #(
		.INIT('h1)
	) name21390 (
		_w31900_,
		_w31901_,
		_w31902_
	);
	LUT2 #(
		.INIT('h8)
	) name21391 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[8]/NET0131 ,
		_w31859_,
		_w31903_
	);
	LUT2 #(
		.INIT('h8)
	) name21392 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[8]/NET0131 ,
		_w31861_,
		_w31904_
	);
	LUT2 #(
		.INIT('h1)
	) name21393 (
		_w31903_,
		_w31904_,
		_w31905_
	);
	LUT2 #(
		.INIT('h8)
	) name21394 (
		\maccontrol1_receivecontrol1_AssembledTimerValue_reg[9]/NET0131 ,
		_w31859_,
		_w31906_
	);
	LUT2 #(
		.INIT('h8)
	) name21395 (
		\maccontrol1_receivecontrol1_LatchedTimerValue_reg[9]/NET0131 ,
		_w31861_,
		_w31907_
	);
	LUT2 #(
		.INIT('h1)
	) name21396 (
		_w31906_,
		_w31907_,
		_w31908_
	);
	LUT2 #(
		.INIT('h4)
	) name21397 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w15143_,
		_w31909_
	);
	LUT2 #(
		.INIT('h1)
	) name21398 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		_w31909_,
		_w31910_
	);
	LUT2 #(
		.INIT('h8)
	) name21399 (
		\wishbone_RxValidBytes_reg[0]/NET0131 ,
		_w31909_,
		_w31911_
	);
	LUT2 #(
		.INIT('h1)
	) name21400 (
		_w31910_,
		_w31911_,
		_w31912_
	);
	LUT2 #(
		.INIT('h1)
	) name21401 (
		_w15138_,
		_w31912_,
		_w31913_
	);
	LUT2 #(
		.INIT('h8)
	) name21402 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		_w15138_,
		_w31914_
	);
	LUT2 #(
		.INIT('h1)
	) name21403 (
		_w31913_,
		_w31914_,
		_w31915_
	);
	LUT2 #(
		.INIT('h2)
	) name21404 (
		\wishbone_RxValidBytes_reg[1]/NET0131 ,
		_w31909_,
		_w31916_
	);
	LUT2 #(
		.INIT('h8)
	) name21405 (
		_w15152_,
		_w31909_,
		_w31917_
	);
	LUT2 #(
		.INIT('h1)
	) name21406 (
		_w31916_,
		_w31917_,
		_w31918_
	);
	LUT2 #(
		.INIT('h1)
	) name21407 (
		_w15138_,
		_w31918_,
		_w31919_
	);
	LUT2 #(
		.INIT('h2)
	) name21408 (
		_w15138_,
		_w31240_,
		_w31920_
	);
	LUT2 #(
		.INIT('h1)
	) name21409 (
		_w31919_,
		_w31920_,
		_w31921_
	);
	LUT2 #(
		.INIT('h2)
	) name21410 (
		\miim1_shftrg_ShiftReg_reg[0]/NET0131 ,
		_w31401_,
		_w31922_
	);
	LUT2 #(
		.INIT('h2)
	) name21411 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[1]/NET0131 ,
		_w31418_,
		_w31923_
	);
	LUT2 #(
		.INIT('h8)
	) name21412 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[0]/NET0131 ,
		_w31428_,
		_w31924_
	);
	LUT2 #(
		.INIT('h8)
	) name21413 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[0]/NET0131 ,
		_w31430_,
		_w31925_
	);
	LUT2 #(
		.INIT('h8)
	) name21414 (
		md_pad_i_pad,
		_w31426_,
		_w31926_
	);
	LUT2 #(
		.INIT('h1)
	) name21415 (
		_w31923_,
		_w31924_,
		_w31927_
	);
	LUT2 #(
		.INIT('h4)
	) name21416 (
		_w31925_,
		_w31927_,
		_w31928_
	);
	LUT2 #(
		.INIT('h4)
	) name21417 (
		_w31926_,
		_w31928_,
		_w31929_
	);
	LUT2 #(
		.INIT('h2)
	) name21418 (
		_w31401_,
		_w31929_,
		_w31930_
	);
	LUT2 #(
		.INIT('h1)
	) name21419 (
		_w31922_,
		_w31930_,
		_w31931_
	);
	LUT2 #(
		.INIT('h8)
	) name21420 (
		\ethreg1_MIITX_DATA_0_DataOut_reg[7]/NET0131 ,
		_w31430_,
		_w31932_
	);
	LUT2 #(
		.INIT('h8)
	) name21421 (
		\ethreg1_MIIADDRESS_0_DataOut_reg[0]/NET0131 ,
		_w31424_,
		_w31933_
	);
	LUT2 #(
		.INIT('h8)
	) name21422 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[7]/NET0131 ,
		_w31428_,
		_w31934_
	);
	LUT2 #(
		.INIT('h8)
	) name21423 (
		\miim1_shftrg_ShiftReg_reg[6]/NET0131 ,
		_w31426_,
		_w31935_
	);
	LUT2 #(
		.INIT('h1)
	) name21424 (
		_w31932_,
		_w31933_,
		_w31936_
	);
	LUT2 #(
		.INIT('h4)
	) name21425 (
		_w31934_,
		_w31936_,
		_w31937_
	);
	LUT2 #(
		.INIT('h4)
	) name21426 (
		_w31935_,
		_w31937_,
		_w31938_
	);
	LUT2 #(
		.INIT('h2)
	) name21427 (
		_w31401_,
		_w31938_,
		_w31939_
	);
	LUT2 #(
		.INIT('h2)
	) name21428 (
		\miim1_shftrg_ShiftReg_reg[7]/NET0131 ,
		_w31401_,
		_w31940_
	);
	LUT2 #(
		.INIT('h1)
	) name21429 (
		_w31939_,
		_w31940_,
		_w31941_
	);
	LUT2 #(
		.INIT('h1)
	) name21430 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		_w12561_,
		_w31942_
	);
	LUT2 #(
		.INIT('h2)
	) name21431 (
		\wishbone_tx_burst_cnt_reg[0]/NET0131 ,
		_w31359_,
		_w31943_
	);
	LUT2 #(
		.INIT('h1)
	) name21432 (
		_w31942_,
		_w31943_,
		_w31944_
	);
	LUT2 #(
		.INIT('h2)
	) name21433 (
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w31360_,
		_w31945_
	);
	LUT2 #(
		.INIT('h1)
	) name21434 (
		_w31361_,
		_w31945_,
		_w31946_
	);
	LUT2 #(
		.INIT('h2)
	) name21435 (
		_w12561_,
		_w31946_,
		_w31947_
	);
	LUT2 #(
		.INIT('h8)
	) name21436 (
		\wishbone_tx_burst_cnt_reg[2]/NET0131 ,
		_w31359_,
		_w31948_
	);
	LUT2 #(
		.INIT('h1)
	) name21437 (
		_w31947_,
		_w31948_,
		_w31949_
	);
	LUT2 #(
		.INIT('h4)
	) name21438 (
		\wishbone_SyncRxStartFrm_q2_reg/NET0131 ,
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		_w31950_
	);
	LUT2 #(
		.INIT('h1)
	) name21439 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w31951_
	);
	LUT2 #(
		.INIT('h1)
	) name21440 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w31952_
	);
	LUT2 #(
		.INIT('h8)
	) name21441 (
		_w31951_,
		_w31952_,
		_w31953_
	);
	LUT2 #(
		.INIT('h1)
	) name21442 (
		_w31950_,
		_w31953_,
		_w31954_
	);
	LUT2 #(
		.INIT('h2)
	) name21443 (
		\wishbone_rx_fifo_fifo_reg[0][0]/P0001 ,
		_w31954_,
		_w31955_
	);
	LUT2 #(
		.INIT('h4)
	) name21444 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w31956_
	);
	LUT2 #(
		.INIT('h2)
	) name21445 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w31957_
	);
	LUT2 #(
		.INIT('h8)
	) name21446 (
		_w31956_,
		_w31957_,
		_w31958_
	);
	LUT2 #(
		.INIT('h8)
	) name21447 (
		\wishbone_rx_fifo_fifo_reg[6][0]/P0001 ,
		_w31958_,
		_w31959_
	);
	LUT2 #(
		.INIT('h4)
	) name21448 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w31960_
	);
	LUT2 #(
		.INIT('h8)
	) name21449 (
		_w31956_,
		_w31960_,
		_w31961_
	);
	LUT2 #(
		.INIT('h8)
	) name21450 (
		\wishbone_rx_fifo_fifo_reg[10][0]/P0001 ,
		_w31961_,
		_w31962_
	);
	LUT2 #(
		.INIT('h8)
	) name21451 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w31963_
	);
	LUT2 #(
		.INIT('h8)
	) name21452 (
		_w31957_,
		_w31963_,
		_w31964_
	);
	LUT2 #(
		.INIT('h8)
	) name21453 (
		\wishbone_rx_fifo_fifo_reg[7][0]/P0001 ,
		_w31964_,
		_w31965_
	);
	LUT2 #(
		.INIT('h8)
	) name21454 (
		_w31951_,
		_w31957_,
		_w31966_
	);
	LUT2 #(
		.INIT('h8)
	) name21455 (
		\wishbone_rx_fifo_fifo_reg[4][0]/P0001 ,
		_w31966_,
		_w31967_
	);
	LUT2 #(
		.INIT('h8)
	) name21456 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w31968_
	);
	LUT2 #(
		.INIT('h8)
	) name21457 (
		_w31963_,
		_w31968_,
		_w31969_
	);
	LUT2 #(
		.INIT('h8)
	) name21458 (
		\wishbone_rx_fifo_fifo_reg[15][0]/P0001 ,
		_w31969_,
		_w31970_
	);
	LUT2 #(
		.INIT('h2)
	) name21459 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w31971_
	);
	LUT2 #(
		.INIT('h8)
	) name21460 (
		_w31960_,
		_w31971_,
		_w31972_
	);
	LUT2 #(
		.INIT('h8)
	) name21461 (
		\wishbone_rx_fifo_fifo_reg[9][0]/P0001 ,
		_w31972_,
		_w31973_
	);
	LUT2 #(
		.INIT('h8)
	) name21462 (
		_w31951_,
		_w31960_,
		_w31974_
	);
	LUT2 #(
		.INIT('h8)
	) name21463 (
		\wishbone_rx_fifo_fifo_reg[8][0]/P0001 ,
		_w31974_,
		_w31975_
	);
	LUT2 #(
		.INIT('h8)
	) name21464 (
		_w31952_,
		_w31971_,
		_w31976_
	);
	LUT2 #(
		.INIT('h8)
	) name21465 (
		\wishbone_rx_fifo_fifo_reg[1][0]/P0001 ,
		_w31976_,
		_w31977_
	);
	LUT2 #(
		.INIT('h8)
	) name21466 (
		_w31952_,
		_w31956_,
		_w31978_
	);
	LUT2 #(
		.INIT('h8)
	) name21467 (
		\wishbone_rx_fifo_fifo_reg[2][0]/P0001 ,
		_w31978_,
		_w31979_
	);
	LUT2 #(
		.INIT('h8)
	) name21468 (
		_w31957_,
		_w31971_,
		_w31980_
	);
	LUT2 #(
		.INIT('h8)
	) name21469 (
		\wishbone_rx_fifo_fifo_reg[5][0]/P0001 ,
		_w31980_,
		_w31981_
	);
	LUT2 #(
		.INIT('h8)
	) name21470 (
		_w31956_,
		_w31968_,
		_w31982_
	);
	LUT2 #(
		.INIT('h8)
	) name21471 (
		\wishbone_rx_fifo_fifo_reg[14][0]/P0001 ,
		_w31982_,
		_w31983_
	);
	LUT2 #(
		.INIT('h8)
	) name21472 (
		_w31951_,
		_w31968_,
		_w31984_
	);
	LUT2 #(
		.INIT('h8)
	) name21473 (
		\wishbone_rx_fifo_fifo_reg[12][0]/P0001 ,
		_w31984_,
		_w31985_
	);
	LUT2 #(
		.INIT('h8)
	) name21474 (
		_w31968_,
		_w31971_,
		_w31986_
	);
	LUT2 #(
		.INIT('h8)
	) name21475 (
		\wishbone_rx_fifo_fifo_reg[13][0]/P0001 ,
		_w31986_,
		_w31987_
	);
	LUT2 #(
		.INIT('h8)
	) name21476 (
		_w31960_,
		_w31963_,
		_w31988_
	);
	LUT2 #(
		.INIT('h8)
	) name21477 (
		\wishbone_rx_fifo_fifo_reg[11][0]/P0001 ,
		_w31988_,
		_w31989_
	);
	LUT2 #(
		.INIT('h8)
	) name21478 (
		_w31952_,
		_w31963_,
		_w31990_
	);
	LUT2 #(
		.INIT('h8)
	) name21479 (
		\wishbone_rx_fifo_fifo_reg[3][0]/P0001 ,
		_w31990_,
		_w31991_
	);
	LUT2 #(
		.INIT('h1)
	) name21480 (
		_w31959_,
		_w31962_,
		_w31992_
	);
	LUT2 #(
		.INIT('h1)
	) name21481 (
		_w31965_,
		_w31967_,
		_w31993_
	);
	LUT2 #(
		.INIT('h1)
	) name21482 (
		_w31970_,
		_w31973_,
		_w31994_
	);
	LUT2 #(
		.INIT('h1)
	) name21483 (
		_w31975_,
		_w31977_,
		_w31995_
	);
	LUT2 #(
		.INIT('h1)
	) name21484 (
		_w31979_,
		_w31981_,
		_w31996_
	);
	LUT2 #(
		.INIT('h1)
	) name21485 (
		_w31983_,
		_w31985_,
		_w31997_
	);
	LUT2 #(
		.INIT('h1)
	) name21486 (
		_w31987_,
		_w31989_,
		_w31998_
	);
	LUT2 #(
		.INIT('h4)
	) name21487 (
		_w31991_,
		_w31998_,
		_w31999_
	);
	LUT2 #(
		.INIT('h8)
	) name21488 (
		_w31996_,
		_w31997_,
		_w32000_
	);
	LUT2 #(
		.INIT('h8)
	) name21489 (
		_w31994_,
		_w31995_,
		_w32001_
	);
	LUT2 #(
		.INIT('h8)
	) name21490 (
		_w31992_,
		_w31993_,
		_w32002_
	);
	LUT2 #(
		.INIT('h8)
	) name21491 (
		_w32001_,
		_w32002_,
		_w32003_
	);
	LUT2 #(
		.INIT('h8)
	) name21492 (
		_w31999_,
		_w32000_,
		_w32004_
	);
	LUT2 #(
		.INIT('h8)
	) name21493 (
		_w32003_,
		_w32004_,
		_w32005_
	);
	LUT2 #(
		.INIT('h1)
	) name21494 (
		_w31950_,
		_w32005_,
		_w32006_
	);
	LUT2 #(
		.INIT('h1)
	) name21495 (
		_w31955_,
		_w32006_,
		_w32007_
	);
	LUT2 #(
		.INIT('h8)
	) name21496 (
		\wishbone_rx_fifo_fifo_reg[5][10]/P0001 ,
		_w31980_,
		_w32008_
	);
	LUT2 #(
		.INIT('h8)
	) name21497 (
		\wishbone_rx_fifo_fifo_reg[7][10]/P0001 ,
		_w31964_,
		_w32009_
	);
	LUT2 #(
		.INIT('h8)
	) name21498 (
		\wishbone_rx_fifo_fifo_reg[1][10]/P0001 ,
		_w31976_,
		_w32010_
	);
	LUT2 #(
		.INIT('h8)
	) name21499 (
		\wishbone_rx_fifo_fifo_reg[11][10]/P0001 ,
		_w31988_,
		_w32011_
	);
	LUT2 #(
		.INIT('h8)
	) name21500 (
		\wishbone_rx_fifo_fifo_reg[3][10]/P0001 ,
		_w31990_,
		_w32012_
	);
	LUT2 #(
		.INIT('h8)
	) name21501 (
		\wishbone_rx_fifo_fifo_reg[6][10]/P0001 ,
		_w31958_,
		_w32013_
	);
	LUT2 #(
		.INIT('h8)
	) name21502 (
		\wishbone_rx_fifo_fifo_reg[15][10]/P0001 ,
		_w31969_,
		_w32014_
	);
	LUT2 #(
		.INIT('h8)
	) name21503 (
		\wishbone_rx_fifo_fifo_reg[14][10]/P0001 ,
		_w31982_,
		_w32015_
	);
	LUT2 #(
		.INIT('h8)
	) name21504 (
		\wishbone_rx_fifo_fifo_reg[2][10]/P0001 ,
		_w31978_,
		_w32016_
	);
	LUT2 #(
		.INIT('h8)
	) name21505 (
		\wishbone_rx_fifo_fifo_reg[8][10]/P0001 ,
		_w31974_,
		_w32017_
	);
	LUT2 #(
		.INIT('h8)
	) name21506 (
		\wishbone_rx_fifo_fifo_reg[4][10]/P0001 ,
		_w31966_,
		_w32018_
	);
	LUT2 #(
		.INIT('h8)
	) name21507 (
		\wishbone_rx_fifo_fifo_reg[12][10]/P0001 ,
		_w31984_,
		_w32019_
	);
	LUT2 #(
		.INIT('h8)
	) name21508 (
		\wishbone_rx_fifo_fifo_reg[10][10]/P0001 ,
		_w31961_,
		_w32020_
	);
	LUT2 #(
		.INIT('h8)
	) name21509 (
		\wishbone_rx_fifo_fifo_reg[9][10]/P0001 ,
		_w31972_,
		_w32021_
	);
	LUT2 #(
		.INIT('h8)
	) name21510 (
		\wishbone_rx_fifo_fifo_reg[13][10]/P0001 ,
		_w31986_,
		_w32022_
	);
	LUT2 #(
		.INIT('h1)
	) name21511 (
		_w31950_,
		_w32008_,
		_w32023_
	);
	LUT2 #(
		.INIT('h1)
	) name21512 (
		_w32009_,
		_w32010_,
		_w32024_
	);
	LUT2 #(
		.INIT('h1)
	) name21513 (
		_w32011_,
		_w32012_,
		_w32025_
	);
	LUT2 #(
		.INIT('h1)
	) name21514 (
		_w32013_,
		_w32014_,
		_w32026_
	);
	LUT2 #(
		.INIT('h1)
	) name21515 (
		_w32015_,
		_w32016_,
		_w32027_
	);
	LUT2 #(
		.INIT('h1)
	) name21516 (
		_w32017_,
		_w32018_,
		_w32028_
	);
	LUT2 #(
		.INIT('h1)
	) name21517 (
		_w32019_,
		_w32020_,
		_w32029_
	);
	LUT2 #(
		.INIT('h1)
	) name21518 (
		_w32021_,
		_w32022_,
		_w32030_
	);
	LUT2 #(
		.INIT('h8)
	) name21519 (
		_w32029_,
		_w32030_,
		_w32031_
	);
	LUT2 #(
		.INIT('h8)
	) name21520 (
		_w32027_,
		_w32028_,
		_w32032_
	);
	LUT2 #(
		.INIT('h8)
	) name21521 (
		_w32025_,
		_w32026_,
		_w32033_
	);
	LUT2 #(
		.INIT('h8)
	) name21522 (
		_w32023_,
		_w32024_,
		_w32034_
	);
	LUT2 #(
		.INIT('h8)
	) name21523 (
		_w32033_,
		_w32034_,
		_w32035_
	);
	LUT2 #(
		.INIT('h8)
	) name21524 (
		_w32031_,
		_w32032_,
		_w32036_
	);
	LUT2 #(
		.INIT('h8)
	) name21525 (
		_w32035_,
		_w32036_,
		_w32037_
	);
	LUT2 #(
		.INIT('h4)
	) name21526 (
		\wishbone_rx_fifo_fifo_reg[0][10]/P0001 ,
		_w31950_,
		_w32038_
	);
	LUT2 #(
		.INIT('h1)
	) name21527 (
		_w32037_,
		_w32038_,
		_w32039_
	);
	LUT2 #(
		.INIT('h8)
	) name21528 (
		\wishbone_rx_fifo_fifo_reg[0][10]/P0001 ,
		_w31953_,
		_w32040_
	);
	LUT2 #(
		.INIT('h1)
	) name21529 (
		_w32039_,
		_w32040_,
		_w32041_
	);
	LUT2 #(
		.INIT('h2)
	) name21530 (
		\wishbone_rx_fifo_fifo_reg[0][11]/P0001 ,
		_w31954_,
		_w32042_
	);
	LUT2 #(
		.INIT('h8)
	) name21531 (
		\wishbone_rx_fifo_fifo_reg[6][11]/P0001 ,
		_w31958_,
		_w32043_
	);
	LUT2 #(
		.INIT('h8)
	) name21532 (
		\wishbone_rx_fifo_fifo_reg[12][11]/P0001 ,
		_w31984_,
		_w32044_
	);
	LUT2 #(
		.INIT('h8)
	) name21533 (
		\wishbone_rx_fifo_fifo_reg[8][11]/P0001 ,
		_w31974_,
		_w32045_
	);
	LUT2 #(
		.INIT('h8)
	) name21534 (
		\wishbone_rx_fifo_fifo_reg[11][11]/P0001 ,
		_w31988_,
		_w32046_
	);
	LUT2 #(
		.INIT('h8)
	) name21535 (
		\wishbone_rx_fifo_fifo_reg[5][11]/P0001 ,
		_w31980_,
		_w32047_
	);
	LUT2 #(
		.INIT('h8)
	) name21536 (
		\wishbone_rx_fifo_fifo_reg[9][11]/P0001 ,
		_w31972_,
		_w32048_
	);
	LUT2 #(
		.INIT('h8)
	) name21537 (
		\wishbone_rx_fifo_fifo_reg[10][11]/P0001 ,
		_w31961_,
		_w32049_
	);
	LUT2 #(
		.INIT('h8)
	) name21538 (
		\wishbone_rx_fifo_fifo_reg[13][11]/P0001 ,
		_w31986_,
		_w32050_
	);
	LUT2 #(
		.INIT('h8)
	) name21539 (
		\wishbone_rx_fifo_fifo_reg[1][11]/P0001 ,
		_w31976_,
		_w32051_
	);
	LUT2 #(
		.INIT('h8)
	) name21540 (
		\wishbone_rx_fifo_fifo_reg[15][11]/P0001 ,
		_w31969_,
		_w32052_
	);
	LUT2 #(
		.INIT('h8)
	) name21541 (
		\wishbone_rx_fifo_fifo_reg[4][11]/P0001 ,
		_w31966_,
		_w32053_
	);
	LUT2 #(
		.INIT('h8)
	) name21542 (
		\wishbone_rx_fifo_fifo_reg[3][11]/P0001 ,
		_w31990_,
		_w32054_
	);
	LUT2 #(
		.INIT('h8)
	) name21543 (
		\wishbone_rx_fifo_fifo_reg[7][11]/P0001 ,
		_w31964_,
		_w32055_
	);
	LUT2 #(
		.INIT('h8)
	) name21544 (
		\wishbone_rx_fifo_fifo_reg[14][11]/P0001 ,
		_w31982_,
		_w32056_
	);
	LUT2 #(
		.INIT('h8)
	) name21545 (
		\wishbone_rx_fifo_fifo_reg[2][11]/P0001 ,
		_w31978_,
		_w32057_
	);
	LUT2 #(
		.INIT('h1)
	) name21546 (
		_w32043_,
		_w32044_,
		_w32058_
	);
	LUT2 #(
		.INIT('h1)
	) name21547 (
		_w32045_,
		_w32046_,
		_w32059_
	);
	LUT2 #(
		.INIT('h1)
	) name21548 (
		_w32047_,
		_w32048_,
		_w32060_
	);
	LUT2 #(
		.INIT('h1)
	) name21549 (
		_w32049_,
		_w32050_,
		_w32061_
	);
	LUT2 #(
		.INIT('h1)
	) name21550 (
		_w32051_,
		_w32052_,
		_w32062_
	);
	LUT2 #(
		.INIT('h1)
	) name21551 (
		_w32053_,
		_w32054_,
		_w32063_
	);
	LUT2 #(
		.INIT('h1)
	) name21552 (
		_w32055_,
		_w32056_,
		_w32064_
	);
	LUT2 #(
		.INIT('h4)
	) name21553 (
		_w32057_,
		_w32064_,
		_w32065_
	);
	LUT2 #(
		.INIT('h8)
	) name21554 (
		_w32062_,
		_w32063_,
		_w32066_
	);
	LUT2 #(
		.INIT('h8)
	) name21555 (
		_w32060_,
		_w32061_,
		_w32067_
	);
	LUT2 #(
		.INIT('h8)
	) name21556 (
		_w32058_,
		_w32059_,
		_w32068_
	);
	LUT2 #(
		.INIT('h8)
	) name21557 (
		_w32067_,
		_w32068_,
		_w32069_
	);
	LUT2 #(
		.INIT('h8)
	) name21558 (
		_w32065_,
		_w32066_,
		_w32070_
	);
	LUT2 #(
		.INIT('h8)
	) name21559 (
		_w32069_,
		_w32070_,
		_w32071_
	);
	LUT2 #(
		.INIT('h1)
	) name21560 (
		_w31950_,
		_w32071_,
		_w32072_
	);
	LUT2 #(
		.INIT('h1)
	) name21561 (
		_w32042_,
		_w32072_,
		_w32073_
	);
	LUT2 #(
		.INIT('h8)
	) name21562 (
		\wishbone_rx_fifo_fifo_reg[3][12]/P0001 ,
		_w31990_,
		_w32074_
	);
	LUT2 #(
		.INIT('h8)
	) name21563 (
		\wishbone_rx_fifo_fifo_reg[14][12]/P0001 ,
		_w31982_,
		_w32075_
	);
	LUT2 #(
		.INIT('h8)
	) name21564 (
		\wishbone_rx_fifo_fifo_reg[2][12]/P0001 ,
		_w31978_,
		_w32076_
	);
	LUT2 #(
		.INIT('h8)
	) name21565 (
		\wishbone_rx_fifo_fifo_reg[5][12]/P0001 ,
		_w31980_,
		_w32077_
	);
	LUT2 #(
		.INIT('h8)
	) name21566 (
		\wishbone_rx_fifo_fifo_reg[11][12]/P0001 ,
		_w31988_,
		_w32078_
	);
	LUT2 #(
		.INIT('h8)
	) name21567 (
		\wishbone_rx_fifo_fifo_reg[10][12]/P0001 ,
		_w31961_,
		_w32079_
	);
	LUT2 #(
		.INIT('h8)
	) name21568 (
		\wishbone_rx_fifo_fifo_reg[1][12]/P0001 ,
		_w31976_,
		_w32080_
	);
	LUT2 #(
		.INIT('h8)
	) name21569 (
		\wishbone_rx_fifo_fifo_reg[4][12]/P0001 ,
		_w31966_,
		_w32081_
	);
	LUT2 #(
		.INIT('h8)
	) name21570 (
		\wishbone_rx_fifo_fifo_reg[8][12]/P0001 ,
		_w31974_,
		_w32082_
	);
	LUT2 #(
		.INIT('h8)
	) name21571 (
		\wishbone_rx_fifo_fifo_reg[15][12]/P0001 ,
		_w31969_,
		_w32083_
	);
	LUT2 #(
		.INIT('h8)
	) name21572 (
		\wishbone_rx_fifo_fifo_reg[7][12]/P0001 ,
		_w31964_,
		_w32084_
	);
	LUT2 #(
		.INIT('h8)
	) name21573 (
		\wishbone_rx_fifo_fifo_reg[9][12]/P0001 ,
		_w31972_,
		_w32085_
	);
	LUT2 #(
		.INIT('h8)
	) name21574 (
		\wishbone_rx_fifo_fifo_reg[12][12]/P0001 ,
		_w31984_,
		_w32086_
	);
	LUT2 #(
		.INIT('h8)
	) name21575 (
		\wishbone_rx_fifo_fifo_reg[6][12]/P0001 ,
		_w31958_,
		_w32087_
	);
	LUT2 #(
		.INIT('h8)
	) name21576 (
		\wishbone_rx_fifo_fifo_reg[13][12]/P0001 ,
		_w31986_,
		_w32088_
	);
	LUT2 #(
		.INIT('h1)
	) name21577 (
		_w31950_,
		_w32074_,
		_w32089_
	);
	LUT2 #(
		.INIT('h1)
	) name21578 (
		_w32075_,
		_w32076_,
		_w32090_
	);
	LUT2 #(
		.INIT('h1)
	) name21579 (
		_w32077_,
		_w32078_,
		_w32091_
	);
	LUT2 #(
		.INIT('h1)
	) name21580 (
		_w32079_,
		_w32080_,
		_w32092_
	);
	LUT2 #(
		.INIT('h1)
	) name21581 (
		_w32081_,
		_w32082_,
		_w32093_
	);
	LUT2 #(
		.INIT('h1)
	) name21582 (
		_w32083_,
		_w32084_,
		_w32094_
	);
	LUT2 #(
		.INIT('h1)
	) name21583 (
		_w32085_,
		_w32086_,
		_w32095_
	);
	LUT2 #(
		.INIT('h1)
	) name21584 (
		_w32087_,
		_w32088_,
		_w32096_
	);
	LUT2 #(
		.INIT('h8)
	) name21585 (
		_w32095_,
		_w32096_,
		_w32097_
	);
	LUT2 #(
		.INIT('h8)
	) name21586 (
		_w32093_,
		_w32094_,
		_w32098_
	);
	LUT2 #(
		.INIT('h8)
	) name21587 (
		_w32091_,
		_w32092_,
		_w32099_
	);
	LUT2 #(
		.INIT('h8)
	) name21588 (
		_w32089_,
		_w32090_,
		_w32100_
	);
	LUT2 #(
		.INIT('h8)
	) name21589 (
		_w32099_,
		_w32100_,
		_w32101_
	);
	LUT2 #(
		.INIT('h8)
	) name21590 (
		_w32097_,
		_w32098_,
		_w32102_
	);
	LUT2 #(
		.INIT('h8)
	) name21591 (
		_w32101_,
		_w32102_,
		_w32103_
	);
	LUT2 #(
		.INIT('h4)
	) name21592 (
		\wishbone_rx_fifo_fifo_reg[0][12]/P0001 ,
		_w31950_,
		_w32104_
	);
	LUT2 #(
		.INIT('h1)
	) name21593 (
		_w32103_,
		_w32104_,
		_w32105_
	);
	LUT2 #(
		.INIT('h8)
	) name21594 (
		\wishbone_rx_fifo_fifo_reg[0][12]/P0001 ,
		_w31953_,
		_w32106_
	);
	LUT2 #(
		.INIT('h1)
	) name21595 (
		_w32105_,
		_w32106_,
		_w32107_
	);
	LUT2 #(
		.INIT('h2)
	) name21596 (
		\wishbone_rx_fifo_fifo_reg[0][13]/P0001 ,
		_w31954_,
		_w32108_
	);
	LUT2 #(
		.INIT('h8)
	) name21597 (
		\wishbone_rx_fifo_fifo_reg[3][13]/P0001 ,
		_w31990_,
		_w32109_
	);
	LUT2 #(
		.INIT('h8)
	) name21598 (
		\wishbone_rx_fifo_fifo_reg[9][13]/P0001 ,
		_w31972_,
		_w32110_
	);
	LUT2 #(
		.INIT('h8)
	) name21599 (
		\wishbone_rx_fifo_fifo_reg[8][13]/P0001 ,
		_w31974_,
		_w32111_
	);
	LUT2 #(
		.INIT('h8)
	) name21600 (
		\wishbone_rx_fifo_fifo_reg[7][13]/P0001 ,
		_w31964_,
		_w32112_
	);
	LUT2 #(
		.INIT('h8)
	) name21601 (
		\wishbone_rx_fifo_fifo_reg[10][13]/P0001 ,
		_w31961_,
		_w32113_
	);
	LUT2 #(
		.INIT('h8)
	) name21602 (
		\wishbone_rx_fifo_fifo_reg[5][13]/P0001 ,
		_w31980_,
		_w32114_
	);
	LUT2 #(
		.INIT('h8)
	) name21603 (
		\wishbone_rx_fifo_fifo_reg[14][13]/P0001 ,
		_w31982_,
		_w32115_
	);
	LUT2 #(
		.INIT('h8)
	) name21604 (
		\wishbone_rx_fifo_fifo_reg[4][13]/P0001 ,
		_w31966_,
		_w32116_
	);
	LUT2 #(
		.INIT('h8)
	) name21605 (
		\wishbone_rx_fifo_fifo_reg[1][13]/P0001 ,
		_w31976_,
		_w32117_
	);
	LUT2 #(
		.INIT('h8)
	) name21606 (
		\wishbone_rx_fifo_fifo_reg[13][13]/P0001 ,
		_w31986_,
		_w32118_
	);
	LUT2 #(
		.INIT('h8)
	) name21607 (
		\wishbone_rx_fifo_fifo_reg[2][13]/P0001 ,
		_w31978_,
		_w32119_
	);
	LUT2 #(
		.INIT('h8)
	) name21608 (
		\wishbone_rx_fifo_fifo_reg[12][13]/P0001 ,
		_w31984_,
		_w32120_
	);
	LUT2 #(
		.INIT('h8)
	) name21609 (
		\wishbone_rx_fifo_fifo_reg[15][13]/P0001 ,
		_w31969_,
		_w32121_
	);
	LUT2 #(
		.INIT('h8)
	) name21610 (
		\wishbone_rx_fifo_fifo_reg[11][13]/P0001 ,
		_w31988_,
		_w32122_
	);
	LUT2 #(
		.INIT('h8)
	) name21611 (
		\wishbone_rx_fifo_fifo_reg[6][13]/P0001 ,
		_w31958_,
		_w32123_
	);
	LUT2 #(
		.INIT('h1)
	) name21612 (
		_w32109_,
		_w32110_,
		_w32124_
	);
	LUT2 #(
		.INIT('h1)
	) name21613 (
		_w32111_,
		_w32112_,
		_w32125_
	);
	LUT2 #(
		.INIT('h1)
	) name21614 (
		_w32113_,
		_w32114_,
		_w32126_
	);
	LUT2 #(
		.INIT('h1)
	) name21615 (
		_w32115_,
		_w32116_,
		_w32127_
	);
	LUT2 #(
		.INIT('h1)
	) name21616 (
		_w32117_,
		_w32118_,
		_w32128_
	);
	LUT2 #(
		.INIT('h1)
	) name21617 (
		_w32119_,
		_w32120_,
		_w32129_
	);
	LUT2 #(
		.INIT('h1)
	) name21618 (
		_w32121_,
		_w32122_,
		_w32130_
	);
	LUT2 #(
		.INIT('h4)
	) name21619 (
		_w32123_,
		_w32130_,
		_w32131_
	);
	LUT2 #(
		.INIT('h8)
	) name21620 (
		_w32128_,
		_w32129_,
		_w32132_
	);
	LUT2 #(
		.INIT('h8)
	) name21621 (
		_w32126_,
		_w32127_,
		_w32133_
	);
	LUT2 #(
		.INIT('h8)
	) name21622 (
		_w32124_,
		_w32125_,
		_w32134_
	);
	LUT2 #(
		.INIT('h8)
	) name21623 (
		_w32133_,
		_w32134_,
		_w32135_
	);
	LUT2 #(
		.INIT('h8)
	) name21624 (
		_w32131_,
		_w32132_,
		_w32136_
	);
	LUT2 #(
		.INIT('h8)
	) name21625 (
		_w32135_,
		_w32136_,
		_w32137_
	);
	LUT2 #(
		.INIT('h1)
	) name21626 (
		_w31950_,
		_w32137_,
		_w32138_
	);
	LUT2 #(
		.INIT('h1)
	) name21627 (
		_w32108_,
		_w32138_,
		_w32139_
	);
	LUT2 #(
		.INIT('h8)
	) name21628 (
		\wishbone_rx_fifo_fifo_reg[12][14]/P0001 ,
		_w31984_,
		_w32140_
	);
	LUT2 #(
		.INIT('h8)
	) name21629 (
		\wishbone_rx_fifo_fifo_reg[5][14]/P0001 ,
		_w31980_,
		_w32141_
	);
	LUT2 #(
		.INIT('h8)
	) name21630 (
		\wishbone_rx_fifo_fifo_reg[2][14]/P0001 ,
		_w31978_,
		_w32142_
	);
	LUT2 #(
		.INIT('h8)
	) name21631 (
		\wishbone_rx_fifo_fifo_reg[11][14]/P0001 ,
		_w31988_,
		_w32143_
	);
	LUT2 #(
		.INIT('h8)
	) name21632 (
		\wishbone_rx_fifo_fifo_reg[3][14]/P0001 ,
		_w31990_,
		_w32144_
	);
	LUT2 #(
		.INIT('h8)
	) name21633 (
		\wishbone_rx_fifo_fifo_reg[6][14]/P0001 ,
		_w31958_,
		_w32145_
	);
	LUT2 #(
		.INIT('h8)
	) name21634 (
		\wishbone_rx_fifo_fifo_reg[8][14]/P0001 ,
		_w31974_,
		_w32146_
	);
	LUT2 #(
		.INIT('h8)
	) name21635 (
		\wishbone_rx_fifo_fifo_reg[15][14]/P0001 ,
		_w31969_,
		_w32147_
	);
	LUT2 #(
		.INIT('h8)
	) name21636 (
		\wishbone_rx_fifo_fifo_reg[13][14]/P0001 ,
		_w31986_,
		_w32148_
	);
	LUT2 #(
		.INIT('h8)
	) name21637 (
		\wishbone_rx_fifo_fifo_reg[7][14]/P0001 ,
		_w31964_,
		_w32149_
	);
	LUT2 #(
		.INIT('h8)
	) name21638 (
		\wishbone_rx_fifo_fifo_reg[14][14]/P0001 ,
		_w31982_,
		_w32150_
	);
	LUT2 #(
		.INIT('h8)
	) name21639 (
		\wishbone_rx_fifo_fifo_reg[1][14]/P0001 ,
		_w31976_,
		_w32151_
	);
	LUT2 #(
		.INIT('h8)
	) name21640 (
		\wishbone_rx_fifo_fifo_reg[10][14]/P0001 ,
		_w31961_,
		_w32152_
	);
	LUT2 #(
		.INIT('h8)
	) name21641 (
		\wishbone_rx_fifo_fifo_reg[9][14]/P0001 ,
		_w31972_,
		_w32153_
	);
	LUT2 #(
		.INIT('h8)
	) name21642 (
		\wishbone_rx_fifo_fifo_reg[4][14]/P0001 ,
		_w31966_,
		_w32154_
	);
	LUT2 #(
		.INIT('h1)
	) name21643 (
		_w31950_,
		_w32140_,
		_w32155_
	);
	LUT2 #(
		.INIT('h1)
	) name21644 (
		_w32141_,
		_w32142_,
		_w32156_
	);
	LUT2 #(
		.INIT('h1)
	) name21645 (
		_w32143_,
		_w32144_,
		_w32157_
	);
	LUT2 #(
		.INIT('h1)
	) name21646 (
		_w32145_,
		_w32146_,
		_w32158_
	);
	LUT2 #(
		.INIT('h1)
	) name21647 (
		_w32147_,
		_w32148_,
		_w32159_
	);
	LUT2 #(
		.INIT('h1)
	) name21648 (
		_w32149_,
		_w32150_,
		_w32160_
	);
	LUT2 #(
		.INIT('h1)
	) name21649 (
		_w32151_,
		_w32152_,
		_w32161_
	);
	LUT2 #(
		.INIT('h1)
	) name21650 (
		_w32153_,
		_w32154_,
		_w32162_
	);
	LUT2 #(
		.INIT('h8)
	) name21651 (
		_w32161_,
		_w32162_,
		_w32163_
	);
	LUT2 #(
		.INIT('h8)
	) name21652 (
		_w32159_,
		_w32160_,
		_w32164_
	);
	LUT2 #(
		.INIT('h8)
	) name21653 (
		_w32157_,
		_w32158_,
		_w32165_
	);
	LUT2 #(
		.INIT('h8)
	) name21654 (
		_w32155_,
		_w32156_,
		_w32166_
	);
	LUT2 #(
		.INIT('h8)
	) name21655 (
		_w32165_,
		_w32166_,
		_w32167_
	);
	LUT2 #(
		.INIT('h8)
	) name21656 (
		_w32163_,
		_w32164_,
		_w32168_
	);
	LUT2 #(
		.INIT('h8)
	) name21657 (
		_w32167_,
		_w32168_,
		_w32169_
	);
	LUT2 #(
		.INIT('h4)
	) name21658 (
		\wishbone_rx_fifo_fifo_reg[0][14]/P0001 ,
		_w31950_,
		_w32170_
	);
	LUT2 #(
		.INIT('h1)
	) name21659 (
		_w32169_,
		_w32170_,
		_w32171_
	);
	LUT2 #(
		.INIT('h8)
	) name21660 (
		\wishbone_rx_fifo_fifo_reg[0][14]/P0001 ,
		_w31953_,
		_w32172_
	);
	LUT2 #(
		.INIT('h1)
	) name21661 (
		_w32171_,
		_w32172_,
		_w32173_
	);
	LUT2 #(
		.INIT('h2)
	) name21662 (
		\wishbone_rx_fifo_fifo_reg[0][15]/P0001 ,
		_w31954_,
		_w32174_
	);
	LUT2 #(
		.INIT('h8)
	) name21663 (
		\wishbone_rx_fifo_fifo_reg[12][15]/P0001 ,
		_w31984_,
		_w32175_
	);
	LUT2 #(
		.INIT('h8)
	) name21664 (
		\wishbone_rx_fifo_fifo_reg[5][15]/P0001 ,
		_w31980_,
		_w32176_
	);
	LUT2 #(
		.INIT('h8)
	) name21665 (
		\wishbone_rx_fifo_fifo_reg[4][15]/P0001 ,
		_w31966_,
		_w32177_
	);
	LUT2 #(
		.INIT('h8)
	) name21666 (
		\wishbone_rx_fifo_fifo_reg[8][15]/P0001 ,
		_w31974_,
		_w32178_
	);
	LUT2 #(
		.INIT('h8)
	) name21667 (
		\wishbone_rx_fifo_fifo_reg[14][15]/P0001 ,
		_w31982_,
		_w32179_
	);
	LUT2 #(
		.INIT('h8)
	) name21668 (
		\wishbone_rx_fifo_fifo_reg[6][15]/P0001 ,
		_w31958_,
		_w32180_
	);
	LUT2 #(
		.INIT('h8)
	) name21669 (
		\wishbone_rx_fifo_fifo_reg[1][15]/P0001 ,
		_w31976_,
		_w32181_
	);
	LUT2 #(
		.INIT('h8)
	) name21670 (
		\wishbone_rx_fifo_fifo_reg[10][15]/P0001 ,
		_w31961_,
		_w32182_
	);
	LUT2 #(
		.INIT('h8)
	) name21671 (
		\wishbone_rx_fifo_fifo_reg[7][15]/P0001 ,
		_w31964_,
		_w32183_
	);
	LUT2 #(
		.INIT('h8)
	) name21672 (
		\wishbone_rx_fifo_fifo_reg[2][15]/P0001 ,
		_w31978_,
		_w32184_
	);
	LUT2 #(
		.INIT('h8)
	) name21673 (
		\wishbone_rx_fifo_fifo_reg[13][15]/P0001 ,
		_w31986_,
		_w32185_
	);
	LUT2 #(
		.INIT('h8)
	) name21674 (
		\wishbone_rx_fifo_fifo_reg[9][15]/P0001 ,
		_w31972_,
		_w32186_
	);
	LUT2 #(
		.INIT('h8)
	) name21675 (
		\wishbone_rx_fifo_fifo_reg[15][15]/P0001 ,
		_w31969_,
		_w32187_
	);
	LUT2 #(
		.INIT('h8)
	) name21676 (
		\wishbone_rx_fifo_fifo_reg[3][15]/P0001 ,
		_w31990_,
		_w32188_
	);
	LUT2 #(
		.INIT('h8)
	) name21677 (
		\wishbone_rx_fifo_fifo_reg[11][15]/P0001 ,
		_w31988_,
		_w32189_
	);
	LUT2 #(
		.INIT('h1)
	) name21678 (
		_w32175_,
		_w32176_,
		_w32190_
	);
	LUT2 #(
		.INIT('h1)
	) name21679 (
		_w32177_,
		_w32178_,
		_w32191_
	);
	LUT2 #(
		.INIT('h1)
	) name21680 (
		_w32179_,
		_w32180_,
		_w32192_
	);
	LUT2 #(
		.INIT('h1)
	) name21681 (
		_w32181_,
		_w32182_,
		_w32193_
	);
	LUT2 #(
		.INIT('h1)
	) name21682 (
		_w32183_,
		_w32184_,
		_w32194_
	);
	LUT2 #(
		.INIT('h1)
	) name21683 (
		_w32185_,
		_w32186_,
		_w32195_
	);
	LUT2 #(
		.INIT('h1)
	) name21684 (
		_w32187_,
		_w32188_,
		_w32196_
	);
	LUT2 #(
		.INIT('h4)
	) name21685 (
		_w32189_,
		_w32196_,
		_w32197_
	);
	LUT2 #(
		.INIT('h8)
	) name21686 (
		_w32194_,
		_w32195_,
		_w32198_
	);
	LUT2 #(
		.INIT('h8)
	) name21687 (
		_w32192_,
		_w32193_,
		_w32199_
	);
	LUT2 #(
		.INIT('h8)
	) name21688 (
		_w32190_,
		_w32191_,
		_w32200_
	);
	LUT2 #(
		.INIT('h8)
	) name21689 (
		_w32199_,
		_w32200_,
		_w32201_
	);
	LUT2 #(
		.INIT('h8)
	) name21690 (
		_w32197_,
		_w32198_,
		_w32202_
	);
	LUT2 #(
		.INIT('h8)
	) name21691 (
		_w32201_,
		_w32202_,
		_w32203_
	);
	LUT2 #(
		.INIT('h1)
	) name21692 (
		_w31950_,
		_w32203_,
		_w32204_
	);
	LUT2 #(
		.INIT('h1)
	) name21693 (
		_w32174_,
		_w32204_,
		_w32205_
	);
	LUT2 #(
		.INIT('h8)
	) name21694 (
		\wishbone_rx_fifo_fifo_reg[12][16]/P0001 ,
		_w31984_,
		_w32206_
	);
	LUT2 #(
		.INIT('h8)
	) name21695 (
		\wishbone_rx_fifo_fifo_reg[3][16]/P0001 ,
		_w31990_,
		_w32207_
	);
	LUT2 #(
		.INIT('h8)
	) name21696 (
		\wishbone_rx_fifo_fifo_reg[1][16]/P0001 ,
		_w31976_,
		_w32208_
	);
	LUT2 #(
		.INIT('h8)
	) name21697 (
		\wishbone_rx_fifo_fifo_reg[11][16]/P0001 ,
		_w31988_,
		_w32209_
	);
	LUT2 #(
		.INIT('h8)
	) name21698 (
		\wishbone_rx_fifo_fifo_reg[9][16]/P0001 ,
		_w31972_,
		_w32210_
	);
	LUT2 #(
		.INIT('h8)
	) name21699 (
		\wishbone_rx_fifo_fifo_reg[6][16]/P0001 ,
		_w31958_,
		_w32211_
	);
	LUT2 #(
		.INIT('h8)
	) name21700 (
		\wishbone_rx_fifo_fifo_reg[15][16]/P0001 ,
		_w31969_,
		_w32212_
	);
	LUT2 #(
		.INIT('h8)
	) name21701 (
		\wishbone_rx_fifo_fifo_reg[7][16]/P0001 ,
		_w31964_,
		_w32213_
	);
	LUT2 #(
		.INIT('h8)
	) name21702 (
		\wishbone_rx_fifo_fifo_reg[8][16]/P0001 ,
		_w31974_,
		_w32214_
	);
	LUT2 #(
		.INIT('h8)
	) name21703 (
		\wishbone_rx_fifo_fifo_reg[13][16]/P0001 ,
		_w31986_,
		_w32215_
	);
	LUT2 #(
		.INIT('h8)
	) name21704 (
		\wishbone_rx_fifo_fifo_reg[14][16]/P0001 ,
		_w31982_,
		_w32216_
	);
	LUT2 #(
		.INIT('h8)
	) name21705 (
		\wishbone_rx_fifo_fifo_reg[5][16]/P0001 ,
		_w31980_,
		_w32217_
	);
	LUT2 #(
		.INIT('h8)
	) name21706 (
		\wishbone_rx_fifo_fifo_reg[10][16]/P0001 ,
		_w31961_,
		_w32218_
	);
	LUT2 #(
		.INIT('h8)
	) name21707 (
		\wishbone_rx_fifo_fifo_reg[2][16]/P0001 ,
		_w31978_,
		_w32219_
	);
	LUT2 #(
		.INIT('h8)
	) name21708 (
		\wishbone_rx_fifo_fifo_reg[4][16]/P0001 ,
		_w31966_,
		_w32220_
	);
	LUT2 #(
		.INIT('h1)
	) name21709 (
		_w31950_,
		_w32206_,
		_w32221_
	);
	LUT2 #(
		.INIT('h1)
	) name21710 (
		_w32207_,
		_w32208_,
		_w32222_
	);
	LUT2 #(
		.INIT('h1)
	) name21711 (
		_w32209_,
		_w32210_,
		_w32223_
	);
	LUT2 #(
		.INIT('h1)
	) name21712 (
		_w32211_,
		_w32212_,
		_w32224_
	);
	LUT2 #(
		.INIT('h1)
	) name21713 (
		_w32213_,
		_w32214_,
		_w32225_
	);
	LUT2 #(
		.INIT('h1)
	) name21714 (
		_w32215_,
		_w32216_,
		_w32226_
	);
	LUT2 #(
		.INIT('h1)
	) name21715 (
		_w32217_,
		_w32218_,
		_w32227_
	);
	LUT2 #(
		.INIT('h1)
	) name21716 (
		_w32219_,
		_w32220_,
		_w32228_
	);
	LUT2 #(
		.INIT('h8)
	) name21717 (
		_w32227_,
		_w32228_,
		_w32229_
	);
	LUT2 #(
		.INIT('h8)
	) name21718 (
		_w32225_,
		_w32226_,
		_w32230_
	);
	LUT2 #(
		.INIT('h8)
	) name21719 (
		_w32223_,
		_w32224_,
		_w32231_
	);
	LUT2 #(
		.INIT('h8)
	) name21720 (
		_w32221_,
		_w32222_,
		_w32232_
	);
	LUT2 #(
		.INIT('h8)
	) name21721 (
		_w32231_,
		_w32232_,
		_w32233_
	);
	LUT2 #(
		.INIT('h8)
	) name21722 (
		_w32229_,
		_w32230_,
		_w32234_
	);
	LUT2 #(
		.INIT('h8)
	) name21723 (
		_w32233_,
		_w32234_,
		_w32235_
	);
	LUT2 #(
		.INIT('h4)
	) name21724 (
		\wishbone_rx_fifo_fifo_reg[0][16]/P0001 ,
		_w31950_,
		_w32236_
	);
	LUT2 #(
		.INIT('h1)
	) name21725 (
		_w32235_,
		_w32236_,
		_w32237_
	);
	LUT2 #(
		.INIT('h8)
	) name21726 (
		\wishbone_rx_fifo_fifo_reg[0][16]/P0001 ,
		_w31953_,
		_w32238_
	);
	LUT2 #(
		.INIT('h1)
	) name21727 (
		_w32237_,
		_w32238_,
		_w32239_
	);
	LUT2 #(
		.INIT('h2)
	) name21728 (
		\wishbone_rx_fifo_fifo_reg[0][17]/P0001 ,
		_w31954_,
		_w32240_
	);
	LUT2 #(
		.INIT('h8)
	) name21729 (
		\wishbone_rx_fifo_fifo_reg[12][17]/P0001 ,
		_w31984_,
		_w32241_
	);
	LUT2 #(
		.INIT('h8)
	) name21730 (
		\wishbone_rx_fifo_fifo_reg[5][17]/P0001 ,
		_w31980_,
		_w32242_
	);
	LUT2 #(
		.INIT('h8)
	) name21731 (
		\wishbone_rx_fifo_fifo_reg[4][17]/P0001 ,
		_w31966_,
		_w32243_
	);
	LUT2 #(
		.INIT('h8)
	) name21732 (
		\wishbone_rx_fifo_fifo_reg[8][17]/P0001 ,
		_w31974_,
		_w32244_
	);
	LUT2 #(
		.INIT('h8)
	) name21733 (
		\wishbone_rx_fifo_fifo_reg[14][17]/P0001 ,
		_w31982_,
		_w32245_
	);
	LUT2 #(
		.INIT('h8)
	) name21734 (
		\wishbone_rx_fifo_fifo_reg[9][17]/P0001 ,
		_w31972_,
		_w32246_
	);
	LUT2 #(
		.INIT('h8)
	) name21735 (
		\wishbone_rx_fifo_fifo_reg[1][17]/P0001 ,
		_w31976_,
		_w32247_
	);
	LUT2 #(
		.INIT('h8)
	) name21736 (
		\wishbone_rx_fifo_fifo_reg[10][17]/P0001 ,
		_w31961_,
		_w32248_
	);
	LUT2 #(
		.INIT('h8)
	) name21737 (
		\wishbone_rx_fifo_fifo_reg[7][17]/P0001 ,
		_w31964_,
		_w32249_
	);
	LUT2 #(
		.INIT('h8)
	) name21738 (
		\wishbone_rx_fifo_fifo_reg[2][17]/P0001 ,
		_w31978_,
		_w32250_
	);
	LUT2 #(
		.INIT('h8)
	) name21739 (
		\wishbone_rx_fifo_fifo_reg[13][17]/P0001 ,
		_w31986_,
		_w32251_
	);
	LUT2 #(
		.INIT('h8)
	) name21740 (
		\wishbone_rx_fifo_fifo_reg[6][17]/P0001 ,
		_w31958_,
		_w32252_
	);
	LUT2 #(
		.INIT('h8)
	) name21741 (
		\wishbone_rx_fifo_fifo_reg[15][17]/P0001 ,
		_w31969_,
		_w32253_
	);
	LUT2 #(
		.INIT('h8)
	) name21742 (
		\wishbone_rx_fifo_fifo_reg[3][17]/P0001 ,
		_w31990_,
		_w32254_
	);
	LUT2 #(
		.INIT('h8)
	) name21743 (
		\wishbone_rx_fifo_fifo_reg[11][17]/P0001 ,
		_w31988_,
		_w32255_
	);
	LUT2 #(
		.INIT('h1)
	) name21744 (
		_w32241_,
		_w32242_,
		_w32256_
	);
	LUT2 #(
		.INIT('h1)
	) name21745 (
		_w32243_,
		_w32244_,
		_w32257_
	);
	LUT2 #(
		.INIT('h1)
	) name21746 (
		_w32245_,
		_w32246_,
		_w32258_
	);
	LUT2 #(
		.INIT('h1)
	) name21747 (
		_w32247_,
		_w32248_,
		_w32259_
	);
	LUT2 #(
		.INIT('h1)
	) name21748 (
		_w32249_,
		_w32250_,
		_w32260_
	);
	LUT2 #(
		.INIT('h1)
	) name21749 (
		_w32251_,
		_w32252_,
		_w32261_
	);
	LUT2 #(
		.INIT('h1)
	) name21750 (
		_w32253_,
		_w32254_,
		_w32262_
	);
	LUT2 #(
		.INIT('h4)
	) name21751 (
		_w32255_,
		_w32262_,
		_w32263_
	);
	LUT2 #(
		.INIT('h8)
	) name21752 (
		_w32260_,
		_w32261_,
		_w32264_
	);
	LUT2 #(
		.INIT('h8)
	) name21753 (
		_w32258_,
		_w32259_,
		_w32265_
	);
	LUT2 #(
		.INIT('h8)
	) name21754 (
		_w32256_,
		_w32257_,
		_w32266_
	);
	LUT2 #(
		.INIT('h8)
	) name21755 (
		_w32265_,
		_w32266_,
		_w32267_
	);
	LUT2 #(
		.INIT('h8)
	) name21756 (
		_w32263_,
		_w32264_,
		_w32268_
	);
	LUT2 #(
		.INIT('h8)
	) name21757 (
		_w32267_,
		_w32268_,
		_w32269_
	);
	LUT2 #(
		.INIT('h1)
	) name21758 (
		_w31950_,
		_w32269_,
		_w32270_
	);
	LUT2 #(
		.INIT('h1)
	) name21759 (
		_w32240_,
		_w32270_,
		_w32271_
	);
	LUT2 #(
		.INIT('h2)
	) name21760 (
		\wishbone_rx_fifo_fifo_reg[0][18]/P0001 ,
		_w31954_,
		_w32272_
	);
	LUT2 #(
		.INIT('h8)
	) name21761 (
		\wishbone_rx_fifo_fifo_reg[3][18]/P0001 ,
		_w31990_,
		_w32273_
	);
	LUT2 #(
		.INIT('h8)
	) name21762 (
		\wishbone_rx_fifo_fifo_reg[9][18]/P0001 ,
		_w31972_,
		_w32274_
	);
	LUT2 #(
		.INIT('h8)
	) name21763 (
		\wishbone_rx_fifo_fifo_reg[5][18]/P0001 ,
		_w31980_,
		_w32275_
	);
	LUT2 #(
		.INIT('h8)
	) name21764 (
		\wishbone_rx_fifo_fifo_reg[7][18]/P0001 ,
		_w31964_,
		_w32276_
	);
	LUT2 #(
		.INIT('h8)
	) name21765 (
		\wishbone_rx_fifo_fifo_reg[10][18]/P0001 ,
		_w31961_,
		_w32277_
	);
	LUT2 #(
		.INIT('h8)
	) name21766 (
		\wishbone_rx_fifo_fifo_reg[6][18]/P0001 ,
		_w31958_,
		_w32278_
	);
	LUT2 #(
		.INIT('h8)
	) name21767 (
		\wishbone_rx_fifo_fifo_reg[12][18]/P0001 ,
		_w31984_,
		_w32279_
	);
	LUT2 #(
		.INIT('h8)
	) name21768 (
		\wishbone_rx_fifo_fifo_reg[4][18]/P0001 ,
		_w31966_,
		_w32280_
	);
	LUT2 #(
		.INIT('h8)
	) name21769 (
		\wishbone_rx_fifo_fifo_reg[1][18]/P0001 ,
		_w31976_,
		_w32281_
	);
	LUT2 #(
		.INIT('h8)
	) name21770 (
		\wishbone_rx_fifo_fifo_reg[13][18]/P0001 ,
		_w31986_,
		_w32282_
	);
	LUT2 #(
		.INIT('h8)
	) name21771 (
		\wishbone_rx_fifo_fifo_reg[2][18]/P0001 ,
		_w31978_,
		_w32283_
	);
	LUT2 #(
		.INIT('h8)
	) name21772 (
		\wishbone_rx_fifo_fifo_reg[14][18]/P0001 ,
		_w31982_,
		_w32284_
	);
	LUT2 #(
		.INIT('h8)
	) name21773 (
		\wishbone_rx_fifo_fifo_reg[8][18]/P0001 ,
		_w31974_,
		_w32285_
	);
	LUT2 #(
		.INIT('h8)
	) name21774 (
		\wishbone_rx_fifo_fifo_reg[11][18]/P0001 ,
		_w31988_,
		_w32286_
	);
	LUT2 #(
		.INIT('h8)
	) name21775 (
		\wishbone_rx_fifo_fifo_reg[15][18]/P0001 ,
		_w31969_,
		_w32287_
	);
	LUT2 #(
		.INIT('h1)
	) name21776 (
		_w32273_,
		_w32274_,
		_w32288_
	);
	LUT2 #(
		.INIT('h1)
	) name21777 (
		_w32275_,
		_w32276_,
		_w32289_
	);
	LUT2 #(
		.INIT('h1)
	) name21778 (
		_w32277_,
		_w32278_,
		_w32290_
	);
	LUT2 #(
		.INIT('h1)
	) name21779 (
		_w32279_,
		_w32280_,
		_w32291_
	);
	LUT2 #(
		.INIT('h1)
	) name21780 (
		_w32281_,
		_w32282_,
		_w32292_
	);
	LUT2 #(
		.INIT('h1)
	) name21781 (
		_w32283_,
		_w32284_,
		_w32293_
	);
	LUT2 #(
		.INIT('h1)
	) name21782 (
		_w32285_,
		_w32286_,
		_w32294_
	);
	LUT2 #(
		.INIT('h4)
	) name21783 (
		_w32287_,
		_w32294_,
		_w32295_
	);
	LUT2 #(
		.INIT('h8)
	) name21784 (
		_w32292_,
		_w32293_,
		_w32296_
	);
	LUT2 #(
		.INIT('h8)
	) name21785 (
		_w32290_,
		_w32291_,
		_w32297_
	);
	LUT2 #(
		.INIT('h8)
	) name21786 (
		_w32288_,
		_w32289_,
		_w32298_
	);
	LUT2 #(
		.INIT('h8)
	) name21787 (
		_w32297_,
		_w32298_,
		_w32299_
	);
	LUT2 #(
		.INIT('h8)
	) name21788 (
		_w32295_,
		_w32296_,
		_w32300_
	);
	LUT2 #(
		.INIT('h8)
	) name21789 (
		_w32299_,
		_w32300_,
		_w32301_
	);
	LUT2 #(
		.INIT('h1)
	) name21790 (
		_w31950_,
		_w32301_,
		_w32302_
	);
	LUT2 #(
		.INIT('h1)
	) name21791 (
		_w32272_,
		_w32302_,
		_w32303_
	);
	LUT2 #(
		.INIT('h2)
	) name21792 (
		\wishbone_rx_fifo_fifo_reg[0][19]/P0001 ,
		_w31954_,
		_w32304_
	);
	LUT2 #(
		.INIT('h8)
	) name21793 (
		\wishbone_rx_fifo_fifo_reg[9][19]/P0001 ,
		_w31972_,
		_w32305_
	);
	LUT2 #(
		.INIT('h8)
	) name21794 (
		\wishbone_rx_fifo_fifo_reg[8][19]/P0001 ,
		_w31974_,
		_w32306_
	);
	LUT2 #(
		.INIT('h8)
	) name21795 (
		\wishbone_rx_fifo_fifo_reg[12][19]/P0001 ,
		_w31984_,
		_w32307_
	);
	LUT2 #(
		.INIT('h8)
	) name21796 (
		\wishbone_rx_fifo_fifo_reg[13][19]/P0001 ,
		_w31986_,
		_w32308_
	);
	LUT2 #(
		.INIT('h8)
	) name21797 (
		\wishbone_rx_fifo_fifo_reg[2][19]/P0001 ,
		_w31978_,
		_w32309_
	);
	LUT2 #(
		.INIT('h8)
	) name21798 (
		\wishbone_rx_fifo_fifo_reg[3][19]/P0001 ,
		_w31990_,
		_w32310_
	);
	LUT2 #(
		.INIT('h8)
	) name21799 (
		\wishbone_rx_fifo_fifo_reg[4][19]/P0001 ,
		_w31966_,
		_w32311_
	);
	LUT2 #(
		.INIT('h8)
	) name21800 (
		\wishbone_rx_fifo_fifo_reg[5][19]/P0001 ,
		_w31980_,
		_w32312_
	);
	LUT2 #(
		.INIT('h8)
	) name21801 (
		\wishbone_rx_fifo_fifo_reg[10][19]/P0001 ,
		_w31961_,
		_w32313_
	);
	LUT2 #(
		.INIT('h8)
	) name21802 (
		\wishbone_rx_fifo_fifo_reg[7][19]/P0001 ,
		_w31964_,
		_w32314_
	);
	LUT2 #(
		.INIT('h8)
	) name21803 (
		\wishbone_rx_fifo_fifo_reg[1][19]/P0001 ,
		_w31976_,
		_w32315_
	);
	LUT2 #(
		.INIT('h8)
	) name21804 (
		\wishbone_rx_fifo_fifo_reg[11][19]/P0001 ,
		_w31988_,
		_w32316_
	);
	LUT2 #(
		.INIT('h8)
	) name21805 (
		\wishbone_rx_fifo_fifo_reg[6][19]/P0001 ,
		_w31958_,
		_w32317_
	);
	LUT2 #(
		.INIT('h8)
	) name21806 (
		\wishbone_rx_fifo_fifo_reg[15][19]/P0001 ,
		_w31969_,
		_w32318_
	);
	LUT2 #(
		.INIT('h8)
	) name21807 (
		\wishbone_rx_fifo_fifo_reg[14][19]/P0001 ,
		_w31982_,
		_w32319_
	);
	LUT2 #(
		.INIT('h1)
	) name21808 (
		_w32305_,
		_w32306_,
		_w32320_
	);
	LUT2 #(
		.INIT('h1)
	) name21809 (
		_w32307_,
		_w32308_,
		_w32321_
	);
	LUT2 #(
		.INIT('h1)
	) name21810 (
		_w32309_,
		_w32310_,
		_w32322_
	);
	LUT2 #(
		.INIT('h1)
	) name21811 (
		_w32311_,
		_w32312_,
		_w32323_
	);
	LUT2 #(
		.INIT('h1)
	) name21812 (
		_w32313_,
		_w32314_,
		_w32324_
	);
	LUT2 #(
		.INIT('h1)
	) name21813 (
		_w32315_,
		_w32316_,
		_w32325_
	);
	LUT2 #(
		.INIT('h1)
	) name21814 (
		_w32317_,
		_w32318_,
		_w32326_
	);
	LUT2 #(
		.INIT('h4)
	) name21815 (
		_w32319_,
		_w32326_,
		_w32327_
	);
	LUT2 #(
		.INIT('h8)
	) name21816 (
		_w32324_,
		_w32325_,
		_w32328_
	);
	LUT2 #(
		.INIT('h8)
	) name21817 (
		_w32322_,
		_w32323_,
		_w32329_
	);
	LUT2 #(
		.INIT('h8)
	) name21818 (
		_w32320_,
		_w32321_,
		_w32330_
	);
	LUT2 #(
		.INIT('h8)
	) name21819 (
		_w32329_,
		_w32330_,
		_w32331_
	);
	LUT2 #(
		.INIT('h8)
	) name21820 (
		_w32327_,
		_w32328_,
		_w32332_
	);
	LUT2 #(
		.INIT('h8)
	) name21821 (
		_w32331_,
		_w32332_,
		_w32333_
	);
	LUT2 #(
		.INIT('h1)
	) name21822 (
		_w31950_,
		_w32333_,
		_w32334_
	);
	LUT2 #(
		.INIT('h1)
	) name21823 (
		_w32304_,
		_w32334_,
		_w32335_
	);
	LUT2 #(
		.INIT('h8)
	) name21824 (
		\wishbone_rx_fifo_fifo_reg[5][1]/P0001 ,
		_w31980_,
		_w32336_
	);
	LUT2 #(
		.INIT('h8)
	) name21825 (
		\wishbone_rx_fifo_fifo_reg[3][1]/P0001 ,
		_w31990_,
		_w32337_
	);
	LUT2 #(
		.INIT('h8)
	) name21826 (
		\wishbone_rx_fifo_fifo_reg[1][1]/P0001 ,
		_w31976_,
		_w32338_
	);
	LUT2 #(
		.INIT('h8)
	) name21827 (
		\wishbone_rx_fifo_fifo_reg[11][1]/P0001 ,
		_w31988_,
		_w32339_
	);
	LUT2 #(
		.INIT('h8)
	) name21828 (
		\wishbone_rx_fifo_fifo_reg[9][1]/P0001 ,
		_w31972_,
		_w32340_
	);
	LUT2 #(
		.INIT('h8)
	) name21829 (
		\wishbone_rx_fifo_fifo_reg[6][1]/P0001 ,
		_w31958_,
		_w32341_
	);
	LUT2 #(
		.INIT('h8)
	) name21830 (
		\wishbone_rx_fifo_fifo_reg[15][1]/P0001 ,
		_w31969_,
		_w32342_
	);
	LUT2 #(
		.INIT('h8)
	) name21831 (
		\wishbone_rx_fifo_fifo_reg[7][1]/P0001 ,
		_w31964_,
		_w32343_
	);
	LUT2 #(
		.INIT('h8)
	) name21832 (
		\wishbone_rx_fifo_fifo_reg[8][1]/P0001 ,
		_w31974_,
		_w32344_
	);
	LUT2 #(
		.INIT('h8)
	) name21833 (
		\wishbone_rx_fifo_fifo_reg[13][1]/P0001 ,
		_w31986_,
		_w32345_
	);
	LUT2 #(
		.INIT('h8)
	) name21834 (
		\wishbone_rx_fifo_fifo_reg[12][1]/P0001 ,
		_w31984_,
		_w32346_
	);
	LUT2 #(
		.INIT('h8)
	) name21835 (
		\wishbone_rx_fifo_fifo_reg[14][1]/P0001 ,
		_w31982_,
		_w32347_
	);
	LUT2 #(
		.INIT('h8)
	) name21836 (
		\wishbone_rx_fifo_fifo_reg[10][1]/P0001 ,
		_w31961_,
		_w32348_
	);
	LUT2 #(
		.INIT('h8)
	) name21837 (
		\wishbone_rx_fifo_fifo_reg[2][1]/P0001 ,
		_w31978_,
		_w32349_
	);
	LUT2 #(
		.INIT('h8)
	) name21838 (
		\wishbone_rx_fifo_fifo_reg[4][1]/P0001 ,
		_w31966_,
		_w32350_
	);
	LUT2 #(
		.INIT('h1)
	) name21839 (
		_w31950_,
		_w32336_,
		_w32351_
	);
	LUT2 #(
		.INIT('h1)
	) name21840 (
		_w32337_,
		_w32338_,
		_w32352_
	);
	LUT2 #(
		.INIT('h1)
	) name21841 (
		_w32339_,
		_w32340_,
		_w32353_
	);
	LUT2 #(
		.INIT('h1)
	) name21842 (
		_w32341_,
		_w32342_,
		_w32354_
	);
	LUT2 #(
		.INIT('h1)
	) name21843 (
		_w32343_,
		_w32344_,
		_w32355_
	);
	LUT2 #(
		.INIT('h1)
	) name21844 (
		_w32345_,
		_w32346_,
		_w32356_
	);
	LUT2 #(
		.INIT('h1)
	) name21845 (
		_w32347_,
		_w32348_,
		_w32357_
	);
	LUT2 #(
		.INIT('h1)
	) name21846 (
		_w32349_,
		_w32350_,
		_w32358_
	);
	LUT2 #(
		.INIT('h8)
	) name21847 (
		_w32357_,
		_w32358_,
		_w32359_
	);
	LUT2 #(
		.INIT('h8)
	) name21848 (
		_w32355_,
		_w32356_,
		_w32360_
	);
	LUT2 #(
		.INIT('h8)
	) name21849 (
		_w32353_,
		_w32354_,
		_w32361_
	);
	LUT2 #(
		.INIT('h8)
	) name21850 (
		_w32351_,
		_w32352_,
		_w32362_
	);
	LUT2 #(
		.INIT('h8)
	) name21851 (
		_w32361_,
		_w32362_,
		_w32363_
	);
	LUT2 #(
		.INIT('h8)
	) name21852 (
		_w32359_,
		_w32360_,
		_w32364_
	);
	LUT2 #(
		.INIT('h8)
	) name21853 (
		_w32363_,
		_w32364_,
		_w32365_
	);
	LUT2 #(
		.INIT('h4)
	) name21854 (
		\wishbone_rx_fifo_fifo_reg[0][1]/P0001 ,
		_w31950_,
		_w32366_
	);
	LUT2 #(
		.INIT('h1)
	) name21855 (
		_w32365_,
		_w32366_,
		_w32367_
	);
	LUT2 #(
		.INIT('h8)
	) name21856 (
		\wishbone_rx_fifo_fifo_reg[0][1]/P0001 ,
		_w31953_,
		_w32368_
	);
	LUT2 #(
		.INIT('h1)
	) name21857 (
		_w32367_,
		_w32368_,
		_w32369_
	);
	LUT2 #(
		.INIT('h8)
	) name21858 (
		\wishbone_rx_fifo_fifo_reg[10][20]/P0001 ,
		_w31961_,
		_w32370_
	);
	LUT2 #(
		.INIT('h8)
	) name21859 (
		\wishbone_rx_fifo_fifo_reg[13][20]/P0001 ,
		_w31986_,
		_w32371_
	);
	LUT2 #(
		.INIT('h8)
	) name21860 (
		\wishbone_rx_fifo_fifo_reg[11][20]/P0001 ,
		_w31988_,
		_w32372_
	);
	LUT2 #(
		.INIT('h8)
	) name21861 (
		\wishbone_rx_fifo_fifo_reg[14][20]/P0001 ,
		_w31982_,
		_w32373_
	);
	LUT2 #(
		.INIT('h8)
	) name21862 (
		\wishbone_rx_fifo_fifo_reg[1][20]/P0001 ,
		_w31976_,
		_w32374_
	);
	LUT2 #(
		.INIT('h8)
	) name21863 (
		\wishbone_rx_fifo_fifo_reg[2][20]/P0001 ,
		_w31978_,
		_w32375_
	);
	LUT2 #(
		.INIT('h8)
	) name21864 (
		\wishbone_rx_fifo_fifo_reg[6][20]/P0001 ,
		_w31958_,
		_w32376_
	);
	LUT2 #(
		.INIT('h8)
	) name21865 (
		\wishbone_rx_fifo_fifo_reg[9][20]/P0001 ,
		_w31972_,
		_w32377_
	);
	LUT2 #(
		.INIT('h8)
	) name21866 (
		\wishbone_rx_fifo_fifo_reg[7][20]/P0001 ,
		_w31964_,
		_w32378_
	);
	LUT2 #(
		.INIT('h8)
	) name21867 (
		\wishbone_rx_fifo_fifo_reg[3][20]/P0001 ,
		_w31990_,
		_w32379_
	);
	LUT2 #(
		.INIT('h8)
	) name21868 (
		\wishbone_rx_fifo_fifo_reg[4][20]/P0001 ,
		_w31966_,
		_w32380_
	);
	LUT2 #(
		.INIT('h8)
	) name21869 (
		\wishbone_rx_fifo_fifo_reg[5][20]/P0001 ,
		_w31980_,
		_w32381_
	);
	LUT2 #(
		.INIT('h8)
	) name21870 (
		\wishbone_rx_fifo_fifo_reg[15][20]/P0001 ,
		_w31969_,
		_w32382_
	);
	LUT2 #(
		.INIT('h8)
	) name21871 (
		\wishbone_rx_fifo_fifo_reg[12][20]/P0001 ,
		_w31984_,
		_w32383_
	);
	LUT2 #(
		.INIT('h8)
	) name21872 (
		\wishbone_rx_fifo_fifo_reg[8][20]/P0001 ,
		_w31974_,
		_w32384_
	);
	LUT2 #(
		.INIT('h1)
	) name21873 (
		_w31950_,
		_w32370_,
		_w32385_
	);
	LUT2 #(
		.INIT('h1)
	) name21874 (
		_w32371_,
		_w32372_,
		_w32386_
	);
	LUT2 #(
		.INIT('h1)
	) name21875 (
		_w32373_,
		_w32374_,
		_w32387_
	);
	LUT2 #(
		.INIT('h1)
	) name21876 (
		_w32375_,
		_w32376_,
		_w32388_
	);
	LUT2 #(
		.INIT('h1)
	) name21877 (
		_w32377_,
		_w32378_,
		_w32389_
	);
	LUT2 #(
		.INIT('h1)
	) name21878 (
		_w32379_,
		_w32380_,
		_w32390_
	);
	LUT2 #(
		.INIT('h1)
	) name21879 (
		_w32381_,
		_w32382_,
		_w32391_
	);
	LUT2 #(
		.INIT('h1)
	) name21880 (
		_w32383_,
		_w32384_,
		_w32392_
	);
	LUT2 #(
		.INIT('h8)
	) name21881 (
		_w32391_,
		_w32392_,
		_w32393_
	);
	LUT2 #(
		.INIT('h8)
	) name21882 (
		_w32389_,
		_w32390_,
		_w32394_
	);
	LUT2 #(
		.INIT('h8)
	) name21883 (
		_w32387_,
		_w32388_,
		_w32395_
	);
	LUT2 #(
		.INIT('h8)
	) name21884 (
		_w32385_,
		_w32386_,
		_w32396_
	);
	LUT2 #(
		.INIT('h8)
	) name21885 (
		_w32395_,
		_w32396_,
		_w32397_
	);
	LUT2 #(
		.INIT('h8)
	) name21886 (
		_w32393_,
		_w32394_,
		_w32398_
	);
	LUT2 #(
		.INIT('h8)
	) name21887 (
		_w32397_,
		_w32398_,
		_w32399_
	);
	LUT2 #(
		.INIT('h4)
	) name21888 (
		\wishbone_rx_fifo_fifo_reg[0][20]/P0001 ,
		_w31950_,
		_w32400_
	);
	LUT2 #(
		.INIT('h1)
	) name21889 (
		_w32399_,
		_w32400_,
		_w32401_
	);
	LUT2 #(
		.INIT('h8)
	) name21890 (
		\wishbone_rx_fifo_fifo_reg[0][20]/P0001 ,
		_w31953_,
		_w32402_
	);
	LUT2 #(
		.INIT('h1)
	) name21891 (
		_w32401_,
		_w32402_,
		_w32403_
	);
	LUT2 #(
		.INIT('h2)
	) name21892 (
		\wishbone_rx_fifo_fifo_reg[0][21]/P0001 ,
		_w31954_,
		_w32404_
	);
	LUT2 #(
		.INIT('h8)
	) name21893 (
		\wishbone_rx_fifo_fifo_reg[6][21]/P0001 ,
		_w31958_,
		_w32405_
	);
	LUT2 #(
		.INIT('h8)
	) name21894 (
		\wishbone_rx_fifo_fifo_reg[12][21]/P0001 ,
		_w31984_,
		_w32406_
	);
	LUT2 #(
		.INIT('h8)
	) name21895 (
		\wishbone_rx_fifo_fifo_reg[9][21]/P0001 ,
		_w31972_,
		_w32407_
	);
	LUT2 #(
		.INIT('h8)
	) name21896 (
		\wishbone_rx_fifo_fifo_reg[11][21]/P0001 ,
		_w31988_,
		_w32408_
	);
	LUT2 #(
		.INIT('h8)
	) name21897 (
		\wishbone_rx_fifo_fifo_reg[7][21]/P0001 ,
		_w31964_,
		_w32409_
	);
	LUT2 #(
		.INIT('h8)
	) name21898 (
		\wishbone_rx_fifo_fifo_reg[5][21]/P0001 ,
		_w31980_,
		_w32410_
	);
	LUT2 #(
		.INIT('h8)
	) name21899 (
		\wishbone_rx_fifo_fifo_reg[2][21]/P0001 ,
		_w31978_,
		_w32411_
	);
	LUT2 #(
		.INIT('h8)
	) name21900 (
		\wishbone_rx_fifo_fifo_reg[13][21]/P0001 ,
		_w31986_,
		_w32412_
	);
	LUT2 #(
		.INIT('h8)
	) name21901 (
		\wishbone_rx_fifo_fifo_reg[4][21]/P0001 ,
		_w31966_,
		_w32413_
	);
	LUT2 #(
		.INIT('h8)
	) name21902 (
		\wishbone_rx_fifo_fifo_reg[15][21]/P0001 ,
		_w31969_,
		_w32414_
	);
	LUT2 #(
		.INIT('h8)
	) name21903 (
		\wishbone_rx_fifo_fifo_reg[8][21]/P0001 ,
		_w31974_,
		_w32415_
	);
	LUT2 #(
		.INIT('h8)
	) name21904 (
		\wishbone_rx_fifo_fifo_reg[14][21]/P0001 ,
		_w31982_,
		_w32416_
	);
	LUT2 #(
		.INIT('h8)
	) name21905 (
		\wishbone_rx_fifo_fifo_reg[10][21]/P0001 ,
		_w31961_,
		_w32417_
	);
	LUT2 #(
		.INIT('h8)
	) name21906 (
		\wishbone_rx_fifo_fifo_reg[1][21]/P0001 ,
		_w31976_,
		_w32418_
	);
	LUT2 #(
		.INIT('h8)
	) name21907 (
		\wishbone_rx_fifo_fifo_reg[3][21]/P0001 ,
		_w31990_,
		_w32419_
	);
	LUT2 #(
		.INIT('h1)
	) name21908 (
		_w32405_,
		_w32406_,
		_w32420_
	);
	LUT2 #(
		.INIT('h1)
	) name21909 (
		_w32407_,
		_w32408_,
		_w32421_
	);
	LUT2 #(
		.INIT('h1)
	) name21910 (
		_w32409_,
		_w32410_,
		_w32422_
	);
	LUT2 #(
		.INIT('h1)
	) name21911 (
		_w32411_,
		_w32412_,
		_w32423_
	);
	LUT2 #(
		.INIT('h1)
	) name21912 (
		_w32413_,
		_w32414_,
		_w32424_
	);
	LUT2 #(
		.INIT('h1)
	) name21913 (
		_w32415_,
		_w32416_,
		_w32425_
	);
	LUT2 #(
		.INIT('h1)
	) name21914 (
		_w32417_,
		_w32418_,
		_w32426_
	);
	LUT2 #(
		.INIT('h4)
	) name21915 (
		_w32419_,
		_w32426_,
		_w32427_
	);
	LUT2 #(
		.INIT('h8)
	) name21916 (
		_w32424_,
		_w32425_,
		_w32428_
	);
	LUT2 #(
		.INIT('h8)
	) name21917 (
		_w32422_,
		_w32423_,
		_w32429_
	);
	LUT2 #(
		.INIT('h8)
	) name21918 (
		_w32420_,
		_w32421_,
		_w32430_
	);
	LUT2 #(
		.INIT('h8)
	) name21919 (
		_w32429_,
		_w32430_,
		_w32431_
	);
	LUT2 #(
		.INIT('h8)
	) name21920 (
		_w32427_,
		_w32428_,
		_w32432_
	);
	LUT2 #(
		.INIT('h8)
	) name21921 (
		_w32431_,
		_w32432_,
		_w32433_
	);
	LUT2 #(
		.INIT('h1)
	) name21922 (
		_w31950_,
		_w32433_,
		_w32434_
	);
	LUT2 #(
		.INIT('h1)
	) name21923 (
		_w32404_,
		_w32434_,
		_w32435_
	);
	LUT2 #(
		.INIT('h2)
	) name21924 (
		\wishbone_rx_fifo_fifo_reg[0][22]/P0001 ,
		_w31954_,
		_w32436_
	);
	LUT2 #(
		.INIT('h8)
	) name21925 (
		\wishbone_rx_fifo_fifo_reg[6][22]/P0001 ,
		_w31958_,
		_w32437_
	);
	LUT2 #(
		.INIT('h8)
	) name21926 (
		\wishbone_rx_fifo_fifo_reg[12][22]/P0001 ,
		_w31984_,
		_w32438_
	);
	LUT2 #(
		.INIT('h8)
	) name21927 (
		\wishbone_rx_fifo_fifo_reg[9][22]/P0001 ,
		_w31972_,
		_w32439_
	);
	LUT2 #(
		.INIT('h8)
	) name21928 (
		\wishbone_rx_fifo_fifo_reg[11][22]/P0001 ,
		_w31988_,
		_w32440_
	);
	LUT2 #(
		.INIT('h8)
	) name21929 (
		\wishbone_rx_fifo_fifo_reg[7][22]/P0001 ,
		_w31964_,
		_w32441_
	);
	LUT2 #(
		.INIT('h8)
	) name21930 (
		\wishbone_rx_fifo_fifo_reg[5][22]/P0001 ,
		_w31980_,
		_w32442_
	);
	LUT2 #(
		.INIT('h8)
	) name21931 (
		\wishbone_rx_fifo_fifo_reg[2][22]/P0001 ,
		_w31978_,
		_w32443_
	);
	LUT2 #(
		.INIT('h8)
	) name21932 (
		\wishbone_rx_fifo_fifo_reg[13][22]/P0001 ,
		_w31986_,
		_w32444_
	);
	LUT2 #(
		.INIT('h8)
	) name21933 (
		\wishbone_rx_fifo_fifo_reg[4][22]/P0001 ,
		_w31966_,
		_w32445_
	);
	LUT2 #(
		.INIT('h8)
	) name21934 (
		\wishbone_rx_fifo_fifo_reg[15][22]/P0001 ,
		_w31969_,
		_w32446_
	);
	LUT2 #(
		.INIT('h8)
	) name21935 (
		\wishbone_rx_fifo_fifo_reg[8][22]/P0001 ,
		_w31974_,
		_w32447_
	);
	LUT2 #(
		.INIT('h8)
	) name21936 (
		\wishbone_rx_fifo_fifo_reg[14][22]/P0001 ,
		_w31982_,
		_w32448_
	);
	LUT2 #(
		.INIT('h8)
	) name21937 (
		\wishbone_rx_fifo_fifo_reg[10][22]/P0001 ,
		_w31961_,
		_w32449_
	);
	LUT2 #(
		.INIT('h8)
	) name21938 (
		\wishbone_rx_fifo_fifo_reg[1][22]/P0001 ,
		_w31976_,
		_w32450_
	);
	LUT2 #(
		.INIT('h8)
	) name21939 (
		\wishbone_rx_fifo_fifo_reg[3][22]/P0001 ,
		_w31990_,
		_w32451_
	);
	LUT2 #(
		.INIT('h1)
	) name21940 (
		_w32437_,
		_w32438_,
		_w32452_
	);
	LUT2 #(
		.INIT('h1)
	) name21941 (
		_w32439_,
		_w32440_,
		_w32453_
	);
	LUT2 #(
		.INIT('h1)
	) name21942 (
		_w32441_,
		_w32442_,
		_w32454_
	);
	LUT2 #(
		.INIT('h1)
	) name21943 (
		_w32443_,
		_w32444_,
		_w32455_
	);
	LUT2 #(
		.INIT('h1)
	) name21944 (
		_w32445_,
		_w32446_,
		_w32456_
	);
	LUT2 #(
		.INIT('h1)
	) name21945 (
		_w32447_,
		_w32448_,
		_w32457_
	);
	LUT2 #(
		.INIT('h1)
	) name21946 (
		_w32449_,
		_w32450_,
		_w32458_
	);
	LUT2 #(
		.INIT('h4)
	) name21947 (
		_w32451_,
		_w32458_,
		_w32459_
	);
	LUT2 #(
		.INIT('h8)
	) name21948 (
		_w32456_,
		_w32457_,
		_w32460_
	);
	LUT2 #(
		.INIT('h8)
	) name21949 (
		_w32454_,
		_w32455_,
		_w32461_
	);
	LUT2 #(
		.INIT('h8)
	) name21950 (
		_w32452_,
		_w32453_,
		_w32462_
	);
	LUT2 #(
		.INIT('h8)
	) name21951 (
		_w32461_,
		_w32462_,
		_w32463_
	);
	LUT2 #(
		.INIT('h8)
	) name21952 (
		_w32459_,
		_w32460_,
		_w32464_
	);
	LUT2 #(
		.INIT('h8)
	) name21953 (
		_w32463_,
		_w32464_,
		_w32465_
	);
	LUT2 #(
		.INIT('h1)
	) name21954 (
		_w31950_,
		_w32465_,
		_w32466_
	);
	LUT2 #(
		.INIT('h1)
	) name21955 (
		_w32436_,
		_w32466_,
		_w32467_
	);
	LUT2 #(
		.INIT('h2)
	) name21956 (
		\wishbone_rx_fifo_fifo_reg[0][23]/P0001 ,
		_w31954_,
		_w32468_
	);
	LUT2 #(
		.INIT('h8)
	) name21957 (
		\wishbone_rx_fifo_fifo_reg[6][23]/P0001 ,
		_w31958_,
		_w32469_
	);
	LUT2 #(
		.INIT('h8)
	) name21958 (
		\wishbone_rx_fifo_fifo_reg[12][23]/P0001 ,
		_w31984_,
		_w32470_
	);
	LUT2 #(
		.INIT('h8)
	) name21959 (
		\wishbone_rx_fifo_fifo_reg[9][23]/P0001 ,
		_w31972_,
		_w32471_
	);
	LUT2 #(
		.INIT('h8)
	) name21960 (
		\wishbone_rx_fifo_fifo_reg[11][23]/P0001 ,
		_w31988_,
		_w32472_
	);
	LUT2 #(
		.INIT('h8)
	) name21961 (
		\wishbone_rx_fifo_fifo_reg[7][23]/P0001 ,
		_w31964_,
		_w32473_
	);
	LUT2 #(
		.INIT('h8)
	) name21962 (
		\wishbone_rx_fifo_fifo_reg[5][23]/P0001 ,
		_w31980_,
		_w32474_
	);
	LUT2 #(
		.INIT('h8)
	) name21963 (
		\wishbone_rx_fifo_fifo_reg[2][23]/P0001 ,
		_w31978_,
		_w32475_
	);
	LUT2 #(
		.INIT('h8)
	) name21964 (
		\wishbone_rx_fifo_fifo_reg[13][23]/P0001 ,
		_w31986_,
		_w32476_
	);
	LUT2 #(
		.INIT('h8)
	) name21965 (
		\wishbone_rx_fifo_fifo_reg[4][23]/P0001 ,
		_w31966_,
		_w32477_
	);
	LUT2 #(
		.INIT('h8)
	) name21966 (
		\wishbone_rx_fifo_fifo_reg[15][23]/P0001 ,
		_w31969_,
		_w32478_
	);
	LUT2 #(
		.INIT('h8)
	) name21967 (
		\wishbone_rx_fifo_fifo_reg[8][23]/P0001 ,
		_w31974_,
		_w32479_
	);
	LUT2 #(
		.INIT('h8)
	) name21968 (
		\wishbone_rx_fifo_fifo_reg[14][23]/P0001 ,
		_w31982_,
		_w32480_
	);
	LUT2 #(
		.INIT('h8)
	) name21969 (
		\wishbone_rx_fifo_fifo_reg[10][23]/P0001 ,
		_w31961_,
		_w32481_
	);
	LUT2 #(
		.INIT('h8)
	) name21970 (
		\wishbone_rx_fifo_fifo_reg[1][23]/P0001 ,
		_w31976_,
		_w32482_
	);
	LUT2 #(
		.INIT('h8)
	) name21971 (
		\wishbone_rx_fifo_fifo_reg[3][23]/P0001 ,
		_w31990_,
		_w32483_
	);
	LUT2 #(
		.INIT('h1)
	) name21972 (
		_w32469_,
		_w32470_,
		_w32484_
	);
	LUT2 #(
		.INIT('h1)
	) name21973 (
		_w32471_,
		_w32472_,
		_w32485_
	);
	LUT2 #(
		.INIT('h1)
	) name21974 (
		_w32473_,
		_w32474_,
		_w32486_
	);
	LUT2 #(
		.INIT('h1)
	) name21975 (
		_w32475_,
		_w32476_,
		_w32487_
	);
	LUT2 #(
		.INIT('h1)
	) name21976 (
		_w32477_,
		_w32478_,
		_w32488_
	);
	LUT2 #(
		.INIT('h1)
	) name21977 (
		_w32479_,
		_w32480_,
		_w32489_
	);
	LUT2 #(
		.INIT('h1)
	) name21978 (
		_w32481_,
		_w32482_,
		_w32490_
	);
	LUT2 #(
		.INIT('h4)
	) name21979 (
		_w32483_,
		_w32490_,
		_w32491_
	);
	LUT2 #(
		.INIT('h8)
	) name21980 (
		_w32488_,
		_w32489_,
		_w32492_
	);
	LUT2 #(
		.INIT('h8)
	) name21981 (
		_w32486_,
		_w32487_,
		_w32493_
	);
	LUT2 #(
		.INIT('h8)
	) name21982 (
		_w32484_,
		_w32485_,
		_w32494_
	);
	LUT2 #(
		.INIT('h8)
	) name21983 (
		_w32493_,
		_w32494_,
		_w32495_
	);
	LUT2 #(
		.INIT('h8)
	) name21984 (
		_w32491_,
		_w32492_,
		_w32496_
	);
	LUT2 #(
		.INIT('h8)
	) name21985 (
		_w32495_,
		_w32496_,
		_w32497_
	);
	LUT2 #(
		.INIT('h1)
	) name21986 (
		_w31950_,
		_w32497_,
		_w32498_
	);
	LUT2 #(
		.INIT('h1)
	) name21987 (
		_w32468_,
		_w32498_,
		_w32499_
	);
	LUT2 #(
		.INIT('h2)
	) name21988 (
		\wishbone_rx_fifo_fifo_reg[0][24]/P0001 ,
		_w31954_,
		_w32500_
	);
	LUT2 #(
		.INIT('h8)
	) name21989 (
		\wishbone_rx_fifo_fifo_reg[9][24]/P0001 ,
		_w31972_,
		_w32501_
	);
	LUT2 #(
		.INIT('h8)
	) name21990 (
		\wishbone_rx_fifo_fifo_reg[8][24]/P0001 ,
		_w31974_,
		_w32502_
	);
	LUT2 #(
		.INIT('h8)
	) name21991 (
		\wishbone_rx_fifo_fifo_reg[12][24]/P0001 ,
		_w31984_,
		_w32503_
	);
	LUT2 #(
		.INIT('h8)
	) name21992 (
		\wishbone_rx_fifo_fifo_reg[13][24]/P0001 ,
		_w31986_,
		_w32504_
	);
	LUT2 #(
		.INIT('h8)
	) name21993 (
		\wishbone_rx_fifo_fifo_reg[2][24]/P0001 ,
		_w31978_,
		_w32505_
	);
	LUT2 #(
		.INIT('h8)
	) name21994 (
		\wishbone_rx_fifo_fifo_reg[3][24]/P0001 ,
		_w31990_,
		_w32506_
	);
	LUT2 #(
		.INIT('h8)
	) name21995 (
		\wishbone_rx_fifo_fifo_reg[4][24]/P0001 ,
		_w31966_,
		_w32507_
	);
	LUT2 #(
		.INIT('h8)
	) name21996 (
		\wishbone_rx_fifo_fifo_reg[5][24]/P0001 ,
		_w31980_,
		_w32508_
	);
	LUT2 #(
		.INIT('h8)
	) name21997 (
		\wishbone_rx_fifo_fifo_reg[10][24]/P0001 ,
		_w31961_,
		_w32509_
	);
	LUT2 #(
		.INIT('h8)
	) name21998 (
		\wishbone_rx_fifo_fifo_reg[7][24]/P0001 ,
		_w31964_,
		_w32510_
	);
	LUT2 #(
		.INIT('h8)
	) name21999 (
		\wishbone_rx_fifo_fifo_reg[1][24]/P0001 ,
		_w31976_,
		_w32511_
	);
	LUT2 #(
		.INIT('h8)
	) name22000 (
		\wishbone_rx_fifo_fifo_reg[11][24]/P0001 ,
		_w31988_,
		_w32512_
	);
	LUT2 #(
		.INIT('h8)
	) name22001 (
		\wishbone_rx_fifo_fifo_reg[6][24]/P0001 ,
		_w31958_,
		_w32513_
	);
	LUT2 #(
		.INIT('h8)
	) name22002 (
		\wishbone_rx_fifo_fifo_reg[15][24]/P0001 ,
		_w31969_,
		_w32514_
	);
	LUT2 #(
		.INIT('h8)
	) name22003 (
		\wishbone_rx_fifo_fifo_reg[14][24]/P0001 ,
		_w31982_,
		_w32515_
	);
	LUT2 #(
		.INIT('h1)
	) name22004 (
		_w32501_,
		_w32502_,
		_w32516_
	);
	LUT2 #(
		.INIT('h1)
	) name22005 (
		_w32503_,
		_w32504_,
		_w32517_
	);
	LUT2 #(
		.INIT('h1)
	) name22006 (
		_w32505_,
		_w32506_,
		_w32518_
	);
	LUT2 #(
		.INIT('h1)
	) name22007 (
		_w32507_,
		_w32508_,
		_w32519_
	);
	LUT2 #(
		.INIT('h1)
	) name22008 (
		_w32509_,
		_w32510_,
		_w32520_
	);
	LUT2 #(
		.INIT('h1)
	) name22009 (
		_w32511_,
		_w32512_,
		_w32521_
	);
	LUT2 #(
		.INIT('h1)
	) name22010 (
		_w32513_,
		_w32514_,
		_w32522_
	);
	LUT2 #(
		.INIT('h4)
	) name22011 (
		_w32515_,
		_w32522_,
		_w32523_
	);
	LUT2 #(
		.INIT('h8)
	) name22012 (
		_w32520_,
		_w32521_,
		_w32524_
	);
	LUT2 #(
		.INIT('h8)
	) name22013 (
		_w32518_,
		_w32519_,
		_w32525_
	);
	LUT2 #(
		.INIT('h8)
	) name22014 (
		_w32516_,
		_w32517_,
		_w32526_
	);
	LUT2 #(
		.INIT('h8)
	) name22015 (
		_w32525_,
		_w32526_,
		_w32527_
	);
	LUT2 #(
		.INIT('h8)
	) name22016 (
		_w32523_,
		_w32524_,
		_w32528_
	);
	LUT2 #(
		.INIT('h8)
	) name22017 (
		_w32527_,
		_w32528_,
		_w32529_
	);
	LUT2 #(
		.INIT('h1)
	) name22018 (
		_w31950_,
		_w32529_,
		_w32530_
	);
	LUT2 #(
		.INIT('h1)
	) name22019 (
		_w32500_,
		_w32530_,
		_w32531_
	);
	LUT2 #(
		.INIT('h2)
	) name22020 (
		\wishbone_rx_fifo_fifo_reg[0][25]/P0001 ,
		_w31954_,
		_w32532_
	);
	LUT2 #(
		.INIT('h8)
	) name22021 (
		\wishbone_rx_fifo_fifo_reg[6][25]/P0001 ,
		_w31958_,
		_w32533_
	);
	LUT2 #(
		.INIT('h8)
	) name22022 (
		\wishbone_rx_fifo_fifo_reg[10][25]/P0001 ,
		_w31961_,
		_w32534_
	);
	LUT2 #(
		.INIT('h8)
	) name22023 (
		\wishbone_rx_fifo_fifo_reg[7][25]/P0001 ,
		_w31964_,
		_w32535_
	);
	LUT2 #(
		.INIT('h8)
	) name22024 (
		\wishbone_rx_fifo_fifo_reg[4][25]/P0001 ,
		_w31966_,
		_w32536_
	);
	LUT2 #(
		.INIT('h8)
	) name22025 (
		\wishbone_rx_fifo_fifo_reg[15][25]/P0001 ,
		_w31969_,
		_w32537_
	);
	LUT2 #(
		.INIT('h8)
	) name22026 (
		\wishbone_rx_fifo_fifo_reg[9][25]/P0001 ,
		_w31972_,
		_w32538_
	);
	LUT2 #(
		.INIT('h8)
	) name22027 (
		\wishbone_rx_fifo_fifo_reg[8][25]/P0001 ,
		_w31974_,
		_w32539_
	);
	LUT2 #(
		.INIT('h8)
	) name22028 (
		\wishbone_rx_fifo_fifo_reg[3][25]/P0001 ,
		_w31990_,
		_w32540_
	);
	LUT2 #(
		.INIT('h8)
	) name22029 (
		\wishbone_rx_fifo_fifo_reg[11][25]/P0001 ,
		_w31988_,
		_w32541_
	);
	LUT2 #(
		.INIT('h8)
	) name22030 (
		\wishbone_rx_fifo_fifo_reg[5][25]/P0001 ,
		_w31980_,
		_w32542_
	);
	LUT2 #(
		.INIT('h8)
	) name22031 (
		\wishbone_rx_fifo_fifo_reg[14][25]/P0001 ,
		_w31982_,
		_w32543_
	);
	LUT2 #(
		.INIT('h8)
	) name22032 (
		\wishbone_rx_fifo_fifo_reg[12][25]/P0001 ,
		_w31984_,
		_w32544_
	);
	LUT2 #(
		.INIT('h8)
	) name22033 (
		\wishbone_rx_fifo_fifo_reg[13][25]/P0001 ,
		_w31986_,
		_w32545_
	);
	LUT2 #(
		.INIT('h8)
	) name22034 (
		\wishbone_rx_fifo_fifo_reg[2][25]/P0001 ,
		_w31978_,
		_w32546_
	);
	LUT2 #(
		.INIT('h8)
	) name22035 (
		\wishbone_rx_fifo_fifo_reg[1][25]/P0001 ,
		_w31976_,
		_w32547_
	);
	LUT2 #(
		.INIT('h1)
	) name22036 (
		_w32533_,
		_w32534_,
		_w32548_
	);
	LUT2 #(
		.INIT('h1)
	) name22037 (
		_w32535_,
		_w32536_,
		_w32549_
	);
	LUT2 #(
		.INIT('h1)
	) name22038 (
		_w32537_,
		_w32538_,
		_w32550_
	);
	LUT2 #(
		.INIT('h1)
	) name22039 (
		_w32539_,
		_w32540_,
		_w32551_
	);
	LUT2 #(
		.INIT('h1)
	) name22040 (
		_w32541_,
		_w32542_,
		_w32552_
	);
	LUT2 #(
		.INIT('h1)
	) name22041 (
		_w32543_,
		_w32544_,
		_w32553_
	);
	LUT2 #(
		.INIT('h1)
	) name22042 (
		_w32545_,
		_w32546_,
		_w32554_
	);
	LUT2 #(
		.INIT('h4)
	) name22043 (
		_w32547_,
		_w32554_,
		_w32555_
	);
	LUT2 #(
		.INIT('h8)
	) name22044 (
		_w32552_,
		_w32553_,
		_w32556_
	);
	LUT2 #(
		.INIT('h8)
	) name22045 (
		_w32550_,
		_w32551_,
		_w32557_
	);
	LUT2 #(
		.INIT('h8)
	) name22046 (
		_w32548_,
		_w32549_,
		_w32558_
	);
	LUT2 #(
		.INIT('h8)
	) name22047 (
		_w32557_,
		_w32558_,
		_w32559_
	);
	LUT2 #(
		.INIT('h8)
	) name22048 (
		_w32555_,
		_w32556_,
		_w32560_
	);
	LUT2 #(
		.INIT('h8)
	) name22049 (
		_w32559_,
		_w32560_,
		_w32561_
	);
	LUT2 #(
		.INIT('h1)
	) name22050 (
		_w31950_,
		_w32561_,
		_w32562_
	);
	LUT2 #(
		.INIT('h1)
	) name22051 (
		_w32532_,
		_w32562_,
		_w32563_
	);
	LUT2 #(
		.INIT('h2)
	) name22052 (
		\wishbone_rx_fifo_fifo_reg[0][26]/P0001 ,
		_w31954_,
		_w32564_
	);
	LUT2 #(
		.INIT('h8)
	) name22053 (
		\wishbone_rx_fifo_fifo_reg[9][26]/P0001 ,
		_w31972_,
		_w32565_
	);
	LUT2 #(
		.INIT('h8)
	) name22054 (
		\wishbone_rx_fifo_fifo_reg[3][26]/P0001 ,
		_w31990_,
		_w32566_
	);
	LUT2 #(
		.INIT('h8)
	) name22055 (
		\wishbone_rx_fifo_fifo_reg[6][26]/P0001 ,
		_w31958_,
		_w32567_
	);
	LUT2 #(
		.INIT('h8)
	) name22056 (
		\wishbone_rx_fifo_fifo_reg[15][26]/P0001 ,
		_w31969_,
		_w32568_
	);
	LUT2 #(
		.INIT('h8)
	) name22057 (
		\wishbone_rx_fifo_fifo_reg[8][26]/P0001 ,
		_w31974_,
		_w32569_
	);
	LUT2 #(
		.INIT('h8)
	) name22058 (
		\wishbone_rx_fifo_fifo_reg[5][26]/P0001 ,
		_w31980_,
		_w32570_
	);
	LUT2 #(
		.INIT('h8)
	) name22059 (
		\wishbone_rx_fifo_fifo_reg[13][26]/P0001 ,
		_w31986_,
		_w32571_
	);
	LUT2 #(
		.INIT('h8)
	) name22060 (
		\wishbone_rx_fifo_fifo_reg[4][26]/P0001 ,
		_w31966_,
		_w32572_
	);
	LUT2 #(
		.INIT('h8)
	) name22061 (
		\wishbone_rx_fifo_fifo_reg[14][26]/P0001 ,
		_w31982_,
		_w32573_
	);
	LUT2 #(
		.INIT('h8)
	) name22062 (
		\wishbone_rx_fifo_fifo_reg[12][26]/P0001 ,
		_w31984_,
		_w32574_
	);
	LUT2 #(
		.INIT('h8)
	) name22063 (
		\wishbone_rx_fifo_fifo_reg[7][26]/P0001 ,
		_w31964_,
		_w32575_
	);
	LUT2 #(
		.INIT('h8)
	) name22064 (
		\wishbone_rx_fifo_fifo_reg[2][26]/P0001 ,
		_w31978_,
		_w32576_
	);
	LUT2 #(
		.INIT('h8)
	) name22065 (
		\wishbone_rx_fifo_fifo_reg[1][26]/P0001 ,
		_w31976_,
		_w32577_
	);
	LUT2 #(
		.INIT('h8)
	) name22066 (
		\wishbone_rx_fifo_fifo_reg[10][26]/P0001 ,
		_w31961_,
		_w32578_
	);
	LUT2 #(
		.INIT('h8)
	) name22067 (
		\wishbone_rx_fifo_fifo_reg[11][26]/P0001 ,
		_w31988_,
		_w32579_
	);
	LUT2 #(
		.INIT('h1)
	) name22068 (
		_w32565_,
		_w32566_,
		_w32580_
	);
	LUT2 #(
		.INIT('h1)
	) name22069 (
		_w32567_,
		_w32568_,
		_w32581_
	);
	LUT2 #(
		.INIT('h1)
	) name22070 (
		_w32569_,
		_w32570_,
		_w32582_
	);
	LUT2 #(
		.INIT('h1)
	) name22071 (
		_w32571_,
		_w32572_,
		_w32583_
	);
	LUT2 #(
		.INIT('h1)
	) name22072 (
		_w32573_,
		_w32574_,
		_w32584_
	);
	LUT2 #(
		.INIT('h1)
	) name22073 (
		_w32575_,
		_w32576_,
		_w32585_
	);
	LUT2 #(
		.INIT('h1)
	) name22074 (
		_w32577_,
		_w32578_,
		_w32586_
	);
	LUT2 #(
		.INIT('h4)
	) name22075 (
		_w32579_,
		_w32586_,
		_w32587_
	);
	LUT2 #(
		.INIT('h8)
	) name22076 (
		_w32584_,
		_w32585_,
		_w32588_
	);
	LUT2 #(
		.INIT('h8)
	) name22077 (
		_w32582_,
		_w32583_,
		_w32589_
	);
	LUT2 #(
		.INIT('h8)
	) name22078 (
		_w32580_,
		_w32581_,
		_w32590_
	);
	LUT2 #(
		.INIT('h8)
	) name22079 (
		_w32589_,
		_w32590_,
		_w32591_
	);
	LUT2 #(
		.INIT('h8)
	) name22080 (
		_w32587_,
		_w32588_,
		_w32592_
	);
	LUT2 #(
		.INIT('h8)
	) name22081 (
		_w32591_,
		_w32592_,
		_w32593_
	);
	LUT2 #(
		.INIT('h1)
	) name22082 (
		_w31950_,
		_w32593_,
		_w32594_
	);
	LUT2 #(
		.INIT('h1)
	) name22083 (
		_w32564_,
		_w32594_,
		_w32595_
	);
	LUT2 #(
		.INIT('h8)
	) name22084 (
		\wishbone_rx_fifo_fifo_reg[12][27]/P0001 ,
		_w31984_,
		_w32596_
	);
	LUT2 #(
		.INIT('h8)
	) name22085 (
		\wishbone_rx_fifo_fifo_reg[3][27]/P0001 ,
		_w31990_,
		_w32597_
	);
	LUT2 #(
		.INIT('h8)
	) name22086 (
		\wishbone_rx_fifo_fifo_reg[1][27]/P0001 ,
		_w31976_,
		_w32598_
	);
	LUT2 #(
		.INIT('h8)
	) name22087 (
		\wishbone_rx_fifo_fifo_reg[11][27]/P0001 ,
		_w31988_,
		_w32599_
	);
	LUT2 #(
		.INIT('h8)
	) name22088 (
		\wishbone_rx_fifo_fifo_reg[9][27]/P0001 ,
		_w31972_,
		_w32600_
	);
	LUT2 #(
		.INIT('h8)
	) name22089 (
		\wishbone_rx_fifo_fifo_reg[6][27]/P0001 ,
		_w31958_,
		_w32601_
	);
	LUT2 #(
		.INIT('h8)
	) name22090 (
		\wishbone_rx_fifo_fifo_reg[15][27]/P0001 ,
		_w31969_,
		_w32602_
	);
	LUT2 #(
		.INIT('h8)
	) name22091 (
		\wishbone_rx_fifo_fifo_reg[7][27]/P0001 ,
		_w31964_,
		_w32603_
	);
	LUT2 #(
		.INIT('h8)
	) name22092 (
		\wishbone_rx_fifo_fifo_reg[8][27]/P0001 ,
		_w31974_,
		_w32604_
	);
	LUT2 #(
		.INIT('h8)
	) name22093 (
		\wishbone_rx_fifo_fifo_reg[13][27]/P0001 ,
		_w31986_,
		_w32605_
	);
	LUT2 #(
		.INIT('h8)
	) name22094 (
		\wishbone_rx_fifo_fifo_reg[14][27]/P0001 ,
		_w31982_,
		_w32606_
	);
	LUT2 #(
		.INIT('h8)
	) name22095 (
		\wishbone_rx_fifo_fifo_reg[5][27]/P0001 ,
		_w31980_,
		_w32607_
	);
	LUT2 #(
		.INIT('h8)
	) name22096 (
		\wishbone_rx_fifo_fifo_reg[10][27]/P0001 ,
		_w31961_,
		_w32608_
	);
	LUT2 #(
		.INIT('h8)
	) name22097 (
		\wishbone_rx_fifo_fifo_reg[2][27]/P0001 ,
		_w31978_,
		_w32609_
	);
	LUT2 #(
		.INIT('h8)
	) name22098 (
		\wishbone_rx_fifo_fifo_reg[4][27]/P0001 ,
		_w31966_,
		_w32610_
	);
	LUT2 #(
		.INIT('h1)
	) name22099 (
		_w31950_,
		_w32596_,
		_w32611_
	);
	LUT2 #(
		.INIT('h1)
	) name22100 (
		_w32597_,
		_w32598_,
		_w32612_
	);
	LUT2 #(
		.INIT('h1)
	) name22101 (
		_w32599_,
		_w32600_,
		_w32613_
	);
	LUT2 #(
		.INIT('h1)
	) name22102 (
		_w32601_,
		_w32602_,
		_w32614_
	);
	LUT2 #(
		.INIT('h1)
	) name22103 (
		_w32603_,
		_w32604_,
		_w32615_
	);
	LUT2 #(
		.INIT('h1)
	) name22104 (
		_w32605_,
		_w32606_,
		_w32616_
	);
	LUT2 #(
		.INIT('h1)
	) name22105 (
		_w32607_,
		_w32608_,
		_w32617_
	);
	LUT2 #(
		.INIT('h1)
	) name22106 (
		_w32609_,
		_w32610_,
		_w32618_
	);
	LUT2 #(
		.INIT('h8)
	) name22107 (
		_w32617_,
		_w32618_,
		_w32619_
	);
	LUT2 #(
		.INIT('h8)
	) name22108 (
		_w32615_,
		_w32616_,
		_w32620_
	);
	LUT2 #(
		.INIT('h8)
	) name22109 (
		_w32613_,
		_w32614_,
		_w32621_
	);
	LUT2 #(
		.INIT('h8)
	) name22110 (
		_w32611_,
		_w32612_,
		_w32622_
	);
	LUT2 #(
		.INIT('h8)
	) name22111 (
		_w32621_,
		_w32622_,
		_w32623_
	);
	LUT2 #(
		.INIT('h8)
	) name22112 (
		_w32619_,
		_w32620_,
		_w32624_
	);
	LUT2 #(
		.INIT('h8)
	) name22113 (
		_w32623_,
		_w32624_,
		_w32625_
	);
	LUT2 #(
		.INIT('h4)
	) name22114 (
		\wishbone_rx_fifo_fifo_reg[0][27]/P0001 ,
		_w31950_,
		_w32626_
	);
	LUT2 #(
		.INIT('h1)
	) name22115 (
		_w32625_,
		_w32626_,
		_w32627_
	);
	LUT2 #(
		.INIT('h8)
	) name22116 (
		\wishbone_rx_fifo_fifo_reg[0][27]/P0001 ,
		_w31953_,
		_w32628_
	);
	LUT2 #(
		.INIT('h1)
	) name22117 (
		_w32627_,
		_w32628_,
		_w32629_
	);
	LUT2 #(
		.INIT('h8)
	) name22118 (
		\wishbone_rx_fifo_fifo_reg[12][28]/P0001 ,
		_w31984_,
		_w32630_
	);
	LUT2 #(
		.INIT('h8)
	) name22119 (
		\wishbone_rx_fifo_fifo_reg[15][28]/P0001 ,
		_w31969_,
		_w32631_
	);
	LUT2 #(
		.INIT('h8)
	) name22120 (
		\wishbone_rx_fifo_fifo_reg[2][28]/P0001 ,
		_w31978_,
		_w32632_
	);
	LUT2 #(
		.INIT('h8)
	) name22121 (
		\wishbone_rx_fifo_fifo_reg[13][28]/P0001 ,
		_w31986_,
		_w32633_
	);
	LUT2 #(
		.INIT('h8)
	) name22122 (
		\wishbone_rx_fifo_fifo_reg[5][28]/P0001 ,
		_w31980_,
		_w32634_
	);
	LUT2 #(
		.INIT('h8)
	) name22123 (
		\wishbone_rx_fifo_fifo_reg[6][28]/P0001 ,
		_w31958_,
		_w32635_
	);
	LUT2 #(
		.INIT('h8)
	) name22124 (
		\wishbone_rx_fifo_fifo_reg[8][28]/P0001 ,
		_w31974_,
		_w32636_
	);
	LUT2 #(
		.INIT('h8)
	) name22125 (
		\wishbone_rx_fifo_fifo_reg[11][28]/P0001 ,
		_w31988_,
		_w32637_
	);
	LUT2 #(
		.INIT('h8)
	) name22126 (
		\wishbone_rx_fifo_fifo_reg[9][28]/P0001 ,
		_w31972_,
		_w32638_
	);
	LUT2 #(
		.INIT('h8)
	) name22127 (
		\wishbone_rx_fifo_fifo_reg[1][28]/P0001 ,
		_w31976_,
		_w32639_
	);
	LUT2 #(
		.INIT('h8)
	) name22128 (
		\wishbone_rx_fifo_fifo_reg[4][28]/P0001 ,
		_w31966_,
		_w32640_
	);
	LUT2 #(
		.INIT('h8)
	) name22129 (
		\wishbone_rx_fifo_fifo_reg[14][28]/P0001 ,
		_w31982_,
		_w32641_
	);
	LUT2 #(
		.INIT('h8)
	) name22130 (
		\wishbone_rx_fifo_fifo_reg[10][28]/P0001 ,
		_w31961_,
		_w32642_
	);
	LUT2 #(
		.INIT('h8)
	) name22131 (
		\wishbone_rx_fifo_fifo_reg[3][28]/P0001 ,
		_w31990_,
		_w32643_
	);
	LUT2 #(
		.INIT('h8)
	) name22132 (
		\wishbone_rx_fifo_fifo_reg[7][28]/P0001 ,
		_w31964_,
		_w32644_
	);
	LUT2 #(
		.INIT('h1)
	) name22133 (
		_w31950_,
		_w32630_,
		_w32645_
	);
	LUT2 #(
		.INIT('h1)
	) name22134 (
		_w32631_,
		_w32632_,
		_w32646_
	);
	LUT2 #(
		.INIT('h1)
	) name22135 (
		_w32633_,
		_w32634_,
		_w32647_
	);
	LUT2 #(
		.INIT('h1)
	) name22136 (
		_w32635_,
		_w32636_,
		_w32648_
	);
	LUT2 #(
		.INIT('h1)
	) name22137 (
		_w32637_,
		_w32638_,
		_w32649_
	);
	LUT2 #(
		.INIT('h1)
	) name22138 (
		_w32639_,
		_w32640_,
		_w32650_
	);
	LUT2 #(
		.INIT('h1)
	) name22139 (
		_w32641_,
		_w32642_,
		_w32651_
	);
	LUT2 #(
		.INIT('h1)
	) name22140 (
		_w32643_,
		_w32644_,
		_w32652_
	);
	LUT2 #(
		.INIT('h8)
	) name22141 (
		_w32651_,
		_w32652_,
		_w32653_
	);
	LUT2 #(
		.INIT('h8)
	) name22142 (
		_w32649_,
		_w32650_,
		_w32654_
	);
	LUT2 #(
		.INIT('h8)
	) name22143 (
		_w32647_,
		_w32648_,
		_w32655_
	);
	LUT2 #(
		.INIT('h8)
	) name22144 (
		_w32645_,
		_w32646_,
		_w32656_
	);
	LUT2 #(
		.INIT('h8)
	) name22145 (
		_w32655_,
		_w32656_,
		_w32657_
	);
	LUT2 #(
		.INIT('h8)
	) name22146 (
		_w32653_,
		_w32654_,
		_w32658_
	);
	LUT2 #(
		.INIT('h8)
	) name22147 (
		_w32657_,
		_w32658_,
		_w32659_
	);
	LUT2 #(
		.INIT('h4)
	) name22148 (
		\wishbone_rx_fifo_fifo_reg[0][28]/P0001 ,
		_w31950_,
		_w32660_
	);
	LUT2 #(
		.INIT('h1)
	) name22149 (
		_w32659_,
		_w32660_,
		_w32661_
	);
	LUT2 #(
		.INIT('h8)
	) name22150 (
		\wishbone_rx_fifo_fifo_reg[0][28]/P0001 ,
		_w31953_,
		_w32662_
	);
	LUT2 #(
		.INIT('h1)
	) name22151 (
		_w32661_,
		_w32662_,
		_w32663_
	);
	LUT2 #(
		.INIT('h8)
	) name22152 (
		\wishbone_rx_fifo_fifo_reg[10][29]/P0001 ,
		_w31961_,
		_w32664_
	);
	LUT2 #(
		.INIT('h8)
	) name22153 (
		\wishbone_rx_fifo_fifo_reg[13][29]/P0001 ,
		_w31986_,
		_w32665_
	);
	LUT2 #(
		.INIT('h8)
	) name22154 (
		\wishbone_rx_fifo_fifo_reg[14][29]/P0001 ,
		_w31982_,
		_w32666_
	);
	LUT2 #(
		.INIT('h8)
	) name22155 (
		\wishbone_rx_fifo_fifo_reg[1][29]/P0001 ,
		_w31976_,
		_w32667_
	);
	LUT2 #(
		.INIT('h8)
	) name22156 (
		\wishbone_rx_fifo_fifo_reg[5][29]/P0001 ,
		_w31980_,
		_w32668_
	);
	LUT2 #(
		.INIT('h8)
	) name22157 (
		\wishbone_rx_fifo_fifo_reg[8][29]/P0001 ,
		_w31974_,
		_w32669_
	);
	LUT2 #(
		.INIT('h8)
	) name22158 (
		\wishbone_rx_fifo_fifo_reg[6][29]/P0001 ,
		_w31958_,
		_w32670_
	);
	LUT2 #(
		.INIT('h8)
	) name22159 (
		\wishbone_rx_fifo_fifo_reg[9][29]/P0001 ,
		_w31972_,
		_w32671_
	);
	LUT2 #(
		.INIT('h8)
	) name22160 (
		\wishbone_rx_fifo_fifo_reg[7][29]/P0001 ,
		_w31964_,
		_w32672_
	);
	LUT2 #(
		.INIT('h8)
	) name22161 (
		\wishbone_rx_fifo_fifo_reg[12][29]/P0001 ,
		_w31984_,
		_w32673_
	);
	LUT2 #(
		.INIT('h8)
	) name22162 (
		\wishbone_rx_fifo_fifo_reg[4][29]/P0001 ,
		_w31966_,
		_w32674_
	);
	LUT2 #(
		.INIT('h8)
	) name22163 (
		\wishbone_rx_fifo_fifo_reg[3][29]/P0001 ,
		_w31990_,
		_w32675_
	);
	LUT2 #(
		.INIT('h8)
	) name22164 (
		\wishbone_rx_fifo_fifo_reg[15][29]/P0001 ,
		_w31969_,
		_w32676_
	);
	LUT2 #(
		.INIT('h8)
	) name22165 (
		\wishbone_rx_fifo_fifo_reg[11][29]/P0001 ,
		_w31988_,
		_w32677_
	);
	LUT2 #(
		.INIT('h8)
	) name22166 (
		\wishbone_rx_fifo_fifo_reg[2][29]/P0001 ,
		_w31978_,
		_w32678_
	);
	LUT2 #(
		.INIT('h1)
	) name22167 (
		_w31950_,
		_w32664_,
		_w32679_
	);
	LUT2 #(
		.INIT('h1)
	) name22168 (
		_w32665_,
		_w32666_,
		_w32680_
	);
	LUT2 #(
		.INIT('h1)
	) name22169 (
		_w32667_,
		_w32668_,
		_w32681_
	);
	LUT2 #(
		.INIT('h1)
	) name22170 (
		_w32669_,
		_w32670_,
		_w32682_
	);
	LUT2 #(
		.INIT('h1)
	) name22171 (
		_w32671_,
		_w32672_,
		_w32683_
	);
	LUT2 #(
		.INIT('h1)
	) name22172 (
		_w32673_,
		_w32674_,
		_w32684_
	);
	LUT2 #(
		.INIT('h1)
	) name22173 (
		_w32675_,
		_w32676_,
		_w32685_
	);
	LUT2 #(
		.INIT('h1)
	) name22174 (
		_w32677_,
		_w32678_,
		_w32686_
	);
	LUT2 #(
		.INIT('h8)
	) name22175 (
		_w32685_,
		_w32686_,
		_w32687_
	);
	LUT2 #(
		.INIT('h8)
	) name22176 (
		_w32683_,
		_w32684_,
		_w32688_
	);
	LUT2 #(
		.INIT('h8)
	) name22177 (
		_w32681_,
		_w32682_,
		_w32689_
	);
	LUT2 #(
		.INIT('h8)
	) name22178 (
		_w32679_,
		_w32680_,
		_w32690_
	);
	LUT2 #(
		.INIT('h8)
	) name22179 (
		_w32689_,
		_w32690_,
		_w32691_
	);
	LUT2 #(
		.INIT('h8)
	) name22180 (
		_w32687_,
		_w32688_,
		_w32692_
	);
	LUT2 #(
		.INIT('h8)
	) name22181 (
		_w32691_,
		_w32692_,
		_w32693_
	);
	LUT2 #(
		.INIT('h4)
	) name22182 (
		\wishbone_rx_fifo_fifo_reg[0][29]/P0001 ,
		_w31950_,
		_w32694_
	);
	LUT2 #(
		.INIT('h1)
	) name22183 (
		_w32693_,
		_w32694_,
		_w32695_
	);
	LUT2 #(
		.INIT('h8)
	) name22184 (
		\wishbone_rx_fifo_fifo_reg[0][29]/P0001 ,
		_w31953_,
		_w32696_
	);
	LUT2 #(
		.INIT('h1)
	) name22185 (
		_w32695_,
		_w32696_,
		_w32697_
	);
	LUT2 #(
		.INIT('h2)
	) name22186 (
		\wishbone_rx_fifo_fifo_reg[0][2]/P0001 ,
		_w31954_,
		_w32698_
	);
	LUT2 #(
		.INIT('h8)
	) name22187 (
		\wishbone_rx_fifo_fifo_reg[3][2]/P0001 ,
		_w31990_,
		_w32699_
	);
	LUT2 #(
		.INIT('h8)
	) name22188 (
		\wishbone_rx_fifo_fifo_reg[9][2]/P0001 ,
		_w31972_,
		_w32700_
	);
	LUT2 #(
		.INIT('h8)
	) name22189 (
		\wishbone_rx_fifo_fifo_reg[5][2]/P0001 ,
		_w31980_,
		_w32701_
	);
	LUT2 #(
		.INIT('h8)
	) name22190 (
		\wishbone_rx_fifo_fifo_reg[7][2]/P0001 ,
		_w31964_,
		_w32702_
	);
	LUT2 #(
		.INIT('h8)
	) name22191 (
		\wishbone_rx_fifo_fifo_reg[10][2]/P0001 ,
		_w31961_,
		_w32703_
	);
	LUT2 #(
		.INIT('h8)
	) name22192 (
		\wishbone_rx_fifo_fifo_reg[6][2]/P0001 ,
		_w31958_,
		_w32704_
	);
	LUT2 #(
		.INIT('h8)
	) name22193 (
		\wishbone_rx_fifo_fifo_reg[12][2]/P0001 ,
		_w31984_,
		_w32705_
	);
	LUT2 #(
		.INIT('h8)
	) name22194 (
		\wishbone_rx_fifo_fifo_reg[4][2]/P0001 ,
		_w31966_,
		_w32706_
	);
	LUT2 #(
		.INIT('h8)
	) name22195 (
		\wishbone_rx_fifo_fifo_reg[1][2]/P0001 ,
		_w31976_,
		_w32707_
	);
	LUT2 #(
		.INIT('h8)
	) name22196 (
		\wishbone_rx_fifo_fifo_reg[13][2]/P0001 ,
		_w31986_,
		_w32708_
	);
	LUT2 #(
		.INIT('h8)
	) name22197 (
		\wishbone_rx_fifo_fifo_reg[2][2]/P0001 ,
		_w31978_,
		_w32709_
	);
	LUT2 #(
		.INIT('h8)
	) name22198 (
		\wishbone_rx_fifo_fifo_reg[14][2]/P0001 ,
		_w31982_,
		_w32710_
	);
	LUT2 #(
		.INIT('h8)
	) name22199 (
		\wishbone_rx_fifo_fifo_reg[8][2]/P0001 ,
		_w31974_,
		_w32711_
	);
	LUT2 #(
		.INIT('h8)
	) name22200 (
		\wishbone_rx_fifo_fifo_reg[11][2]/P0001 ,
		_w31988_,
		_w32712_
	);
	LUT2 #(
		.INIT('h8)
	) name22201 (
		\wishbone_rx_fifo_fifo_reg[15][2]/P0001 ,
		_w31969_,
		_w32713_
	);
	LUT2 #(
		.INIT('h1)
	) name22202 (
		_w32699_,
		_w32700_,
		_w32714_
	);
	LUT2 #(
		.INIT('h1)
	) name22203 (
		_w32701_,
		_w32702_,
		_w32715_
	);
	LUT2 #(
		.INIT('h1)
	) name22204 (
		_w32703_,
		_w32704_,
		_w32716_
	);
	LUT2 #(
		.INIT('h1)
	) name22205 (
		_w32705_,
		_w32706_,
		_w32717_
	);
	LUT2 #(
		.INIT('h1)
	) name22206 (
		_w32707_,
		_w32708_,
		_w32718_
	);
	LUT2 #(
		.INIT('h1)
	) name22207 (
		_w32709_,
		_w32710_,
		_w32719_
	);
	LUT2 #(
		.INIT('h1)
	) name22208 (
		_w32711_,
		_w32712_,
		_w32720_
	);
	LUT2 #(
		.INIT('h4)
	) name22209 (
		_w32713_,
		_w32720_,
		_w32721_
	);
	LUT2 #(
		.INIT('h8)
	) name22210 (
		_w32718_,
		_w32719_,
		_w32722_
	);
	LUT2 #(
		.INIT('h8)
	) name22211 (
		_w32716_,
		_w32717_,
		_w32723_
	);
	LUT2 #(
		.INIT('h8)
	) name22212 (
		_w32714_,
		_w32715_,
		_w32724_
	);
	LUT2 #(
		.INIT('h8)
	) name22213 (
		_w32723_,
		_w32724_,
		_w32725_
	);
	LUT2 #(
		.INIT('h8)
	) name22214 (
		_w32721_,
		_w32722_,
		_w32726_
	);
	LUT2 #(
		.INIT('h8)
	) name22215 (
		_w32725_,
		_w32726_,
		_w32727_
	);
	LUT2 #(
		.INIT('h1)
	) name22216 (
		_w31950_,
		_w32727_,
		_w32728_
	);
	LUT2 #(
		.INIT('h1)
	) name22217 (
		_w32698_,
		_w32728_,
		_w32729_
	);
	LUT2 #(
		.INIT('h2)
	) name22218 (
		\wishbone_rx_fifo_fifo_reg[0][30]/P0001 ,
		_w31954_,
		_w32730_
	);
	LUT2 #(
		.INIT('h8)
	) name22219 (
		\wishbone_rx_fifo_fifo_reg[3][30]/P0001 ,
		_w31990_,
		_w32731_
	);
	LUT2 #(
		.INIT('h8)
	) name22220 (
		\wishbone_rx_fifo_fifo_reg[5][30]/P0001 ,
		_w31980_,
		_w32732_
	);
	LUT2 #(
		.INIT('h8)
	) name22221 (
		\wishbone_rx_fifo_fifo_reg[15][30]/P0001 ,
		_w31969_,
		_w32733_
	);
	LUT2 #(
		.INIT('h8)
	) name22222 (
		\wishbone_rx_fifo_fifo_reg[2][30]/P0001 ,
		_w31978_,
		_w32734_
	);
	LUT2 #(
		.INIT('h8)
	) name22223 (
		\wishbone_rx_fifo_fifo_reg[13][30]/P0001 ,
		_w31986_,
		_w32735_
	);
	LUT2 #(
		.INIT('h8)
	) name22224 (
		\wishbone_rx_fifo_fifo_reg[9][30]/P0001 ,
		_w31972_,
		_w32736_
	);
	LUT2 #(
		.INIT('h8)
	) name22225 (
		\wishbone_rx_fifo_fifo_reg[8][30]/P0001 ,
		_w31974_,
		_w32737_
	);
	LUT2 #(
		.INIT('h8)
	) name22226 (
		\wishbone_rx_fifo_fifo_reg[14][30]/P0001 ,
		_w31982_,
		_w32738_
	);
	LUT2 #(
		.INIT('h8)
	) name22227 (
		\wishbone_rx_fifo_fifo_reg[7][30]/P0001 ,
		_w31964_,
		_w32739_
	);
	LUT2 #(
		.INIT('h8)
	) name22228 (
		\wishbone_rx_fifo_fifo_reg[10][30]/P0001 ,
		_w31961_,
		_w32740_
	);
	LUT2 #(
		.INIT('h8)
	) name22229 (
		\wishbone_rx_fifo_fifo_reg[11][30]/P0001 ,
		_w31988_,
		_w32741_
	);
	LUT2 #(
		.INIT('h8)
	) name22230 (
		\wishbone_rx_fifo_fifo_reg[12][30]/P0001 ,
		_w31984_,
		_w32742_
	);
	LUT2 #(
		.INIT('h8)
	) name22231 (
		\wishbone_rx_fifo_fifo_reg[4][30]/P0001 ,
		_w31966_,
		_w32743_
	);
	LUT2 #(
		.INIT('h8)
	) name22232 (
		\wishbone_rx_fifo_fifo_reg[6][30]/P0001 ,
		_w31958_,
		_w32744_
	);
	LUT2 #(
		.INIT('h8)
	) name22233 (
		\wishbone_rx_fifo_fifo_reg[1][30]/P0001 ,
		_w31976_,
		_w32745_
	);
	LUT2 #(
		.INIT('h1)
	) name22234 (
		_w32731_,
		_w32732_,
		_w32746_
	);
	LUT2 #(
		.INIT('h1)
	) name22235 (
		_w32733_,
		_w32734_,
		_w32747_
	);
	LUT2 #(
		.INIT('h1)
	) name22236 (
		_w32735_,
		_w32736_,
		_w32748_
	);
	LUT2 #(
		.INIT('h1)
	) name22237 (
		_w32737_,
		_w32738_,
		_w32749_
	);
	LUT2 #(
		.INIT('h1)
	) name22238 (
		_w32739_,
		_w32740_,
		_w32750_
	);
	LUT2 #(
		.INIT('h1)
	) name22239 (
		_w32741_,
		_w32742_,
		_w32751_
	);
	LUT2 #(
		.INIT('h1)
	) name22240 (
		_w32743_,
		_w32744_,
		_w32752_
	);
	LUT2 #(
		.INIT('h4)
	) name22241 (
		_w32745_,
		_w32752_,
		_w32753_
	);
	LUT2 #(
		.INIT('h8)
	) name22242 (
		_w32750_,
		_w32751_,
		_w32754_
	);
	LUT2 #(
		.INIT('h8)
	) name22243 (
		_w32748_,
		_w32749_,
		_w32755_
	);
	LUT2 #(
		.INIT('h8)
	) name22244 (
		_w32746_,
		_w32747_,
		_w32756_
	);
	LUT2 #(
		.INIT('h8)
	) name22245 (
		_w32755_,
		_w32756_,
		_w32757_
	);
	LUT2 #(
		.INIT('h8)
	) name22246 (
		_w32753_,
		_w32754_,
		_w32758_
	);
	LUT2 #(
		.INIT('h8)
	) name22247 (
		_w32757_,
		_w32758_,
		_w32759_
	);
	LUT2 #(
		.INIT('h1)
	) name22248 (
		_w31950_,
		_w32759_,
		_w32760_
	);
	LUT2 #(
		.INIT('h1)
	) name22249 (
		_w32730_,
		_w32760_,
		_w32761_
	);
	LUT2 #(
		.INIT('h8)
	) name22250 (
		\wishbone_rx_fifo_fifo_reg[12][31]/P0001 ,
		_w31984_,
		_w32762_
	);
	LUT2 #(
		.INIT('h8)
	) name22251 (
		\wishbone_rx_fifo_fifo_reg[5][31]/P0001 ,
		_w31980_,
		_w32763_
	);
	LUT2 #(
		.INIT('h8)
	) name22252 (
		\wishbone_rx_fifo_fifo_reg[2][31]/P0001 ,
		_w31978_,
		_w32764_
	);
	LUT2 #(
		.INIT('h8)
	) name22253 (
		\wishbone_rx_fifo_fifo_reg[11][31]/P0001 ,
		_w31988_,
		_w32765_
	);
	LUT2 #(
		.INIT('h8)
	) name22254 (
		\wishbone_rx_fifo_fifo_reg[3][31]/P0001 ,
		_w31990_,
		_w32766_
	);
	LUT2 #(
		.INIT('h8)
	) name22255 (
		\wishbone_rx_fifo_fifo_reg[6][31]/P0001 ,
		_w31958_,
		_w32767_
	);
	LUT2 #(
		.INIT('h8)
	) name22256 (
		\wishbone_rx_fifo_fifo_reg[8][31]/P0001 ,
		_w31974_,
		_w32768_
	);
	LUT2 #(
		.INIT('h8)
	) name22257 (
		\wishbone_rx_fifo_fifo_reg[15][31]/P0001 ,
		_w31969_,
		_w32769_
	);
	LUT2 #(
		.INIT('h8)
	) name22258 (
		\wishbone_rx_fifo_fifo_reg[13][31]/P0001 ,
		_w31986_,
		_w32770_
	);
	LUT2 #(
		.INIT('h8)
	) name22259 (
		\wishbone_rx_fifo_fifo_reg[7][31]/P0001 ,
		_w31964_,
		_w32771_
	);
	LUT2 #(
		.INIT('h8)
	) name22260 (
		\wishbone_rx_fifo_fifo_reg[14][31]/P0001 ,
		_w31982_,
		_w32772_
	);
	LUT2 #(
		.INIT('h8)
	) name22261 (
		\wishbone_rx_fifo_fifo_reg[1][31]/P0001 ,
		_w31976_,
		_w32773_
	);
	LUT2 #(
		.INIT('h8)
	) name22262 (
		\wishbone_rx_fifo_fifo_reg[10][31]/P0001 ,
		_w31961_,
		_w32774_
	);
	LUT2 #(
		.INIT('h8)
	) name22263 (
		\wishbone_rx_fifo_fifo_reg[9][31]/P0001 ,
		_w31972_,
		_w32775_
	);
	LUT2 #(
		.INIT('h8)
	) name22264 (
		\wishbone_rx_fifo_fifo_reg[4][31]/P0001 ,
		_w31966_,
		_w32776_
	);
	LUT2 #(
		.INIT('h1)
	) name22265 (
		_w31950_,
		_w32762_,
		_w32777_
	);
	LUT2 #(
		.INIT('h1)
	) name22266 (
		_w32763_,
		_w32764_,
		_w32778_
	);
	LUT2 #(
		.INIT('h1)
	) name22267 (
		_w32765_,
		_w32766_,
		_w32779_
	);
	LUT2 #(
		.INIT('h1)
	) name22268 (
		_w32767_,
		_w32768_,
		_w32780_
	);
	LUT2 #(
		.INIT('h1)
	) name22269 (
		_w32769_,
		_w32770_,
		_w32781_
	);
	LUT2 #(
		.INIT('h1)
	) name22270 (
		_w32771_,
		_w32772_,
		_w32782_
	);
	LUT2 #(
		.INIT('h1)
	) name22271 (
		_w32773_,
		_w32774_,
		_w32783_
	);
	LUT2 #(
		.INIT('h1)
	) name22272 (
		_w32775_,
		_w32776_,
		_w32784_
	);
	LUT2 #(
		.INIT('h8)
	) name22273 (
		_w32783_,
		_w32784_,
		_w32785_
	);
	LUT2 #(
		.INIT('h8)
	) name22274 (
		_w32781_,
		_w32782_,
		_w32786_
	);
	LUT2 #(
		.INIT('h8)
	) name22275 (
		_w32779_,
		_w32780_,
		_w32787_
	);
	LUT2 #(
		.INIT('h8)
	) name22276 (
		_w32777_,
		_w32778_,
		_w32788_
	);
	LUT2 #(
		.INIT('h8)
	) name22277 (
		_w32787_,
		_w32788_,
		_w32789_
	);
	LUT2 #(
		.INIT('h8)
	) name22278 (
		_w32785_,
		_w32786_,
		_w32790_
	);
	LUT2 #(
		.INIT('h8)
	) name22279 (
		_w32789_,
		_w32790_,
		_w32791_
	);
	LUT2 #(
		.INIT('h4)
	) name22280 (
		\wishbone_rx_fifo_fifo_reg[0][31]/P0001 ,
		_w31950_,
		_w32792_
	);
	LUT2 #(
		.INIT('h1)
	) name22281 (
		_w32791_,
		_w32792_,
		_w32793_
	);
	LUT2 #(
		.INIT('h8)
	) name22282 (
		\wishbone_rx_fifo_fifo_reg[0][31]/P0001 ,
		_w31953_,
		_w32794_
	);
	LUT2 #(
		.INIT('h1)
	) name22283 (
		_w32793_,
		_w32794_,
		_w32795_
	);
	LUT2 #(
		.INIT('h2)
	) name22284 (
		\wishbone_rx_fifo_fifo_reg[0][3]/P0001 ,
		_w31954_,
		_w32796_
	);
	LUT2 #(
		.INIT('h8)
	) name22285 (
		\wishbone_rx_fifo_fifo_reg[8][3]/P0001 ,
		_w31974_,
		_w32797_
	);
	LUT2 #(
		.INIT('h8)
	) name22286 (
		\wishbone_rx_fifo_fifo_reg[7][3]/P0001 ,
		_w31964_,
		_w32798_
	);
	LUT2 #(
		.INIT('h8)
	) name22287 (
		\wishbone_rx_fifo_fifo_reg[10][3]/P0001 ,
		_w31961_,
		_w32799_
	);
	LUT2 #(
		.INIT('h8)
	) name22288 (
		\wishbone_rx_fifo_fifo_reg[12][3]/P0001 ,
		_w31984_,
		_w32800_
	);
	LUT2 #(
		.INIT('h8)
	) name22289 (
		\wishbone_rx_fifo_fifo_reg[5][3]/P0001 ,
		_w31980_,
		_w32801_
	);
	LUT2 #(
		.INIT('h8)
	) name22290 (
		\wishbone_rx_fifo_fifo_reg[1][3]/P0001 ,
		_w31976_,
		_w32802_
	);
	LUT2 #(
		.INIT('h8)
	) name22291 (
		\wishbone_rx_fifo_fifo_reg[11][3]/P0001 ,
		_w31988_,
		_w32803_
	);
	LUT2 #(
		.INIT('h8)
	) name22292 (
		\wishbone_rx_fifo_fifo_reg[4][3]/P0001 ,
		_w31966_,
		_w32804_
	);
	LUT2 #(
		.INIT('h8)
	) name22293 (
		\wishbone_rx_fifo_fifo_reg[13][3]/P0001 ,
		_w31986_,
		_w32805_
	);
	LUT2 #(
		.INIT('h8)
	) name22294 (
		\wishbone_rx_fifo_fifo_reg[6][3]/P0001 ,
		_w31958_,
		_w32806_
	);
	LUT2 #(
		.INIT('h8)
	) name22295 (
		\wishbone_rx_fifo_fifo_reg[14][3]/P0001 ,
		_w31982_,
		_w32807_
	);
	LUT2 #(
		.INIT('h8)
	) name22296 (
		\wishbone_rx_fifo_fifo_reg[15][3]/P0001 ,
		_w31969_,
		_w32808_
	);
	LUT2 #(
		.INIT('h8)
	) name22297 (
		\wishbone_rx_fifo_fifo_reg[9][3]/P0001 ,
		_w31972_,
		_w32809_
	);
	LUT2 #(
		.INIT('h8)
	) name22298 (
		\wishbone_rx_fifo_fifo_reg[2][3]/P0001 ,
		_w31978_,
		_w32810_
	);
	LUT2 #(
		.INIT('h8)
	) name22299 (
		\wishbone_rx_fifo_fifo_reg[3][3]/P0001 ,
		_w31990_,
		_w32811_
	);
	LUT2 #(
		.INIT('h1)
	) name22300 (
		_w32797_,
		_w32798_,
		_w32812_
	);
	LUT2 #(
		.INIT('h1)
	) name22301 (
		_w32799_,
		_w32800_,
		_w32813_
	);
	LUT2 #(
		.INIT('h1)
	) name22302 (
		_w32801_,
		_w32802_,
		_w32814_
	);
	LUT2 #(
		.INIT('h1)
	) name22303 (
		_w32803_,
		_w32804_,
		_w32815_
	);
	LUT2 #(
		.INIT('h1)
	) name22304 (
		_w32805_,
		_w32806_,
		_w32816_
	);
	LUT2 #(
		.INIT('h1)
	) name22305 (
		_w32807_,
		_w32808_,
		_w32817_
	);
	LUT2 #(
		.INIT('h1)
	) name22306 (
		_w32809_,
		_w32810_,
		_w32818_
	);
	LUT2 #(
		.INIT('h4)
	) name22307 (
		_w32811_,
		_w32818_,
		_w32819_
	);
	LUT2 #(
		.INIT('h8)
	) name22308 (
		_w32816_,
		_w32817_,
		_w32820_
	);
	LUT2 #(
		.INIT('h8)
	) name22309 (
		_w32814_,
		_w32815_,
		_w32821_
	);
	LUT2 #(
		.INIT('h8)
	) name22310 (
		_w32812_,
		_w32813_,
		_w32822_
	);
	LUT2 #(
		.INIT('h8)
	) name22311 (
		_w32821_,
		_w32822_,
		_w32823_
	);
	LUT2 #(
		.INIT('h8)
	) name22312 (
		_w32819_,
		_w32820_,
		_w32824_
	);
	LUT2 #(
		.INIT('h8)
	) name22313 (
		_w32823_,
		_w32824_,
		_w32825_
	);
	LUT2 #(
		.INIT('h1)
	) name22314 (
		_w31950_,
		_w32825_,
		_w32826_
	);
	LUT2 #(
		.INIT('h1)
	) name22315 (
		_w32796_,
		_w32826_,
		_w32827_
	);
	LUT2 #(
		.INIT('h8)
	) name22316 (
		\wishbone_rx_fifo_fifo_reg[12][4]/P0001 ,
		_w31984_,
		_w32828_
	);
	LUT2 #(
		.INIT('h8)
	) name22317 (
		\wishbone_rx_fifo_fifo_reg[5][4]/P0001 ,
		_w31980_,
		_w32829_
	);
	LUT2 #(
		.INIT('h8)
	) name22318 (
		\wishbone_rx_fifo_fifo_reg[2][4]/P0001 ,
		_w31978_,
		_w32830_
	);
	LUT2 #(
		.INIT('h8)
	) name22319 (
		\wishbone_rx_fifo_fifo_reg[11][4]/P0001 ,
		_w31988_,
		_w32831_
	);
	LUT2 #(
		.INIT('h8)
	) name22320 (
		\wishbone_rx_fifo_fifo_reg[3][4]/P0001 ,
		_w31990_,
		_w32832_
	);
	LUT2 #(
		.INIT('h8)
	) name22321 (
		\wishbone_rx_fifo_fifo_reg[9][4]/P0001 ,
		_w31972_,
		_w32833_
	);
	LUT2 #(
		.INIT('h8)
	) name22322 (
		\wishbone_rx_fifo_fifo_reg[8][4]/P0001 ,
		_w31974_,
		_w32834_
	);
	LUT2 #(
		.INIT('h8)
	) name22323 (
		\wishbone_rx_fifo_fifo_reg[15][4]/P0001 ,
		_w31969_,
		_w32835_
	);
	LUT2 #(
		.INIT('h8)
	) name22324 (
		\wishbone_rx_fifo_fifo_reg[13][4]/P0001 ,
		_w31986_,
		_w32836_
	);
	LUT2 #(
		.INIT('h8)
	) name22325 (
		\wishbone_rx_fifo_fifo_reg[7][4]/P0001 ,
		_w31964_,
		_w32837_
	);
	LUT2 #(
		.INIT('h8)
	) name22326 (
		\wishbone_rx_fifo_fifo_reg[14][4]/P0001 ,
		_w31982_,
		_w32838_
	);
	LUT2 #(
		.INIT('h8)
	) name22327 (
		\wishbone_rx_fifo_fifo_reg[1][4]/P0001 ,
		_w31976_,
		_w32839_
	);
	LUT2 #(
		.INIT('h8)
	) name22328 (
		\wishbone_rx_fifo_fifo_reg[10][4]/P0001 ,
		_w31961_,
		_w32840_
	);
	LUT2 #(
		.INIT('h8)
	) name22329 (
		\wishbone_rx_fifo_fifo_reg[6][4]/P0001 ,
		_w31958_,
		_w32841_
	);
	LUT2 #(
		.INIT('h8)
	) name22330 (
		\wishbone_rx_fifo_fifo_reg[4][4]/P0001 ,
		_w31966_,
		_w32842_
	);
	LUT2 #(
		.INIT('h1)
	) name22331 (
		_w31950_,
		_w32828_,
		_w32843_
	);
	LUT2 #(
		.INIT('h1)
	) name22332 (
		_w32829_,
		_w32830_,
		_w32844_
	);
	LUT2 #(
		.INIT('h1)
	) name22333 (
		_w32831_,
		_w32832_,
		_w32845_
	);
	LUT2 #(
		.INIT('h1)
	) name22334 (
		_w32833_,
		_w32834_,
		_w32846_
	);
	LUT2 #(
		.INIT('h1)
	) name22335 (
		_w32835_,
		_w32836_,
		_w32847_
	);
	LUT2 #(
		.INIT('h1)
	) name22336 (
		_w32837_,
		_w32838_,
		_w32848_
	);
	LUT2 #(
		.INIT('h1)
	) name22337 (
		_w32839_,
		_w32840_,
		_w32849_
	);
	LUT2 #(
		.INIT('h1)
	) name22338 (
		_w32841_,
		_w32842_,
		_w32850_
	);
	LUT2 #(
		.INIT('h8)
	) name22339 (
		_w32849_,
		_w32850_,
		_w32851_
	);
	LUT2 #(
		.INIT('h8)
	) name22340 (
		_w32847_,
		_w32848_,
		_w32852_
	);
	LUT2 #(
		.INIT('h8)
	) name22341 (
		_w32845_,
		_w32846_,
		_w32853_
	);
	LUT2 #(
		.INIT('h8)
	) name22342 (
		_w32843_,
		_w32844_,
		_w32854_
	);
	LUT2 #(
		.INIT('h8)
	) name22343 (
		_w32853_,
		_w32854_,
		_w32855_
	);
	LUT2 #(
		.INIT('h8)
	) name22344 (
		_w32851_,
		_w32852_,
		_w32856_
	);
	LUT2 #(
		.INIT('h8)
	) name22345 (
		_w32855_,
		_w32856_,
		_w32857_
	);
	LUT2 #(
		.INIT('h4)
	) name22346 (
		\wishbone_rx_fifo_fifo_reg[0][4]/P0001 ,
		_w31950_,
		_w32858_
	);
	LUT2 #(
		.INIT('h1)
	) name22347 (
		_w32857_,
		_w32858_,
		_w32859_
	);
	LUT2 #(
		.INIT('h8)
	) name22348 (
		\wishbone_rx_fifo_fifo_reg[0][4]/P0001 ,
		_w31953_,
		_w32860_
	);
	LUT2 #(
		.INIT('h1)
	) name22349 (
		_w32859_,
		_w32860_,
		_w32861_
	);
	LUT2 #(
		.INIT('h8)
	) name22350 (
		\wishbone_rx_fifo_fifo_reg[10][5]/P0001 ,
		_w31961_,
		_w32862_
	);
	LUT2 #(
		.INIT('h8)
	) name22351 (
		\wishbone_rx_fifo_fifo_reg[1][5]/P0001 ,
		_w31976_,
		_w32863_
	);
	LUT2 #(
		.INIT('h8)
	) name22352 (
		\wishbone_rx_fifo_fifo_reg[8][5]/P0001 ,
		_w31974_,
		_w32864_
	);
	LUT2 #(
		.INIT('h8)
	) name22353 (
		\wishbone_rx_fifo_fifo_reg[4][5]/P0001 ,
		_w31966_,
		_w32865_
	);
	LUT2 #(
		.INIT('h8)
	) name22354 (
		\wishbone_rx_fifo_fifo_reg[13][5]/P0001 ,
		_w31986_,
		_w32866_
	);
	LUT2 #(
		.INIT('h8)
	) name22355 (
		\wishbone_rx_fifo_fifo_reg[2][5]/P0001 ,
		_w31978_,
		_w32867_
	);
	LUT2 #(
		.INIT('h8)
	) name22356 (
		\wishbone_rx_fifo_fifo_reg[12][5]/P0001 ,
		_w31984_,
		_w32868_
	);
	LUT2 #(
		.INIT('h8)
	) name22357 (
		\wishbone_rx_fifo_fifo_reg[15][5]/P0001 ,
		_w31969_,
		_w32869_
	);
	LUT2 #(
		.INIT('h8)
	) name22358 (
		\wishbone_rx_fifo_fifo_reg[3][5]/P0001 ,
		_w31990_,
		_w32870_
	);
	LUT2 #(
		.INIT('h8)
	) name22359 (
		\wishbone_rx_fifo_fifo_reg[14][5]/P0001 ,
		_w31982_,
		_w32871_
	);
	LUT2 #(
		.INIT('h8)
	) name22360 (
		\wishbone_rx_fifo_fifo_reg[11][5]/P0001 ,
		_w31988_,
		_w32872_
	);
	LUT2 #(
		.INIT('h8)
	) name22361 (
		\wishbone_rx_fifo_fifo_reg[6][5]/P0001 ,
		_w31958_,
		_w32873_
	);
	LUT2 #(
		.INIT('h8)
	) name22362 (
		\wishbone_rx_fifo_fifo_reg[7][5]/P0001 ,
		_w31964_,
		_w32874_
	);
	LUT2 #(
		.INIT('h8)
	) name22363 (
		\wishbone_rx_fifo_fifo_reg[9][5]/P0001 ,
		_w31972_,
		_w32875_
	);
	LUT2 #(
		.INIT('h8)
	) name22364 (
		\wishbone_rx_fifo_fifo_reg[5][5]/P0001 ,
		_w31980_,
		_w32876_
	);
	LUT2 #(
		.INIT('h1)
	) name22365 (
		_w31950_,
		_w32862_,
		_w32877_
	);
	LUT2 #(
		.INIT('h1)
	) name22366 (
		_w32863_,
		_w32864_,
		_w32878_
	);
	LUT2 #(
		.INIT('h1)
	) name22367 (
		_w32865_,
		_w32866_,
		_w32879_
	);
	LUT2 #(
		.INIT('h1)
	) name22368 (
		_w32867_,
		_w32868_,
		_w32880_
	);
	LUT2 #(
		.INIT('h1)
	) name22369 (
		_w32869_,
		_w32870_,
		_w32881_
	);
	LUT2 #(
		.INIT('h1)
	) name22370 (
		_w32871_,
		_w32872_,
		_w32882_
	);
	LUT2 #(
		.INIT('h1)
	) name22371 (
		_w32873_,
		_w32874_,
		_w32883_
	);
	LUT2 #(
		.INIT('h1)
	) name22372 (
		_w32875_,
		_w32876_,
		_w32884_
	);
	LUT2 #(
		.INIT('h8)
	) name22373 (
		_w32883_,
		_w32884_,
		_w32885_
	);
	LUT2 #(
		.INIT('h8)
	) name22374 (
		_w32881_,
		_w32882_,
		_w32886_
	);
	LUT2 #(
		.INIT('h8)
	) name22375 (
		_w32879_,
		_w32880_,
		_w32887_
	);
	LUT2 #(
		.INIT('h8)
	) name22376 (
		_w32877_,
		_w32878_,
		_w32888_
	);
	LUT2 #(
		.INIT('h8)
	) name22377 (
		_w32887_,
		_w32888_,
		_w32889_
	);
	LUT2 #(
		.INIT('h8)
	) name22378 (
		_w32885_,
		_w32886_,
		_w32890_
	);
	LUT2 #(
		.INIT('h8)
	) name22379 (
		_w32889_,
		_w32890_,
		_w32891_
	);
	LUT2 #(
		.INIT('h4)
	) name22380 (
		_w31953_,
		_w32891_,
		_w32892_
	);
	LUT2 #(
		.INIT('h2)
	) name22381 (
		\wishbone_rx_fifo_fifo_reg[0][5]/P0001 ,
		_w32892_,
		_w32893_
	);
	LUT2 #(
		.INIT('h1)
	) name22382 (
		_w31950_,
		_w32891_,
		_w32894_
	);
	LUT2 #(
		.INIT('h1)
	) name22383 (
		_w32893_,
		_w32894_,
		_w32895_
	);
	LUT2 #(
		.INIT('h2)
	) name22384 (
		\wishbone_rx_fifo_fifo_reg[0][6]/P0001 ,
		_w31954_,
		_w32896_
	);
	LUT2 #(
		.INIT('h8)
	) name22385 (
		\wishbone_rx_fifo_fifo_reg[5][6]/P0001 ,
		_w31980_,
		_w32897_
	);
	LUT2 #(
		.INIT('h8)
	) name22386 (
		\wishbone_rx_fifo_fifo_reg[14][6]/P0001 ,
		_w31982_,
		_w32898_
	);
	LUT2 #(
		.INIT('h8)
	) name22387 (
		\wishbone_rx_fifo_fifo_reg[12][6]/P0001 ,
		_w31984_,
		_w32899_
	);
	LUT2 #(
		.INIT('h8)
	) name22388 (
		\wishbone_rx_fifo_fifo_reg[3][6]/P0001 ,
		_w31990_,
		_w32900_
	);
	LUT2 #(
		.INIT('h8)
	) name22389 (
		\wishbone_rx_fifo_fifo_reg[9][6]/P0001 ,
		_w31972_,
		_w32901_
	);
	LUT2 #(
		.INIT('h8)
	) name22390 (
		\wishbone_rx_fifo_fifo_reg[6][6]/P0001 ,
		_w31958_,
		_w32902_
	);
	LUT2 #(
		.INIT('h8)
	) name22391 (
		\wishbone_rx_fifo_fifo_reg[2][6]/P0001 ,
		_w31978_,
		_w32903_
	);
	LUT2 #(
		.INIT('h8)
	) name22392 (
		\wishbone_rx_fifo_fifo_reg[1][6]/P0001 ,
		_w31976_,
		_w32904_
	);
	LUT2 #(
		.INIT('h8)
	) name22393 (
		\wishbone_rx_fifo_fifo_reg[4][6]/P0001 ,
		_w31966_,
		_w32905_
	);
	LUT2 #(
		.INIT('h8)
	) name22394 (
		\wishbone_rx_fifo_fifo_reg[11][6]/P0001 ,
		_w31988_,
		_w32906_
	);
	LUT2 #(
		.INIT('h8)
	) name22395 (
		\wishbone_rx_fifo_fifo_reg[15][6]/P0001 ,
		_w31969_,
		_w32907_
	);
	LUT2 #(
		.INIT('h8)
	) name22396 (
		\wishbone_rx_fifo_fifo_reg[13][6]/P0001 ,
		_w31986_,
		_w32908_
	);
	LUT2 #(
		.INIT('h8)
	) name22397 (
		\wishbone_rx_fifo_fifo_reg[10][6]/P0001 ,
		_w31961_,
		_w32909_
	);
	LUT2 #(
		.INIT('h8)
	) name22398 (
		\wishbone_rx_fifo_fifo_reg[8][6]/P0001 ,
		_w31974_,
		_w32910_
	);
	LUT2 #(
		.INIT('h8)
	) name22399 (
		\wishbone_rx_fifo_fifo_reg[7][6]/P0001 ,
		_w31964_,
		_w32911_
	);
	LUT2 #(
		.INIT('h1)
	) name22400 (
		_w32897_,
		_w32898_,
		_w32912_
	);
	LUT2 #(
		.INIT('h1)
	) name22401 (
		_w32899_,
		_w32900_,
		_w32913_
	);
	LUT2 #(
		.INIT('h1)
	) name22402 (
		_w32901_,
		_w32902_,
		_w32914_
	);
	LUT2 #(
		.INIT('h1)
	) name22403 (
		_w32903_,
		_w32904_,
		_w32915_
	);
	LUT2 #(
		.INIT('h1)
	) name22404 (
		_w32905_,
		_w32906_,
		_w32916_
	);
	LUT2 #(
		.INIT('h1)
	) name22405 (
		_w32907_,
		_w32908_,
		_w32917_
	);
	LUT2 #(
		.INIT('h1)
	) name22406 (
		_w32909_,
		_w32910_,
		_w32918_
	);
	LUT2 #(
		.INIT('h4)
	) name22407 (
		_w32911_,
		_w32918_,
		_w32919_
	);
	LUT2 #(
		.INIT('h8)
	) name22408 (
		_w32916_,
		_w32917_,
		_w32920_
	);
	LUT2 #(
		.INIT('h8)
	) name22409 (
		_w32914_,
		_w32915_,
		_w32921_
	);
	LUT2 #(
		.INIT('h8)
	) name22410 (
		_w32912_,
		_w32913_,
		_w32922_
	);
	LUT2 #(
		.INIT('h8)
	) name22411 (
		_w32921_,
		_w32922_,
		_w32923_
	);
	LUT2 #(
		.INIT('h8)
	) name22412 (
		_w32919_,
		_w32920_,
		_w32924_
	);
	LUT2 #(
		.INIT('h8)
	) name22413 (
		_w32923_,
		_w32924_,
		_w32925_
	);
	LUT2 #(
		.INIT('h1)
	) name22414 (
		_w31950_,
		_w32925_,
		_w32926_
	);
	LUT2 #(
		.INIT('h1)
	) name22415 (
		_w32896_,
		_w32926_,
		_w32927_
	);
	LUT2 #(
		.INIT('h8)
	) name22416 (
		\wishbone_rx_fifo_fifo_reg[3][7]/P0001 ,
		_w31990_,
		_w32928_
	);
	LUT2 #(
		.INIT('h8)
	) name22417 (
		\wishbone_rx_fifo_fifo_reg[2][7]/P0001 ,
		_w31978_,
		_w32929_
	);
	LUT2 #(
		.INIT('h8)
	) name22418 (
		\wishbone_rx_fifo_fifo_reg[15][7]/P0001 ,
		_w31969_,
		_w32930_
	);
	LUT2 #(
		.INIT('h8)
	) name22419 (
		\wishbone_rx_fifo_fifo_reg[13][7]/P0001 ,
		_w31986_,
		_w32931_
	);
	LUT2 #(
		.INIT('h8)
	) name22420 (
		\wishbone_rx_fifo_fifo_reg[9][7]/P0001 ,
		_w31972_,
		_w32932_
	);
	LUT2 #(
		.INIT('h8)
	) name22421 (
		\wishbone_rx_fifo_fifo_reg[6][7]/P0001 ,
		_w31958_,
		_w32933_
	);
	LUT2 #(
		.INIT('h8)
	) name22422 (
		\wishbone_rx_fifo_fifo_reg[12][7]/P0001 ,
		_w31984_,
		_w32934_
	);
	LUT2 #(
		.INIT('h8)
	) name22423 (
		\wishbone_rx_fifo_fifo_reg[14][7]/P0001 ,
		_w31982_,
		_w32935_
	);
	LUT2 #(
		.INIT('h8)
	) name22424 (
		\wishbone_rx_fifo_fifo_reg[10][7]/P0001 ,
		_w31961_,
		_w32936_
	);
	LUT2 #(
		.INIT('h8)
	) name22425 (
		\wishbone_rx_fifo_fifo_reg[1][7]/P0001 ,
		_w31976_,
		_w32937_
	);
	LUT2 #(
		.INIT('h8)
	) name22426 (
		\wishbone_rx_fifo_fifo_reg[4][7]/P0001 ,
		_w31966_,
		_w32938_
	);
	LUT2 #(
		.INIT('h8)
	) name22427 (
		\wishbone_rx_fifo_fifo_reg[8][7]/P0001 ,
		_w31974_,
		_w32939_
	);
	LUT2 #(
		.INIT('h8)
	) name22428 (
		\wishbone_rx_fifo_fifo_reg[5][7]/P0001 ,
		_w31980_,
		_w32940_
	);
	LUT2 #(
		.INIT('h8)
	) name22429 (
		\wishbone_rx_fifo_fifo_reg[11][7]/P0001 ,
		_w31988_,
		_w32941_
	);
	LUT2 #(
		.INIT('h8)
	) name22430 (
		\wishbone_rx_fifo_fifo_reg[7][7]/P0001 ,
		_w31964_,
		_w32942_
	);
	LUT2 #(
		.INIT('h1)
	) name22431 (
		_w31950_,
		_w32928_,
		_w32943_
	);
	LUT2 #(
		.INIT('h1)
	) name22432 (
		_w32929_,
		_w32930_,
		_w32944_
	);
	LUT2 #(
		.INIT('h1)
	) name22433 (
		_w32931_,
		_w32932_,
		_w32945_
	);
	LUT2 #(
		.INIT('h1)
	) name22434 (
		_w32933_,
		_w32934_,
		_w32946_
	);
	LUT2 #(
		.INIT('h1)
	) name22435 (
		_w32935_,
		_w32936_,
		_w32947_
	);
	LUT2 #(
		.INIT('h1)
	) name22436 (
		_w32937_,
		_w32938_,
		_w32948_
	);
	LUT2 #(
		.INIT('h1)
	) name22437 (
		_w32939_,
		_w32940_,
		_w32949_
	);
	LUT2 #(
		.INIT('h1)
	) name22438 (
		_w32941_,
		_w32942_,
		_w32950_
	);
	LUT2 #(
		.INIT('h8)
	) name22439 (
		_w32949_,
		_w32950_,
		_w32951_
	);
	LUT2 #(
		.INIT('h8)
	) name22440 (
		_w32947_,
		_w32948_,
		_w32952_
	);
	LUT2 #(
		.INIT('h8)
	) name22441 (
		_w32945_,
		_w32946_,
		_w32953_
	);
	LUT2 #(
		.INIT('h8)
	) name22442 (
		_w32943_,
		_w32944_,
		_w32954_
	);
	LUT2 #(
		.INIT('h8)
	) name22443 (
		_w32953_,
		_w32954_,
		_w32955_
	);
	LUT2 #(
		.INIT('h8)
	) name22444 (
		_w32951_,
		_w32952_,
		_w32956_
	);
	LUT2 #(
		.INIT('h8)
	) name22445 (
		_w32955_,
		_w32956_,
		_w32957_
	);
	LUT2 #(
		.INIT('h4)
	) name22446 (
		\wishbone_rx_fifo_fifo_reg[0][7]/P0001 ,
		_w31950_,
		_w32958_
	);
	LUT2 #(
		.INIT('h1)
	) name22447 (
		_w32957_,
		_w32958_,
		_w32959_
	);
	LUT2 #(
		.INIT('h8)
	) name22448 (
		\wishbone_rx_fifo_fifo_reg[0][7]/P0001 ,
		_w31953_,
		_w32960_
	);
	LUT2 #(
		.INIT('h1)
	) name22449 (
		_w32959_,
		_w32960_,
		_w32961_
	);
	LUT2 #(
		.INIT('h2)
	) name22450 (
		\wishbone_rx_fifo_fifo_reg[0][8]/P0001 ,
		_w31954_,
		_w32962_
	);
	LUT2 #(
		.INIT('h8)
	) name22451 (
		\wishbone_rx_fifo_fifo_reg[3][8]/P0001 ,
		_w31990_,
		_w32963_
	);
	LUT2 #(
		.INIT('h8)
	) name22452 (
		\wishbone_rx_fifo_fifo_reg[6][8]/P0001 ,
		_w31958_,
		_w32964_
	);
	LUT2 #(
		.INIT('h8)
	) name22453 (
		\wishbone_rx_fifo_fifo_reg[12][8]/P0001 ,
		_w31984_,
		_w32965_
	);
	LUT2 #(
		.INIT('h8)
	) name22454 (
		\wishbone_rx_fifo_fifo_reg[2][8]/P0001 ,
		_w31978_,
		_w32966_
	);
	LUT2 #(
		.INIT('h8)
	) name22455 (
		\wishbone_rx_fifo_fifo_reg[13][8]/P0001 ,
		_w31986_,
		_w32967_
	);
	LUT2 #(
		.INIT('h8)
	) name22456 (
		\wishbone_rx_fifo_fifo_reg[5][8]/P0001 ,
		_w31980_,
		_w32968_
	);
	LUT2 #(
		.INIT('h8)
	) name22457 (
		\wishbone_rx_fifo_fifo_reg[9][8]/P0001 ,
		_w31972_,
		_w32969_
	);
	LUT2 #(
		.INIT('h8)
	) name22458 (
		\wishbone_rx_fifo_fifo_reg[7][8]/P0001 ,
		_w31964_,
		_w32970_
	);
	LUT2 #(
		.INIT('h8)
	) name22459 (
		\wishbone_rx_fifo_fifo_reg[14][8]/P0001 ,
		_w31982_,
		_w32971_
	);
	LUT2 #(
		.INIT('h8)
	) name22460 (
		\wishbone_rx_fifo_fifo_reg[10][8]/P0001 ,
		_w31961_,
		_w32972_
	);
	LUT2 #(
		.INIT('h8)
	) name22461 (
		\wishbone_rx_fifo_fifo_reg[11][8]/P0001 ,
		_w31988_,
		_w32973_
	);
	LUT2 #(
		.INIT('h8)
	) name22462 (
		\wishbone_rx_fifo_fifo_reg[15][8]/P0001 ,
		_w31969_,
		_w32974_
	);
	LUT2 #(
		.INIT('h8)
	) name22463 (
		\wishbone_rx_fifo_fifo_reg[4][8]/P0001 ,
		_w31966_,
		_w32975_
	);
	LUT2 #(
		.INIT('h8)
	) name22464 (
		\wishbone_rx_fifo_fifo_reg[8][8]/P0001 ,
		_w31974_,
		_w32976_
	);
	LUT2 #(
		.INIT('h8)
	) name22465 (
		\wishbone_rx_fifo_fifo_reg[1][8]/P0001 ,
		_w31976_,
		_w32977_
	);
	LUT2 #(
		.INIT('h1)
	) name22466 (
		_w32963_,
		_w32964_,
		_w32978_
	);
	LUT2 #(
		.INIT('h1)
	) name22467 (
		_w32965_,
		_w32966_,
		_w32979_
	);
	LUT2 #(
		.INIT('h1)
	) name22468 (
		_w32967_,
		_w32968_,
		_w32980_
	);
	LUT2 #(
		.INIT('h1)
	) name22469 (
		_w32969_,
		_w32970_,
		_w32981_
	);
	LUT2 #(
		.INIT('h1)
	) name22470 (
		_w32971_,
		_w32972_,
		_w32982_
	);
	LUT2 #(
		.INIT('h1)
	) name22471 (
		_w32973_,
		_w32974_,
		_w32983_
	);
	LUT2 #(
		.INIT('h1)
	) name22472 (
		_w32975_,
		_w32976_,
		_w32984_
	);
	LUT2 #(
		.INIT('h4)
	) name22473 (
		_w32977_,
		_w32984_,
		_w32985_
	);
	LUT2 #(
		.INIT('h8)
	) name22474 (
		_w32982_,
		_w32983_,
		_w32986_
	);
	LUT2 #(
		.INIT('h8)
	) name22475 (
		_w32980_,
		_w32981_,
		_w32987_
	);
	LUT2 #(
		.INIT('h8)
	) name22476 (
		_w32978_,
		_w32979_,
		_w32988_
	);
	LUT2 #(
		.INIT('h8)
	) name22477 (
		_w32987_,
		_w32988_,
		_w32989_
	);
	LUT2 #(
		.INIT('h8)
	) name22478 (
		_w32985_,
		_w32986_,
		_w32990_
	);
	LUT2 #(
		.INIT('h8)
	) name22479 (
		_w32989_,
		_w32990_,
		_w32991_
	);
	LUT2 #(
		.INIT('h1)
	) name22480 (
		_w31950_,
		_w32991_,
		_w32992_
	);
	LUT2 #(
		.INIT('h1)
	) name22481 (
		_w32962_,
		_w32992_,
		_w32993_
	);
	LUT2 #(
		.INIT('h8)
	) name22482 (
		\wishbone_rx_fifo_fifo_reg[3][9]/P0001 ,
		_w31990_,
		_w32994_
	);
	LUT2 #(
		.INIT('h8)
	) name22483 (
		\wishbone_rx_fifo_fifo_reg[12][9]/P0001 ,
		_w31984_,
		_w32995_
	);
	LUT2 #(
		.INIT('h8)
	) name22484 (
		\wishbone_rx_fifo_fifo_reg[5][9]/P0001 ,
		_w31980_,
		_w32996_
	);
	LUT2 #(
		.INIT('h8)
	) name22485 (
		\wishbone_rx_fifo_fifo_reg[14][9]/P0001 ,
		_w31982_,
		_w32997_
	);
	LUT2 #(
		.INIT('h8)
	) name22486 (
		\wishbone_rx_fifo_fifo_reg[9][9]/P0001 ,
		_w31972_,
		_w32998_
	);
	LUT2 #(
		.INIT('h8)
	) name22487 (
		\wishbone_rx_fifo_fifo_reg[6][9]/P0001 ,
		_w31958_,
		_w32999_
	);
	LUT2 #(
		.INIT('h8)
	) name22488 (
		\wishbone_rx_fifo_fifo_reg[15][9]/P0001 ,
		_w31969_,
		_w33000_
	);
	LUT2 #(
		.INIT('h8)
	) name22489 (
		\wishbone_rx_fifo_fifo_reg[7][9]/P0001 ,
		_w31964_,
		_w33001_
	);
	LUT2 #(
		.INIT('h8)
	) name22490 (
		\wishbone_rx_fifo_fifo_reg[2][9]/P0001 ,
		_w31978_,
		_w33002_
	);
	LUT2 #(
		.INIT('h8)
	) name22491 (
		\wishbone_rx_fifo_fifo_reg[13][9]/P0001 ,
		_w31986_,
		_w33003_
	);
	LUT2 #(
		.INIT('h8)
	) name22492 (
		\wishbone_rx_fifo_fifo_reg[11][9]/P0001 ,
		_w31988_,
		_w33004_
	);
	LUT2 #(
		.INIT('h8)
	) name22493 (
		\wishbone_rx_fifo_fifo_reg[1][9]/P0001 ,
		_w31976_,
		_w33005_
	);
	LUT2 #(
		.INIT('h8)
	) name22494 (
		\wishbone_rx_fifo_fifo_reg[10][9]/P0001 ,
		_w31961_,
		_w33006_
	);
	LUT2 #(
		.INIT('h8)
	) name22495 (
		\wishbone_rx_fifo_fifo_reg[8][9]/P0001 ,
		_w31974_,
		_w33007_
	);
	LUT2 #(
		.INIT('h8)
	) name22496 (
		\wishbone_rx_fifo_fifo_reg[4][9]/P0001 ,
		_w31966_,
		_w33008_
	);
	LUT2 #(
		.INIT('h1)
	) name22497 (
		_w31950_,
		_w32994_,
		_w33009_
	);
	LUT2 #(
		.INIT('h1)
	) name22498 (
		_w32995_,
		_w32996_,
		_w33010_
	);
	LUT2 #(
		.INIT('h1)
	) name22499 (
		_w32997_,
		_w32998_,
		_w33011_
	);
	LUT2 #(
		.INIT('h1)
	) name22500 (
		_w32999_,
		_w33000_,
		_w33012_
	);
	LUT2 #(
		.INIT('h1)
	) name22501 (
		_w33001_,
		_w33002_,
		_w33013_
	);
	LUT2 #(
		.INIT('h1)
	) name22502 (
		_w33003_,
		_w33004_,
		_w33014_
	);
	LUT2 #(
		.INIT('h1)
	) name22503 (
		_w33005_,
		_w33006_,
		_w33015_
	);
	LUT2 #(
		.INIT('h1)
	) name22504 (
		_w33007_,
		_w33008_,
		_w33016_
	);
	LUT2 #(
		.INIT('h8)
	) name22505 (
		_w33015_,
		_w33016_,
		_w33017_
	);
	LUT2 #(
		.INIT('h8)
	) name22506 (
		_w33013_,
		_w33014_,
		_w33018_
	);
	LUT2 #(
		.INIT('h8)
	) name22507 (
		_w33011_,
		_w33012_,
		_w33019_
	);
	LUT2 #(
		.INIT('h8)
	) name22508 (
		_w33009_,
		_w33010_,
		_w33020_
	);
	LUT2 #(
		.INIT('h8)
	) name22509 (
		_w33019_,
		_w33020_,
		_w33021_
	);
	LUT2 #(
		.INIT('h8)
	) name22510 (
		_w33017_,
		_w33018_,
		_w33022_
	);
	LUT2 #(
		.INIT('h8)
	) name22511 (
		_w33021_,
		_w33022_,
		_w33023_
	);
	LUT2 #(
		.INIT('h4)
	) name22512 (
		\wishbone_rx_fifo_fifo_reg[0][9]/P0001 ,
		_w31950_,
		_w33024_
	);
	LUT2 #(
		.INIT('h1)
	) name22513 (
		_w33023_,
		_w33024_,
		_w33025_
	);
	LUT2 #(
		.INIT('h8)
	) name22514 (
		\wishbone_rx_fifo_fifo_reg[0][9]/P0001 ,
		_w31953_,
		_w33026_
	);
	LUT2 #(
		.INIT('h1)
	) name22515 (
		_w33025_,
		_w33026_,
		_w33027_
	);
	LUT2 #(
		.INIT('h1)
	) name22516 (
		\wishbone_TxAbortPacket_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w33028_
	);
	LUT2 #(
		.INIT('h1)
	) name22517 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w33029_
	);
	LUT2 #(
		.INIT('h1)
	) name22518 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w33030_
	);
	LUT2 #(
		.INIT('h8)
	) name22519 (
		_w33029_,
		_w33030_,
		_w33031_
	);
	LUT2 #(
		.INIT('h2)
	) name22520 (
		_w33028_,
		_w33031_,
		_w33032_
	);
	LUT2 #(
		.INIT('h2)
	) name22521 (
		\wishbone_tx_fifo_fifo_reg[0][0]/P0001 ,
		_w33032_,
		_w33033_
	);
	LUT2 #(
		.INIT('h8)
	) name22522 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w33034_
	);
	LUT2 #(
		.INIT('h4)
	) name22523 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w33035_
	);
	LUT2 #(
		.INIT('h8)
	) name22524 (
		_w33034_,
		_w33035_,
		_w33036_
	);
	LUT2 #(
		.INIT('h8)
	) name22525 (
		\wishbone_tx_fifo_fifo_reg[11][0]/P0001 ,
		_w33036_,
		_w33037_
	);
	LUT2 #(
		.INIT('h2)
	) name22526 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w33038_
	);
	LUT2 #(
		.INIT('h2)
	) name22527 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w33039_
	);
	LUT2 #(
		.INIT('h8)
	) name22528 (
		_w33038_,
		_w33039_,
		_w33040_
	);
	LUT2 #(
		.INIT('h8)
	) name22529 (
		\wishbone_tx_fifo_fifo_reg[5][0]/P0001 ,
		_w33040_,
		_w33041_
	);
	LUT2 #(
		.INIT('h8)
	) name22530 (
		_w33029_,
		_w33035_,
		_w33042_
	);
	LUT2 #(
		.INIT('h8)
	) name22531 (
		\wishbone_tx_fifo_fifo_reg[8][0]/P0001 ,
		_w33042_,
		_w33043_
	);
	LUT2 #(
		.INIT('h8)
	) name22532 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w33044_
	);
	LUT2 #(
		.INIT('h8)
	) name22533 (
		_w33034_,
		_w33044_,
		_w33045_
	);
	LUT2 #(
		.INIT('h8)
	) name22534 (
		\wishbone_tx_fifo_fifo_reg[15][0]/P0001 ,
		_w33045_,
		_w33046_
	);
	LUT2 #(
		.INIT('h8)
	) name22535 (
		_w33039_,
		_w33044_,
		_w33047_
	);
	LUT2 #(
		.INIT('h8)
	) name22536 (
		\wishbone_tx_fifo_fifo_reg[13][0]/P0001 ,
		_w33047_,
		_w33048_
	);
	LUT2 #(
		.INIT('h4)
	) name22537 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w33049_
	);
	LUT2 #(
		.INIT('h8)
	) name22538 (
		_w33044_,
		_w33049_,
		_w33050_
	);
	LUT2 #(
		.INIT('h8)
	) name22539 (
		\wishbone_tx_fifo_fifo_reg[14][0]/P0001 ,
		_w33050_,
		_w33051_
	);
	LUT2 #(
		.INIT('h8)
	) name22540 (
		_w33035_,
		_w33039_,
		_w33052_
	);
	LUT2 #(
		.INIT('h8)
	) name22541 (
		\wishbone_tx_fifo_fifo_reg[9][0]/P0001 ,
		_w33052_,
		_w33053_
	);
	LUT2 #(
		.INIT('h8)
	) name22542 (
		_w33034_,
		_w33038_,
		_w33054_
	);
	LUT2 #(
		.INIT('h8)
	) name22543 (
		\wishbone_tx_fifo_fifo_reg[7][0]/P0001 ,
		_w33054_,
		_w33055_
	);
	LUT2 #(
		.INIT('h8)
	) name22544 (
		_w33038_,
		_w33049_,
		_w33056_
	);
	LUT2 #(
		.INIT('h8)
	) name22545 (
		\wishbone_tx_fifo_fifo_reg[6][0]/P0001 ,
		_w33056_,
		_w33057_
	);
	LUT2 #(
		.INIT('h8)
	) name22546 (
		_w33029_,
		_w33044_,
		_w33058_
	);
	LUT2 #(
		.INIT('h8)
	) name22547 (
		\wishbone_tx_fifo_fifo_reg[12][0]/P0001 ,
		_w33058_,
		_w33059_
	);
	LUT2 #(
		.INIT('h8)
	) name22548 (
		_w33030_,
		_w33039_,
		_w33060_
	);
	LUT2 #(
		.INIT('h8)
	) name22549 (
		\wishbone_tx_fifo_fifo_reg[1][0]/P0001 ,
		_w33060_,
		_w33061_
	);
	LUT2 #(
		.INIT('h8)
	) name22550 (
		_w33030_,
		_w33034_,
		_w33062_
	);
	LUT2 #(
		.INIT('h8)
	) name22551 (
		\wishbone_tx_fifo_fifo_reg[3][0]/P0001 ,
		_w33062_,
		_w33063_
	);
	LUT2 #(
		.INIT('h8)
	) name22552 (
		_w33029_,
		_w33038_,
		_w33064_
	);
	LUT2 #(
		.INIT('h8)
	) name22553 (
		\wishbone_tx_fifo_fifo_reg[4][0]/P0001 ,
		_w33064_,
		_w33065_
	);
	LUT2 #(
		.INIT('h8)
	) name22554 (
		_w33035_,
		_w33049_,
		_w33066_
	);
	LUT2 #(
		.INIT('h8)
	) name22555 (
		\wishbone_tx_fifo_fifo_reg[10][0]/P0001 ,
		_w33066_,
		_w33067_
	);
	LUT2 #(
		.INIT('h8)
	) name22556 (
		_w33030_,
		_w33049_,
		_w33068_
	);
	LUT2 #(
		.INIT('h8)
	) name22557 (
		\wishbone_tx_fifo_fifo_reg[2][0]/P0001 ,
		_w33068_,
		_w33069_
	);
	LUT2 #(
		.INIT('h1)
	) name22558 (
		_w33037_,
		_w33041_,
		_w33070_
	);
	LUT2 #(
		.INIT('h1)
	) name22559 (
		_w33043_,
		_w33046_,
		_w33071_
	);
	LUT2 #(
		.INIT('h1)
	) name22560 (
		_w33048_,
		_w33051_,
		_w33072_
	);
	LUT2 #(
		.INIT('h1)
	) name22561 (
		_w33053_,
		_w33055_,
		_w33073_
	);
	LUT2 #(
		.INIT('h1)
	) name22562 (
		_w33057_,
		_w33059_,
		_w33074_
	);
	LUT2 #(
		.INIT('h1)
	) name22563 (
		_w33061_,
		_w33063_,
		_w33075_
	);
	LUT2 #(
		.INIT('h1)
	) name22564 (
		_w33065_,
		_w33067_,
		_w33076_
	);
	LUT2 #(
		.INIT('h4)
	) name22565 (
		_w33069_,
		_w33076_,
		_w33077_
	);
	LUT2 #(
		.INIT('h8)
	) name22566 (
		_w33074_,
		_w33075_,
		_w33078_
	);
	LUT2 #(
		.INIT('h8)
	) name22567 (
		_w33072_,
		_w33073_,
		_w33079_
	);
	LUT2 #(
		.INIT('h8)
	) name22568 (
		_w33070_,
		_w33071_,
		_w33080_
	);
	LUT2 #(
		.INIT('h8)
	) name22569 (
		_w33079_,
		_w33080_,
		_w33081_
	);
	LUT2 #(
		.INIT('h8)
	) name22570 (
		_w33077_,
		_w33078_,
		_w33082_
	);
	LUT2 #(
		.INIT('h8)
	) name22571 (
		_w33081_,
		_w33082_,
		_w33083_
	);
	LUT2 #(
		.INIT('h2)
	) name22572 (
		_w33028_,
		_w33083_,
		_w33084_
	);
	LUT2 #(
		.INIT('h1)
	) name22573 (
		_w33033_,
		_w33084_,
		_w33085_
	);
	LUT2 #(
		.INIT('h2)
	) name22574 (
		\wishbone_tx_fifo_fifo_reg[0][10]/P0001 ,
		_w33032_,
		_w33086_
	);
	LUT2 #(
		.INIT('h8)
	) name22575 (
		\wishbone_tx_fifo_fifo_reg[2][10]/P0001 ,
		_w33068_,
		_w33087_
	);
	LUT2 #(
		.INIT('h8)
	) name22576 (
		\wishbone_tx_fifo_fifo_reg[13][10]/P0001 ,
		_w33047_,
		_w33088_
	);
	LUT2 #(
		.INIT('h8)
	) name22577 (
		\wishbone_tx_fifo_fifo_reg[5][10]/P0001 ,
		_w33040_,
		_w33089_
	);
	LUT2 #(
		.INIT('h8)
	) name22578 (
		\wishbone_tx_fifo_fifo_reg[11][10]/P0001 ,
		_w33036_,
		_w33090_
	);
	LUT2 #(
		.INIT('h8)
	) name22579 (
		\wishbone_tx_fifo_fifo_reg[3][10]/P0001 ,
		_w33062_,
		_w33091_
	);
	LUT2 #(
		.INIT('h8)
	) name22580 (
		\wishbone_tx_fifo_fifo_reg[7][10]/P0001 ,
		_w33054_,
		_w33092_
	);
	LUT2 #(
		.INIT('h8)
	) name22581 (
		\wishbone_tx_fifo_fifo_reg[15][10]/P0001 ,
		_w33045_,
		_w33093_
	);
	LUT2 #(
		.INIT('h8)
	) name22582 (
		\wishbone_tx_fifo_fifo_reg[14][10]/P0001 ,
		_w33050_,
		_w33094_
	);
	LUT2 #(
		.INIT('h8)
	) name22583 (
		\wishbone_tx_fifo_fifo_reg[12][10]/P0001 ,
		_w33058_,
		_w33095_
	);
	LUT2 #(
		.INIT('h8)
	) name22584 (
		\wishbone_tx_fifo_fifo_reg[4][10]/P0001 ,
		_w33064_,
		_w33096_
	);
	LUT2 #(
		.INIT('h8)
	) name22585 (
		\wishbone_tx_fifo_fifo_reg[1][10]/P0001 ,
		_w33060_,
		_w33097_
	);
	LUT2 #(
		.INIT('h8)
	) name22586 (
		\wishbone_tx_fifo_fifo_reg[9][10]/P0001 ,
		_w33052_,
		_w33098_
	);
	LUT2 #(
		.INIT('h8)
	) name22587 (
		\wishbone_tx_fifo_fifo_reg[10][10]/P0001 ,
		_w33066_,
		_w33099_
	);
	LUT2 #(
		.INIT('h8)
	) name22588 (
		\wishbone_tx_fifo_fifo_reg[6][10]/P0001 ,
		_w33056_,
		_w33100_
	);
	LUT2 #(
		.INIT('h8)
	) name22589 (
		\wishbone_tx_fifo_fifo_reg[8][10]/P0001 ,
		_w33042_,
		_w33101_
	);
	LUT2 #(
		.INIT('h1)
	) name22590 (
		_w33087_,
		_w33088_,
		_w33102_
	);
	LUT2 #(
		.INIT('h1)
	) name22591 (
		_w33089_,
		_w33090_,
		_w33103_
	);
	LUT2 #(
		.INIT('h1)
	) name22592 (
		_w33091_,
		_w33092_,
		_w33104_
	);
	LUT2 #(
		.INIT('h1)
	) name22593 (
		_w33093_,
		_w33094_,
		_w33105_
	);
	LUT2 #(
		.INIT('h1)
	) name22594 (
		_w33095_,
		_w33096_,
		_w33106_
	);
	LUT2 #(
		.INIT('h1)
	) name22595 (
		_w33097_,
		_w33098_,
		_w33107_
	);
	LUT2 #(
		.INIT('h1)
	) name22596 (
		_w33099_,
		_w33100_,
		_w33108_
	);
	LUT2 #(
		.INIT('h4)
	) name22597 (
		_w33101_,
		_w33108_,
		_w33109_
	);
	LUT2 #(
		.INIT('h8)
	) name22598 (
		_w33106_,
		_w33107_,
		_w33110_
	);
	LUT2 #(
		.INIT('h8)
	) name22599 (
		_w33104_,
		_w33105_,
		_w33111_
	);
	LUT2 #(
		.INIT('h8)
	) name22600 (
		_w33102_,
		_w33103_,
		_w33112_
	);
	LUT2 #(
		.INIT('h8)
	) name22601 (
		_w33111_,
		_w33112_,
		_w33113_
	);
	LUT2 #(
		.INIT('h8)
	) name22602 (
		_w33109_,
		_w33110_,
		_w33114_
	);
	LUT2 #(
		.INIT('h8)
	) name22603 (
		_w33113_,
		_w33114_,
		_w33115_
	);
	LUT2 #(
		.INIT('h2)
	) name22604 (
		_w33028_,
		_w33115_,
		_w33116_
	);
	LUT2 #(
		.INIT('h1)
	) name22605 (
		_w33086_,
		_w33116_,
		_w33117_
	);
	LUT2 #(
		.INIT('h2)
	) name22606 (
		\wishbone_tx_fifo_fifo_reg[0][11]/P0001 ,
		_w33032_,
		_w33118_
	);
	LUT2 #(
		.INIT('h8)
	) name22607 (
		\wishbone_tx_fifo_fifo_reg[3][11]/P0001 ,
		_w33062_,
		_w33119_
	);
	LUT2 #(
		.INIT('h8)
	) name22608 (
		\wishbone_tx_fifo_fifo_reg[6][11]/P0001 ,
		_w33056_,
		_w33120_
	);
	LUT2 #(
		.INIT('h8)
	) name22609 (
		\wishbone_tx_fifo_fifo_reg[8][11]/P0001 ,
		_w33042_,
		_w33121_
	);
	LUT2 #(
		.INIT('h8)
	) name22610 (
		\wishbone_tx_fifo_fifo_reg[7][11]/P0001 ,
		_w33054_,
		_w33122_
	);
	LUT2 #(
		.INIT('h8)
	) name22611 (
		\wishbone_tx_fifo_fifo_reg[10][11]/P0001 ,
		_w33066_,
		_w33123_
	);
	LUT2 #(
		.INIT('h8)
	) name22612 (
		\wishbone_tx_fifo_fifo_reg[5][11]/P0001 ,
		_w33040_,
		_w33124_
	);
	LUT2 #(
		.INIT('h8)
	) name22613 (
		\wishbone_tx_fifo_fifo_reg[14][11]/P0001 ,
		_w33050_,
		_w33125_
	);
	LUT2 #(
		.INIT('h8)
	) name22614 (
		\wishbone_tx_fifo_fifo_reg[4][11]/P0001 ,
		_w33064_,
		_w33126_
	);
	LUT2 #(
		.INIT('h8)
	) name22615 (
		\wishbone_tx_fifo_fifo_reg[1][11]/P0001 ,
		_w33060_,
		_w33127_
	);
	LUT2 #(
		.INIT('h8)
	) name22616 (
		\wishbone_tx_fifo_fifo_reg[13][11]/P0001 ,
		_w33047_,
		_w33128_
	);
	LUT2 #(
		.INIT('h8)
	) name22617 (
		\wishbone_tx_fifo_fifo_reg[2][11]/P0001 ,
		_w33068_,
		_w33129_
	);
	LUT2 #(
		.INIT('h8)
	) name22618 (
		\wishbone_tx_fifo_fifo_reg[12][11]/P0001 ,
		_w33058_,
		_w33130_
	);
	LUT2 #(
		.INIT('h8)
	) name22619 (
		\wishbone_tx_fifo_fifo_reg[15][11]/P0001 ,
		_w33045_,
		_w33131_
	);
	LUT2 #(
		.INIT('h8)
	) name22620 (
		\wishbone_tx_fifo_fifo_reg[11][11]/P0001 ,
		_w33036_,
		_w33132_
	);
	LUT2 #(
		.INIT('h8)
	) name22621 (
		\wishbone_tx_fifo_fifo_reg[9][11]/P0001 ,
		_w33052_,
		_w33133_
	);
	LUT2 #(
		.INIT('h1)
	) name22622 (
		_w33119_,
		_w33120_,
		_w33134_
	);
	LUT2 #(
		.INIT('h1)
	) name22623 (
		_w33121_,
		_w33122_,
		_w33135_
	);
	LUT2 #(
		.INIT('h1)
	) name22624 (
		_w33123_,
		_w33124_,
		_w33136_
	);
	LUT2 #(
		.INIT('h1)
	) name22625 (
		_w33125_,
		_w33126_,
		_w33137_
	);
	LUT2 #(
		.INIT('h1)
	) name22626 (
		_w33127_,
		_w33128_,
		_w33138_
	);
	LUT2 #(
		.INIT('h1)
	) name22627 (
		_w33129_,
		_w33130_,
		_w33139_
	);
	LUT2 #(
		.INIT('h1)
	) name22628 (
		_w33131_,
		_w33132_,
		_w33140_
	);
	LUT2 #(
		.INIT('h4)
	) name22629 (
		_w33133_,
		_w33140_,
		_w33141_
	);
	LUT2 #(
		.INIT('h8)
	) name22630 (
		_w33138_,
		_w33139_,
		_w33142_
	);
	LUT2 #(
		.INIT('h8)
	) name22631 (
		_w33136_,
		_w33137_,
		_w33143_
	);
	LUT2 #(
		.INIT('h8)
	) name22632 (
		_w33134_,
		_w33135_,
		_w33144_
	);
	LUT2 #(
		.INIT('h8)
	) name22633 (
		_w33143_,
		_w33144_,
		_w33145_
	);
	LUT2 #(
		.INIT('h8)
	) name22634 (
		_w33141_,
		_w33142_,
		_w33146_
	);
	LUT2 #(
		.INIT('h8)
	) name22635 (
		_w33145_,
		_w33146_,
		_w33147_
	);
	LUT2 #(
		.INIT('h2)
	) name22636 (
		_w33028_,
		_w33147_,
		_w33148_
	);
	LUT2 #(
		.INIT('h1)
	) name22637 (
		_w33118_,
		_w33148_,
		_w33149_
	);
	LUT2 #(
		.INIT('h2)
	) name22638 (
		\wishbone_tx_fifo_fifo_reg[0][12]/P0001 ,
		_w33032_,
		_w33150_
	);
	LUT2 #(
		.INIT('h8)
	) name22639 (
		\wishbone_tx_fifo_fifo_reg[6][12]/P0001 ,
		_w33056_,
		_w33151_
	);
	LUT2 #(
		.INIT('h8)
	) name22640 (
		\wishbone_tx_fifo_fifo_reg[12][12]/P0001 ,
		_w33058_,
		_w33152_
	);
	LUT2 #(
		.INIT('h8)
	) name22641 (
		\wishbone_tx_fifo_fifo_reg[8][12]/P0001 ,
		_w33042_,
		_w33153_
	);
	LUT2 #(
		.INIT('h8)
	) name22642 (
		\wishbone_tx_fifo_fifo_reg[11][12]/P0001 ,
		_w33036_,
		_w33154_
	);
	LUT2 #(
		.INIT('h8)
	) name22643 (
		\wishbone_tx_fifo_fifo_reg[5][12]/P0001 ,
		_w33040_,
		_w33155_
	);
	LUT2 #(
		.INIT('h8)
	) name22644 (
		\wishbone_tx_fifo_fifo_reg[9][12]/P0001 ,
		_w33052_,
		_w33156_
	);
	LUT2 #(
		.INIT('h8)
	) name22645 (
		\wishbone_tx_fifo_fifo_reg[10][12]/P0001 ,
		_w33066_,
		_w33157_
	);
	LUT2 #(
		.INIT('h8)
	) name22646 (
		\wishbone_tx_fifo_fifo_reg[13][12]/P0001 ,
		_w33047_,
		_w33158_
	);
	LUT2 #(
		.INIT('h8)
	) name22647 (
		\wishbone_tx_fifo_fifo_reg[1][12]/P0001 ,
		_w33060_,
		_w33159_
	);
	LUT2 #(
		.INIT('h8)
	) name22648 (
		\wishbone_tx_fifo_fifo_reg[15][12]/P0001 ,
		_w33045_,
		_w33160_
	);
	LUT2 #(
		.INIT('h8)
	) name22649 (
		\wishbone_tx_fifo_fifo_reg[4][12]/P0001 ,
		_w33064_,
		_w33161_
	);
	LUT2 #(
		.INIT('h8)
	) name22650 (
		\wishbone_tx_fifo_fifo_reg[3][12]/P0001 ,
		_w33062_,
		_w33162_
	);
	LUT2 #(
		.INIT('h8)
	) name22651 (
		\wishbone_tx_fifo_fifo_reg[7][12]/P0001 ,
		_w33054_,
		_w33163_
	);
	LUT2 #(
		.INIT('h8)
	) name22652 (
		\wishbone_tx_fifo_fifo_reg[14][12]/P0001 ,
		_w33050_,
		_w33164_
	);
	LUT2 #(
		.INIT('h8)
	) name22653 (
		\wishbone_tx_fifo_fifo_reg[2][12]/P0001 ,
		_w33068_,
		_w33165_
	);
	LUT2 #(
		.INIT('h1)
	) name22654 (
		_w33151_,
		_w33152_,
		_w33166_
	);
	LUT2 #(
		.INIT('h1)
	) name22655 (
		_w33153_,
		_w33154_,
		_w33167_
	);
	LUT2 #(
		.INIT('h1)
	) name22656 (
		_w33155_,
		_w33156_,
		_w33168_
	);
	LUT2 #(
		.INIT('h1)
	) name22657 (
		_w33157_,
		_w33158_,
		_w33169_
	);
	LUT2 #(
		.INIT('h1)
	) name22658 (
		_w33159_,
		_w33160_,
		_w33170_
	);
	LUT2 #(
		.INIT('h1)
	) name22659 (
		_w33161_,
		_w33162_,
		_w33171_
	);
	LUT2 #(
		.INIT('h1)
	) name22660 (
		_w33163_,
		_w33164_,
		_w33172_
	);
	LUT2 #(
		.INIT('h4)
	) name22661 (
		_w33165_,
		_w33172_,
		_w33173_
	);
	LUT2 #(
		.INIT('h8)
	) name22662 (
		_w33170_,
		_w33171_,
		_w33174_
	);
	LUT2 #(
		.INIT('h8)
	) name22663 (
		_w33168_,
		_w33169_,
		_w33175_
	);
	LUT2 #(
		.INIT('h8)
	) name22664 (
		_w33166_,
		_w33167_,
		_w33176_
	);
	LUT2 #(
		.INIT('h8)
	) name22665 (
		_w33175_,
		_w33176_,
		_w33177_
	);
	LUT2 #(
		.INIT('h8)
	) name22666 (
		_w33173_,
		_w33174_,
		_w33178_
	);
	LUT2 #(
		.INIT('h8)
	) name22667 (
		_w33177_,
		_w33178_,
		_w33179_
	);
	LUT2 #(
		.INIT('h2)
	) name22668 (
		_w33028_,
		_w33179_,
		_w33180_
	);
	LUT2 #(
		.INIT('h1)
	) name22669 (
		_w33150_,
		_w33180_,
		_w33181_
	);
	LUT2 #(
		.INIT('h2)
	) name22670 (
		\wishbone_tx_fifo_fifo_reg[0][13]/P0001 ,
		_w33032_,
		_w33182_
	);
	LUT2 #(
		.INIT('h8)
	) name22671 (
		\wishbone_tx_fifo_fifo_reg[3][13]/P0001 ,
		_w33062_,
		_w33183_
	);
	LUT2 #(
		.INIT('h8)
	) name22672 (
		\wishbone_tx_fifo_fifo_reg[5][13]/P0001 ,
		_w33040_,
		_w33184_
	);
	LUT2 #(
		.INIT('h8)
	) name22673 (
		\wishbone_tx_fifo_fifo_reg[15][13]/P0001 ,
		_w33045_,
		_w33185_
	);
	LUT2 #(
		.INIT('h8)
	) name22674 (
		\wishbone_tx_fifo_fifo_reg[2][13]/P0001 ,
		_w33068_,
		_w33186_
	);
	LUT2 #(
		.INIT('h8)
	) name22675 (
		\wishbone_tx_fifo_fifo_reg[13][13]/P0001 ,
		_w33047_,
		_w33187_
	);
	LUT2 #(
		.INIT('h8)
	) name22676 (
		\wishbone_tx_fifo_fifo_reg[9][13]/P0001 ,
		_w33052_,
		_w33188_
	);
	LUT2 #(
		.INIT('h8)
	) name22677 (
		\wishbone_tx_fifo_fifo_reg[8][13]/P0001 ,
		_w33042_,
		_w33189_
	);
	LUT2 #(
		.INIT('h8)
	) name22678 (
		\wishbone_tx_fifo_fifo_reg[14][13]/P0001 ,
		_w33050_,
		_w33190_
	);
	LUT2 #(
		.INIT('h8)
	) name22679 (
		\wishbone_tx_fifo_fifo_reg[7][13]/P0001 ,
		_w33054_,
		_w33191_
	);
	LUT2 #(
		.INIT('h8)
	) name22680 (
		\wishbone_tx_fifo_fifo_reg[10][13]/P0001 ,
		_w33066_,
		_w33192_
	);
	LUT2 #(
		.INIT('h8)
	) name22681 (
		\wishbone_tx_fifo_fifo_reg[11][13]/P0001 ,
		_w33036_,
		_w33193_
	);
	LUT2 #(
		.INIT('h8)
	) name22682 (
		\wishbone_tx_fifo_fifo_reg[12][13]/P0001 ,
		_w33058_,
		_w33194_
	);
	LUT2 #(
		.INIT('h8)
	) name22683 (
		\wishbone_tx_fifo_fifo_reg[4][13]/P0001 ,
		_w33064_,
		_w33195_
	);
	LUT2 #(
		.INIT('h8)
	) name22684 (
		\wishbone_tx_fifo_fifo_reg[6][13]/P0001 ,
		_w33056_,
		_w33196_
	);
	LUT2 #(
		.INIT('h8)
	) name22685 (
		\wishbone_tx_fifo_fifo_reg[1][13]/P0001 ,
		_w33060_,
		_w33197_
	);
	LUT2 #(
		.INIT('h1)
	) name22686 (
		_w33183_,
		_w33184_,
		_w33198_
	);
	LUT2 #(
		.INIT('h1)
	) name22687 (
		_w33185_,
		_w33186_,
		_w33199_
	);
	LUT2 #(
		.INIT('h1)
	) name22688 (
		_w33187_,
		_w33188_,
		_w33200_
	);
	LUT2 #(
		.INIT('h1)
	) name22689 (
		_w33189_,
		_w33190_,
		_w33201_
	);
	LUT2 #(
		.INIT('h1)
	) name22690 (
		_w33191_,
		_w33192_,
		_w33202_
	);
	LUT2 #(
		.INIT('h1)
	) name22691 (
		_w33193_,
		_w33194_,
		_w33203_
	);
	LUT2 #(
		.INIT('h1)
	) name22692 (
		_w33195_,
		_w33196_,
		_w33204_
	);
	LUT2 #(
		.INIT('h4)
	) name22693 (
		_w33197_,
		_w33204_,
		_w33205_
	);
	LUT2 #(
		.INIT('h8)
	) name22694 (
		_w33202_,
		_w33203_,
		_w33206_
	);
	LUT2 #(
		.INIT('h8)
	) name22695 (
		_w33200_,
		_w33201_,
		_w33207_
	);
	LUT2 #(
		.INIT('h8)
	) name22696 (
		_w33198_,
		_w33199_,
		_w33208_
	);
	LUT2 #(
		.INIT('h8)
	) name22697 (
		_w33207_,
		_w33208_,
		_w33209_
	);
	LUT2 #(
		.INIT('h8)
	) name22698 (
		_w33205_,
		_w33206_,
		_w33210_
	);
	LUT2 #(
		.INIT('h8)
	) name22699 (
		_w33209_,
		_w33210_,
		_w33211_
	);
	LUT2 #(
		.INIT('h2)
	) name22700 (
		_w33028_,
		_w33211_,
		_w33212_
	);
	LUT2 #(
		.INIT('h1)
	) name22701 (
		_w33182_,
		_w33212_,
		_w33213_
	);
	LUT2 #(
		.INIT('h2)
	) name22702 (
		\wishbone_tx_fifo_fifo_reg[0][14]/P0001 ,
		_w33032_,
		_w33214_
	);
	LUT2 #(
		.INIT('h8)
	) name22703 (
		\wishbone_tx_fifo_fifo_reg[10][14]/P0001 ,
		_w33066_,
		_w33215_
	);
	LUT2 #(
		.INIT('h8)
	) name22704 (
		\wishbone_tx_fifo_fifo_reg[9][14]/P0001 ,
		_w33052_,
		_w33216_
	);
	LUT2 #(
		.INIT('h8)
	) name22705 (
		\wishbone_tx_fifo_fifo_reg[12][14]/P0001 ,
		_w33058_,
		_w33217_
	);
	LUT2 #(
		.INIT('h8)
	) name22706 (
		\wishbone_tx_fifo_fifo_reg[8][14]/P0001 ,
		_w33042_,
		_w33218_
	);
	LUT2 #(
		.INIT('h8)
	) name22707 (
		\wishbone_tx_fifo_fifo_reg[15][14]/P0001 ,
		_w33045_,
		_w33219_
	);
	LUT2 #(
		.INIT('h8)
	) name22708 (
		\wishbone_tx_fifo_fifo_reg[6][14]/P0001 ,
		_w33056_,
		_w33220_
	);
	LUT2 #(
		.INIT('h8)
	) name22709 (
		\wishbone_tx_fifo_fifo_reg[3][14]/P0001 ,
		_w33062_,
		_w33221_
	);
	LUT2 #(
		.INIT('h8)
	) name22710 (
		\wishbone_tx_fifo_fifo_reg[11][14]/P0001 ,
		_w33036_,
		_w33222_
	);
	LUT2 #(
		.INIT('h8)
	) name22711 (
		\wishbone_tx_fifo_fifo_reg[5][14]/P0001 ,
		_w33040_,
		_w33223_
	);
	LUT2 #(
		.INIT('h8)
	) name22712 (
		\wishbone_tx_fifo_fifo_reg[14][14]/P0001 ,
		_w33050_,
		_w33224_
	);
	LUT2 #(
		.INIT('h8)
	) name22713 (
		\wishbone_tx_fifo_fifo_reg[7][14]/P0001 ,
		_w33054_,
		_w33225_
	);
	LUT2 #(
		.INIT('h8)
	) name22714 (
		\wishbone_tx_fifo_fifo_reg[13][14]/P0001 ,
		_w33047_,
		_w33226_
	);
	LUT2 #(
		.INIT('h8)
	) name22715 (
		\wishbone_tx_fifo_fifo_reg[4][14]/P0001 ,
		_w33064_,
		_w33227_
	);
	LUT2 #(
		.INIT('h8)
	) name22716 (
		\wishbone_tx_fifo_fifo_reg[1][14]/P0001 ,
		_w33060_,
		_w33228_
	);
	LUT2 #(
		.INIT('h8)
	) name22717 (
		\wishbone_tx_fifo_fifo_reg[2][14]/P0001 ,
		_w33068_,
		_w33229_
	);
	LUT2 #(
		.INIT('h1)
	) name22718 (
		_w33215_,
		_w33216_,
		_w33230_
	);
	LUT2 #(
		.INIT('h1)
	) name22719 (
		_w33217_,
		_w33218_,
		_w33231_
	);
	LUT2 #(
		.INIT('h1)
	) name22720 (
		_w33219_,
		_w33220_,
		_w33232_
	);
	LUT2 #(
		.INIT('h1)
	) name22721 (
		_w33221_,
		_w33222_,
		_w33233_
	);
	LUT2 #(
		.INIT('h1)
	) name22722 (
		_w33223_,
		_w33224_,
		_w33234_
	);
	LUT2 #(
		.INIT('h1)
	) name22723 (
		_w33225_,
		_w33226_,
		_w33235_
	);
	LUT2 #(
		.INIT('h1)
	) name22724 (
		_w33227_,
		_w33228_,
		_w33236_
	);
	LUT2 #(
		.INIT('h4)
	) name22725 (
		_w33229_,
		_w33236_,
		_w33237_
	);
	LUT2 #(
		.INIT('h8)
	) name22726 (
		_w33234_,
		_w33235_,
		_w33238_
	);
	LUT2 #(
		.INIT('h8)
	) name22727 (
		_w33232_,
		_w33233_,
		_w33239_
	);
	LUT2 #(
		.INIT('h8)
	) name22728 (
		_w33230_,
		_w33231_,
		_w33240_
	);
	LUT2 #(
		.INIT('h8)
	) name22729 (
		_w33239_,
		_w33240_,
		_w33241_
	);
	LUT2 #(
		.INIT('h8)
	) name22730 (
		_w33237_,
		_w33238_,
		_w33242_
	);
	LUT2 #(
		.INIT('h8)
	) name22731 (
		_w33241_,
		_w33242_,
		_w33243_
	);
	LUT2 #(
		.INIT('h2)
	) name22732 (
		_w33028_,
		_w33243_,
		_w33244_
	);
	LUT2 #(
		.INIT('h1)
	) name22733 (
		_w33214_,
		_w33244_,
		_w33245_
	);
	LUT2 #(
		.INIT('h2)
	) name22734 (
		\wishbone_tx_fifo_fifo_reg[0][15]/P0001 ,
		_w33032_,
		_w33246_
	);
	LUT2 #(
		.INIT('h8)
	) name22735 (
		\wishbone_tx_fifo_fifo_reg[1][15]/P0001 ,
		_w33060_,
		_w33247_
	);
	LUT2 #(
		.INIT('h8)
	) name22736 (
		\wishbone_tx_fifo_fifo_reg[13][15]/P0001 ,
		_w33047_,
		_w33248_
	);
	LUT2 #(
		.INIT('h8)
	) name22737 (
		\wishbone_tx_fifo_fifo_reg[5][15]/P0001 ,
		_w33040_,
		_w33249_
	);
	LUT2 #(
		.INIT('h8)
	) name22738 (
		\wishbone_tx_fifo_fifo_reg[3][15]/P0001 ,
		_w33062_,
		_w33250_
	);
	LUT2 #(
		.INIT('h8)
	) name22739 (
		\wishbone_tx_fifo_fifo_reg[2][15]/P0001 ,
		_w33068_,
		_w33251_
	);
	LUT2 #(
		.INIT('h8)
	) name22740 (
		\wishbone_tx_fifo_fifo_reg[7][15]/P0001 ,
		_w33054_,
		_w33252_
	);
	LUT2 #(
		.INIT('h8)
	) name22741 (
		\wishbone_tx_fifo_fifo_reg[15][15]/P0001 ,
		_w33045_,
		_w33253_
	);
	LUT2 #(
		.INIT('h8)
	) name22742 (
		\wishbone_tx_fifo_fifo_reg[14][15]/P0001 ,
		_w33050_,
		_w33254_
	);
	LUT2 #(
		.INIT('h8)
	) name22743 (
		\wishbone_tx_fifo_fifo_reg[12][15]/P0001 ,
		_w33058_,
		_w33255_
	);
	LUT2 #(
		.INIT('h8)
	) name22744 (
		\wishbone_tx_fifo_fifo_reg[4][15]/P0001 ,
		_w33064_,
		_w33256_
	);
	LUT2 #(
		.INIT('h8)
	) name22745 (
		\wishbone_tx_fifo_fifo_reg[11][15]/P0001 ,
		_w33036_,
		_w33257_
	);
	LUT2 #(
		.INIT('h8)
	) name22746 (
		\wishbone_tx_fifo_fifo_reg[9][15]/P0001 ,
		_w33052_,
		_w33258_
	);
	LUT2 #(
		.INIT('h8)
	) name22747 (
		\wishbone_tx_fifo_fifo_reg[10][15]/P0001 ,
		_w33066_,
		_w33259_
	);
	LUT2 #(
		.INIT('h8)
	) name22748 (
		\wishbone_tx_fifo_fifo_reg[6][15]/P0001 ,
		_w33056_,
		_w33260_
	);
	LUT2 #(
		.INIT('h8)
	) name22749 (
		\wishbone_tx_fifo_fifo_reg[8][15]/P0001 ,
		_w33042_,
		_w33261_
	);
	LUT2 #(
		.INIT('h1)
	) name22750 (
		_w33247_,
		_w33248_,
		_w33262_
	);
	LUT2 #(
		.INIT('h1)
	) name22751 (
		_w33249_,
		_w33250_,
		_w33263_
	);
	LUT2 #(
		.INIT('h1)
	) name22752 (
		_w33251_,
		_w33252_,
		_w33264_
	);
	LUT2 #(
		.INIT('h1)
	) name22753 (
		_w33253_,
		_w33254_,
		_w33265_
	);
	LUT2 #(
		.INIT('h1)
	) name22754 (
		_w33255_,
		_w33256_,
		_w33266_
	);
	LUT2 #(
		.INIT('h1)
	) name22755 (
		_w33257_,
		_w33258_,
		_w33267_
	);
	LUT2 #(
		.INIT('h1)
	) name22756 (
		_w33259_,
		_w33260_,
		_w33268_
	);
	LUT2 #(
		.INIT('h4)
	) name22757 (
		_w33261_,
		_w33268_,
		_w33269_
	);
	LUT2 #(
		.INIT('h8)
	) name22758 (
		_w33266_,
		_w33267_,
		_w33270_
	);
	LUT2 #(
		.INIT('h8)
	) name22759 (
		_w33264_,
		_w33265_,
		_w33271_
	);
	LUT2 #(
		.INIT('h8)
	) name22760 (
		_w33262_,
		_w33263_,
		_w33272_
	);
	LUT2 #(
		.INIT('h8)
	) name22761 (
		_w33271_,
		_w33272_,
		_w33273_
	);
	LUT2 #(
		.INIT('h8)
	) name22762 (
		_w33269_,
		_w33270_,
		_w33274_
	);
	LUT2 #(
		.INIT('h8)
	) name22763 (
		_w33273_,
		_w33274_,
		_w33275_
	);
	LUT2 #(
		.INIT('h2)
	) name22764 (
		_w33028_,
		_w33275_,
		_w33276_
	);
	LUT2 #(
		.INIT('h1)
	) name22765 (
		_w33246_,
		_w33276_,
		_w33277_
	);
	LUT2 #(
		.INIT('h2)
	) name22766 (
		\wishbone_tx_fifo_fifo_reg[0][16]/P0001 ,
		_w33032_,
		_w33278_
	);
	LUT2 #(
		.INIT('h8)
	) name22767 (
		\wishbone_tx_fifo_fifo_reg[2][16]/P0001 ,
		_w33068_,
		_w33279_
	);
	LUT2 #(
		.INIT('h8)
	) name22768 (
		\wishbone_tx_fifo_fifo_reg[5][16]/P0001 ,
		_w33040_,
		_w33280_
	);
	LUT2 #(
		.INIT('h8)
	) name22769 (
		\wishbone_tx_fifo_fifo_reg[15][16]/P0001 ,
		_w33045_,
		_w33281_
	);
	LUT2 #(
		.INIT('h8)
	) name22770 (
		\wishbone_tx_fifo_fifo_reg[1][16]/P0001 ,
		_w33060_,
		_w33282_
	);
	LUT2 #(
		.INIT('h8)
	) name22771 (
		\wishbone_tx_fifo_fifo_reg[13][16]/P0001 ,
		_w33047_,
		_w33283_
	);
	LUT2 #(
		.INIT('h8)
	) name22772 (
		\wishbone_tx_fifo_fifo_reg[6][16]/P0001 ,
		_w33056_,
		_w33284_
	);
	LUT2 #(
		.INIT('h8)
	) name22773 (
		\wishbone_tx_fifo_fifo_reg[8][16]/P0001 ,
		_w33042_,
		_w33285_
	);
	LUT2 #(
		.INIT('h8)
	) name22774 (
		\wishbone_tx_fifo_fifo_reg[14][16]/P0001 ,
		_w33050_,
		_w33286_
	);
	LUT2 #(
		.INIT('h8)
	) name22775 (
		\wishbone_tx_fifo_fifo_reg[7][16]/P0001 ,
		_w33054_,
		_w33287_
	);
	LUT2 #(
		.INIT('h8)
	) name22776 (
		\wishbone_tx_fifo_fifo_reg[10][16]/P0001 ,
		_w33066_,
		_w33288_
	);
	LUT2 #(
		.INIT('h8)
	) name22777 (
		\wishbone_tx_fifo_fifo_reg[3][16]/P0001 ,
		_w33062_,
		_w33289_
	);
	LUT2 #(
		.INIT('h8)
	) name22778 (
		\wishbone_tx_fifo_fifo_reg[12][16]/P0001 ,
		_w33058_,
		_w33290_
	);
	LUT2 #(
		.INIT('h8)
	) name22779 (
		\wishbone_tx_fifo_fifo_reg[4][16]/P0001 ,
		_w33064_,
		_w33291_
	);
	LUT2 #(
		.INIT('h8)
	) name22780 (
		\wishbone_tx_fifo_fifo_reg[9][16]/P0001 ,
		_w33052_,
		_w33292_
	);
	LUT2 #(
		.INIT('h8)
	) name22781 (
		\wishbone_tx_fifo_fifo_reg[11][16]/P0001 ,
		_w33036_,
		_w33293_
	);
	LUT2 #(
		.INIT('h1)
	) name22782 (
		_w33279_,
		_w33280_,
		_w33294_
	);
	LUT2 #(
		.INIT('h1)
	) name22783 (
		_w33281_,
		_w33282_,
		_w33295_
	);
	LUT2 #(
		.INIT('h1)
	) name22784 (
		_w33283_,
		_w33284_,
		_w33296_
	);
	LUT2 #(
		.INIT('h1)
	) name22785 (
		_w33285_,
		_w33286_,
		_w33297_
	);
	LUT2 #(
		.INIT('h1)
	) name22786 (
		_w33287_,
		_w33288_,
		_w33298_
	);
	LUT2 #(
		.INIT('h1)
	) name22787 (
		_w33289_,
		_w33290_,
		_w33299_
	);
	LUT2 #(
		.INIT('h1)
	) name22788 (
		_w33291_,
		_w33292_,
		_w33300_
	);
	LUT2 #(
		.INIT('h4)
	) name22789 (
		_w33293_,
		_w33300_,
		_w33301_
	);
	LUT2 #(
		.INIT('h8)
	) name22790 (
		_w33298_,
		_w33299_,
		_w33302_
	);
	LUT2 #(
		.INIT('h8)
	) name22791 (
		_w33296_,
		_w33297_,
		_w33303_
	);
	LUT2 #(
		.INIT('h8)
	) name22792 (
		_w33294_,
		_w33295_,
		_w33304_
	);
	LUT2 #(
		.INIT('h8)
	) name22793 (
		_w33303_,
		_w33304_,
		_w33305_
	);
	LUT2 #(
		.INIT('h8)
	) name22794 (
		_w33301_,
		_w33302_,
		_w33306_
	);
	LUT2 #(
		.INIT('h8)
	) name22795 (
		_w33305_,
		_w33306_,
		_w33307_
	);
	LUT2 #(
		.INIT('h2)
	) name22796 (
		_w33028_,
		_w33307_,
		_w33308_
	);
	LUT2 #(
		.INIT('h1)
	) name22797 (
		_w33278_,
		_w33308_,
		_w33309_
	);
	LUT2 #(
		.INIT('h2)
	) name22798 (
		\wishbone_tx_fifo_fifo_reg[0][17]/P0001 ,
		_w33032_,
		_w33310_
	);
	LUT2 #(
		.INIT('h8)
	) name22799 (
		\wishbone_tx_fifo_fifo_reg[1][17]/P0001 ,
		_w33060_,
		_w33311_
	);
	LUT2 #(
		.INIT('h8)
	) name22800 (
		\wishbone_tx_fifo_fifo_reg[13][17]/P0001 ,
		_w33047_,
		_w33312_
	);
	LUT2 #(
		.INIT('h8)
	) name22801 (
		\wishbone_tx_fifo_fifo_reg[5][17]/P0001 ,
		_w33040_,
		_w33313_
	);
	LUT2 #(
		.INIT('h8)
	) name22802 (
		\wishbone_tx_fifo_fifo_reg[3][17]/P0001 ,
		_w33062_,
		_w33314_
	);
	LUT2 #(
		.INIT('h8)
	) name22803 (
		\wishbone_tx_fifo_fifo_reg[2][17]/P0001 ,
		_w33068_,
		_w33315_
	);
	LUT2 #(
		.INIT('h8)
	) name22804 (
		\wishbone_tx_fifo_fifo_reg[7][17]/P0001 ,
		_w33054_,
		_w33316_
	);
	LUT2 #(
		.INIT('h8)
	) name22805 (
		\wishbone_tx_fifo_fifo_reg[15][17]/P0001 ,
		_w33045_,
		_w33317_
	);
	LUT2 #(
		.INIT('h8)
	) name22806 (
		\wishbone_tx_fifo_fifo_reg[14][17]/P0001 ,
		_w33050_,
		_w33318_
	);
	LUT2 #(
		.INIT('h8)
	) name22807 (
		\wishbone_tx_fifo_fifo_reg[12][17]/P0001 ,
		_w33058_,
		_w33319_
	);
	LUT2 #(
		.INIT('h8)
	) name22808 (
		\wishbone_tx_fifo_fifo_reg[4][17]/P0001 ,
		_w33064_,
		_w33320_
	);
	LUT2 #(
		.INIT('h8)
	) name22809 (
		\wishbone_tx_fifo_fifo_reg[11][17]/P0001 ,
		_w33036_,
		_w33321_
	);
	LUT2 #(
		.INIT('h8)
	) name22810 (
		\wishbone_tx_fifo_fifo_reg[9][17]/P0001 ,
		_w33052_,
		_w33322_
	);
	LUT2 #(
		.INIT('h8)
	) name22811 (
		\wishbone_tx_fifo_fifo_reg[10][17]/P0001 ,
		_w33066_,
		_w33323_
	);
	LUT2 #(
		.INIT('h8)
	) name22812 (
		\wishbone_tx_fifo_fifo_reg[6][17]/P0001 ,
		_w33056_,
		_w33324_
	);
	LUT2 #(
		.INIT('h8)
	) name22813 (
		\wishbone_tx_fifo_fifo_reg[8][17]/P0001 ,
		_w33042_,
		_w33325_
	);
	LUT2 #(
		.INIT('h1)
	) name22814 (
		_w33311_,
		_w33312_,
		_w33326_
	);
	LUT2 #(
		.INIT('h1)
	) name22815 (
		_w33313_,
		_w33314_,
		_w33327_
	);
	LUT2 #(
		.INIT('h1)
	) name22816 (
		_w33315_,
		_w33316_,
		_w33328_
	);
	LUT2 #(
		.INIT('h1)
	) name22817 (
		_w33317_,
		_w33318_,
		_w33329_
	);
	LUT2 #(
		.INIT('h1)
	) name22818 (
		_w33319_,
		_w33320_,
		_w33330_
	);
	LUT2 #(
		.INIT('h1)
	) name22819 (
		_w33321_,
		_w33322_,
		_w33331_
	);
	LUT2 #(
		.INIT('h1)
	) name22820 (
		_w33323_,
		_w33324_,
		_w33332_
	);
	LUT2 #(
		.INIT('h4)
	) name22821 (
		_w33325_,
		_w33332_,
		_w33333_
	);
	LUT2 #(
		.INIT('h8)
	) name22822 (
		_w33330_,
		_w33331_,
		_w33334_
	);
	LUT2 #(
		.INIT('h8)
	) name22823 (
		_w33328_,
		_w33329_,
		_w33335_
	);
	LUT2 #(
		.INIT('h8)
	) name22824 (
		_w33326_,
		_w33327_,
		_w33336_
	);
	LUT2 #(
		.INIT('h8)
	) name22825 (
		_w33335_,
		_w33336_,
		_w33337_
	);
	LUT2 #(
		.INIT('h8)
	) name22826 (
		_w33333_,
		_w33334_,
		_w33338_
	);
	LUT2 #(
		.INIT('h8)
	) name22827 (
		_w33337_,
		_w33338_,
		_w33339_
	);
	LUT2 #(
		.INIT('h2)
	) name22828 (
		_w33028_,
		_w33339_,
		_w33340_
	);
	LUT2 #(
		.INIT('h1)
	) name22829 (
		_w33310_,
		_w33340_,
		_w33341_
	);
	LUT2 #(
		.INIT('h2)
	) name22830 (
		\wishbone_tx_fifo_fifo_reg[0][18]/P0001 ,
		_w33032_,
		_w33342_
	);
	LUT2 #(
		.INIT('h8)
	) name22831 (
		\wishbone_tx_fifo_fifo_reg[10][18]/P0001 ,
		_w33066_,
		_w33343_
	);
	LUT2 #(
		.INIT('h8)
	) name22832 (
		\wishbone_tx_fifo_fifo_reg[4][18]/P0001 ,
		_w33064_,
		_w33344_
	);
	LUT2 #(
		.INIT('h8)
	) name22833 (
		\wishbone_tx_fifo_fifo_reg[3][18]/P0001 ,
		_w33062_,
		_w33345_
	);
	LUT2 #(
		.INIT('h8)
	) name22834 (
		\wishbone_tx_fifo_fifo_reg[11][18]/P0001 ,
		_w33036_,
		_w33346_
	);
	LUT2 #(
		.INIT('h8)
	) name22835 (
		\wishbone_tx_fifo_fifo_reg[2][18]/P0001 ,
		_w33068_,
		_w33347_
	);
	LUT2 #(
		.INIT('h8)
	) name22836 (
		\wishbone_tx_fifo_fifo_reg[5][18]/P0001 ,
		_w33040_,
		_w33348_
	);
	LUT2 #(
		.INIT('h8)
	) name22837 (
		\wishbone_tx_fifo_fifo_reg[14][18]/P0001 ,
		_w33050_,
		_w33349_
	);
	LUT2 #(
		.INIT('h8)
	) name22838 (
		\wishbone_tx_fifo_fifo_reg[12][18]/P0001 ,
		_w33058_,
		_w33350_
	);
	LUT2 #(
		.INIT('h8)
	) name22839 (
		\wishbone_tx_fifo_fifo_reg[15][18]/P0001 ,
		_w33045_,
		_w33351_
	);
	LUT2 #(
		.INIT('h8)
	) name22840 (
		\wishbone_tx_fifo_fifo_reg[1][18]/P0001 ,
		_w33060_,
		_w33352_
	);
	LUT2 #(
		.INIT('h8)
	) name22841 (
		\wishbone_tx_fifo_fifo_reg[13][18]/P0001 ,
		_w33047_,
		_w33353_
	);
	LUT2 #(
		.INIT('h8)
	) name22842 (
		\wishbone_tx_fifo_fifo_reg[9][18]/P0001 ,
		_w33052_,
		_w33354_
	);
	LUT2 #(
		.INIT('h8)
	) name22843 (
		\wishbone_tx_fifo_fifo_reg[6][18]/P0001 ,
		_w33056_,
		_w33355_
	);
	LUT2 #(
		.INIT('h8)
	) name22844 (
		\wishbone_tx_fifo_fifo_reg[7][18]/P0001 ,
		_w33054_,
		_w33356_
	);
	LUT2 #(
		.INIT('h8)
	) name22845 (
		\wishbone_tx_fifo_fifo_reg[8][18]/P0001 ,
		_w33042_,
		_w33357_
	);
	LUT2 #(
		.INIT('h1)
	) name22846 (
		_w33343_,
		_w33344_,
		_w33358_
	);
	LUT2 #(
		.INIT('h1)
	) name22847 (
		_w33345_,
		_w33346_,
		_w33359_
	);
	LUT2 #(
		.INIT('h1)
	) name22848 (
		_w33347_,
		_w33348_,
		_w33360_
	);
	LUT2 #(
		.INIT('h1)
	) name22849 (
		_w33349_,
		_w33350_,
		_w33361_
	);
	LUT2 #(
		.INIT('h1)
	) name22850 (
		_w33351_,
		_w33352_,
		_w33362_
	);
	LUT2 #(
		.INIT('h1)
	) name22851 (
		_w33353_,
		_w33354_,
		_w33363_
	);
	LUT2 #(
		.INIT('h1)
	) name22852 (
		_w33355_,
		_w33356_,
		_w33364_
	);
	LUT2 #(
		.INIT('h4)
	) name22853 (
		_w33357_,
		_w33364_,
		_w33365_
	);
	LUT2 #(
		.INIT('h8)
	) name22854 (
		_w33362_,
		_w33363_,
		_w33366_
	);
	LUT2 #(
		.INIT('h8)
	) name22855 (
		_w33360_,
		_w33361_,
		_w33367_
	);
	LUT2 #(
		.INIT('h8)
	) name22856 (
		_w33358_,
		_w33359_,
		_w33368_
	);
	LUT2 #(
		.INIT('h8)
	) name22857 (
		_w33367_,
		_w33368_,
		_w33369_
	);
	LUT2 #(
		.INIT('h8)
	) name22858 (
		_w33365_,
		_w33366_,
		_w33370_
	);
	LUT2 #(
		.INIT('h8)
	) name22859 (
		_w33369_,
		_w33370_,
		_w33371_
	);
	LUT2 #(
		.INIT('h2)
	) name22860 (
		_w33028_,
		_w33371_,
		_w33372_
	);
	LUT2 #(
		.INIT('h1)
	) name22861 (
		_w33342_,
		_w33372_,
		_w33373_
	);
	LUT2 #(
		.INIT('h2)
	) name22862 (
		\wishbone_tx_fifo_fifo_reg[0][19]/P0001 ,
		_w33032_,
		_w33374_
	);
	LUT2 #(
		.INIT('h8)
	) name22863 (
		\wishbone_tx_fifo_fifo_reg[3][19]/P0001 ,
		_w33062_,
		_w33375_
	);
	LUT2 #(
		.INIT('h8)
	) name22864 (
		\wishbone_tx_fifo_fifo_reg[6][19]/P0001 ,
		_w33056_,
		_w33376_
	);
	LUT2 #(
		.INIT('h8)
	) name22865 (
		\wishbone_tx_fifo_fifo_reg[12][19]/P0001 ,
		_w33058_,
		_w33377_
	);
	LUT2 #(
		.INIT('h8)
	) name22866 (
		\wishbone_tx_fifo_fifo_reg[2][19]/P0001 ,
		_w33068_,
		_w33378_
	);
	LUT2 #(
		.INIT('h8)
	) name22867 (
		\wishbone_tx_fifo_fifo_reg[13][19]/P0001 ,
		_w33047_,
		_w33379_
	);
	LUT2 #(
		.INIT('h8)
	) name22868 (
		\wishbone_tx_fifo_fifo_reg[5][19]/P0001 ,
		_w33040_,
		_w33380_
	);
	LUT2 #(
		.INIT('h8)
	) name22869 (
		\wishbone_tx_fifo_fifo_reg[9][19]/P0001 ,
		_w33052_,
		_w33381_
	);
	LUT2 #(
		.INIT('h8)
	) name22870 (
		\wishbone_tx_fifo_fifo_reg[7][19]/P0001 ,
		_w33054_,
		_w33382_
	);
	LUT2 #(
		.INIT('h8)
	) name22871 (
		\wishbone_tx_fifo_fifo_reg[14][19]/P0001 ,
		_w33050_,
		_w33383_
	);
	LUT2 #(
		.INIT('h8)
	) name22872 (
		\wishbone_tx_fifo_fifo_reg[10][19]/P0001 ,
		_w33066_,
		_w33384_
	);
	LUT2 #(
		.INIT('h8)
	) name22873 (
		\wishbone_tx_fifo_fifo_reg[11][19]/P0001 ,
		_w33036_,
		_w33385_
	);
	LUT2 #(
		.INIT('h8)
	) name22874 (
		\wishbone_tx_fifo_fifo_reg[15][19]/P0001 ,
		_w33045_,
		_w33386_
	);
	LUT2 #(
		.INIT('h8)
	) name22875 (
		\wishbone_tx_fifo_fifo_reg[4][19]/P0001 ,
		_w33064_,
		_w33387_
	);
	LUT2 #(
		.INIT('h8)
	) name22876 (
		\wishbone_tx_fifo_fifo_reg[8][19]/P0001 ,
		_w33042_,
		_w33388_
	);
	LUT2 #(
		.INIT('h8)
	) name22877 (
		\wishbone_tx_fifo_fifo_reg[1][19]/P0001 ,
		_w33060_,
		_w33389_
	);
	LUT2 #(
		.INIT('h1)
	) name22878 (
		_w33375_,
		_w33376_,
		_w33390_
	);
	LUT2 #(
		.INIT('h1)
	) name22879 (
		_w33377_,
		_w33378_,
		_w33391_
	);
	LUT2 #(
		.INIT('h1)
	) name22880 (
		_w33379_,
		_w33380_,
		_w33392_
	);
	LUT2 #(
		.INIT('h1)
	) name22881 (
		_w33381_,
		_w33382_,
		_w33393_
	);
	LUT2 #(
		.INIT('h1)
	) name22882 (
		_w33383_,
		_w33384_,
		_w33394_
	);
	LUT2 #(
		.INIT('h1)
	) name22883 (
		_w33385_,
		_w33386_,
		_w33395_
	);
	LUT2 #(
		.INIT('h1)
	) name22884 (
		_w33387_,
		_w33388_,
		_w33396_
	);
	LUT2 #(
		.INIT('h4)
	) name22885 (
		_w33389_,
		_w33396_,
		_w33397_
	);
	LUT2 #(
		.INIT('h8)
	) name22886 (
		_w33394_,
		_w33395_,
		_w33398_
	);
	LUT2 #(
		.INIT('h8)
	) name22887 (
		_w33392_,
		_w33393_,
		_w33399_
	);
	LUT2 #(
		.INIT('h8)
	) name22888 (
		_w33390_,
		_w33391_,
		_w33400_
	);
	LUT2 #(
		.INIT('h8)
	) name22889 (
		_w33399_,
		_w33400_,
		_w33401_
	);
	LUT2 #(
		.INIT('h8)
	) name22890 (
		_w33397_,
		_w33398_,
		_w33402_
	);
	LUT2 #(
		.INIT('h8)
	) name22891 (
		_w33401_,
		_w33402_,
		_w33403_
	);
	LUT2 #(
		.INIT('h2)
	) name22892 (
		_w33028_,
		_w33403_,
		_w33404_
	);
	LUT2 #(
		.INIT('h1)
	) name22893 (
		_w33374_,
		_w33404_,
		_w33405_
	);
	LUT2 #(
		.INIT('h2)
	) name22894 (
		\wishbone_tx_fifo_fifo_reg[0][1]/P0001 ,
		_w33032_,
		_w33406_
	);
	LUT2 #(
		.INIT('h8)
	) name22895 (
		\wishbone_tx_fifo_fifo_reg[5][1]/P0001 ,
		_w33040_,
		_w33407_
	);
	LUT2 #(
		.INIT('h8)
	) name22896 (
		\wishbone_tx_fifo_fifo_reg[14][1]/P0001 ,
		_w33050_,
		_w33408_
	);
	LUT2 #(
		.INIT('h8)
	) name22897 (
		\wishbone_tx_fifo_fifo_reg[12][1]/P0001 ,
		_w33058_,
		_w33409_
	);
	LUT2 #(
		.INIT('h8)
	) name22898 (
		\wishbone_tx_fifo_fifo_reg[3][1]/P0001 ,
		_w33062_,
		_w33410_
	);
	LUT2 #(
		.INIT('h8)
	) name22899 (
		\wishbone_tx_fifo_fifo_reg[9][1]/P0001 ,
		_w33052_,
		_w33411_
	);
	LUT2 #(
		.INIT('h8)
	) name22900 (
		\wishbone_tx_fifo_fifo_reg[6][1]/P0001 ,
		_w33056_,
		_w33412_
	);
	LUT2 #(
		.INIT('h8)
	) name22901 (
		\wishbone_tx_fifo_fifo_reg[2][1]/P0001 ,
		_w33068_,
		_w33413_
	);
	LUT2 #(
		.INIT('h8)
	) name22902 (
		\wishbone_tx_fifo_fifo_reg[1][1]/P0001 ,
		_w33060_,
		_w33414_
	);
	LUT2 #(
		.INIT('h8)
	) name22903 (
		\wishbone_tx_fifo_fifo_reg[4][1]/P0001 ,
		_w33064_,
		_w33415_
	);
	LUT2 #(
		.INIT('h8)
	) name22904 (
		\wishbone_tx_fifo_fifo_reg[11][1]/P0001 ,
		_w33036_,
		_w33416_
	);
	LUT2 #(
		.INIT('h8)
	) name22905 (
		\wishbone_tx_fifo_fifo_reg[15][1]/P0001 ,
		_w33045_,
		_w33417_
	);
	LUT2 #(
		.INIT('h8)
	) name22906 (
		\wishbone_tx_fifo_fifo_reg[13][1]/P0001 ,
		_w33047_,
		_w33418_
	);
	LUT2 #(
		.INIT('h8)
	) name22907 (
		\wishbone_tx_fifo_fifo_reg[10][1]/P0001 ,
		_w33066_,
		_w33419_
	);
	LUT2 #(
		.INIT('h8)
	) name22908 (
		\wishbone_tx_fifo_fifo_reg[8][1]/P0001 ,
		_w33042_,
		_w33420_
	);
	LUT2 #(
		.INIT('h8)
	) name22909 (
		\wishbone_tx_fifo_fifo_reg[7][1]/P0001 ,
		_w33054_,
		_w33421_
	);
	LUT2 #(
		.INIT('h1)
	) name22910 (
		_w33407_,
		_w33408_,
		_w33422_
	);
	LUT2 #(
		.INIT('h1)
	) name22911 (
		_w33409_,
		_w33410_,
		_w33423_
	);
	LUT2 #(
		.INIT('h1)
	) name22912 (
		_w33411_,
		_w33412_,
		_w33424_
	);
	LUT2 #(
		.INIT('h1)
	) name22913 (
		_w33413_,
		_w33414_,
		_w33425_
	);
	LUT2 #(
		.INIT('h1)
	) name22914 (
		_w33415_,
		_w33416_,
		_w33426_
	);
	LUT2 #(
		.INIT('h1)
	) name22915 (
		_w33417_,
		_w33418_,
		_w33427_
	);
	LUT2 #(
		.INIT('h1)
	) name22916 (
		_w33419_,
		_w33420_,
		_w33428_
	);
	LUT2 #(
		.INIT('h4)
	) name22917 (
		_w33421_,
		_w33428_,
		_w33429_
	);
	LUT2 #(
		.INIT('h8)
	) name22918 (
		_w33426_,
		_w33427_,
		_w33430_
	);
	LUT2 #(
		.INIT('h8)
	) name22919 (
		_w33424_,
		_w33425_,
		_w33431_
	);
	LUT2 #(
		.INIT('h8)
	) name22920 (
		_w33422_,
		_w33423_,
		_w33432_
	);
	LUT2 #(
		.INIT('h8)
	) name22921 (
		_w33431_,
		_w33432_,
		_w33433_
	);
	LUT2 #(
		.INIT('h8)
	) name22922 (
		_w33429_,
		_w33430_,
		_w33434_
	);
	LUT2 #(
		.INIT('h8)
	) name22923 (
		_w33433_,
		_w33434_,
		_w33435_
	);
	LUT2 #(
		.INIT('h2)
	) name22924 (
		_w33028_,
		_w33435_,
		_w33436_
	);
	LUT2 #(
		.INIT('h1)
	) name22925 (
		_w33406_,
		_w33436_,
		_w33437_
	);
	LUT2 #(
		.INIT('h2)
	) name22926 (
		\wishbone_tx_fifo_fifo_reg[0][20]/P0001 ,
		_w33032_,
		_w33438_
	);
	LUT2 #(
		.INIT('h8)
	) name22927 (
		\wishbone_tx_fifo_fifo_reg[6][20]/P0001 ,
		_w33056_,
		_w33439_
	);
	LUT2 #(
		.INIT('h8)
	) name22928 (
		\wishbone_tx_fifo_fifo_reg[10][20]/P0001 ,
		_w33066_,
		_w33440_
	);
	LUT2 #(
		.INIT('h8)
	) name22929 (
		\wishbone_tx_fifo_fifo_reg[7][20]/P0001 ,
		_w33054_,
		_w33441_
	);
	LUT2 #(
		.INIT('h8)
	) name22930 (
		\wishbone_tx_fifo_fifo_reg[4][20]/P0001 ,
		_w33064_,
		_w33442_
	);
	LUT2 #(
		.INIT('h8)
	) name22931 (
		\wishbone_tx_fifo_fifo_reg[15][20]/P0001 ,
		_w33045_,
		_w33443_
	);
	LUT2 #(
		.INIT('h8)
	) name22932 (
		\wishbone_tx_fifo_fifo_reg[9][20]/P0001 ,
		_w33052_,
		_w33444_
	);
	LUT2 #(
		.INIT('h8)
	) name22933 (
		\wishbone_tx_fifo_fifo_reg[8][20]/P0001 ,
		_w33042_,
		_w33445_
	);
	LUT2 #(
		.INIT('h8)
	) name22934 (
		\wishbone_tx_fifo_fifo_reg[3][20]/P0001 ,
		_w33062_,
		_w33446_
	);
	LUT2 #(
		.INIT('h8)
	) name22935 (
		\wishbone_tx_fifo_fifo_reg[11][20]/P0001 ,
		_w33036_,
		_w33447_
	);
	LUT2 #(
		.INIT('h8)
	) name22936 (
		\wishbone_tx_fifo_fifo_reg[5][20]/P0001 ,
		_w33040_,
		_w33448_
	);
	LUT2 #(
		.INIT('h8)
	) name22937 (
		\wishbone_tx_fifo_fifo_reg[14][20]/P0001 ,
		_w33050_,
		_w33449_
	);
	LUT2 #(
		.INIT('h8)
	) name22938 (
		\wishbone_tx_fifo_fifo_reg[12][20]/P0001 ,
		_w33058_,
		_w33450_
	);
	LUT2 #(
		.INIT('h8)
	) name22939 (
		\wishbone_tx_fifo_fifo_reg[13][20]/P0001 ,
		_w33047_,
		_w33451_
	);
	LUT2 #(
		.INIT('h8)
	) name22940 (
		\wishbone_tx_fifo_fifo_reg[2][20]/P0001 ,
		_w33068_,
		_w33452_
	);
	LUT2 #(
		.INIT('h8)
	) name22941 (
		\wishbone_tx_fifo_fifo_reg[1][20]/P0001 ,
		_w33060_,
		_w33453_
	);
	LUT2 #(
		.INIT('h1)
	) name22942 (
		_w33439_,
		_w33440_,
		_w33454_
	);
	LUT2 #(
		.INIT('h1)
	) name22943 (
		_w33441_,
		_w33442_,
		_w33455_
	);
	LUT2 #(
		.INIT('h1)
	) name22944 (
		_w33443_,
		_w33444_,
		_w33456_
	);
	LUT2 #(
		.INIT('h1)
	) name22945 (
		_w33445_,
		_w33446_,
		_w33457_
	);
	LUT2 #(
		.INIT('h1)
	) name22946 (
		_w33447_,
		_w33448_,
		_w33458_
	);
	LUT2 #(
		.INIT('h1)
	) name22947 (
		_w33449_,
		_w33450_,
		_w33459_
	);
	LUT2 #(
		.INIT('h1)
	) name22948 (
		_w33451_,
		_w33452_,
		_w33460_
	);
	LUT2 #(
		.INIT('h4)
	) name22949 (
		_w33453_,
		_w33460_,
		_w33461_
	);
	LUT2 #(
		.INIT('h8)
	) name22950 (
		_w33458_,
		_w33459_,
		_w33462_
	);
	LUT2 #(
		.INIT('h8)
	) name22951 (
		_w33456_,
		_w33457_,
		_w33463_
	);
	LUT2 #(
		.INIT('h8)
	) name22952 (
		_w33454_,
		_w33455_,
		_w33464_
	);
	LUT2 #(
		.INIT('h8)
	) name22953 (
		_w33463_,
		_w33464_,
		_w33465_
	);
	LUT2 #(
		.INIT('h8)
	) name22954 (
		_w33461_,
		_w33462_,
		_w33466_
	);
	LUT2 #(
		.INIT('h8)
	) name22955 (
		_w33465_,
		_w33466_,
		_w33467_
	);
	LUT2 #(
		.INIT('h2)
	) name22956 (
		_w33028_,
		_w33467_,
		_w33468_
	);
	LUT2 #(
		.INIT('h1)
	) name22957 (
		_w33438_,
		_w33468_,
		_w33469_
	);
	LUT2 #(
		.INIT('h2)
	) name22958 (
		\wishbone_tx_fifo_fifo_reg[0][21]/P0001 ,
		_w33032_,
		_w33470_
	);
	LUT2 #(
		.INIT('h8)
	) name22959 (
		\wishbone_tx_fifo_fifo_reg[11][21]/P0001 ,
		_w33036_,
		_w33471_
	);
	LUT2 #(
		.INIT('h8)
	) name22960 (
		\wishbone_tx_fifo_fifo_reg[5][21]/P0001 ,
		_w33040_,
		_w33472_
	);
	LUT2 #(
		.INIT('h8)
	) name22961 (
		\wishbone_tx_fifo_fifo_reg[8][21]/P0001 ,
		_w33042_,
		_w33473_
	);
	LUT2 #(
		.INIT('h8)
	) name22962 (
		\wishbone_tx_fifo_fifo_reg[15][21]/P0001 ,
		_w33045_,
		_w33474_
	);
	LUT2 #(
		.INIT('h8)
	) name22963 (
		\wishbone_tx_fifo_fifo_reg[13][21]/P0001 ,
		_w33047_,
		_w33475_
	);
	LUT2 #(
		.INIT('h8)
	) name22964 (
		\wishbone_tx_fifo_fifo_reg[14][21]/P0001 ,
		_w33050_,
		_w33476_
	);
	LUT2 #(
		.INIT('h8)
	) name22965 (
		\wishbone_tx_fifo_fifo_reg[9][21]/P0001 ,
		_w33052_,
		_w33477_
	);
	LUT2 #(
		.INIT('h8)
	) name22966 (
		\wishbone_tx_fifo_fifo_reg[7][21]/P0001 ,
		_w33054_,
		_w33478_
	);
	LUT2 #(
		.INIT('h8)
	) name22967 (
		\wishbone_tx_fifo_fifo_reg[6][21]/P0001 ,
		_w33056_,
		_w33479_
	);
	LUT2 #(
		.INIT('h8)
	) name22968 (
		\wishbone_tx_fifo_fifo_reg[12][21]/P0001 ,
		_w33058_,
		_w33480_
	);
	LUT2 #(
		.INIT('h8)
	) name22969 (
		\wishbone_tx_fifo_fifo_reg[1][21]/P0001 ,
		_w33060_,
		_w33481_
	);
	LUT2 #(
		.INIT('h8)
	) name22970 (
		\wishbone_tx_fifo_fifo_reg[3][21]/P0001 ,
		_w33062_,
		_w33482_
	);
	LUT2 #(
		.INIT('h8)
	) name22971 (
		\wishbone_tx_fifo_fifo_reg[4][21]/P0001 ,
		_w33064_,
		_w33483_
	);
	LUT2 #(
		.INIT('h8)
	) name22972 (
		\wishbone_tx_fifo_fifo_reg[10][21]/P0001 ,
		_w33066_,
		_w33484_
	);
	LUT2 #(
		.INIT('h8)
	) name22973 (
		\wishbone_tx_fifo_fifo_reg[2][21]/P0001 ,
		_w33068_,
		_w33485_
	);
	LUT2 #(
		.INIT('h1)
	) name22974 (
		_w33471_,
		_w33472_,
		_w33486_
	);
	LUT2 #(
		.INIT('h1)
	) name22975 (
		_w33473_,
		_w33474_,
		_w33487_
	);
	LUT2 #(
		.INIT('h1)
	) name22976 (
		_w33475_,
		_w33476_,
		_w33488_
	);
	LUT2 #(
		.INIT('h1)
	) name22977 (
		_w33477_,
		_w33478_,
		_w33489_
	);
	LUT2 #(
		.INIT('h1)
	) name22978 (
		_w33479_,
		_w33480_,
		_w33490_
	);
	LUT2 #(
		.INIT('h1)
	) name22979 (
		_w33481_,
		_w33482_,
		_w33491_
	);
	LUT2 #(
		.INIT('h1)
	) name22980 (
		_w33483_,
		_w33484_,
		_w33492_
	);
	LUT2 #(
		.INIT('h4)
	) name22981 (
		_w33485_,
		_w33492_,
		_w33493_
	);
	LUT2 #(
		.INIT('h8)
	) name22982 (
		_w33490_,
		_w33491_,
		_w33494_
	);
	LUT2 #(
		.INIT('h8)
	) name22983 (
		_w33488_,
		_w33489_,
		_w33495_
	);
	LUT2 #(
		.INIT('h8)
	) name22984 (
		_w33486_,
		_w33487_,
		_w33496_
	);
	LUT2 #(
		.INIT('h8)
	) name22985 (
		_w33495_,
		_w33496_,
		_w33497_
	);
	LUT2 #(
		.INIT('h8)
	) name22986 (
		_w33493_,
		_w33494_,
		_w33498_
	);
	LUT2 #(
		.INIT('h8)
	) name22987 (
		_w33497_,
		_w33498_,
		_w33499_
	);
	LUT2 #(
		.INIT('h2)
	) name22988 (
		_w33028_,
		_w33499_,
		_w33500_
	);
	LUT2 #(
		.INIT('h1)
	) name22989 (
		_w33470_,
		_w33500_,
		_w33501_
	);
	LUT2 #(
		.INIT('h2)
	) name22990 (
		\wishbone_tx_fifo_fifo_reg[0][22]/P0001 ,
		_w33032_,
		_w33502_
	);
	LUT2 #(
		.INIT('h8)
	) name22991 (
		\wishbone_tx_fifo_fifo_reg[2][22]/P0001 ,
		_w33068_,
		_w33503_
	);
	LUT2 #(
		.INIT('h8)
	) name22992 (
		\wishbone_tx_fifo_fifo_reg[6][22]/P0001 ,
		_w33056_,
		_w33504_
	);
	LUT2 #(
		.INIT('h8)
	) name22993 (
		\wishbone_tx_fifo_fifo_reg[14][22]/P0001 ,
		_w33050_,
		_w33505_
	);
	LUT2 #(
		.INIT('h8)
	) name22994 (
		\wishbone_tx_fifo_fifo_reg[1][22]/P0001 ,
		_w33060_,
		_w33506_
	);
	LUT2 #(
		.INIT('h8)
	) name22995 (
		\wishbone_tx_fifo_fifo_reg[13][22]/P0001 ,
		_w33047_,
		_w33507_
	);
	LUT2 #(
		.INIT('h8)
	) name22996 (
		\wishbone_tx_fifo_fifo_reg[12][22]/P0001 ,
		_w33058_,
		_w33508_
	);
	LUT2 #(
		.INIT('h8)
	) name22997 (
		\wishbone_tx_fifo_fifo_reg[9][22]/P0001 ,
		_w33052_,
		_w33509_
	);
	LUT2 #(
		.INIT('h8)
	) name22998 (
		\wishbone_tx_fifo_fifo_reg[7][22]/P0001 ,
		_w33054_,
		_w33510_
	);
	LUT2 #(
		.INIT('h8)
	) name22999 (
		\wishbone_tx_fifo_fifo_reg[5][22]/P0001 ,
		_w33040_,
		_w33511_
	);
	LUT2 #(
		.INIT('h8)
	) name23000 (
		\wishbone_tx_fifo_fifo_reg[10][22]/P0001 ,
		_w33066_,
		_w33512_
	);
	LUT2 #(
		.INIT('h8)
	) name23001 (
		\wishbone_tx_fifo_fifo_reg[3][22]/P0001 ,
		_w33062_,
		_w33513_
	);
	LUT2 #(
		.INIT('h8)
	) name23002 (
		\wishbone_tx_fifo_fifo_reg[15][22]/P0001 ,
		_w33045_,
		_w33514_
	);
	LUT2 #(
		.INIT('h8)
	) name23003 (
		\wishbone_tx_fifo_fifo_reg[4][22]/P0001 ,
		_w33064_,
		_w33515_
	);
	LUT2 #(
		.INIT('h8)
	) name23004 (
		\wishbone_tx_fifo_fifo_reg[8][22]/P0001 ,
		_w33042_,
		_w33516_
	);
	LUT2 #(
		.INIT('h8)
	) name23005 (
		\wishbone_tx_fifo_fifo_reg[11][22]/P0001 ,
		_w33036_,
		_w33517_
	);
	LUT2 #(
		.INIT('h1)
	) name23006 (
		_w33503_,
		_w33504_,
		_w33518_
	);
	LUT2 #(
		.INIT('h1)
	) name23007 (
		_w33505_,
		_w33506_,
		_w33519_
	);
	LUT2 #(
		.INIT('h1)
	) name23008 (
		_w33507_,
		_w33508_,
		_w33520_
	);
	LUT2 #(
		.INIT('h1)
	) name23009 (
		_w33509_,
		_w33510_,
		_w33521_
	);
	LUT2 #(
		.INIT('h1)
	) name23010 (
		_w33511_,
		_w33512_,
		_w33522_
	);
	LUT2 #(
		.INIT('h1)
	) name23011 (
		_w33513_,
		_w33514_,
		_w33523_
	);
	LUT2 #(
		.INIT('h1)
	) name23012 (
		_w33515_,
		_w33516_,
		_w33524_
	);
	LUT2 #(
		.INIT('h4)
	) name23013 (
		_w33517_,
		_w33524_,
		_w33525_
	);
	LUT2 #(
		.INIT('h8)
	) name23014 (
		_w33522_,
		_w33523_,
		_w33526_
	);
	LUT2 #(
		.INIT('h8)
	) name23015 (
		_w33520_,
		_w33521_,
		_w33527_
	);
	LUT2 #(
		.INIT('h8)
	) name23016 (
		_w33518_,
		_w33519_,
		_w33528_
	);
	LUT2 #(
		.INIT('h8)
	) name23017 (
		_w33527_,
		_w33528_,
		_w33529_
	);
	LUT2 #(
		.INIT('h8)
	) name23018 (
		_w33525_,
		_w33526_,
		_w33530_
	);
	LUT2 #(
		.INIT('h8)
	) name23019 (
		_w33529_,
		_w33530_,
		_w33531_
	);
	LUT2 #(
		.INIT('h2)
	) name23020 (
		_w33028_,
		_w33531_,
		_w33532_
	);
	LUT2 #(
		.INIT('h1)
	) name23021 (
		_w33502_,
		_w33532_,
		_w33533_
	);
	LUT2 #(
		.INIT('h2)
	) name23022 (
		\wishbone_tx_fifo_fifo_reg[0][23]/P0001 ,
		_w33032_,
		_w33534_
	);
	LUT2 #(
		.INIT('h8)
	) name23023 (
		\wishbone_tx_fifo_fifo_reg[2][23]/P0001 ,
		_w33068_,
		_w33535_
	);
	LUT2 #(
		.INIT('h8)
	) name23024 (
		\wishbone_tx_fifo_fifo_reg[6][23]/P0001 ,
		_w33056_,
		_w33536_
	);
	LUT2 #(
		.INIT('h8)
	) name23025 (
		\wishbone_tx_fifo_fifo_reg[8][23]/P0001 ,
		_w33042_,
		_w33537_
	);
	LUT2 #(
		.INIT('h8)
	) name23026 (
		\wishbone_tx_fifo_fifo_reg[7][23]/P0001 ,
		_w33054_,
		_w33538_
	);
	LUT2 #(
		.INIT('h8)
	) name23027 (
		\wishbone_tx_fifo_fifo_reg[10][23]/P0001 ,
		_w33066_,
		_w33539_
	);
	LUT2 #(
		.INIT('h8)
	) name23028 (
		\wishbone_tx_fifo_fifo_reg[5][23]/P0001 ,
		_w33040_,
		_w33540_
	);
	LUT2 #(
		.INIT('h8)
	) name23029 (
		\wishbone_tx_fifo_fifo_reg[14][23]/P0001 ,
		_w33050_,
		_w33541_
	);
	LUT2 #(
		.INIT('h8)
	) name23030 (
		\wishbone_tx_fifo_fifo_reg[4][23]/P0001 ,
		_w33064_,
		_w33542_
	);
	LUT2 #(
		.INIT('h8)
	) name23031 (
		\wishbone_tx_fifo_fifo_reg[11][23]/P0001 ,
		_w33036_,
		_w33543_
	);
	LUT2 #(
		.INIT('h8)
	) name23032 (
		\wishbone_tx_fifo_fifo_reg[13][23]/P0001 ,
		_w33047_,
		_w33544_
	);
	LUT2 #(
		.INIT('h8)
	) name23033 (
		\wishbone_tx_fifo_fifo_reg[1][23]/P0001 ,
		_w33060_,
		_w33545_
	);
	LUT2 #(
		.INIT('h8)
	) name23034 (
		\wishbone_tx_fifo_fifo_reg[12][23]/P0001 ,
		_w33058_,
		_w33546_
	);
	LUT2 #(
		.INIT('h8)
	) name23035 (
		\wishbone_tx_fifo_fifo_reg[15][23]/P0001 ,
		_w33045_,
		_w33547_
	);
	LUT2 #(
		.INIT('h8)
	) name23036 (
		\wishbone_tx_fifo_fifo_reg[3][23]/P0001 ,
		_w33062_,
		_w33548_
	);
	LUT2 #(
		.INIT('h8)
	) name23037 (
		\wishbone_tx_fifo_fifo_reg[9][23]/P0001 ,
		_w33052_,
		_w33549_
	);
	LUT2 #(
		.INIT('h1)
	) name23038 (
		_w33535_,
		_w33536_,
		_w33550_
	);
	LUT2 #(
		.INIT('h1)
	) name23039 (
		_w33537_,
		_w33538_,
		_w33551_
	);
	LUT2 #(
		.INIT('h1)
	) name23040 (
		_w33539_,
		_w33540_,
		_w33552_
	);
	LUT2 #(
		.INIT('h1)
	) name23041 (
		_w33541_,
		_w33542_,
		_w33553_
	);
	LUT2 #(
		.INIT('h1)
	) name23042 (
		_w33543_,
		_w33544_,
		_w33554_
	);
	LUT2 #(
		.INIT('h1)
	) name23043 (
		_w33545_,
		_w33546_,
		_w33555_
	);
	LUT2 #(
		.INIT('h1)
	) name23044 (
		_w33547_,
		_w33548_,
		_w33556_
	);
	LUT2 #(
		.INIT('h4)
	) name23045 (
		_w33549_,
		_w33556_,
		_w33557_
	);
	LUT2 #(
		.INIT('h8)
	) name23046 (
		_w33554_,
		_w33555_,
		_w33558_
	);
	LUT2 #(
		.INIT('h8)
	) name23047 (
		_w33552_,
		_w33553_,
		_w33559_
	);
	LUT2 #(
		.INIT('h8)
	) name23048 (
		_w33550_,
		_w33551_,
		_w33560_
	);
	LUT2 #(
		.INIT('h8)
	) name23049 (
		_w33559_,
		_w33560_,
		_w33561_
	);
	LUT2 #(
		.INIT('h8)
	) name23050 (
		_w33557_,
		_w33558_,
		_w33562_
	);
	LUT2 #(
		.INIT('h8)
	) name23051 (
		_w33561_,
		_w33562_,
		_w33563_
	);
	LUT2 #(
		.INIT('h2)
	) name23052 (
		_w33028_,
		_w33563_,
		_w33564_
	);
	LUT2 #(
		.INIT('h1)
	) name23053 (
		_w33534_,
		_w33564_,
		_w33565_
	);
	LUT2 #(
		.INIT('h2)
	) name23054 (
		\wishbone_tx_fifo_fifo_reg[0][24]/P0001 ,
		_w33032_,
		_w33566_
	);
	LUT2 #(
		.INIT('h8)
	) name23055 (
		\wishbone_tx_fifo_fifo_reg[8][24]/P0001 ,
		_w33042_,
		_w33567_
	);
	LUT2 #(
		.INIT('h8)
	) name23056 (
		\wishbone_tx_fifo_fifo_reg[7][24]/P0001 ,
		_w33054_,
		_w33568_
	);
	LUT2 #(
		.INIT('h8)
	) name23057 (
		\wishbone_tx_fifo_fifo_reg[10][24]/P0001 ,
		_w33066_,
		_w33569_
	);
	LUT2 #(
		.INIT('h8)
	) name23058 (
		\wishbone_tx_fifo_fifo_reg[12][24]/P0001 ,
		_w33058_,
		_w33570_
	);
	LUT2 #(
		.INIT('h8)
	) name23059 (
		\wishbone_tx_fifo_fifo_reg[5][24]/P0001 ,
		_w33040_,
		_w33571_
	);
	LUT2 #(
		.INIT('h8)
	) name23060 (
		\wishbone_tx_fifo_fifo_reg[3][24]/P0001 ,
		_w33062_,
		_w33572_
	);
	LUT2 #(
		.INIT('h8)
	) name23061 (
		\wishbone_tx_fifo_fifo_reg[2][24]/P0001 ,
		_w33068_,
		_w33573_
	);
	LUT2 #(
		.INIT('h8)
	) name23062 (
		\wishbone_tx_fifo_fifo_reg[4][24]/P0001 ,
		_w33064_,
		_w33574_
	);
	LUT2 #(
		.INIT('h8)
	) name23063 (
		\wishbone_tx_fifo_fifo_reg[13][24]/P0001 ,
		_w33047_,
		_w33575_
	);
	LUT2 #(
		.INIT('h8)
	) name23064 (
		\wishbone_tx_fifo_fifo_reg[6][24]/P0001 ,
		_w33056_,
		_w33576_
	);
	LUT2 #(
		.INIT('h8)
	) name23065 (
		\wishbone_tx_fifo_fifo_reg[14][24]/P0001 ,
		_w33050_,
		_w33577_
	);
	LUT2 #(
		.INIT('h8)
	) name23066 (
		\wishbone_tx_fifo_fifo_reg[15][24]/P0001 ,
		_w33045_,
		_w33578_
	);
	LUT2 #(
		.INIT('h8)
	) name23067 (
		\wishbone_tx_fifo_fifo_reg[9][24]/P0001 ,
		_w33052_,
		_w33579_
	);
	LUT2 #(
		.INIT('h8)
	) name23068 (
		\wishbone_tx_fifo_fifo_reg[11][24]/P0001 ,
		_w33036_,
		_w33580_
	);
	LUT2 #(
		.INIT('h8)
	) name23069 (
		\wishbone_tx_fifo_fifo_reg[1][24]/P0001 ,
		_w33060_,
		_w33581_
	);
	LUT2 #(
		.INIT('h1)
	) name23070 (
		_w33567_,
		_w33568_,
		_w33582_
	);
	LUT2 #(
		.INIT('h1)
	) name23071 (
		_w33569_,
		_w33570_,
		_w33583_
	);
	LUT2 #(
		.INIT('h1)
	) name23072 (
		_w33571_,
		_w33572_,
		_w33584_
	);
	LUT2 #(
		.INIT('h1)
	) name23073 (
		_w33573_,
		_w33574_,
		_w33585_
	);
	LUT2 #(
		.INIT('h1)
	) name23074 (
		_w33575_,
		_w33576_,
		_w33586_
	);
	LUT2 #(
		.INIT('h1)
	) name23075 (
		_w33577_,
		_w33578_,
		_w33587_
	);
	LUT2 #(
		.INIT('h1)
	) name23076 (
		_w33579_,
		_w33580_,
		_w33588_
	);
	LUT2 #(
		.INIT('h4)
	) name23077 (
		_w33581_,
		_w33588_,
		_w33589_
	);
	LUT2 #(
		.INIT('h8)
	) name23078 (
		_w33586_,
		_w33587_,
		_w33590_
	);
	LUT2 #(
		.INIT('h8)
	) name23079 (
		_w33584_,
		_w33585_,
		_w33591_
	);
	LUT2 #(
		.INIT('h8)
	) name23080 (
		_w33582_,
		_w33583_,
		_w33592_
	);
	LUT2 #(
		.INIT('h8)
	) name23081 (
		_w33591_,
		_w33592_,
		_w33593_
	);
	LUT2 #(
		.INIT('h8)
	) name23082 (
		_w33589_,
		_w33590_,
		_w33594_
	);
	LUT2 #(
		.INIT('h8)
	) name23083 (
		_w33593_,
		_w33594_,
		_w33595_
	);
	LUT2 #(
		.INIT('h2)
	) name23084 (
		_w33028_,
		_w33595_,
		_w33596_
	);
	LUT2 #(
		.INIT('h1)
	) name23085 (
		_w33566_,
		_w33596_,
		_w33597_
	);
	LUT2 #(
		.INIT('h2)
	) name23086 (
		\wishbone_tx_fifo_fifo_reg[0][25]/P0001 ,
		_w33032_,
		_w33598_
	);
	LUT2 #(
		.INIT('h8)
	) name23087 (
		\wishbone_tx_fifo_fifo_reg[6][25]/P0001 ,
		_w33056_,
		_w33599_
	);
	LUT2 #(
		.INIT('h8)
	) name23088 (
		\wishbone_tx_fifo_fifo_reg[10][25]/P0001 ,
		_w33066_,
		_w33600_
	);
	LUT2 #(
		.INIT('h8)
	) name23089 (
		\wishbone_tx_fifo_fifo_reg[12][25]/P0001 ,
		_w33058_,
		_w33601_
	);
	LUT2 #(
		.INIT('h8)
	) name23090 (
		\wishbone_tx_fifo_fifo_reg[14][25]/P0001 ,
		_w33050_,
		_w33602_
	);
	LUT2 #(
		.INIT('h8)
	) name23091 (
		\wishbone_tx_fifo_fifo_reg[13][25]/P0001 ,
		_w33047_,
		_w33603_
	);
	LUT2 #(
		.INIT('h8)
	) name23092 (
		\wishbone_tx_fifo_fifo_reg[3][25]/P0001 ,
		_w33062_,
		_w33604_
	);
	LUT2 #(
		.INIT('h8)
	) name23093 (
		\wishbone_tx_fifo_fifo_reg[11][25]/P0001 ,
		_w33036_,
		_w33605_
	);
	LUT2 #(
		.INIT('h8)
	) name23094 (
		\wishbone_tx_fifo_fifo_reg[5][25]/P0001 ,
		_w33040_,
		_w33606_
	);
	LUT2 #(
		.INIT('h8)
	) name23095 (
		\wishbone_tx_fifo_fifo_reg[1][25]/P0001 ,
		_w33060_,
		_w33607_
	);
	LUT2 #(
		.INIT('h8)
	) name23096 (
		\wishbone_tx_fifo_fifo_reg[4][25]/P0001 ,
		_w33064_,
		_w33608_
	);
	LUT2 #(
		.INIT('h8)
	) name23097 (
		\wishbone_tx_fifo_fifo_reg[8][25]/P0001 ,
		_w33042_,
		_w33609_
	);
	LUT2 #(
		.INIT('h8)
	) name23098 (
		\wishbone_tx_fifo_fifo_reg[7][25]/P0001 ,
		_w33054_,
		_w33610_
	);
	LUT2 #(
		.INIT('h8)
	) name23099 (
		\wishbone_tx_fifo_fifo_reg[2][25]/P0001 ,
		_w33068_,
		_w33611_
	);
	LUT2 #(
		.INIT('h8)
	) name23100 (
		\wishbone_tx_fifo_fifo_reg[9][25]/P0001 ,
		_w33052_,
		_w33612_
	);
	LUT2 #(
		.INIT('h8)
	) name23101 (
		\wishbone_tx_fifo_fifo_reg[15][25]/P0001 ,
		_w33045_,
		_w33613_
	);
	LUT2 #(
		.INIT('h1)
	) name23102 (
		_w33599_,
		_w33600_,
		_w33614_
	);
	LUT2 #(
		.INIT('h1)
	) name23103 (
		_w33601_,
		_w33602_,
		_w33615_
	);
	LUT2 #(
		.INIT('h1)
	) name23104 (
		_w33603_,
		_w33604_,
		_w33616_
	);
	LUT2 #(
		.INIT('h1)
	) name23105 (
		_w33605_,
		_w33606_,
		_w33617_
	);
	LUT2 #(
		.INIT('h1)
	) name23106 (
		_w33607_,
		_w33608_,
		_w33618_
	);
	LUT2 #(
		.INIT('h1)
	) name23107 (
		_w33609_,
		_w33610_,
		_w33619_
	);
	LUT2 #(
		.INIT('h1)
	) name23108 (
		_w33611_,
		_w33612_,
		_w33620_
	);
	LUT2 #(
		.INIT('h4)
	) name23109 (
		_w33613_,
		_w33620_,
		_w33621_
	);
	LUT2 #(
		.INIT('h8)
	) name23110 (
		_w33618_,
		_w33619_,
		_w33622_
	);
	LUT2 #(
		.INIT('h8)
	) name23111 (
		_w33616_,
		_w33617_,
		_w33623_
	);
	LUT2 #(
		.INIT('h8)
	) name23112 (
		_w33614_,
		_w33615_,
		_w33624_
	);
	LUT2 #(
		.INIT('h8)
	) name23113 (
		_w33623_,
		_w33624_,
		_w33625_
	);
	LUT2 #(
		.INIT('h8)
	) name23114 (
		_w33621_,
		_w33622_,
		_w33626_
	);
	LUT2 #(
		.INIT('h8)
	) name23115 (
		_w33625_,
		_w33626_,
		_w33627_
	);
	LUT2 #(
		.INIT('h2)
	) name23116 (
		_w33028_,
		_w33627_,
		_w33628_
	);
	LUT2 #(
		.INIT('h1)
	) name23117 (
		_w33598_,
		_w33628_,
		_w33629_
	);
	LUT2 #(
		.INIT('h2)
	) name23118 (
		\wishbone_tx_fifo_fifo_reg[0][26]/P0001 ,
		_w33032_,
		_w33630_
	);
	LUT2 #(
		.INIT('h8)
	) name23119 (
		\wishbone_tx_fifo_fifo_reg[5][26]/P0001 ,
		_w33040_,
		_w33631_
	);
	LUT2 #(
		.INIT('h8)
	) name23120 (
		\wishbone_tx_fifo_fifo_reg[14][26]/P0001 ,
		_w33050_,
		_w33632_
	);
	LUT2 #(
		.INIT('h8)
	) name23121 (
		\wishbone_tx_fifo_fifo_reg[12][26]/P0001 ,
		_w33058_,
		_w33633_
	);
	LUT2 #(
		.INIT('h8)
	) name23122 (
		\wishbone_tx_fifo_fifo_reg[3][26]/P0001 ,
		_w33062_,
		_w33634_
	);
	LUT2 #(
		.INIT('h8)
	) name23123 (
		\wishbone_tx_fifo_fifo_reg[6][26]/P0001 ,
		_w33056_,
		_w33635_
	);
	LUT2 #(
		.INIT('h8)
	) name23124 (
		\wishbone_tx_fifo_fifo_reg[9][26]/P0001 ,
		_w33052_,
		_w33636_
	);
	LUT2 #(
		.INIT('h8)
	) name23125 (
		\wishbone_tx_fifo_fifo_reg[2][26]/P0001 ,
		_w33068_,
		_w33637_
	);
	LUT2 #(
		.INIT('h8)
	) name23126 (
		\wishbone_tx_fifo_fifo_reg[1][26]/P0001 ,
		_w33060_,
		_w33638_
	);
	LUT2 #(
		.INIT('h8)
	) name23127 (
		\wishbone_tx_fifo_fifo_reg[4][26]/P0001 ,
		_w33064_,
		_w33639_
	);
	LUT2 #(
		.INIT('h8)
	) name23128 (
		\wishbone_tx_fifo_fifo_reg[11][26]/P0001 ,
		_w33036_,
		_w33640_
	);
	LUT2 #(
		.INIT('h8)
	) name23129 (
		\wishbone_tx_fifo_fifo_reg[15][26]/P0001 ,
		_w33045_,
		_w33641_
	);
	LUT2 #(
		.INIT('h8)
	) name23130 (
		\wishbone_tx_fifo_fifo_reg[13][26]/P0001 ,
		_w33047_,
		_w33642_
	);
	LUT2 #(
		.INIT('h8)
	) name23131 (
		\wishbone_tx_fifo_fifo_reg[10][26]/P0001 ,
		_w33066_,
		_w33643_
	);
	LUT2 #(
		.INIT('h8)
	) name23132 (
		\wishbone_tx_fifo_fifo_reg[8][26]/P0001 ,
		_w33042_,
		_w33644_
	);
	LUT2 #(
		.INIT('h8)
	) name23133 (
		\wishbone_tx_fifo_fifo_reg[7][26]/P0001 ,
		_w33054_,
		_w33645_
	);
	LUT2 #(
		.INIT('h1)
	) name23134 (
		_w33631_,
		_w33632_,
		_w33646_
	);
	LUT2 #(
		.INIT('h1)
	) name23135 (
		_w33633_,
		_w33634_,
		_w33647_
	);
	LUT2 #(
		.INIT('h1)
	) name23136 (
		_w33635_,
		_w33636_,
		_w33648_
	);
	LUT2 #(
		.INIT('h1)
	) name23137 (
		_w33637_,
		_w33638_,
		_w33649_
	);
	LUT2 #(
		.INIT('h1)
	) name23138 (
		_w33639_,
		_w33640_,
		_w33650_
	);
	LUT2 #(
		.INIT('h1)
	) name23139 (
		_w33641_,
		_w33642_,
		_w33651_
	);
	LUT2 #(
		.INIT('h1)
	) name23140 (
		_w33643_,
		_w33644_,
		_w33652_
	);
	LUT2 #(
		.INIT('h4)
	) name23141 (
		_w33645_,
		_w33652_,
		_w33653_
	);
	LUT2 #(
		.INIT('h8)
	) name23142 (
		_w33650_,
		_w33651_,
		_w33654_
	);
	LUT2 #(
		.INIT('h8)
	) name23143 (
		_w33648_,
		_w33649_,
		_w33655_
	);
	LUT2 #(
		.INIT('h8)
	) name23144 (
		_w33646_,
		_w33647_,
		_w33656_
	);
	LUT2 #(
		.INIT('h8)
	) name23145 (
		_w33655_,
		_w33656_,
		_w33657_
	);
	LUT2 #(
		.INIT('h8)
	) name23146 (
		_w33653_,
		_w33654_,
		_w33658_
	);
	LUT2 #(
		.INIT('h8)
	) name23147 (
		_w33657_,
		_w33658_,
		_w33659_
	);
	LUT2 #(
		.INIT('h2)
	) name23148 (
		_w33028_,
		_w33659_,
		_w33660_
	);
	LUT2 #(
		.INIT('h1)
	) name23149 (
		_w33630_,
		_w33660_,
		_w33661_
	);
	LUT2 #(
		.INIT('h2)
	) name23150 (
		\wishbone_tx_fifo_fifo_reg[0][27]/P0001 ,
		_w33032_,
		_w33662_
	);
	LUT2 #(
		.INIT('h8)
	) name23151 (
		\wishbone_tx_fifo_fifo_reg[6][27]/P0001 ,
		_w33056_,
		_w33663_
	);
	LUT2 #(
		.INIT('h8)
	) name23152 (
		\wishbone_tx_fifo_fifo_reg[10][27]/P0001 ,
		_w33066_,
		_w33664_
	);
	LUT2 #(
		.INIT('h8)
	) name23153 (
		\wishbone_tx_fifo_fifo_reg[5][27]/P0001 ,
		_w33040_,
		_w33665_
	);
	LUT2 #(
		.INIT('h8)
	) name23154 (
		\wishbone_tx_fifo_fifo_reg[7][27]/P0001 ,
		_w33054_,
		_w33666_
	);
	LUT2 #(
		.INIT('h8)
	) name23155 (
		\wishbone_tx_fifo_fifo_reg[1][27]/P0001 ,
		_w33060_,
		_w33667_
	);
	LUT2 #(
		.INIT('h8)
	) name23156 (
		\wishbone_tx_fifo_fifo_reg[12][27]/P0001 ,
		_w33058_,
		_w33668_
	);
	LUT2 #(
		.INIT('h8)
	) name23157 (
		\wishbone_tx_fifo_fifo_reg[9][27]/P0001 ,
		_w33052_,
		_w33669_
	);
	LUT2 #(
		.INIT('h8)
	) name23158 (
		\wishbone_tx_fifo_fifo_reg[11][27]/P0001 ,
		_w33036_,
		_w33670_
	);
	LUT2 #(
		.INIT('h8)
	) name23159 (
		\wishbone_tx_fifo_fifo_reg[4][27]/P0001 ,
		_w33064_,
		_w33671_
	);
	LUT2 #(
		.INIT('h8)
	) name23160 (
		\wishbone_tx_fifo_fifo_reg[3][27]/P0001 ,
		_w33062_,
		_w33672_
	);
	LUT2 #(
		.INIT('h8)
	) name23161 (
		\wishbone_tx_fifo_fifo_reg[13][27]/P0001 ,
		_w33047_,
		_w33673_
	);
	LUT2 #(
		.INIT('h8)
	) name23162 (
		\wishbone_tx_fifo_fifo_reg[14][27]/P0001 ,
		_w33050_,
		_w33674_
	);
	LUT2 #(
		.INIT('h8)
	) name23163 (
		\wishbone_tx_fifo_fifo_reg[15][27]/P0001 ,
		_w33045_,
		_w33675_
	);
	LUT2 #(
		.INIT('h8)
	) name23164 (
		\wishbone_tx_fifo_fifo_reg[2][27]/P0001 ,
		_w33068_,
		_w33676_
	);
	LUT2 #(
		.INIT('h8)
	) name23165 (
		\wishbone_tx_fifo_fifo_reg[8][27]/P0001 ,
		_w33042_,
		_w33677_
	);
	LUT2 #(
		.INIT('h1)
	) name23166 (
		_w33663_,
		_w33664_,
		_w33678_
	);
	LUT2 #(
		.INIT('h1)
	) name23167 (
		_w33665_,
		_w33666_,
		_w33679_
	);
	LUT2 #(
		.INIT('h1)
	) name23168 (
		_w33667_,
		_w33668_,
		_w33680_
	);
	LUT2 #(
		.INIT('h1)
	) name23169 (
		_w33669_,
		_w33670_,
		_w33681_
	);
	LUT2 #(
		.INIT('h1)
	) name23170 (
		_w33671_,
		_w33672_,
		_w33682_
	);
	LUT2 #(
		.INIT('h1)
	) name23171 (
		_w33673_,
		_w33674_,
		_w33683_
	);
	LUT2 #(
		.INIT('h1)
	) name23172 (
		_w33675_,
		_w33676_,
		_w33684_
	);
	LUT2 #(
		.INIT('h4)
	) name23173 (
		_w33677_,
		_w33684_,
		_w33685_
	);
	LUT2 #(
		.INIT('h8)
	) name23174 (
		_w33682_,
		_w33683_,
		_w33686_
	);
	LUT2 #(
		.INIT('h8)
	) name23175 (
		_w33680_,
		_w33681_,
		_w33687_
	);
	LUT2 #(
		.INIT('h8)
	) name23176 (
		_w33678_,
		_w33679_,
		_w33688_
	);
	LUT2 #(
		.INIT('h8)
	) name23177 (
		_w33687_,
		_w33688_,
		_w33689_
	);
	LUT2 #(
		.INIT('h8)
	) name23178 (
		_w33685_,
		_w33686_,
		_w33690_
	);
	LUT2 #(
		.INIT('h8)
	) name23179 (
		_w33689_,
		_w33690_,
		_w33691_
	);
	LUT2 #(
		.INIT('h2)
	) name23180 (
		_w33028_,
		_w33691_,
		_w33692_
	);
	LUT2 #(
		.INIT('h1)
	) name23181 (
		_w33662_,
		_w33692_,
		_w33693_
	);
	LUT2 #(
		.INIT('h2)
	) name23182 (
		\wishbone_tx_fifo_fifo_reg[0][28]/P0001 ,
		_w33032_,
		_w33694_
	);
	LUT2 #(
		.INIT('h8)
	) name23183 (
		\wishbone_tx_fifo_fifo_reg[12][28]/P0001 ,
		_w33058_,
		_w33695_
	);
	LUT2 #(
		.INIT('h8)
	) name23184 (
		\wishbone_tx_fifo_fifo_reg[5][28]/P0001 ,
		_w33040_,
		_w33696_
	);
	LUT2 #(
		.INIT('h8)
	) name23185 (
		\wishbone_tx_fifo_fifo_reg[4][28]/P0001 ,
		_w33064_,
		_w33697_
	);
	LUT2 #(
		.INIT('h8)
	) name23186 (
		\wishbone_tx_fifo_fifo_reg[8][28]/P0001 ,
		_w33042_,
		_w33698_
	);
	LUT2 #(
		.INIT('h8)
	) name23187 (
		\wishbone_tx_fifo_fifo_reg[14][28]/P0001 ,
		_w33050_,
		_w33699_
	);
	LUT2 #(
		.INIT('h8)
	) name23188 (
		\wishbone_tx_fifo_fifo_reg[6][28]/P0001 ,
		_w33056_,
		_w33700_
	);
	LUT2 #(
		.INIT('h8)
	) name23189 (
		\wishbone_tx_fifo_fifo_reg[1][28]/P0001 ,
		_w33060_,
		_w33701_
	);
	LUT2 #(
		.INIT('h8)
	) name23190 (
		\wishbone_tx_fifo_fifo_reg[10][28]/P0001 ,
		_w33066_,
		_w33702_
	);
	LUT2 #(
		.INIT('h8)
	) name23191 (
		\wishbone_tx_fifo_fifo_reg[7][28]/P0001 ,
		_w33054_,
		_w33703_
	);
	LUT2 #(
		.INIT('h8)
	) name23192 (
		\wishbone_tx_fifo_fifo_reg[2][28]/P0001 ,
		_w33068_,
		_w33704_
	);
	LUT2 #(
		.INIT('h8)
	) name23193 (
		\wishbone_tx_fifo_fifo_reg[13][28]/P0001 ,
		_w33047_,
		_w33705_
	);
	LUT2 #(
		.INIT('h8)
	) name23194 (
		\wishbone_tx_fifo_fifo_reg[9][28]/P0001 ,
		_w33052_,
		_w33706_
	);
	LUT2 #(
		.INIT('h8)
	) name23195 (
		\wishbone_tx_fifo_fifo_reg[15][28]/P0001 ,
		_w33045_,
		_w33707_
	);
	LUT2 #(
		.INIT('h8)
	) name23196 (
		\wishbone_tx_fifo_fifo_reg[3][28]/P0001 ,
		_w33062_,
		_w33708_
	);
	LUT2 #(
		.INIT('h8)
	) name23197 (
		\wishbone_tx_fifo_fifo_reg[11][28]/P0001 ,
		_w33036_,
		_w33709_
	);
	LUT2 #(
		.INIT('h1)
	) name23198 (
		_w33695_,
		_w33696_,
		_w33710_
	);
	LUT2 #(
		.INIT('h1)
	) name23199 (
		_w33697_,
		_w33698_,
		_w33711_
	);
	LUT2 #(
		.INIT('h1)
	) name23200 (
		_w33699_,
		_w33700_,
		_w33712_
	);
	LUT2 #(
		.INIT('h1)
	) name23201 (
		_w33701_,
		_w33702_,
		_w33713_
	);
	LUT2 #(
		.INIT('h1)
	) name23202 (
		_w33703_,
		_w33704_,
		_w33714_
	);
	LUT2 #(
		.INIT('h1)
	) name23203 (
		_w33705_,
		_w33706_,
		_w33715_
	);
	LUT2 #(
		.INIT('h1)
	) name23204 (
		_w33707_,
		_w33708_,
		_w33716_
	);
	LUT2 #(
		.INIT('h4)
	) name23205 (
		_w33709_,
		_w33716_,
		_w33717_
	);
	LUT2 #(
		.INIT('h8)
	) name23206 (
		_w33714_,
		_w33715_,
		_w33718_
	);
	LUT2 #(
		.INIT('h8)
	) name23207 (
		_w33712_,
		_w33713_,
		_w33719_
	);
	LUT2 #(
		.INIT('h8)
	) name23208 (
		_w33710_,
		_w33711_,
		_w33720_
	);
	LUT2 #(
		.INIT('h8)
	) name23209 (
		_w33719_,
		_w33720_,
		_w33721_
	);
	LUT2 #(
		.INIT('h8)
	) name23210 (
		_w33717_,
		_w33718_,
		_w33722_
	);
	LUT2 #(
		.INIT('h8)
	) name23211 (
		_w33721_,
		_w33722_,
		_w33723_
	);
	LUT2 #(
		.INIT('h2)
	) name23212 (
		_w33028_,
		_w33723_,
		_w33724_
	);
	LUT2 #(
		.INIT('h1)
	) name23213 (
		_w33694_,
		_w33724_,
		_w33725_
	);
	LUT2 #(
		.INIT('h2)
	) name23214 (
		\wishbone_tx_fifo_fifo_reg[0][29]/P0001 ,
		_w33032_,
		_w33726_
	);
	LUT2 #(
		.INIT('h8)
	) name23215 (
		\wishbone_tx_fifo_fifo_reg[3][29]/P0001 ,
		_w33062_,
		_w33727_
	);
	LUT2 #(
		.INIT('h8)
	) name23216 (
		\wishbone_tx_fifo_fifo_reg[13][29]/P0001 ,
		_w33047_,
		_w33728_
	);
	LUT2 #(
		.INIT('h8)
	) name23217 (
		\wishbone_tx_fifo_fifo_reg[1][29]/P0001 ,
		_w33060_,
		_w33729_
	);
	LUT2 #(
		.INIT('h8)
	) name23218 (
		\wishbone_tx_fifo_fifo_reg[12][29]/P0001 ,
		_w33058_,
		_w33730_
	);
	LUT2 #(
		.INIT('h8)
	) name23219 (
		\wishbone_tx_fifo_fifo_reg[11][29]/P0001 ,
		_w33036_,
		_w33731_
	);
	LUT2 #(
		.INIT('h8)
	) name23220 (
		\wishbone_tx_fifo_fifo_reg[10][29]/P0001 ,
		_w33066_,
		_w33732_
	);
	LUT2 #(
		.INIT('h8)
	) name23221 (
		\wishbone_tx_fifo_fifo_reg[8][29]/P0001 ,
		_w33042_,
		_w33733_
	);
	LUT2 #(
		.INIT('h8)
	) name23222 (
		\wishbone_tx_fifo_fifo_reg[4][29]/P0001 ,
		_w33064_,
		_w33734_
	);
	LUT2 #(
		.INIT('h8)
	) name23223 (
		\wishbone_tx_fifo_fifo_reg[6][29]/P0001 ,
		_w33056_,
		_w33735_
	);
	LUT2 #(
		.INIT('h8)
	) name23224 (
		\wishbone_tx_fifo_fifo_reg[7][29]/P0001 ,
		_w33054_,
		_w33736_
	);
	LUT2 #(
		.INIT('h8)
	) name23225 (
		\wishbone_tx_fifo_fifo_reg[5][29]/P0001 ,
		_w33040_,
		_w33737_
	);
	LUT2 #(
		.INIT('h8)
	) name23226 (
		\wishbone_tx_fifo_fifo_reg[2][29]/P0001 ,
		_w33068_,
		_w33738_
	);
	LUT2 #(
		.INIT('h8)
	) name23227 (
		\wishbone_tx_fifo_fifo_reg[9][29]/P0001 ,
		_w33052_,
		_w33739_
	);
	LUT2 #(
		.INIT('h8)
	) name23228 (
		\wishbone_tx_fifo_fifo_reg[14][29]/P0001 ,
		_w33050_,
		_w33740_
	);
	LUT2 #(
		.INIT('h8)
	) name23229 (
		\wishbone_tx_fifo_fifo_reg[15][29]/P0001 ,
		_w33045_,
		_w33741_
	);
	LUT2 #(
		.INIT('h1)
	) name23230 (
		_w33727_,
		_w33728_,
		_w33742_
	);
	LUT2 #(
		.INIT('h1)
	) name23231 (
		_w33729_,
		_w33730_,
		_w33743_
	);
	LUT2 #(
		.INIT('h1)
	) name23232 (
		_w33731_,
		_w33732_,
		_w33744_
	);
	LUT2 #(
		.INIT('h1)
	) name23233 (
		_w33733_,
		_w33734_,
		_w33745_
	);
	LUT2 #(
		.INIT('h1)
	) name23234 (
		_w33735_,
		_w33736_,
		_w33746_
	);
	LUT2 #(
		.INIT('h1)
	) name23235 (
		_w33737_,
		_w33738_,
		_w33747_
	);
	LUT2 #(
		.INIT('h1)
	) name23236 (
		_w33739_,
		_w33740_,
		_w33748_
	);
	LUT2 #(
		.INIT('h4)
	) name23237 (
		_w33741_,
		_w33748_,
		_w33749_
	);
	LUT2 #(
		.INIT('h8)
	) name23238 (
		_w33746_,
		_w33747_,
		_w33750_
	);
	LUT2 #(
		.INIT('h8)
	) name23239 (
		_w33744_,
		_w33745_,
		_w33751_
	);
	LUT2 #(
		.INIT('h8)
	) name23240 (
		_w33742_,
		_w33743_,
		_w33752_
	);
	LUT2 #(
		.INIT('h8)
	) name23241 (
		_w33751_,
		_w33752_,
		_w33753_
	);
	LUT2 #(
		.INIT('h8)
	) name23242 (
		_w33749_,
		_w33750_,
		_w33754_
	);
	LUT2 #(
		.INIT('h8)
	) name23243 (
		_w33753_,
		_w33754_,
		_w33755_
	);
	LUT2 #(
		.INIT('h2)
	) name23244 (
		_w33028_,
		_w33755_,
		_w33756_
	);
	LUT2 #(
		.INIT('h1)
	) name23245 (
		_w33726_,
		_w33756_,
		_w33757_
	);
	LUT2 #(
		.INIT('h2)
	) name23246 (
		\wishbone_tx_fifo_fifo_reg[0][2]/P0001 ,
		_w33032_,
		_w33758_
	);
	LUT2 #(
		.INIT('h8)
	) name23247 (
		\wishbone_tx_fifo_fifo_reg[1][2]/P0001 ,
		_w33060_,
		_w33759_
	);
	LUT2 #(
		.INIT('h8)
	) name23248 (
		\wishbone_tx_fifo_fifo_reg[13][2]/P0001 ,
		_w33047_,
		_w33760_
	);
	LUT2 #(
		.INIT('h8)
	) name23249 (
		\wishbone_tx_fifo_fifo_reg[5][2]/P0001 ,
		_w33040_,
		_w33761_
	);
	LUT2 #(
		.INIT('h8)
	) name23250 (
		\wishbone_tx_fifo_fifo_reg[3][2]/P0001 ,
		_w33062_,
		_w33762_
	);
	LUT2 #(
		.INIT('h8)
	) name23251 (
		\wishbone_tx_fifo_fifo_reg[2][2]/P0001 ,
		_w33068_,
		_w33763_
	);
	LUT2 #(
		.INIT('h8)
	) name23252 (
		\wishbone_tx_fifo_fifo_reg[7][2]/P0001 ,
		_w33054_,
		_w33764_
	);
	LUT2 #(
		.INIT('h8)
	) name23253 (
		\wishbone_tx_fifo_fifo_reg[15][2]/P0001 ,
		_w33045_,
		_w33765_
	);
	LUT2 #(
		.INIT('h8)
	) name23254 (
		\wishbone_tx_fifo_fifo_reg[14][2]/P0001 ,
		_w33050_,
		_w33766_
	);
	LUT2 #(
		.INIT('h8)
	) name23255 (
		\wishbone_tx_fifo_fifo_reg[12][2]/P0001 ,
		_w33058_,
		_w33767_
	);
	LUT2 #(
		.INIT('h8)
	) name23256 (
		\wishbone_tx_fifo_fifo_reg[4][2]/P0001 ,
		_w33064_,
		_w33768_
	);
	LUT2 #(
		.INIT('h8)
	) name23257 (
		\wishbone_tx_fifo_fifo_reg[11][2]/P0001 ,
		_w33036_,
		_w33769_
	);
	LUT2 #(
		.INIT('h8)
	) name23258 (
		\wishbone_tx_fifo_fifo_reg[9][2]/P0001 ,
		_w33052_,
		_w33770_
	);
	LUT2 #(
		.INIT('h8)
	) name23259 (
		\wishbone_tx_fifo_fifo_reg[10][2]/P0001 ,
		_w33066_,
		_w33771_
	);
	LUT2 #(
		.INIT('h8)
	) name23260 (
		\wishbone_tx_fifo_fifo_reg[6][2]/P0001 ,
		_w33056_,
		_w33772_
	);
	LUT2 #(
		.INIT('h8)
	) name23261 (
		\wishbone_tx_fifo_fifo_reg[8][2]/P0001 ,
		_w33042_,
		_w33773_
	);
	LUT2 #(
		.INIT('h1)
	) name23262 (
		_w33759_,
		_w33760_,
		_w33774_
	);
	LUT2 #(
		.INIT('h1)
	) name23263 (
		_w33761_,
		_w33762_,
		_w33775_
	);
	LUT2 #(
		.INIT('h1)
	) name23264 (
		_w33763_,
		_w33764_,
		_w33776_
	);
	LUT2 #(
		.INIT('h1)
	) name23265 (
		_w33765_,
		_w33766_,
		_w33777_
	);
	LUT2 #(
		.INIT('h1)
	) name23266 (
		_w33767_,
		_w33768_,
		_w33778_
	);
	LUT2 #(
		.INIT('h1)
	) name23267 (
		_w33769_,
		_w33770_,
		_w33779_
	);
	LUT2 #(
		.INIT('h1)
	) name23268 (
		_w33771_,
		_w33772_,
		_w33780_
	);
	LUT2 #(
		.INIT('h4)
	) name23269 (
		_w33773_,
		_w33780_,
		_w33781_
	);
	LUT2 #(
		.INIT('h8)
	) name23270 (
		_w33778_,
		_w33779_,
		_w33782_
	);
	LUT2 #(
		.INIT('h8)
	) name23271 (
		_w33776_,
		_w33777_,
		_w33783_
	);
	LUT2 #(
		.INIT('h8)
	) name23272 (
		_w33774_,
		_w33775_,
		_w33784_
	);
	LUT2 #(
		.INIT('h8)
	) name23273 (
		_w33783_,
		_w33784_,
		_w33785_
	);
	LUT2 #(
		.INIT('h8)
	) name23274 (
		_w33781_,
		_w33782_,
		_w33786_
	);
	LUT2 #(
		.INIT('h8)
	) name23275 (
		_w33785_,
		_w33786_,
		_w33787_
	);
	LUT2 #(
		.INIT('h2)
	) name23276 (
		_w33028_,
		_w33787_,
		_w33788_
	);
	LUT2 #(
		.INIT('h1)
	) name23277 (
		_w33758_,
		_w33788_,
		_w33789_
	);
	LUT2 #(
		.INIT('h2)
	) name23278 (
		\wishbone_tx_fifo_fifo_reg[0][30]/P0001 ,
		_w33032_,
		_w33790_
	);
	LUT2 #(
		.INIT('h8)
	) name23279 (
		\wishbone_tx_fifo_fifo_reg[6][30]/P0001 ,
		_w33056_,
		_w33791_
	);
	LUT2 #(
		.INIT('h8)
	) name23280 (
		\wishbone_tx_fifo_fifo_reg[12][30]/P0001 ,
		_w33058_,
		_w33792_
	);
	LUT2 #(
		.INIT('h8)
	) name23281 (
		\wishbone_tx_fifo_fifo_reg[8][30]/P0001 ,
		_w33042_,
		_w33793_
	);
	LUT2 #(
		.INIT('h8)
	) name23282 (
		\wishbone_tx_fifo_fifo_reg[11][30]/P0001 ,
		_w33036_,
		_w33794_
	);
	LUT2 #(
		.INIT('h8)
	) name23283 (
		\wishbone_tx_fifo_fifo_reg[5][30]/P0001 ,
		_w33040_,
		_w33795_
	);
	LUT2 #(
		.INIT('h8)
	) name23284 (
		\wishbone_tx_fifo_fifo_reg[9][30]/P0001 ,
		_w33052_,
		_w33796_
	);
	LUT2 #(
		.INIT('h8)
	) name23285 (
		\wishbone_tx_fifo_fifo_reg[10][30]/P0001 ,
		_w33066_,
		_w33797_
	);
	LUT2 #(
		.INIT('h8)
	) name23286 (
		\wishbone_tx_fifo_fifo_reg[13][30]/P0001 ,
		_w33047_,
		_w33798_
	);
	LUT2 #(
		.INIT('h8)
	) name23287 (
		\wishbone_tx_fifo_fifo_reg[1][30]/P0001 ,
		_w33060_,
		_w33799_
	);
	LUT2 #(
		.INIT('h8)
	) name23288 (
		\wishbone_tx_fifo_fifo_reg[15][30]/P0001 ,
		_w33045_,
		_w33800_
	);
	LUT2 #(
		.INIT('h8)
	) name23289 (
		\wishbone_tx_fifo_fifo_reg[4][30]/P0001 ,
		_w33064_,
		_w33801_
	);
	LUT2 #(
		.INIT('h8)
	) name23290 (
		\wishbone_tx_fifo_fifo_reg[3][30]/P0001 ,
		_w33062_,
		_w33802_
	);
	LUT2 #(
		.INIT('h8)
	) name23291 (
		\wishbone_tx_fifo_fifo_reg[7][30]/P0001 ,
		_w33054_,
		_w33803_
	);
	LUT2 #(
		.INIT('h8)
	) name23292 (
		\wishbone_tx_fifo_fifo_reg[14][30]/P0001 ,
		_w33050_,
		_w33804_
	);
	LUT2 #(
		.INIT('h8)
	) name23293 (
		\wishbone_tx_fifo_fifo_reg[2][30]/P0001 ,
		_w33068_,
		_w33805_
	);
	LUT2 #(
		.INIT('h1)
	) name23294 (
		_w33791_,
		_w33792_,
		_w33806_
	);
	LUT2 #(
		.INIT('h1)
	) name23295 (
		_w33793_,
		_w33794_,
		_w33807_
	);
	LUT2 #(
		.INIT('h1)
	) name23296 (
		_w33795_,
		_w33796_,
		_w33808_
	);
	LUT2 #(
		.INIT('h1)
	) name23297 (
		_w33797_,
		_w33798_,
		_w33809_
	);
	LUT2 #(
		.INIT('h1)
	) name23298 (
		_w33799_,
		_w33800_,
		_w33810_
	);
	LUT2 #(
		.INIT('h1)
	) name23299 (
		_w33801_,
		_w33802_,
		_w33811_
	);
	LUT2 #(
		.INIT('h1)
	) name23300 (
		_w33803_,
		_w33804_,
		_w33812_
	);
	LUT2 #(
		.INIT('h4)
	) name23301 (
		_w33805_,
		_w33812_,
		_w33813_
	);
	LUT2 #(
		.INIT('h8)
	) name23302 (
		_w33810_,
		_w33811_,
		_w33814_
	);
	LUT2 #(
		.INIT('h8)
	) name23303 (
		_w33808_,
		_w33809_,
		_w33815_
	);
	LUT2 #(
		.INIT('h8)
	) name23304 (
		_w33806_,
		_w33807_,
		_w33816_
	);
	LUT2 #(
		.INIT('h8)
	) name23305 (
		_w33815_,
		_w33816_,
		_w33817_
	);
	LUT2 #(
		.INIT('h8)
	) name23306 (
		_w33813_,
		_w33814_,
		_w33818_
	);
	LUT2 #(
		.INIT('h8)
	) name23307 (
		_w33817_,
		_w33818_,
		_w33819_
	);
	LUT2 #(
		.INIT('h2)
	) name23308 (
		_w33028_,
		_w33819_,
		_w33820_
	);
	LUT2 #(
		.INIT('h1)
	) name23309 (
		_w33790_,
		_w33820_,
		_w33821_
	);
	LUT2 #(
		.INIT('h2)
	) name23310 (
		\wishbone_tx_fifo_fifo_reg[0][31]/P0001 ,
		_w33032_,
		_w33822_
	);
	LUT2 #(
		.INIT('h8)
	) name23311 (
		\wishbone_tx_fifo_fifo_reg[2][31]/P0001 ,
		_w33068_,
		_w33823_
	);
	LUT2 #(
		.INIT('h8)
	) name23312 (
		\wishbone_tx_fifo_fifo_reg[13][31]/P0001 ,
		_w33047_,
		_w33824_
	);
	LUT2 #(
		.INIT('h8)
	) name23313 (
		\wishbone_tx_fifo_fifo_reg[5][31]/P0001 ,
		_w33040_,
		_w33825_
	);
	LUT2 #(
		.INIT('h8)
	) name23314 (
		\wishbone_tx_fifo_fifo_reg[11][31]/P0001 ,
		_w33036_,
		_w33826_
	);
	LUT2 #(
		.INIT('h8)
	) name23315 (
		\wishbone_tx_fifo_fifo_reg[3][31]/P0001 ,
		_w33062_,
		_w33827_
	);
	LUT2 #(
		.INIT('h8)
	) name23316 (
		\wishbone_tx_fifo_fifo_reg[7][31]/P0001 ,
		_w33054_,
		_w33828_
	);
	LUT2 #(
		.INIT('h8)
	) name23317 (
		\wishbone_tx_fifo_fifo_reg[15][31]/P0001 ,
		_w33045_,
		_w33829_
	);
	LUT2 #(
		.INIT('h8)
	) name23318 (
		\wishbone_tx_fifo_fifo_reg[14][31]/P0001 ,
		_w33050_,
		_w33830_
	);
	LUT2 #(
		.INIT('h8)
	) name23319 (
		\wishbone_tx_fifo_fifo_reg[12][31]/P0001 ,
		_w33058_,
		_w33831_
	);
	LUT2 #(
		.INIT('h8)
	) name23320 (
		\wishbone_tx_fifo_fifo_reg[4][31]/P0001 ,
		_w33064_,
		_w33832_
	);
	LUT2 #(
		.INIT('h8)
	) name23321 (
		\wishbone_tx_fifo_fifo_reg[1][31]/P0001 ,
		_w33060_,
		_w33833_
	);
	LUT2 #(
		.INIT('h8)
	) name23322 (
		\wishbone_tx_fifo_fifo_reg[9][31]/P0001 ,
		_w33052_,
		_w33834_
	);
	LUT2 #(
		.INIT('h8)
	) name23323 (
		\wishbone_tx_fifo_fifo_reg[10][31]/P0001 ,
		_w33066_,
		_w33835_
	);
	LUT2 #(
		.INIT('h8)
	) name23324 (
		\wishbone_tx_fifo_fifo_reg[6][31]/P0001 ,
		_w33056_,
		_w33836_
	);
	LUT2 #(
		.INIT('h8)
	) name23325 (
		\wishbone_tx_fifo_fifo_reg[8][31]/P0001 ,
		_w33042_,
		_w33837_
	);
	LUT2 #(
		.INIT('h1)
	) name23326 (
		_w33823_,
		_w33824_,
		_w33838_
	);
	LUT2 #(
		.INIT('h1)
	) name23327 (
		_w33825_,
		_w33826_,
		_w33839_
	);
	LUT2 #(
		.INIT('h1)
	) name23328 (
		_w33827_,
		_w33828_,
		_w33840_
	);
	LUT2 #(
		.INIT('h1)
	) name23329 (
		_w33829_,
		_w33830_,
		_w33841_
	);
	LUT2 #(
		.INIT('h1)
	) name23330 (
		_w33831_,
		_w33832_,
		_w33842_
	);
	LUT2 #(
		.INIT('h1)
	) name23331 (
		_w33833_,
		_w33834_,
		_w33843_
	);
	LUT2 #(
		.INIT('h1)
	) name23332 (
		_w33835_,
		_w33836_,
		_w33844_
	);
	LUT2 #(
		.INIT('h4)
	) name23333 (
		_w33837_,
		_w33844_,
		_w33845_
	);
	LUT2 #(
		.INIT('h8)
	) name23334 (
		_w33842_,
		_w33843_,
		_w33846_
	);
	LUT2 #(
		.INIT('h8)
	) name23335 (
		_w33840_,
		_w33841_,
		_w33847_
	);
	LUT2 #(
		.INIT('h8)
	) name23336 (
		_w33838_,
		_w33839_,
		_w33848_
	);
	LUT2 #(
		.INIT('h8)
	) name23337 (
		_w33847_,
		_w33848_,
		_w33849_
	);
	LUT2 #(
		.INIT('h8)
	) name23338 (
		_w33845_,
		_w33846_,
		_w33850_
	);
	LUT2 #(
		.INIT('h8)
	) name23339 (
		_w33849_,
		_w33850_,
		_w33851_
	);
	LUT2 #(
		.INIT('h2)
	) name23340 (
		_w33028_,
		_w33851_,
		_w33852_
	);
	LUT2 #(
		.INIT('h1)
	) name23341 (
		_w33822_,
		_w33852_,
		_w33853_
	);
	LUT2 #(
		.INIT('h2)
	) name23342 (
		\wishbone_tx_fifo_fifo_reg[0][3]/P0001 ,
		_w33032_,
		_w33854_
	);
	LUT2 #(
		.INIT('h8)
	) name23343 (
		\wishbone_tx_fifo_fifo_reg[12][3]/P0001 ,
		_w33058_,
		_w33855_
	);
	LUT2 #(
		.INIT('h8)
	) name23344 (
		\wishbone_tx_fifo_fifo_reg[10][3]/P0001 ,
		_w33066_,
		_w33856_
	);
	LUT2 #(
		.INIT('h8)
	) name23345 (
		\wishbone_tx_fifo_fifo_reg[5][3]/P0001 ,
		_w33040_,
		_w33857_
	);
	LUT2 #(
		.INIT('h8)
	) name23346 (
		\wishbone_tx_fifo_fifo_reg[8][3]/P0001 ,
		_w33042_,
		_w33858_
	);
	LUT2 #(
		.INIT('h8)
	) name23347 (
		\wishbone_tx_fifo_fifo_reg[15][3]/P0001 ,
		_w33045_,
		_w33859_
	);
	LUT2 #(
		.INIT('h8)
	) name23348 (
		\wishbone_tx_fifo_fifo_reg[6][3]/P0001 ,
		_w33056_,
		_w33860_
	);
	LUT2 #(
		.INIT('h8)
	) name23349 (
		\wishbone_tx_fifo_fifo_reg[3][3]/P0001 ,
		_w33062_,
		_w33861_
	);
	LUT2 #(
		.INIT('h8)
	) name23350 (
		\wishbone_tx_fifo_fifo_reg[11][3]/P0001 ,
		_w33036_,
		_w33862_
	);
	LUT2 #(
		.INIT('h8)
	) name23351 (
		\wishbone_tx_fifo_fifo_reg[13][3]/P0001 ,
		_w33047_,
		_w33863_
	);
	LUT2 #(
		.INIT('h8)
	) name23352 (
		\wishbone_tx_fifo_fifo_reg[9][3]/P0001 ,
		_w33052_,
		_w33864_
	);
	LUT2 #(
		.INIT('h8)
	) name23353 (
		\wishbone_tx_fifo_fifo_reg[7][3]/P0001 ,
		_w33054_,
		_w33865_
	);
	LUT2 #(
		.INIT('h8)
	) name23354 (
		\wishbone_tx_fifo_fifo_reg[4][3]/P0001 ,
		_w33064_,
		_w33866_
	);
	LUT2 #(
		.INIT('h8)
	) name23355 (
		\wishbone_tx_fifo_fifo_reg[14][3]/P0001 ,
		_w33050_,
		_w33867_
	);
	LUT2 #(
		.INIT('h8)
	) name23356 (
		\wishbone_tx_fifo_fifo_reg[1][3]/P0001 ,
		_w33060_,
		_w33868_
	);
	LUT2 #(
		.INIT('h8)
	) name23357 (
		\wishbone_tx_fifo_fifo_reg[2][3]/P0001 ,
		_w33068_,
		_w33869_
	);
	LUT2 #(
		.INIT('h1)
	) name23358 (
		_w33855_,
		_w33856_,
		_w33870_
	);
	LUT2 #(
		.INIT('h1)
	) name23359 (
		_w33857_,
		_w33858_,
		_w33871_
	);
	LUT2 #(
		.INIT('h1)
	) name23360 (
		_w33859_,
		_w33860_,
		_w33872_
	);
	LUT2 #(
		.INIT('h1)
	) name23361 (
		_w33861_,
		_w33862_,
		_w33873_
	);
	LUT2 #(
		.INIT('h1)
	) name23362 (
		_w33863_,
		_w33864_,
		_w33874_
	);
	LUT2 #(
		.INIT('h1)
	) name23363 (
		_w33865_,
		_w33866_,
		_w33875_
	);
	LUT2 #(
		.INIT('h1)
	) name23364 (
		_w33867_,
		_w33868_,
		_w33876_
	);
	LUT2 #(
		.INIT('h4)
	) name23365 (
		_w33869_,
		_w33876_,
		_w33877_
	);
	LUT2 #(
		.INIT('h8)
	) name23366 (
		_w33874_,
		_w33875_,
		_w33878_
	);
	LUT2 #(
		.INIT('h8)
	) name23367 (
		_w33872_,
		_w33873_,
		_w33879_
	);
	LUT2 #(
		.INIT('h8)
	) name23368 (
		_w33870_,
		_w33871_,
		_w33880_
	);
	LUT2 #(
		.INIT('h8)
	) name23369 (
		_w33879_,
		_w33880_,
		_w33881_
	);
	LUT2 #(
		.INIT('h8)
	) name23370 (
		_w33877_,
		_w33878_,
		_w33882_
	);
	LUT2 #(
		.INIT('h8)
	) name23371 (
		_w33881_,
		_w33882_,
		_w33883_
	);
	LUT2 #(
		.INIT('h2)
	) name23372 (
		_w33028_,
		_w33883_,
		_w33884_
	);
	LUT2 #(
		.INIT('h1)
	) name23373 (
		_w33854_,
		_w33884_,
		_w33885_
	);
	LUT2 #(
		.INIT('h2)
	) name23374 (
		\wishbone_tx_fifo_fifo_reg[0][4]/P0001 ,
		_w33032_,
		_w33886_
	);
	LUT2 #(
		.INIT('h8)
	) name23375 (
		\wishbone_tx_fifo_fifo_reg[3][4]/P0001 ,
		_w33062_,
		_w33887_
	);
	LUT2 #(
		.INIT('h8)
	) name23376 (
		\wishbone_tx_fifo_fifo_reg[5][4]/P0001 ,
		_w33040_,
		_w33888_
	);
	LUT2 #(
		.INIT('h8)
	) name23377 (
		\wishbone_tx_fifo_fifo_reg[15][4]/P0001 ,
		_w33045_,
		_w33889_
	);
	LUT2 #(
		.INIT('h8)
	) name23378 (
		\wishbone_tx_fifo_fifo_reg[2][4]/P0001 ,
		_w33068_,
		_w33890_
	);
	LUT2 #(
		.INIT('h8)
	) name23379 (
		\wishbone_tx_fifo_fifo_reg[13][4]/P0001 ,
		_w33047_,
		_w33891_
	);
	LUT2 #(
		.INIT('h8)
	) name23380 (
		\wishbone_tx_fifo_fifo_reg[6][4]/P0001 ,
		_w33056_,
		_w33892_
	);
	LUT2 #(
		.INIT('h8)
	) name23381 (
		\wishbone_tx_fifo_fifo_reg[8][4]/P0001 ,
		_w33042_,
		_w33893_
	);
	LUT2 #(
		.INIT('h8)
	) name23382 (
		\wishbone_tx_fifo_fifo_reg[14][4]/P0001 ,
		_w33050_,
		_w33894_
	);
	LUT2 #(
		.INIT('h8)
	) name23383 (
		\wishbone_tx_fifo_fifo_reg[7][4]/P0001 ,
		_w33054_,
		_w33895_
	);
	LUT2 #(
		.INIT('h8)
	) name23384 (
		\wishbone_tx_fifo_fifo_reg[10][4]/P0001 ,
		_w33066_,
		_w33896_
	);
	LUT2 #(
		.INIT('h8)
	) name23385 (
		\wishbone_tx_fifo_fifo_reg[11][4]/P0001 ,
		_w33036_,
		_w33897_
	);
	LUT2 #(
		.INIT('h8)
	) name23386 (
		\wishbone_tx_fifo_fifo_reg[12][4]/P0001 ,
		_w33058_,
		_w33898_
	);
	LUT2 #(
		.INIT('h8)
	) name23387 (
		\wishbone_tx_fifo_fifo_reg[4][4]/P0001 ,
		_w33064_,
		_w33899_
	);
	LUT2 #(
		.INIT('h8)
	) name23388 (
		\wishbone_tx_fifo_fifo_reg[9][4]/P0001 ,
		_w33052_,
		_w33900_
	);
	LUT2 #(
		.INIT('h8)
	) name23389 (
		\wishbone_tx_fifo_fifo_reg[1][4]/P0001 ,
		_w33060_,
		_w33901_
	);
	LUT2 #(
		.INIT('h1)
	) name23390 (
		_w33887_,
		_w33888_,
		_w33902_
	);
	LUT2 #(
		.INIT('h1)
	) name23391 (
		_w33889_,
		_w33890_,
		_w33903_
	);
	LUT2 #(
		.INIT('h1)
	) name23392 (
		_w33891_,
		_w33892_,
		_w33904_
	);
	LUT2 #(
		.INIT('h1)
	) name23393 (
		_w33893_,
		_w33894_,
		_w33905_
	);
	LUT2 #(
		.INIT('h1)
	) name23394 (
		_w33895_,
		_w33896_,
		_w33906_
	);
	LUT2 #(
		.INIT('h1)
	) name23395 (
		_w33897_,
		_w33898_,
		_w33907_
	);
	LUT2 #(
		.INIT('h1)
	) name23396 (
		_w33899_,
		_w33900_,
		_w33908_
	);
	LUT2 #(
		.INIT('h4)
	) name23397 (
		_w33901_,
		_w33908_,
		_w33909_
	);
	LUT2 #(
		.INIT('h8)
	) name23398 (
		_w33906_,
		_w33907_,
		_w33910_
	);
	LUT2 #(
		.INIT('h8)
	) name23399 (
		_w33904_,
		_w33905_,
		_w33911_
	);
	LUT2 #(
		.INIT('h8)
	) name23400 (
		_w33902_,
		_w33903_,
		_w33912_
	);
	LUT2 #(
		.INIT('h8)
	) name23401 (
		_w33911_,
		_w33912_,
		_w33913_
	);
	LUT2 #(
		.INIT('h8)
	) name23402 (
		_w33909_,
		_w33910_,
		_w33914_
	);
	LUT2 #(
		.INIT('h8)
	) name23403 (
		_w33913_,
		_w33914_,
		_w33915_
	);
	LUT2 #(
		.INIT('h2)
	) name23404 (
		_w33028_,
		_w33915_,
		_w33916_
	);
	LUT2 #(
		.INIT('h1)
	) name23405 (
		_w33886_,
		_w33916_,
		_w33917_
	);
	LUT2 #(
		.INIT('h2)
	) name23406 (
		\wishbone_tx_fifo_fifo_reg[0][5]/P0001 ,
		_w33032_,
		_w33918_
	);
	LUT2 #(
		.INIT('h8)
	) name23407 (
		\wishbone_tx_fifo_fifo_reg[3][5]/P0001 ,
		_w33062_,
		_w33919_
	);
	LUT2 #(
		.INIT('h8)
	) name23408 (
		\wishbone_tx_fifo_fifo_reg[9][5]/P0001 ,
		_w33052_,
		_w33920_
	);
	LUT2 #(
		.INIT('h8)
	) name23409 (
		\wishbone_tx_fifo_fifo_reg[5][5]/P0001 ,
		_w33040_,
		_w33921_
	);
	LUT2 #(
		.INIT('h8)
	) name23410 (
		\wishbone_tx_fifo_fifo_reg[7][5]/P0001 ,
		_w33054_,
		_w33922_
	);
	LUT2 #(
		.INIT('h8)
	) name23411 (
		\wishbone_tx_fifo_fifo_reg[10][5]/P0001 ,
		_w33066_,
		_w33923_
	);
	LUT2 #(
		.INIT('h8)
	) name23412 (
		\wishbone_tx_fifo_fifo_reg[6][5]/P0001 ,
		_w33056_,
		_w33924_
	);
	LUT2 #(
		.INIT('h8)
	) name23413 (
		\wishbone_tx_fifo_fifo_reg[12][5]/P0001 ,
		_w33058_,
		_w33925_
	);
	LUT2 #(
		.INIT('h8)
	) name23414 (
		\wishbone_tx_fifo_fifo_reg[4][5]/P0001 ,
		_w33064_,
		_w33926_
	);
	LUT2 #(
		.INIT('h8)
	) name23415 (
		\wishbone_tx_fifo_fifo_reg[1][5]/P0001 ,
		_w33060_,
		_w33927_
	);
	LUT2 #(
		.INIT('h8)
	) name23416 (
		\wishbone_tx_fifo_fifo_reg[13][5]/P0001 ,
		_w33047_,
		_w33928_
	);
	LUT2 #(
		.INIT('h8)
	) name23417 (
		\wishbone_tx_fifo_fifo_reg[2][5]/P0001 ,
		_w33068_,
		_w33929_
	);
	LUT2 #(
		.INIT('h8)
	) name23418 (
		\wishbone_tx_fifo_fifo_reg[14][5]/P0001 ,
		_w33050_,
		_w33930_
	);
	LUT2 #(
		.INIT('h8)
	) name23419 (
		\wishbone_tx_fifo_fifo_reg[8][5]/P0001 ,
		_w33042_,
		_w33931_
	);
	LUT2 #(
		.INIT('h8)
	) name23420 (
		\wishbone_tx_fifo_fifo_reg[11][5]/P0001 ,
		_w33036_,
		_w33932_
	);
	LUT2 #(
		.INIT('h8)
	) name23421 (
		\wishbone_tx_fifo_fifo_reg[15][5]/P0001 ,
		_w33045_,
		_w33933_
	);
	LUT2 #(
		.INIT('h1)
	) name23422 (
		_w33919_,
		_w33920_,
		_w33934_
	);
	LUT2 #(
		.INIT('h1)
	) name23423 (
		_w33921_,
		_w33922_,
		_w33935_
	);
	LUT2 #(
		.INIT('h1)
	) name23424 (
		_w33923_,
		_w33924_,
		_w33936_
	);
	LUT2 #(
		.INIT('h1)
	) name23425 (
		_w33925_,
		_w33926_,
		_w33937_
	);
	LUT2 #(
		.INIT('h1)
	) name23426 (
		_w33927_,
		_w33928_,
		_w33938_
	);
	LUT2 #(
		.INIT('h1)
	) name23427 (
		_w33929_,
		_w33930_,
		_w33939_
	);
	LUT2 #(
		.INIT('h1)
	) name23428 (
		_w33931_,
		_w33932_,
		_w33940_
	);
	LUT2 #(
		.INIT('h4)
	) name23429 (
		_w33933_,
		_w33940_,
		_w33941_
	);
	LUT2 #(
		.INIT('h8)
	) name23430 (
		_w33938_,
		_w33939_,
		_w33942_
	);
	LUT2 #(
		.INIT('h8)
	) name23431 (
		_w33936_,
		_w33937_,
		_w33943_
	);
	LUT2 #(
		.INIT('h8)
	) name23432 (
		_w33934_,
		_w33935_,
		_w33944_
	);
	LUT2 #(
		.INIT('h8)
	) name23433 (
		_w33943_,
		_w33944_,
		_w33945_
	);
	LUT2 #(
		.INIT('h8)
	) name23434 (
		_w33941_,
		_w33942_,
		_w33946_
	);
	LUT2 #(
		.INIT('h8)
	) name23435 (
		_w33945_,
		_w33946_,
		_w33947_
	);
	LUT2 #(
		.INIT('h2)
	) name23436 (
		_w33028_,
		_w33947_,
		_w33948_
	);
	LUT2 #(
		.INIT('h1)
	) name23437 (
		_w33918_,
		_w33948_,
		_w33949_
	);
	LUT2 #(
		.INIT('h2)
	) name23438 (
		\wishbone_tx_fifo_fifo_reg[0][6]/P0001 ,
		_w33032_,
		_w33950_
	);
	LUT2 #(
		.INIT('h8)
	) name23439 (
		\wishbone_tx_fifo_fifo_reg[12][6]/P0001 ,
		_w33058_,
		_w33951_
	);
	LUT2 #(
		.INIT('h8)
	) name23440 (
		\wishbone_tx_fifo_fifo_reg[5][6]/P0001 ,
		_w33040_,
		_w33952_
	);
	LUT2 #(
		.INIT('h8)
	) name23441 (
		\wishbone_tx_fifo_fifo_reg[14][6]/P0001 ,
		_w33050_,
		_w33953_
	);
	LUT2 #(
		.INIT('h8)
	) name23442 (
		\wishbone_tx_fifo_fifo_reg[3][6]/P0001 ,
		_w33062_,
		_w33954_
	);
	LUT2 #(
		.INIT('h8)
	) name23443 (
		\wishbone_tx_fifo_fifo_reg[9][6]/P0001 ,
		_w33052_,
		_w33955_
	);
	LUT2 #(
		.INIT('h8)
	) name23444 (
		\wishbone_tx_fifo_fifo_reg[6][6]/P0001 ,
		_w33056_,
		_w33956_
	);
	LUT2 #(
		.INIT('h8)
	) name23445 (
		\wishbone_tx_fifo_fifo_reg[2][6]/P0001 ,
		_w33068_,
		_w33957_
	);
	LUT2 #(
		.INIT('h8)
	) name23446 (
		\wishbone_tx_fifo_fifo_reg[1][6]/P0001 ,
		_w33060_,
		_w33958_
	);
	LUT2 #(
		.INIT('h8)
	) name23447 (
		\wishbone_tx_fifo_fifo_reg[4][6]/P0001 ,
		_w33064_,
		_w33959_
	);
	LUT2 #(
		.INIT('h8)
	) name23448 (
		\wishbone_tx_fifo_fifo_reg[11][6]/P0001 ,
		_w33036_,
		_w33960_
	);
	LUT2 #(
		.INIT('h8)
	) name23449 (
		\wishbone_tx_fifo_fifo_reg[15][6]/P0001 ,
		_w33045_,
		_w33961_
	);
	LUT2 #(
		.INIT('h8)
	) name23450 (
		\wishbone_tx_fifo_fifo_reg[13][6]/P0001 ,
		_w33047_,
		_w33962_
	);
	LUT2 #(
		.INIT('h8)
	) name23451 (
		\wishbone_tx_fifo_fifo_reg[10][6]/P0001 ,
		_w33066_,
		_w33963_
	);
	LUT2 #(
		.INIT('h8)
	) name23452 (
		\wishbone_tx_fifo_fifo_reg[8][6]/P0001 ,
		_w33042_,
		_w33964_
	);
	LUT2 #(
		.INIT('h8)
	) name23453 (
		\wishbone_tx_fifo_fifo_reg[7][6]/P0001 ,
		_w33054_,
		_w33965_
	);
	LUT2 #(
		.INIT('h1)
	) name23454 (
		_w33951_,
		_w33952_,
		_w33966_
	);
	LUT2 #(
		.INIT('h1)
	) name23455 (
		_w33953_,
		_w33954_,
		_w33967_
	);
	LUT2 #(
		.INIT('h1)
	) name23456 (
		_w33955_,
		_w33956_,
		_w33968_
	);
	LUT2 #(
		.INIT('h1)
	) name23457 (
		_w33957_,
		_w33958_,
		_w33969_
	);
	LUT2 #(
		.INIT('h1)
	) name23458 (
		_w33959_,
		_w33960_,
		_w33970_
	);
	LUT2 #(
		.INIT('h1)
	) name23459 (
		_w33961_,
		_w33962_,
		_w33971_
	);
	LUT2 #(
		.INIT('h1)
	) name23460 (
		_w33963_,
		_w33964_,
		_w33972_
	);
	LUT2 #(
		.INIT('h4)
	) name23461 (
		_w33965_,
		_w33972_,
		_w33973_
	);
	LUT2 #(
		.INIT('h8)
	) name23462 (
		_w33970_,
		_w33971_,
		_w33974_
	);
	LUT2 #(
		.INIT('h8)
	) name23463 (
		_w33968_,
		_w33969_,
		_w33975_
	);
	LUT2 #(
		.INIT('h8)
	) name23464 (
		_w33966_,
		_w33967_,
		_w33976_
	);
	LUT2 #(
		.INIT('h8)
	) name23465 (
		_w33975_,
		_w33976_,
		_w33977_
	);
	LUT2 #(
		.INIT('h8)
	) name23466 (
		_w33973_,
		_w33974_,
		_w33978_
	);
	LUT2 #(
		.INIT('h8)
	) name23467 (
		_w33977_,
		_w33978_,
		_w33979_
	);
	LUT2 #(
		.INIT('h2)
	) name23468 (
		_w33028_,
		_w33979_,
		_w33980_
	);
	LUT2 #(
		.INIT('h1)
	) name23469 (
		_w33950_,
		_w33980_,
		_w33981_
	);
	LUT2 #(
		.INIT('h2)
	) name23470 (
		\wishbone_tx_fifo_fifo_reg[0][7]/P0001 ,
		_w33032_,
		_w33982_
	);
	LUT2 #(
		.INIT('h8)
	) name23471 (
		\wishbone_tx_fifo_fifo_reg[9][7]/P0001 ,
		_w33052_,
		_w33983_
	);
	LUT2 #(
		.INIT('h8)
	) name23472 (
		\wishbone_tx_fifo_fifo_reg[14][7]/P0001 ,
		_w33050_,
		_w33984_
	);
	LUT2 #(
		.INIT('h8)
	) name23473 (
		\wishbone_tx_fifo_fifo_reg[10][7]/P0001 ,
		_w33066_,
		_w33985_
	);
	LUT2 #(
		.INIT('h8)
	) name23474 (
		\wishbone_tx_fifo_fifo_reg[15][7]/P0001 ,
		_w33045_,
		_w33986_
	);
	LUT2 #(
		.INIT('h8)
	) name23475 (
		\wishbone_tx_fifo_fifo_reg[6][7]/P0001 ,
		_w33056_,
		_w33987_
	);
	LUT2 #(
		.INIT('h8)
	) name23476 (
		\wishbone_tx_fifo_fifo_reg[1][7]/P0001 ,
		_w33060_,
		_w33988_
	);
	LUT2 #(
		.INIT('h8)
	) name23477 (
		\wishbone_tx_fifo_fifo_reg[11][7]/P0001 ,
		_w33036_,
		_w33989_
	);
	LUT2 #(
		.INIT('h8)
	) name23478 (
		\wishbone_tx_fifo_fifo_reg[4][7]/P0001 ,
		_w33064_,
		_w33990_
	);
	LUT2 #(
		.INIT('h8)
	) name23479 (
		\wishbone_tx_fifo_fifo_reg[13][7]/P0001 ,
		_w33047_,
		_w33991_
	);
	LUT2 #(
		.INIT('h8)
	) name23480 (
		\wishbone_tx_fifo_fifo_reg[5][7]/P0001 ,
		_w33040_,
		_w33992_
	);
	LUT2 #(
		.INIT('h8)
	) name23481 (
		\wishbone_tx_fifo_fifo_reg[7][7]/P0001 ,
		_w33054_,
		_w33993_
	);
	LUT2 #(
		.INIT('h8)
	) name23482 (
		\wishbone_tx_fifo_fifo_reg[12][7]/P0001 ,
		_w33058_,
		_w33994_
	);
	LUT2 #(
		.INIT('h8)
	) name23483 (
		\wishbone_tx_fifo_fifo_reg[8][7]/P0001 ,
		_w33042_,
		_w33995_
	);
	LUT2 #(
		.INIT('h8)
	) name23484 (
		\wishbone_tx_fifo_fifo_reg[2][7]/P0001 ,
		_w33068_,
		_w33996_
	);
	LUT2 #(
		.INIT('h8)
	) name23485 (
		\wishbone_tx_fifo_fifo_reg[3][7]/P0001 ,
		_w33062_,
		_w33997_
	);
	LUT2 #(
		.INIT('h1)
	) name23486 (
		_w33983_,
		_w33984_,
		_w33998_
	);
	LUT2 #(
		.INIT('h1)
	) name23487 (
		_w33985_,
		_w33986_,
		_w33999_
	);
	LUT2 #(
		.INIT('h1)
	) name23488 (
		_w33987_,
		_w33988_,
		_w34000_
	);
	LUT2 #(
		.INIT('h1)
	) name23489 (
		_w33989_,
		_w33990_,
		_w34001_
	);
	LUT2 #(
		.INIT('h1)
	) name23490 (
		_w33991_,
		_w33992_,
		_w34002_
	);
	LUT2 #(
		.INIT('h1)
	) name23491 (
		_w33993_,
		_w33994_,
		_w34003_
	);
	LUT2 #(
		.INIT('h1)
	) name23492 (
		_w33995_,
		_w33996_,
		_w34004_
	);
	LUT2 #(
		.INIT('h4)
	) name23493 (
		_w33997_,
		_w34004_,
		_w34005_
	);
	LUT2 #(
		.INIT('h8)
	) name23494 (
		_w34002_,
		_w34003_,
		_w34006_
	);
	LUT2 #(
		.INIT('h8)
	) name23495 (
		_w34000_,
		_w34001_,
		_w34007_
	);
	LUT2 #(
		.INIT('h8)
	) name23496 (
		_w33998_,
		_w33999_,
		_w34008_
	);
	LUT2 #(
		.INIT('h8)
	) name23497 (
		_w34007_,
		_w34008_,
		_w34009_
	);
	LUT2 #(
		.INIT('h8)
	) name23498 (
		_w34005_,
		_w34006_,
		_w34010_
	);
	LUT2 #(
		.INIT('h8)
	) name23499 (
		_w34009_,
		_w34010_,
		_w34011_
	);
	LUT2 #(
		.INIT('h2)
	) name23500 (
		_w33028_,
		_w34011_,
		_w34012_
	);
	LUT2 #(
		.INIT('h1)
	) name23501 (
		_w33982_,
		_w34012_,
		_w34013_
	);
	LUT2 #(
		.INIT('h2)
	) name23502 (
		\wishbone_tx_fifo_fifo_reg[0][8]/P0001 ,
		_w33032_,
		_w34014_
	);
	LUT2 #(
		.INIT('h8)
	) name23503 (
		\wishbone_tx_fifo_fifo_reg[9][8]/P0001 ,
		_w33052_,
		_w34015_
	);
	LUT2 #(
		.INIT('h8)
	) name23504 (
		\wishbone_tx_fifo_fifo_reg[3][8]/P0001 ,
		_w33062_,
		_w34016_
	);
	LUT2 #(
		.INIT('h8)
	) name23505 (
		\wishbone_tx_fifo_fifo_reg[6][8]/P0001 ,
		_w33056_,
		_w34017_
	);
	LUT2 #(
		.INIT('h8)
	) name23506 (
		\wishbone_tx_fifo_fifo_reg[15][8]/P0001 ,
		_w33045_,
		_w34018_
	);
	LUT2 #(
		.INIT('h8)
	) name23507 (
		\wishbone_tx_fifo_fifo_reg[8][8]/P0001 ,
		_w33042_,
		_w34019_
	);
	LUT2 #(
		.INIT('h8)
	) name23508 (
		\wishbone_tx_fifo_fifo_reg[5][8]/P0001 ,
		_w33040_,
		_w34020_
	);
	LUT2 #(
		.INIT('h8)
	) name23509 (
		\wishbone_tx_fifo_fifo_reg[13][8]/P0001 ,
		_w33047_,
		_w34021_
	);
	LUT2 #(
		.INIT('h8)
	) name23510 (
		\wishbone_tx_fifo_fifo_reg[4][8]/P0001 ,
		_w33064_,
		_w34022_
	);
	LUT2 #(
		.INIT('h8)
	) name23511 (
		\wishbone_tx_fifo_fifo_reg[14][8]/P0001 ,
		_w33050_,
		_w34023_
	);
	LUT2 #(
		.INIT('h8)
	) name23512 (
		\wishbone_tx_fifo_fifo_reg[12][8]/P0001 ,
		_w33058_,
		_w34024_
	);
	LUT2 #(
		.INIT('h8)
	) name23513 (
		\wishbone_tx_fifo_fifo_reg[7][8]/P0001 ,
		_w33054_,
		_w34025_
	);
	LUT2 #(
		.INIT('h8)
	) name23514 (
		\wishbone_tx_fifo_fifo_reg[2][8]/P0001 ,
		_w33068_,
		_w34026_
	);
	LUT2 #(
		.INIT('h8)
	) name23515 (
		\wishbone_tx_fifo_fifo_reg[1][8]/P0001 ,
		_w33060_,
		_w34027_
	);
	LUT2 #(
		.INIT('h8)
	) name23516 (
		\wishbone_tx_fifo_fifo_reg[10][8]/P0001 ,
		_w33066_,
		_w34028_
	);
	LUT2 #(
		.INIT('h8)
	) name23517 (
		\wishbone_tx_fifo_fifo_reg[11][8]/P0001 ,
		_w33036_,
		_w34029_
	);
	LUT2 #(
		.INIT('h1)
	) name23518 (
		_w34015_,
		_w34016_,
		_w34030_
	);
	LUT2 #(
		.INIT('h1)
	) name23519 (
		_w34017_,
		_w34018_,
		_w34031_
	);
	LUT2 #(
		.INIT('h1)
	) name23520 (
		_w34019_,
		_w34020_,
		_w34032_
	);
	LUT2 #(
		.INIT('h1)
	) name23521 (
		_w34021_,
		_w34022_,
		_w34033_
	);
	LUT2 #(
		.INIT('h1)
	) name23522 (
		_w34023_,
		_w34024_,
		_w34034_
	);
	LUT2 #(
		.INIT('h1)
	) name23523 (
		_w34025_,
		_w34026_,
		_w34035_
	);
	LUT2 #(
		.INIT('h1)
	) name23524 (
		_w34027_,
		_w34028_,
		_w34036_
	);
	LUT2 #(
		.INIT('h4)
	) name23525 (
		_w34029_,
		_w34036_,
		_w34037_
	);
	LUT2 #(
		.INIT('h8)
	) name23526 (
		_w34034_,
		_w34035_,
		_w34038_
	);
	LUT2 #(
		.INIT('h8)
	) name23527 (
		_w34032_,
		_w34033_,
		_w34039_
	);
	LUT2 #(
		.INIT('h8)
	) name23528 (
		_w34030_,
		_w34031_,
		_w34040_
	);
	LUT2 #(
		.INIT('h8)
	) name23529 (
		_w34039_,
		_w34040_,
		_w34041_
	);
	LUT2 #(
		.INIT('h8)
	) name23530 (
		_w34037_,
		_w34038_,
		_w34042_
	);
	LUT2 #(
		.INIT('h8)
	) name23531 (
		_w34041_,
		_w34042_,
		_w34043_
	);
	LUT2 #(
		.INIT('h2)
	) name23532 (
		_w33028_,
		_w34043_,
		_w34044_
	);
	LUT2 #(
		.INIT('h1)
	) name23533 (
		_w34014_,
		_w34044_,
		_w34045_
	);
	LUT2 #(
		.INIT('h2)
	) name23534 (
		\wishbone_tx_fifo_fifo_reg[0][9]/P0001 ,
		_w33032_,
		_w34046_
	);
	LUT2 #(
		.INIT('h8)
	) name23535 (
		\wishbone_tx_fifo_fifo_reg[11][9]/P0001 ,
		_w33036_,
		_w34047_
	);
	LUT2 #(
		.INIT('h8)
	) name23536 (
		\wishbone_tx_fifo_fifo_reg[5][9]/P0001 ,
		_w33040_,
		_w34048_
	);
	LUT2 #(
		.INIT('h8)
	) name23537 (
		\wishbone_tx_fifo_fifo_reg[8][9]/P0001 ,
		_w33042_,
		_w34049_
	);
	LUT2 #(
		.INIT('h8)
	) name23538 (
		\wishbone_tx_fifo_fifo_reg[15][9]/P0001 ,
		_w33045_,
		_w34050_
	);
	LUT2 #(
		.INIT('h8)
	) name23539 (
		\wishbone_tx_fifo_fifo_reg[13][9]/P0001 ,
		_w33047_,
		_w34051_
	);
	LUT2 #(
		.INIT('h8)
	) name23540 (
		\wishbone_tx_fifo_fifo_reg[14][9]/P0001 ,
		_w33050_,
		_w34052_
	);
	LUT2 #(
		.INIT('h8)
	) name23541 (
		\wishbone_tx_fifo_fifo_reg[9][9]/P0001 ,
		_w33052_,
		_w34053_
	);
	LUT2 #(
		.INIT('h8)
	) name23542 (
		\wishbone_tx_fifo_fifo_reg[7][9]/P0001 ,
		_w33054_,
		_w34054_
	);
	LUT2 #(
		.INIT('h8)
	) name23543 (
		\wishbone_tx_fifo_fifo_reg[6][9]/P0001 ,
		_w33056_,
		_w34055_
	);
	LUT2 #(
		.INIT('h8)
	) name23544 (
		\wishbone_tx_fifo_fifo_reg[12][9]/P0001 ,
		_w33058_,
		_w34056_
	);
	LUT2 #(
		.INIT('h8)
	) name23545 (
		\wishbone_tx_fifo_fifo_reg[1][9]/P0001 ,
		_w33060_,
		_w34057_
	);
	LUT2 #(
		.INIT('h8)
	) name23546 (
		\wishbone_tx_fifo_fifo_reg[3][9]/P0001 ,
		_w33062_,
		_w34058_
	);
	LUT2 #(
		.INIT('h8)
	) name23547 (
		\wishbone_tx_fifo_fifo_reg[4][9]/P0001 ,
		_w33064_,
		_w34059_
	);
	LUT2 #(
		.INIT('h8)
	) name23548 (
		\wishbone_tx_fifo_fifo_reg[10][9]/P0001 ,
		_w33066_,
		_w34060_
	);
	LUT2 #(
		.INIT('h8)
	) name23549 (
		\wishbone_tx_fifo_fifo_reg[2][9]/P0001 ,
		_w33068_,
		_w34061_
	);
	LUT2 #(
		.INIT('h1)
	) name23550 (
		_w34047_,
		_w34048_,
		_w34062_
	);
	LUT2 #(
		.INIT('h1)
	) name23551 (
		_w34049_,
		_w34050_,
		_w34063_
	);
	LUT2 #(
		.INIT('h1)
	) name23552 (
		_w34051_,
		_w34052_,
		_w34064_
	);
	LUT2 #(
		.INIT('h1)
	) name23553 (
		_w34053_,
		_w34054_,
		_w34065_
	);
	LUT2 #(
		.INIT('h1)
	) name23554 (
		_w34055_,
		_w34056_,
		_w34066_
	);
	LUT2 #(
		.INIT('h1)
	) name23555 (
		_w34057_,
		_w34058_,
		_w34067_
	);
	LUT2 #(
		.INIT('h1)
	) name23556 (
		_w34059_,
		_w34060_,
		_w34068_
	);
	LUT2 #(
		.INIT('h4)
	) name23557 (
		_w34061_,
		_w34068_,
		_w34069_
	);
	LUT2 #(
		.INIT('h8)
	) name23558 (
		_w34066_,
		_w34067_,
		_w34070_
	);
	LUT2 #(
		.INIT('h8)
	) name23559 (
		_w34064_,
		_w34065_,
		_w34071_
	);
	LUT2 #(
		.INIT('h8)
	) name23560 (
		_w34062_,
		_w34063_,
		_w34072_
	);
	LUT2 #(
		.INIT('h8)
	) name23561 (
		_w34071_,
		_w34072_,
		_w34073_
	);
	LUT2 #(
		.INIT('h8)
	) name23562 (
		_w34069_,
		_w34070_,
		_w34074_
	);
	LUT2 #(
		.INIT('h8)
	) name23563 (
		_w34073_,
		_w34074_,
		_w34075_
	);
	LUT2 #(
		.INIT('h2)
	) name23564 (
		_w33028_,
		_w34075_,
		_w34076_
	);
	LUT2 #(
		.INIT('h1)
	) name23565 (
		_w34046_,
		_w34076_,
		_w34077_
	);
	LUT2 #(
		.INIT('h8)
	) name23566 (
		\wishbone_tx_burst_cnt_reg[1]/NET0131 ,
		_w31359_,
		_w34078_
	);
	LUT2 #(
		.INIT('h1)
	) name23567 (
		_w12574_,
		_w31360_,
		_w34079_
	);
	LUT2 #(
		.INIT('h8)
	) name23568 (
		_w12561_,
		_w34079_,
		_w34080_
	);
	LUT2 #(
		.INIT('h1)
	) name23569 (
		_w34078_,
		_w34080_,
		_w34081_
	);
	LUT2 #(
		.INIT('h8)
	) name23570 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w34082_
	);
	LUT2 #(
		.INIT('h8)
	) name23571 (
		_w31365_,
		_w34082_,
		_w34083_
	);
	LUT2 #(
		.INIT('h2)
	) name23572 (
		_w12657_,
		_w34083_,
		_w34084_
	);
	LUT2 #(
		.INIT('h2)
	) name23573 (
		\wishbone_ReadTxDataFromFifo_sync2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_sync3_reg/NET0131 ,
		_w34085_
	);
	LUT2 #(
		.INIT('h1)
	) name23574 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w34086_
	);
	LUT2 #(
		.INIT('h4)
	) name23575 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w34086_,
		_w34087_
	);
	LUT2 #(
		.INIT('h1)
	) name23576 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w34088_
	);
	LUT2 #(
		.INIT('h8)
	) name23577 (
		_w34087_,
		_w34088_,
		_w34089_
	);
	LUT2 #(
		.INIT('h2)
	) name23578 (
		_w34085_,
		_w34089_,
		_w34090_
	);
	LUT2 #(
		.INIT('h2)
	) name23579 (
		_w12657_,
		_w34090_,
		_w34091_
	);
	LUT2 #(
		.INIT('h4)
	) name23580 (
		_w12657_,
		_w34090_,
		_w34092_
	);
	LUT2 #(
		.INIT('h1)
	) name23581 (
		_w34091_,
		_w34092_,
		_w34093_
	);
	LUT2 #(
		.INIT('h4)
	) name23582 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w34087_,
		_w34094_
	);
	LUT2 #(
		.INIT('h2)
	) name23583 (
		_w34085_,
		_w34094_,
		_w34095_
	);
	LUT2 #(
		.INIT('h1)
	) name23584 (
		_w34084_,
		_w34095_,
		_w34096_
	);
	LUT2 #(
		.INIT('h4)
	) name23585 (
		_w34093_,
		_w34096_,
		_w34097_
	);
	LUT2 #(
		.INIT('h8)
	) name23586 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w34097_,
		_w34098_
	);
	LUT2 #(
		.INIT('h1)
	) name23587 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w34097_,
		_w34099_
	);
	LUT2 #(
		.INIT('h2)
	) name23588 (
		_w33028_,
		_w34098_,
		_w34100_
	);
	LUT2 #(
		.INIT('h4)
	) name23589 (
		_w34099_,
		_w34100_,
		_w34101_
	);
	LUT2 #(
		.INIT('h8)
	) name23590 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\wishbone_RxStatusWriteLatched_sync2_reg/NET0131 ,
		_w34102_
	);
	LUT2 #(
		.INIT('h1)
	) name23591 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		_w31730_,
		_w34103_
	);
	LUT2 #(
		.INIT('h1)
	) name23592 (
		_w12532_,
		_w34102_,
		_w34104_
	);
	LUT2 #(
		.INIT('h4)
	) name23593 (
		_w34103_,
		_w34104_,
		_w34105_
	);
	LUT2 #(
		.INIT('h4)
	) name23594 (
		mdc_pad_o_pad,
		_w31208_,
		_w34106_
	);
	LUT2 #(
		.INIT('h2)
	) name23595 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w34106_,
		_w34107_
	);
	LUT2 #(
		.INIT('h8)
	) name23596 (
		_w31410_,
		_w34106_,
		_w34108_
	);
	LUT2 #(
		.INIT('h8)
	) name23597 (
		\miim1_InProgress_reg/NET0131 ,
		_w34106_,
		_w34109_
	);
	LUT2 #(
		.INIT('h8)
	) name23598 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[1]/NET0131 ,
		_w34110_
	);
	LUT2 #(
		.INIT('h8)
	) name23599 (
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w34110_,
		_w34111_
	);
	LUT2 #(
		.INIT('h8)
	) name23600 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w34111_,
		_w34112_
	);
	LUT2 #(
		.INIT('h8)
	) name23601 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w34112_,
		_w34113_
	);
	LUT2 #(
		.INIT('h1)
	) name23602 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w34113_,
		_w34114_
	);
	LUT2 #(
		.INIT('h8)
	) name23603 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w34113_,
		_w34115_
	);
	LUT2 #(
		.INIT('h1)
	) name23604 (
		_w34114_,
		_w34115_,
		_w34116_
	);
	LUT2 #(
		.INIT('h8)
	) name23605 (
		_w34109_,
		_w34116_,
		_w34117_
	);
	LUT2 #(
		.INIT('h1)
	) name23606 (
		_w34107_,
		_w34108_,
		_w34118_
	);
	LUT2 #(
		.INIT('h4)
	) name23607 (
		_w34117_,
		_w34118_,
		_w34119_
	);
	LUT2 #(
		.INIT('h4)
	) name23608 (
		_w12621_,
		_w31329_,
		_w34120_
	);
	LUT2 #(
		.INIT('h8)
	) name23609 (
		\wishbone_rx_burst_en_reg/NET0131 ,
		_w34120_,
		_w34121_
	);
	LUT2 #(
		.INIT('h8)
	) name23610 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		_w34122_
	);
	LUT2 #(
		.INIT('h4)
	) name23611 (
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w34122_,
		_w34123_
	);
	LUT2 #(
		.INIT('h2)
	) name23612 (
		_w12621_,
		_w34123_,
		_w34124_
	);
	LUT2 #(
		.INIT('h8)
	) name23613 (
		\wishbone_MasterWbRX_reg/NET0131 ,
		_w12551_,
		_w34125_
	);
	LUT2 #(
		.INIT('h2)
	) name23614 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w34125_,
		_w34126_
	);
	LUT2 #(
		.INIT('h2)
	) name23615 (
		_w12553_,
		_w34126_,
		_w34127_
	);
	LUT2 #(
		.INIT('h1)
	) name23616 (
		_w31329_,
		_w34127_,
		_w34128_
	);
	LUT2 #(
		.INIT('h1)
	) name23617 (
		_w34124_,
		_w34128_,
		_w34129_
	);
	LUT2 #(
		.INIT('h4)
	) name23618 (
		_w34121_,
		_w34129_,
		_w34130_
	);
	LUT2 #(
		.INIT('h8)
	) name23619 (
		_w12552_,
		_w15698_,
		_w34131_
	);
	LUT2 #(
		.INIT('h1)
	) name23620 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w34131_,
		_w34132_
	);
	LUT2 #(
		.INIT('h2)
	) name23621 (
		\wishbone_WriteRxDataToFifoSync2_reg/NET0131 ,
		\wishbone_WriteRxDataToFifoSync3_reg/NET0131 ,
		_w34133_
	);
	LUT2 #(
		.INIT('h4)
	) name23622 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w34134_
	);
	LUT2 #(
		.INIT('h8)
	) name23623 (
		_w12552_,
		_w34134_,
		_w34135_
	);
	LUT2 #(
		.INIT('h2)
	) name23624 (
		_w34133_,
		_w34135_,
		_w34136_
	);
	LUT2 #(
		.INIT('h2)
	) name23625 (
		_w15698_,
		_w34136_,
		_w34137_
	);
	LUT2 #(
		.INIT('h4)
	) name23626 (
		_w15698_,
		_w34136_,
		_w34138_
	);
	LUT2 #(
		.INIT('h1)
	) name23627 (
		_w34137_,
		_w34138_,
		_w34139_
	);
	LUT2 #(
		.INIT('h8)
	) name23628 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w34140_
	);
	LUT2 #(
		.INIT('h2)
	) name23629 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w15698_,
		_w34141_
	);
	LUT2 #(
		.INIT('h8)
	) name23630 (
		_w34140_,
		_w34141_,
		_w34142_
	);
	LUT2 #(
		.INIT('h2)
	) name23631 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w34142_,
		_w34143_
	);
	LUT2 #(
		.INIT('h1)
	) name23632 (
		_w34132_,
		_w34143_,
		_w34144_
	);
	LUT2 #(
		.INIT('h4)
	) name23633 (
		_w34139_,
		_w34144_,
		_w34145_
	);
	LUT2 #(
		.INIT('h1)
	) name23634 (
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w34145_,
		_w34146_
	);
	LUT2 #(
		.INIT('h8)
	) name23635 (
		\wishbone_rx_fifo_cnt_reg[4]/NET0131 ,
		_w34145_,
		_w34147_
	);
	LUT2 #(
		.INIT('h1)
	) name23636 (
		_w31950_,
		_w34146_,
		_w34148_
	);
	LUT2 #(
		.INIT('h4)
	) name23637 (
		_w34147_,
		_w34148_,
		_w34149_
	);
	LUT2 #(
		.INIT('h1)
	) name23638 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w34150_
	);
	LUT2 #(
		.INIT('h8)
	) name23639 (
		\rxethmac1_RxValid_reg/NET0131 ,
		_w34150_,
		_w34151_
	);
	LUT2 #(
		.INIT('h8)
	) name23640 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		_w34151_,
		_w34152_
	);
	LUT2 #(
		.INIT('h8)
	) name23641 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34152_,
		_w34153_
	);
	LUT2 #(
		.INIT('h1)
	) name23642 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34152_,
		_w34154_
	);
	LUT2 #(
		.INIT('h1)
	) name23643 (
		_w31346_,
		_w34153_,
		_w34155_
	);
	LUT2 #(
		.INIT('h4)
	) name23644 (
		_w34154_,
		_w34155_,
		_w34156_
	);
	LUT2 #(
		.INIT('h1)
	) name23645 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		_w34151_,
		_w34157_
	);
	LUT2 #(
		.INIT('h1)
	) name23646 (
		_w31346_,
		_w34152_,
		_w34158_
	);
	LUT2 #(
		.INIT('h4)
	) name23647 (
		_w34157_,
		_w34158_,
		_w34159_
	);
	LUT2 #(
		.INIT('h1)
	) name23648 (
		\maccontrol1_receivecontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		_w34153_,
		_w34160_
	);
	LUT2 #(
		.INIT('h1)
	) name23649 (
		_w31346_,
		_w34160_,
		_w34161_
	);
	LUT2 #(
		.INIT('h4)
	) name23650 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w34162_
	);
	LUT2 #(
		.INIT('h4)
	) name23651 (
		\txethmac1_txcrc_Crc_reg[28]/NET0131 ,
		_w34162_,
		_w34163_
	);
	LUT2 #(
		.INIT('h1)
	) name23652 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		\txethmac1_txstatem1_StateFCS_reg/NET0131 ,
		_w34164_
	);
	LUT2 #(
		.INIT('h1)
	) name23653 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w11071_,
		_w34165_
	);
	LUT2 #(
		.INIT('h2)
	) name23654 (
		_w34164_,
		_w34165_,
		_w34166_
	);
	LUT2 #(
		.INIT('h1)
	) name23655 (
		_w34163_,
		_w34166_,
		_w34167_
	);
	LUT2 #(
		.INIT('h1)
	) name23656 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w34167_,
		_w34168_
	);
	LUT2 #(
		.INIT('h2)
	) name23657 (
		_w11295_,
		_w34168_,
		_w34169_
	);
	LUT2 #(
		.INIT('h2)
	) name23658 (
		\txethmac1_txcrc_Crc_reg[1]/NET0131 ,
		_w12472_,
		_w34170_
	);
	LUT2 #(
		.INIT('h4)
	) name23659 (
		\txethmac1_txcrc_Crc_reg[1]/NET0131 ,
		_w12472_,
		_w34171_
	);
	LUT2 #(
		.INIT('h2)
	) name23660 (
		_w11181_,
		_w34170_,
		_w34172_
	);
	LUT2 #(
		.INIT('h4)
	) name23661 (
		_w34171_,
		_w34172_,
		_w34173_
	);
	LUT2 #(
		.INIT('h2)
	) name23662 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w15136_,
		_w34174_
	);
	LUT2 #(
		.INIT('h2)
	) name23663 (
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w15135_,
		_w34175_
	);
	LUT2 #(
		.INIT('h8)
	) name23664 (
		_w31214_,
		_w34175_,
		_w34176_
	);
	LUT2 #(
		.INIT('h1)
	) name23665 (
		_w34174_,
		_w34176_,
		_w34177_
	);
	LUT2 #(
		.INIT('h1)
	) name23666 (
		\RxAbort_wb_reg/NET0131 ,
		_w34177_,
		_w34178_
	);
	LUT2 #(
		.INIT('h8)
	) name23667 (
		\rxethmac1_LatchedByte_reg[4]/NET0131 ,
		_w31852_,
		_w34179_
	);
	LUT2 #(
		.INIT('h8)
	) name23668 (
		\rxethmac1_RxData_d_reg[4]/NET0131 ,
		_w31853_,
		_w34180_
	);
	LUT2 #(
		.INIT('h1)
	) name23669 (
		_w34179_,
		_w34180_,
		_w34181_
	);
	LUT2 #(
		.INIT('h4)
	) name23670 (
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w34115_,
		_w34182_
	);
	LUT2 #(
		.INIT('h1)
	) name23671 (
		\miim1_InProgress_q1_reg/NET0131 ,
		\miim1_InProgress_q2_reg/NET0131 ,
		_w34183_
	);
	LUT2 #(
		.INIT('h4)
	) name23672 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w34184_
	);
	LUT2 #(
		.INIT('h8)
	) name23673 (
		_w34183_,
		_w34184_,
		_w34185_
	);
	LUT2 #(
		.INIT('h2)
	) name23674 (
		\miim1_WCtrlDataStart_q1_reg/NET0131 ,
		\miim1_WCtrlDataStart_q2_reg/NET0131 ,
		_w34186_
	);
	LUT2 #(
		.INIT('h2)
	) name23675 (
		\miim1_RStatStart_q1_reg/NET0131 ,
		\miim1_RStatStart_q2_reg/NET0131 ,
		_w34187_
	);
	LUT2 #(
		.INIT('h1)
	) name23676 (
		_w34186_,
		_w34187_,
		_w34188_
	);
	LUT2 #(
		.INIT('h4)
	) name23677 (
		_w34185_,
		_w34188_,
		_w34189_
	);
	LUT2 #(
		.INIT('h4)
	) name23678 (
		_w34182_,
		_w34189_,
		_w34190_
	);
	LUT2 #(
		.INIT('h2)
	) name23679 (
		_w34106_,
		_w34190_,
		_w34191_
	);
	LUT2 #(
		.INIT('h2)
	) name23680 (
		\miim1_WriteOp_reg/NET0131 ,
		_w34191_,
		_w34192_
	);
	LUT2 #(
		.INIT('h2)
	) name23681 (
		_w34106_,
		_w34189_,
		_w34193_
	);
	LUT2 #(
		.INIT('h2)
	) name23682 (
		\miim1_InProgress_reg/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w34194_
	);
	LUT2 #(
		.INIT('h1)
	) name23683 (
		\miim1_InProgress_reg/NET0131 ,
		_w34186_,
		_w34195_
	);
	LUT2 #(
		.INIT('h1)
	) name23684 (
		_w34194_,
		_w34195_,
		_w34196_
	);
	LUT2 #(
		.INIT('h8)
	) name23685 (
		_w34193_,
		_w34196_,
		_w34197_
	);
	LUT2 #(
		.INIT('h1)
	) name23686 (
		_w34192_,
		_w34197_,
		_w34198_
	);
	LUT2 #(
		.INIT('h2)
	) name23687 (
		\ethreg1_MODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w34199_
	);
	LUT2 #(
		.INIT('h4)
	) name23688 (
		\wishbone_r_RxEn_q_reg/NET0131 ,
		_w34199_,
		_w34200_
	);
	LUT2 #(
		.INIT('h8)
	) name23689 (
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w15175_,
		_w34201_
	);
	LUT2 #(
		.INIT('h1)
	) name23690 (
		_w34200_,
		_w34201_,
		_w34202_
	);
	LUT2 #(
		.INIT('h1)
	) name23691 (
		\wishbone_RxStatus_reg[13]/NET0131 ,
		_w34200_,
		_w34203_
	);
	LUT2 #(
		.INIT('h1)
	) name23692 (
		_w34202_,
		_w34203_,
		_w34204_
	);
	LUT2 #(
		.INIT('h8)
	) name23693 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w34204_,
		_w34205_
	);
	LUT2 #(
		.INIT('h8)
	) name23694 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w34206_
	);
	LUT2 #(
		.INIT('h8)
	) name23695 (
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w34206_,
		_w34207_
	);
	LUT2 #(
		.INIT('h8)
	) name23696 (
		_w34201_,
		_w34207_,
		_w34208_
	);
	LUT2 #(
		.INIT('h1)
	) name23697 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		_w34208_,
		_w34209_
	);
	LUT2 #(
		.INIT('h8)
	) name23698 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		_w34208_,
		_w34210_
	);
	LUT2 #(
		.INIT('h1)
	) name23699 (
		_w34204_,
		_w34209_,
		_w34211_
	);
	LUT2 #(
		.INIT('h4)
	) name23700 (
		_w34210_,
		_w34211_,
		_w34212_
	);
	LUT2 #(
		.INIT('h1)
	) name23701 (
		_w34205_,
		_w34212_,
		_w34213_
	);
	LUT2 #(
		.INIT('h4)
	) name23702 (
		\wishbone_ShiftWillEnd_reg/NET0131 ,
		_w31349_,
		_w34214_
	);
	LUT2 #(
		.INIT('h2)
	) name23703 (
		_w31212_,
		_w34214_,
		_w34215_
	);
	LUT2 #(
		.INIT('h2)
	) name23704 (
		\miim1_BitCounter_reg[1]/NET0131 ,
		_w34106_,
		_w34216_
	);
	LUT2 #(
		.INIT('h4)
	) name23705 (
		_w31409_,
		_w34109_,
		_w34217_
	);
	LUT2 #(
		.INIT('h1)
	) name23706 (
		_w31403_,
		_w34110_,
		_w34218_
	);
	LUT2 #(
		.INIT('h8)
	) name23707 (
		_w34217_,
		_w34218_,
		_w34219_
	);
	LUT2 #(
		.INIT('h1)
	) name23708 (
		_w34216_,
		_w34219_,
		_w34220_
	);
	LUT2 #(
		.INIT('h2)
	) name23709 (
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w34106_,
		_w34221_
	);
	LUT2 #(
		.INIT('h1)
	) name23710 (
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w34110_,
		_w34222_
	);
	LUT2 #(
		.INIT('h1)
	) name23711 (
		_w34111_,
		_w34222_,
		_w34223_
	);
	LUT2 #(
		.INIT('h8)
	) name23712 (
		_w34217_,
		_w34223_,
		_w34224_
	);
	LUT2 #(
		.INIT('h1)
	) name23713 (
		_w34221_,
		_w34224_,
		_w34225_
	);
	LUT2 #(
		.INIT('h2)
	) name23714 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w34106_,
		_w34226_
	);
	LUT2 #(
		.INIT('h1)
	) name23715 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w34111_,
		_w34227_
	);
	LUT2 #(
		.INIT('h1)
	) name23716 (
		_w34112_,
		_w34227_,
		_w34228_
	);
	LUT2 #(
		.INIT('h8)
	) name23717 (
		_w34217_,
		_w34228_,
		_w34229_
	);
	LUT2 #(
		.INIT('h1)
	) name23718 (
		_w34226_,
		_w34229_,
		_w34230_
	);
	LUT2 #(
		.INIT('h2)
	) name23719 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w34106_,
		_w34231_
	);
	LUT2 #(
		.INIT('h1)
	) name23720 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		_w34112_,
		_w34232_
	);
	LUT2 #(
		.INIT('h1)
	) name23721 (
		_w34113_,
		_w34232_,
		_w34233_
	);
	LUT2 #(
		.INIT('h8)
	) name23722 (
		_w34217_,
		_w34233_,
		_w34234_
	);
	LUT2 #(
		.INIT('h1)
	) name23723 (
		_w34231_,
		_w34234_,
		_w34235_
	);
	LUT2 #(
		.INIT('h2)
	) name23724 (
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w34106_,
		_w34236_
	);
	LUT2 #(
		.INIT('h2)
	) name23725 (
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w34115_,
		_w34237_
	);
	LUT2 #(
		.INIT('h1)
	) name23726 (
		_w34182_,
		_w34237_,
		_w34238_
	);
	LUT2 #(
		.INIT('h2)
	) name23727 (
		_w34217_,
		_w34238_,
		_w34239_
	);
	LUT2 #(
		.INIT('h1)
	) name23728 (
		_w34236_,
		_w34239_,
		_w34240_
	);
	LUT2 #(
		.INIT('h2)
	) name23729 (
		\miim1_clkgen_Counter_reg[6]/NET0131 ,
		_w31207_,
		_w34241_
	);
	LUT2 #(
		.INIT('h4)
	) name23730 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		_w31206_,
		_w34242_
	);
	LUT2 #(
		.INIT('h1)
	) name23731 (
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w34242_,
		_w34243_
	);
	LUT2 #(
		.INIT('h8)
	) name23732 (
		\ethreg1_MIIMODER_0_DataOut_reg[7]/NET0131 ,
		_w34242_,
		_w34244_
	);
	LUT2 #(
		.INIT('h2)
	) name23733 (
		_w31208_,
		_w34243_,
		_w34245_
	);
	LUT2 #(
		.INIT('h4)
	) name23734 (
		_w34244_,
		_w34245_,
		_w34246_
	);
	LUT2 #(
		.INIT('h1)
	) name23735 (
		_w34241_,
		_w34246_,
		_w34247_
	);
	LUT2 #(
		.INIT('h8)
	) name23736 (
		\rxethmac1_Multicast_reg/NET0131 ,
		_w12477_,
		_w34248_
	);
	LUT2 #(
		.INIT('h8)
	) name23737 (
		\rxethmac1_LatchedByte_reg[0]/NET0131 ,
		_w12484_,
		_w34249_
	);
	LUT2 #(
		.INIT('h1)
	) name23738 (
		_w34248_,
		_w34249_,
		_w34250_
	);
	LUT2 #(
		.INIT('h1)
	) name23739 (
		\maccontrol1_receivecontrol1_DetectionWindow_reg/NET0131 ,
		\macstatus1_ReceiveEnd_reg/NET0131 ,
		_w34251_
	);
	LUT2 #(
		.INIT('h1)
	) name23740 (
		_w31227_,
		_w34251_,
		_w34252_
	);
	LUT2 #(
		.INIT('h2)
	) name23741 (
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		_w10659_,
		_w34253_
	);
	LUT2 #(
		.INIT('h4)
	) name23742 (
		\rxethmac1_crcrx_Crc_reg[13]/NET0131 ,
		_w10659_,
		_w34254_
	);
	LUT2 #(
		.INIT('h2)
	) name23743 (
		_w10580_,
		_w34253_,
		_w34255_
	);
	LUT2 #(
		.INIT('h4)
	) name23744 (
		_w34254_,
		_w34255_,
		_w34256_
	);
	LUT2 #(
		.INIT('h1)
	) name23745 (
		\txethmac1_TxAbort_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w34257_
	);
	LUT2 #(
		.INIT('h1)
	) name23746 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w34257_,
		_w34258_
	);
	LUT2 #(
		.INIT('h1)
	) name23747 (
		wb_rst_i_pad,
		_w34258_,
		_w34259_
	);
	LUT2 #(
		.INIT('h4)
	) name23748 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_q_reg/P0001 ,
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w34260_
	);
	LUT2 #(
		.INIT('h1)
	) name23749 (
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w34260_,
		_w34261_
	);
	LUT2 #(
		.INIT('h1)
	) name23750 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w34262_
	);
	LUT2 #(
		.INIT('h8)
	) name23751 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34262_,
		_w34263_
	);
	LUT2 #(
		.INIT('h4)
	) name23752 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w34264_
	);
	LUT2 #(
		.INIT('h4)
	) name23753 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34264_,
		_w34265_
	);
	LUT2 #(
		.INIT('h8)
	) name23754 (
		_w34263_,
		_w34265_,
		_w34266_
	);
	LUT2 #(
		.INIT('h8)
	) name23755 (
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w34266_,
		_w34267_
	);
	LUT2 #(
		.INIT('h8)
	) name23756 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34268_
	);
	LUT2 #(
		.INIT('h2)
	) name23757 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w34268_,
		_w34269_
	);
	LUT2 #(
		.INIT('h2)
	) name23758 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w34269_,
		_w34270_
	);
	LUT2 #(
		.INIT('h4)
	) name23759 (
		_w34261_,
		_w34270_,
		_w34271_
	);
	LUT2 #(
		.INIT('h4)
	) name23760 (
		_w34267_,
		_w34271_,
		_w34272_
	);
	LUT2 #(
		.INIT('h8)
	) name23761 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w34272_,
		_w34273_
	);
	LUT2 #(
		.INIT('h8)
	) name23762 (
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w34260_,
		_w34274_
	);
	LUT2 #(
		.INIT('h8)
	) name23763 (
		_w34270_,
		_w34274_,
		_w34275_
	);
	LUT2 #(
		.INIT('h1)
	) name23764 (
		_w34273_,
		_w34275_,
		_w34276_
	);
	LUT2 #(
		.INIT('h2)
	) name23765 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w34276_,
		_w34277_
	);
	LUT2 #(
		.INIT('h8)
	) name23766 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34277_,
		_w34278_
	);
	LUT2 #(
		.INIT('h1)
	) name23767 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		_w34278_,
		_w34279_
	);
	LUT2 #(
		.INIT('h8)
	) name23768 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		_w34278_,
		_w34280_
	);
	LUT2 #(
		.INIT('h2)
	) name23769 (
		_w34259_,
		_w34279_,
		_w34281_
	);
	LUT2 #(
		.INIT('h4)
	) name23770 (
		_w34280_,
		_w34281_,
		_w34282_
	);
	LUT2 #(
		.INIT('h4)
	) name23771 (
		\wishbone_LatchValidBytes_q_reg/NET0131 ,
		\wishbone_LatchValidBytes_reg/NET0131 ,
		_w34283_
	);
	LUT2 #(
		.INIT('h8)
	) name23772 (
		_w13499_,
		_w34283_,
		_w34284_
	);
	LUT2 #(
		.INIT('h8)
	) name23773 (
		\wishbone_TxLength_reg[0]/NET0131 ,
		_w34284_,
		_w34285_
	);
	LUT2 #(
		.INIT('h4)
	) name23774 (
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w34286_
	);
	LUT2 #(
		.INIT('h4)
	) name23775 (
		\wishbone_TxAbort_wb_q_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w34287_
	);
	LUT2 #(
		.INIT('h4)
	) name23776 (
		\wishbone_TxRetry_wb_q_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w34288_
	);
	LUT2 #(
		.INIT('h1)
	) name23777 (
		_w34287_,
		_w34288_,
		_w34289_
	);
	LUT2 #(
		.INIT('h4)
	) name23778 (
		_w34286_,
		_w34289_,
		_w34290_
	);
	LUT2 #(
		.INIT('h4)
	) name23779 (
		_w34283_,
		_w34290_,
		_w34291_
	);
	LUT2 #(
		.INIT('h8)
	) name23780 (
		\wishbone_TxValidBytesLatched_reg[0]/NET0131 ,
		_w34291_,
		_w34292_
	);
	LUT2 #(
		.INIT('h1)
	) name23781 (
		_w34285_,
		_w34292_,
		_w34293_
	);
	LUT2 #(
		.INIT('h8)
	) name23782 (
		\wishbone_TxLength_reg[1]/NET0131 ,
		_w34284_,
		_w34294_
	);
	LUT2 #(
		.INIT('h8)
	) name23783 (
		\wishbone_TxValidBytesLatched_reg[1]/NET0131 ,
		_w34291_,
		_w34295_
	);
	LUT2 #(
		.INIT('h1)
	) name23784 (
		_w34294_,
		_w34295_,
		_w34296_
	);
	LUT2 #(
		.INIT('h2)
	) name23785 (
		_w11181_,
		_w12107_,
		_w34297_
	);
	LUT2 #(
		.INIT('h2)
	) name23786 (
		_w11181_,
		_w12210_,
		_w34298_
	);
	LUT2 #(
		.INIT('h4)
	) name23787 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		_w34109_,
		_w34299_
	);
	LUT2 #(
		.INIT('h2)
	) name23788 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		_w34106_,
		_w34300_
	);
	LUT2 #(
		.INIT('h1)
	) name23789 (
		_w34108_,
		_w34300_,
		_w34301_
	);
	LUT2 #(
		.INIT('h4)
	) name23790 (
		_w34299_,
		_w34301_,
		_w34302_
	);
	LUT2 #(
		.INIT('h1)
	) name23791 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w11222_,
		_w34303_
	);
	LUT2 #(
		.INIT('h8)
	) name23792 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w10683_,
		_w34304_
	);
	LUT2 #(
		.INIT('h1)
	) name23793 (
		_w11071_,
		_w34304_,
		_w34305_
	);
	LUT2 #(
		.INIT('h1)
	) name23794 (
		_w10684_,
		_w34305_,
		_w34306_
	);
	LUT2 #(
		.INIT('h1)
	) name23795 (
		_w11074_,
		_w34303_,
		_w34307_
	);
	LUT2 #(
		.INIT('h4)
	) name23796 (
		_w34306_,
		_w34307_,
		_w34308_
	);
	LUT2 #(
		.INIT('h8)
	) name23797 (
		_w34106_,
		_w34182_,
		_w34309_
	);
	LUT2 #(
		.INIT('h2)
	) name23798 (
		\miim1_InProgress_reg/NET0131 ,
		_w34309_,
		_w34310_
	);
	LUT2 #(
		.INIT('h1)
	) name23799 (
		_w34193_,
		_w34310_,
		_w34311_
	);
	LUT2 #(
		.INIT('h2)
	) name23800 (
		\ethreg1_MIIMODER_0_DataOut_reg[3]/NET0131 ,
		_w31202_,
		_w34312_
	);
	LUT2 #(
		.INIT('h4)
	) name23801 (
		_w31203_,
		_w31208_,
		_w34313_
	);
	LUT2 #(
		.INIT('h4)
	) name23802 (
		_w34312_,
		_w34313_,
		_w34314_
	);
	LUT2 #(
		.INIT('h2)
	) name23803 (
		\miim1_clkgen_Counter_reg[2]/NET0131 ,
		_w31190_,
		_w34315_
	);
	LUT2 #(
		.INIT('h1)
	) name23804 (
		_w31191_,
		_w34315_,
		_w34316_
	);
	LUT2 #(
		.INIT('h4)
	) name23805 (
		_w31208_,
		_w34316_,
		_w34317_
	);
	LUT2 #(
		.INIT('h1)
	) name23806 (
		_w34314_,
		_w34317_,
		_w34318_
	);
	LUT2 #(
		.INIT('h2)
	) name23807 (
		\miim1_LatchByte1_d_reg/NET0131 ,
		_w34106_,
		_w34319_
	);
	LUT2 #(
		.INIT('h8)
	) name23808 (
		\miim1_BitCounter_reg[1]/NET0131 ,
		\miim1_BitCounter_reg[2]/NET0131 ,
		_w34320_
	);
	LUT2 #(
		.INIT('h2)
	) name23809 (
		\miim1_BitCounter_reg[0]/NET0131 ,
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w34321_
	);
	LUT2 #(
		.INIT('h2)
	) name23810 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		\miim1_WriteOp_reg/NET0131 ,
		_w34322_
	);
	LUT2 #(
		.INIT('h8)
	) name23811 (
		_w34321_,
		_w34322_,
		_w34323_
	);
	LUT2 #(
		.INIT('h8)
	) name23812 (
		_w34320_,
		_w34323_,
		_w34324_
	);
	LUT2 #(
		.INIT('h8)
	) name23813 (
		_w31420_,
		_w34324_,
		_w34325_
	);
	LUT2 #(
		.INIT('h8)
	) name23814 (
		_w34106_,
		_w34325_,
		_w34326_
	);
	LUT2 #(
		.INIT('h1)
	) name23815 (
		_w34319_,
		_w34326_,
		_w34327_
	);
	LUT2 #(
		.INIT('h8)
	) name23816 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		_w34204_,
		_w34328_
	);
	LUT2 #(
		.INIT('h8)
	) name23817 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w34329_
	);
	LUT2 #(
		.INIT('h8)
	) name23818 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w34329_,
		_w34330_
	);
	LUT2 #(
		.INIT('h8)
	) name23819 (
		_w34208_,
		_w34330_,
		_w34331_
	);
	LUT2 #(
		.INIT('h1)
	) name23820 (
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w34331_,
		_w34332_
	);
	LUT2 #(
		.INIT('h8)
	) name23821 (
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w34331_,
		_w34333_
	);
	LUT2 #(
		.INIT('h1)
	) name23822 (
		_w34204_,
		_w34332_,
		_w34334_
	);
	LUT2 #(
		.INIT('h4)
	) name23823 (
		_w34333_,
		_w34334_,
		_w34335_
	);
	LUT2 #(
		.INIT('h1)
	) name23824 (
		_w34328_,
		_w34335_,
		_w34336_
	);
	LUT2 #(
		.INIT('h4)
	) name23825 (
		\wishbone_LastByteIn_reg/NET0131 ,
		_w31213_,
		_w34337_
	);
	LUT2 #(
		.INIT('h8)
	) name23826 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31239_,
		_w34338_
	);
	LUT2 #(
		.INIT('h1)
	) name23827 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w34339_
	);
	LUT2 #(
		.INIT('h8)
	) name23828 (
		_w31345_,
		_w34339_,
		_w34340_
	);
	LUT2 #(
		.INIT('h1)
	) name23829 (
		_w34338_,
		_w34340_,
		_w34341_
	);
	LUT2 #(
		.INIT('h2)
	) name23830 (
		_w34337_,
		_w34341_,
		_w34342_
	);
	LUT2 #(
		.INIT('h1)
	) name23831 (
		\wishbone_RxDataLatched1_reg[10]/NET0131 ,
		_w34342_,
		_w34343_
	);
	LUT2 #(
		.INIT('h4)
	) name23832 (
		\rxethmac1_RxData_reg[2]/NET0131 ,
		_w34337_,
		_w34344_
	);
	LUT2 #(
		.INIT('h4)
	) name23833 (
		_w34341_,
		_w34344_,
		_w34345_
	);
	LUT2 #(
		.INIT('h1)
	) name23834 (
		_w34343_,
		_w34345_,
		_w34346_
	);
	LUT2 #(
		.INIT('h1)
	) name23835 (
		\wishbone_RxDataLatched1_reg[11]/NET0131 ,
		_w34342_,
		_w34347_
	);
	LUT2 #(
		.INIT('h4)
	) name23836 (
		\rxethmac1_RxData_reg[3]/NET0131 ,
		_w34337_,
		_w34348_
	);
	LUT2 #(
		.INIT('h4)
	) name23837 (
		_w34341_,
		_w34348_,
		_w34349_
	);
	LUT2 #(
		.INIT('h1)
	) name23838 (
		_w34347_,
		_w34349_,
		_w34350_
	);
	LUT2 #(
		.INIT('h1)
	) name23839 (
		\wishbone_RxDataLatched1_reg[12]/NET0131 ,
		_w34342_,
		_w34351_
	);
	LUT2 #(
		.INIT('h4)
	) name23840 (
		\rxethmac1_RxData_reg[4]/NET0131 ,
		_w34337_,
		_w34352_
	);
	LUT2 #(
		.INIT('h4)
	) name23841 (
		_w34341_,
		_w34352_,
		_w34353_
	);
	LUT2 #(
		.INIT('h1)
	) name23842 (
		_w34351_,
		_w34353_,
		_w34354_
	);
	LUT2 #(
		.INIT('h1)
	) name23843 (
		\wishbone_RxDataLatched1_reg[13]/NET0131 ,
		_w34342_,
		_w34355_
	);
	LUT2 #(
		.INIT('h4)
	) name23844 (
		\rxethmac1_RxData_reg[5]/NET0131 ,
		_w34337_,
		_w34356_
	);
	LUT2 #(
		.INIT('h4)
	) name23845 (
		_w34341_,
		_w34356_,
		_w34357_
	);
	LUT2 #(
		.INIT('h1)
	) name23846 (
		_w34355_,
		_w34357_,
		_w34358_
	);
	LUT2 #(
		.INIT('h1)
	) name23847 (
		\wishbone_RxDataLatched1_reg[14]/NET0131 ,
		_w34342_,
		_w34359_
	);
	LUT2 #(
		.INIT('h4)
	) name23848 (
		\rxethmac1_RxData_reg[6]/NET0131 ,
		_w34337_,
		_w34360_
	);
	LUT2 #(
		.INIT('h4)
	) name23849 (
		_w34341_,
		_w34360_,
		_w34361_
	);
	LUT2 #(
		.INIT('h1)
	) name23850 (
		_w34359_,
		_w34361_,
		_w34362_
	);
	LUT2 #(
		.INIT('h1)
	) name23851 (
		\wishbone_RxDataLatched1_reg[15]/NET0131 ,
		_w34342_,
		_w34363_
	);
	LUT2 #(
		.INIT('h4)
	) name23852 (
		\rxethmac1_RxData_reg[7]/NET0131 ,
		_w34337_,
		_w34364_
	);
	LUT2 #(
		.INIT('h4)
	) name23853 (
		_w34341_,
		_w34364_,
		_w34365_
	);
	LUT2 #(
		.INIT('h1)
	) name23854 (
		_w34363_,
		_w34365_,
		_w34366_
	);
	LUT2 #(
		.INIT('h8)
	) name23855 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31238_,
		_w34367_
	);
	LUT2 #(
		.INIT('h4)
	) name23856 (
		\wishbone_RxByteCnt_reg[1]/NET0131 ,
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w34368_
	);
	LUT2 #(
		.INIT('h4)
	) name23857 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_RxByteCnt_reg[0]/NET0131 ,
		_w34369_
	);
	LUT2 #(
		.INIT('h8)
	) name23858 (
		_w34368_,
		_w34369_,
		_w34370_
	);
	LUT2 #(
		.INIT('h1)
	) name23859 (
		_w34367_,
		_w34370_,
		_w34371_
	);
	LUT2 #(
		.INIT('h2)
	) name23860 (
		_w34337_,
		_w34371_,
		_w34372_
	);
	LUT2 #(
		.INIT('h1)
	) name23861 (
		\wishbone_RxDataLatched1_reg[16]/NET0131 ,
		_w34372_,
		_w34373_
	);
	LUT2 #(
		.INIT('h4)
	) name23862 (
		\rxethmac1_RxData_reg[0]/NET0131 ,
		_w34337_,
		_w34374_
	);
	LUT2 #(
		.INIT('h4)
	) name23863 (
		_w34371_,
		_w34374_,
		_w34375_
	);
	LUT2 #(
		.INIT('h1)
	) name23864 (
		_w34373_,
		_w34375_,
		_w34376_
	);
	LUT2 #(
		.INIT('h1)
	) name23865 (
		\wishbone_RxDataLatched1_reg[17]/NET0131 ,
		_w34372_,
		_w34377_
	);
	LUT2 #(
		.INIT('h4)
	) name23866 (
		\rxethmac1_RxData_reg[1]/NET0131 ,
		_w34337_,
		_w34378_
	);
	LUT2 #(
		.INIT('h4)
	) name23867 (
		_w34371_,
		_w34378_,
		_w34379_
	);
	LUT2 #(
		.INIT('h1)
	) name23868 (
		_w34377_,
		_w34379_,
		_w34380_
	);
	LUT2 #(
		.INIT('h1)
	) name23869 (
		\wishbone_RxDataLatched1_reg[18]/NET0131 ,
		_w34372_,
		_w34381_
	);
	LUT2 #(
		.INIT('h2)
	) name23870 (
		_w34344_,
		_w34371_,
		_w34382_
	);
	LUT2 #(
		.INIT('h1)
	) name23871 (
		_w34381_,
		_w34382_,
		_w34383_
	);
	LUT2 #(
		.INIT('h1)
	) name23872 (
		\wishbone_RxDataLatched1_reg[19]/NET0131 ,
		_w34372_,
		_w34384_
	);
	LUT2 #(
		.INIT('h2)
	) name23873 (
		_w34348_,
		_w34371_,
		_w34385_
	);
	LUT2 #(
		.INIT('h1)
	) name23874 (
		_w34384_,
		_w34385_,
		_w34386_
	);
	LUT2 #(
		.INIT('h1)
	) name23875 (
		\wishbone_RxDataLatched1_reg[20]/NET0131 ,
		_w34372_,
		_w34387_
	);
	LUT2 #(
		.INIT('h2)
	) name23876 (
		_w34352_,
		_w34371_,
		_w34388_
	);
	LUT2 #(
		.INIT('h1)
	) name23877 (
		_w34387_,
		_w34388_,
		_w34389_
	);
	LUT2 #(
		.INIT('h1)
	) name23878 (
		\wishbone_RxDataLatched1_reg[21]/NET0131 ,
		_w34372_,
		_w34390_
	);
	LUT2 #(
		.INIT('h2)
	) name23879 (
		_w34356_,
		_w34371_,
		_w34391_
	);
	LUT2 #(
		.INIT('h1)
	) name23880 (
		_w34390_,
		_w34391_,
		_w34392_
	);
	LUT2 #(
		.INIT('h1)
	) name23881 (
		\wishbone_RxDataLatched1_reg[22]/NET0131 ,
		_w34372_,
		_w34393_
	);
	LUT2 #(
		.INIT('h2)
	) name23882 (
		_w34360_,
		_w34371_,
		_w34394_
	);
	LUT2 #(
		.INIT('h1)
	) name23883 (
		_w34393_,
		_w34394_,
		_w34395_
	);
	LUT2 #(
		.INIT('h1)
	) name23884 (
		\wishbone_RxDataLatched1_reg[23]/NET0131 ,
		_w34372_,
		_w34396_
	);
	LUT2 #(
		.INIT('h2)
	) name23885 (
		_w34364_,
		_w34371_,
		_w34397_
	);
	LUT2 #(
		.INIT('h1)
	) name23886 (
		_w34396_,
		_w34397_,
		_w34398_
	);
	LUT2 #(
		.INIT('h8)
	) name23887 (
		_w34339_,
		_w34368_,
		_w34399_
	);
	LUT2 #(
		.INIT('h8)
	) name23888 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w31813_,
		_w34400_
	);
	LUT2 #(
		.INIT('h1)
	) name23889 (
		_w34399_,
		_w34400_,
		_w34401_
	);
	LUT2 #(
		.INIT('h2)
	) name23890 (
		_w34337_,
		_w34401_,
		_w34402_
	);
	LUT2 #(
		.INIT('h1)
	) name23891 (
		\wishbone_RxDataLatched1_reg[24]/NET0131 ,
		_w34402_,
		_w34403_
	);
	LUT2 #(
		.INIT('h2)
	) name23892 (
		_w34374_,
		_w34401_,
		_w34404_
	);
	LUT2 #(
		.INIT('h1)
	) name23893 (
		_w34403_,
		_w34404_,
		_w34405_
	);
	LUT2 #(
		.INIT('h1)
	) name23894 (
		\wishbone_RxDataLatched1_reg[25]/NET0131 ,
		_w34402_,
		_w34406_
	);
	LUT2 #(
		.INIT('h2)
	) name23895 (
		_w34378_,
		_w34401_,
		_w34407_
	);
	LUT2 #(
		.INIT('h1)
	) name23896 (
		_w34406_,
		_w34407_,
		_w34408_
	);
	LUT2 #(
		.INIT('h1)
	) name23897 (
		\wishbone_RxDataLatched1_reg[26]/NET0131 ,
		_w34402_,
		_w34409_
	);
	LUT2 #(
		.INIT('h2)
	) name23898 (
		_w34344_,
		_w34401_,
		_w34410_
	);
	LUT2 #(
		.INIT('h1)
	) name23899 (
		_w34409_,
		_w34410_,
		_w34411_
	);
	LUT2 #(
		.INIT('h1)
	) name23900 (
		\wishbone_RxDataLatched1_reg[27]/NET0131 ,
		_w34402_,
		_w34412_
	);
	LUT2 #(
		.INIT('h2)
	) name23901 (
		_w34348_,
		_w34401_,
		_w34413_
	);
	LUT2 #(
		.INIT('h1)
	) name23902 (
		_w34412_,
		_w34413_,
		_w34414_
	);
	LUT2 #(
		.INIT('h1)
	) name23903 (
		\wishbone_RxDataLatched1_reg[28]/NET0131 ,
		_w34402_,
		_w34415_
	);
	LUT2 #(
		.INIT('h2)
	) name23904 (
		_w34352_,
		_w34401_,
		_w34416_
	);
	LUT2 #(
		.INIT('h1)
	) name23905 (
		_w34415_,
		_w34416_,
		_w34417_
	);
	LUT2 #(
		.INIT('h1)
	) name23906 (
		\wishbone_RxDataLatched1_reg[29]/NET0131 ,
		_w34402_,
		_w34418_
	);
	LUT2 #(
		.INIT('h2)
	) name23907 (
		_w34356_,
		_w34401_,
		_w34419_
	);
	LUT2 #(
		.INIT('h1)
	) name23908 (
		_w34418_,
		_w34419_,
		_w34420_
	);
	LUT2 #(
		.INIT('h1)
	) name23909 (
		\wishbone_RxDataLatched1_reg[30]/NET0131 ,
		_w34402_,
		_w34421_
	);
	LUT2 #(
		.INIT('h2)
	) name23910 (
		_w34360_,
		_w34401_,
		_w34422_
	);
	LUT2 #(
		.INIT('h1)
	) name23911 (
		_w34421_,
		_w34422_,
		_w34423_
	);
	LUT2 #(
		.INIT('h1)
	) name23912 (
		\wishbone_RxDataLatched1_reg[31]/NET0131 ,
		_w34402_,
		_w34424_
	);
	LUT2 #(
		.INIT('h2)
	) name23913 (
		_w34364_,
		_w34401_,
		_w34425_
	);
	LUT2 #(
		.INIT('h1)
	) name23914 (
		_w34424_,
		_w34425_,
		_w34426_
	);
	LUT2 #(
		.INIT('h1)
	) name23915 (
		\wishbone_RxDataLatched1_reg[8]/NET0131 ,
		_w34342_,
		_w34427_
	);
	LUT2 #(
		.INIT('h4)
	) name23916 (
		_w34341_,
		_w34374_,
		_w34428_
	);
	LUT2 #(
		.INIT('h1)
	) name23917 (
		_w34427_,
		_w34428_,
		_w34429_
	);
	LUT2 #(
		.INIT('h1)
	) name23918 (
		\wishbone_RxDataLatched1_reg[9]/NET0131 ,
		_w34342_,
		_w34430_
	);
	LUT2 #(
		.INIT('h4)
	) name23919 (
		_w34341_,
		_w34378_,
		_w34431_
	);
	LUT2 #(
		.INIT('h1)
	) name23920 (
		_w34430_,
		_w34431_,
		_w34432_
	);
	LUT2 #(
		.INIT('h2)
	) name23921 (
		\miim1_LatchByte0_d_reg/NET0131 ,
		_w34106_,
		_w34433_
	);
	LUT2 #(
		.INIT('h8)
	) name23922 (
		_w34194_,
		_w34309_,
		_w34434_
	);
	LUT2 #(
		.INIT('h1)
	) name23923 (
		_w34433_,
		_w34434_,
		_w34435_
	);
	LUT2 #(
		.INIT('h8)
	) name23924 (
		\wishbone_rx_burst_cnt_reg[1]/NET0131 ,
		_w34120_,
		_w34436_
	);
	LUT2 #(
		.INIT('h1)
	) name23925 (
		_w12607_,
		_w34122_,
		_w34437_
	);
	LUT2 #(
		.INIT('h8)
	) name23926 (
		_w12621_,
		_w34437_,
		_w34438_
	);
	LUT2 #(
		.INIT('h1)
	) name23927 (
		_w34436_,
		_w34438_,
		_w34439_
	);
	LUT2 #(
		.INIT('h8)
	) name23928 (
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w34120_,
		_w34440_
	);
	LUT2 #(
		.INIT('h2)
	) name23929 (
		\wishbone_rx_burst_cnt_reg[2]/NET0131 ,
		_w34122_,
		_w34441_
	);
	LUT2 #(
		.INIT('h1)
	) name23930 (
		_w34123_,
		_w34441_,
		_w34442_
	);
	LUT2 #(
		.INIT('h2)
	) name23931 (
		_w12621_,
		_w34442_,
		_w34443_
	);
	LUT2 #(
		.INIT('h1)
	) name23932 (
		_w34440_,
		_w34443_,
		_w34444_
	);
	LUT2 #(
		.INIT('h4)
	) name23933 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34445_
	);
	LUT2 #(
		.INIT('h8)
	) name23934 (
		\wishbone_tx_fifo_cnt_reg[4]/NET0131 ,
		_w34094_,
		_w34446_
	);
	LUT2 #(
		.INIT('h2)
	) name23935 (
		_w12657_,
		_w34446_,
		_w34447_
	);
	LUT2 #(
		.INIT('h2)
	) name23936 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34448_
	);
	LUT2 #(
		.INIT('h8)
	) name23937 (
		_w34447_,
		_w34448_,
		_w34449_
	);
	LUT2 #(
		.INIT('h8)
	) name23938 (
		_w33028_,
		_w34449_,
		_w34450_
	);
	LUT2 #(
		.INIT('h8)
	) name23939 (
		_w34445_,
		_w34450_,
		_w34451_
	);
	LUT2 #(
		.INIT('h4)
	) name23940 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34452_
	);
	LUT2 #(
		.INIT('h8)
	) name23941 (
		_w34447_,
		_w34452_,
		_w34453_
	);
	LUT2 #(
		.INIT('h8)
	) name23942 (
		_w33028_,
		_w34453_,
		_w34454_
	);
	LUT2 #(
		.INIT('h8)
	) name23943 (
		_w34445_,
		_w34454_,
		_w34455_
	);
	LUT2 #(
		.INIT('h8)
	) name23944 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34456_
	);
	LUT2 #(
		.INIT('h8)
	) name23945 (
		_w34454_,
		_w34456_,
		_w34457_
	);
	LUT2 #(
		.INIT('h8)
	) name23946 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		_w34447_,
		_w34458_
	);
	LUT2 #(
		.INIT('h1)
	) name23947 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34459_
	);
	LUT2 #(
		.INIT('h8)
	) name23948 (
		_w34458_,
		_w34459_,
		_w34460_
	);
	LUT2 #(
		.INIT('h4)
	) name23949 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w33028_,
		_w34461_
	);
	LUT2 #(
		.INIT('h8)
	) name23950 (
		_w34460_,
		_w34461_,
		_w34462_
	);
	LUT2 #(
		.INIT('h1)
	) name23951 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34463_
	);
	LUT2 #(
		.INIT('h8)
	) name23952 (
		_w34450_,
		_w34463_,
		_w34464_
	);
	LUT2 #(
		.INIT('h2)
	) name23953 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34465_
	);
	LUT2 #(
		.INIT('h8)
	) name23954 (
		_w34450_,
		_w34465_,
		_w34466_
	);
	LUT2 #(
		.INIT('h8)
	) name23955 (
		_w34454_,
		_w34463_,
		_w34467_
	);
	LUT2 #(
		.INIT('h8)
	) name23956 (
		_w34454_,
		_w34465_,
		_w34468_
	);
	LUT2 #(
		.INIT('h8)
	) name23957 (
		_w34447_,
		_w34463_,
		_w34469_
	);
	LUT2 #(
		.INIT('h8)
	) name23958 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34470_
	);
	LUT2 #(
		.INIT('h8)
	) name23959 (
		_w33028_,
		_w34470_,
		_w34471_
	);
	LUT2 #(
		.INIT('h8)
	) name23960 (
		_w34469_,
		_w34471_,
		_w34472_
	);
	LUT2 #(
		.INIT('h8)
	) name23961 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		_w34458_,
		_w34473_
	);
	LUT2 #(
		.INIT('h8)
	) name23962 (
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34473_,
		_w34474_
	);
	LUT2 #(
		.INIT('h4)
	) name23963 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34474_,
		_w34475_
	);
	LUT2 #(
		.INIT('h8)
	) name23964 (
		_w33028_,
		_w34475_,
		_w34476_
	);
	LUT2 #(
		.INIT('h8)
	) name23965 (
		_w33028_,
		_w34459_,
		_w34477_
	);
	LUT2 #(
		.INIT('h8)
	) name23966 (
		_w34447_,
		_w34456_,
		_w34478_
	);
	LUT2 #(
		.INIT('h8)
	) name23967 (
		_w34477_,
		_w34478_,
		_w34479_
	);
	LUT2 #(
		.INIT('h1)
	) name23968 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		_w12621_,
		_w34480_
	);
	LUT2 #(
		.INIT('h2)
	) name23969 (
		\wishbone_rx_burst_cnt_reg[0]/NET0131 ,
		_w34120_,
		_w34481_
	);
	LUT2 #(
		.INIT('h1)
	) name23970 (
		_w34480_,
		_w34481_,
		_w34482_
	);
	LUT2 #(
		.INIT('h8)
	) name23971 (
		_w34087_,
		_w34090_,
		_w34483_
	);
	LUT2 #(
		.INIT('h8)
	) name23972 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w34082_,
		_w34484_
	);
	LUT2 #(
		.INIT('h4)
	) name23973 (
		_w34085_,
		_w34484_,
		_w34485_
	);
	LUT2 #(
		.INIT('h1)
	) name23974 (
		_w34483_,
		_w34485_,
		_w34486_
	);
	LUT2 #(
		.INIT('h1)
	) name23975 (
		_w34093_,
		_w34486_,
		_w34487_
	);
	LUT2 #(
		.INIT('h1)
	) name23976 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w34487_,
		_w34488_
	);
	LUT2 #(
		.INIT('h8)
	) name23977 (
		\wishbone_tx_fifo_cnt_reg[3]/NET0131 ,
		_w34487_,
		_w34489_
	);
	LUT2 #(
		.INIT('h2)
	) name23978 (
		_w33028_,
		_w34488_,
		_w34490_
	);
	LUT2 #(
		.INIT('h4)
	) name23979 (
		_w34489_,
		_w34490_,
		_w34491_
	);
	LUT2 #(
		.INIT('h4)
	) name23980 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w34276_,
		_w34492_
	);
	LUT2 #(
		.INIT('h2)
	) name23981 (
		_w34259_,
		_w34277_,
		_w34493_
	);
	LUT2 #(
		.INIT('h4)
	) name23982 (
		_w34492_,
		_w34493_,
		_w34494_
	);
	LUT2 #(
		.INIT('h1)
	) name23983 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34277_,
		_w34495_
	);
	LUT2 #(
		.INIT('h2)
	) name23984 (
		_w34259_,
		_w34278_,
		_w34496_
	);
	LUT2 #(
		.INIT('h4)
	) name23985 (
		_w34495_,
		_w34496_,
		_w34497_
	);
	LUT2 #(
		.INIT('h1)
	) name23986 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w34280_,
		_w34498_
	);
	LUT2 #(
		.INIT('h8)
	) name23987 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w34499_
	);
	LUT2 #(
		.INIT('h8)
	) name23988 (
		_w34278_,
		_w34499_,
		_w34500_
	);
	LUT2 #(
		.INIT('h2)
	) name23989 (
		_w34259_,
		_w34500_,
		_w34501_
	);
	LUT2 #(
		.INIT('h4)
	) name23990 (
		_w34498_,
		_w34501_,
		_w34502_
	);
	LUT2 #(
		.INIT('h2)
	) name23991 (
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w11179_,
		_w34503_
	);
	LUT2 #(
		.INIT('h1)
	) name23992 (
		_w11071_,
		_w34503_,
		_w34504_
	);
	LUT2 #(
		.INIT('h2)
	) name23993 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w34504_,
		_w34505_
	);
	LUT2 #(
		.INIT('h8)
	) name23994 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w34505_,
		_w34506_
	);
	LUT2 #(
		.INIT('h1)
	) name23995 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w34505_,
		_w34507_
	);
	LUT2 #(
		.INIT('h8)
	) name23996 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\txethmac1_txstatem1_StateData_reg[1]/NET0131 ,
		_w34508_
	);
	LUT2 #(
		.INIT('h8)
	) name23997 (
		_w11178_,
		_w34508_,
		_w34509_
	);
	LUT2 #(
		.INIT('h1)
	) name23998 (
		\txethmac1_PacketFinished_q_reg/NET0131 ,
		_w34509_,
		_w34510_
	);
	LUT2 #(
		.INIT('h4)
	) name23999 (
		_w11074_,
		_w34510_,
		_w34511_
	);
	LUT2 #(
		.INIT('h1)
	) name24000 (
		_w34506_,
		_w34507_,
		_w34512_
	);
	LUT2 #(
		.INIT('h8)
	) name24001 (
		_w34511_,
		_w34512_,
		_w34513_
	);
	LUT2 #(
		.INIT('h8)
	) name24002 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34506_,
		_w34514_
	);
	LUT2 #(
		.INIT('h1)
	) name24003 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w34514_,
		_w34515_
	);
	LUT2 #(
		.INIT('h8)
	) name24004 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w34514_,
		_w34516_
	);
	LUT2 #(
		.INIT('h2)
	) name24005 (
		_w34511_,
		_w34515_,
		_w34517_
	);
	LUT2 #(
		.INIT('h4)
	) name24006 (
		_w34516_,
		_w34517_,
		_w34518_
	);
	LUT2 #(
		.INIT('h1)
	) name24007 (
		_w34131_,
		_w34142_,
		_w34519_
	);
	LUT2 #(
		.INIT('h1)
	) name24008 (
		_w34139_,
		_w34519_,
		_w34520_
	);
	LUT2 #(
		.INIT('h1)
	) name24009 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w34520_,
		_w34521_
	);
	LUT2 #(
		.INIT('h8)
	) name24010 (
		\wishbone_rx_fifo_cnt_reg[3]/NET0131 ,
		_w34520_,
		_w34522_
	);
	LUT2 #(
		.INIT('h1)
	) name24011 (
		_w31950_,
		_w34521_,
		_w34523_
	);
	LUT2 #(
		.INIT('h4)
	) name24012 (
		_w34522_,
		_w34523_,
		_w34524_
	);
	LUT2 #(
		.INIT('h8)
	) name24013 (
		_w22963_,
		_w31684_,
		_w34525_
	);
	LUT2 #(
		.INIT('h8)
	) name24014 (
		_w31686_,
		_w34525_,
		_w34526_
	);
	LUT2 #(
		.INIT('h8)
	) name24015 (
		_w24728_,
		_w34526_,
		_w34527_
	);
	LUT2 #(
		.INIT('h1)
	) name24016 (
		\ethreg1_MIICOMMAND1_DataOut_reg[0]/NET0131 ,
		_w34527_,
		_w34528_
	);
	LUT2 #(
		.INIT('h4)
	) name24017 (
		\wb_dat_i[1]_pad ,
		_w34527_,
		_w34529_
	);
	LUT2 #(
		.INIT('h1)
	) name24018 (
		\miim1_RStatStart_reg/NET0131 ,
		_w34528_,
		_w34530_
	);
	LUT2 #(
		.INIT('h4)
	) name24019 (
		_w34529_,
		_w34530_,
		_w34531_
	);
	LUT2 #(
		.INIT('h1)
	) name24020 (
		\ethreg1_MIICOMMAND2_DataOut_reg[0]/NET0131 ,
		_w34527_,
		_w34532_
	);
	LUT2 #(
		.INIT('h4)
	) name24021 (
		\wb_dat_i[2]_pad ,
		_w34527_,
		_w34533_
	);
	LUT2 #(
		.INIT('h1)
	) name24022 (
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w34532_,
		_w34534_
	);
	LUT2 #(
		.INIT('h4)
	) name24023 (
		_w34533_,
		_w34534_,
		_w34535_
	);
	LUT2 #(
		.INIT('h2)
	) name24024 (
		_w34272_,
		_w34275_,
		_w34536_
	);
	LUT2 #(
		.INIT('h1)
	) name24025 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w34536_,
		_w34537_
	);
	LUT2 #(
		.INIT('h8)
	) name24026 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		_w34536_,
		_w34538_
	);
	LUT2 #(
		.INIT('h2)
	) name24027 (
		_w34259_,
		_w34537_,
		_w34539_
	);
	LUT2 #(
		.INIT('h4)
	) name24028 (
		_w34538_,
		_w34539_,
		_w34540_
	);
	LUT2 #(
		.INIT('h1)
	) name24029 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34500_,
		_w34541_
	);
	LUT2 #(
		.INIT('h8)
	) name24030 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34500_,
		_w34542_
	);
	LUT2 #(
		.INIT('h2)
	) name24031 (
		_w34259_,
		_w34541_,
		_w34543_
	);
	LUT2 #(
		.INIT('h4)
	) name24032 (
		_w34542_,
		_w34543_,
		_w34544_
	);
	LUT2 #(
		.INIT('h2)
	) name24033 (
		_w10861_,
		_w10926_,
		_w34545_
	);
	LUT2 #(
		.INIT('h1)
	) name24034 (
		_w34306_,
		_w34545_,
		_w34546_
	);
	LUT2 #(
		.INIT('h1)
	) name24035 (
		\txethmac1_txcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34506_,
		_w34547_
	);
	LUT2 #(
		.INIT('h2)
	) name24036 (
		_w34511_,
		_w34514_,
		_w34548_
	);
	LUT2 #(
		.INIT('h4)
	) name24037 (
		_w34547_,
		_w34548_,
		_w34549_
	);
	LUT2 #(
		.INIT('h4)
	) name24038 (
		\wishbone_TxLength_reg[4]/NET0131 ,
		_w31367_,
		_w34550_
	);
	LUT2 #(
		.INIT('h8)
	) name24039 (
		_w31370_,
		_w34550_,
		_w34551_
	);
	LUT2 #(
		.INIT('h1)
	) name24040 (
		_w34083_,
		_w34551_,
		_w34552_
	);
	LUT2 #(
		.INIT('h2)
	) name24041 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		_w34553_
	);
	LUT2 #(
		.INIT('h1)
	) name24042 (
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		\wishbone_cyc_cleared_reg/NET0131 ,
		_w34554_
	);
	LUT2 #(
		.INIT('h8)
	) name24043 (
		_w34553_,
		_w34554_,
		_w34555_
	);
	LUT2 #(
		.INIT('h4)
	) name24044 (
		_w34552_,
		_w34555_,
		_w34556_
	);
	LUT2 #(
		.INIT('h2)
	) name24045 (
		\wishbone_BlockReadTxDataFromMemory_reg/NET0131 ,
		\wishbone_TxDonePacket_reg/NET0131 ,
		_w34557_
	);
	LUT2 #(
		.INIT('h8)
	) name24046 (
		_w33028_,
		_w34557_,
		_w34558_
	);
	LUT2 #(
		.INIT('h4)
	) name24047 (
		_w34085_,
		_w34558_,
		_w34559_
	);
	LUT2 #(
		.INIT('h1)
	) name24048 (
		_w34556_,
		_w34559_,
		_w34560_
	);
	LUT2 #(
		.INIT('h2)
	) name24049 (
		\miim1_InProgress_q1_reg/NET0131 ,
		_w34106_,
		_w34561_
	);
	LUT2 #(
		.INIT('h1)
	) name24050 (
		_w34109_,
		_w34561_,
		_w34562_
	);
	LUT2 #(
		.INIT('h2)
	) name24051 (
		_w10526_,
		_w12133_,
		_w34563_
	);
	LUT2 #(
		.INIT('h2)
	) name24052 (
		_w11757_,
		_w34563_,
		_w34564_
	);
	LUT2 #(
		.INIT('h1)
	) name24053 (
		\rxethmac1_RxEndFrm_d_reg/NET0131 ,
		_w34564_,
		_w34565_
	);
	LUT2 #(
		.INIT('h8)
	) name24054 (
		\wb_adr_i[2]_pad ,
		_w34525_,
		_w34566_
	);
	LUT2 #(
		.INIT('h8)
	) name24055 (
		_w22958_,
		_w34566_,
		_w34567_
	);
	LUT2 #(
		.INIT('h8)
	) name24056 (
		\wb_dat_i[2]_pad ,
		_w34567_,
		_w34568_
	);
	LUT2 #(
		.INIT('h2)
	) name24057 (
		\ethreg1_irq_rxb_reg/NET0131 ,
		_w34568_,
		_w34569_
	);
	LUT2 #(
		.INIT('h1)
	) name24058 (
		\wishbone_RxB_IRQ_reg/NET0131 ,
		_w34569_,
		_w34570_
	);
	LUT2 #(
		.INIT('h8)
	) name24059 (
		\wb_dat_i[6]_pad ,
		_w34567_,
		_w34571_
	);
	LUT2 #(
		.INIT('h2)
	) name24060 (
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w34571_,
		_w34572_
	);
	LUT2 #(
		.INIT('h1)
	) name24061 (
		\ethreg1_SetRxCIrq_reg/NET0131 ,
		_w34572_,
		_w34573_
	);
	LUT2 #(
		.INIT('h8)
	) name24062 (
		\wb_dat_i[3]_pad ,
		_w34567_,
		_w34574_
	);
	LUT2 #(
		.INIT('h2)
	) name24063 (
		\ethreg1_irq_rxe_reg/NET0131 ,
		_w34574_,
		_w34575_
	);
	LUT2 #(
		.INIT('h1)
	) name24064 (
		\wishbone_RxE_IRQ_reg/NET0131 ,
		_w34575_,
		_w34576_
	);
	LUT2 #(
		.INIT('h8)
	) name24065 (
		\wb_dat_i[0]_pad ,
		_w34567_,
		_w34577_
	);
	LUT2 #(
		.INIT('h2)
	) name24066 (
		\ethreg1_irq_txb_reg/NET0131 ,
		_w34577_,
		_w34578_
	);
	LUT2 #(
		.INIT('h1)
	) name24067 (
		\wishbone_TxB_IRQ_reg/NET0131 ,
		_w34578_,
		_w34579_
	);
	LUT2 #(
		.INIT('h8)
	) name24068 (
		\wb_dat_i[5]_pad ,
		_w34567_,
		_w34580_
	);
	LUT2 #(
		.INIT('h2)
	) name24069 (
		\ethreg1_irq_txc_reg/NET0131 ,
		_w34580_,
		_w34581_
	);
	LUT2 #(
		.INIT('h1)
	) name24070 (
		\ethreg1_SetTxCIrq_reg/NET0131 ,
		_w34581_,
		_w34582_
	);
	LUT2 #(
		.INIT('h8)
	) name24071 (
		\wb_dat_i[1]_pad ,
		_w34567_,
		_w34583_
	);
	LUT2 #(
		.INIT('h2)
	) name24072 (
		\ethreg1_irq_txe_reg/NET0131 ,
		_w34583_,
		_w34584_
	);
	LUT2 #(
		.INIT('h1)
	) name24073 (
		\wishbone_TxE_IRQ_reg/NET0131 ,
		_w34584_,
		_w34585_
	);
	LUT2 #(
		.INIT('h2)
	) name24074 (
		_w11002_,
		_w11067_,
		_w34586_
	);
	LUT2 #(
		.INIT('h8)
	) name24075 (
		_w11074_,
		_w34586_,
		_w34587_
	);
	LUT2 #(
		.INIT('h1)
	) name24076 (
		\txethmac1_TxRetry_reg/NET0131 ,
		_w34587_,
		_w34588_
	);
	LUT2 #(
		.INIT('h1)
	) name24077 (
		_w11388_,
		_w34588_,
		_w34589_
	);
	LUT2 #(
		.INIT('h4)
	) name24078 (
		\wishbone_RxReady_reg/NET0131 ,
		_w15138_,
		_w34590_
	);
	LUT2 #(
		.INIT('h2)
	) name24079 (
		\wishbone_Busy_IRQ_rck_reg/NET0131 ,
		\wishbone_Busy_IRQ_syncb2_reg/P0001 ,
		_w34591_
	);
	LUT2 #(
		.INIT('h1)
	) name24080 (
		_w34590_,
		_w34591_,
		_w34592_
	);
	LUT2 #(
		.INIT('h8)
	) name24081 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		_w34201_,
		_w34593_
	);
	LUT2 #(
		.INIT('h8)
	) name24082 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w34593_,
		_w34594_
	);
	LUT2 #(
		.INIT('h1)
	) name24083 (
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w34594_,
		_w34595_
	);
	LUT2 #(
		.INIT('h1)
	) name24084 (
		_w34204_,
		_w34208_,
		_w34596_
	);
	LUT2 #(
		.INIT('h4)
	) name24085 (
		_w34595_,
		_w34596_,
		_w34597_
	);
	LUT2 #(
		.INIT('h8)
	) name24086 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		_w34204_,
		_w34598_
	);
	LUT2 #(
		.INIT('h1)
	) name24087 (
		_w34597_,
		_w34598_,
		_w34599_
	);
	LUT2 #(
		.INIT('h8)
	) name24088 (
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w34210_,
		_w34600_
	);
	LUT2 #(
		.INIT('h1)
	) name24089 (
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w34210_,
		_w34601_
	);
	LUT2 #(
		.INIT('h1)
	) name24090 (
		_w34204_,
		_w34600_,
		_w34602_
	);
	LUT2 #(
		.INIT('h4)
	) name24091 (
		_w34601_,
		_w34602_,
		_w34603_
	);
	LUT2 #(
		.INIT('h8)
	) name24092 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		_w34204_,
		_w34604_
	);
	LUT2 #(
		.INIT('h1)
	) name24093 (
		_w34603_,
		_w34604_,
		_w34605_
	);
	LUT2 #(
		.INIT('h8)
	) name24094 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		_w34204_,
		_w34606_
	);
	LUT2 #(
		.INIT('h2)
	) name24095 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w34201_,
		_w34607_
	);
	LUT2 #(
		.INIT('h8)
	) name24096 (
		_w34207_,
		_w34330_,
		_w34608_
	);
	LUT2 #(
		.INIT('h1)
	) name24097 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w34600_,
		_w34609_
	);
	LUT2 #(
		.INIT('h1)
	) name24098 (
		\wishbone_RxStatus_reg[13]/NET0131 ,
		_w34608_,
		_w34610_
	);
	LUT2 #(
		.INIT('h4)
	) name24099 (
		_w34609_,
		_w34610_,
		_w34611_
	);
	LUT2 #(
		.INIT('h1)
	) name24100 (
		_w34607_,
		_w34611_,
		_w34612_
	);
	LUT2 #(
		.INIT('h1)
	) name24101 (
		_w34200_,
		_w34612_,
		_w34613_
	);
	LUT2 #(
		.INIT('h1)
	) name24102 (
		_w34606_,
		_w34613_,
		_w34614_
	);
	LUT2 #(
		.INIT('h2)
	) name24103 (
		\miim1_clkgen_Counter_reg[5]/NET0131 ,
		_w31193_,
		_w34615_
	);
	LUT2 #(
		.INIT('h1)
	) name24104 (
		_w31207_,
		_w34615_,
		_w34616_
	);
	LUT2 #(
		.INIT('h2)
	) name24105 (
		\ethreg1_MIIMODER_0_DataOut_reg[6]/NET0131 ,
		_w31206_,
		_w34617_
	);
	LUT2 #(
		.INIT('h2)
	) name24106 (
		_w31208_,
		_w34242_,
		_w34618_
	);
	LUT2 #(
		.INIT('h4)
	) name24107 (
		_w34617_,
		_w34618_,
		_w34619_
	);
	LUT2 #(
		.INIT('h1)
	) name24108 (
		_w34616_,
		_w34619_,
		_w34620_
	);
	LUT2 #(
		.INIT('h2)
	) name24109 (
		_w12657_,
		_w33028_,
		_w34621_
	);
	LUT2 #(
		.INIT('h2)
	) name24110 (
		_w34445_,
		_w34621_,
		_w34622_
	);
	LUT2 #(
		.INIT('h8)
	) name24111 (
		_w34449_,
		_w34622_,
		_w34623_
	);
	LUT2 #(
		.INIT('h2)
	) name24112 (
		\wishbone_tx_fifo_fifo_reg[10][14]/P0001 ,
		_w34623_,
		_w34624_
	);
	LUT2 #(
		.INIT('h8)
	) name24113 (
		\m_wb_dat_i[14]_pad ,
		_w34623_,
		_w34625_
	);
	LUT2 #(
		.INIT('h1)
	) name24114 (
		_w34624_,
		_w34625_,
		_w34626_
	);
	LUT2 #(
		.INIT('h2)
	) name24115 (
		\wishbone_tx_fifo_fifo_reg[10][18]/P0001 ,
		_w34623_,
		_w34627_
	);
	LUT2 #(
		.INIT('h8)
	) name24116 (
		\m_wb_dat_i[18]_pad ,
		_w34623_,
		_w34628_
	);
	LUT2 #(
		.INIT('h1)
	) name24117 (
		_w34627_,
		_w34628_,
		_w34629_
	);
	LUT2 #(
		.INIT('h2)
	) name24118 (
		\wishbone_tx_fifo_fifo_reg[10][27]/P0001 ,
		_w34623_,
		_w34630_
	);
	LUT2 #(
		.INIT('h8)
	) name24119 (
		\m_wb_dat_i[27]_pad ,
		_w34623_,
		_w34631_
	);
	LUT2 #(
		.INIT('h1)
	) name24120 (
		_w34630_,
		_w34631_,
		_w34632_
	);
	LUT2 #(
		.INIT('h2)
	) name24121 (
		\wishbone_tx_fifo_fifo_reg[10][29]/P0001 ,
		_w34623_,
		_w34633_
	);
	LUT2 #(
		.INIT('h8)
	) name24122 (
		\m_wb_dat_i[29]_pad ,
		_w34623_,
		_w34634_
	);
	LUT2 #(
		.INIT('h1)
	) name24123 (
		_w34633_,
		_w34634_,
		_w34635_
	);
	LUT2 #(
		.INIT('h2)
	) name24124 (
		\wishbone_tx_fifo_fifo_reg[10][3]/P0001 ,
		_w34623_,
		_w34636_
	);
	LUT2 #(
		.INIT('h8)
	) name24125 (
		\m_wb_dat_i[3]_pad ,
		_w34623_,
		_w34637_
	);
	LUT2 #(
		.INIT('h1)
	) name24126 (
		_w34636_,
		_w34637_,
		_w34638_
	);
	LUT2 #(
		.INIT('h8)
	) name24127 (
		_w34453_,
		_w34622_,
		_w34639_
	);
	LUT2 #(
		.INIT('h2)
	) name24128 (
		\wishbone_tx_fifo_fifo_reg[12][12]/P0001 ,
		_w34639_,
		_w34640_
	);
	LUT2 #(
		.INIT('h8)
	) name24129 (
		\m_wb_dat_i[12]_pad ,
		_w34639_,
		_w34641_
	);
	LUT2 #(
		.INIT('h1)
	) name24130 (
		_w34640_,
		_w34641_,
		_w34642_
	);
	LUT2 #(
		.INIT('h2)
	) name24131 (
		\wishbone_tx_fifo_fifo_reg[12][14]/P0001 ,
		_w34639_,
		_w34643_
	);
	LUT2 #(
		.INIT('h8)
	) name24132 (
		\m_wb_dat_i[14]_pad ,
		_w34639_,
		_w34644_
	);
	LUT2 #(
		.INIT('h1)
	) name24133 (
		_w34643_,
		_w34644_,
		_w34645_
	);
	LUT2 #(
		.INIT('h2)
	) name24134 (
		\wishbone_tx_fifo_fifo_reg[12][18]/P0001 ,
		_w34639_,
		_w34646_
	);
	LUT2 #(
		.INIT('h8)
	) name24135 (
		\m_wb_dat_i[18]_pad ,
		_w34639_,
		_w34647_
	);
	LUT2 #(
		.INIT('h1)
	) name24136 (
		_w34646_,
		_w34647_,
		_w34648_
	);
	LUT2 #(
		.INIT('h2)
	) name24137 (
		\wishbone_tx_fifo_fifo_reg[12][22]/P0001 ,
		_w34639_,
		_w34649_
	);
	LUT2 #(
		.INIT('h8)
	) name24138 (
		\m_wb_dat_i[22]_pad ,
		_w34639_,
		_w34650_
	);
	LUT2 #(
		.INIT('h1)
	) name24139 (
		_w34649_,
		_w34650_,
		_w34651_
	);
	LUT2 #(
		.INIT('h2)
	) name24140 (
		\wishbone_tx_fifo_fifo_reg[12][25]/P0001 ,
		_w34639_,
		_w34652_
	);
	LUT2 #(
		.INIT('h8)
	) name24141 (
		\m_wb_dat_i[25]_pad ,
		_w34639_,
		_w34653_
	);
	LUT2 #(
		.INIT('h1)
	) name24142 (
		_w34652_,
		_w34653_,
		_w34654_
	);
	LUT2 #(
		.INIT('h2)
	) name24143 (
		\wishbone_tx_fifo_fifo_reg[12][27]/P0001 ,
		_w34639_,
		_w34655_
	);
	LUT2 #(
		.INIT('h8)
	) name24144 (
		\m_wb_dat_i[27]_pad ,
		_w34639_,
		_w34656_
	);
	LUT2 #(
		.INIT('h1)
	) name24145 (
		_w34655_,
		_w34656_,
		_w34657_
	);
	LUT2 #(
		.INIT('h2)
	) name24146 (
		\wishbone_tx_fifo_fifo_reg[12][28]/P0001 ,
		_w34639_,
		_w34658_
	);
	LUT2 #(
		.INIT('h8)
	) name24147 (
		\m_wb_dat_i[28]_pad ,
		_w34639_,
		_w34659_
	);
	LUT2 #(
		.INIT('h1)
	) name24148 (
		_w34658_,
		_w34659_,
		_w34660_
	);
	LUT2 #(
		.INIT('h2)
	) name24149 (
		\wishbone_tx_fifo_fifo_reg[12][30]/P0001 ,
		_w34639_,
		_w34661_
	);
	LUT2 #(
		.INIT('h8)
	) name24150 (
		\m_wb_dat_i[30]_pad ,
		_w34639_,
		_w34662_
	);
	LUT2 #(
		.INIT('h1)
	) name24151 (
		_w34661_,
		_w34662_,
		_w34663_
	);
	LUT2 #(
		.INIT('h2)
	) name24152 (
		\wishbone_tx_fifo_fifo_reg[12][3]/P0001 ,
		_w34639_,
		_w34664_
	);
	LUT2 #(
		.INIT('h8)
	) name24153 (
		\m_wb_dat_i[3]_pad ,
		_w34639_,
		_w34665_
	);
	LUT2 #(
		.INIT('h1)
	) name24154 (
		_w34664_,
		_w34665_,
		_w34666_
	);
	LUT2 #(
		.INIT('h2)
	) name24155 (
		\wishbone_tx_fifo_fifo_reg[12][6]/P0001 ,
		_w34639_,
		_w34667_
	);
	LUT2 #(
		.INIT('h8)
	) name24156 (
		\m_wb_dat_i[6]_pad ,
		_w34639_,
		_w34668_
	);
	LUT2 #(
		.INIT('h1)
	) name24157 (
		_w34667_,
		_w34668_,
		_w34669_
	);
	LUT2 #(
		.INIT('h2)
	) name24158 (
		_w34465_,
		_w34621_,
		_w34670_
	);
	LUT2 #(
		.INIT('h8)
	) name24159 (
		_w34449_,
		_w34670_,
		_w34671_
	);
	LUT2 #(
		.INIT('h2)
	) name24160 (
		\wishbone_tx_fifo_fifo_reg[3][10]/P0001 ,
		_w34671_,
		_w34672_
	);
	LUT2 #(
		.INIT('h8)
	) name24161 (
		\m_wb_dat_i[10]_pad ,
		_w34671_,
		_w34673_
	);
	LUT2 #(
		.INIT('h1)
	) name24162 (
		_w34672_,
		_w34673_,
		_w34674_
	);
	LUT2 #(
		.INIT('h2)
	) name24163 (
		\wishbone_tx_fifo_fifo_reg[3][11]/P0001 ,
		_w34671_,
		_w34675_
	);
	LUT2 #(
		.INIT('h8)
	) name24164 (
		\m_wb_dat_i[11]_pad ,
		_w34671_,
		_w34676_
	);
	LUT2 #(
		.INIT('h1)
	) name24165 (
		_w34675_,
		_w34676_,
		_w34677_
	);
	LUT2 #(
		.INIT('h2)
	) name24166 (
		\wishbone_tx_fifo_fifo_reg[3][13]/P0001 ,
		_w34671_,
		_w34678_
	);
	LUT2 #(
		.INIT('h8)
	) name24167 (
		\m_wb_dat_i[13]_pad ,
		_w34671_,
		_w34679_
	);
	LUT2 #(
		.INIT('h1)
	) name24168 (
		_w34678_,
		_w34679_,
		_w34680_
	);
	LUT2 #(
		.INIT('h2)
	) name24169 (
		\wishbone_tx_fifo_fifo_reg[3][18]/P0001 ,
		_w34671_,
		_w34681_
	);
	LUT2 #(
		.INIT('h8)
	) name24170 (
		\m_wb_dat_i[18]_pad ,
		_w34671_,
		_w34682_
	);
	LUT2 #(
		.INIT('h1)
	) name24171 (
		_w34681_,
		_w34682_,
		_w34683_
	);
	LUT2 #(
		.INIT('h2)
	) name24172 (
		\wishbone_tx_fifo_fifo_reg[3][19]/P0001 ,
		_w34671_,
		_w34684_
	);
	LUT2 #(
		.INIT('h8)
	) name24173 (
		\m_wb_dat_i[19]_pad ,
		_w34671_,
		_w34685_
	);
	LUT2 #(
		.INIT('h1)
	) name24174 (
		_w34684_,
		_w34685_,
		_w34686_
	);
	LUT2 #(
		.INIT('h2)
	) name24175 (
		\wishbone_tx_fifo_fifo_reg[3][25]/P0001 ,
		_w34671_,
		_w34687_
	);
	LUT2 #(
		.INIT('h8)
	) name24176 (
		\m_wb_dat_i[25]_pad ,
		_w34671_,
		_w34688_
	);
	LUT2 #(
		.INIT('h1)
	) name24177 (
		_w34687_,
		_w34688_,
		_w34689_
	);
	LUT2 #(
		.INIT('h2)
	) name24178 (
		\wishbone_tx_fifo_fifo_reg[3][29]/P0001 ,
		_w34671_,
		_w34690_
	);
	LUT2 #(
		.INIT('h8)
	) name24179 (
		\m_wb_dat_i[29]_pad ,
		_w34671_,
		_w34691_
	);
	LUT2 #(
		.INIT('h1)
	) name24180 (
		_w34690_,
		_w34691_,
		_w34692_
	);
	LUT2 #(
		.INIT('h2)
	) name24181 (
		\wishbone_tx_fifo_fifo_reg[3][31]/P0001 ,
		_w34671_,
		_w34693_
	);
	LUT2 #(
		.INIT('h8)
	) name24182 (
		\m_wb_dat_i[31]_pad ,
		_w34671_,
		_w34694_
	);
	LUT2 #(
		.INIT('h1)
	) name24183 (
		_w34693_,
		_w34694_,
		_w34695_
	);
	LUT2 #(
		.INIT('h2)
	) name24184 (
		\wishbone_tx_fifo_fifo_reg[3][4]/P0001 ,
		_w34671_,
		_w34696_
	);
	LUT2 #(
		.INIT('h8)
	) name24185 (
		\m_wb_dat_i[4]_pad ,
		_w34671_,
		_w34697_
	);
	LUT2 #(
		.INIT('h1)
	) name24186 (
		_w34696_,
		_w34697_,
		_w34698_
	);
	LUT2 #(
		.INIT('h2)
	) name24187 (
		\wishbone_tx_fifo_fifo_reg[3][5]/P0001 ,
		_w34671_,
		_w34699_
	);
	LUT2 #(
		.INIT('h8)
	) name24188 (
		\m_wb_dat_i[5]_pad ,
		_w34671_,
		_w34700_
	);
	LUT2 #(
		.INIT('h1)
	) name24189 (
		_w34699_,
		_w34700_,
		_w34701_
	);
	LUT2 #(
		.INIT('h2)
	) name24190 (
		\wishbone_tx_fifo_fifo_reg[3][8]/P0001 ,
		_w34671_,
		_w34702_
	);
	LUT2 #(
		.INIT('h8)
	) name24191 (
		\m_wb_dat_i[8]_pad ,
		_w34671_,
		_w34703_
	);
	LUT2 #(
		.INIT('h1)
	) name24192 (
		_w34702_,
		_w34703_,
		_w34704_
	);
	LUT2 #(
		.INIT('h8)
	) name24193 (
		_w34453_,
		_w34670_,
		_w34705_
	);
	LUT2 #(
		.INIT('h2)
	) name24194 (
		\wishbone_tx_fifo_fifo_reg[5][11]/P0001 ,
		_w34705_,
		_w34706_
	);
	LUT2 #(
		.INIT('h8)
	) name24195 (
		\m_wb_dat_i[11]_pad ,
		_w34705_,
		_w34707_
	);
	LUT2 #(
		.INIT('h1)
	) name24196 (
		_w34706_,
		_w34707_,
		_w34708_
	);
	LUT2 #(
		.INIT('h2)
	) name24197 (
		\wishbone_tx_fifo_fifo_reg[5][18]/P0001 ,
		_w34705_,
		_w34709_
	);
	LUT2 #(
		.INIT('h8)
	) name24198 (
		\m_wb_dat_i[18]_pad ,
		_w34705_,
		_w34710_
	);
	LUT2 #(
		.INIT('h1)
	) name24199 (
		_w34709_,
		_w34710_,
		_w34711_
	);
	LUT2 #(
		.INIT('h2)
	) name24200 (
		\wishbone_tx_fifo_fifo_reg[5][19]/P0001 ,
		_w34705_,
		_w34712_
	);
	LUT2 #(
		.INIT('h8)
	) name24201 (
		\m_wb_dat_i[19]_pad ,
		_w34705_,
		_w34713_
	);
	LUT2 #(
		.INIT('h1)
	) name24202 (
		_w34712_,
		_w34713_,
		_w34714_
	);
	LUT2 #(
		.INIT('h2)
	) name24203 (
		\wishbone_tx_fifo_fifo_reg[5][1]/P0001 ,
		_w34705_,
		_w34715_
	);
	LUT2 #(
		.INIT('h8)
	) name24204 (
		\m_wb_dat_i[1]_pad ,
		_w34705_,
		_w34716_
	);
	LUT2 #(
		.INIT('h1)
	) name24205 (
		_w34715_,
		_w34716_,
		_w34717_
	);
	LUT2 #(
		.INIT('h2)
	) name24206 (
		\wishbone_tx_fifo_fifo_reg[5][23]/P0001 ,
		_w34705_,
		_w34718_
	);
	LUT2 #(
		.INIT('h8)
	) name24207 (
		\m_wb_dat_i[23]_pad ,
		_w34705_,
		_w34719_
	);
	LUT2 #(
		.INIT('h1)
	) name24208 (
		_w34718_,
		_w34719_,
		_w34720_
	);
	LUT2 #(
		.INIT('h2)
	) name24209 (
		\wishbone_tx_fifo_fifo_reg[5][24]/P0001 ,
		_w34705_,
		_w34721_
	);
	LUT2 #(
		.INIT('h8)
	) name24210 (
		\m_wb_dat_i[24]_pad ,
		_w34705_,
		_w34722_
	);
	LUT2 #(
		.INIT('h1)
	) name24211 (
		_w34721_,
		_w34722_,
		_w34723_
	);
	LUT2 #(
		.INIT('h2)
	) name24212 (
		\wishbone_tx_fifo_fifo_reg[5][25]/P0001 ,
		_w34705_,
		_w34724_
	);
	LUT2 #(
		.INIT('h8)
	) name24213 (
		\m_wb_dat_i[25]_pad ,
		_w34705_,
		_w34725_
	);
	LUT2 #(
		.INIT('h1)
	) name24214 (
		_w34724_,
		_w34725_,
		_w34726_
	);
	LUT2 #(
		.INIT('h2)
	) name24215 (
		\wishbone_tx_fifo_fifo_reg[5][26]/P0001 ,
		_w34705_,
		_w34727_
	);
	LUT2 #(
		.INIT('h8)
	) name24216 (
		\m_wb_dat_i[26]_pad ,
		_w34705_,
		_w34728_
	);
	LUT2 #(
		.INIT('h1)
	) name24217 (
		_w34727_,
		_w34728_,
		_w34729_
	);
	LUT2 #(
		.INIT('h2)
	) name24218 (
		\wishbone_tx_fifo_fifo_reg[5][28]/P0001 ,
		_w34705_,
		_w34730_
	);
	LUT2 #(
		.INIT('h8)
	) name24219 (
		\m_wb_dat_i[28]_pad ,
		_w34705_,
		_w34731_
	);
	LUT2 #(
		.INIT('h1)
	) name24220 (
		_w34730_,
		_w34731_,
		_w34732_
	);
	LUT2 #(
		.INIT('h2)
	) name24221 (
		\wishbone_tx_fifo_fifo_reg[5][3]/P0001 ,
		_w34705_,
		_w34733_
	);
	LUT2 #(
		.INIT('h8)
	) name24222 (
		\m_wb_dat_i[3]_pad ,
		_w34705_,
		_w34734_
	);
	LUT2 #(
		.INIT('h1)
	) name24223 (
		_w34733_,
		_w34734_,
		_w34735_
	);
	LUT2 #(
		.INIT('h2)
	) name24224 (
		\wishbone_tx_fifo_fifo_reg[5][8]/P0001 ,
		_w34705_,
		_w34736_
	);
	LUT2 #(
		.INIT('h8)
	) name24225 (
		\m_wb_dat_i[8]_pad ,
		_w34705_,
		_w34737_
	);
	LUT2 #(
		.INIT('h1)
	) name24226 (
		_w34736_,
		_w34737_,
		_w34738_
	);
	LUT2 #(
		.INIT('h2)
	) name24227 (
		_w34470_,
		_w34621_,
		_w34739_
	);
	LUT2 #(
		.INIT('h8)
	) name24228 (
		_w34469_,
		_w34739_,
		_w34740_
	);
	LUT2 #(
		.INIT('h2)
	) name24229 (
		\wishbone_tx_fifo_fifo_reg[6][11]/P0001 ,
		_w34740_,
		_w34741_
	);
	LUT2 #(
		.INIT('h8)
	) name24230 (
		\m_wb_dat_i[11]_pad ,
		_w34740_,
		_w34742_
	);
	LUT2 #(
		.INIT('h1)
	) name24231 (
		_w34741_,
		_w34742_,
		_w34743_
	);
	LUT2 #(
		.INIT('h2)
	) name24232 (
		\wishbone_tx_fifo_fifo_reg[6][12]/P0001 ,
		_w34740_,
		_w34744_
	);
	LUT2 #(
		.INIT('h8)
	) name24233 (
		\m_wb_dat_i[12]_pad ,
		_w34740_,
		_w34745_
	);
	LUT2 #(
		.INIT('h1)
	) name24234 (
		_w34744_,
		_w34745_,
		_w34746_
	);
	LUT2 #(
		.INIT('h2)
	) name24235 (
		\wishbone_tx_fifo_fifo_reg[6][14]/P0001 ,
		_w34740_,
		_w34747_
	);
	LUT2 #(
		.INIT('h8)
	) name24236 (
		\m_wb_dat_i[14]_pad ,
		_w34740_,
		_w34748_
	);
	LUT2 #(
		.INIT('h1)
	) name24237 (
		_w34747_,
		_w34748_,
		_w34749_
	);
	LUT2 #(
		.INIT('h2)
	) name24238 (
		\wishbone_tx_fifo_fifo_reg[6][16]/P0001 ,
		_w34740_,
		_w34750_
	);
	LUT2 #(
		.INIT('h8)
	) name24239 (
		\m_wb_dat_i[16]_pad ,
		_w34740_,
		_w34751_
	);
	LUT2 #(
		.INIT('h1)
	) name24240 (
		_w34750_,
		_w34751_,
		_w34752_
	);
	LUT2 #(
		.INIT('h2)
	) name24241 (
		\wishbone_tx_fifo_fifo_reg[6][18]/P0001 ,
		_w34740_,
		_w34753_
	);
	LUT2 #(
		.INIT('h8)
	) name24242 (
		\m_wb_dat_i[18]_pad ,
		_w34740_,
		_w34754_
	);
	LUT2 #(
		.INIT('h1)
	) name24243 (
		_w34753_,
		_w34754_,
		_w34755_
	);
	LUT2 #(
		.INIT('h2)
	) name24244 (
		\wishbone_tx_fifo_fifo_reg[6][1]/P0001 ,
		_w34740_,
		_w34756_
	);
	LUT2 #(
		.INIT('h8)
	) name24245 (
		\m_wb_dat_i[1]_pad ,
		_w34740_,
		_w34757_
	);
	LUT2 #(
		.INIT('h1)
	) name24246 (
		_w34756_,
		_w34757_,
		_w34758_
	);
	LUT2 #(
		.INIT('h2)
	) name24247 (
		\wishbone_tx_fifo_fifo_reg[6][20]/P0001 ,
		_w34740_,
		_w34759_
	);
	LUT2 #(
		.INIT('h8)
	) name24248 (
		\m_wb_dat_i[20]_pad ,
		_w34740_,
		_w34760_
	);
	LUT2 #(
		.INIT('h1)
	) name24249 (
		_w34759_,
		_w34760_,
		_w34761_
	);
	LUT2 #(
		.INIT('h2)
	) name24250 (
		\wishbone_tx_fifo_fifo_reg[6][25]/P0001 ,
		_w34740_,
		_w34762_
	);
	LUT2 #(
		.INIT('h8)
	) name24251 (
		\m_wb_dat_i[25]_pad ,
		_w34740_,
		_w34763_
	);
	LUT2 #(
		.INIT('h1)
	) name24252 (
		_w34762_,
		_w34763_,
		_w34764_
	);
	LUT2 #(
		.INIT('h2)
	) name24253 (
		\wishbone_tx_fifo_fifo_reg[6][27]/P0001 ,
		_w34740_,
		_w34765_
	);
	LUT2 #(
		.INIT('h8)
	) name24254 (
		\m_wb_dat_i[27]_pad ,
		_w34740_,
		_w34766_
	);
	LUT2 #(
		.INIT('h1)
	) name24255 (
		_w34765_,
		_w34766_,
		_w34767_
	);
	LUT2 #(
		.INIT('h2)
	) name24256 (
		\wishbone_tx_fifo_fifo_reg[6][28]/P0001 ,
		_w34740_,
		_w34768_
	);
	LUT2 #(
		.INIT('h8)
	) name24257 (
		\m_wb_dat_i[28]_pad ,
		_w34740_,
		_w34769_
	);
	LUT2 #(
		.INIT('h1)
	) name24258 (
		_w34768_,
		_w34769_,
		_w34770_
	);
	LUT2 #(
		.INIT('h2)
	) name24259 (
		\wishbone_tx_fifo_fifo_reg[6][30]/P0001 ,
		_w34740_,
		_w34771_
	);
	LUT2 #(
		.INIT('h8)
	) name24260 (
		\m_wb_dat_i[30]_pad ,
		_w34740_,
		_w34772_
	);
	LUT2 #(
		.INIT('h1)
	) name24261 (
		_w34771_,
		_w34772_,
		_w34773_
	);
	LUT2 #(
		.INIT('h2)
	) name24262 (
		\wishbone_tx_fifo_fifo_reg[6][3]/P0001 ,
		_w34740_,
		_w34774_
	);
	LUT2 #(
		.INIT('h8)
	) name24263 (
		\m_wb_dat_i[3]_pad ,
		_w34740_,
		_w34775_
	);
	LUT2 #(
		.INIT('h1)
	) name24264 (
		_w34774_,
		_w34775_,
		_w34776_
	);
	LUT2 #(
		.INIT('h2)
	) name24265 (
		\wishbone_tx_fifo_fifo_reg[6][4]/P0001 ,
		_w34740_,
		_w34777_
	);
	LUT2 #(
		.INIT('h8)
	) name24266 (
		\m_wb_dat_i[4]_pad ,
		_w34740_,
		_w34778_
	);
	LUT2 #(
		.INIT('h1)
	) name24267 (
		_w34777_,
		_w34778_,
		_w34779_
	);
	LUT2 #(
		.INIT('h2)
	) name24268 (
		\wishbone_tx_fifo_fifo_reg[6][5]/P0001 ,
		_w34740_,
		_w34780_
	);
	LUT2 #(
		.INIT('h8)
	) name24269 (
		\m_wb_dat_i[5]_pad ,
		_w34740_,
		_w34781_
	);
	LUT2 #(
		.INIT('h1)
	) name24270 (
		_w34780_,
		_w34781_,
		_w34782_
	);
	LUT2 #(
		.INIT('h2)
	) name24271 (
		\wishbone_tx_fifo_fifo_reg[6][6]/P0001 ,
		_w34740_,
		_w34783_
	);
	LUT2 #(
		.INIT('h8)
	) name24272 (
		\m_wb_dat_i[6]_pad ,
		_w34740_,
		_w34784_
	);
	LUT2 #(
		.INIT('h1)
	) name24273 (
		_w34783_,
		_w34784_,
		_w34785_
	);
	LUT2 #(
		.INIT('h2)
	) name24274 (
		\wishbone_tx_fifo_fifo_reg[6][7]/P0001 ,
		_w34740_,
		_w34786_
	);
	LUT2 #(
		.INIT('h8)
	) name24275 (
		\m_wb_dat_i[7]_pad ,
		_w34740_,
		_w34787_
	);
	LUT2 #(
		.INIT('h1)
	) name24276 (
		_w34786_,
		_w34787_,
		_w34788_
	);
	LUT2 #(
		.INIT('h2)
	) name24277 (
		\wishbone_tx_fifo_fifo_reg[6][8]/P0001 ,
		_w34740_,
		_w34789_
	);
	LUT2 #(
		.INIT('h8)
	) name24278 (
		\m_wb_dat_i[8]_pad ,
		_w34740_,
		_w34790_
	);
	LUT2 #(
		.INIT('h1)
	) name24279 (
		_w34789_,
		_w34790_,
		_w34791_
	);
	LUT2 #(
		.INIT('h2)
	) name24280 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34621_,
		_w34792_
	);
	LUT2 #(
		.INIT('h8)
	) name24281 (
		_w34460_,
		_w34792_,
		_w34793_
	);
	LUT2 #(
		.INIT('h2)
	) name24282 (
		\wishbone_tx_fifo_fifo_reg[9][12]/P0001 ,
		_w34793_,
		_w34794_
	);
	LUT2 #(
		.INIT('h8)
	) name24283 (
		\m_wb_dat_i[12]_pad ,
		_w34793_,
		_w34795_
	);
	LUT2 #(
		.INIT('h1)
	) name24284 (
		_w34794_,
		_w34795_,
		_w34796_
	);
	LUT2 #(
		.INIT('h2)
	) name24285 (
		\wishbone_tx_fifo_fifo_reg[9][13]/P0001 ,
		_w34793_,
		_w34797_
	);
	LUT2 #(
		.INIT('h8)
	) name24286 (
		\m_wb_dat_i[13]_pad ,
		_w34793_,
		_w34798_
	);
	LUT2 #(
		.INIT('h1)
	) name24287 (
		_w34797_,
		_w34798_,
		_w34799_
	);
	LUT2 #(
		.INIT('h2)
	) name24288 (
		\wishbone_tx_fifo_fifo_reg[9][14]/P0001 ,
		_w34793_,
		_w34800_
	);
	LUT2 #(
		.INIT('h8)
	) name24289 (
		\m_wb_dat_i[14]_pad ,
		_w34793_,
		_w34801_
	);
	LUT2 #(
		.INIT('h1)
	) name24290 (
		_w34800_,
		_w34801_,
		_w34802_
	);
	LUT2 #(
		.INIT('h2)
	) name24291 (
		\wishbone_tx_fifo_fifo_reg[9][20]/P0001 ,
		_w34793_,
		_w34803_
	);
	LUT2 #(
		.INIT('h8)
	) name24292 (
		\m_wb_dat_i[20]_pad ,
		_w34793_,
		_w34804_
	);
	LUT2 #(
		.INIT('h1)
	) name24293 (
		_w34803_,
		_w34804_,
		_w34805_
	);
	LUT2 #(
		.INIT('h2)
	) name24294 (
		\wishbone_tx_fifo_fifo_reg[9][25]/P0001 ,
		_w34793_,
		_w34806_
	);
	LUT2 #(
		.INIT('h8)
	) name24295 (
		\m_wb_dat_i[25]_pad ,
		_w34793_,
		_w34807_
	);
	LUT2 #(
		.INIT('h1)
	) name24296 (
		_w34806_,
		_w34807_,
		_w34808_
	);
	LUT2 #(
		.INIT('h2)
	) name24297 (
		\wishbone_tx_fifo_fifo_reg[9][26]/P0001 ,
		_w34793_,
		_w34809_
	);
	LUT2 #(
		.INIT('h8)
	) name24298 (
		\m_wb_dat_i[26]_pad ,
		_w34793_,
		_w34810_
	);
	LUT2 #(
		.INIT('h1)
	) name24299 (
		_w34809_,
		_w34810_,
		_w34811_
	);
	LUT2 #(
		.INIT('h2)
	) name24300 (
		\wishbone_tx_fifo_fifo_reg[9][30]/P0001 ,
		_w34793_,
		_w34812_
	);
	LUT2 #(
		.INIT('h8)
	) name24301 (
		\m_wb_dat_i[30]_pad ,
		_w34793_,
		_w34813_
	);
	LUT2 #(
		.INIT('h1)
	) name24302 (
		_w34812_,
		_w34813_,
		_w34814_
	);
	LUT2 #(
		.INIT('h2)
	) name24303 (
		\wishbone_tx_fifo_fifo_reg[9][5]/P0001 ,
		_w34793_,
		_w34815_
	);
	LUT2 #(
		.INIT('h8)
	) name24304 (
		\m_wb_dat_i[5]_pad ,
		_w34793_,
		_w34816_
	);
	LUT2 #(
		.INIT('h1)
	) name24305 (
		_w34815_,
		_w34816_,
		_w34817_
	);
	LUT2 #(
		.INIT('h2)
	) name24306 (
		\wishbone_tx_fifo_fifo_reg[9][8]/P0001 ,
		_w34793_,
		_w34818_
	);
	LUT2 #(
		.INIT('h8)
	) name24307 (
		\m_wb_dat_i[8]_pad ,
		_w34793_,
		_w34819_
	);
	LUT2 #(
		.INIT('h1)
	) name24308 (
		_w34818_,
		_w34819_,
		_w34820_
	);
	LUT2 #(
		.INIT('h2)
	) name24309 (
		\wishbone_tx_fifo_fifo_reg[6][23]/P0001 ,
		_w34740_,
		_w34821_
	);
	LUT2 #(
		.INIT('h8)
	) name24310 (
		\m_wb_dat_i[23]_pad ,
		_w34740_,
		_w34822_
	);
	LUT2 #(
		.INIT('h1)
	) name24311 (
		_w34821_,
		_w34822_,
		_w34823_
	);
	LUT2 #(
		.INIT('h8)
	) name24312 (
		_w34459_,
		_w34469_,
		_w34824_
	);
	LUT2 #(
		.INIT('h1)
	) name24313 (
		_w34621_,
		_w34824_,
		_w34825_
	);
	LUT2 #(
		.INIT('h8)
	) name24314 (
		_w34450_,
		_w34456_,
		_w34826_
	);
	LUT2 #(
		.INIT('h8)
	) name24315 (
		_w34445_,
		_w34447_,
		_w34827_
	);
	LUT2 #(
		.INIT('h8)
	) name24316 (
		_w34471_,
		_w34827_,
		_w34828_
	);
	LUT2 #(
		.INIT('h8)
	) name24317 (
		_w34471_,
		_w34478_,
		_w34829_
	);
	LUT2 #(
		.INIT('h8)
	) name24318 (
		_w34477_,
		_w34827_,
		_w34830_
	);
	LUT2 #(
		.INIT('h2)
	) name24319 (
		\wishbone_Busy_IRQ_sync2_reg/P0001 ,
		\wishbone_Busy_IRQ_sync3_reg/P0001 ,
		_w34831_
	);
	LUT2 #(
		.INIT('h8)
	) name24320 (
		\wb_dat_i[4]_pad ,
		_w34567_,
		_w34832_
	);
	LUT2 #(
		.INIT('h2)
	) name24321 (
		\ethreg1_irq_busy_reg/NET0131 ,
		_w34832_,
		_w34833_
	);
	LUT2 #(
		.INIT('h1)
	) name24322 (
		_w34831_,
		_w34833_,
		_w34834_
	);
	LUT2 #(
		.INIT('h4)
	) name24323 (
		\miim1_LatchByte_reg[0]/NET0131 ,
		\miim1_LatchByte_reg[1]/NET0131 ,
		_w34835_
	);
	LUT2 #(
		.INIT('h8)
	) name24324 (
		_w31426_,
		_w34835_,
		_w34836_
	);
	LUT2 #(
		.INIT('h8)
	) name24325 (
		_w31401_,
		_w34836_,
		_w34837_
	);
	LUT2 #(
		.INIT('h2)
	) name24326 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		_w31950_,
		_w34838_
	);
	LUT2 #(
		.INIT('h2)
	) name24327 (
		_w34139_,
		_w34838_,
		_w34839_
	);
	LUT2 #(
		.INIT('h4)
	) name24328 (
		_w34139_,
		_w34838_,
		_w34840_
	);
	LUT2 #(
		.INIT('h1)
	) name24329 (
		_w34839_,
		_w34840_,
		_w34841_
	);
	LUT2 #(
		.INIT('h2)
	) name24330 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11472_,
		_w34842_
	);
	LUT2 #(
		.INIT('h1)
	) name24331 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[13]/NET0131 ,
		_w34843_
	);
	LUT2 #(
		.INIT('h1)
	) name24332 (
		_w34842_,
		_w34843_,
		_w34844_
	);
	LUT2 #(
		.INIT('h2)
	) name24333 (
		_w10580_,
		_w11767_,
		_w34845_
	);
	LUT2 #(
		.INIT('h2)
	) name24334 (
		_w10580_,
		_w11427_,
		_w34846_
	);
	LUT2 #(
		.INIT('h2)
	) name24335 (
		_w10580_,
		_w11236_,
		_w34847_
	);
	LUT2 #(
		.INIT('h1)
	) name24336 (
		_w34137_,
		_w34140_,
		_w34848_
	);
	LUT2 #(
		.INIT('h1)
	) name24337 (
		_w12551_,
		_w34138_,
		_w34849_
	);
	LUT2 #(
		.INIT('h1)
	) name24338 (
		_w34848_,
		_w34849_,
		_w34850_
	);
	LUT2 #(
		.INIT('h1)
	) name24339 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w34850_,
		_w34851_
	);
	LUT2 #(
		.INIT('h8)
	) name24340 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w34850_,
		_w34852_
	);
	LUT2 #(
		.INIT('h1)
	) name24341 (
		_w31950_,
		_w34851_,
		_w34853_
	);
	LUT2 #(
		.INIT('h4)
	) name24342 (
		_w34852_,
		_w34853_,
		_w34854_
	);
	LUT2 #(
		.INIT('h1)
	) name24343 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		\wishbone_LatchedRxStartFrm_reg/NET0131 ,
		_w34855_
	);
	LUT2 #(
		.INIT('h1)
	) name24344 (
		\wishbone_SyncRxStartFrm_q_reg/NET0131 ,
		_w34855_,
		_w34856_
	);
	LUT2 #(
		.INIT('h8)
	) name24345 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w34857_
	);
	LUT2 #(
		.INIT('h2)
	) name24346 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34858_
	);
	LUT2 #(
		.INIT('h4)
	) name24347 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w34859_
	);
	LUT2 #(
		.INIT('h8)
	) name24348 (
		_w34858_,
		_w34859_,
		_w34860_
	);
	LUT2 #(
		.INIT('h1)
	) name24349 (
		_w34857_,
		_w34860_,
		_w34861_
	);
	LUT2 #(
		.INIT('h8)
	) name24350 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w34862_
	);
	LUT2 #(
		.INIT('h8)
	) name24351 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34862_,
		_w34863_
	);
	LUT2 #(
		.INIT('h8)
	) name24352 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w34863_,
		_w34864_
	);
	LUT2 #(
		.INIT('h1)
	) name24353 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w34864_,
		_w34865_
	);
	LUT2 #(
		.INIT('h8)
	) name24354 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[3]/NET0131 ,
		_w34864_,
		_w34866_
	);
	LUT2 #(
		.INIT('h2)
	) name24355 (
		_w34861_,
		_w34865_,
		_w34867_
	);
	LUT2 #(
		.INIT('h4)
	) name24356 (
		_w34866_,
		_w34867_,
		_w34868_
	);
	LUT2 #(
		.INIT('h8)
	) name24357 (
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w34139_,
		_w34869_
	);
	LUT2 #(
		.INIT('h1)
	) name24358 (
		_w12551_,
		_w34140_,
		_w34870_
	);
	LUT2 #(
		.INIT('h2)
	) name24359 (
		_w34137_,
		_w34870_,
		_w34871_
	);
	LUT2 #(
		.INIT('h8)
	) name24360 (
		_w34138_,
		_w34870_,
		_w34872_
	);
	LUT2 #(
		.INIT('h1)
	) name24361 (
		_w34871_,
		_w34872_,
		_w34873_
	);
	LUT2 #(
		.INIT('h4)
	) name24362 (
		_w34869_,
		_w34873_,
		_w34874_
	);
	LUT2 #(
		.INIT('h1)
	) name24363 (
		_w31950_,
		_w34874_,
		_w34875_
	);
	LUT2 #(
		.INIT('h1)
	) name24364 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[3]/NET0131 ,
		_w11622_,
		_w34876_
	);
	LUT2 #(
		.INIT('h1)
	) name24365 (
		wb_rst_i_pad,
		_w11623_,
		_w34877_
	);
	LUT2 #(
		.INIT('h4)
	) name24366 (
		_w34876_,
		_w34877_,
		_w34878_
	);
	LUT2 #(
		.INIT('h8)
	) name24367 (
		\wishbone_StartOccured_reg/NET0131 ,
		_w34290_,
		_w34879_
	);
	LUT2 #(
		.INIT('h1)
	) name24368 (
		\wishbone_TxStartFrm_wb_reg/NET0131 ,
		_w34879_,
		_w34880_
	);
	LUT2 #(
		.INIT('h1)
	) name24369 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		_w34881_
	);
	LUT2 #(
		.INIT('h1)
	) name24370 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[3]/NET0131 ,
		_w34882_
	);
	LUT2 #(
		.INIT('h1)
	) name24371 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[5]/NET0131 ,
		_w34883_
	);
	LUT2 #(
		.INIT('h1)
	) name24372 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_TX_BD_NUM_0_DataOut_reg[7]/NET0131 ,
		_w34884_
	);
	LUT2 #(
		.INIT('h8)
	) name24373 (
		_w34883_,
		_w34884_,
		_w34885_
	);
	LUT2 #(
		.INIT('h8)
	) name24374 (
		_w34881_,
		_w34882_,
		_w34886_
	);
	LUT2 #(
		.INIT('h8)
	) name24375 (
		_w34885_,
		_w34886_,
		_w34887_
	);
	LUT2 #(
		.INIT('h2)
	) name24376 (
		\ethreg1_MODER_0_DataOut_reg[1]/NET0131 ,
		_w34887_,
		_w34888_
	);
	LUT2 #(
		.INIT('h4)
	) name24377 (
		\wishbone_r_TxEn_q_reg/NET0131 ,
		_w34888_,
		_w34889_
	);
	LUT2 #(
		.INIT('h1)
	) name24378 (
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		_w34890_
	);
	LUT2 #(
		.INIT('h2)
	) name24379 (
		_w12655_,
		_w34890_,
		_w34891_
	);
	LUT2 #(
		.INIT('h4)
	) name24380 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w34891_,
		_w34892_
	);
	LUT2 #(
		.INIT('h1)
	) name24381 (
		_w34889_,
		_w34892_,
		_w34893_
	);
	LUT2 #(
		.INIT('h8)
	) name24382 (
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w34893_,
		_w34894_
	);
	LUT2 #(
		.INIT('h4)
	) name24383 (
		\wishbone_TxStatus_reg[13]/NET0131 ,
		_w34892_,
		_w34895_
	);
	LUT2 #(
		.INIT('h4)
	) name24384 (
		_w34889_,
		_w34895_,
		_w34896_
	);
	LUT2 #(
		.INIT('h8)
	) name24385 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w34897_
	);
	LUT2 #(
		.INIT('h8)
	) name24386 (
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w34897_,
		_w34898_
	);
	LUT2 #(
		.INIT('h1)
	) name24387 (
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w34898_,
		_w34899_
	);
	LUT2 #(
		.INIT('h8)
	) name24388 (
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w34898_,
		_w34900_
	);
	LUT2 #(
		.INIT('h1)
	) name24389 (
		_w34899_,
		_w34900_,
		_w34901_
	);
	LUT2 #(
		.INIT('h8)
	) name24390 (
		_w34896_,
		_w34901_,
		_w34902_
	);
	LUT2 #(
		.INIT('h1)
	) name24391 (
		_w34894_,
		_w34902_,
		_w34903_
	);
	LUT2 #(
		.INIT('h8)
	) name24392 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w34900_,
		_w34904_
	);
	LUT2 #(
		.INIT('h8)
	) name24393 (
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		_w34904_,
		_w34905_
	);
	LUT2 #(
		.INIT('h2)
	) name24394 (
		_w34896_,
		_w34905_,
		_w34906_
	);
	LUT2 #(
		.INIT('h1)
	) name24395 (
		_w34893_,
		_w34906_,
		_w34907_
	);
	LUT2 #(
		.INIT('h2)
	) name24396 (
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		_w34907_,
		_w34908_
	);
	LUT2 #(
		.INIT('h8)
	) name24397 (
		_w34904_,
		_w34906_,
		_w34909_
	);
	LUT2 #(
		.INIT('h1)
	) name24398 (
		_w34908_,
		_w34909_,
		_w34910_
	);
	LUT2 #(
		.INIT('h2)
	) name24399 (
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		_w34907_,
		_w34911_
	);
	LUT2 #(
		.INIT('h4)
	) name24400 (
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		_w34905_,
		_w34912_
	);
	LUT2 #(
		.INIT('h8)
	) name24401 (
		_w34896_,
		_w34912_,
		_w34913_
	);
	LUT2 #(
		.INIT('h1)
	) name24402 (
		_w34911_,
		_w34913_,
		_w34914_
	);
	LUT2 #(
		.INIT('h8)
	) name24403 (
		\wishbone_TxEndFrm_wb_reg/NET0131 ,
		_w34290_,
		_w34915_
	);
	LUT2 #(
		.INIT('h8)
	) name24404 (
		_w13499_,
		_w16763_,
		_w34916_
	);
	LUT2 #(
		.INIT('h2)
	) name24405 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w34917_
	);
	LUT2 #(
		.INIT('h4)
	) name24406 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w34917_,
		_w34918_
	);
	LUT2 #(
		.INIT('h8)
	) name24407 (
		_w12240_,
		_w34088_,
		_w34919_
	);
	LUT2 #(
		.INIT('h8)
	) name24408 (
		_w34918_,
		_w34919_,
		_w34920_
	);
	LUT2 #(
		.INIT('h8)
	) name24409 (
		_w34916_,
		_w34920_,
		_w34921_
	);
	LUT2 #(
		.INIT('h1)
	) name24410 (
		_w34915_,
		_w34921_,
		_w34922_
	);
	LUT2 #(
		.INIT('h2)
	) name24411 (
		\miim1_outctrl_Mdo_2d_reg/NET0131 ,
		_w31401_,
		_w34923_
	);
	LUT2 #(
		.INIT('h8)
	) name24412 (
		\miim1_BitCounter_reg[3]/NET0131 ,
		_w34320_,
		_w34924_
	);
	LUT2 #(
		.INIT('h1)
	) name24413 (
		\miim1_BitCounter_reg[4]/NET0131 ,
		\miim1_BitCounter_reg[6]/NET0131 ,
		_w34925_
	);
	LUT2 #(
		.INIT('h4)
	) name24414 (
		_w34924_,
		_w34925_,
		_w34926_
	);
	LUT2 #(
		.INIT('h1)
	) name24415 (
		\miim1_WriteOp_reg/NET0131 ,
		_w34926_,
		_w34927_
	);
	LUT2 #(
		.INIT('h1)
	) name24416 (
		_w31404_,
		_w34927_,
		_w34928_
	);
	LUT2 #(
		.INIT('h1)
	) name24417 (
		_w31409_,
		_w34928_,
		_w34929_
	);
	LUT2 #(
		.INIT('h2)
	) name24418 (
		\miim1_InProgress_reg/NET0131 ,
		_w34929_,
		_w34930_
	);
	LUT2 #(
		.INIT('h8)
	) name24419 (
		_w31401_,
		_w31404_,
		_w34931_
	);
	LUT2 #(
		.INIT('h4)
	) name24420 (
		_w34930_,
		_w34931_,
		_w34932_
	);
	LUT2 #(
		.INIT('h1)
	) name24421 (
		_w34923_,
		_w34932_,
		_w34933_
	);
	LUT2 #(
		.INIT('h2)
	) name24422 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w34934_
	);
	LUT2 #(
		.INIT('h4)
	) name24423 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34934_,
		_w34935_
	);
	LUT2 #(
		.INIT('h1)
	) name24424 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[1]/NET0131 ,
		_w34936_
	);
	LUT2 #(
		.INIT('h8)
	) name24425 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34936_,
		_w34937_
	);
	LUT2 #(
		.INIT('h8)
	) name24426 (
		_w34935_,
		_w34937_,
		_w34938_
	);
	LUT2 #(
		.INIT('h8)
	) name24427 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[0]/NET0131 ,
		_w34938_,
		_w34939_
	);
	LUT2 #(
		.INIT('h4)
	) name24428 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[3]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[4]/NET0131 ,
		_w34940_
	);
	LUT2 #(
		.INIT('h4)
	) name24429 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34940_,
		_w34941_
	);
	LUT2 #(
		.INIT('h8)
	) name24430 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[0]/NET0131 ,
		_w34941_,
		_w34942_
	);
	LUT2 #(
		.INIT('h8)
	) name24431 (
		\ethreg1_TXCTRL_0_DataOut_reg[0]/NET0131 ,
		_w34263_,
		_w34943_
	);
	LUT2 #(
		.INIT('h1)
	) name24432 (
		_w34935_,
		_w34942_,
		_w34944_
	);
	LUT2 #(
		.INIT('h4)
	) name24433 (
		_w34943_,
		_w34944_,
		_w34945_
	);
	LUT2 #(
		.INIT('h2)
	) name24434 (
		_w34265_,
		_w34945_,
		_w34946_
	);
	LUT2 #(
		.INIT('h4)
	) name24435 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34936_,
		_w34947_
	);
	LUT2 #(
		.INIT('h8)
	) name24436 (
		\ethreg1_TXCTRL_1_DataOut_reg[0]/NET0131 ,
		_w34263_,
		_w34948_
	);
	LUT2 #(
		.INIT('h4)
	) name24437 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34262_,
		_w34949_
	);
	LUT2 #(
		.INIT('h4)
	) name24438 (
		_w34269_,
		_w34949_,
		_w34950_
	);
	LUT2 #(
		.INIT('h8)
	) name24439 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[0]/NET0131 ,
		_w34941_,
		_w34951_
	);
	LUT2 #(
		.INIT('h1)
	) name24440 (
		_w34948_,
		_w34950_,
		_w34952_
	);
	LUT2 #(
		.INIT('h4)
	) name24441 (
		_w34951_,
		_w34952_,
		_w34953_
	);
	LUT2 #(
		.INIT('h2)
	) name24442 (
		_w34947_,
		_w34953_,
		_w34954_
	);
	LUT2 #(
		.INIT('h8)
	) name24443 (
		_w34937_,
		_w34941_,
		_w34955_
	);
	LUT2 #(
		.INIT('h8)
	) name24444 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[0]/NET0131 ,
		_w34955_,
		_w34956_
	);
	LUT2 #(
		.INIT('h8)
	) name24445 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w34264_,
		_w34957_
	);
	LUT2 #(
		.INIT('h8)
	) name24446 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[0]/NET0131 ,
		_w34941_,
		_w34958_
	);
	LUT2 #(
		.INIT('h8)
	) name24447 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[0]/NET0131 ,
		_w34935_,
		_w34959_
	);
	LUT2 #(
		.INIT('h4)
	) name24448 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[5]/NET0131 ,
		_w34499_,
		_w34960_
	);
	LUT2 #(
		.INIT('h1)
	) name24449 (
		_w34958_,
		_w34960_,
		_w34961_
	);
	LUT2 #(
		.INIT('h4)
	) name24450 (
		_w34959_,
		_w34961_,
		_w34962_
	);
	LUT2 #(
		.INIT('h2)
	) name24451 (
		_w34957_,
		_w34962_,
		_w34963_
	);
	LUT2 #(
		.INIT('h1)
	) name24452 (
		_w34939_,
		_w34956_,
		_w34964_
	);
	LUT2 #(
		.INIT('h4)
	) name24453 (
		_w34946_,
		_w34964_,
		_w34965_
	);
	LUT2 #(
		.INIT('h1)
	) name24454 (
		_w34954_,
		_w34963_,
		_w34966_
	);
	LUT2 #(
		.INIT('h8)
	) name24455 (
		_w34965_,
		_w34966_,
		_w34967_
	);
	LUT2 #(
		.INIT('h8)
	) name24456 (
		\txethmac1_txstatem1_StateJam_q_reg/NET0131 ,
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		_w34968_
	);
	LUT2 #(
		.INIT('h2)
	) name24457 (
		\txethmac1_random1_RandomLatched_reg[9]/NET0131 ,
		_w34968_,
		_w34969_
	);
	LUT2 #(
		.INIT('h1)
	) name24458 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w34970_
	);
	LUT2 #(
		.INIT('h8)
	) name24459 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[9]/NET0131 ,
		_w34971_
	);
	LUT2 #(
		.INIT('h8)
	) name24460 (
		_w34968_,
		_w34971_,
		_w34972_
	);
	LUT2 #(
		.INIT('h4)
	) name24461 (
		_w34970_,
		_w34972_,
		_w34973_
	);
	LUT2 #(
		.INIT('h1)
	) name24462 (
		_w34969_,
		_w34973_,
		_w34974_
	);
	LUT2 #(
		.INIT('h4)
	) name24463 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_WbEn_q_reg/NET0131 ,
		_w34975_
	);
	LUT2 #(
		.INIT('h1)
	) name24464 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		_w34976_
	);
	LUT2 #(
		.INIT('h8)
	) name24465 (
		_w34975_,
		_w34976_,
		_w34977_
	);
	LUT2 #(
		.INIT('h2)
	) name24466 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w34978_
	);
	LUT2 #(
		.INIT('h4)
	) name24467 (
		\wishbone_WbEn_q_reg/NET0131 ,
		_w34978_,
		_w34979_
	);
	LUT2 #(
		.INIT('h1)
	) name24468 (
		_w34977_,
		_w34979_,
		_w34980_
	);
	LUT2 #(
		.INIT('h2)
	) name24469 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w34980_,
		_w34981_
	);
	LUT2 #(
		.INIT('h8)
	) name24470 (
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w34981_,
		_w34982_
	);
	LUT2 #(
		.INIT('h2)
	) name24471 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		\wishbone_RxEn_q_reg/NET0131 ,
		_w34983_
	);
	LUT2 #(
		.INIT('h8)
	) name24472 (
		_w34975_,
		_w34983_,
		_w34984_
	);
	LUT2 #(
		.INIT('h1)
	) name24473 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w34983_,
		_w34985_
	);
	LUT2 #(
		.INIT('h1)
	) name24474 (
		\wishbone_TxEn_q_reg/NET0131 ,
		_w34985_,
		_w34986_
	);
	LUT2 #(
		.INIT('h8)
	) name24475 (
		\wishbone_RxEn_q_reg/NET0131 ,
		\wishbone_TxEn_q_reg/NET0131 ,
		_w34987_
	);
	LUT2 #(
		.INIT('h1)
	) name24476 (
		\wishbone_WbEn_q_reg/NET0131 ,
		_w34987_,
		_w34988_
	);
	LUT2 #(
		.INIT('h4)
	) name24477 (
		_w34986_,
		_w34988_,
		_w34989_
	);
	LUT2 #(
		.INIT('h1)
	) name24478 (
		_w34981_,
		_w34989_,
		_w34990_
	);
	LUT2 #(
		.INIT('h4)
	) name24479 (
		_w34984_,
		_w34990_,
		_w34991_
	);
	LUT2 #(
		.INIT('h8)
	) name24480 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		_w34991_,
		_w34992_
	);
	LUT2 #(
		.INIT('h8)
	) name24481 (
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w34984_,
		_w34993_
	);
	LUT2 #(
		.INIT('h8)
	) name24482 (
		\wb_adr_i[2]_pad ,
		_w34989_,
		_w34994_
	);
	LUT2 #(
		.INIT('h1)
	) name24483 (
		_w34982_,
		_w34993_,
		_w34995_
	);
	LUT2 #(
		.INIT('h4)
	) name24484 (
		_w34994_,
		_w34995_,
		_w34996_
	);
	LUT2 #(
		.INIT('h4)
	) name24485 (
		_w34992_,
		_w34996_,
		_w34997_
	);
	LUT2 #(
		.INIT('h8)
	) name24486 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		_w34981_,
		_w34998_
	);
	LUT2 #(
		.INIT('h8)
	) name24487 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		_w34991_,
		_w34999_
	);
	LUT2 #(
		.INIT('h8)
	) name24488 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		_w34984_,
		_w35000_
	);
	LUT2 #(
		.INIT('h8)
	) name24489 (
		\wb_adr_i[3]_pad ,
		_w34989_,
		_w35001_
	);
	LUT2 #(
		.INIT('h1)
	) name24490 (
		_w34998_,
		_w35000_,
		_w35002_
	);
	LUT2 #(
		.INIT('h4)
	) name24491 (
		_w35001_,
		_w35002_,
		_w35003_
	);
	LUT2 #(
		.INIT('h4)
	) name24492 (
		_w34999_,
		_w35003_,
		_w35004_
	);
	LUT2 #(
		.INIT('h8)
	) name24493 (
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w34981_,
		_w35005_
	);
	LUT2 #(
		.INIT('h8)
	) name24494 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		_w34991_,
		_w35006_
	);
	LUT2 #(
		.INIT('h8)
	) name24495 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w34984_,
		_w35007_
	);
	LUT2 #(
		.INIT('h8)
	) name24496 (
		\wb_adr_i[4]_pad ,
		_w34989_,
		_w35008_
	);
	LUT2 #(
		.INIT('h1)
	) name24497 (
		_w35005_,
		_w35007_,
		_w35009_
	);
	LUT2 #(
		.INIT('h4)
	) name24498 (
		_w35008_,
		_w35009_,
		_w35010_
	);
	LUT2 #(
		.INIT('h4)
	) name24499 (
		_w35006_,
		_w35010_,
		_w35011_
	);
	LUT2 #(
		.INIT('h8)
	) name24500 (
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w34981_,
		_w35012_
	);
	LUT2 #(
		.INIT('h8)
	) name24501 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		_w34991_,
		_w35013_
	);
	LUT2 #(
		.INIT('h8)
	) name24502 (
		\wishbone_RxBDAddress_reg[3]/NET0131 ,
		_w34984_,
		_w35014_
	);
	LUT2 #(
		.INIT('h8)
	) name24503 (
		\wb_adr_i[5]_pad ,
		_w34989_,
		_w35015_
	);
	LUT2 #(
		.INIT('h1)
	) name24504 (
		_w35012_,
		_w35014_,
		_w35016_
	);
	LUT2 #(
		.INIT('h4)
	) name24505 (
		_w35015_,
		_w35016_,
		_w35017_
	);
	LUT2 #(
		.INIT('h4)
	) name24506 (
		_w35013_,
		_w35017_,
		_w35018_
	);
	LUT2 #(
		.INIT('h8)
	) name24507 (
		\wishbone_TxBDAddress_reg[4]/NET0131 ,
		_w34981_,
		_w35019_
	);
	LUT2 #(
		.INIT('h8)
	) name24508 (
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w34991_,
		_w35020_
	);
	LUT2 #(
		.INIT('h8)
	) name24509 (
		\wishbone_RxBDAddress_reg[4]/NET0131 ,
		_w34984_,
		_w35021_
	);
	LUT2 #(
		.INIT('h8)
	) name24510 (
		\wb_adr_i[6]_pad ,
		_w34989_,
		_w35022_
	);
	LUT2 #(
		.INIT('h1)
	) name24511 (
		_w35019_,
		_w35021_,
		_w35023_
	);
	LUT2 #(
		.INIT('h4)
	) name24512 (
		_w35022_,
		_w35023_,
		_w35024_
	);
	LUT2 #(
		.INIT('h4)
	) name24513 (
		_w35020_,
		_w35024_,
		_w35025_
	);
	LUT2 #(
		.INIT('h8)
	) name24514 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w34981_,
		_w35026_
	);
	LUT2 #(
		.INIT('h8)
	) name24515 (
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w34991_,
		_w35027_
	);
	LUT2 #(
		.INIT('h8)
	) name24516 (
		\wishbone_RxBDAddress_reg[5]/NET0131 ,
		_w34984_,
		_w35028_
	);
	LUT2 #(
		.INIT('h8)
	) name24517 (
		\wb_adr_i[7]_pad ,
		_w34989_,
		_w35029_
	);
	LUT2 #(
		.INIT('h1)
	) name24518 (
		_w35026_,
		_w35028_,
		_w35030_
	);
	LUT2 #(
		.INIT('h4)
	) name24519 (
		_w35029_,
		_w35030_,
		_w35031_
	);
	LUT2 #(
		.INIT('h4)
	) name24520 (
		_w35027_,
		_w35031_,
		_w35032_
	);
	LUT2 #(
		.INIT('h8)
	) name24521 (
		\wishbone_TxBDAddress_reg[6]/NET0131 ,
		_w34981_,
		_w35033_
	);
	LUT2 #(
		.INIT('h8)
	) name24522 (
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w34991_,
		_w35034_
	);
	LUT2 #(
		.INIT('h8)
	) name24523 (
		\wishbone_RxBDAddress_reg[6]/NET0131 ,
		_w34984_,
		_w35035_
	);
	LUT2 #(
		.INIT('h8)
	) name24524 (
		\wb_adr_i[8]_pad ,
		_w34989_,
		_w35036_
	);
	LUT2 #(
		.INIT('h1)
	) name24525 (
		_w35033_,
		_w35035_,
		_w35037_
	);
	LUT2 #(
		.INIT('h4)
	) name24526 (
		_w35036_,
		_w35037_,
		_w35038_
	);
	LUT2 #(
		.INIT('h4)
	) name24527 (
		_w35034_,
		_w35038_,
		_w35039_
	);
	LUT2 #(
		.INIT('h8)
	) name24528 (
		\wishbone_TxBDAddress_reg[7]/NET0131 ,
		_w34981_,
		_w35040_
	);
	LUT2 #(
		.INIT('h8)
	) name24529 (
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w34991_,
		_w35041_
	);
	LUT2 #(
		.INIT('h8)
	) name24530 (
		\wishbone_RxBDAddress_reg[7]/NET0131 ,
		_w34984_,
		_w35042_
	);
	LUT2 #(
		.INIT('h8)
	) name24531 (
		\wb_adr_i[9]_pad ,
		_w34989_,
		_w35043_
	);
	LUT2 #(
		.INIT('h1)
	) name24532 (
		_w35040_,
		_w35042_,
		_w35044_
	);
	LUT2 #(
		.INIT('h4)
	) name24533 (
		_w35043_,
		_w35044_,
		_w35045_
	);
	LUT2 #(
		.INIT('h4)
	) name24534 (
		_w35041_,
		_w35045_,
		_w35046_
	);
	LUT2 #(
		.INIT('h8)
	) name24535 (
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		_w34981_,
		_w35047_
	);
	LUT2 #(
		.INIT('h8)
	) name24536 (
		\wishbone_ram_di_reg[0]/NET0131 ,
		_w34991_,
		_w35048_
	);
	LUT2 #(
		.INIT('h8)
	) name24537 (
		\wishbone_RxStatusInLatched_reg[0]/NET0131 ,
		_w34984_,
		_w35049_
	);
	LUT2 #(
		.INIT('h8)
	) name24538 (
		\wb_dat_i[0]_pad ,
		_w34989_,
		_w35050_
	);
	LUT2 #(
		.INIT('h1)
	) name24539 (
		_w35047_,
		_w35049_,
		_w35051_
	);
	LUT2 #(
		.INIT('h4)
	) name24540 (
		_w35050_,
		_w35051_,
		_w35052_
	);
	LUT2 #(
		.INIT('h4)
	) name24541 (
		_w35048_,
		_w35052_,
		_w35053_
	);
	LUT2 #(
		.INIT('h8)
	) name24542 (
		\wishbone_TxStatus_reg[13]/NET0131 ,
		_w34981_,
		_w35054_
	);
	LUT2 #(
		.INIT('h8)
	) name24543 (
		\wishbone_ram_di_reg[13]/NET0131 ,
		_w34991_,
		_w35055_
	);
	LUT2 #(
		.INIT('h8)
	) name24544 (
		\wishbone_RxStatus_reg[13]/NET0131 ,
		_w34984_,
		_w35056_
	);
	LUT2 #(
		.INIT('h8)
	) name24545 (
		\wb_dat_i[13]_pad ,
		_w34989_,
		_w35057_
	);
	LUT2 #(
		.INIT('h1)
	) name24546 (
		_w35054_,
		_w35056_,
		_w35058_
	);
	LUT2 #(
		.INIT('h4)
	) name24547 (
		_w35057_,
		_w35058_,
		_w35059_
	);
	LUT2 #(
		.INIT('h4)
	) name24548 (
		_w35055_,
		_w35059_,
		_w35060_
	);
	LUT2 #(
		.INIT('h8)
	) name24549 (
		\wishbone_TxStatus_reg[14]/NET0131 ,
		_w34981_,
		_w35061_
	);
	LUT2 #(
		.INIT('h8)
	) name24550 (
		\wishbone_ram_di_reg[14]/NET0131 ,
		_w34991_,
		_w35062_
	);
	LUT2 #(
		.INIT('h8)
	) name24551 (
		\wishbone_RxStatus_reg[14]/NET0131 ,
		_w34984_,
		_w35063_
	);
	LUT2 #(
		.INIT('h8)
	) name24552 (
		\wb_dat_i[14]_pad ,
		_w34989_,
		_w35064_
	);
	LUT2 #(
		.INIT('h1)
	) name24553 (
		_w35061_,
		_w35063_,
		_w35065_
	);
	LUT2 #(
		.INIT('h4)
	) name24554 (
		_w35064_,
		_w35065_,
		_w35066_
	);
	LUT2 #(
		.INIT('h4)
	) name24555 (
		_w35062_,
		_w35066_,
		_w35067_
	);
	LUT2 #(
		.INIT('h8)
	) name24556 (
		\wb_dat_i[16]_pad ,
		_w34989_,
		_w35068_
	);
	LUT2 #(
		.INIT('h8)
	) name24557 (
		\wishbone_ram_di_reg[16]/NET0131 ,
		_w34991_,
		_w35069_
	);
	LUT2 #(
		.INIT('h8)
	) name24558 (
		\wishbone_LatchedRxLength_reg[0]/NET0131 ,
		_w34984_,
		_w35070_
	);
	LUT2 #(
		.INIT('h8)
	) name24559 (
		\wishbone_LatchedTxLength_reg[0]/NET0131 ,
		_w34981_,
		_w35071_
	);
	LUT2 #(
		.INIT('h1)
	) name24560 (
		_w35068_,
		_w35070_,
		_w35072_
	);
	LUT2 #(
		.INIT('h4)
	) name24561 (
		_w35071_,
		_w35072_,
		_w35073_
	);
	LUT2 #(
		.INIT('h4)
	) name24562 (
		_w35069_,
		_w35073_,
		_w35074_
	);
	LUT2 #(
		.INIT('h8)
	) name24563 (
		\wb_dat_i[17]_pad ,
		_w34989_,
		_w35075_
	);
	LUT2 #(
		.INIT('h8)
	) name24564 (
		\wishbone_ram_di_reg[17]/NET0131 ,
		_w34991_,
		_w35076_
	);
	LUT2 #(
		.INIT('h8)
	) name24565 (
		\wishbone_LatchedRxLength_reg[1]/NET0131 ,
		_w34984_,
		_w35077_
	);
	LUT2 #(
		.INIT('h8)
	) name24566 (
		\wishbone_LatchedTxLength_reg[1]/NET0131 ,
		_w34981_,
		_w35078_
	);
	LUT2 #(
		.INIT('h1)
	) name24567 (
		_w35075_,
		_w35077_,
		_w35079_
	);
	LUT2 #(
		.INIT('h4)
	) name24568 (
		_w35078_,
		_w35079_,
		_w35080_
	);
	LUT2 #(
		.INIT('h4)
	) name24569 (
		_w35076_,
		_w35080_,
		_w35081_
	);
	LUT2 #(
		.INIT('h8)
	) name24570 (
		\wb_dat_i[18]_pad ,
		_w34989_,
		_w35082_
	);
	LUT2 #(
		.INIT('h8)
	) name24571 (
		\wishbone_ram_di_reg[18]/NET0131 ,
		_w34991_,
		_w35083_
	);
	LUT2 #(
		.INIT('h8)
	) name24572 (
		\wishbone_LatchedRxLength_reg[2]/NET0131 ,
		_w34984_,
		_w35084_
	);
	LUT2 #(
		.INIT('h8)
	) name24573 (
		\wishbone_LatchedTxLength_reg[2]/NET0131 ,
		_w34981_,
		_w35085_
	);
	LUT2 #(
		.INIT('h1)
	) name24574 (
		_w35082_,
		_w35084_,
		_w35086_
	);
	LUT2 #(
		.INIT('h4)
	) name24575 (
		_w35085_,
		_w35086_,
		_w35087_
	);
	LUT2 #(
		.INIT('h4)
	) name24576 (
		_w35083_,
		_w35087_,
		_w35088_
	);
	LUT2 #(
		.INIT('h8)
	) name24577 (
		\wb_dat_i[19]_pad ,
		_w34989_,
		_w35089_
	);
	LUT2 #(
		.INIT('h8)
	) name24578 (
		\wishbone_ram_di_reg[19]/NET0131 ,
		_w34991_,
		_w35090_
	);
	LUT2 #(
		.INIT('h8)
	) name24579 (
		\wishbone_LatchedRxLength_reg[3]/NET0131 ,
		_w34984_,
		_w35091_
	);
	LUT2 #(
		.INIT('h8)
	) name24580 (
		\wishbone_LatchedTxLength_reg[3]/NET0131 ,
		_w34981_,
		_w35092_
	);
	LUT2 #(
		.INIT('h1)
	) name24581 (
		_w35089_,
		_w35091_,
		_w35093_
	);
	LUT2 #(
		.INIT('h4)
	) name24582 (
		_w35092_,
		_w35093_,
		_w35094_
	);
	LUT2 #(
		.INIT('h4)
	) name24583 (
		_w35090_,
		_w35094_,
		_w35095_
	);
	LUT2 #(
		.INIT('h8)
	) name24584 (
		\macstatus1_DeferLatched_reg/NET0131 ,
		_w34981_,
		_w35096_
	);
	LUT2 #(
		.INIT('h8)
	) name24585 (
		\wishbone_ram_di_reg[1]/NET0131 ,
		_w34991_,
		_w35097_
	);
	LUT2 #(
		.INIT('h8)
	) name24586 (
		\wishbone_RxStatusInLatched_reg[1]/NET0131 ,
		_w34984_,
		_w35098_
	);
	LUT2 #(
		.INIT('h8)
	) name24587 (
		\wb_dat_i[1]_pad ,
		_w34989_,
		_w35099_
	);
	LUT2 #(
		.INIT('h1)
	) name24588 (
		_w35096_,
		_w35098_,
		_w35100_
	);
	LUT2 #(
		.INIT('h4)
	) name24589 (
		_w35099_,
		_w35100_,
		_w35101_
	);
	LUT2 #(
		.INIT('h4)
	) name24590 (
		_w35097_,
		_w35101_,
		_w35102_
	);
	LUT2 #(
		.INIT('h8)
	) name24591 (
		\wb_dat_i[20]_pad ,
		_w34989_,
		_w35103_
	);
	LUT2 #(
		.INIT('h8)
	) name24592 (
		\wishbone_ram_di_reg[20]/NET0131 ,
		_w34991_,
		_w35104_
	);
	LUT2 #(
		.INIT('h8)
	) name24593 (
		\wishbone_LatchedRxLength_reg[4]/NET0131 ,
		_w34984_,
		_w35105_
	);
	LUT2 #(
		.INIT('h8)
	) name24594 (
		\wishbone_LatchedTxLength_reg[4]/NET0131 ,
		_w34981_,
		_w35106_
	);
	LUT2 #(
		.INIT('h1)
	) name24595 (
		_w35103_,
		_w35105_,
		_w35107_
	);
	LUT2 #(
		.INIT('h4)
	) name24596 (
		_w35106_,
		_w35107_,
		_w35108_
	);
	LUT2 #(
		.INIT('h4)
	) name24597 (
		_w35104_,
		_w35108_,
		_w35109_
	);
	LUT2 #(
		.INIT('h8)
	) name24598 (
		\wb_dat_i[21]_pad ,
		_w34989_,
		_w35110_
	);
	LUT2 #(
		.INIT('h8)
	) name24599 (
		\wishbone_ram_di_reg[21]/NET0131 ,
		_w34991_,
		_w35111_
	);
	LUT2 #(
		.INIT('h8)
	) name24600 (
		\wishbone_LatchedRxLength_reg[5]/NET0131 ,
		_w34984_,
		_w35112_
	);
	LUT2 #(
		.INIT('h8)
	) name24601 (
		\wishbone_LatchedTxLength_reg[5]/NET0131 ,
		_w34981_,
		_w35113_
	);
	LUT2 #(
		.INIT('h1)
	) name24602 (
		_w35110_,
		_w35112_,
		_w35114_
	);
	LUT2 #(
		.INIT('h4)
	) name24603 (
		_w35113_,
		_w35114_,
		_w35115_
	);
	LUT2 #(
		.INIT('h4)
	) name24604 (
		_w35111_,
		_w35115_,
		_w35116_
	);
	LUT2 #(
		.INIT('h8)
	) name24605 (
		\wb_dat_i[22]_pad ,
		_w34989_,
		_w35117_
	);
	LUT2 #(
		.INIT('h8)
	) name24606 (
		\wishbone_ram_di_reg[22]/NET0131 ,
		_w34991_,
		_w35118_
	);
	LUT2 #(
		.INIT('h8)
	) name24607 (
		\wishbone_LatchedRxLength_reg[6]/NET0131 ,
		_w34984_,
		_w35119_
	);
	LUT2 #(
		.INIT('h8)
	) name24608 (
		\wishbone_LatchedTxLength_reg[6]/NET0131 ,
		_w34981_,
		_w35120_
	);
	LUT2 #(
		.INIT('h1)
	) name24609 (
		_w35117_,
		_w35119_,
		_w35121_
	);
	LUT2 #(
		.INIT('h4)
	) name24610 (
		_w35120_,
		_w35121_,
		_w35122_
	);
	LUT2 #(
		.INIT('h4)
	) name24611 (
		_w35118_,
		_w35122_,
		_w35123_
	);
	LUT2 #(
		.INIT('h8)
	) name24612 (
		\wishbone_LatchedTxLength_reg[7]/NET0131 ,
		_w34981_,
		_w35124_
	);
	LUT2 #(
		.INIT('h8)
	) name24613 (
		\wishbone_ram_di_reg[23]/NET0131 ,
		_w34991_,
		_w35125_
	);
	LUT2 #(
		.INIT('h8)
	) name24614 (
		\wishbone_LatchedRxLength_reg[7]/NET0131 ,
		_w34984_,
		_w35126_
	);
	LUT2 #(
		.INIT('h8)
	) name24615 (
		\wb_dat_i[23]_pad ,
		_w34989_,
		_w35127_
	);
	LUT2 #(
		.INIT('h1)
	) name24616 (
		_w35124_,
		_w35126_,
		_w35128_
	);
	LUT2 #(
		.INIT('h4)
	) name24617 (
		_w35127_,
		_w35128_,
		_w35129_
	);
	LUT2 #(
		.INIT('h4)
	) name24618 (
		_w35125_,
		_w35129_,
		_w35130_
	);
	LUT2 #(
		.INIT('h8)
	) name24619 (
		\wishbone_LatchedTxLength_reg[8]/NET0131 ,
		_w34981_,
		_w35131_
	);
	LUT2 #(
		.INIT('h8)
	) name24620 (
		\wishbone_ram_di_reg[24]/NET0131 ,
		_w34991_,
		_w35132_
	);
	LUT2 #(
		.INIT('h8)
	) name24621 (
		\wishbone_LatchedRxLength_reg[8]/NET0131 ,
		_w34984_,
		_w35133_
	);
	LUT2 #(
		.INIT('h8)
	) name24622 (
		\wb_dat_i[24]_pad ,
		_w34989_,
		_w35134_
	);
	LUT2 #(
		.INIT('h1)
	) name24623 (
		_w35131_,
		_w35133_,
		_w35135_
	);
	LUT2 #(
		.INIT('h4)
	) name24624 (
		_w35134_,
		_w35135_,
		_w35136_
	);
	LUT2 #(
		.INIT('h4)
	) name24625 (
		_w35132_,
		_w35136_,
		_w35137_
	);
	LUT2 #(
		.INIT('h8)
	) name24626 (
		\wb_dat_i[25]_pad ,
		_w34989_,
		_w35138_
	);
	LUT2 #(
		.INIT('h8)
	) name24627 (
		\wishbone_ram_di_reg[25]/NET0131 ,
		_w34991_,
		_w35139_
	);
	LUT2 #(
		.INIT('h8)
	) name24628 (
		\wishbone_LatchedRxLength_reg[9]/NET0131 ,
		_w34984_,
		_w35140_
	);
	LUT2 #(
		.INIT('h8)
	) name24629 (
		\wishbone_LatchedTxLength_reg[9]/NET0131 ,
		_w34981_,
		_w35141_
	);
	LUT2 #(
		.INIT('h1)
	) name24630 (
		_w35138_,
		_w35140_,
		_w35142_
	);
	LUT2 #(
		.INIT('h4)
	) name24631 (
		_w35141_,
		_w35142_,
		_w35143_
	);
	LUT2 #(
		.INIT('h4)
	) name24632 (
		_w35139_,
		_w35143_,
		_w35144_
	);
	LUT2 #(
		.INIT('h8)
	) name24633 (
		\wb_dat_i[26]_pad ,
		_w34989_,
		_w35145_
	);
	LUT2 #(
		.INIT('h8)
	) name24634 (
		\wishbone_ram_di_reg[26]/NET0131 ,
		_w34991_,
		_w35146_
	);
	LUT2 #(
		.INIT('h8)
	) name24635 (
		\wishbone_LatchedRxLength_reg[10]/NET0131 ,
		_w34984_,
		_w35147_
	);
	LUT2 #(
		.INIT('h8)
	) name24636 (
		\wishbone_LatchedTxLength_reg[10]/NET0131 ,
		_w34981_,
		_w35148_
	);
	LUT2 #(
		.INIT('h1)
	) name24637 (
		_w35145_,
		_w35147_,
		_w35149_
	);
	LUT2 #(
		.INIT('h4)
	) name24638 (
		_w35148_,
		_w35149_,
		_w35150_
	);
	LUT2 #(
		.INIT('h4)
	) name24639 (
		_w35146_,
		_w35150_,
		_w35151_
	);
	LUT2 #(
		.INIT('h8)
	) name24640 (
		\wishbone_LatchedTxLength_reg[11]/NET0131 ,
		_w34981_,
		_w35152_
	);
	LUT2 #(
		.INIT('h8)
	) name24641 (
		\wishbone_ram_di_reg[27]/NET0131 ,
		_w34991_,
		_w35153_
	);
	LUT2 #(
		.INIT('h8)
	) name24642 (
		\wishbone_LatchedRxLength_reg[11]/NET0131 ,
		_w34984_,
		_w35154_
	);
	LUT2 #(
		.INIT('h8)
	) name24643 (
		\wb_dat_i[27]_pad ,
		_w34989_,
		_w35155_
	);
	LUT2 #(
		.INIT('h1)
	) name24644 (
		_w35152_,
		_w35154_,
		_w35156_
	);
	LUT2 #(
		.INIT('h4)
	) name24645 (
		_w35155_,
		_w35156_,
		_w35157_
	);
	LUT2 #(
		.INIT('h4)
	) name24646 (
		_w35153_,
		_w35157_,
		_w35158_
	);
	LUT2 #(
		.INIT('h8)
	) name24647 (
		\wb_dat_i[28]_pad ,
		_w34989_,
		_w35159_
	);
	LUT2 #(
		.INIT('h8)
	) name24648 (
		\wishbone_ram_di_reg[28]/NET0131 ,
		_w34991_,
		_w35160_
	);
	LUT2 #(
		.INIT('h8)
	) name24649 (
		\wishbone_LatchedRxLength_reg[12]/NET0131 ,
		_w34984_,
		_w35161_
	);
	LUT2 #(
		.INIT('h8)
	) name24650 (
		\wishbone_LatchedTxLength_reg[12]/NET0131 ,
		_w34981_,
		_w35162_
	);
	LUT2 #(
		.INIT('h1)
	) name24651 (
		_w35159_,
		_w35161_,
		_w35163_
	);
	LUT2 #(
		.INIT('h4)
	) name24652 (
		_w35162_,
		_w35163_,
		_w35164_
	);
	LUT2 #(
		.INIT('h4)
	) name24653 (
		_w35160_,
		_w35164_,
		_w35165_
	);
	LUT2 #(
		.INIT('h8)
	) name24654 (
		\wishbone_LatchedTxLength_reg[13]/NET0131 ,
		_w34981_,
		_w35166_
	);
	LUT2 #(
		.INIT('h8)
	) name24655 (
		\wishbone_ram_di_reg[29]/NET0131 ,
		_w34991_,
		_w35167_
	);
	LUT2 #(
		.INIT('h8)
	) name24656 (
		\wishbone_LatchedRxLength_reg[13]/NET0131 ,
		_w34984_,
		_w35168_
	);
	LUT2 #(
		.INIT('h8)
	) name24657 (
		\wb_dat_i[29]_pad ,
		_w34989_,
		_w35169_
	);
	LUT2 #(
		.INIT('h1)
	) name24658 (
		_w35166_,
		_w35168_,
		_w35170_
	);
	LUT2 #(
		.INIT('h4)
	) name24659 (
		_w35169_,
		_w35170_,
		_w35171_
	);
	LUT2 #(
		.INIT('h4)
	) name24660 (
		_w35167_,
		_w35171_,
		_w35172_
	);
	LUT2 #(
		.INIT('h8)
	) name24661 (
		\wb_dat_i[2]_pad ,
		_w34989_,
		_w35173_
	);
	LUT2 #(
		.INIT('h8)
	) name24662 (
		\wishbone_ram_di_reg[2]/NET0131 ,
		_w34991_,
		_w35174_
	);
	LUT2 #(
		.INIT('h8)
	) name24663 (
		\wishbone_RxStatusInLatched_reg[2]/NET0131 ,
		_w34984_,
		_w35175_
	);
	LUT2 #(
		.INIT('h8)
	) name24664 (
		\macstatus1_LateCollLatched_reg/P0002 ,
		_w34981_,
		_w35176_
	);
	LUT2 #(
		.INIT('h1)
	) name24665 (
		_w35173_,
		_w35175_,
		_w35177_
	);
	LUT2 #(
		.INIT('h4)
	) name24666 (
		_w35176_,
		_w35177_,
		_w35178_
	);
	LUT2 #(
		.INIT('h4)
	) name24667 (
		_w35174_,
		_w35178_,
		_w35179_
	);
	LUT2 #(
		.INIT('h8)
	) name24668 (
		\wb_dat_i[30]_pad ,
		_w34989_,
		_w35180_
	);
	LUT2 #(
		.INIT('h8)
	) name24669 (
		\wishbone_ram_di_reg[30]/NET0131 ,
		_w34991_,
		_w35181_
	);
	LUT2 #(
		.INIT('h8)
	) name24670 (
		\wishbone_LatchedRxLength_reg[14]/NET0131 ,
		_w34984_,
		_w35182_
	);
	LUT2 #(
		.INIT('h8)
	) name24671 (
		\wishbone_LatchedTxLength_reg[14]/NET0131 ,
		_w34981_,
		_w35183_
	);
	LUT2 #(
		.INIT('h1)
	) name24672 (
		_w35180_,
		_w35182_,
		_w35184_
	);
	LUT2 #(
		.INIT('h4)
	) name24673 (
		_w35183_,
		_w35184_,
		_w35185_
	);
	LUT2 #(
		.INIT('h4)
	) name24674 (
		_w35181_,
		_w35185_,
		_w35186_
	);
	LUT2 #(
		.INIT('h8)
	) name24675 (
		\wb_dat_i[31]_pad ,
		_w34989_,
		_w35187_
	);
	LUT2 #(
		.INIT('h8)
	) name24676 (
		\wishbone_ram_di_reg[31]/NET0131 ,
		_w34991_,
		_w35188_
	);
	LUT2 #(
		.INIT('h8)
	) name24677 (
		\wishbone_LatchedRxLength_reg[15]/NET0131 ,
		_w34984_,
		_w35189_
	);
	LUT2 #(
		.INIT('h8)
	) name24678 (
		\wishbone_LatchedTxLength_reg[15]/NET0131 ,
		_w34981_,
		_w35190_
	);
	LUT2 #(
		.INIT('h1)
	) name24679 (
		_w35187_,
		_w35189_,
		_w35191_
	);
	LUT2 #(
		.INIT('h4)
	) name24680 (
		_w35190_,
		_w35191_,
		_w35192_
	);
	LUT2 #(
		.INIT('h4)
	) name24681 (
		_w35188_,
		_w35192_,
		_w35193_
	);
	LUT2 #(
		.INIT('h8)
	) name24682 (
		\macstatus1_RetryLimit_reg/P0002 ,
		_w34981_,
		_w35194_
	);
	LUT2 #(
		.INIT('h8)
	) name24683 (
		\wishbone_ram_di_reg[3]/NET0131 ,
		_w34991_,
		_w35195_
	);
	LUT2 #(
		.INIT('h8)
	) name24684 (
		\wishbone_RxStatusInLatched_reg[3]/NET0131 ,
		_w34984_,
		_w35196_
	);
	LUT2 #(
		.INIT('h8)
	) name24685 (
		\wb_dat_i[3]_pad ,
		_w34989_,
		_w35197_
	);
	LUT2 #(
		.INIT('h1)
	) name24686 (
		_w35194_,
		_w35196_,
		_w35198_
	);
	LUT2 #(
		.INIT('h4)
	) name24687 (
		_w35197_,
		_w35198_,
		_w35199_
	);
	LUT2 #(
		.INIT('h4)
	) name24688 (
		_w35195_,
		_w35199_,
		_w35200_
	);
	LUT2 #(
		.INIT('h8)
	) name24689 (
		\wb_dat_i[4]_pad ,
		_w34989_,
		_w35201_
	);
	LUT2 #(
		.INIT('h8)
	) name24690 (
		\wishbone_ram_di_reg[4]/NET0131 ,
		_w34991_,
		_w35202_
	);
	LUT2 #(
		.INIT('h8)
	) name24691 (
		\wishbone_RxStatusInLatched_reg[4]/NET0131 ,
		_w34984_,
		_w35203_
	);
	LUT2 #(
		.INIT('h8)
	) name24692 (
		\macstatus1_RetryCntLatched_reg[0]/P0002 ,
		_w34981_,
		_w35204_
	);
	LUT2 #(
		.INIT('h1)
	) name24693 (
		_w35201_,
		_w35203_,
		_w35205_
	);
	LUT2 #(
		.INIT('h4)
	) name24694 (
		_w35204_,
		_w35205_,
		_w35206_
	);
	LUT2 #(
		.INIT('h4)
	) name24695 (
		_w35202_,
		_w35206_,
		_w35207_
	);
	LUT2 #(
		.INIT('h8)
	) name24696 (
		\wb_dat_i[5]_pad ,
		_w34989_,
		_w35208_
	);
	LUT2 #(
		.INIT('h8)
	) name24697 (
		\wishbone_ram_di_reg[5]/NET0131 ,
		_w34991_,
		_w35209_
	);
	LUT2 #(
		.INIT('h8)
	) name24698 (
		\wishbone_RxStatusInLatched_reg[5]/NET0131 ,
		_w34984_,
		_w35210_
	);
	LUT2 #(
		.INIT('h8)
	) name24699 (
		\macstatus1_RetryCntLatched_reg[1]/P0002 ,
		_w34981_,
		_w35211_
	);
	LUT2 #(
		.INIT('h1)
	) name24700 (
		_w35208_,
		_w35210_,
		_w35212_
	);
	LUT2 #(
		.INIT('h4)
	) name24701 (
		_w35211_,
		_w35212_,
		_w35213_
	);
	LUT2 #(
		.INIT('h4)
	) name24702 (
		_w35209_,
		_w35213_,
		_w35214_
	);
	LUT2 #(
		.INIT('h8)
	) name24703 (
		\wb_dat_i[6]_pad ,
		_w34989_,
		_w35215_
	);
	LUT2 #(
		.INIT('h8)
	) name24704 (
		\wishbone_ram_di_reg[6]/NET0131 ,
		_w34991_,
		_w35216_
	);
	LUT2 #(
		.INIT('h8)
	) name24705 (
		\wishbone_RxStatusInLatched_reg[6]/NET0131 ,
		_w34984_,
		_w35217_
	);
	LUT2 #(
		.INIT('h8)
	) name24706 (
		\macstatus1_RetryCntLatched_reg[2]/P0002 ,
		_w34981_,
		_w35218_
	);
	LUT2 #(
		.INIT('h1)
	) name24707 (
		_w35215_,
		_w35217_,
		_w35219_
	);
	LUT2 #(
		.INIT('h4)
	) name24708 (
		_w35218_,
		_w35219_,
		_w35220_
	);
	LUT2 #(
		.INIT('h4)
	) name24709 (
		_w35216_,
		_w35220_,
		_w35221_
	);
	LUT2 #(
		.INIT('h8)
	) name24710 (
		\wb_dat_i[7]_pad ,
		_w34989_,
		_w35222_
	);
	LUT2 #(
		.INIT('h8)
	) name24711 (
		\wishbone_ram_di_reg[7]/NET0131 ,
		_w34991_,
		_w35223_
	);
	LUT2 #(
		.INIT('h8)
	) name24712 (
		\wishbone_RxStatusInLatched_reg[7]/NET0131 ,
		_w34984_,
		_w35224_
	);
	LUT2 #(
		.INIT('h8)
	) name24713 (
		\macstatus1_RetryCntLatched_reg[3]/P0002 ,
		_w34981_,
		_w35225_
	);
	LUT2 #(
		.INIT('h1)
	) name24714 (
		_w35222_,
		_w35224_,
		_w35226_
	);
	LUT2 #(
		.INIT('h4)
	) name24715 (
		_w35225_,
		_w35226_,
		_w35227_
	);
	LUT2 #(
		.INIT('h4)
	) name24716 (
		_w35223_,
		_w35227_,
		_w35228_
	);
	LUT2 #(
		.INIT('h8)
	) name24717 (
		\wb_dat_i[8]_pad ,
		_w34989_,
		_w35229_
	);
	LUT2 #(
		.INIT('h8)
	) name24718 (
		\wishbone_ram_di_reg[8]/NET0131 ,
		_w34991_,
		_w35230_
	);
	LUT2 #(
		.INIT('h8)
	) name24719 (
		\wishbone_RxStatusInLatched_reg[8]/NET0131 ,
		_w34984_,
		_w35231_
	);
	LUT2 #(
		.INIT('h8)
	) name24720 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w34981_,
		_w35232_
	);
	LUT2 #(
		.INIT('h1)
	) name24721 (
		_w35229_,
		_w35231_,
		_w35233_
	);
	LUT2 #(
		.INIT('h4)
	) name24722 (
		_w35232_,
		_w35233_,
		_w35234_
	);
	LUT2 #(
		.INIT('h4)
	) name24723 (
		_w35230_,
		_w35234_,
		_w35235_
	);
	LUT2 #(
		.INIT('h2)
	) name24724 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		_w31950_,
		_w35236_
	);
	LUT2 #(
		.INIT('h4)
	) name24725 (
		_w34136_,
		_w35236_,
		_w35237_
	);
	LUT2 #(
		.INIT('h2)
	) name24726 (
		_w34136_,
		_w35236_,
		_w35238_
	);
	LUT2 #(
		.INIT('h1)
	) name24727 (
		_w35237_,
		_w35238_,
		_w35239_
	);
	LUT2 #(
		.INIT('h1)
	) name24728 (
		\wishbone_tx_fifo_write_pointer_reg[0]/NET0131 ,
		_w34447_,
		_w35240_
	);
	LUT2 #(
		.INIT('h2)
	) name24729 (
		_w33028_,
		_w34458_,
		_w35241_
	);
	LUT2 #(
		.INIT('h4)
	) name24730 (
		_w35240_,
		_w35241_,
		_w35242_
	);
	LUT2 #(
		.INIT('h1)
	) name24731 (
		_w34621_,
		_w35242_,
		_w35243_
	);
	LUT2 #(
		.INIT('h4)
	) name24732 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35244_
	);
	LUT2 #(
		.INIT('h4)
	) name24733 (
		_w31950_,
		_w34136_,
		_w35245_
	);
	LUT2 #(
		.INIT('h2)
	) name24734 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w35246_
	);
	LUT2 #(
		.INIT('h8)
	) name24735 (
		_w35245_,
		_w35246_,
		_w35247_
	);
	LUT2 #(
		.INIT('h8)
	) name24736 (
		_w35244_,
		_w35247_,
		_w35248_
	);
	LUT2 #(
		.INIT('h2)
	) name24737 (
		\wishbone_rx_fifo_fifo_reg[10][10]/P0001 ,
		_w35248_,
		_w35249_
	);
	LUT2 #(
		.INIT('h8)
	) name24738 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w35248_,
		_w35250_
	);
	LUT2 #(
		.INIT('h1)
	) name24739 (
		_w35249_,
		_w35250_,
		_w35251_
	);
	LUT2 #(
		.INIT('h2)
	) name24740 (
		\wishbone_rx_fifo_fifo_reg[10][12]/P0001 ,
		_w35248_,
		_w35252_
	);
	LUT2 #(
		.INIT('h8)
	) name24741 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		_w35248_,
		_w35253_
	);
	LUT2 #(
		.INIT('h1)
	) name24742 (
		_w35252_,
		_w35253_,
		_w35254_
	);
	LUT2 #(
		.INIT('h2)
	) name24743 (
		\wishbone_rx_fifo_fifo_reg[10][14]/P0001 ,
		_w35248_,
		_w35255_
	);
	LUT2 #(
		.INIT('h8)
	) name24744 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w35248_,
		_w35256_
	);
	LUT2 #(
		.INIT('h1)
	) name24745 (
		_w35255_,
		_w35256_,
		_w35257_
	);
	LUT2 #(
		.INIT('h2)
	) name24746 (
		\wishbone_rx_fifo_fifo_reg[10][16]/P0001 ,
		_w35248_,
		_w35258_
	);
	LUT2 #(
		.INIT('h8)
	) name24747 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w35248_,
		_w35259_
	);
	LUT2 #(
		.INIT('h1)
	) name24748 (
		_w35258_,
		_w35259_,
		_w35260_
	);
	LUT2 #(
		.INIT('h2)
	) name24749 (
		\wishbone_rx_fifo_fifo_reg[10][1]/P0001 ,
		_w35248_,
		_w35261_
	);
	LUT2 #(
		.INIT('h8)
	) name24750 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w35248_,
		_w35262_
	);
	LUT2 #(
		.INIT('h1)
	) name24751 (
		_w35261_,
		_w35262_,
		_w35263_
	);
	LUT2 #(
		.INIT('h2)
	) name24752 (
		\wishbone_rx_fifo_fifo_reg[10][20]/P0001 ,
		_w35248_,
		_w35264_
	);
	LUT2 #(
		.INIT('h8)
	) name24753 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		_w35248_,
		_w35265_
	);
	LUT2 #(
		.INIT('h1)
	) name24754 (
		_w35264_,
		_w35265_,
		_w35266_
	);
	LUT2 #(
		.INIT('h2)
	) name24755 (
		\wishbone_rx_fifo_fifo_reg[10][27]/P0001 ,
		_w35248_,
		_w35267_
	);
	LUT2 #(
		.INIT('h8)
	) name24756 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		_w35248_,
		_w35268_
	);
	LUT2 #(
		.INIT('h1)
	) name24757 (
		_w35267_,
		_w35268_,
		_w35269_
	);
	LUT2 #(
		.INIT('h2)
	) name24758 (
		\wishbone_rx_fifo_fifo_reg[10][28]/P0001 ,
		_w35248_,
		_w35270_
	);
	LUT2 #(
		.INIT('h8)
	) name24759 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		_w35248_,
		_w35271_
	);
	LUT2 #(
		.INIT('h1)
	) name24760 (
		_w35270_,
		_w35271_,
		_w35272_
	);
	LUT2 #(
		.INIT('h2)
	) name24761 (
		\wishbone_rx_fifo_fifo_reg[10][29]/P0001 ,
		_w35248_,
		_w35273_
	);
	LUT2 #(
		.INIT('h8)
	) name24762 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		_w35248_,
		_w35274_
	);
	LUT2 #(
		.INIT('h1)
	) name24763 (
		_w35273_,
		_w35274_,
		_w35275_
	);
	LUT2 #(
		.INIT('h2)
	) name24764 (
		\wishbone_rx_fifo_fifo_reg[10][31]/P0001 ,
		_w35248_,
		_w35276_
	);
	LUT2 #(
		.INIT('h8)
	) name24765 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		_w35248_,
		_w35277_
	);
	LUT2 #(
		.INIT('h1)
	) name24766 (
		_w35276_,
		_w35277_,
		_w35278_
	);
	LUT2 #(
		.INIT('h2)
	) name24767 (
		\wishbone_rx_fifo_fifo_reg[10][4]/P0001 ,
		_w35248_,
		_w35279_
	);
	LUT2 #(
		.INIT('h8)
	) name24768 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w35248_,
		_w35280_
	);
	LUT2 #(
		.INIT('h1)
	) name24769 (
		_w35279_,
		_w35280_,
		_w35281_
	);
	LUT2 #(
		.INIT('h2)
	) name24770 (
		\wishbone_rx_fifo_fifo_reg[10][5]/P0001 ,
		_w35248_,
		_w35282_
	);
	LUT2 #(
		.INIT('h8)
	) name24771 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		_w35248_,
		_w35283_
	);
	LUT2 #(
		.INIT('h1)
	) name24772 (
		_w35282_,
		_w35283_,
		_w35284_
	);
	LUT2 #(
		.INIT('h2)
	) name24773 (
		\wishbone_rx_fifo_fifo_reg[10][7]/P0001 ,
		_w35248_,
		_w35285_
	);
	LUT2 #(
		.INIT('h8)
	) name24774 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w35248_,
		_w35286_
	);
	LUT2 #(
		.INIT('h1)
	) name24775 (
		_w35285_,
		_w35286_,
		_w35287_
	);
	LUT2 #(
		.INIT('h2)
	) name24776 (
		\wishbone_rx_fifo_fifo_reg[10][9]/P0001 ,
		_w35248_,
		_w35288_
	);
	LUT2 #(
		.INIT('h8)
	) name24777 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w35248_,
		_w35289_
	);
	LUT2 #(
		.INIT('h1)
	) name24778 (
		_w35288_,
		_w35289_,
		_w35290_
	);
	LUT2 #(
		.INIT('h8)
	) name24779 (
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w35245_,
		_w35291_
	);
	LUT2 #(
		.INIT('h4)
	) name24780 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w35291_,
		_w35292_
	);
	LUT2 #(
		.INIT('h8)
	) name24781 (
		_w35244_,
		_w35292_,
		_w35293_
	);
	LUT2 #(
		.INIT('h2)
	) name24782 (
		\wishbone_rx_fifo_fifo_reg[12][11]/P0001 ,
		_w35293_,
		_w35294_
	);
	LUT2 #(
		.INIT('h8)
	) name24783 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		_w35293_,
		_w35295_
	);
	LUT2 #(
		.INIT('h1)
	) name24784 (
		_w35294_,
		_w35295_,
		_w35296_
	);
	LUT2 #(
		.INIT('h2)
	) name24785 (
		\wishbone_rx_fifo_fifo_reg[12][12]/P0001 ,
		_w35293_,
		_w35297_
	);
	LUT2 #(
		.INIT('h8)
	) name24786 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		_w35293_,
		_w35298_
	);
	LUT2 #(
		.INIT('h1)
	) name24787 (
		_w35297_,
		_w35298_,
		_w35299_
	);
	LUT2 #(
		.INIT('h2)
	) name24788 (
		\wishbone_rx_fifo_fifo_reg[12][14]/P0001 ,
		_w35293_,
		_w35300_
	);
	LUT2 #(
		.INIT('h8)
	) name24789 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w35293_,
		_w35301_
	);
	LUT2 #(
		.INIT('h1)
	) name24790 (
		_w35300_,
		_w35301_,
		_w35302_
	);
	LUT2 #(
		.INIT('h2)
	) name24791 (
		\wishbone_rx_fifo_fifo_reg[12][15]/P0001 ,
		_w35293_,
		_w35303_
	);
	LUT2 #(
		.INIT('h8)
	) name24792 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		_w35293_,
		_w35304_
	);
	LUT2 #(
		.INIT('h1)
	) name24793 (
		_w35303_,
		_w35304_,
		_w35305_
	);
	LUT2 #(
		.INIT('h2)
	) name24794 (
		\wishbone_rx_fifo_fifo_reg[12][16]/P0001 ,
		_w35293_,
		_w35306_
	);
	LUT2 #(
		.INIT('h8)
	) name24795 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w35293_,
		_w35307_
	);
	LUT2 #(
		.INIT('h1)
	) name24796 (
		_w35306_,
		_w35307_,
		_w35308_
	);
	LUT2 #(
		.INIT('h2)
	) name24797 (
		\wishbone_rx_fifo_fifo_reg[12][17]/P0001 ,
		_w35293_,
		_w35309_
	);
	LUT2 #(
		.INIT('h8)
	) name24798 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		_w35293_,
		_w35310_
	);
	LUT2 #(
		.INIT('h1)
	) name24799 (
		_w35309_,
		_w35310_,
		_w35311_
	);
	LUT2 #(
		.INIT('h2)
	) name24800 (
		\wishbone_rx_fifo_fifo_reg[12][19]/P0001 ,
		_w35293_,
		_w35312_
	);
	LUT2 #(
		.INIT('h8)
	) name24801 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w35293_,
		_w35313_
	);
	LUT2 #(
		.INIT('h1)
	) name24802 (
		_w35312_,
		_w35313_,
		_w35314_
	);
	LUT2 #(
		.INIT('h2)
	) name24803 (
		\wishbone_rx_fifo_fifo_reg[12][21]/P0001 ,
		_w35293_,
		_w35315_
	);
	LUT2 #(
		.INIT('h8)
	) name24804 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w35293_,
		_w35316_
	);
	LUT2 #(
		.INIT('h1)
	) name24805 (
		_w35315_,
		_w35316_,
		_w35317_
	);
	LUT2 #(
		.INIT('h2)
	) name24806 (
		\wishbone_rx_fifo_fifo_reg[12][22]/P0001 ,
		_w35293_,
		_w35318_
	);
	LUT2 #(
		.INIT('h8)
	) name24807 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w35293_,
		_w35319_
	);
	LUT2 #(
		.INIT('h1)
	) name24808 (
		_w35318_,
		_w35319_,
		_w35320_
	);
	LUT2 #(
		.INIT('h2)
	) name24809 (
		\wishbone_rx_fifo_fifo_reg[12][23]/P0001 ,
		_w35293_,
		_w35321_
	);
	LUT2 #(
		.INIT('h8)
	) name24810 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w35293_,
		_w35322_
	);
	LUT2 #(
		.INIT('h1)
	) name24811 (
		_w35321_,
		_w35322_,
		_w35323_
	);
	LUT2 #(
		.INIT('h2)
	) name24812 (
		\wishbone_rx_fifo_fifo_reg[12][24]/P0001 ,
		_w35293_,
		_w35324_
	);
	LUT2 #(
		.INIT('h8)
	) name24813 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		_w35293_,
		_w35325_
	);
	LUT2 #(
		.INIT('h1)
	) name24814 (
		_w35324_,
		_w35325_,
		_w35326_
	);
	LUT2 #(
		.INIT('h2)
	) name24815 (
		\wishbone_rx_fifo_fifo_reg[12][27]/P0001 ,
		_w35293_,
		_w35327_
	);
	LUT2 #(
		.INIT('h8)
	) name24816 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		_w35293_,
		_w35328_
	);
	LUT2 #(
		.INIT('h1)
	) name24817 (
		_w35327_,
		_w35328_,
		_w35329_
	);
	LUT2 #(
		.INIT('h2)
	) name24818 (
		\wishbone_rx_fifo_fifo_reg[12][28]/P0001 ,
		_w35293_,
		_w35330_
	);
	LUT2 #(
		.INIT('h8)
	) name24819 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		_w35293_,
		_w35331_
	);
	LUT2 #(
		.INIT('h1)
	) name24820 (
		_w35330_,
		_w35331_,
		_w35332_
	);
	LUT2 #(
		.INIT('h2)
	) name24821 (
		\wishbone_rx_fifo_fifo_reg[12][31]/P0001 ,
		_w35293_,
		_w35333_
	);
	LUT2 #(
		.INIT('h8)
	) name24822 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		_w35293_,
		_w35334_
	);
	LUT2 #(
		.INIT('h1)
	) name24823 (
		_w35333_,
		_w35334_,
		_w35335_
	);
	LUT2 #(
		.INIT('h2)
	) name24824 (
		\wishbone_rx_fifo_fifo_reg[12][4]/P0001 ,
		_w35293_,
		_w35336_
	);
	LUT2 #(
		.INIT('h8)
	) name24825 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w35293_,
		_w35337_
	);
	LUT2 #(
		.INIT('h1)
	) name24826 (
		_w35336_,
		_w35337_,
		_w35338_
	);
	LUT2 #(
		.INIT('h2)
	) name24827 (
		\wishbone_rx_fifo_fifo_reg[12][7]/P0001 ,
		_w35293_,
		_w35339_
	);
	LUT2 #(
		.INIT('h8)
	) name24828 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w35293_,
		_w35340_
	);
	LUT2 #(
		.INIT('h1)
	) name24829 (
		_w35339_,
		_w35340_,
		_w35341_
	);
	LUT2 #(
		.INIT('h2)
	) name24830 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35342_
	);
	LUT2 #(
		.INIT('h8)
	) name24831 (
		_w35247_,
		_w35342_,
		_w35343_
	);
	LUT2 #(
		.INIT('h2)
	) name24832 (
		\wishbone_rx_fifo_fifo_reg[3][10]/P0001 ,
		_w35343_,
		_w35344_
	);
	LUT2 #(
		.INIT('h8)
	) name24833 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w35343_,
		_w35345_
	);
	LUT2 #(
		.INIT('h1)
	) name24834 (
		_w35344_,
		_w35345_,
		_w35346_
	);
	LUT2 #(
		.INIT('h2)
	) name24835 (
		\wishbone_rx_fifo_fifo_reg[3][12]/P0001 ,
		_w35343_,
		_w35347_
	);
	LUT2 #(
		.INIT('h8)
	) name24836 (
		\wishbone_RxDataLatched2_reg[12]/NET0131 ,
		_w35343_,
		_w35348_
	);
	LUT2 #(
		.INIT('h1)
	) name24837 (
		_w35347_,
		_w35348_,
		_w35349_
	);
	LUT2 #(
		.INIT('h2)
	) name24838 (
		\wishbone_rx_fifo_fifo_reg[3][13]/P0001 ,
		_w35343_,
		_w35350_
	);
	LUT2 #(
		.INIT('h8)
	) name24839 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		_w35343_,
		_w35351_
	);
	LUT2 #(
		.INIT('h1)
	) name24840 (
		_w35350_,
		_w35351_,
		_w35352_
	);
	LUT2 #(
		.INIT('h2)
	) name24841 (
		\wishbone_rx_fifo_fifo_reg[3][14]/P0001 ,
		_w35343_,
		_w35353_
	);
	LUT2 #(
		.INIT('h8)
	) name24842 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w35343_,
		_w35354_
	);
	LUT2 #(
		.INIT('h1)
	) name24843 (
		_w35353_,
		_w35354_,
		_w35355_
	);
	LUT2 #(
		.INIT('h2)
	) name24844 (
		\wishbone_rx_fifo_fifo_reg[3][18]/P0001 ,
		_w35343_,
		_w35356_
	);
	LUT2 #(
		.INIT('h8)
	) name24845 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		_w35343_,
		_w35357_
	);
	LUT2 #(
		.INIT('h1)
	) name24846 (
		_w35356_,
		_w35357_,
		_w35358_
	);
	LUT2 #(
		.INIT('h2)
	) name24847 (
		\wishbone_rx_fifo_fifo_reg[3][19]/P0001 ,
		_w35343_,
		_w35359_
	);
	LUT2 #(
		.INIT('h8)
	) name24848 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w35343_,
		_w35360_
	);
	LUT2 #(
		.INIT('h1)
	) name24849 (
		_w35359_,
		_w35360_,
		_w35361_
	);
	LUT2 #(
		.INIT('h2)
	) name24850 (
		\wishbone_rx_fifo_fifo_reg[3][24]/P0001 ,
		_w35343_,
		_w35362_
	);
	LUT2 #(
		.INIT('h8)
	) name24851 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		_w35343_,
		_w35363_
	);
	LUT2 #(
		.INIT('h1)
	) name24852 (
		_w35362_,
		_w35363_,
		_w35364_
	);
	LUT2 #(
		.INIT('h2)
	) name24853 (
		\wishbone_rx_fifo_fifo_reg[3][26]/P0001 ,
		_w35343_,
		_w35365_
	);
	LUT2 #(
		.INIT('h8)
	) name24854 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		_w35343_,
		_w35366_
	);
	LUT2 #(
		.INIT('h1)
	) name24855 (
		_w35365_,
		_w35366_,
		_w35367_
	);
	LUT2 #(
		.INIT('h2)
	) name24856 (
		\wishbone_rx_fifo_fifo_reg[3][29]/P0001 ,
		_w35343_,
		_w35368_
	);
	LUT2 #(
		.INIT('h8)
	) name24857 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		_w35343_,
		_w35369_
	);
	LUT2 #(
		.INIT('h1)
	) name24858 (
		_w35368_,
		_w35369_,
		_w35370_
	);
	LUT2 #(
		.INIT('h2)
	) name24859 (
		\wishbone_rx_fifo_fifo_reg[3][28]/P0001 ,
		_w35343_,
		_w35371_
	);
	LUT2 #(
		.INIT('h8)
	) name24860 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		_w35343_,
		_w35372_
	);
	LUT2 #(
		.INIT('h1)
	) name24861 (
		_w35371_,
		_w35372_,
		_w35373_
	);
	LUT2 #(
		.INIT('h2)
	) name24862 (
		\wishbone_rx_fifo_fifo_reg[3][2]/P0001 ,
		_w35343_,
		_w35374_
	);
	LUT2 #(
		.INIT('h8)
	) name24863 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		_w35343_,
		_w35375_
	);
	LUT2 #(
		.INIT('h1)
	) name24864 (
		_w35374_,
		_w35375_,
		_w35376_
	);
	LUT2 #(
		.INIT('h2)
	) name24865 (
		\wishbone_rx_fifo_fifo_reg[3][30]/P0001 ,
		_w35343_,
		_w35377_
	);
	LUT2 #(
		.INIT('h8)
	) name24866 (
		\wishbone_RxDataLatched2_reg[30]/NET0131 ,
		_w35343_,
		_w35378_
	);
	LUT2 #(
		.INIT('h1)
	) name24867 (
		_w35377_,
		_w35378_,
		_w35379_
	);
	LUT2 #(
		.INIT('h2)
	) name24868 (
		\wishbone_rx_fifo_fifo_reg[3][31]/P0001 ,
		_w35343_,
		_w35380_
	);
	LUT2 #(
		.INIT('h8)
	) name24869 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		_w35343_,
		_w35381_
	);
	LUT2 #(
		.INIT('h1)
	) name24870 (
		_w35380_,
		_w35381_,
		_w35382_
	);
	LUT2 #(
		.INIT('h2)
	) name24871 (
		\wishbone_rx_fifo_fifo_reg[3][4]/P0001 ,
		_w35343_,
		_w35383_
	);
	LUT2 #(
		.INIT('h8)
	) name24872 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w35343_,
		_w35384_
	);
	LUT2 #(
		.INIT('h1)
	) name24873 (
		_w35383_,
		_w35384_,
		_w35385_
	);
	LUT2 #(
		.INIT('h2)
	) name24874 (
		\wishbone_rx_fifo_fifo_reg[3][7]/P0001 ,
		_w35343_,
		_w35386_
	);
	LUT2 #(
		.INIT('h8)
	) name24875 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w35343_,
		_w35387_
	);
	LUT2 #(
		.INIT('h1)
	) name24876 (
		_w35386_,
		_w35387_,
		_w35388_
	);
	LUT2 #(
		.INIT('h2)
	) name24877 (
		\wishbone_rx_fifo_fifo_reg[3][8]/P0001 ,
		_w35343_,
		_w35389_
	);
	LUT2 #(
		.INIT('h8)
	) name24878 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		_w35343_,
		_w35390_
	);
	LUT2 #(
		.INIT('h1)
	) name24879 (
		_w35389_,
		_w35390_,
		_w35391_
	);
	LUT2 #(
		.INIT('h2)
	) name24880 (
		\wishbone_rx_fifo_fifo_reg[3][9]/P0001 ,
		_w35343_,
		_w35392_
	);
	LUT2 #(
		.INIT('h8)
	) name24881 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w35343_,
		_w35393_
	);
	LUT2 #(
		.INIT('h1)
	) name24882 (
		_w35392_,
		_w35393_,
		_w35394_
	);
	LUT2 #(
		.INIT('h8)
	) name24883 (
		_w35292_,
		_w35342_,
		_w35395_
	);
	LUT2 #(
		.INIT('h2)
	) name24884 (
		\wishbone_rx_fifo_fifo_reg[5][10]/P0001 ,
		_w35395_,
		_w35396_
	);
	LUT2 #(
		.INIT('h8)
	) name24885 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w35395_,
		_w35397_
	);
	LUT2 #(
		.INIT('h1)
	) name24886 (
		_w35396_,
		_w35397_,
		_w35398_
	);
	LUT2 #(
		.INIT('h2)
	) name24887 (
		\wishbone_rx_fifo_fifo_reg[5][13]/P0001 ,
		_w35395_,
		_w35399_
	);
	LUT2 #(
		.INIT('h8)
	) name24888 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		_w35395_,
		_w35400_
	);
	LUT2 #(
		.INIT('h1)
	) name24889 (
		_w35399_,
		_w35400_,
		_w35401_
	);
	LUT2 #(
		.INIT('h2)
	) name24890 (
		\wishbone_rx_fifo_fifo_reg[5][15]/P0001 ,
		_w35395_,
		_w35402_
	);
	LUT2 #(
		.INIT('h8)
	) name24891 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		_w35395_,
		_w35403_
	);
	LUT2 #(
		.INIT('h1)
	) name24892 (
		_w35402_,
		_w35403_,
		_w35404_
	);
	LUT2 #(
		.INIT('h2)
	) name24893 (
		\wishbone_rx_fifo_fifo_reg[5][17]/P0001 ,
		_w35395_,
		_w35405_
	);
	LUT2 #(
		.INIT('h8)
	) name24894 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		_w35395_,
		_w35406_
	);
	LUT2 #(
		.INIT('h1)
	) name24895 (
		_w35405_,
		_w35406_,
		_w35407_
	);
	LUT2 #(
		.INIT('h2)
	) name24896 (
		\wishbone_rx_fifo_fifo_reg[5][19]/P0001 ,
		_w35395_,
		_w35408_
	);
	LUT2 #(
		.INIT('h8)
	) name24897 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w35395_,
		_w35409_
	);
	LUT2 #(
		.INIT('h1)
	) name24898 (
		_w35408_,
		_w35409_,
		_w35410_
	);
	LUT2 #(
		.INIT('h2)
	) name24899 (
		\wishbone_rx_fifo_fifo_reg[5][1]/P0001 ,
		_w35395_,
		_w35411_
	);
	LUT2 #(
		.INIT('h8)
	) name24900 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w35395_,
		_w35412_
	);
	LUT2 #(
		.INIT('h1)
	) name24901 (
		_w35411_,
		_w35412_,
		_w35413_
	);
	LUT2 #(
		.INIT('h2)
	) name24902 (
		\wishbone_rx_fifo_fifo_reg[5][21]/P0001 ,
		_w35395_,
		_w35414_
	);
	LUT2 #(
		.INIT('h8)
	) name24903 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w35395_,
		_w35415_
	);
	LUT2 #(
		.INIT('h1)
	) name24904 (
		_w35414_,
		_w35415_,
		_w35416_
	);
	LUT2 #(
		.INIT('h2)
	) name24905 (
		\wishbone_rx_fifo_fifo_reg[5][22]/P0001 ,
		_w35395_,
		_w35417_
	);
	LUT2 #(
		.INIT('h8)
	) name24906 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w35395_,
		_w35418_
	);
	LUT2 #(
		.INIT('h1)
	) name24907 (
		_w35417_,
		_w35418_,
		_w35419_
	);
	LUT2 #(
		.INIT('h2)
	) name24908 (
		\wishbone_rx_fifo_fifo_reg[5][20]/P0001 ,
		_w35395_,
		_w35420_
	);
	LUT2 #(
		.INIT('h8)
	) name24909 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		_w35395_,
		_w35421_
	);
	LUT2 #(
		.INIT('h1)
	) name24910 (
		_w35420_,
		_w35421_,
		_w35422_
	);
	LUT2 #(
		.INIT('h2)
	) name24911 (
		\wishbone_rx_fifo_fifo_reg[5][23]/P0001 ,
		_w35395_,
		_w35423_
	);
	LUT2 #(
		.INIT('h8)
	) name24912 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w35395_,
		_w35424_
	);
	LUT2 #(
		.INIT('h1)
	) name24913 (
		_w35423_,
		_w35424_,
		_w35425_
	);
	LUT2 #(
		.INIT('h2)
	) name24914 (
		\wishbone_rx_fifo_fifo_reg[5][24]/P0001 ,
		_w35395_,
		_w35426_
	);
	LUT2 #(
		.INIT('h8)
	) name24915 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		_w35395_,
		_w35427_
	);
	LUT2 #(
		.INIT('h1)
	) name24916 (
		_w35426_,
		_w35427_,
		_w35428_
	);
	LUT2 #(
		.INIT('h2)
	) name24917 (
		\wishbone_rx_fifo_fifo_reg[5][26]/P0001 ,
		_w35395_,
		_w35429_
	);
	LUT2 #(
		.INIT('h8)
	) name24918 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		_w35395_,
		_w35430_
	);
	LUT2 #(
		.INIT('h1)
	) name24919 (
		_w35429_,
		_w35430_,
		_w35431_
	);
	LUT2 #(
		.INIT('h2)
	) name24920 (
		\wishbone_rx_fifo_fifo_reg[5][28]/P0001 ,
		_w35395_,
		_w35432_
	);
	LUT2 #(
		.INIT('h8)
	) name24921 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		_w35395_,
		_w35433_
	);
	LUT2 #(
		.INIT('h1)
	) name24922 (
		_w35432_,
		_w35433_,
		_w35434_
	);
	LUT2 #(
		.INIT('h2)
	) name24923 (
		\wishbone_rx_fifo_fifo_reg[5][3]/P0001 ,
		_w35395_,
		_w35435_
	);
	LUT2 #(
		.INIT('h8)
	) name24924 (
		\wishbone_RxDataLatched2_reg[3]/NET0131 ,
		_w35395_,
		_w35436_
	);
	LUT2 #(
		.INIT('h1)
	) name24925 (
		_w35435_,
		_w35436_,
		_w35437_
	);
	LUT2 #(
		.INIT('h2)
	) name24926 (
		\wishbone_rx_fifo_fifo_reg[5][6]/P0001 ,
		_w35395_,
		_w35438_
	);
	LUT2 #(
		.INIT('h8)
	) name24927 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		_w35395_,
		_w35439_
	);
	LUT2 #(
		.INIT('h1)
	) name24928 (
		_w35438_,
		_w35439_,
		_w35440_
	);
	LUT2 #(
		.INIT('h2)
	) name24929 (
		\wishbone_rx_fifo_fifo_reg[5][8]/P0001 ,
		_w35395_,
		_w35441_
	);
	LUT2 #(
		.INIT('h8)
	) name24930 (
		\wishbone_RxDataLatched2_reg[8]/NET0131 ,
		_w35395_,
		_w35442_
	);
	LUT2 #(
		.INIT('h1)
	) name24931 (
		_w35441_,
		_w35442_,
		_w35443_
	);
	LUT2 #(
		.INIT('h1)
	) name24932 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35444_
	);
	LUT2 #(
		.INIT('h8)
	) name24933 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w35291_,
		_w35445_
	);
	LUT2 #(
		.INIT('h8)
	) name24934 (
		_w35444_,
		_w35445_,
		_w35446_
	);
	LUT2 #(
		.INIT('h2)
	) name24935 (
		\wishbone_rx_fifo_fifo_reg[6][0]/P0001 ,
		_w35446_,
		_w35447_
	);
	LUT2 #(
		.INIT('h8)
	) name24936 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		_w35446_,
		_w35448_
	);
	LUT2 #(
		.INIT('h1)
	) name24937 (
		_w35447_,
		_w35448_,
		_w35449_
	);
	LUT2 #(
		.INIT('h2)
	) name24938 (
		\wishbone_rx_fifo_fifo_reg[6][10]/P0001 ,
		_w35446_,
		_w35450_
	);
	LUT2 #(
		.INIT('h8)
	) name24939 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w35446_,
		_w35451_
	);
	LUT2 #(
		.INIT('h1)
	) name24940 (
		_w35450_,
		_w35451_,
		_w35452_
	);
	LUT2 #(
		.INIT('h2)
	) name24941 (
		\wishbone_rx_fifo_fifo_reg[6][11]/P0001 ,
		_w35446_,
		_w35453_
	);
	LUT2 #(
		.INIT('h8)
	) name24942 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		_w35446_,
		_w35454_
	);
	LUT2 #(
		.INIT('h1)
	) name24943 (
		_w35453_,
		_w35454_,
		_w35455_
	);
	LUT2 #(
		.INIT('h2)
	) name24944 (
		\wishbone_rx_fifo_fifo_reg[6][14]/P0001 ,
		_w35446_,
		_w35456_
	);
	LUT2 #(
		.INIT('h8)
	) name24945 (
		\wishbone_RxDataLatched2_reg[14]/NET0131 ,
		_w35446_,
		_w35457_
	);
	LUT2 #(
		.INIT('h1)
	) name24946 (
		_w35456_,
		_w35457_,
		_w35458_
	);
	LUT2 #(
		.INIT('h2)
	) name24947 (
		\wishbone_rx_fifo_fifo_reg[6][15]/P0001 ,
		_w35446_,
		_w35459_
	);
	LUT2 #(
		.INIT('h8)
	) name24948 (
		\wishbone_RxDataLatched2_reg[15]/NET0131 ,
		_w35446_,
		_w35460_
	);
	LUT2 #(
		.INIT('h1)
	) name24949 (
		_w35459_,
		_w35460_,
		_w35461_
	);
	LUT2 #(
		.INIT('h2)
	) name24950 (
		\wishbone_rx_fifo_fifo_reg[6][16]/P0001 ,
		_w35446_,
		_w35462_
	);
	LUT2 #(
		.INIT('h8)
	) name24951 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w35446_,
		_w35463_
	);
	LUT2 #(
		.INIT('h1)
	) name24952 (
		_w35462_,
		_w35463_,
		_w35464_
	);
	LUT2 #(
		.INIT('h2)
	) name24953 (
		\wishbone_rx_fifo_fifo_reg[6][18]/P0001 ,
		_w35446_,
		_w35465_
	);
	LUT2 #(
		.INIT('h8)
	) name24954 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		_w35446_,
		_w35466_
	);
	LUT2 #(
		.INIT('h1)
	) name24955 (
		_w35465_,
		_w35466_,
		_w35467_
	);
	LUT2 #(
		.INIT('h2)
	) name24956 (
		\wishbone_rx_fifo_fifo_reg[6][19]/P0001 ,
		_w35446_,
		_w35468_
	);
	LUT2 #(
		.INIT('h8)
	) name24957 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w35446_,
		_w35469_
	);
	LUT2 #(
		.INIT('h1)
	) name24958 (
		_w35468_,
		_w35469_,
		_w35470_
	);
	LUT2 #(
		.INIT('h2)
	) name24959 (
		\wishbone_rx_fifo_fifo_reg[6][1]/P0001 ,
		_w35446_,
		_w35471_
	);
	LUT2 #(
		.INIT('h8)
	) name24960 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w35446_,
		_w35472_
	);
	LUT2 #(
		.INIT('h1)
	) name24961 (
		_w35471_,
		_w35472_,
		_w35473_
	);
	LUT2 #(
		.INIT('h2)
	) name24962 (
		\wishbone_rx_fifo_fifo_reg[6][21]/P0001 ,
		_w35446_,
		_w35474_
	);
	LUT2 #(
		.INIT('h8)
	) name24963 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w35446_,
		_w35475_
	);
	LUT2 #(
		.INIT('h1)
	) name24964 (
		_w35474_,
		_w35475_,
		_w35476_
	);
	LUT2 #(
		.INIT('h2)
	) name24965 (
		\wishbone_rx_fifo_fifo_reg[6][22]/P0001 ,
		_w35446_,
		_w35477_
	);
	LUT2 #(
		.INIT('h8)
	) name24966 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w35446_,
		_w35478_
	);
	LUT2 #(
		.INIT('h1)
	) name24967 (
		_w35477_,
		_w35478_,
		_w35479_
	);
	LUT2 #(
		.INIT('h2)
	) name24968 (
		\wishbone_rx_fifo_fifo_reg[6][23]/P0001 ,
		_w35446_,
		_w35480_
	);
	LUT2 #(
		.INIT('h8)
	) name24969 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w35446_,
		_w35481_
	);
	LUT2 #(
		.INIT('h1)
	) name24970 (
		_w35480_,
		_w35481_,
		_w35482_
	);
	LUT2 #(
		.INIT('h2)
	) name24971 (
		\wishbone_rx_fifo_fifo_reg[6][25]/P0001 ,
		_w35446_,
		_w35483_
	);
	LUT2 #(
		.INIT('h8)
	) name24972 (
		\wishbone_RxDataLatched2_reg[25]/NET0131 ,
		_w35446_,
		_w35484_
	);
	LUT2 #(
		.INIT('h1)
	) name24973 (
		_w35483_,
		_w35484_,
		_w35485_
	);
	LUT2 #(
		.INIT('h2)
	) name24974 (
		\wishbone_rx_fifo_fifo_reg[6][26]/P0001 ,
		_w35446_,
		_w35486_
	);
	LUT2 #(
		.INIT('h8)
	) name24975 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		_w35446_,
		_w35487_
	);
	LUT2 #(
		.INIT('h1)
	) name24976 (
		_w35486_,
		_w35487_,
		_w35488_
	);
	LUT2 #(
		.INIT('h2)
	) name24977 (
		\wishbone_rx_fifo_fifo_reg[6][24]/P0001 ,
		_w35446_,
		_w35489_
	);
	LUT2 #(
		.INIT('h8)
	) name24978 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		_w35446_,
		_w35490_
	);
	LUT2 #(
		.INIT('h1)
	) name24979 (
		_w35489_,
		_w35490_,
		_w35491_
	);
	LUT2 #(
		.INIT('h2)
	) name24980 (
		\wishbone_rx_fifo_fifo_reg[6][27]/P0001 ,
		_w35446_,
		_w35492_
	);
	LUT2 #(
		.INIT('h8)
	) name24981 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		_w35446_,
		_w35493_
	);
	LUT2 #(
		.INIT('h1)
	) name24982 (
		_w35492_,
		_w35493_,
		_w35494_
	);
	LUT2 #(
		.INIT('h2)
	) name24983 (
		\wishbone_rx_fifo_fifo_reg[6][28]/P0001 ,
		_w35446_,
		_w35495_
	);
	LUT2 #(
		.INIT('h8)
	) name24984 (
		\wishbone_RxDataLatched2_reg[28]/NET0131 ,
		_w35446_,
		_w35496_
	);
	LUT2 #(
		.INIT('h1)
	) name24985 (
		_w35495_,
		_w35496_,
		_w35497_
	);
	LUT2 #(
		.INIT('h2)
	) name24986 (
		\wishbone_rx_fifo_fifo_reg[6][2]/P0001 ,
		_w35446_,
		_w35498_
	);
	LUT2 #(
		.INIT('h8)
	) name24987 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		_w35446_,
		_w35499_
	);
	LUT2 #(
		.INIT('h1)
	) name24988 (
		_w35498_,
		_w35499_,
		_w35500_
	);
	LUT2 #(
		.INIT('h2)
	) name24989 (
		\wishbone_rx_fifo_fifo_reg[6][31]/P0001 ,
		_w35446_,
		_w35501_
	);
	LUT2 #(
		.INIT('h8)
	) name24990 (
		\wishbone_RxDataLatched2_reg[31]/NET0131 ,
		_w35446_,
		_w35502_
	);
	LUT2 #(
		.INIT('h1)
	) name24991 (
		_w35501_,
		_w35502_,
		_w35503_
	);
	LUT2 #(
		.INIT('h2)
	) name24992 (
		\wishbone_rx_fifo_fifo_reg[6][5]/P0001 ,
		_w35446_,
		_w35504_
	);
	LUT2 #(
		.INIT('h8)
	) name24993 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		_w35446_,
		_w35505_
	);
	LUT2 #(
		.INIT('h1)
	) name24994 (
		_w35504_,
		_w35505_,
		_w35506_
	);
	LUT2 #(
		.INIT('h2)
	) name24995 (
		\wishbone_rx_fifo_fifo_reg[6][6]/P0001 ,
		_w35446_,
		_w35507_
	);
	LUT2 #(
		.INIT('h8)
	) name24996 (
		\wishbone_RxDataLatched2_reg[6]/NET0131 ,
		_w35446_,
		_w35508_
	);
	LUT2 #(
		.INIT('h1)
	) name24997 (
		_w35507_,
		_w35508_,
		_w35509_
	);
	LUT2 #(
		.INIT('h2)
	) name24998 (
		\wishbone_rx_fifo_fifo_reg[6][7]/P0001 ,
		_w35446_,
		_w35510_
	);
	LUT2 #(
		.INIT('h8)
	) name24999 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w35446_,
		_w35511_
	);
	LUT2 #(
		.INIT('h1)
	) name25000 (
		_w35510_,
		_w35511_,
		_w35512_
	);
	LUT2 #(
		.INIT('h2)
	) name25001 (
		\wishbone_rx_fifo_fifo_reg[6][9]/P0001 ,
		_w35446_,
		_w35513_
	);
	LUT2 #(
		.INIT('h8)
	) name25002 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w35446_,
		_w35514_
	);
	LUT2 #(
		.INIT('h1)
	) name25003 (
		_w35513_,
		_w35514_,
		_w35515_
	);
	LUT2 #(
		.INIT('h1)
	) name25004 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w35516_
	);
	LUT2 #(
		.INIT('h8)
	) name25005 (
		_w34136_,
		_w35516_,
		_w35517_
	);
	LUT2 #(
		.INIT('h8)
	) name25006 (
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35236_,
		_w35518_
	);
	LUT2 #(
		.INIT('h8)
	) name25007 (
		_w35517_,
		_w35518_,
		_w35519_
	);
	LUT2 #(
		.INIT('h2)
	) name25008 (
		\wishbone_rx_fifo_fifo_reg[9][0]/P0001 ,
		_w35519_,
		_w35520_
	);
	LUT2 #(
		.INIT('h8)
	) name25009 (
		\wishbone_RxDataLatched2_reg[0]/NET0131 ,
		_w35519_,
		_w35521_
	);
	LUT2 #(
		.INIT('h1)
	) name25010 (
		_w35520_,
		_w35521_,
		_w35522_
	);
	LUT2 #(
		.INIT('h2)
	) name25011 (
		\wishbone_rx_fifo_fifo_reg[9][10]/P0001 ,
		_w35519_,
		_w35523_
	);
	LUT2 #(
		.INIT('h8)
	) name25012 (
		\wishbone_RxDataLatched2_reg[10]/NET0131 ,
		_w35519_,
		_w35524_
	);
	LUT2 #(
		.INIT('h1)
	) name25013 (
		_w35523_,
		_w35524_,
		_w35525_
	);
	LUT2 #(
		.INIT('h2)
	) name25014 (
		\wishbone_rx_fifo_fifo_reg[9][11]/P0001 ,
		_w35519_,
		_w35526_
	);
	LUT2 #(
		.INIT('h8)
	) name25015 (
		\wishbone_RxDataLatched2_reg[11]/NET0131 ,
		_w35519_,
		_w35527_
	);
	LUT2 #(
		.INIT('h1)
	) name25016 (
		_w35526_,
		_w35527_,
		_w35528_
	);
	LUT2 #(
		.INIT('h2)
	) name25017 (
		\wishbone_rx_fifo_fifo_reg[9][13]/P0001 ,
		_w35519_,
		_w35529_
	);
	LUT2 #(
		.INIT('h8)
	) name25018 (
		\wishbone_RxDataLatched2_reg[13]/NET0131 ,
		_w35519_,
		_w35530_
	);
	LUT2 #(
		.INIT('h1)
	) name25019 (
		_w35529_,
		_w35530_,
		_w35531_
	);
	LUT2 #(
		.INIT('h2)
	) name25020 (
		\wishbone_rx_fifo_fifo_reg[9][16]/P0001 ,
		_w35519_,
		_w35532_
	);
	LUT2 #(
		.INIT('h8)
	) name25021 (
		\wishbone_RxDataLatched2_reg[16]/NET0131 ,
		_w35519_,
		_w35533_
	);
	LUT2 #(
		.INIT('h1)
	) name25022 (
		_w35532_,
		_w35533_,
		_w35534_
	);
	LUT2 #(
		.INIT('h2)
	) name25023 (
		\wishbone_rx_fifo_fifo_reg[9][17]/P0001 ,
		_w35519_,
		_w35535_
	);
	LUT2 #(
		.INIT('h8)
	) name25024 (
		\wishbone_RxDataLatched2_reg[17]/NET0131 ,
		_w35519_,
		_w35536_
	);
	LUT2 #(
		.INIT('h1)
	) name25025 (
		_w35535_,
		_w35536_,
		_w35537_
	);
	LUT2 #(
		.INIT('h2)
	) name25026 (
		\wishbone_rx_fifo_fifo_reg[9][18]/P0001 ,
		_w35519_,
		_w35538_
	);
	LUT2 #(
		.INIT('h8)
	) name25027 (
		\wishbone_RxDataLatched2_reg[18]/NET0131 ,
		_w35519_,
		_w35539_
	);
	LUT2 #(
		.INIT('h1)
	) name25028 (
		_w35538_,
		_w35539_,
		_w35540_
	);
	LUT2 #(
		.INIT('h2)
	) name25029 (
		\wishbone_rx_fifo_fifo_reg[9][19]/P0001 ,
		_w35519_,
		_w35541_
	);
	LUT2 #(
		.INIT('h8)
	) name25030 (
		\wishbone_RxDataLatched2_reg[19]/NET0131 ,
		_w35519_,
		_w35542_
	);
	LUT2 #(
		.INIT('h1)
	) name25031 (
		_w35541_,
		_w35542_,
		_w35543_
	);
	LUT2 #(
		.INIT('h2)
	) name25032 (
		\wishbone_rx_fifo_fifo_reg[9][1]/P0001 ,
		_w35519_,
		_w35544_
	);
	LUT2 #(
		.INIT('h8)
	) name25033 (
		\wishbone_RxDataLatched2_reg[1]/NET0131 ,
		_w35519_,
		_w35545_
	);
	LUT2 #(
		.INIT('h1)
	) name25034 (
		_w35544_,
		_w35545_,
		_w35546_
	);
	LUT2 #(
		.INIT('h2)
	) name25035 (
		\wishbone_rx_fifo_fifo_reg[9][20]/P0001 ,
		_w35519_,
		_w35547_
	);
	LUT2 #(
		.INIT('h8)
	) name25036 (
		\wishbone_RxDataLatched2_reg[20]/NET0131 ,
		_w35519_,
		_w35548_
	);
	LUT2 #(
		.INIT('h1)
	) name25037 (
		_w35547_,
		_w35548_,
		_w35549_
	);
	LUT2 #(
		.INIT('h2)
	) name25038 (
		\wishbone_rx_fifo_fifo_reg[9][21]/P0001 ,
		_w35519_,
		_w35550_
	);
	LUT2 #(
		.INIT('h8)
	) name25039 (
		\wishbone_RxDataLatched2_reg[21]/NET0131 ,
		_w35519_,
		_w35551_
	);
	LUT2 #(
		.INIT('h1)
	) name25040 (
		_w35550_,
		_w35551_,
		_w35552_
	);
	LUT2 #(
		.INIT('h2)
	) name25041 (
		\wishbone_rx_fifo_fifo_reg[9][22]/P0001 ,
		_w35519_,
		_w35553_
	);
	LUT2 #(
		.INIT('h8)
	) name25042 (
		\wishbone_RxDataLatched2_reg[22]/NET0131 ,
		_w35519_,
		_w35554_
	);
	LUT2 #(
		.INIT('h1)
	) name25043 (
		_w35553_,
		_w35554_,
		_w35555_
	);
	LUT2 #(
		.INIT('h2)
	) name25044 (
		\wishbone_rx_fifo_fifo_reg[9][23]/P0001 ,
		_w35519_,
		_w35556_
	);
	LUT2 #(
		.INIT('h8)
	) name25045 (
		\wishbone_RxDataLatched2_reg[23]/NET0131 ,
		_w35519_,
		_w35557_
	);
	LUT2 #(
		.INIT('h1)
	) name25046 (
		_w35556_,
		_w35557_,
		_w35558_
	);
	LUT2 #(
		.INIT('h2)
	) name25047 (
		\wishbone_rx_fifo_fifo_reg[9][24]/P0001 ,
		_w35519_,
		_w35559_
	);
	LUT2 #(
		.INIT('h8)
	) name25048 (
		\wishbone_RxDataLatched2_reg[24]/NET0131 ,
		_w35519_,
		_w35560_
	);
	LUT2 #(
		.INIT('h1)
	) name25049 (
		_w35559_,
		_w35560_,
		_w35561_
	);
	LUT2 #(
		.INIT('h2)
	) name25050 (
		\wishbone_rx_fifo_fifo_reg[9][25]/P0001 ,
		_w35519_,
		_w35562_
	);
	LUT2 #(
		.INIT('h8)
	) name25051 (
		\wishbone_RxDataLatched2_reg[25]/NET0131 ,
		_w35519_,
		_w35563_
	);
	LUT2 #(
		.INIT('h1)
	) name25052 (
		_w35562_,
		_w35563_,
		_w35564_
	);
	LUT2 #(
		.INIT('h2)
	) name25053 (
		\wishbone_rx_fifo_fifo_reg[9][26]/P0001 ,
		_w35519_,
		_w35565_
	);
	LUT2 #(
		.INIT('h8)
	) name25054 (
		\wishbone_RxDataLatched2_reg[26]/NET0131 ,
		_w35519_,
		_w35566_
	);
	LUT2 #(
		.INIT('h1)
	) name25055 (
		_w35565_,
		_w35566_,
		_w35567_
	);
	LUT2 #(
		.INIT('h2)
	) name25056 (
		\wishbone_rx_fifo_fifo_reg[9][27]/P0001 ,
		_w35519_,
		_w35568_
	);
	LUT2 #(
		.INIT('h8)
	) name25057 (
		\wishbone_RxDataLatched2_reg[27]/NET0131 ,
		_w35519_,
		_w35569_
	);
	LUT2 #(
		.INIT('h1)
	) name25058 (
		_w35568_,
		_w35569_,
		_w35570_
	);
	LUT2 #(
		.INIT('h2)
	) name25059 (
		\wishbone_rx_fifo_fifo_reg[9][29]/P0001 ,
		_w35519_,
		_w35571_
	);
	LUT2 #(
		.INIT('h8)
	) name25060 (
		\wishbone_RxDataLatched2_reg[29]/NET0131 ,
		_w35519_,
		_w35572_
	);
	LUT2 #(
		.INIT('h1)
	) name25061 (
		_w35571_,
		_w35572_,
		_w35573_
	);
	LUT2 #(
		.INIT('h2)
	) name25062 (
		\wishbone_rx_fifo_fifo_reg[9][2]/P0001 ,
		_w35519_,
		_w35574_
	);
	LUT2 #(
		.INIT('h8)
	) name25063 (
		\wishbone_RxDataLatched2_reg[2]/NET0131 ,
		_w35519_,
		_w35575_
	);
	LUT2 #(
		.INIT('h1)
	) name25064 (
		_w35574_,
		_w35575_,
		_w35576_
	);
	LUT2 #(
		.INIT('h2)
	) name25065 (
		\wishbone_rx_fifo_fifo_reg[9][30]/P0001 ,
		_w35519_,
		_w35577_
	);
	LUT2 #(
		.INIT('h8)
	) name25066 (
		\wishbone_RxDataLatched2_reg[30]/NET0131 ,
		_w35519_,
		_w35578_
	);
	LUT2 #(
		.INIT('h1)
	) name25067 (
		_w35577_,
		_w35578_,
		_w35579_
	);
	LUT2 #(
		.INIT('h2)
	) name25068 (
		\wishbone_rx_fifo_fifo_reg[9][4]/P0001 ,
		_w35519_,
		_w35580_
	);
	LUT2 #(
		.INIT('h8)
	) name25069 (
		\wishbone_RxDataLatched2_reg[4]/NET0131 ,
		_w35519_,
		_w35581_
	);
	LUT2 #(
		.INIT('h1)
	) name25070 (
		_w35580_,
		_w35581_,
		_w35582_
	);
	LUT2 #(
		.INIT('h2)
	) name25071 (
		\wishbone_rx_fifo_fifo_reg[9][5]/P0001 ,
		_w35519_,
		_w35583_
	);
	LUT2 #(
		.INIT('h8)
	) name25072 (
		\wishbone_RxDataLatched2_reg[5]/NET0131 ,
		_w35519_,
		_w35584_
	);
	LUT2 #(
		.INIT('h1)
	) name25073 (
		_w35583_,
		_w35584_,
		_w35585_
	);
	LUT2 #(
		.INIT('h2)
	) name25074 (
		\wishbone_rx_fifo_fifo_reg[9][7]/P0001 ,
		_w35519_,
		_w35586_
	);
	LUT2 #(
		.INIT('h8)
	) name25075 (
		\wishbone_RxDataLatched2_reg[7]/NET0131 ,
		_w35519_,
		_w35587_
	);
	LUT2 #(
		.INIT('h1)
	) name25076 (
		_w35586_,
		_w35587_,
		_w35588_
	);
	LUT2 #(
		.INIT('h2)
	) name25077 (
		\wishbone_rx_fifo_fifo_reg[9][9]/P0001 ,
		_w35519_,
		_w35589_
	);
	LUT2 #(
		.INIT('h8)
	) name25078 (
		\wishbone_RxDataLatched2_reg[9]/NET0131 ,
		_w35519_,
		_w35590_
	);
	LUT2 #(
		.INIT('h1)
	) name25079 (
		_w35589_,
		_w35590_,
		_w35591_
	);
	LUT2 #(
		.INIT('h8)
	) name25080 (
		\wishbone_tx_fifo_cnt_reg[0]/NET0131 ,
		_w33028_,
		_w35592_
	);
	LUT2 #(
		.INIT('h8)
	) name25081 (
		_w34093_,
		_w35592_,
		_w35593_
	);
	LUT2 #(
		.INIT('h1)
	) name25082 (
		_w34093_,
		_w35592_,
		_w35594_
	);
	LUT2 #(
		.INIT('h1)
	) name25083 (
		_w35593_,
		_w35594_,
		_w35595_
	);
	LUT2 #(
		.INIT('h8)
	) name25084 (
		_w35444_,
		_w35516_,
		_w35596_
	);
	LUT2 #(
		.INIT('h1)
	) name25085 (
		_w31950_,
		_w35596_,
		_w35597_
	);
	LUT2 #(
		.INIT('h2)
	) name25086 (
		_w34136_,
		_w35597_,
		_w35598_
	);
	LUT2 #(
		.INIT('h8)
	) name25087 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35599_
	);
	LUT2 #(
		.INIT('h8)
	) name25088 (
		_w35247_,
		_w35599_,
		_w35600_
	);
	LUT2 #(
		.INIT('h8)
	) name25089 (
		_w35292_,
		_w35599_,
		_w35601_
	);
	LUT2 #(
		.INIT('h8)
	) name25090 (
		_w35244_,
		_w35445_,
		_w35602_
	);
	LUT2 #(
		.INIT('h8)
	) name25091 (
		_w35445_,
		_w35599_,
		_w35603_
	);
	LUT2 #(
		.INIT('h4)
	) name25092 (
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35236_,
		_w35604_
	);
	LUT2 #(
		.INIT('h8)
	) name25093 (
		_w35517_,
		_w35604_,
		_w35605_
	);
	LUT2 #(
		.INIT('h8)
	) name25094 (
		_w35247_,
		_w35444_,
		_w35606_
	);
	LUT2 #(
		.INIT('h8)
	) name25095 (
		_w35292_,
		_w35444_,
		_w35607_
	);
	LUT2 #(
		.INIT('h8)
	) name25096 (
		_w35342_,
		_w35445_,
		_w35608_
	);
	LUT2 #(
		.INIT('h8)
	) name25097 (
		_w35244_,
		_w35516_,
		_w35609_
	);
	LUT2 #(
		.INIT('h8)
	) name25098 (
		_w35245_,
		_w35609_,
		_w35610_
	);
	LUT2 #(
		.INIT('h8)
	) name25099 (
		\miim1_LatchByte_reg[0]/NET0131 ,
		_w31426_,
		_w35611_
	);
	LUT2 #(
		.INIT('h8)
	) name25100 (
		_w31401_,
		_w35611_,
		_w35612_
	);
	LUT2 #(
		.INIT('h8)
	) name25101 (
		\wishbone_tx_fifo_read_pointer_reg[0]/NET0131 ,
		_w33028_,
		_w35613_
	);
	LUT2 #(
		.INIT('h4)
	) name25102 (
		_w34090_,
		_w35613_,
		_w35614_
	);
	LUT2 #(
		.INIT('h2)
	) name25103 (
		_w34090_,
		_w35613_,
		_w35615_
	);
	LUT2 #(
		.INIT('h1)
	) name25104 (
		_w35614_,
		_w35615_,
		_w35616_
	);
	LUT2 #(
		.INIT('h8)
	) name25105 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[7]/NET0131 ,
		_w34941_,
		_w35617_
	);
	LUT2 #(
		.INIT('h8)
	) name25106 (
		\ethreg1_TXCTRL_1_DataOut_reg[7]/NET0131 ,
		_w34263_,
		_w35618_
	);
	LUT2 #(
		.INIT('h1)
	) name25107 (
		_w34960_,
		_w35617_,
		_w35619_
	);
	LUT2 #(
		.INIT('h4)
	) name25108 (
		_w35618_,
		_w35619_,
		_w35620_
	);
	LUT2 #(
		.INIT('h2)
	) name25109 (
		_w34947_,
		_w35620_,
		_w35621_
	);
	LUT2 #(
		.INIT('h8)
	) name25110 (
		_w34935_,
		_w34957_,
		_w35622_
	);
	LUT2 #(
		.INIT('h8)
	) name25111 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[7]/NET0131 ,
		_w35622_,
		_w35623_
	);
	LUT2 #(
		.INIT('h8)
	) name25112 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[7]/NET0131 ,
		_w34955_,
		_w35624_
	);
	LUT2 #(
		.INIT('h8)
	) name25113 (
		_w34265_,
		_w34941_,
		_w35625_
	);
	LUT2 #(
		.INIT('h8)
	) name25114 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[7]/NET0131 ,
		_w35625_,
		_w35626_
	);
	LUT2 #(
		.INIT('h8)
	) name25115 (
		_w34941_,
		_w34957_,
		_w35627_
	);
	LUT2 #(
		.INIT('h8)
	) name25116 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[7]/NET0131 ,
		_w35627_,
		_w35628_
	);
	LUT2 #(
		.INIT('h8)
	) name25117 (
		\ethreg1_TXCTRL_0_DataOut_reg[7]/NET0131 ,
		_w34266_,
		_w35629_
	);
	LUT2 #(
		.INIT('h8)
	) name25118 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[7]/NET0131 ,
		_w34938_,
		_w35630_
	);
	LUT2 #(
		.INIT('h1)
	) name25119 (
		_w34265_,
		_w34937_,
		_w35631_
	);
	LUT2 #(
		.INIT('h2)
	) name25120 (
		_w34949_,
		_w35631_,
		_w35632_
	);
	LUT2 #(
		.INIT('h1)
	) name25121 (
		_w35623_,
		_w35624_,
		_w35633_
	);
	LUT2 #(
		.INIT('h1)
	) name25122 (
		_w35626_,
		_w35628_,
		_w35634_
	);
	LUT2 #(
		.INIT('h1)
	) name25123 (
		_w35629_,
		_w35630_,
		_w35635_
	);
	LUT2 #(
		.INIT('h4)
	) name25124 (
		_w35632_,
		_w35635_,
		_w35636_
	);
	LUT2 #(
		.INIT('h8)
	) name25125 (
		_w35633_,
		_w35634_,
		_w35637_
	);
	LUT2 #(
		.INIT('h8)
	) name25126 (
		_w35636_,
		_w35637_,
		_w35638_
	);
	LUT2 #(
		.INIT('h4)
	) name25127 (
		_w35621_,
		_w35638_,
		_w35639_
	);
	LUT2 #(
		.INIT('h4)
	) name25128 (
		_w12554_,
		_w15698_,
		_w35640_
	);
	LUT2 #(
		.INIT('h8)
	) name25129 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		_w35640_,
		_w35641_
	);
	LUT2 #(
		.INIT('h8)
	) name25130 (
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w35641_,
		_w35642_
	);
	LUT2 #(
		.INIT('h8)
	) name25131 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		_w35642_,
		_w35643_
	);
	LUT2 #(
		.INIT('h2)
	) name25132 (
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w35643_,
		_w35644_
	);
	LUT2 #(
		.INIT('h4)
	) name25133 (
		\wishbone_rx_fifo_read_pointer_reg[3]/NET0131 ,
		_w35643_,
		_w35645_
	);
	LUT2 #(
		.INIT('h1)
	) name25134 (
		_w35644_,
		_w35645_,
		_w35646_
	);
	LUT2 #(
		.INIT('h1)
	) name25135 (
		_w31950_,
		_w35646_,
		_w35647_
	);
	LUT2 #(
		.INIT('h1)
	) name25136 (
		_w34082_,
		_w34092_,
		_w35648_
	);
	LUT2 #(
		.INIT('h1)
	) name25137 (
		_w34086_,
		_w34091_,
		_w35649_
	);
	LUT2 #(
		.INIT('h1)
	) name25138 (
		_w35648_,
		_w35649_,
		_w35650_
	);
	LUT2 #(
		.INIT('h8)
	) name25139 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w35650_,
		_w35651_
	);
	LUT2 #(
		.INIT('h1)
	) name25140 (
		\wishbone_tx_fifo_cnt_reg[2]/NET0131 ,
		_w35650_,
		_w35652_
	);
	LUT2 #(
		.INIT('h2)
	) name25141 (
		_w33028_,
		_w35651_,
		_w35653_
	);
	LUT2 #(
		.INIT('h4)
	) name25142 (
		_w35652_,
		_w35653_,
		_w35654_
	);
	LUT2 #(
		.INIT('h1)
	) name25143 (
		_w33039_,
		_w33049_,
		_w35655_
	);
	LUT2 #(
		.INIT('h8)
	) name25144 (
		_w34090_,
		_w35655_,
		_w35656_
	);
	LUT2 #(
		.INIT('h1)
	) name25145 (
		\wishbone_tx_fifo_read_pointer_reg[1]/NET0131 ,
		_w34090_,
		_w35657_
	);
	LUT2 #(
		.INIT('h2)
	) name25146 (
		_w33028_,
		_w35656_,
		_w35658_
	);
	LUT2 #(
		.INIT('h4)
	) name25147 (
		_w35657_,
		_w35658_,
		_w35659_
	);
	LUT2 #(
		.INIT('h8)
	) name25148 (
		_w33045_,
		_w34090_,
		_w35660_
	);
	LUT2 #(
		.INIT('h8)
	) name25149 (
		_w33034_,
		_w34090_,
		_w35661_
	);
	LUT2 #(
		.INIT('h8)
	) name25150 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		_w35661_,
		_w35662_
	);
	LUT2 #(
		.INIT('h1)
	) name25151 (
		\wishbone_tx_fifo_read_pointer_reg[3]/NET0131 ,
		_w35662_,
		_w35663_
	);
	LUT2 #(
		.INIT('h2)
	) name25152 (
		_w33028_,
		_w35660_,
		_w35664_
	);
	LUT2 #(
		.INIT('h4)
	) name25153 (
		_w35663_,
		_w35664_,
		_w35665_
	);
	LUT2 #(
		.INIT('h8)
	) name25154 (
		\wishbone_rx_fifo_write_pointer_reg[0]/NET0131 ,
		_w34136_,
		_w35666_
	);
	LUT2 #(
		.INIT('h8)
	) name25155 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w35666_,
		_w35667_
	);
	LUT2 #(
		.INIT('h1)
	) name25156 (
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w35667_,
		_w35668_
	);
	LUT2 #(
		.INIT('h8)
	) name25157 (
		\wishbone_rx_fifo_write_pointer_reg[2]/NET0131 ,
		_w35667_,
		_w35669_
	);
	LUT2 #(
		.INIT('h1)
	) name25158 (
		_w31950_,
		_w35668_,
		_w35670_
	);
	LUT2 #(
		.INIT('h4)
	) name25159 (
		_w35669_,
		_w35670_,
		_w35671_
	);
	LUT2 #(
		.INIT('h1)
	) name25160 (
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35669_,
		_w35672_
	);
	LUT2 #(
		.INIT('h8)
	) name25161 (
		\wishbone_rx_fifo_write_pointer_reg[3]/NET0131 ,
		_w35669_,
		_w35673_
	);
	LUT2 #(
		.INIT('h1)
	) name25162 (
		_w31950_,
		_w35672_,
		_w35674_
	);
	LUT2 #(
		.INIT('h4)
	) name25163 (
		_w35673_,
		_w35674_,
		_w35675_
	);
	LUT2 #(
		.INIT('h1)
	) name25164 (
		\wishbone_tx_fifo_write_pointer_reg[2]/NET0131 ,
		_w34473_,
		_w35676_
	);
	LUT2 #(
		.INIT('h2)
	) name25165 (
		_w33028_,
		_w34474_,
		_w35677_
	);
	LUT2 #(
		.INIT('h4)
	) name25166 (
		_w35676_,
		_w35677_,
		_w35678_
	);
	LUT2 #(
		.INIT('h2)
	) name25167 (
		\wishbone_tx_fifo_write_pointer_reg[3]/NET0131 ,
		_w34474_,
		_w35679_
	);
	LUT2 #(
		.INIT('h1)
	) name25168 (
		_w34475_,
		_w35679_,
		_w35680_
	);
	LUT2 #(
		.INIT('h2)
	) name25169 (
		_w33028_,
		_w35680_,
		_w35681_
	);
	LUT2 #(
		.INIT('h8)
	) name25170 (
		\wishbone_TxEn_reg/NET0131 ,
		_w34991_,
		_w35682_
	);
	LUT2 #(
		.INIT('h1)
	) name25171 (
		_w34981_,
		_w35682_,
		_w35683_
	);
	LUT2 #(
		.INIT('h4)
	) name25172 (
		_w10650_,
		_w34563_,
		_w35684_
	);
	LUT2 #(
		.INIT('h2)
	) name25173 (
		_w11758_,
		_w35684_,
		_w35685_
	);
	LUT2 #(
		.INIT('h1)
	) name25174 (
		\wishbone_rx_fifo_write_pointer_reg[1]/NET0131 ,
		_w35666_,
		_w35686_
	);
	LUT2 #(
		.INIT('h1)
	) name25175 (
		_w31950_,
		_w35667_,
		_w35687_
	);
	LUT2 #(
		.INIT('h4)
	) name25176 (
		_w35686_,
		_w35687_,
		_w35688_
	);
	LUT2 #(
		.INIT('h8)
	) name25177 (
		\wishbone_tx_fifo_cnt_reg[1]/NET0131 ,
		_w34093_,
		_w35689_
	);
	LUT2 #(
		.INIT('h1)
	) name25178 (
		_w34082_,
		_w34086_,
		_w35690_
	);
	LUT2 #(
		.INIT('h2)
	) name25179 (
		_w34092_,
		_w35690_,
		_w35691_
	);
	LUT2 #(
		.INIT('h8)
	) name25180 (
		_w34091_,
		_w35690_,
		_w35692_
	);
	LUT2 #(
		.INIT('h1)
	) name25181 (
		_w35691_,
		_w35692_,
		_w35693_
	);
	LUT2 #(
		.INIT('h4)
	) name25182 (
		_w35689_,
		_w35693_,
		_w35694_
	);
	LUT2 #(
		.INIT('h2)
	) name25183 (
		_w33028_,
		_w35694_,
		_w35695_
	);
	LUT2 #(
		.INIT('h1)
	) name25184 (
		\wishbone_tx_fifo_read_pointer_reg[2]/NET0131 ,
		_w35661_,
		_w35696_
	);
	LUT2 #(
		.INIT('h2)
	) name25185 (
		_w33028_,
		_w35662_,
		_w35697_
	);
	LUT2 #(
		.INIT('h4)
	) name25186 (
		_w35696_,
		_w35697_,
		_w35698_
	);
	LUT2 #(
		.INIT('h1)
	) name25187 (
		\wishbone_tx_fifo_write_pointer_reg[1]/NET0131 ,
		_w34458_,
		_w35699_
	);
	LUT2 #(
		.INIT('h2)
	) name25188 (
		_w33028_,
		_w34473_,
		_w35700_
	);
	LUT2 #(
		.INIT('h4)
	) name25189 (
		_w35699_,
		_w35700_,
		_w35701_
	);
	LUT2 #(
		.INIT('h2)
	) name25190 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_PauseTimerEq0_sync2_reg/NET0131 ,
		_w35702_
	);
	LUT2 #(
		.INIT('h2)
	) name25191 (
		_w11181_,
		_w11414_,
		_w35703_
	);
	LUT2 #(
		.INIT('h8)
	) name25192 (
		\wb_sel_i[2]_pad ,
		_w22942_,
		_w35704_
	);
	LUT2 #(
		.INIT('h8)
	) name25193 (
		_w31683_,
		_w35704_,
		_w35705_
	);
	LUT2 #(
		.INIT('h8)
	) name25194 (
		_w23499_,
		_w35705_,
		_w35706_
	);
	LUT2 #(
		.INIT('h4)
	) name25195 (
		\wb_dat_i[16]_pad ,
		_w35706_,
		_w35707_
	);
	LUT2 #(
		.INIT('h1)
	) name25196 (
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		_w35706_,
		_w35708_
	);
	LUT2 #(
		.INIT('h1)
	) name25197 (
		\RstTxPauseRq_reg/NET0131 ,
		_w35707_,
		_w35709_
	);
	LUT2 #(
		.INIT('h4)
	) name25198 (
		_w35708_,
		_w35709_,
		_w35710_
	);
	LUT2 #(
		.INIT('h1)
	) name25199 (
		\RxAbort_wb_reg/NET0131 ,
		\rxethmac1_RxEndFrm_reg/NET0131 ,
		_w35711_
	);
	LUT2 #(
		.INIT('h8)
	) name25200 (
		\wishbone_RxEnableWindow_reg/NET0131 ,
		_w35711_,
		_w35712_
	);
	LUT2 #(
		.INIT('h1)
	) name25201 (
		\rxethmac1_RxStartFrm_reg/NET0131 ,
		_w35712_,
		_w35713_
	);
	LUT2 #(
		.INIT('h8)
	) name25202 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		\miim1_clkgen_Counter_reg[1]/NET0131 ,
		_w35714_
	);
	LUT2 #(
		.INIT('h1)
	) name25203 (
		_w31190_,
		_w35714_,
		_w35715_
	);
	LUT2 #(
		.INIT('h4)
	) name25204 (
		_w31208_,
		_w35715_,
		_w35716_
	);
	LUT2 #(
		.INIT('h8)
	) name25205 (
		\ethreg1_MIIMODER_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_MIIMODER_0_DataOut_reg[2]/NET0131 ,
		_w35717_
	);
	LUT2 #(
		.INIT('h1)
	) name25206 (
		_w31202_,
		_w35717_,
		_w35718_
	);
	LUT2 #(
		.INIT('h8)
	) name25207 (
		_w31208_,
		_w35718_,
		_w35719_
	);
	LUT2 #(
		.INIT('h1)
	) name25208 (
		_w35716_,
		_w35719_,
		_w35720_
	);
	LUT2 #(
		.INIT('h2)
	) name25209 (
		\rxethmac1_rxaddrcheck1_AddressMiss_reg/NET0131 ,
		_w12512_,
		_w35721_
	);
	LUT2 #(
		.INIT('h4)
	) name25210 (
		\ethreg1_MODER_0_DataOut_reg[3]/NET0131 ,
		\rxethmac1_Broadcast_reg/NET0131 ,
		_w35722_
	);
	LUT2 #(
		.INIT('h1)
	) name25211 (
		\rxethmac1_rxaddrcheck1_MulticastOK_reg/NET0131 ,
		\rxethmac1_rxaddrcheck1_UnicastOK_reg/NET0131 ,
		_w35723_
	);
	LUT2 #(
		.INIT('h4)
	) name25212 (
		_w35722_,
		_w35723_,
		_w35724_
	);
	LUT2 #(
		.INIT('h8)
	) name25213 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\maccontrol1_receivecontrol1_AddressOK_reg/NET0131 ,
		_w35725_
	);
	LUT2 #(
		.INIT('h2)
	) name25214 (
		_w35724_,
		_w35725_,
		_w35726_
	);
	LUT2 #(
		.INIT('h8)
	) name25215 (
		_w12512_,
		_w35726_,
		_w35727_
	);
	LUT2 #(
		.INIT('h1)
	) name25216 (
		_w35721_,
		_w35727_,
		_w35728_
	);
	LUT2 #(
		.INIT('h8)
	) name25217 (
		\wb_dat_i[11]_pad ,
		_w34989_,
		_w35729_
	);
	LUT2 #(
		.INIT('h8)
	) name25218 (
		\wishbone_TxStatus_reg[11]/NET0131 ,
		_w34981_,
		_w35730_
	);
	LUT2 #(
		.INIT('h8)
	) name25219 (
		\wishbone_ram_di_reg[11]/NET0131 ,
		_w34991_,
		_w35731_
	);
	LUT2 #(
		.INIT('h1)
	) name25220 (
		_w35729_,
		_w35730_,
		_w35732_
	);
	LUT2 #(
		.INIT('h4)
	) name25221 (
		_w35731_,
		_w35732_,
		_w35733_
	);
	LUT2 #(
		.INIT('h8)
	) name25222 (
		\wb_dat_i[12]_pad ,
		_w34989_,
		_w35734_
	);
	LUT2 #(
		.INIT('h8)
	) name25223 (
		\wishbone_TxStatus_reg[12]/NET0131 ,
		_w34981_,
		_w35735_
	);
	LUT2 #(
		.INIT('h8)
	) name25224 (
		\wishbone_ram_di_reg[12]/NET0131 ,
		_w34991_,
		_w35736_
	);
	LUT2 #(
		.INIT('h1)
	) name25225 (
		_w35734_,
		_w35735_,
		_w35737_
	);
	LUT2 #(
		.INIT('h4)
	) name25226 (
		_w35736_,
		_w35737_,
		_w35738_
	);
	LUT2 #(
		.INIT('h2)
	) name25227 (
		\txethmac1_random1_RandomLatched_reg[8]/NET0131 ,
		_w34968_,
		_w35739_
	);
	LUT2 #(
		.INIT('h1)
	) name25228 (
		\txethmac1_RetryCnt_reg[0]/NET0131 ,
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w35740_
	);
	LUT2 #(
		.INIT('h4)
	) name25229 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w35740_,
		_w35741_
	);
	LUT2 #(
		.INIT('h8)
	) name25230 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[8]/NET0131 ,
		_w35742_
	);
	LUT2 #(
		.INIT('h8)
	) name25231 (
		_w34968_,
		_w35742_,
		_w35743_
	);
	LUT2 #(
		.INIT('h4)
	) name25232 (
		_w35741_,
		_w35743_,
		_w35744_
	);
	LUT2 #(
		.INIT('h1)
	) name25233 (
		_w35739_,
		_w35744_,
		_w35745_
	);
	LUT2 #(
		.INIT('h2)
	) name25234 (
		\wishbone_BDRead_reg/NET0131 ,
		_w34989_,
		_w35746_
	);
	LUT2 #(
		.INIT('h2)
	) name25235 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w35747_
	);
	LUT2 #(
		.INIT('h8)
	) name25236 (
		_w22942_,
		_w35747_,
		_w35748_
	);
	LUT2 #(
		.INIT('h8)
	) name25237 (
		_w34989_,
		_w35748_,
		_w35749_
	);
	LUT2 #(
		.INIT('h1)
	) name25238 (
		_w35746_,
		_w35749_,
		_w35750_
	);
	LUT2 #(
		.INIT('h2)
	) name25239 (
		\wishbone_TxAbort_wb_q_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w35751_
	);
	LUT2 #(
		.INIT('h1)
	) name25240 (
		\wishbone_TxAbortPacketBlocked_reg/NET0131 ,
		\wishbone_TxAbortPacket_reg/NET0131 ,
		_w35752_
	);
	LUT2 #(
		.INIT('h1)
	) name25241 (
		_w35751_,
		_w35752_,
		_w35753_
	);
	LUT2 #(
		.INIT('h2)
	) name25242 (
		\wishbone_TxDone_wb_q_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w35754_
	);
	LUT2 #(
		.INIT('h1)
	) name25243 (
		\wishbone_TxDonePacketBlocked_reg/NET0131 ,
		\wishbone_TxDonePacket_reg/NET0131 ,
		_w35755_
	);
	LUT2 #(
		.INIT('h1)
	) name25244 (
		_w35754_,
		_w35755_,
		_w35756_
	);
	LUT2 #(
		.INIT('h1)
	) name25245 (
		\txethmac1_random1_x_reg[2]/NET0131 ,
		\txethmac1_random1_x_reg[9]/NET0131 ,
		_w35757_
	);
	LUT2 #(
		.INIT('h8)
	) name25246 (
		\txethmac1_random1_x_reg[2]/NET0131 ,
		\txethmac1_random1_x_reg[9]/NET0131 ,
		_w35758_
	);
	LUT2 #(
		.INIT('h1)
	) name25247 (
		_w35757_,
		_w35758_,
		_w35759_
	);
	LUT2 #(
		.INIT('h2)
	) name25248 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11481_,
		_w35760_
	);
	LUT2 #(
		.INIT('h1)
	) name25249 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[11]/NET0131 ,
		_w35761_
	);
	LUT2 #(
		.INIT('h1)
	) name25250 (
		_w35760_,
		_w35761_,
		_w35762_
	);
	LUT2 #(
		.INIT('h8)
	) name25251 (
		\TPauseRq_reg/NET0131 ,
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		_w35763_
	);
	LUT2 #(
		.INIT('h1)
	) name25252 (
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		_w35763_,
		_w35764_
	);
	LUT2 #(
		.INIT('h1)
	) name25253 (
		_w10682_,
		_w35764_,
		_w35765_
	);
	LUT2 #(
		.INIT('h1)
	) name25254 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[4]/NET0131 ,
		_w11623_,
		_w35766_
	);
	LUT2 #(
		.INIT('h1)
	) name25255 (
		wb_rst_i_pad,
		_w11624_,
		_w35767_
	);
	LUT2 #(
		.INIT('h4)
	) name25256 (
		_w35766_,
		_w35767_,
		_w35768_
	);
	LUT2 #(
		.INIT('h8)
	) name25257 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		_w34892_,
		_w35769_
	);
	LUT2 #(
		.INIT('h1)
	) name25258 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		_w34895_,
		_w35770_
	);
	LUT2 #(
		.INIT('h1)
	) name25259 (
		_w34889_,
		_w35769_,
		_w35771_
	);
	LUT2 #(
		.INIT('h4)
	) name25260 (
		_w35770_,
		_w35771_,
		_w35772_
	);
	LUT2 #(
		.INIT('h2)
	) name25261 (
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w34892_,
		_w35773_
	);
	LUT2 #(
		.INIT('h1)
	) name25262 (
		\wishbone_TxBDAddress_reg[1]/NET0131 ,
		\wishbone_TxBDAddress_reg[2]/NET0131 ,
		_w35774_
	);
	LUT2 #(
		.INIT('h1)
	) name25263 (
		_w34897_,
		_w35774_,
		_w35775_
	);
	LUT2 #(
		.INIT('h8)
	) name25264 (
		_w34895_,
		_w35775_,
		_w35776_
	);
	LUT2 #(
		.INIT('h1)
	) name25265 (
		_w35773_,
		_w35776_,
		_w35777_
	);
	LUT2 #(
		.INIT('h1)
	) name25266 (
		_w34889_,
		_w35777_,
		_w35778_
	);
	LUT2 #(
		.INIT('h2)
	) name25267 (
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w34892_,
		_w35779_
	);
	LUT2 #(
		.INIT('h1)
	) name25268 (
		\wishbone_TxBDAddress_reg[3]/NET0131 ,
		_w34897_,
		_w35780_
	);
	LUT2 #(
		.INIT('h1)
	) name25269 (
		_w34898_,
		_w35780_,
		_w35781_
	);
	LUT2 #(
		.INIT('h8)
	) name25270 (
		_w34895_,
		_w35781_,
		_w35782_
	);
	LUT2 #(
		.INIT('h1)
	) name25271 (
		_w35779_,
		_w35782_,
		_w35783_
	);
	LUT2 #(
		.INIT('h1)
	) name25272 (
		_w34889_,
		_w35783_,
		_w35784_
	);
	LUT2 #(
		.INIT('h2)
	) name25273 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w34892_,
		_w35785_
	);
	LUT2 #(
		.INIT('h1)
	) name25274 (
		\wishbone_TxBDAddress_reg[5]/NET0131 ,
		_w34900_,
		_w35786_
	);
	LUT2 #(
		.INIT('h2)
	) name25275 (
		_w34895_,
		_w34904_,
		_w35787_
	);
	LUT2 #(
		.INIT('h4)
	) name25276 (
		_w35786_,
		_w35787_,
		_w35788_
	);
	LUT2 #(
		.INIT('h1)
	) name25277 (
		_w35785_,
		_w35788_,
		_w35789_
	);
	LUT2 #(
		.INIT('h1)
	) name25278 (
		_w34889_,
		_w35789_,
		_w35790_
	);
	LUT2 #(
		.INIT('h2)
	) name25279 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w12240_,
		_w35791_
	);
	LUT2 #(
		.INIT('h8)
	) name25280 (
		\wishbone_TxPointerLSB_reg[0]/NET0131 ,
		_w35791_,
		_w35792_
	);
	LUT2 #(
		.INIT('h1)
	) name25281 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		_w12246_,
		_w35793_
	);
	LUT2 #(
		.INIT('h8)
	) name25282 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		_w12246_,
		_w35794_
	);
	LUT2 #(
		.INIT('h1)
	) name25283 (
		_w35793_,
		_w35794_,
		_w35795_
	);
	LUT2 #(
		.INIT('h1)
	) name25284 (
		_w35791_,
		_w35795_,
		_w35796_
	);
	LUT2 #(
		.INIT('h1)
	) name25285 (
		\wishbone_TxAbort_q_reg/NET0131 ,
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w35797_
	);
	LUT2 #(
		.INIT('h4)
	) name25286 (
		_w35792_,
		_w35797_,
		_w35798_
	);
	LUT2 #(
		.INIT('h4)
	) name25287 (
		_w35796_,
		_w35798_,
		_w35799_
	);
	LUT2 #(
		.INIT('h1)
	) name25288 (
		_w12267_,
		_w12269_,
		_w35800_
	);
	LUT2 #(
		.INIT('h2)
	) name25289 (
		_w35791_,
		_w35800_,
		_w35801_
	);
	LUT2 #(
		.INIT('h1)
	) name25290 (
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w35794_,
		_w35802_
	);
	LUT2 #(
		.INIT('h8)
	) name25291 (
		\wishbone_TxByteCnt_reg[1]/NET0131 ,
		_w35794_,
		_w35803_
	);
	LUT2 #(
		.INIT('h1)
	) name25292 (
		_w35791_,
		_w35802_,
		_w35804_
	);
	LUT2 #(
		.INIT('h4)
	) name25293 (
		_w35803_,
		_w35804_,
		_w35805_
	);
	LUT2 #(
		.INIT('h1)
	) name25294 (
		_w35801_,
		_w35805_,
		_w35806_
	);
	LUT2 #(
		.INIT('h2)
	) name25295 (
		_w35797_,
		_w35806_,
		_w35807_
	);
	LUT2 #(
		.INIT('h4)
	) name25296 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w34977_,
		_w35808_
	);
	LUT2 #(
		.INIT('h2)
	) name25297 (
		\wishbone_WbEn_reg/NET0131 ,
		_w35808_,
		_w35809_
	);
	LUT2 #(
		.INIT('h8)
	) name25298 (
		_w34991_,
		_w35809_,
		_w35810_
	);
	LUT2 #(
		.INIT('h1)
	) name25299 (
		_w34989_,
		_w35810_,
		_w35811_
	);
	LUT2 #(
		.INIT('h4)
	) name25300 (
		\miim1_BitCounter_reg[5]/NET0131 ,
		_w31411_,
		_w35812_
	);
	LUT2 #(
		.INIT('h1)
	) name25301 (
		_w34930_,
		_w35812_,
		_w35813_
	);
	LUT2 #(
		.INIT('h1)
	) name25302 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[2]/NET0131 ,
		_w34863_,
		_w35814_
	);
	LUT2 #(
		.INIT('h2)
	) name25303 (
		_w34861_,
		_w34864_,
		_w35815_
	);
	LUT2 #(
		.INIT('h4)
	) name25304 (
		_w35814_,
		_w35815_,
		_w35816_
	);
	LUT2 #(
		.INIT('h1)
	) name25305 (
		\wishbone_WB_ACK_O_reg/P0001 ,
		_w22943_,
		_w35817_
	);
	LUT2 #(
		.INIT('h1)
	) name25306 (
		wb_ack_o_pad,
		_w35817_,
		_w35818_
	);
	LUT2 #(
		.INIT('h1)
	) name25307 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[2]/NET0131 ,
		_w11621_,
		_w35819_
	);
	LUT2 #(
		.INIT('h1)
	) name25308 (
		wb_rst_i_pad,
		_w11622_,
		_w35820_
	);
	LUT2 #(
		.INIT('h4)
	) name25309 (
		_w35819_,
		_w35820_,
		_w35821_
	);
	LUT2 #(
		.INIT('h8)
	) name25310 (
		_w23498_,
		_w34566_,
		_w35822_
	);
	LUT2 #(
		.INIT('h8)
	) name25311 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[3]/NET0131 ,
		_w34938_,
		_w35823_
	);
	LUT2 #(
		.INIT('h8)
	) name25312 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[3]/NET0131 ,
		_w35627_,
		_w35824_
	);
	LUT2 #(
		.INIT('h8)
	) name25313 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[3]/NET0131 ,
		_w34955_,
		_w35825_
	);
	LUT2 #(
		.INIT('h8)
	) name25314 (
		\ethreg1_TXCTRL_0_DataOut_reg[3]/NET0131 ,
		_w34266_,
		_w35826_
	);
	LUT2 #(
		.INIT('h8)
	) name25315 (
		_w34941_,
		_w34947_,
		_w35827_
	);
	LUT2 #(
		.INIT('h8)
	) name25316 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[3]/NET0131 ,
		_w35827_,
		_w35828_
	);
	LUT2 #(
		.INIT('h8)
	) name25317 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[3]/NET0131 ,
		_w35622_,
		_w35829_
	);
	LUT2 #(
		.INIT('h8)
	) name25318 (
		_w34263_,
		_w34947_,
		_w35830_
	);
	LUT2 #(
		.INIT('h8)
	) name25319 (
		\ethreg1_TXCTRL_1_DataOut_reg[3]/NET0131 ,
		_w35830_,
		_w35831_
	);
	LUT2 #(
		.INIT('h8)
	) name25320 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[3]/NET0131 ,
		_w35625_,
		_w35832_
	);
	LUT2 #(
		.INIT('h1)
	) name25321 (
		\maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ,
		\maccontrol1_transmitcontrol1_ByteCnt_reg[2]/NET0131 ,
		_w35833_
	);
	LUT2 #(
		.INIT('h8)
	) name25322 (
		_w34960_,
		_w35833_,
		_w35834_
	);
	LUT2 #(
		.INIT('h1)
	) name25323 (
		_w35823_,
		_w35834_,
		_w35835_
	);
	LUT2 #(
		.INIT('h1)
	) name25324 (
		_w35824_,
		_w35825_,
		_w35836_
	);
	LUT2 #(
		.INIT('h1)
	) name25325 (
		_w35826_,
		_w35828_,
		_w35837_
	);
	LUT2 #(
		.INIT('h1)
	) name25326 (
		_w35829_,
		_w35831_,
		_w35838_
	);
	LUT2 #(
		.INIT('h4)
	) name25327 (
		_w35832_,
		_w35838_,
		_w35839_
	);
	LUT2 #(
		.INIT('h8)
	) name25328 (
		_w35836_,
		_w35837_,
		_w35840_
	);
	LUT2 #(
		.INIT('h8)
	) name25329 (
		_w35835_,
		_w35840_,
		_w35841_
	);
	LUT2 #(
		.INIT('h8)
	) name25330 (
		_w35839_,
		_w35841_,
		_w35842_
	);
	LUT2 #(
		.INIT('h1)
	) name25331 (
		\macstatus1_DribbleNibble_reg/NET0131 ,
		_w11757_,
		_w35843_
	);
	LUT2 #(
		.INIT('h1)
	) name25332 (
		\rxethmac1_rxstatem1_StateSFD_reg/NET0131 ,
		_w35843_,
		_w35844_
	);
	LUT2 #(
		.INIT('h1)
	) name25333 (
		\rxethmac1_CrcHash_reg[2]/P0001 ,
		_w10568_,
		_w35845_
	);
	LUT2 #(
		.INIT('h4)
	) name25334 (
		\rxethmac1_crcrx_Crc_reg[28]/NET0131 ,
		_w10568_,
		_w35846_
	);
	LUT2 #(
		.INIT('h2)
	) name25335 (
		_w10563_,
		_w35845_,
		_w35847_
	);
	LUT2 #(
		.INIT('h4)
	) name25336 (
		_w35846_,
		_w35847_,
		_w35848_
	);
	LUT2 #(
		.INIT('h1)
	) name25337 (
		\rxethmac1_CrcHash_reg[3]/P0001 ,
		_w10568_,
		_w35849_
	);
	LUT2 #(
		.INIT('h4)
	) name25338 (
		\rxethmac1_crcrx_Crc_reg[29]/NET0131 ,
		_w10568_,
		_w35850_
	);
	LUT2 #(
		.INIT('h2)
	) name25339 (
		_w10563_,
		_w35849_,
		_w35851_
	);
	LUT2 #(
		.INIT('h4)
	) name25340 (
		_w35850_,
		_w35851_,
		_w35852_
	);
	LUT2 #(
		.INIT('h1)
	) name25341 (
		\rxethmac1_CrcHash_reg[4]/P0001 ,
		_w10568_,
		_w35853_
	);
	LUT2 #(
		.INIT('h4)
	) name25342 (
		\rxethmac1_crcrx_Crc_reg[30]/NET0131 ,
		_w10568_,
		_w35854_
	);
	LUT2 #(
		.INIT('h2)
	) name25343 (
		_w10563_,
		_w35853_,
		_w35855_
	);
	LUT2 #(
		.INIT('h4)
	) name25344 (
		_w35854_,
		_w35855_,
		_w35856_
	);
	LUT2 #(
		.INIT('h1)
	) name25345 (
		\rxethmac1_CrcHash_reg[5]/P0001 ,
		_w10568_,
		_w35857_
	);
	LUT2 #(
		.INIT('h4)
	) name25346 (
		\rxethmac1_crcrx_Crc_reg[31]/NET0131 ,
		_w10568_,
		_w35858_
	);
	LUT2 #(
		.INIT('h2)
	) name25347 (
		_w10563_,
		_w35857_,
		_w35859_
	);
	LUT2 #(
		.INIT('h4)
	) name25348 (
		_w35858_,
		_w35859_,
		_w35860_
	);
	LUT2 #(
		.INIT('h1)
	) name25349 (
		\wishbone_ReadTxDataFromMemory_reg/NET0131 ,
		_w17883_,
		_w35861_
	);
	LUT2 #(
		.INIT('h2)
	) name25350 (
		_w34289_,
		_w35861_,
		_w35862_
	);
	LUT2 #(
		.INIT('h4)
	) name25351 (
		_w34916_,
		_w35862_,
		_w35863_
	);
	LUT2 #(
		.INIT('h8)
	) name25352 (
		\wishbone_RxEn_reg/NET0131 ,
		_w34990_,
		_w35864_
	);
	LUT2 #(
		.INIT('h1)
	) name25353 (
		_w34984_,
		_w35864_,
		_w35865_
	);
	LUT2 #(
		.INIT('h2)
	) name25354 (
		mdc_pad_o_pad,
		_w31208_,
		_w35866_
	);
	LUT2 #(
		.INIT('h1)
	) name25355 (
		_w34106_,
		_w35866_,
		_w35867_
	);
	LUT2 #(
		.INIT('h8)
	) name25356 (
		\rxethmac1_LatchedByte_reg[1]/NET0131 ,
		_w31852_,
		_w35868_
	);
	LUT2 #(
		.INIT('h8)
	) name25357 (
		\rxethmac1_RxData_d_reg[1]/NET0131 ,
		_w31853_,
		_w35869_
	);
	LUT2 #(
		.INIT('h1)
	) name25358 (
		_w35868_,
		_w35869_,
		_w35870_
	);
	LUT2 #(
		.INIT('h8)
	) name25359 (
		\rxethmac1_LatchedByte_reg[2]/NET0131 ,
		_w31852_,
		_w35871_
	);
	LUT2 #(
		.INIT('h8)
	) name25360 (
		\rxethmac1_RxData_d_reg[2]/NET0131 ,
		_w31853_,
		_w35872_
	);
	LUT2 #(
		.INIT('h1)
	) name25361 (
		_w35871_,
		_w35872_,
		_w35873_
	);
	LUT2 #(
		.INIT('h8)
	) name25362 (
		\rxethmac1_LatchedByte_reg[3]/NET0131 ,
		_w31852_,
		_w35874_
	);
	LUT2 #(
		.INIT('h8)
	) name25363 (
		\rxethmac1_RxData_d_reg[3]/NET0131 ,
		_w31853_,
		_w35875_
	);
	LUT2 #(
		.INIT('h1)
	) name25364 (
		_w35874_,
		_w35875_,
		_w35876_
	);
	LUT2 #(
		.INIT('h8)
	) name25365 (
		\rxethmac1_LatchedByte_reg[5]/NET0131 ,
		_w31852_,
		_w35877_
	);
	LUT2 #(
		.INIT('h8)
	) name25366 (
		\rxethmac1_RxData_d_reg[5]/NET0131 ,
		_w31853_,
		_w35878_
	);
	LUT2 #(
		.INIT('h1)
	) name25367 (
		_w35877_,
		_w35878_,
		_w35879_
	);
	LUT2 #(
		.INIT('h8)
	) name25368 (
		\rxethmac1_LatchedByte_reg[6]/NET0131 ,
		_w31852_,
		_w35880_
	);
	LUT2 #(
		.INIT('h8)
	) name25369 (
		\rxethmac1_RxData_d_reg[6]/NET0131 ,
		_w31853_,
		_w35881_
	);
	LUT2 #(
		.INIT('h1)
	) name25370 (
		_w35880_,
		_w35881_,
		_w35882_
	);
	LUT2 #(
		.INIT('h8)
	) name25371 (
		\rxethmac1_LatchedByte_reg[7]/NET0131 ,
		_w31852_,
		_w35883_
	);
	LUT2 #(
		.INIT('h8)
	) name25372 (
		\rxethmac1_RxData_d_reg[7]/NET0131 ,
		_w31853_,
		_w35884_
	);
	LUT2 #(
		.INIT('h1)
	) name25373 (
		_w35883_,
		_w35884_,
		_w35885_
	);
	LUT2 #(
		.INIT('h1)
	) name25374 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[0]/NET0131 ,
		_w10578_,
		_w35886_
	);
	LUT2 #(
		.INIT('h1)
	) name25375 (
		_w34862_,
		_w35886_,
		_w35887_
	);
	LUT2 #(
		.INIT('h1)
	) name25376 (
		_w34857_,
		_w35887_,
		_w35888_
	);
	LUT2 #(
		.INIT('h1)
	) name25377 (
		_w34860_,
		_w35888_,
		_w35889_
	);
	LUT2 #(
		.INIT('h2)
	) name25378 (
		\wb_adr_i[2]_pad ,
		\wb_adr_i[3]_pad ,
		_w35890_
	);
	LUT2 #(
		.INIT('h8)
	) name25379 (
		_w34526_,
		_w35890_,
		_w35891_
	);
	LUT2 #(
		.INIT('h4)
	) name25380 (
		\wb_adr_i[4]_pad ,
		_w31684_,
		_w35892_
	);
	LUT2 #(
		.INIT('h8)
	) name25381 (
		_w22965_,
		_w35892_,
		_w35893_
	);
	LUT2 #(
		.INIT('h1)
	) name25382 (
		\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w35894_
	);
	LUT2 #(
		.INIT('h1)
	) name25383 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxAbort_reg/NET0131 ,
		_w35895_
	);
	LUT2 #(
		.INIT('h4)
	) name25384 (
		\maccontrol1_MuxedAbort_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w35896_
	);
	LUT2 #(
		.INIT('h2)
	) name25385 (
		_w35894_,
		_w35895_,
		_w35897_
	);
	LUT2 #(
		.INIT('h4)
	) name25386 (
		_w35896_,
		_w35897_,
		_w35898_
	);
	LUT2 #(
		.INIT('h1)
	) name25387 (
		\txethmac1_TxRetry_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w35899_
	);
	LUT2 #(
		.INIT('h4)
	) name25388 (
		_w35898_,
		_w35899_,
		_w35900_
	);
	LUT2 #(
		.INIT('h2)
	) name25389 (
		\wishbone_Flop_reg/NET0131 ,
		_w35900_,
		_w35901_
	);
	LUT2 #(
		.INIT('h1)
	) name25390 (
		\wishbone_LastWord_reg/NET0131 ,
		_w35803_,
		_w35902_
	);
	LUT2 #(
		.INIT('h4)
	) name25391 (
		\wishbone_TxEndFrm_wb_reg/NET0131 ,
		_w35803_,
		_w35903_
	);
	LUT2 #(
		.INIT('h1)
	) name25392 (
		_w35901_,
		_w35902_,
		_w35904_
	);
	LUT2 #(
		.INIT('h4)
	) name25393 (
		_w35903_,
		_w35904_,
		_w35905_
	);
	LUT2 #(
		.INIT('h2)
	) name25394 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		_w34989_,
		_w35906_
	);
	LUT2 #(
		.INIT('h8)
	) name25395 (
		\wb_adr_i[10]_pad ,
		wb_we_i_pad,
		_w35907_
	);
	LUT2 #(
		.INIT('h8)
	) name25396 (
		_w34989_,
		_w35907_,
		_w35908_
	);
	LUT2 #(
		.INIT('h8)
	) name25397 (
		_w31682_,
		_w35908_,
		_w35909_
	);
	LUT2 #(
		.INIT('h1)
	) name25398 (
		_w35906_,
		_w35909_,
		_w35910_
	);
	LUT2 #(
		.INIT('h2)
	) name25399 (
		\wishbone_BDWrite_reg[1]/NET0131 ,
		_w34989_,
		_w35911_
	);
	LUT2 #(
		.INIT('h8)
	) name25400 (
		\wb_sel_i[1]_pad ,
		_w22942_,
		_w35912_
	);
	LUT2 #(
		.INIT('h8)
	) name25401 (
		_w35908_,
		_w35912_,
		_w35913_
	);
	LUT2 #(
		.INIT('h1)
	) name25402 (
		_w35911_,
		_w35913_,
		_w35914_
	);
	LUT2 #(
		.INIT('h2)
	) name25403 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		_w34989_,
		_w35915_
	);
	LUT2 #(
		.INIT('h8)
	) name25404 (
		_w35704_,
		_w35908_,
		_w35916_
	);
	LUT2 #(
		.INIT('h1)
	) name25405 (
		_w35915_,
		_w35916_,
		_w35917_
	);
	LUT2 #(
		.INIT('h4)
	) name25406 (
		\wishbone_LastWord_reg/NET0131 ,
		_w35803_,
		_w35918_
	);
	LUT2 #(
		.INIT('h2)
	) name25407 (
		\wishbone_ReadTxDataFromFifo_syncb2_reg/NET0131 ,
		\wishbone_ReadTxDataFromFifo_syncb3_reg/NET0131 ,
		_w35919_
	);
	LUT2 #(
		.INIT('h2)
	) name25408 (
		\wishbone_ReadTxDataFromFifo_tck_reg/NET0131 ,
		_w35919_,
		_w35920_
	);
	LUT2 #(
		.INIT('h8)
	) name25409 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w12253_,
		_w35921_
	);
	LUT2 #(
		.INIT('h8)
	) name25410 (
		_w12246_,
		_w35921_,
		_w35922_
	);
	LUT2 #(
		.INIT('h1)
	) name25411 (
		_w12245_,
		_w35922_,
		_w35923_
	);
	LUT2 #(
		.INIT('h4)
	) name25412 (
		_w35920_,
		_w35923_,
		_w35924_
	);
	LUT2 #(
		.INIT('h4)
	) name25413 (
		_w35918_,
		_w35924_,
		_w35925_
	);
	LUT2 #(
		.INIT('h4)
	) name25414 (
		_w31201_,
		_w31208_,
		_w35926_
	);
	LUT2 #(
		.INIT('h2)
	) name25415 (
		\miim1_clkgen_Counter_reg[0]/NET0131 ,
		_w31208_,
		_w35927_
	);
	LUT2 #(
		.INIT('h1)
	) name25416 (
		_w35926_,
		_w35927_,
		_w35928_
	);
	LUT2 #(
		.INIT('h2)
	) name25417 (
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		_w12655_,
		_w35929_
	);
	LUT2 #(
		.INIT('h1)
	) name25418 (
		\wishbone_tx_burst_en_reg/NET0131 ,
		_w12540_,
		_w35930_
	);
	LUT2 #(
		.INIT('h2)
	) name25419 (
		\wishbone_MasterWbTX_reg/NET0131 ,
		_w35930_,
		_w35931_
	);
	LUT2 #(
		.INIT('h4)
	) name25420 (
		\wishbone_TxAbortPacketBlocked_reg/NET0131 ,
		\wishbone_TxAbort_wb_reg/NET0131 ,
		_w35932_
	);
	LUT2 #(
		.INIT('h4)
	) name25421 (
		_w35931_,
		_w35932_,
		_w35933_
	);
	LUT2 #(
		.INIT('h4)
	) name25422 (
		\wishbone_TxAbortPacket_NotCleared_reg/NET0131 ,
		_w35933_,
		_w35934_
	);
	LUT2 #(
		.INIT('h1)
	) name25423 (
		_w35929_,
		_w35934_,
		_w35935_
	);
	LUT2 #(
		.INIT('h2)
	) name25424 (
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		_w12655_,
		_w35936_
	);
	LUT2 #(
		.INIT('h4)
	) name25425 (
		\wishbone_TxDonePacketBlocked_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w35937_
	);
	LUT2 #(
		.INIT('h4)
	) name25426 (
		_w35931_,
		_w35937_,
		_w35938_
	);
	LUT2 #(
		.INIT('h4)
	) name25427 (
		\wishbone_TxDonePacket_NotCleared_reg/NET0131 ,
		_w35938_,
		_w35939_
	);
	LUT2 #(
		.INIT('h1)
	) name25428 (
		_w35936_,
		_w35939_,
		_w35940_
	);
	LUT2 #(
		.INIT('h8)
	) name25429 (
		_w15698_,
		_w31950_,
		_w35941_
	);
	LUT2 #(
		.INIT('h1)
	) name25430 (
		\wishbone_rx_fifo_read_pointer_reg[0]/NET0131 ,
		_w35640_,
		_w35942_
	);
	LUT2 #(
		.INIT('h1)
	) name25431 (
		_w31950_,
		_w35641_,
		_w35943_
	);
	LUT2 #(
		.INIT('h4)
	) name25432 (
		_w35942_,
		_w35943_,
		_w35944_
	);
	LUT2 #(
		.INIT('h1)
	) name25433 (
		_w35941_,
		_w35944_,
		_w35945_
	);
	LUT2 #(
		.INIT('h8)
	) name25434 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[1]/NET0131 ,
		_w34204_,
		_w35946_
	);
	LUT2 #(
		.INIT('h1)
	) name25435 (
		\wishbone_RxBDAddress_reg[2]/NET0131 ,
		_w34593_,
		_w35947_
	);
	LUT2 #(
		.INIT('h1)
	) name25436 (
		_w34204_,
		_w34594_,
		_w35948_
	);
	LUT2 #(
		.INIT('h4)
	) name25437 (
		_w35947_,
		_w35948_,
		_w35949_
	);
	LUT2 #(
		.INIT('h1)
	) name25438 (
		_w35946_,
		_w35949_,
		_w35950_
	);
	LUT2 #(
		.INIT('h8)
	) name25439 (
		\wb_dat_i[10]_pad ,
		_w34989_,
		_w35951_
	);
	LUT2 #(
		.INIT('h8)
	) name25440 (
		\wishbone_ram_di_reg[10]/NET0131 ,
		_w34991_,
		_w35952_
	);
	LUT2 #(
		.INIT('h1)
	) name25441 (
		_w35951_,
		_w35952_,
		_w35953_
	);
	LUT2 #(
		.INIT('h8)
	) name25442 (
		\wb_dat_i[15]_pad ,
		_w34989_,
		_w35954_
	);
	LUT2 #(
		.INIT('h8)
	) name25443 (
		\wishbone_ram_di_reg[15]/NET0131 ,
		_w34991_,
		_w35955_
	);
	LUT2 #(
		.INIT('h1)
	) name25444 (
		_w35954_,
		_w35955_,
		_w35956_
	);
	LUT2 #(
		.INIT('h8)
	) name25445 (
		\wb_dat_i[9]_pad ,
		_w34989_,
		_w35957_
	);
	LUT2 #(
		.INIT('h8)
	) name25446 (
		\wishbone_ram_di_reg[9]/NET0131 ,
		_w34991_,
		_w35958_
	);
	LUT2 #(
		.INIT('h1)
	) name25447 (
		_w35957_,
		_w35958_,
		_w35959_
	);
	LUT2 #(
		.INIT('h8)
	) name25448 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11525_,
		_w35960_
	);
	LUT2 #(
		.INIT('h4)
	) name25449 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[8]/NET0131 ,
		_w35961_
	);
	LUT2 #(
		.INIT('h1)
	) name25450 (
		_w35960_,
		_w35961_,
		_w35962_
	);
	LUT2 #(
		.INIT('h2)
	) name25451 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w11518_,
		_w35963_
	);
	LUT2 #(
		.INIT('h1)
	) name25452 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		\wishbone_LatchedRxLength_reg[7]/NET0131 ,
		_w35964_
	);
	LUT2 #(
		.INIT('h1)
	) name25453 (
		_w35963_,
		_w35964_,
		_w35965_
	);
	LUT2 #(
		.INIT('h2)
	) name25454 (
		\txethmac1_TxRetry_reg/NET0131 ,
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w35966_
	);
	LUT2 #(
		.INIT('h2)
	) name25455 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		\wishbone_TxUsedData_q_reg/NET0131 ,
		_w35967_
	);
	LUT2 #(
		.INIT('h4)
	) name25456 (
		_w35966_,
		_w35967_,
		_w35968_
	);
	LUT2 #(
		.INIT('h1)
	) name25457 (
		\wishbone_TxStartFrm_sync2_reg/NET0131 ,
		_w35968_,
		_w35969_
	);
	LUT2 #(
		.INIT('h1)
	) name25458 (
		\wishbone_rx_fifo_read_pointer_reg[1]/NET0131 ,
		_w35641_,
		_w35970_
	);
	LUT2 #(
		.INIT('h1)
	) name25459 (
		_w31950_,
		_w35642_,
		_w35971_
	);
	LUT2 #(
		.INIT('h4)
	) name25460 (
		_w35970_,
		_w35971_,
		_w35972_
	);
	LUT2 #(
		.INIT('h8)
	) name25461 (
		\wb_adr_i[4]_pad ,
		\wb_adr_i[5]_pad ,
		_w35973_
	);
	LUT2 #(
		.INIT('h8)
	) name25462 (
		_w35890_,
		_w35973_,
		_w35974_
	);
	LUT2 #(
		.INIT('h8)
	) name25463 (
		_w34525_,
		_w35974_,
		_w35975_
	);
	LUT2 #(
		.INIT('h8)
	) name25464 (
		_w31683_,
		_w35912_,
		_w35976_
	);
	LUT2 #(
		.INIT('h8)
	) name25465 (
		_w22963_,
		_w35976_,
		_w35977_
	);
	LUT2 #(
		.INIT('h8)
	) name25466 (
		_w35974_,
		_w35977_,
		_w35978_
	);
	LUT2 #(
		.INIT('h8)
	) name25467 (
		_w34133_,
		_w34135_,
		_w35979_
	);
	LUT2 #(
		.INIT('h1)
	) name25468 (
		\wishbone_RxOverrun_reg/NET0131 ,
		_w35979_,
		_w35980_
	);
	LUT2 #(
		.INIT('h1)
	) name25469 (
		_w34201_,
		_w35980_,
		_w35981_
	);
	LUT2 #(
		.INIT('h8)
	) name25470 (
		_w34085_,
		_w34089_,
		_w35982_
	);
	LUT2 #(
		.INIT('h1)
	) name25471 (
		\wishbone_TxUnderRun_wb_reg/NET0131 ,
		_w35982_,
		_w35983_
	);
	LUT2 #(
		.INIT('h1)
	) name25472 (
		_w34287_,
		_w35983_,
		_w35984_
	);
	LUT2 #(
		.INIT('h8)
	) name25473 (
		_w24730_,
		_w31684_,
		_w35985_
	);
	LUT2 #(
		.INIT('h8)
	) name25474 (
		_w24730_,
		_w35705_,
		_w35986_
	);
	LUT2 #(
		.INIT('h4)
	) name25475 (
		\ethreg1_MODER_0_DataOut_reg[5]/NET0131 ,
		_w35724_,
		_w35987_
	);
	LUT2 #(
		.INIT('h8)
	) name25476 (
		_w12512_,
		_w35987_,
		_w35988_
	);
	LUT2 #(
		.INIT('h8)
	) name25477 (
		_w23501_,
		_w31684_,
		_w35989_
	);
	LUT2 #(
		.INIT('h1)
	) name25478 (
		\rxethmac1_rxcounters1_DlyCrcCnt_reg[1]/NET0131 ,
		_w34862_,
		_w35990_
	);
	LUT2 #(
		.INIT('h1)
	) name25479 (
		_w34863_,
		_w35990_,
		_w35991_
	);
	LUT2 #(
		.INIT('h8)
	) name25480 (
		_w34861_,
		_w35991_,
		_w35992_
	);
	LUT2 #(
		.INIT('h8)
	) name25481 (
		_w23501_,
		_w35976_,
		_w35993_
	);
	LUT2 #(
		.INIT('h2)
	) name25482 (
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		\maccontrol1_receivecontrol1_Divider2_reg/NET0131 ,
		_w35994_
	);
	LUT2 #(
		.INIT('h4)
	) name25483 (
		_w11640_,
		_w35994_,
		_w35995_
	);
	LUT2 #(
		.INIT('h1)
	) name25484 (
		\wishbone_rx_fifo_read_pointer_reg[2]/NET0131 ,
		_w35642_,
		_w35996_
	);
	LUT2 #(
		.INIT('h1)
	) name25485 (
		_w31950_,
		_w35643_,
		_w35997_
	);
	LUT2 #(
		.INIT('h4)
	) name25486 (
		_w35996_,
		_w35997_,
		_w35998_
	);
	LUT2 #(
		.INIT('h4)
	) name25487 (
		\wb_adr_i[2]_pad ,
		_w23498_,
		_w35999_
	);
	LUT2 #(
		.INIT('h8)
	) name25488 (
		_w34525_,
		_w35999_,
		_w36000_
	);
	LUT2 #(
		.INIT('h1)
	) name25489 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[5]/NET0131 ,
		_w11624_,
		_w36001_
	);
	LUT2 #(
		.INIT('h1)
	) name25490 (
		wb_rst_i_pad,
		_w11625_,
		_w36002_
	);
	LUT2 #(
		.INIT('h4)
	) name25491 (
		_w36001_,
		_w36002_,
		_w36003_
	);
	LUT2 #(
		.INIT('h2)
	) name25492 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		_w36004_
	);
	LUT2 #(
		.INIT('h8)
	) name25493 (
		\txethmac1_TxUsedData_reg/NET0131 ,
		_w36004_,
		_w36005_
	);
	LUT2 #(
		.INIT('h8)
	) name25494 (
		_w34268_,
		_w36005_,
		_w36006_
	);
	LUT2 #(
		.INIT('h1)
	) name25495 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[2]/NET0131 ,
		_w36006_,
		_w36007_
	);
	LUT2 #(
		.INIT('h2)
	) name25496 (
		_w34259_,
		_w36007_,
		_w36008_
	);
	LUT2 #(
		.INIT('h2)
	) name25497 (
		_w11110_,
		_w11222_,
		_w36009_
	);
	LUT2 #(
		.INIT('h2)
	) name25498 (
		\txethmac1_random1_RandomLatched_reg[5]/NET0131 ,
		_w34968_,
		_w36010_
	);
	LUT2 #(
		.INIT('h8)
	) name25499 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w36011_
	);
	LUT2 #(
		.INIT('h1)
	) name25500 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w36011_,
		_w36012_
	);
	LUT2 #(
		.INIT('h8)
	) name25501 (
		\txethmac1_random1_x_reg[5]/NET0131 ,
		_w34968_,
		_w36013_
	);
	LUT2 #(
		.INIT('h4)
	) name25502 (
		_w36012_,
		_w36013_,
		_w36014_
	);
	LUT2 #(
		.INIT('h1)
	) name25503 (
		_w36010_,
		_w36014_,
		_w36015_
	);
	LUT2 #(
		.INIT('h8)
	) name25504 (
		_w24729_,
		_w35892_,
		_w36016_
	);
	LUT2 #(
		.INIT('h2)
	) name25505 (
		_w11181_,
		_w11400_,
		_w36017_
	);
	LUT2 #(
		.INIT('h2)
	) name25506 (
		\wishbone_BDWrite_reg[3]/NET0131 ,
		_w34989_,
		_w36018_
	);
	LUT2 #(
		.INIT('h8)
	) name25507 (
		\wb_sel_i[3]_pad ,
		_w22942_,
		_w36019_
	);
	LUT2 #(
		.INIT('h8)
	) name25508 (
		_w35908_,
		_w36019_,
		_w36020_
	);
	LUT2 #(
		.INIT('h1)
	) name25509 (
		_w36018_,
		_w36020_,
		_w36021_
	);
	LUT2 #(
		.INIT('h8)
	) name25510 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		_w36022_
	);
	LUT2 #(
		.INIT('h1)
	) name25511 (
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		_w34892_,
		_w36023_
	);
	LUT2 #(
		.INIT('h1)
	) name25512 (
		\wishbone_BlockingTxBDRead_reg/NET0131 ,
		_w36023_,
		_w36024_
	);
	LUT2 #(
		.INIT('h4)
	) name25513 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w36024_,
		_w36025_
	);
	LUT2 #(
		.INIT('h1)
	) name25514 (
		_w36022_,
		_w36025_,
		_w36026_
	);
	LUT2 #(
		.INIT('h4)
	) name25515 (
		\wishbone_TxStartFrm_syncb2_reg/NET0131 ,
		\wishbone_TxStartFrm_wb_reg/NET0131 ,
		_w36027_
	);
	LUT2 #(
		.INIT('h1)
	) name25516 (
		_w34446_,
		_w34916_,
		_w36028_
	);
	LUT2 #(
		.INIT('h4)
	) name25517 (
		\wishbone_StartOccured_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		_w36029_
	);
	LUT2 #(
		.INIT('h4)
	) name25518 (
		_w36028_,
		_w36029_,
		_w36030_
	);
	LUT2 #(
		.INIT('h1)
	) name25519 (
		_w36027_,
		_w36030_,
		_w36031_
	);
	LUT2 #(
		.INIT('h8)
	) name25520 (
		_w31685_,
		_w35973_,
		_w36032_
	);
	LUT2 #(
		.INIT('h8)
	) name25521 (
		_w34525_,
		_w36032_,
		_w36033_
	);
	LUT2 #(
		.INIT('h8)
	) name25522 (
		_w35977_,
		_w36032_,
		_w36034_
	);
	LUT2 #(
		.INIT('h8)
	) name25523 (
		_w22961_,
		_w31686_,
		_w36035_
	);
	LUT2 #(
		.INIT('h8)
	) name25524 (
		_w34525_,
		_w36035_,
		_w36036_
	);
	LUT2 #(
		.INIT('h8)
	) name25525 (
		_w35977_,
		_w36035_,
		_w36037_
	);
	LUT2 #(
		.INIT('h8)
	) name25526 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[1]/NET0131 ,
		_w35622_,
		_w36038_
	);
	LUT2 #(
		.INIT('h8)
	) name25527 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[1]/NET0131 ,
		_w35827_,
		_w36039_
	);
	LUT2 #(
		.INIT('h8)
	) name25528 (
		\ethreg1_TXCTRL_0_DataOut_reg[1]/NET0131 ,
		_w34266_,
		_w36040_
	);
	LUT2 #(
		.INIT('h8)
	) name25529 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[1]/NET0131 ,
		_w35625_,
		_w36041_
	);
	LUT2 #(
		.INIT('h8)
	) name25530 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[1]/NET0131 ,
		_w35627_,
		_w36042_
	);
	LUT2 #(
		.INIT('h8)
	) name25531 (
		\ethreg1_TXCTRL_1_DataOut_reg[1]/NET0131 ,
		_w35830_,
		_w36043_
	);
	LUT2 #(
		.INIT('h8)
	) name25532 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[1]/NET0131 ,
		_w34938_,
		_w36044_
	);
	LUT2 #(
		.INIT('h8)
	) name25533 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[1]/NET0131 ,
		_w34955_,
		_w36045_
	);
	LUT2 #(
		.INIT('h8)
	) name25534 (
		_w34937_,
		_w34949_,
		_w36046_
	);
	LUT2 #(
		.INIT('h1)
	) name25535 (
		_w36038_,
		_w36046_,
		_w36047_
	);
	LUT2 #(
		.INIT('h1)
	) name25536 (
		_w36039_,
		_w36040_,
		_w36048_
	);
	LUT2 #(
		.INIT('h1)
	) name25537 (
		_w36041_,
		_w36042_,
		_w36049_
	);
	LUT2 #(
		.INIT('h1)
	) name25538 (
		_w36043_,
		_w36044_,
		_w36050_
	);
	LUT2 #(
		.INIT('h4)
	) name25539 (
		_w36045_,
		_w36050_,
		_w36051_
	);
	LUT2 #(
		.INIT('h8)
	) name25540 (
		_w36048_,
		_w36049_,
		_w36052_
	);
	LUT2 #(
		.INIT('h8)
	) name25541 (
		_w36047_,
		_w36052_,
		_w36053_
	);
	LUT2 #(
		.INIT('h8)
	) name25542 (
		_w36051_,
		_w36053_,
		_w36054_
	);
	LUT2 #(
		.INIT('h8)
	) name25543 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[6]/NET0131 ,
		_w35622_,
		_w36055_
	);
	LUT2 #(
		.INIT('h8)
	) name25544 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[6]/NET0131 ,
		_w35827_,
		_w36056_
	);
	LUT2 #(
		.INIT('h8)
	) name25545 (
		\ethreg1_TXCTRL_0_DataOut_reg[6]/NET0131 ,
		_w34266_,
		_w36057_
	);
	LUT2 #(
		.INIT('h8)
	) name25546 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[6]/NET0131 ,
		_w35625_,
		_w36058_
	);
	LUT2 #(
		.INIT('h8)
	) name25547 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[6]/NET0131 ,
		_w35627_,
		_w36059_
	);
	LUT2 #(
		.INIT('h8)
	) name25548 (
		\ethreg1_TXCTRL_1_DataOut_reg[6]/NET0131 ,
		_w35830_,
		_w36060_
	);
	LUT2 #(
		.INIT('h8)
	) name25549 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[6]/NET0131 ,
		_w34938_,
		_w36061_
	);
	LUT2 #(
		.INIT('h8)
	) name25550 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[6]/NET0131 ,
		_w34955_,
		_w36062_
	);
	LUT2 #(
		.INIT('h1)
	) name25551 (
		_w36046_,
		_w36055_,
		_w36063_
	);
	LUT2 #(
		.INIT('h1)
	) name25552 (
		_w36056_,
		_w36057_,
		_w36064_
	);
	LUT2 #(
		.INIT('h1)
	) name25553 (
		_w36058_,
		_w36059_,
		_w36065_
	);
	LUT2 #(
		.INIT('h1)
	) name25554 (
		_w36060_,
		_w36061_,
		_w36066_
	);
	LUT2 #(
		.INIT('h4)
	) name25555 (
		_w36062_,
		_w36066_,
		_w36067_
	);
	LUT2 #(
		.INIT('h8)
	) name25556 (
		_w36064_,
		_w36065_,
		_w36068_
	);
	LUT2 #(
		.INIT('h8)
	) name25557 (
		_w36063_,
		_w36068_,
		_w36069_
	);
	LUT2 #(
		.INIT('h8)
	) name25558 (
		_w36067_,
		_w36069_,
		_w36070_
	);
	LUT2 #(
		.INIT('h8)
	) name25559 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w11273_,
		_w36071_
	);
	LUT2 #(
		.INIT('h1)
	) name25560 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w36071_,
		_w36072_
	);
	LUT2 #(
		.INIT('h2)
	) name25561 (
		\txethmac1_random1_x_reg[6]/NET0131 ,
		_w36072_,
		_w36073_
	);
	LUT2 #(
		.INIT('h2)
	) name25562 (
		_w34968_,
		_w36073_,
		_w36074_
	);
	LUT2 #(
		.INIT('h1)
	) name25563 (
		\txethmac1_random1_RandomLatched_reg[6]/NET0131 ,
		_w34968_,
		_w36075_
	);
	LUT2 #(
		.INIT('h1)
	) name25564 (
		_w36074_,
		_w36075_,
		_w36076_
	);
	LUT2 #(
		.INIT('h1)
	) name25565 (
		\wishbone_TxBDRead_reg/NET0131 ,
		_w36024_,
		_w36077_
	);
	LUT2 #(
		.INIT('h1)
	) name25566 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w36077_,
		_w36078_
	);
	LUT2 #(
		.INIT('h4)
	) name25567 (
		\wishbone_TxRetryPacketBlocked_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w36079_
	);
	LUT2 #(
		.INIT('h4)
	) name25568 (
		_w35931_,
		_w36079_,
		_w36080_
	);
	LUT2 #(
		.INIT('h1)
	) name25569 (
		\wishbone_TxRetryPacket_NotCleared_reg/NET0131 ,
		_w36080_,
		_w36081_
	);
	LUT2 #(
		.INIT('h1)
	) name25570 (
		_w36025_,
		_w36081_,
		_w36082_
	);
	LUT2 #(
		.INIT('h1)
	) name25571 (
		\wishbone_Flop_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w36083_
	);
	LUT2 #(
		.INIT('h1)
	) name25572 (
		\wishbone_TxRetry_q_reg/NET0131 ,
		_w35898_,
		_w36084_
	);
	LUT2 #(
		.INIT('h1)
	) name25573 (
		_w12249_,
		_w12251_,
		_w36085_
	);
	LUT2 #(
		.INIT('h1)
	) name25574 (
		\wishbone_TxValidBytesLatched_reg[1]/NET0131 ,
		_w36085_,
		_w36086_
	);
	LUT2 #(
		.INIT('h8)
	) name25575 (
		\wishbone_TxValidBytesLatched_reg[1]/NET0131 ,
		_w36085_,
		_w36087_
	);
	LUT2 #(
		.INIT('h2)
	) name25576 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxValidBytesLatched_reg[0]/NET0131 ,
		_w36088_
	);
	LUT2 #(
		.INIT('h4)
	) name25577 (
		\wishbone_TxByteCnt_reg[0]/NET0131 ,
		\wishbone_TxValidBytesLatched_reg[0]/NET0131 ,
		_w36089_
	);
	LUT2 #(
		.INIT('h1)
	) name25578 (
		_w36088_,
		_w36089_,
		_w36090_
	);
	LUT2 #(
		.INIT('h2)
	) name25579 (
		\wishbone_LastWord_reg/NET0131 ,
		\wishbone_TxEndFrm_reg/NET0131 ,
		_w36091_
	);
	LUT2 #(
		.INIT('h4)
	) name25580 (
		_w36090_,
		_w36091_,
		_w36092_
	);
	LUT2 #(
		.INIT('h4)
	) name25581 (
		_w36086_,
		_w36092_,
		_w36093_
	);
	LUT2 #(
		.INIT('h4)
	) name25582 (
		_w36087_,
		_w36093_,
		_w36094_
	);
	LUT2 #(
		.INIT('h2)
	) name25583 (
		\wishbone_Flop_reg/NET0131 ,
		_w36094_,
		_w36095_
	);
	LUT2 #(
		.INIT('h4)
	) name25584 (
		_w36083_,
		_w36084_,
		_w36096_
	);
	LUT2 #(
		.INIT('h4)
	) name25585 (
		_w36095_,
		_w36096_,
		_w36097_
	);
	LUT2 #(
		.INIT('h8)
	) name25586 (
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w36098_
	);
	LUT2 #(
		.INIT('h8)
	) name25587 (
		\wishbone_BDWrite_reg[1]/NET0131 ,
		_w36098_,
		_w36099_
	);
	LUT2 #(
		.INIT('h1)
	) name25588 (
		_w34201_,
		_w34892_,
		_w36100_
	);
	LUT2 #(
		.INIT('h4)
	) name25589 (
		_w36099_,
		_w36100_,
		_w36101_
	);
	LUT2 #(
		.INIT('h1)
	) name25590 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w36102_
	);
	LUT2 #(
		.INIT('h8)
	) name25591 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w36103_
	);
	LUT2 #(
		.INIT('h8)
	) name25592 (
		_w36102_,
		_w36103_,
		_w36104_
	);
	LUT2 #(
		.INIT('h2)
	) name25593 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w36105_
	);
	LUT2 #(
		.INIT('h4)
	) name25594 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w36106_
	);
	LUT2 #(
		.INIT('h8)
	) name25595 (
		_w36105_,
		_w36106_,
		_w36107_
	);
	LUT2 #(
		.INIT('h8)
	) name25596 (
		_w36104_,
		_w36107_,
		_w36108_
	);
	LUT2 #(
		.INIT('h4)
	) name25597 (
		_w36101_,
		_w36108_,
		_w36109_
	);
	LUT2 #(
		.INIT('h8)
	) name25598 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		_w36098_,
		_w36110_
	);
	LUT2 #(
		.INIT('h2)
	) name25599 (
		_w36100_,
		_w36110_,
		_w36111_
	);
	LUT2 #(
		.INIT('h8)
	) name25600 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w36112_
	);
	LUT2 #(
		.INIT('h1)
	) name25601 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w36113_
	);
	LUT2 #(
		.INIT('h8)
	) name25602 (
		_w36112_,
		_w36113_,
		_w36114_
	);
	LUT2 #(
		.INIT('h8)
	) name25603 (
		_w36104_,
		_w36114_,
		_w36115_
	);
	LUT2 #(
		.INIT('h4)
	) name25604 (
		_w36111_,
		_w36115_,
		_w36116_
	);
	LUT2 #(
		.INIT('h8)
	) name25605 (
		_w36105_,
		_w36112_,
		_w36117_
	);
	LUT2 #(
		.INIT('h4)
	) name25606 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w36118_
	);
	LUT2 #(
		.INIT('h8)
	) name25607 (
		_w36102_,
		_w36118_,
		_w36119_
	);
	LUT2 #(
		.INIT('h8)
	) name25608 (
		_w36117_,
		_w36119_,
		_w36120_
	);
	LUT2 #(
		.INIT('h4)
	) name25609 (
		_w36111_,
		_w36120_,
		_w36121_
	);
	LUT2 #(
		.INIT('h2)
	) name25610 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w36122_
	);
	LUT2 #(
		.INIT('h8)
	) name25611 (
		_w36103_,
		_w36122_,
		_w36123_
	);
	LUT2 #(
		.INIT('h8)
	) name25612 (
		_w36106_,
		_w36113_,
		_w36124_
	);
	LUT2 #(
		.INIT('h8)
	) name25613 (
		_w36123_,
		_w36124_,
		_w36125_
	);
	LUT2 #(
		.INIT('h4)
	) name25614 (
		_w36111_,
		_w36125_,
		_w36126_
	);
	LUT2 #(
		.INIT('h8)
	) name25615 (
		_w36118_,
		_w36122_,
		_w36127_
	);
	LUT2 #(
		.INIT('h8)
	) name25616 (
		_w36107_,
		_w36127_,
		_w36128_
	);
	LUT2 #(
		.INIT('h4)
	) name25617 (
		_w36111_,
		_w36128_,
		_w36129_
	);
	LUT2 #(
		.INIT('h8)
	) name25618 (
		_w36114_,
		_w36127_,
		_w36130_
	);
	LUT2 #(
		.INIT('h4)
	) name25619 (
		_w36111_,
		_w36130_,
		_w36131_
	);
	LUT2 #(
		.INIT('h8)
	) name25620 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		_w36098_,
		_w36132_
	);
	LUT2 #(
		.INIT('h2)
	) name25621 (
		_w36100_,
		_w36132_,
		_w36133_
	);
	LUT2 #(
		.INIT('h1)
	) name25622 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w36134_
	);
	LUT2 #(
		.INIT('h8)
	) name25623 (
		_w36105_,
		_w36134_,
		_w36135_
	);
	LUT2 #(
		.INIT('h8)
	) name25624 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w36136_
	);
	LUT2 #(
		.INIT('h8)
	) name25625 (
		_w36103_,
		_w36136_,
		_w36137_
	);
	LUT2 #(
		.INIT('h8)
	) name25626 (
		_w36135_,
		_w36137_,
		_w36138_
	);
	LUT2 #(
		.INIT('h4)
	) name25627 (
		_w36133_,
		_w36138_,
		_w36139_
	);
	LUT2 #(
		.INIT('h4)
	) name25628 (
		\wishbone_ram_addr_reg[3]/NET0131 ,
		\wishbone_ram_addr_reg[4]/NET0131 ,
		_w36140_
	);
	LUT2 #(
		.INIT('h8)
	) name25629 (
		_w36103_,
		_w36140_,
		_w36141_
	);
	LUT2 #(
		.INIT('h8)
	) name25630 (
		_w36124_,
		_w36141_,
		_w36142_
	);
	LUT2 #(
		.INIT('h4)
	) name25631 (
		_w36111_,
		_w36142_,
		_w36143_
	);
	LUT2 #(
		.INIT('h8)
	) name25632 (
		_w36118_,
		_w36140_,
		_w36144_
	);
	LUT2 #(
		.INIT('h8)
	) name25633 (
		_w36107_,
		_w36144_,
		_w36145_
	);
	LUT2 #(
		.INIT('h4)
	) name25634 (
		_w36111_,
		_w36145_,
		_w36146_
	);
	LUT2 #(
		.INIT('h8)
	) name25635 (
		_w36114_,
		_w36144_,
		_w36147_
	);
	LUT2 #(
		.INIT('h4)
	) name25636 (
		_w36111_,
		_w36147_,
		_w36148_
	);
	LUT2 #(
		.INIT('h8)
	) name25637 (
		_w36118_,
		_w36136_,
		_w36149_
	);
	LUT2 #(
		.INIT('h8)
	) name25638 (
		_w36124_,
		_w36149_,
		_w36150_
	);
	LUT2 #(
		.INIT('h4)
	) name25639 (
		_w36111_,
		_w36150_,
		_w36151_
	);
	LUT2 #(
		.INIT('h8)
	) name25640 (
		_w36124_,
		_w36137_,
		_w36152_
	);
	LUT2 #(
		.INIT('h4)
	) name25641 (
		_w36111_,
		_w36152_,
		_w36153_
	);
	LUT2 #(
		.INIT('h8)
	) name25642 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w36154_
	);
	LUT2 #(
		.INIT('h2)
	) name25643 (
		\wishbone_ram_addr_reg[2]/NET0131 ,
		\wishbone_ram_addr_reg[5]/NET0131 ,
		_w36155_
	);
	LUT2 #(
		.INIT('h8)
	) name25644 (
		_w36154_,
		_w36155_,
		_w36156_
	);
	LUT2 #(
		.INIT('h1)
	) name25645 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w36157_
	);
	LUT2 #(
		.INIT('h8)
	) name25646 (
		_w36102_,
		_w36157_,
		_w36158_
	);
	LUT2 #(
		.INIT('h8)
	) name25647 (
		_w36156_,
		_w36158_,
		_w36159_
	);
	LUT2 #(
		.INIT('h4)
	) name25648 (
		_w36111_,
		_w36159_,
		_w36160_
	);
	LUT2 #(
		.INIT('h2)
	) name25649 (
		\wishbone_ram_addr_reg[0]/NET0131 ,
		\wishbone_ram_addr_reg[6]/NET0131 ,
		_w36161_
	);
	LUT2 #(
		.INIT('h8)
	) name25650 (
		_w36102_,
		_w36161_,
		_w36162_
	);
	LUT2 #(
		.INIT('h8)
	) name25651 (
		_w36156_,
		_w36162_,
		_w36163_
	);
	LUT2 #(
		.INIT('h4)
	) name25652 (
		_w36111_,
		_w36163_,
		_w36164_
	);
	LUT2 #(
		.INIT('h8)
	) name25653 (
		_w36134_,
		_w36154_,
		_w36165_
	);
	LUT2 #(
		.INIT('h8)
	) name25654 (
		_w36122_,
		_w36161_,
		_w36166_
	);
	LUT2 #(
		.INIT('h8)
	) name25655 (
		_w36165_,
		_w36166_,
		_w36167_
	);
	LUT2 #(
		.INIT('h4)
	) name25656 (
		_w36111_,
		_w36167_,
		_w36168_
	);
	LUT2 #(
		.INIT('h4)
	) name25657 (
		\wishbone_ram_addr_reg[1]/NET0131 ,
		\wishbone_ram_addr_reg[7]/NET0131 ,
		_w36169_
	);
	LUT2 #(
		.INIT('h8)
	) name25658 (
		_w36155_,
		_w36169_,
		_w36170_
	);
	LUT2 #(
		.INIT('h8)
	) name25659 (
		_w36166_,
		_w36170_,
		_w36171_
	);
	LUT2 #(
		.INIT('h4)
	) name25660 (
		_w36111_,
		_w36171_,
		_w36172_
	);
	LUT2 #(
		.INIT('h8)
	) name25661 (
		_w36122_,
		_w36157_,
		_w36173_
	);
	LUT2 #(
		.INIT('h8)
	) name25662 (
		_w36156_,
		_w36173_,
		_w36174_
	);
	LUT2 #(
		.INIT('h4)
	) name25663 (
		_w36111_,
		_w36174_,
		_w36175_
	);
	LUT2 #(
		.INIT('h8)
	) name25664 (
		_w36140_,
		_w36161_,
		_w36176_
	);
	LUT2 #(
		.INIT('h8)
	) name25665 (
		_w36165_,
		_w36176_,
		_w36177_
	);
	LUT2 #(
		.INIT('h4)
	) name25666 (
		_w36111_,
		_w36177_,
		_w36178_
	);
	LUT2 #(
		.INIT('h8)
	) name25667 (
		_w36170_,
		_w36176_,
		_w36179_
	);
	LUT2 #(
		.INIT('h4)
	) name25668 (
		_w36111_,
		_w36179_,
		_w36180_
	);
	LUT2 #(
		.INIT('h8)
	) name25669 (
		_w36140_,
		_w36157_,
		_w36181_
	);
	LUT2 #(
		.INIT('h8)
	) name25670 (
		_w36156_,
		_w36181_,
		_w36182_
	);
	LUT2 #(
		.INIT('h4)
	) name25671 (
		_w36111_,
		_w36182_,
		_w36183_
	);
	LUT2 #(
		.INIT('h4)
	) name25672 (
		_w36101_,
		_w36159_,
		_w36184_
	);
	LUT2 #(
		.INIT('h8)
	) name25673 (
		_w36134_,
		_w36169_,
		_w36185_
	);
	LUT2 #(
		.INIT('h8)
	) name25674 (
		_w36136_,
		_w36161_,
		_w36186_
	);
	LUT2 #(
		.INIT('h8)
	) name25675 (
		_w36185_,
		_w36186_,
		_w36187_
	);
	LUT2 #(
		.INIT('h4)
	) name25676 (
		_w36111_,
		_w36187_,
		_w36188_
	);
	LUT2 #(
		.INIT('h8)
	) name25677 (
		_w36136_,
		_w36157_,
		_w36189_
	);
	LUT2 #(
		.INIT('h8)
	) name25678 (
		_w36165_,
		_w36189_,
		_w36190_
	);
	LUT2 #(
		.INIT('h4)
	) name25679 (
		_w36111_,
		_w36190_,
		_w36191_
	);
	LUT2 #(
		.INIT('h8)
	) name25680 (
		_w36170_,
		_w36189_,
		_w36192_
	);
	LUT2 #(
		.INIT('h4)
	) name25681 (
		_w36111_,
		_w36192_,
		_w36193_
	);
	LUT2 #(
		.INIT('h8)
	) name25682 (
		_w36105_,
		_w36155_,
		_w36194_
	);
	LUT2 #(
		.INIT('h8)
	) name25683 (
		_w36166_,
		_w36194_,
		_w36195_
	);
	LUT2 #(
		.INIT('h4)
	) name25684 (
		_w36111_,
		_w36195_,
		_w36196_
	);
	LUT2 #(
		.INIT('h8)
	) name25685 (
		_w36106_,
		_w36154_,
		_w36197_
	);
	LUT2 #(
		.INIT('h8)
	) name25686 (
		_w36158_,
		_w36197_,
		_w36198_
	);
	LUT2 #(
		.INIT('h4)
	) name25687 (
		_w36111_,
		_w36198_,
		_w36199_
	);
	LUT2 #(
		.INIT('h8)
	) name25688 (
		_w36162_,
		_w36197_,
		_w36200_
	);
	LUT2 #(
		.INIT('h4)
	) name25689 (
		_w36111_,
		_w36200_,
		_w36201_
	);
	LUT2 #(
		.INIT('h8)
	) name25690 (
		_w36112_,
		_w36169_,
		_w36202_
	);
	LUT2 #(
		.INIT('h8)
	) name25691 (
		_w36158_,
		_w36202_,
		_w36203_
	);
	LUT2 #(
		.INIT('h4)
	) name25692 (
		_w36111_,
		_w36203_,
		_w36204_
	);
	LUT2 #(
		.INIT('h8)
	) name25693 (
		_w36162_,
		_w36202_,
		_w36205_
	);
	LUT2 #(
		.INIT('h4)
	) name25694 (
		_w36111_,
		_w36205_,
		_w36206_
	);
	LUT2 #(
		.INIT('h8)
	) name25695 (
		_w36112_,
		_w36154_,
		_w36207_
	);
	LUT2 #(
		.INIT('h8)
	) name25696 (
		_w36158_,
		_w36207_,
		_w36208_
	);
	LUT2 #(
		.INIT('h4)
	) name25697 (
		_w36111_,
		_w36208_,
		_w36209_
	);
	LUT2 #(
		.INIT('h8)
	) name25698 (
		_w36162_,
		_w36207_,
		_w36210_
	);
	LUT2 #(
		.INIT('h4)
	) name25699 (
		_w36111_,
		_w36210_,
		_w36211_
	);
	LUT2 #(
		.INIT('h8)
	) name25700 (
		_w36106_,
		_w36169_,
		_w36212_
	);
	LUT2 #(
		.INIT('h8)
	) name25701 (
		_w36166_,
		_w36212_,
		_w36213_
	);
	LUT2 #(
		.INIT('h4)
	) name25702 (
		_w36111_,
		_w36213_,
		_w36214_
	);
	LUT2 #(
		.INIT('h8)
	) name25703 (
		_w36173_,
		_w36197_,
		_w36215_
	);
	LUT2 #(
		.INIT('h4)
	) name25704 (
		_w36111_,
		_w36215_,
		_w36216_
	);
	LUT2 #(
		.INIT('h8)
	) name25705 (
		_w36173_,
		_w36202_,
		_w36217_
	);
	LUT2 #(
		.INIT('h4)
	) name25706 (
		_w36111_,
		_w36217_,
		_w36218_
	);
	LUT2 #(
		.INIT('h8)
	) name25707 (
		_w36173_,
		_w36207_,
		_w36219_
	);
	LUT2 #(
		.INIT('h4)
	) name25708 (
		_w36111_,
		_w36219_,
		_w36220_
	);
	LUT2 #(
		.INIT('h8)
	) name25709 (
		_w36176_,
		_w36212_,
		_w36221_
	);
	LUT2 #(
		.INIT('h4)
	) name25710 (
		_w36111_,
		_w36221_,
		_w36222_
	);
	LUT2 #(
		.INIT('h8)
	) name25711 (
		_w36181_,
		_w36197_,
		_w36223_
	);
	LUT2 #(
		.INIT('h4)
	) name25712 (
		_w36111_,
		_w36223_,
		_w36224_
	);
	LUT2 #(
		.INIT('h8)
	) name25713 (
		_w36181_,
		_w36202_,
		_w36225_
	);
	LUT2 #(
		.INIT('h4)
	) name25714 (
		_w36111_,
		_w36225_,
		_w36226_
	);
	LUT2 #(
		.INIT('h8)
	) name25715 (
		_w36181_,
		_w36207_,
		_w36227_
	);
	LUT2 #(
		.INIT('h4)
	) name25716 (
		_w36111_,
		_w36227_,
		_w36228_
	);
	LUT2 #(
		.INIT('h8)
	) name25717 (
		_w36189_,
		_w36212_,
		_w36229_
	);
	LUT2 #(
		.INIT('h4)
	) name25718 (
		_w36111_,
		_w36229_,
		_w36230_
	);
	LUT2 #(
		.INIT('h8)
	) name25719 (
		_w36104_,
		_w36165_,
		_w36231_
	);
	LUT2 #(
		.INIT('h4)
	) name25720 (
		_w36111_,
		_w36231_,
		_w36232_
	);
	LUT2 #(
		.INIT('h8)
	) name25721 (
		_w36104_,
		_w36170_,
		_w36233_
	);
	LUT2 #(
		.INIT('h4)
	) name25722 (
		_w36111_,
		_w36233_,
		_w36234_
	);
	LUT2 #(
		.INIT('h8)
	) name25723 (
		_w36119_,
		_w36156_,
		_w36235_
	);
	LUT2 #(
		.INIT('h4)
	) name25724 (
		_w36111_,
		_w36235_,
		_w36236_
	);
	LUT2 #(
		.INIT('h8)
	) name25725 (
		_w36123_,
		_w36185_,
		_w36237_
	);
	LUT2 #(
		.INIT('h4)
	) name25726 (
		_w36111_,
		_w36237_,
		_w36238_
	);
	LUT2 #(
		.INIT('h8)
	) name25727 (
		_w36127_,
		_w36165_,
		_w36239_
	);
	LUT2 #(
		.INIT('h4)
	) name25728 (
		_w36111_,
		_w36239_,
		_w36240_
	);
	LUT2 #(
		.INIT('h8)
	) name25729 (
		_w36127_,
		_w36170_,
		_w36241_
	);
	LUT2 #(
		.INIT('h4)
	) name25730 (
		_w36111_,
		_w36241_,
		_w36242_
	);
	LUT2 #(
		.INIT('h8)
	) name25731 (
		_w36141_,
		_w36185_,
		_w36243_
	);
	LUT2 #(
		.INIT('h4)
	) name25732 (
		_w36111_,
		_w36243_,
		_w36244_
	);
	LUT2 #(
		.INIT('h8)
	) name25733 (
		_w36144_,
		_w36165_,
		_w36245_
	);
	LUT2 #(
		.INIT('h4)
	) name25734 (
		_w36111_,
		_w36245_,
		_w36246_
	);
	LUT2 #(
		.INIT('h8)
	) name25735 (
		_w36144_,
		_w36170_,
		_w36247_
	);
	LUT2 #(
		.INIT('h4)
	) name25736 (
		_w36111_,
		_w36247_,
		_w36248_
	);
	LUT2 #(
		.INIT('h8)
	) name25737 (
		_w36149_,
		_w36185_,
		_w36249_
	);
	LUT2 #(
		.INIT('h4)
	) name25738 (
		_w36111_,
		_w36249_,
		_w36250_
	);
	LUT2 #(
		.INIT('h8)
	) name25739 (
		_w36137_,
		_w36185_,
		_w36251_
	);
	LUT2 #(
		.INIT('h4)
	) name25740 (
		_w36111_,
		_w36251_,
		_w36252_
	);
	LUT2 #(
		.INIT('h4)
	) name25741 (
		_w36101_,
		_w36163_,
		_w36253_
	);
	LUT2 #(
		.INIT('h8)
	) name25742 (
		_w36104_,
		_w36212_,
		_w36254_
	);
	LUT2 #(
		.INIT('h4)
	) name25743 (
		_w36111_,
		_w36254_,
		_w36255_
	);
	LUT2 #(
		.INIT('h8)
	) name25744 (
		_w36119_,
		_w36197_,
		_w36256_
	);
	LUT2 #(
		.INIT('h4)
	) name25745 (
		_w36111_,
		_w36256_,
		_w36257_
	);
	LUT2 #(
		.INIT('h2)
	) name25746 (
		_w36115_,
		_w36133_,
		_w36258_
	);
	LUT2 #(
		.INIT('h8)
	) name25747 (
		_w36119_,
		_w36202_,
		_w36259_
	);
	LUT2 #(
		.INIT('h4)
	) name25748 (
		_w36111_,
		_w36259_,
		_w36260_
	);
	LUT2 #(
		.INIT('h2)
	) name25749 (
		_w36120_,
		_w36133_,
		_w36261_
	);
	LUT2 #(
		.INIT('h8)
	) name25750 (
		_w36119_,
		_w36207_,
		_w36262_
	);
	LUT2 #(
		.INIT('h4)
	) name25751 (
		_w36111_,
		_w36262_,
		_w36263_
	);
	LUT2 #(
		.INIT('h8)
	) name25752 (
		_w36127_,
		_w36212_,
		_w36264_
	);
	LUT2 #(
		.INIT('h4)
	) name25753 (
		_w36111_,
		_w36264_,
		_w36265_
	);
	LUT2 #(
		.INIT('h2)
	) name25754 (
		_w36125_,
		_w36133_,
		_w36266_
	);
	LUT2 #(
		.INIT('h2)
	) name25755 (
		_w36128_,
		_w36133_,
		_w36267_
	);
	LUT2 #(
		.INIT('h8)
	) name25756 (
		_w36176_,
		_w36194_,
		_w36268_
	);
	LUT2 #(
		.INIT('h4)
	) name25757 (
		_w36111_,
		_w36268_,
		_w36269_
	);
	LUT2 #(
		.INIT('h2)
	) name25758 (
		_w36130_,
		_w36133_,
		_w36270_
	);
	LUT2 #(
		.INIT('h8)
	) name25759 (
		_w36144_,
		_w36212_,
		_w36271_
	);
	LUT2 #(
		.INIT('h4)
	) name25760 (
		_w36111_,
		_w36271_,
		_w36272_
	);
	LUT2 #(
		.INIT('h4)
	) name25761 (
		_w36133_,
		_w36142_,
		_w36273_
	);
	LUT2 #(
		.INIT('h8)
	) name25762 (
		_w36113_,
		_w36155_,
		_w36274_
	);
	LUT2 #(
		.INIT('h8)
	) name25763 (
		_w36123_,
		_w36274_,
		_w36275_
	);
	LUT2 #(
		.INIT('h4)
	) name25764 (
		_w36133_,
		_w36275_,
		_w36276_
	);
	LUT2 #(
		.INIT('h4)
	) name25765 (
		_w36133_,
		_w36145_,
		_w36277_
	);
	LUT2 #(
		.INIT('h8)
	) name25766 (
		_w36113_,
		_w36134_,
		_w36278_
	);
	LUT2 #(
		.INIT('h8)
	) name25767 (
		_w36186_,
		_w36278_,
		_w36279_
	);
	LUT2 #(
		.INIT('h4)
	) name25768 (
		_w36111_,
		_w36279_,
		_w36280_
	);
	LUT2 #(
		.INIT('h4)
	) name25769 (
		_w36133_,
		_w36147_,
		_w36281_
	);
	LUT2 #(
		.INIT('h8)
	) name25770 (
		_w36135_,
		_w36186_,
		_w36282_
	);
	LUT2 #(
		.INIT('h4)
	) name25771 (
		_w36111_,
		_w36282_,
		_w36283_
	);
	LUT2 #(
		.INIT('h8)
	) name25772 (
		_w36186_,
		_w36274_,
		_w36284_
	);
	LUT2 #(
		.INIT('h4)
	) name25773 (
		_w36111_,
		_w36284_,
		_w36285_
	);
	LUT2 #(
		.INIT('h8)
	) name25774 (
		_w36189_,
		_w36194_,
		_w36286_
	);
	LUT2 #(
		.INIT('h4)
	) name25775 (
		_w36111_,
		_w36286_,
		_w36287_
	);
	LUT2 #(
		.INIT('h4)
	) name25776 (
		_w36133_,
		_w36150_,
		_w36288_
	);
	LUT2 #(
		.INIT('h4)
	) name25777 (
		_w36133_,
		_w36152_,
		_w36289_
	);
	LUT2 #(
		.INIT('h8)
	) name25778 (
		_w36117_,
		_w36158_,
		_w36290_
	);
	LUT2 #(
		.INIT('h4)
	) name25779 (
		_w36111_,
		_w36290_,
		_w36291_
	);
	LUT2 #(
		.INIT('h8)
	) name25780 (
		_w36117_,
		_w36162_,
		_w36292_
	);
	LUT2 #(
		.INIT('h4)
	) name25781 (
		_w36111_,
		_w36292_,
		_w36293_
	);
	LUT2 #(
		.INIT('h8)
	) name25782 (
		_w36107_,
		_w36166_,
		_w36294_
	);
	LUT2 #(
		.INIT('h4)
	) name25783 (
		_w36111_,
		_w36294_,
		_w36295_
	);
	LUT2 #(
		.INIT('h8)
	) name25784 (
		_w36114_,
		_w36166_,
		_w36296_
	);
	LUT2 #(
		.INIT('h4)
	) name25785 (
		_w36111_,
		_w36296_,
		_w36297_
	);
	LUT2 #(
		.INIT('h8)
	) name25786 (
		_w36117_,
		_w36173_,
		_w36298_
	);
	LUT2 #(
		.INIT('h4)
	) name25787 (
		_w36111_,
		_w36298_,
		_w36299_
	);
	LUT2 #(
		.INIT('h8)
	) name25788 (
		_w36107_,
		_w36176_,
		_w36300_
	);
	LUT2 #(
		.INIT('h4)
	) name25789 (
		_w36111_,
		_w36300_,
		_w36301_
	);
	LUT2 #(
		.INIT('h8)
	) name25790 (
		_w36114_,
		_w36176_,
		_w36302_
	);
	LUT2 #(
		.INIT('h4)
	) name25791 (
		_w36111_,
		_w36302_,
		_w36303_
	);
	LUT2 #(
		.INIT('h8)
	) name25792 (
		_w36117_,
		_w36181_,
		_w36304_
	);
	LUT2 #(
		.INIT('h4)
	) name25793 (
		_w36111_,
		_w36304_,
		_w36305_
	);
	LUT2 #(
		.INIT('h8)
	) name25794 (
		_w36124_,
		_w36186_,
		_w36306_
	);
	LUT2 #(
		.INIT('h4)
	) name25795 (
		_w36111_,
		_w36306_,
		_w36307_
	);
	LUT2 #(
		.INIT('h8)
	) name25796 (
		_w36107_,
		_w36189_,
		_w36308_
	);
	LUT2 #(
		.INIT('h4)
	) name25797 (
		_w36111_,
		_w36308_,
		_w36309_
	);
	LUT2 #(
		.INIT('h8)
	) name25798 (
		_w36114_,
		_w36189_,
		_w36310_
	);
	LUT2 #(
		.INIT('h4)
	) name25799 (
		_w36111_,
		_w36310_,
		_w36311_
	);
	LUT2 #(
		.INIT('h4)
	) name25800 (
		_w36133_,
		_w36159_,
		_w36312_
	);
	LUT2 #(
		.INIT('h4)
	) name25801 (
		_w36133_,
		_w36163_,
		_w36313_
	);
	LUT2 #(
		.INIT('h8)
	) name25802 (
		_w36104_,
		_w36194_,
		_w36314_
	);
	LUT2 #(
		.INIT('h4)
	) name25803 (
		_w36111_,
		_w36314_,
		_w36315_
	);
	LUT2 #(
		.INIT('h4)
	) name25804 (
		_w36133_,
		_w36167_,
		_w36316_
	);
	LUT2 #(
		.INIT('h8)
	) name25805 (
		_w36123_,
		_w36278_,
		_w36317_
	);
	LUT2 #(
		.INIT('h4)
	) name25806 (
		_w36111_,
		_w36317_,
		_w36318_
	);
	LUT2 #(
		.INIT('h8)
	) name25807 (
		_w36123_,
		_w36135_,
		_w36319_
	);
	LUT2 #(
		.INIT('h4)
	) name25808 (
		_w36111_,
		_w36319_,
		_w36320_
	);
	LUT2 #(
		.INIT('h4)
	) name25809 (
		_w36111_,
		_w36275_,
		_w36321_
	);
	LUT2 #(
		.INIT('h8)
	) name25810 (
		_w36127_,
		_w36194_,
		_w36322_
	);
	LUT2 #(
		.INIT('h4)
	) name25811 (
		_w36111_,
		_w36322_,
		_w36323_
	);
	LUT2 #(
		.INIT('h4)
	) name25812 (
		_w36133_,
		_w36171_,
		_w36324_
	);
	LUT2 #(
		.INIT('h4)
	) name25813 (
		_w36133_,
		_w36174_,
		_w36325_
	);
	LUT2 #(
		.INIT('h8)
	) name25814 (
		_w36141_,
		_w36278_,
		_w36326_
	);
	LUT2 #(
		.INIT('h4)
	) name25815 (
		_w36111_,
		_w36326_,
		_w36327_
	);
	LUT2 #(
		.INIT('h8)
	) name25816 (
		_w36135_,
		_w36141_,
		_w36328_
	);
	LUT2 #(
		.INIT('h4)
	) name25817 (
		_w36111_,
		_w36328_,
		_w36329_
	);
	LUT2 #(
		.INIT('h8)
	) name25818 (
		_w36141_,
		_w36274_,
		_w36330_
	);
	LUT2 #(
		.INIT('h4)
	) name25819 (
		_w36111_,
		_w36330_,
		_w36331_
	);
	LUT2 #(
		.INIT('h8)
	) name25820 (
		_w36144_,
		_w36194_,
		_w36332_
	);
	LUT2 #(
		.INIT('h4)
	) name25821 (
		_w36111_,
		_w36332_,
		_w36333_
	);
	LUT2 #(
		.INIT('h8)
	) name25822 (
		_w36149_,
		_w36278_,
		_w36334_
	);
	LUT2 #(
		.INIT('h4)
	) name25823 (
		_w36111_,
		_w36334_,
		_w36335_
	);
	LUT2 #(
		.INIT('h8)
	) name25824 (
		_w36137_,
		_w36278_,
		_w36336_
	);
	LUT2 #(
		.INIT('h4)
	) name25825 (
		_w36111_,
		_w36336_,
		_w36337_
	);
	LUT2 #(
		.INIT('h4)
	) name25826 (
		_w36133_,
		_w36177_,
		_w36338_
	);
	LUT2 #(
		.INIT('h8)
	) name25827 (
		_w36135_,
		_w36149_,
		_w36339_
	);
	LUT2 #(
		.INIT('h4)
	) name25828 (
		_w36111_,
		_w36339_,
		_w36340_
	);
	LUT2 #(
		.INIT('h4)
	) name25829 (
		_w36111_,
		_w36138_,
		_w36341_
	);
	LUT2 #(
		.INIT('h8)
	) name25830 (
		_w36149_,
		_w36274_,
		_w36342_
	);
	LUT2 #(
		.INIT('h4)
	) name25831 (
		_w36111_,
		_w36342_,
		_w36343_
	);
	LUT2 #(
		.INIT('h4)
	) name25832 (
		_w36133_,
		_w36179_,
		_w36344_
	);
	LUT2 #(
		.INIT('h8)
	) name25833 (
		_w36137_,
		_w36274_,
		_w36345_
	);
	LUT2 #(
		.INIT('h4)
	) name25834 (
		_w36111_,
		_w36345_,
		_w36346_
	);
	LUT2 #(
		.INIT('h4)
	) name25835 (
		_w36133_,
		_w36182_,
		_w36347_
	);
	LUT2 #(
		.INIT('h2)
	) name25836 (
		_w36108_,
		_w36111_,
		_w36348_
	);
	LUT2 #(
		.INIT('h4)
	) name25837 (
		_w36133_,
		_w36187_,
		_w36349_
	);
	LUT2 #(
		.INIT('h8)
	) name25838 (
		\wishbone_BDWrite_reg[3]/NET0131 ,
		_w36098_,
		_w36350_
	);
	LUT2 #(
		.INIT('h2)
	) name25839 (
		_w36100_,
		_w36350_,
		_w36351_
	);
	LUT2 #(
		.INIT('h2)
	) name25840 (
		_w36115_,
		_w36351_,
		_w36352_
	);
	LUT2 #(
		.INIT('h2)
	) name25841 (
		_w36120_,
		_w36351_,
		_w36353_
	);
	LUT2 #(
		.INIT('h4)
	) name25842 (
		_w36133_,
		_w36190_,
		_w36354_
	);
	LUT2 #(
		.INIT('h2)
	) name25843 (
		_w36125_,
		_w36351_,
		_w36355_
	);
	LUT2 #(
		.INIT('h2)
	) name25844 (
		_w36128_,
		_w36351_,
		_w36356_
	);
	LUT2 #(
		.INIT('h4)
	) name25845 (
		_w36133_,
		_w36192_,
		_w36357_
	);
	LUT2 #(
		.INIT('h2)
	) name25846 (
		_w36130_,
		_w36351_,
		_w36358_
	);
	LUT2 #(
		.INIT('h2)
	) name25847 (
		_w36142_,
		_w36351_,
		_w36359_
	);
	LUT2 #(
		.INIT('h4)
	) name25848 (
		_w36133_,
		_w36195_,
		_w36360_
	);
	LUT2 #(
		.INIT('h2)
	) name25849 (
		_w36145_,
		_w36351_,
		_w36361_
	);
	LUT2 #(
		.INIT('h2)
	) name25850 (
		_w36147_,
		_w36351_,
		_w36362_
	);
	LUT2 #(
		.INIT('h4)
	) name25851 (
		_w36133_,
		_w36198_,
		_w36363_
	);
	LUT2 #(
		.INIT('h2)
	) name25852 (
		_w36150_,
		_w36351_,
		_w36364_
	);
	LUT2 #(
		.INIT('h2)
	) name25853 (
		_w36152_,
		_w36351_,
		_w36365_
	);
	LUT2 #(
		.INIT('h4)
	) name25854 (
		_w36133_,
		_w36200_,
		_w36366_
	);
	LUT2 #(
		.INIT('h4)
	) name25855 (
		_w36133_,
		_w36203_,
		_w36367_
	);
	LUT2 #(
		.INIT('h4)
	) name25856 (
		_w36133_,
		_w36205_,
		_w36368_
	);
	LUT2 #(
		.INIT('h4)
	) name25857 (
		_w36133_,
		_w36208_,
		_w36369_
	);
	LUT2 #(
		.INIT('h4)
	) name25858 (
		_w36133_,
		_w36210_,
		_w36370_
	);
	LUT2 #(
		.INIT('h4)
	) name25859 (
		_w36133_,
		_w36213_,
		_w36371_
	);
	LUT2 #(
		.INIT('h2)
	) name25860 (
		_w36159_,
		_w36351_,
		_w36372_
	);
	LUT2 #(
		.INIT('h2)
	) name25861 (
		_w36163_,
		_w36351_,
		_w36373_
	);
	LUT2 #(
		.INIT('h4)
	) name25862 (
		_w36133_,
		_w36215_,
		_w36374_
	);
	LUT2 #(
		.INIT('h2)
	) name25863 (
		_w36167_,
		_w36351_,
		_w36375_
	);
	LUT2 #(
		.INIT('h4)
	) name25864 (
		_w36133_,
		_w36217_,
		_w36376_
	);
	LUT2 #(
		.INIT('h2)
	) name25865 (
		_w36171_,
		_w36351_,
		_w36377_
	);
	LUT2 #(
		.INIT('h2)
	) name25866 (
		_w36174_,
		_w36351_,
		_w36378_
	);
	LUT2 #(
		.INIT('h4)
	) name25867 (
		_w36133_,
		_w36219_,
		_w36379_
	);
	LUT2 #(
		.INIT('h2)
	) name25868 (
		_w36177_,
		_w36351_,
		_w36380_
	);
	LUT2 #(
		.INIT('h2)
	) name25869 (
		_w36179_,
		_w36351_,
		_w36381_
	);
	LUT2 #(
		.INIT('h4)
	) name25870 (
		_w36133_,
		_w36221_,
		_w36382_
	);
	LUT2 #(
		.INIT('h2)
	) name25871 (
		_w36182_,
		_w36351_,
		_w36383_
	);
	LUT2 #(
		.INIT('h4)
	) name25872 (
		_w36133_,
		_w36223_,
		_w36384_
	);
	LUT2 #(
		.INIT('h2)
	) name25873 (
		_w36187_,
		_w36351_,
		_w36385_
	);
	LUT2 #(
		.INIT('h2)
	) name25874 (
		_w36190_,
		_w36351_,
		_w36386_
	);
	LUT2 #(
		.INIT('h2)
	) name25875 (
		_w36192_,
		_w36351_,
		_w36387_
	);
	LUT2 #(
		.INIT('h4)
	) name25876 (
		_w36133_,
		_w36225_,
		_w36388_
	);
	LUT2 #(
		.INIT('h2)
	) name25877 (
		_w36195_,
		_w36351_,
		_w36389_
	);
	LUT2 #(
		.INIT('h4)
	) name25878 (
		_w36133_,
		_w36227_,
		_w36390_
	);
	LUT2 #(
		.INIT('h2)
	) name25879 (
		_w36198_,
		_w36351_,
		_w36391_
	);
	LUT2 #(
		.INIT('h2)
	) name25880 (
		_w36200_,
		_w36351_,
		_w36392_
	);
	LUT2 #(
		.INIT('h2)
	) name25881 (
		_w36203_,
		_w36351_,
		_w36393_
	);
	LUT2 #(
		.INIT('h4)
	) name25882 (
		_w36133_,
		_w36229_,
		_w36394_
	);
	LUT2 #(
		.INIT('h2)
	) name25883 (
		_w36205_,
		_w36351_,
		_w36395_
	);
	LUT2 #(
		.INIT('h2)
	) name25884 (
		_w36208_,
		_w36351_,
		_w36396_
	);
	LUT2 #(
		.INIT('h2)
	) name25885 (
		_w36210_,
		_w36351_,
		_w36397_
	);
	LUT2 #(
		.INIT('h2)
	) name25886 (
		_w36213_,
		_w36351_,
		_w36398_
	);
	LUT2 #(
		.INIT('h2)
	) name25887 (
		_w36215_,
		_w36351_,
		_w36399_
	);
	LUT2 #(
		.INIT('h2)
	) name25888 (
		_w36217_,
		_w36351_,
		_w36400_
	);
	LUT2 #(
		.INIT('h2)
	) name25889 (
		_w36219_,
		_w36351_,
		_w36401_
	);
	LUT2 #(
		.INIT('h2)
	) name25890 (
		_w36221_,
		_w36351_,
		_w36402_
	);
	LUT2 #(
		.INIT('h2)
	) name25891 (
		_w36223_,
		_w36351_,
		_w36403_
	);
	LUT2 #(
		.INIT('h2)
	) name25892 (
		_w36225_,
		_w36351_,
		_w36404_
	);
	LUT2 #(
		.INIT('h2)
	) name25893 (
		_w36227_,
		_w36351_,
		_w36405_
	);
	LUT2 #(
		.INIT('h2)
	) name25894 (
		_w36229_,
		_w36351_,
		_w36406_
	);
	LUT2 #(
		.INIT('h4)
	) name25895 (
		_w36133_,
		_w36231_,
		_w36407_
	);
	LUT2 #(
		.INIT('h4)
	) name25896 (
		_w36133_,
		_w36233_,
		_w36408_
	);
	LUT2 #(
		.INIT('h4)
	) name25897 (
		_w36133_,
		_w36235_,
		_w36409_
	);
	LUT2 #(
		.INIT('h2)
	) name25898 (
		_w36231_,
		_w36351_,
		_w36410_
	);
	LUT2 #(
		.INIT('h2)
	) name25899 (
		_w36233_,
		_w36351_,
		_w36411_
	);
	LUT2 #(
		.INIT('h2)
	) name25900 (
		_w36235_,
		_w36351_,
		_w36412_
	);
	LUT2 #(
		.INIT('h4)
	) name25901 (
		_w36133_,
		_w36237_,
		_w36413_
	);
	LUT2 #(
		.INIT('h2)
	) name25902 (
		_w36237_,
		_w36351_,
		_w36414_
	);
	LUT2 #(
		.INIT('h4)
	) name25903 (
		_w36133_,
		_w36239_,
		_w36415_
	);
	LUT2 #(
		.INIT('h2)
	) name25904 (
		_w36239_,
		_w36351_,
		_w36416_
	);
	LUT2 #(
		.INIT('h2)
	) name25905 (
		_w36241_,
		_w36351_,
		_w36417_
	);
	LUT2 #(
		.INIT('h4)
	) name25906 (
		_w36133_,
		_w36241_,
		_w36418_
	);
	LUT2 #(
		.INIT('h2)
	) name25907 (
		_w36243_,
		_w36351_,
		_w36419_
	);
	LUT2 #(
		.INIT('h2)
	) name25908 (
		_w36245_,
		_w36351_,
		_w36420_
	);
	LUT2 #(
		.INIT('h2)
	) name25909 (
		_w36247_,
		_w36351_,
		_w36421_
	);
	LUT2 #(
		.INIT('h4)
	) name25910 (
		_w36133_,
		_w36243_,
		_w36422_
	);
	LUT2 #(
		.INIT('h2)
	) name25911 (
		_w36249_,
		_w36351_,
		_w36423_
	);
	LUT2 #(
		.INIT('h2)
	) name25912 (
		_w36251_,
		_w36351_,
		_w36424_
	);
	LUT2 #(
		.INIT('h4)
	) name25913 (
		_w36133_,
		_w36245_,
		_w36425_
	);
	LUT2 #(
		.INIT('h4)
	) name25914 (
		_w36133_,
		_w36247_,
		_w36426_
	);
	LUT2 #(
		.INIT('h2)
	) name25915 (
		_w36254_,
		_w36351_,
		_w36427_
	);
	LUT2 #(
		.INIT('h2)
	) name25916 (
		_w36256_,
		_w36351_,
		_w36428_
	);
	LUT2 #(
		.INIT('h2)
	) name25917 (
		_w36259_,
		_w36351_,
		_w36429_
	);
	LUT2 #(
		.INIT('h4)
	) name25918 (
		_w36133_,
		_w36249_,
		_w36430_
	);
	LUT2 #(
		.INIT('h2)
	) name25919 (
		_w36262_,
		_w36351_,
		_w36431_
	);
	LUT2 #(
		.INIT('h4)
	) name25920 (
		_w36133_,
		_w36251_,
		_w36432_
	);
	LUT2 #(
		.INIT('h2)
	) name25921 (
		_w36264_,
		_w36351_,
		_w36433_
	);
	LUT2 #(
		.INIT('h2)
	) name25922 (
		_w36268_,
		_w36351_,
		_w36434_
	);
	LUT2 #(
		.INIT('h2)
	) name25923 (
		_w36271_,
		_w36351_,
		_w36435_
	);
	LUT2 #(
		.INIT('h4)
	) name25924 (
		_w36133_,
		_w36254_,
		_w36436_
	);
	LUT2 #(
		.INIT('h4)
	) name25925 (
		_w36133_,
		_w36256_,
		_w36437_
	);
	LUT2 #(
		.INIT('h4)
	) name25926 (
		_w36133_,
		_w36259_,
		_w36438_
	);
	LUT2 #(
		.INIT('h2)
	) name25927 (
		_w36279_,
		_w36351_,
		_w36439_
	);
	LUT2 #(
		.INIT('h2)
	) name25928 (
		_w36282_,
		_w36351_,
		_w36440_
	);
	LUT2 #(
		.INIT('h4)
	) name25929 (
		_w36133_,
		_w36262_,
		_w36441_
	);
	LUT2 #(
		.INIT('h2)
	) name25930 (
		_w36284_,
		_w36351_,
		_w36442_
	);
	LUT2 #(
		.INIT('h2)
	) name25931 (
		_w36286_,
		_w36351_,
		_w36443_
	);
	LUT2 #(
		.INIT('h4)
	) name25932 (
		_w36133_,
		_w36264_,
		_w36444_
	);
	LUT2 #(
		.INIT('h2)
	) name25933 (
		_w36290_,
		_w36351_,
		_w36445_
	);
	LUT2 #(
		.INIT('h2)
	) name25934 (
		_w36292_,
		_w36351_,
		_w36446_
	);
	LUT2 #(
		.INIT('h2)
	) name25935 (
		_w36294_,
		_w36351_,
		_w36447_
	);
	LUT2 #(
		.INIT('h2)
	) name25936 (
		_w36296_,
		_w36351_,
		_w36448_
	);
	LUT2 #(
		.INIT('h2)
	) name25937 (
		_w36298_,
		_w36351_,
		_w36449_
	);
	LUT2 #(
		.INIT('h4)
	) name25938 (
		_w36133_,
		_w36268_,
		_w36450_
	);
	LUT2 #(
		.INIT('h4)
	) name25939 (
		_w36133_,
		_w36271_,
		_w36451_
	);
	LUT2 #(
		.INIT('h2)
	) name25940 (
		_w36300_,
		_w36351_,
		_w36452_
	);
	LUT2 #(
		.INIT('h2)
	) name25941 (
		_w36302_,
		_w36351_,
		_w36453_
	);
	LUT2 #(
		.INIT('h2)
	) name25942 (
		_w36304_,
		_w36351_,
		_w36454_
	);
	LUT2 #(
		.INIT('h2)
	) name25943 (
		_w36306_,
		_w36351_,
		_w36455_
	);
	LUT2 #(
		.INIT('h2)
	) name25944 (
		_w36308_,
		_w36351_,
		_w36456_
	);
	LUT2 #(
		.INIT('h2)
	) name25945 (
		_w36310_,
		_w36351_,
		_w36457_
	);
	LUT2 #(
		.INIT('h2)
	) name25946 (
		_w36314_,
		_w36351_,
		_w36458_
	);
	LUT2 #(
		.INIT('h2)
	) name25947 (
		_w36317_,
		_w36351_,
		_w36459_
	);
	LUT2 #(
		.INIT('h2)
	) name25948 (
		_w36319_,
		_w36351_,
		_w36460_
	);
	LUT2 #(
		.INIT('h2)
	) name25949 (
		_w36275_,
		_w36351_,
		_w36461_
	);
	LUT2 #(
		.INIT('h2)
	) name25950 (
		_w36322_,
		_w36351_,
		_w36462_
	);
	LUT2 #(
		.INIT('h4)
	) name25951 (
		_w36133_,
		_w36279_,
		_w36463_
	);
	LUT2 #(
		.INIT('h2)
	) name25952 (
		_w36326_,
		_w36351_,
		_w36464_
	);
	LUT2 #(
		.INIT('h2)
	) name25953 (
		_w36328_,
		_w36351_,
		_w36465_
	);
	LUT2 #(
		.INIT('h4)
	) name25954 (
		_w36133_,
		_w36282_,
		_w36466_
	);
	LUT2 #(
		.INIT('h2)
	) name25955 (
		_w36330_,
		_w36351_,
		_w36467_
	);
	LUT2 #(
		.INIT('h2)
	) name25956 (
		_w36332_,
		_w36351_,
		_w36468_
	);
	LUT2 #(
		.INIT('h2)
	) name25957 (
		_w36334_,
		_w36351_,
		_w36469_
	);
	LUT2 #(
		.INIT('h4)
	) name25958 (
		_w36133_,
		_w36284_,
		_w36470_
	);
	LUT2 #(
		.INIT('h2)
	) name25959 (
		_w36336_,
		_w36351_,
		_w36471_
	);
	LUT2 #(
		.INIT('h2)
	) name25960 (
		_w36339_,
		_w36351_,
		_w36472_
	);
	LUT2 #(
		.INIT('h2)
	) name25961 (
		_w36138_,
		_w36351_,
		_w36473_
	);
	LUT2 #(
		.INIT('h4)
	) name25962 (
		_w36133_,
		_w36286_,
		_w36474_
	);
	LUT2 #(
		.INIT('h2)
	) name25963 (
		_w36342_,
		_w36351_,
		_w36475_
	);
	LUT2 #(
		.INIT('h2)
	) name25964 (
		_w36345_,
		_w36351_,
		_w36476_
	);
	LUT2 #(
		.INIT('h2)
	) name25965 (
		_w36108_,
		_w36351_,
		_w36477_
	);
	LUT2 #(
		.INIT('h4)
	) name25966 (
		_w36133_,
		_w36290_,
		_w36478_
	);
	LUT2 #(
		.INIT('h4)
	) name25967 (
		_w36133_,
		_w36292_,
		_w36479_
	);
	LUT2 #(
		.INIT('h4)
	) name25968 (
		_w36133_,
		_w36330_,
		_w36480_
	);
	LUT2 #(
		.INIT('h4)
	) name25969 (
		_w36133_,
		_w36294_,
		_w36481_
	);
	LUT2 #(
		.INIT('h4)
	) name25970 (
		_w36133_,
		_w36296_,
		_w36482_
	);
	LUT2 #(
		.INIT('h4)
	) name25971 (
		_w36133_,
		_w36298_,
		_w36483_
	);
	LUT2 #(
		.INIT('h4)
	) name25972 (
		_w36101_,
		_w36152_,
		_w36484_
	);
	LUT2 #(
		.INIT('h4)
	) name25973 (
		_w36133_,
		_w36300_,
		_w36485_
	);
	LUT2 #(
		.INIT('h4)
	) name25974 (
		_w36133_,
		_w36302_,
		_w36486_
	);
	LUT2 #(
		.INIT('h4)
	) name25975 (
		_w36133_,
		_w36304_,
		_w36487_
	);
	LUT2 #(
		.INIT('h4)
	) name25976 (
		_w36133_,
		_w36306_,
		_w36488_
	);
	LUT2 #(
		.INIT('h4)
	) name25977 (
		_w36133_,
		_w36308_,
		_w36489_
	);
	LUT2 #(
		.INIT('h4)
	) name25978 (
		_w36133_,
		_w36310_,
		_w36490_
	);
	LUT2 #(
		.INIT('h4)
	) name25979 (
		_w36133_,
		_w36314_,
		_w36491_
	);
	LUT2 #(
		.INIT('h4)
	) name25980 (
		_w36133_,
		_w36317_,
		_w36492_
	);
	LUT2 #(
		.INIT('h4)
	) name25981 (
		_w36133_,
		_w36342_,
		_w36493_
	);
	LUT2 #(
		.INIT('h4)
	) name25982 (
		_w36133_,
		_w36319_,
		_w36494_
	);
	LUT2 #(
		.INIT('h4)
	) name25983 (
		_w36133_,
		_w36322_,
		_w36495_
	);
	LUT2 #(
		.INIT('h4)
	) name25984 (
		_w36133_,
		_w36326_,
		_w36496_
	);
	LUT2 #(
		.INIT('h4)
	) name25985 (
		_w36133_,
		_w36328_,
		_w36497_
	);
	LUT2 #(
		.INIT('h4)
	) name25986 (
		_w36133_,
		_w36332_,
		_w36498_
	);
	LUT2 #(
		.INIT('h4)
	) name25987 (
		_w36133_,
		_w36334_,
		_w36499_
	);
	LUT2 #(
		.INIT('h4)
	) name25988 (
		_w36133_,
		_w36336_,
		_w36500_
	);
	LUT2 #(
		.INIT('h4)
	) name25989 (
		_w36133_,
		_w36339_,
		_w36501_
	);
	LUT2 #(
		.INIT('h4)
	) name25990 (
		_w36133_,
		_w36345_,
		_w36502_
	);
	LUT2 #(
		.INIT('h2)
	) name25991 (
		_w36108_,
		_w36133_,
		_w36503_
	);
	LUT2 #(
		.INIT('h4)
	) name25992 (
		_w36101_,
		_w36115_,
		_w36504_
	);
	LUT2 #(
		.INIT('h4)
	) name25993 (
		_w36101_,
		_w36120_,
		_w36505_
	);
	LUT2 #(
		.INIT('h4)
	) name25994 (
		_w36101_,
		_w36125_,
		_w36506_
	);
	LUT2 #(
		.INIT('h4)
	) name25995 (
		_w36101_,
		_w36128_,
		_w36507_
	);
	LUT2 #(
		.INIT('h4)
	) name25996 (
		_w36101_,
		_w36130_,
		_w36508_
	);
	LUT2 #(
		.INIT('h4)
	) name25997 (
		_w36101_,
		_w36150_,
		_w36509_
	);
	LUT2 #(
		.INIT('h4)
	) name25998 (
		_w36101_,
		_w36142_,
		_w36510_
	);
	LUT2 #(
		.INIT('h4)
	) name25999 (
		_w36101_,
		_w36145_,
		_w36511_
	);
	LUT2 #(
		.INIT('h4)
	) name26000 (
		_w36101_,
		_w36147_,
		_w36512_
	);
	LUT2 #(
		.INIT('h4)
	) name26001 (
		_w36101_,
		_w36167_,
		_w36513_
	);
	LUT2 #(
		.INIT('h4)
	) name26002 (
		_w36101_,
		_w36171_,
		_w36514_
	);
	LUT2 #(
		.INIT('h4)
	) name26003 (
		_w36101_,
		_w36174_,
		_w36515_
	);
	LUT2 #(
		.INIT('h4)
	) name26004 (
		_w36101_,
		_w36177_,
		_w36516_
	);
	LUT2 #(
		.INIT('h4)
	) name26005 (
		_w36101_,
		_w36179_,
		_w36517_
	);
	LUT2 #(
		.INIT('h4)
	) name26006 (
		_w36101_,
		_w36182_,
		_w36518_
	);
	LUT2 #(
		.INIT('h4)
	) name26007 (
		_w36101_,
		_w36187_,
		_w36519_
	);
	LUT2 #(
		.INIT('h4)
	) name26008 (
		_w36101_,
		_w36190_,
		_w36520_
	);
	LUT2 #(
		.INIT('h4)
	) name26009 (
		_w36101_,
		_w36192_,
		_w36521_
	);
	LUT2 #(
		.INIT('h4)
	) name26010 (
		_w36101_,
		_w36195_,
		_w36522_
	);
	LUT2 #(
		.INIT('h4)
	) name26011 (
		_w36101_,
		_w36198_,
		_w36523_
	);
	LUT2 #(
		.INIT('h4)
	) name26012 (
		_w36101_,
		_w36200_,
		_w36524_
	);
	LUT2 #(
		.INIT('h4)
	) name26013 (
		_w36101_,
		_w36203_,
		_w36525_
	);
	LUT2 #(
		.INIT('h4)
	) name26014 (
		_w36101_,
		_w36205_,
		_w36526_
	);
	LUT2 #(
		.INIT('h4)
	) name26015 (
		_w36101_,
		_w36208_,
		_w36527_
	);
	LUT2 #(
		.INIT('h4)
	) name26016 (
		_w36101_,
		_w36210_,
		_w36528_
	);
	LUT2 #(
		.INIT('h4)
	) name26017 (
		_w36101_,
		_w36213_,
		_w36529_
	);
	LUT2 #(
		.INIT('h4)
	) name26018 (
		_w36101_,
		_w36215_,
		_w36530_
	);
	LUT2 #(
		.INIT('h4)
	) name26019 (
		_w36101_,
		_w36217_,
		_w36531_
	);
	LUT2 #(
		.INIT('h4)
	) name26020 (
		_w36101_,
		_w36219_,
		_w36532_
	);
	LUT2 #(
		.INIT('h4)
	) name26021 (
		_w36101_,
		_w36221_,
		_w36533_
	);
	LUT2 #(
		.INIT('h4)
	) name26022 (
		_w36101_,
		_w36223_,
		_w36534_
	);
	LUT2 #(
		.INIT('h4)
	) name26023 (
		_w36101_,
		_w36225_,
		_w36535_
	);
	LUT2 #(
		.INIT('h4)
	) name26024 (
		_w36101_,
		_w36227_,
		_w36536_
	);
	LUT2 #(
		.INIT('h4)
	) name26025 (
		_w36101_,
		_w36229_,
		_w36537_
	);
	LUT2 #(
		.INIT('h4)
	) name26026 (
		_w36101_,
		_w36231_,
		_w36538_
	);
	LUT2 #(
		.INIT('h4)
	) name26027 (
		_w36101_,
		_w36233_,
		_w36539_
	);
	LUT2 #(
		.INIT('h4)
	) name26028 (
		_w36101_,
		_w36235_,
		_w36540_
	);
	LUT2 #(
		.INIT('h4)
	) name26029 (
		_w36101_,
		_w36237_,
		_w36541_
	);
	LUT2 #(
		.INIT('h4)
	) name26030 (
		_w36101_,
		_w36239_,
		_w36542_
	);
	LUT2 #(
		.INIT('h4)
	) name26031 (
		_w36101_,
		_w36241_,
		_w36543_
	);
	LUT2 #(
		.INIT('h4)
	) name26032 (
		_w36101_,
		_w36243_,
		_w36544_
	);
	LUT2 #(
		.INIT('h4)
	) name26033 (
		_w36101_,
		_w36245_,
		_w36545_
	);
	LUT2 #(
		.INIT('h4)
	) name26034 (
		_w36101_,
		_w36247_,
		_w36546_
	);
	LUT2 #(
		.INIT('h4)
	) name26035 (
		_w36101_,
		_w36249_,
		_w36547_
	);
	LUT2 #(
		.INIT('h4)
	) name26036 (
		_w36101_,
		_w36251_,
		_w36548_
	);
	LUT2 #(
		.INIT('h4)
	) name26037 (
		_w36101_,
		_w36254_,
		_w36549_
	);
	LUT2 #(
		.INIT('h4)
	) name26038 (
		_w36101_,
		_w36256_,
		_w36550_
	);
	LUT2 #(
		.INIT('h4)
	) name26039 (
		_w36101_,
		_w36259_,
		_w36551_
	);
	LUT2 #(
		.INIT('h4)
	) name26040 (
		_w36101_,
		_w36262_,
		_w36552_
	);
	LUT2 #(
		.INIT('h4)
	) name26041 (
		_w36101_,
		_w36264_,
		_w36553_
	);
	LUT2 #(
		.INIT('h4)
	) name26042 (
		_w36101_,
		_w36268_,
		_w36554_
	);
	LUT2 #(
		.INIT('h4)
	) name26043 (
		_w36101_,
		_w36271_,
		_w36555_
	);
	LUT2 #(
		.INIT('h4)
	) name26044 (
		_w36101_,
		_w36279_,
		_w36556_
	);
	LUT2 #(
		.INIT('h4)
	) name26045 (
		_w36101_,
		_w36282_,
		_w36557_
	);
	LUT2 #(
		.INIT('h4)
	) name26046 (
		_w36101_,
		_w36284_,
		_w36558_
	);
	LUT2 #(
		.INIT('h4)
	) name26047 (
		_w36101_,
		_w36286_,
		_w36559_
	);
	LUT2 #(
		.INIT('h4)
	) name26048 (
		_w36101_,
		_w36290_,
		_w36560_
	);
	LUT2 #(
		.INIT('h4)
	) name26049 (
		_w36101_,
		_w36292_,
		_w36561_
	);
	LUT2 #(
		.INIT('h4)
	) name26050 (
		_w36101_,
		_w36294_,
		_w36562_
	);
	LUT2 #(
		.INIT('h4)
	) name26051 (
		_w36101_,
		_w36296_,
		_w36563_
	);
	LUT2 #(
		.INIT('h4)
	) name26052 (
		_w36101_,
		_w36298_,
		_w36564_
	);
	LUT2 #(
		.INIT('h4)
	) name26053 (
		_w36101_,
		_w36300_,
		_w36565_
	);
	LUT2 #(
		.INIT('h4)
	) name26054 (
		_w36101_,
		_w36302_,
		_w36566_
	);
	LUT2 #(
		.INIT('h4)
	) name26055 (
		_w36101_,
		_w36304_,
		_w36567_
	);
	LUT2 #(
		.INIT('h4)
	) name26056 (
		_w36101_,
		_w36306_,
		_w36568_
	);
	LUT2 #(
		.INIT('h4)
	) name26057 (
		_w36101_,
		_w36308_,
		_w36569_
	);
	LUT2 #(
		.INIT('h4)
	) name26058 (
		_w36101_,
		_w36310_,
		_w36570_
	);
	LUT2 #(
		.INIT('h4)
	) name26059 (
		_w36101_,
		_w36314_,
		_w36571_
	);
	LUT2 #(
		.INIT('h4)
	) name26060 (
		_w36101_,
		_w36317_,
		_w36572_
	);
	LUT2 #(
		.INIT('h4)
	) name26061 (
		_w36101_,
		_w36319_,
		_w36573_
	);
	LUT2 #(
		.INIT('h4)
	) name26062 (
		_w36101_,
		_w36275_,
		_w36574_
	);
	LUT2 #(
		.INIT('h4)
	) name26063 (
		_w36101_,
		_w36322_,
		_w36575_
	);
	LUT2 #(
		.INIT('h4)
	) name26064 (
		_w36101_,
		_w36326_,
		_w36576_
	);
	LUT2 #(
		.INIT('h4)
	) name26065 (
		_w36101_,
		_w36328_,
		_w36577_
	);
	LUT2 #(
		.INIT('h4)
	) name26066 (
		_w36101_,
		_w36330_,
		_w36578_
	);
	LUT2 #(
		.INIT('h4)
	) name26067 (
		_w36101_,
		_w36332_,
		_w36579_
	);
	LUT2 #(
		.INIT('h4)
	) name26068 (
		_w36101_,
		_w36334_,
		_w36580_
	);
	LUT2 #(
		.INIT('h4)
	) name26069 (
		_w36101_,
		_w36336_,
		_w36581_
	);
	LUT2 #(
		.INIT('h4)
	) name26070 (
		_w36101_,
		_w36339_,
		_w36582_
	);
	LUT2 #(
		.INIT('h4)
	) name26071 (
		_w36101_,
		_w36138_,
		_w36583_
	);
	LUT2 #(
		.INIT('h4)
	) name26072 (
		_w36101_,
		_w36342_,
		_w36584_
	);
	LUT2 #(
		.INIT('h4)
	) name26073 (
		_w36101_,
		_w36345_,
		_w36585_
	);
	LUT2 #(
		.INIT('h8)
	) name26074 (
		_w36166_,
		_w36278_,
		_w36586_
	);
	LUT2 #(
		.INIT('h4)
	) name26075 (
		_w36101_,
		_w36586_,
		_w36587_
	);
	LUT2 #(
		.INIT('h8)
	) name26076 (
		_w36107_,
		_w36141_,
		_w36588_
	);
	LUT2 #(
		.INIT('h4)
	) name26077 (
		_w36101_,
		_w36588_,
		_w36589_
	);
	LUT2 #(
		.INIT('h8)
	) name26078 (
		_w36158_,
		_w36278_,
		_w36590_
	);
	LUT2 #(
		.INIT('h4)
	) name26079 (
		_w36111_,
		_w36590_,
		_w36591_
	);
	LUT2 #(
		.INIT('h8)
	) name26080 (
		_w36114_,
		_w36119_,
		_w36592_
	);
	LUT2 #(
		.INIT('h4)
	) name26081 (
		_w36111_,
		_w36592_,
		_w36593_
	);
	LUT2 #(
		.INIT('h8)
	) name26082 (
		_w36104_,
		_w36117_,
		_w36594_
	);
	LUT2 #(
		.INIT('h4)
	) name26083 (
		_w36111_,
		_w36594_,
		_w36595_
	);
	LUT2 #(
		.INIT('h8)
	) name26084 (
		_w36124_,
		_w36127_,
		_w36596_
	);
	LUT2 #(
		.INIT('h4)
	) name26085 (
		_w36111_,
		_w36596_,
		_w36597_
	);
	LUT2 #(
		.INIT('h8)
	) name26086 (
		_w36107_,
		_w36123_,
		_w36598_
	);
	LUT2 #(
		.INIT('h4)
	) name26087 (
		_w36111_,
		_w36598_,
		_w36599_
	);
	LUT2 #(
		.INIT('h8)
	) name26088 (
		_w36114_,
		_w36123_,
		_w36600_
	);
	LUT2 #(
		.INIT('h4)
	) name26089 (
		_w36111_,
		_w36600_,
		_w36601_
	);
	LUT2 #(
		.INIT('h8)
	) name26090 (
		_w36135_,
		_w36173_,
		_w36602_
	);
	LUT2 #(
		.INIT('h4)
	) name26091 (
		_w36111_,
		_w36602_,
		_w36603_
	);
	LUT2 #(
		.INIT('h8)
	) name26092 (
		_w36117_,
		_w36127_,
		_w36604_
	);
	LUT2 #(
		.INIT('h4)
	) name26093 (
		_w36111_,
		_w36604_,
		_w36605_
	);
	LUT2 #(
		.INIT('h8)
	) name26094 (
		_w36117_,
		_w36123_,
		_w36606_
	);
	LUT2 #(
		.INIT('h4)
	) name26095 (
		_w36111_,
		_w36606_,
		_w36607_
	);
	LUT2 #(
		.INIT('h8)
	) name26096 (
		_w36124_,
		_w36144_,
		_w36608_
	);
	LUT2 #(
		.INIT('h4)
	) name26097 (
		_w36111_,
		_w36608_,
		_w36609_
	);
	LUT2 #(
		.INIT('h4)
	) name26098 (
		_w36111_,
		_w36588_,
		_w36610_
	);
	LUT2 #(
		.INIT('h8)
	) name26099 (
		_w36114_,
		_w36141_,
		_w36611_
	);
	LUT2 #(
		.INIT('h4)
	) name26100 (
		_w36111_,
		_w36611_,
		_w36612_
	);
	LUT2 #(
		.INIT('h8)
	) name26101 (
		_w36117_,
		_w36144_,
		_w36613_
	);
	LUT2 #(
		.INIT('h4)
	) name26102 (
		_w36111_,
		_w36613_,
		_w36614_
	);
	LUT2 #(
		.INIT('h8)
	) name26103 (
		_w36114_,
		_w36173_,
		_w36615_
	);
	LUT2 #(
		.INIT('h4)
	) name26104 (
		_w36133_,
		_w36615_,
		_w36616_
	);
	LUT2 #(
		.INIT('h8)
	) name26105 (
		_w36117_,
		_w36141_,
		_w36617_
	);
	LUT2 #(
		.INIT('h4)
	) name26106 (
		_w36111_,
		_w36617_,
		_w36618_
	);
	LUT2 #(
		.INIT('h8)
	) name26107 (
		_w36135_,
		_w36166_,
		_w36619_
	);
	LUT2 #(
		.INIT('h4)
	) name26108 (
		_w36111_,
		_w36619_,
		_w36620_
	);
	LUT2 #(
		.INIT('h8)
	) name26109 (
		_w36107_,
		_w36149_,
		_w36621_
	);
	LUT2 #(
		.INIT('h4)
	) name26110 (
		_w36111_,
		_w36621_,
		_w36622_
	);
	LUT2 #(
		.INIT('h8)
	) name26111 (
		_w36107_,
		_w36137_,
		_w36623_
	);
	LUT2 #(
		.INIT('h4)
	) name26112 (
		_w36111_,
		_w36623_,
		_w36624_
	);
	LUT2 #(
		.INIT('h8)
	) name26113 (
		_w36114_,
		_w36149_,
		_w36625_
	);
	LUT2 #(
		.INIT('h4)
	) name26114 (
		_w36111_,
		_w36625_,
		_w36626_
	);
	LUT2 #(
		.INIT('h8)
	) name26115 (
		_w36114_,
		_w36137_,
		_w36627_
	);
	LUT2 #(
		.INIT('h4)
	) name26116 (
		_w36111_,
		_w36627_,
		_w36628_
	);
	LUT2 #(
		.INIT('h8)
	) name26117 (
		_w36117_,
		_w36149_,
		_w36629_
	);
	LUT2 #(
		.INIT('h4)
	) name26118 (
		_w36111_,
		_w36629_,
		_w36630_
	);
	LUT2 #(
		.INIT('h8)
	) name26119 (
		_w36117_,
		_w36137_,
		_w36631_
	);
	LUT2 #(
		.INIT('h4)
	) name26120 (
		_w36111_,
		_w36631_,
		_w36632_
	);
	LUT2 #(
		.INIT('h8)
	) name26121 (
		_w36158_,
		_w36185_,
		_w36633_
	);
	LUT2 #(
		.INIT('h4)
	) name26122 (
		_w36111_,
		_w36633_,
		_w36634_
	);
	LUT2 #(
		.INIT('h8)
	) name26123 (
		_w36162_,
		_w36185_,
		_w36635_
	);
	LUT2 #(
		.INIT('h4)
	) name26124 (
		_w36111_,
		_w36635_,
		_w36636_
	);
	LUT2 #(
		.INIT('h8)
	) name26125 (
		_w36173_,
		_w36274_,
		_w36637_
	);
	LUT2 #(
		.INIT('h4)
	) name26126 (
		_w36111_,
		_w36637_,
		_w36638_
	);
	LUT2 #(
		.INIT('h8)
	) name26127 (
		_w36158_,
		_w36165_,
		_w36639_
	);
	LUT2 #(
		.INIT('h4)
	) name26128 (
		_w36111_,
		_w36639_,
		_w36640_
	);
	LUT2 #(
		.INIT('h8)
	) name26129 (
		_w36162_,
		_w36165_,
		_w36641_
	);
	LUT2 #(
		.INIT('h4)
	) name26130 (
		_w36111_,
		_w36641_,
		_w36642_
	);
	LUT2 #(
		.INIT('h8)
	) name26131 (
		_w36158_,
		_w36170_,
		_w36643_
	);
	LUT2 #(
		.INIT('h4)
	) name26132 (
		_w36111_,
		_w36643_,
		_w36644_
	);
	LUT2 #(
		.INIT('h8)
	) name26133 (
		_w36162_,
		_w36170_,
		_w36645_
	);
	LUT2 #(
		.INIT('h4)
	) name26134 (
		_w36111_,
		_w36645_,
		_w36646_
	);
	LUT2 #(
		.INIT('h8)
	) name26135 (
		_w36173_,
		_w36185_,
		_w36647_
	);
	LUT2 #(
		.INIT('h4)
	) name26136 (
		_w36111_,
		_w36647_,
		_w36648_
	);
	LUT2 #(
		.INIT('h8)
	) name26137 (
		_w36166_,
		_w36185_,
		_w36649_
	);
	LUT2 #(
		.INIT('h4)
	) name26138 (
		_w36111_,
		_w36649_,
		_w36650_
	);
	LUT2 #(
		.INIT('h8)
	) name26139 (
		_w36165_,
		_w36173_,
		_w36651_
	);
	LUT2 #(
		.INIT('h4)
	) name26140 (
		_w36111_,
		_w36651_,
		_w36652_
	);
	LUT2 #(
		.INIT('h8)
	) name26141 (
		_w36166_,
		_w36274_,
		_w36653_
	);
	LUT2 #(
		.INIT('h4)
	) name26142 (
		_w36111_,
		_w36653_,
		_w36654_
	);
	LUT2 #(
		.INIT('h8)
	) name26143 (
		_w36170_,
		_w36173_,
		_w36655_
	);
	LUT2 #(
		.INIT('h4)
	) name26144 (
		_w36111_,
		_w36655_,
		_w36656_
	);
	LUT2 #(
		.INIT('h8)
	) name26145 (
		_w36156_,
		_w36166_,
		_w36657_
	);
	LUT2 #(
		.INIT('h4)
	) name26146 (
		_w36111_,
		_w36657_,
		_w36658_
	);
	LUT2 #(
		.INIT('h8)
	) name26147 (
		_w36181_,
		_w36185_,
		_w36659_
	);
	LUT2 #(
		.INIT('h4)
	) name26148 (
		_w36111_,
		_w36659_,
		_w36660_
	);
	LUT2 #(
		.INIT('h4)
	) name26149 (
		_w36101_,
		_w36635_,
		_w36661_
	);
	LUT2 #(
		.INIT('h4)
	) name26150 (
		_w36101_,
		_w36645_,
		_w36662_
	);
	LUT2 #(
		.INIT('h8)
	) name26151 (
		_w36176_,
		_w36185_,
		_w36663_
	);
	LUT2 #(
		.INIT('h4)
	) name26152 (
		_w36111_,
		_w36663_,
		_w36664_
	);
	LUT2 #(
		.INIT('h8)
	) name26153 (
		_w36165_,
		_w36181_,
		_w36665_
	);
	LUT2 #(
		.INIT('h4)
	) name26154 (
		_w36111_,
		_w36665_,
		_w36666_
	);
	LUT2 #(
		.INIT('h4)
	) name26155 (
		_w36101_,
		_w36631_,
		_w36667_
	);
	LUT2 #(
		.INIT('h8)
	) name26156 (
		_w36170_,
		_w36181_,
		_w36668_
	);
	LUT2 #(
		.INIT('h4)
	) name26157 (
		_w36111_,
		_w36668_,
		_w36669_
	);
	LUT2 #(
		.INIT('h8)
	) name26158 (
		_w36173_,
		_w36194_,
		_w36670_
	);
	LUT2 #(
		.INIT('h4)
	) name26159 (
		_w36111_,
		_w36670_,
		_w36671_
	);
	LUT2 #(
		.INIT('h4)
	) name26160 (
		_w36101_,
		_w36647_,
		_w36672_
	);
	LUT2 #(
		.INIT('h8)
	) name26161 (
		_w36156_,
		_w36176_,
		_w36673_
	);
	LUT2 #(
		.INIT('h4)
	) name26162 (
		_w36111_,
		_w36673_,
		_w36674_
	);
	LUT2 #(
		.INIT('h8)
	) name26163 (
		_w36185_,
		_w36189_,
		_w36675_
	);
	LUT2 #(
		.INIT('h4)
	) name26164 (
		_w36111_,
		_w36675_,
		_w36676_
	);
	LUT2 #(
		.INIT('h8)
	) name26165 (
		_w36165_,
		_w36186_,
		_w36677_
	);
	LUT2 #(
		.INIT('h4)
	) name26166 (
		_w36111_,
		_w36677_,
		_w36678_
	);
	LUT2 #(
		.INIT('h8)
	) name26167 (
		_w36170_,
		_w36186_,
		_w36679_
	);
	LUT2 #(
		.INIT('h4)
	) name26168 (
		_w36111_,
		_w36679_,
		_w36680_
	);
	LUT2 #(
		.INIT('h8)
	) name26169 (
		_w36156_,
		_w36189_,
		_w36681_
	);
	LUT2 #(
		.INIT('h4)
	) name26170 (
		_w36111_,
		_w36681_,
		_w36682_
	);
	LUT2 #(
		.INIT('h4)
	) name26171 (
		_w36101_,
		_w36639_,
		_w36683_
	);
	LUT2 #(
		.INIT('h8)
	) name26172 (
		_w36156_,
		_w36186_,
		_w36684_
	);
	LUT2 #(
		.INIT('h4)
	) name26173 (
		_w36111_,
		_w36684_,
		_w36685_
	);
	LUT2 #(
		.INIT('h8)
	) name26174 (
		_w36158_,
		_w36212_,
		_w36686_
	);
	LUT2 #(
		.INIT('h4)
	) name26175 (
		_w36111_,
		_w36686_,
		_w36687_
	);
	LUT2 #(
		.INIT('h8)
	) name26176 (
		_w36162_,
		_w36212_,
		_w36688_
	);
	LUT2 #(
		.INIT('h4)
	) name26177 (
		_w36111_,
		_w36688_,
		_w36689_
	);
	LUT2 #(
		.INIT('h4)
	) name26178 (
		_w36101_,
		_w36637_,
		_w36690_
	);
	LUT2 #(
		.INIT('h4)
	) name26179 (
		_w36101_,
		_w36653_,
		_w36691_
	);
	LUT2 #(
		.INIT('h8)
	) name26180 (
		_w36173_,
		_w36212_,
		_w36692_
	);
	LUT2 #(
		.INIT('h4)
	) name26181 (
		_w36111_,
		_w36692_,
		_w36693_
	);
	LUT2 #(
		.INIT('h8)
	) name26182 (
		_w36181_,
		_w36278_,
		_w36694_
	);
	LUT2 #(
		.INIT('h4)
	) name26183 (
		_w36111_,
		_w36694_,
		_w36695_
	);
	LUT2 #(
		.INIT('h8)
	) name26184 (
		_w36166_,
		_w36197_,
		_w36696_
	);
	LUT2 #(
		.INIT('h4)
	) name26185 (
		_w36111_,
		_w36696_,
		_w36697_
	);
	LUT2 #(
		.INIT('h8)
	) name26186 (
		_w36166_,
		_w36202_,
		_w36698_
	);
	LUT2 #(
		.INIT('h4)
	) name26187 (
		_w36111_,
		_w36698_,
		_w36699_
	);
	LUT2 #(
		.INIT('h4)
	) name26188 (
		_w36101_,
		_w36651_,
		_w36700_
	);
	LUT2 #(
		.INIT('h8)
	) name26189 (
		_w36166_,
		_w36207_,
		_w36701_
	);
	LUT2 #(
		.INIT('h4)
	) name26190 (
		_w36111_,
		_w36701_,
		_w36702_
	);
	LUT2 #(
		.INIT('h8)
	) name26191 (
		_w36181_,
		_w36212_,
		_w36703_
	);
	LUT2 #(
		.INIT('h4)
	) name26192 (
		_w36111_,
		_w36703_,
		_w36704_
	);
	LUT2 #(
		.INIT('h4)
	) name26193 (
		_w36101_,
		_w36643_,
		_w36705_
	);
	LUT2 #(
		.INIT('h8)
	) name26194 (
		_w36176_,
		_w36197_,
		_w36706_
	);
	LUT2 #(
		.INIT('h4)
	) name26195 (
		_w36111_,
		_w36706_,
		_w36707_
	);
	LUT2 #(
		.INIT('h8)
	) name26196 (
		_w36176_,
		_w36278_,
		_w36708_
	);
	LUT2 #(
		.INIT('h4)
	) name26197 (
		_w36111_,
		_w36708_,
		_w36709_
	);
	LUT2 #(
		.INIT('h4)
	) name26198 (
		_w36101_,
		_w36629_,
		_w36710_
	);
	LUT2 #(
		.INIT('h8)
	) name26199 (
		_w36119_,
		_w36278_,
		_w36711_
	);
	LUT2 #(
		.INIT('h4)
	) name26200 (
		_w36133_,
		_w36711_,
		_w36712_
	);
	LUT2 #(
		.INIT('h8)
	) name26201 (
		_w36176_,
		_w36202_,
		_w36713_
	);
	LUT2 #(
		.INIT('h4)
	) name26202 (
		_w36111_,
		_w36713_,
		_w36714_
	);
	LUT2 #(
		.INIT('h8)
	) name26203 (
		_w36176_,
		_w36207_,
		_w36715_
	);
	LUT2 #(
		.INIT('h4)
	) name26204 (
		_w36111_,
		_w36715_,
		_w36716_
	);
	LUT2 #(
		.INIT('h8)
	) name26205 (
		_w36186_,
		_w36212_,
		_w36717_
	);
	LUT2 #(
		.INIT('h4)
	) name26206 (
		_w36111_,
		_w36717_,
		_w36718_
	);
	LUT2 #(
		.INIT('h8)
	) name26207 (
		_w36189_,
		_w36197_,
		_w36719_
	);
	LUT2 #(
		.INIT('h4)
	) name26208 (
		_w36111_,
		_w36719_,
		_w36720_
	);
	LUT2 #(
		.INIT('h8)
	) name26209 (
		_w36186_,
		_w36197_,
		_w36721_
	);
	LUT2 #(
		.INIT('h4)
	) name26210 (
		_w36111_,
		_w36721_,
		_w36722_
	);
	LUT2 #(
		.INIT('h8)
	) name26211 (
		_w36189_,
		_w36202_,
		_w36723_
	);
	LUT2 #(
		.INIT('h4)
	) name26212 (
		_w36111_,
		_w36723_,
		_w36724_
	);
	LUT2 #(
		.INIT('h8)
	) name26213 (
		_w36186_,
		_w36202_,
		_w36725_
	);
	LUT2 #(
		.INIT('h4)
	) name26214 (
		_w36111_,
		_w36725_,
		_w36726_
	);
	LUT2 #(
		.INIT('h4)
	) name26215 (
		_w36101_,
		_w36592_,
		_w36727_
	);
	LUT2 #(
		.INIT('h8)
	) name26216 (
		_w36135_,
		_w36181_,
		_w36728_
	);
	LUT2 #(
		.INIT('h4)
	) name26217 (
		_w36111_,
		_w36728_,
		_w36729_
	);
	LUT2 #(
		.INIT('h8)
	) name26218 (
		_w36189_,
		_w36207_,
		_w36730_
	);
	LUT2 #(
		.INIT('h4)
	) name26219 (
		_w36111_,
		_w36730_,
		_w36731_
	);
	LUT2 #(
		.INIT('h8)
	) name26220 (
		_w36186_,
		_w36207_,
		_w36732_
	);
	LUT2 #(
		.INIT('h4)
	) name26221 (
		_w36111_,
		_w36732_,
		_w36733_
	);
	LUT2 #(
		.INIT('h8)
	) name26222 (
		_w36119_,
		_w36185_,
		_w36734_
	);
	LUT2 #(
		.INIT('h4)
	) name26223 (
		_w36111_,
		_w36734_,
		_w36735_
	);
	LUT2 #(
		.INIT('h8)
	) name26224 (
		_w36104_,
		_w36185_,
		_w36736_
	);
	LUT2 #(
		.INIT('h4)
	) name26225 (
		_w36111_,
		_w36736_,
		_w36737_
	);
	LUT2 #(
		.INIT('h8)
	) name26226 (
		_w36119_,
		_w36165_,
		_w36738_
	);
	LUT2 #(
		.INIT('h4)
	) name26227 (
		_w36111_,
		_w36738_,
		_w36739_
	);
	LUT2 #(
		.INIT('h8)
	) name26228 (
		_w36119_,
		_w36170_,
		_w36740_
	);
	LUT2 #(
		.INIT('h4)
	) name26229 (
		_w36111_,
		_w36740_,
		_w36741_
	);
	LUT2 #(
		.INIT('h8)
	) name26230 (
		_w36104_,
		_w36156_,
		_w36742_
	);
	LUT2 #(
		.INIT('h4)
	) name26231 (
		_w36111_,
		_w36742_,
		_w36743_
	);
	LUT2 #(
		.INIT('h8)
	) name26232 (
		_w36135_,
		_w36176_,
		_w36744_
	);
	LUT2 #(
		.INIT('h4)
	) name26233 (
		_w36111_,
		_w36744_,
		_w36745_
	);
	LUT2 #(
		.INIT('h8)
	) name26234 (
		_w36162_,
		_w36278_,
		_w36746_
	);
	LUT2 #(
		.INIT('h4)
	) name26235 (
		_w36111_,
		_w36746_,
		_w36747_
	);
	LUT2 #(
		.INIT('h8)
	) name26236 (
		_w36127_,
		_w36185_,
		_w36748_
	);
	LUT2 #(
		.INIT('h4)
	) name26237 (
		_w36111_,
		_w36748_,
		_w36749_
	);
	LUT2 #(
		.INIT('h4)
	) name26238 (
		_w36101_,
		_w36627_,
		_w36750_
	);
	LUT2 #(
		.INIT('h8)
	) name26239 (
		_w36123_,
		_w36165_,
		_w36751_
	);
	LUT2 #(
		.INIT('h4)
	) name26240 (
		_w36111_,
		_w36751_,
		_w36752_
	);
	LUT2 #(
		.INIT('h8)
	) name26241 (
		_w36123_,
		_w36170_,
		_w36753_
	);
	LUT2 #(
		.INIT('h4)
	) name26242 (
		_w36111_,
		_w36753_,
		_w36754_
	);
	LUT2 #(
		.INIT('h8)
	) name26243 (
		_w36127_,
		_w36156_,
		_w36755_
	);
	LUT2 #(
		.INIT('h4)
	) name26244 (
		_w36111_,
		_w36755_,
		_w36756_
	);
	LUT2 #(
		.INIT('h8)
	) name26245 (
		_w36123_,
		_w36156_,
		_w36757_
	);
	LUT2 #(
		.INIT('h4)
	) name26246 (
		_w36111_,
		_w36757_,
		_w36758_
	);
	LUT2 #(
		.INIT('h8)
	) name26247 (
		_w36144_,
		_w36185_,
		_w36759_
	);
	LUT2 #(
		.INIT('h4)
	) name26248 (
		_w36111_,
		_w36759_,
		_w36760_
	);
	LUT2 #(
		.INIT('h8)
	) name26249 (
		_w36181_,
		_w36274_,
		_w36761_
	);
	LUT2 #(
		.INIT('h4)
	) name26250 (
		_w36111_,
		_w36761_,
		_w36762_
	);
	LUT2 #(
		.INIT('h8)
	) name26251 (
		_w36141_,
		_w36165_,
		_w36763_
	);
	LUT2 #(
		.INIT('h4)
	) name26252 (
		_w36111_,
		_w36763_,
		_w36764_
	);
	LUT2 #(
		.INIT('h8)
	) name26253 (
		_w36141_,
		_w36170_,
		_w36765_
	);
	LUT2 #(
		.INIT('h4)
	) name26254 (
		_w36111_,
		_w36765_,
		_w36766_
	);
	LUT2 #(
		.INIT('h8)
	) name26255 (
		_w36144_,
		_w36156_,
		_w36767_
	);
	LUT2 #(
		.INIT('h4)
	) name26256 (
		_w36111_,
		_w36767_,
		_w36768_
	);
	LUT2 #(
		.INIT('h8)
	) name26257 (
		_w36141_,
		_w36156_,
		_w36769_
	);
	LUT2 #(
		.INIT('h4)
	) name26258 (
		_w36111_,
		_w36769_,
		_w36770_
	);
	LUT2 #(
		.INIT('h8)
	) name26259 (
		_w36135_,
		_w36144_,
		_w36771_
	);
	LUT2 #(
		.INIT('h4)
	) name26260 (
		_w36133_,
		_w36771_,
		_w36772_
	);
	LUT2 #(
		.INIT('h8)
	) name26261 (
		_w36149_,
		_w36165_,
		_w36773_
	);
	LUT2 #(
		.INIT('h4)
	) name26262 (
		_w36111_,
		_w36773_,
		_w36774_
	);
	LUT2 #(
		.INIT('h8)
	) name26263 (
		_w36137_,
		_w36165_,
		_w36775_
	);
	LUT2 #(
		.INIT('h4)
	) name26264 (
		_w36111_,
		_w36775_,
		_w36776_
	);
	LUT2 #(
		.INIT('h8)
	) name26265 (
		_w36176_,
		_w36274_,
		_w36777_
	);
	LUT2 #(
		.INIT('h4)
	) name26266 (
		_w36111_,
		_w36777_,
		_w36778_
	);
	LUT2 #(
		.INIT('h8)
	) name26267 (
		_w36149_,
		_w36170_,
		_w36779_
	);
	LUT2 #(
		.INIT('h4)
	) name26268 (
		_w36111_,
		_w36779_,
		_w36780_
	);
	LUT2 #(
		.INIT('h8)
	) name26269 (
		_w36137_,
		_w36170_,
		_w36781_
	);
	LUT2 #(
		.INIT('h4)
	) name26270 (
		_w36111_,
		_w36781_,
		_w36782_
	);
	LUT2 #(
		.INIT('h4)
	) name26271 (
		_w36133_,
		_w36590_,
		_w36783_
	);
	LUT2 #(
		.INIT('h8)
	) name26272 (
		_w36149_,
		_w36156_,
		_w36784_
	);
	LUT2 #(
		.INIT('h4)
	) name26273 (
		_w36111_,
		_w36784_,
		_w36785_
	);
	LUT2 #(
		.INIT('h8)
	) name26274 (
		_w36137_,
		_w36156_,
		_w36786_
	);
	LUT2 #(
		.INIT('h4)
	) name26275 (
		_w36111_,
		_w36786_,
		_w36787_
	);
	LUT2 #(
		.INIT('h8)
	) name26276 (
		_w36119_,
		_w36212_,
		_w36788_
	);
	LUT2 #(
		.INIT('h4)
	) name26277 (
		_w36111_,
		_w36788_,
		_w36789_
	);
	LUT2 #(
		.INIT('h4)
	) name26278 (
		_w36133_,
		_w36592_,
		_w36790_
	);
	LUT2 #(
		.INIT('h8)
	) name26279 (
		_w36104_,
		_w36197_,
		_w36791_
	);
	LUT2 #(
		.INIT('h4)
	) name26280 (
		_w36111_,
		_w36791_,
		_w36792_
	);
	LUT2 #(
		.INIT('h8)
	) name26281 (
		_w36104_,
		_w36202_,
		_w36793_
	);
	LUT2 #(
		.INIT('h4)
	) name26282 (
		_w36111_,
		_w36793_,
		_w36794_
	);
	LUT2 #(
		.INIT('h8)
	) name26283 (
		_w36181_,
		_w36194_,
		_w36795_
	);
	LUT2 #(
		.INIT('h4)
	) name26284 (
		_w36111_,
		_w36795_,
		_w36796_
	);
	LUT2 #(
		.INIT('h4)
	) name26285 (
		_w36133_,
		_w36594_,
		_w36797_
	);
	LUT2 #(
		.INIT('h8)
	) name26286 (
		_w36104_,
		_w36207_,
		_w36798_
	);
	LUT2 #(
		.INIT('h4)
	) name26287 (
		_w36111_,
		_w36798_,
		_w36799_
	);
	LUT2 #(
		.INIT('h4)
	) name26288 (
		_w36133_,
		_w36596_,
		_w36800_
	);
	LUT2 #(
		.INIT('h8)
	) name26289 (
		_w36123_,
		_w36212_,
		_w36801_
	);
	LUT2 #(
		.INIT('h4)
	) name26290 (
		_w36111_,
		_w36801_,
		_w36802_
	);
	LUT2 #(
		.INIT('h8)
	) name26291 (
		_w36127_,
		_w36197_,
		_w36803_
	);
	LUT2 #(
		.INIT('h4)
	) name26292 (
		_w36111_,
		_w36803_,
		_w36804_
	);
	LUT2 #(
		.INIT('h8)
	) name26293 (
		_w36123_,
		_w36197_,
		_w36805_
	);
	LUT2 #(
		.INIT('h4)
	) name26294 (
		_w36111_,
		_w36805_,
		_w36806_
	);
	LUT2 #(
		.INIT('h8)
	) name26295 (
		_w36127_,
		_w36202_,
		_w36807_
	);
	LUT2 #(
		.INIT('h4)
	) name26296 (
		_w36111_,
		_w36807_,
		_w36808_
	);
	LUT2 #(
		.INIT('h8)
	) name26297 (
		_w36123_,
		_w36202_,
		_w36809_
	);
	LUT2 #(
		.INIT('h4)
	) name26298 (
		_w36111_,
		_w36809_,
		_w36810_
	);
	LUT2 #(
		.INIT('h8)
	) name26299 (
		_w36127_,
		_w36207_,
		_w36811_
	);
	LUT2 #(
		.INIT('h4)
	) name26300 (
		_w36111_,
		_w36811_,
		_w36812_
	);
	LUT2 #(
		.INIT('h4)
	) name26301 (
		_w36133_,
		_w36598_,
		_w36813_
	);
	LUT2 #(
		.INIT('h8)
	) name26302 (
		_w36123_,
		_w36207_,
		_w36814_
	);
	LUT2 #(
		.INIT('h4)
	) name26303 (
		_w36111_,
		_w36814_,
		_w36815_
	);
	LUT2 #(
		.INIT('h8)
	) name26304 (
		_w36162_,
		_w36194_,
		_w36816_
	);
	LUT2 #(
		.INIT('h4)
	) name26305 (
		_w36133_,
		_w36816_,
		_w36817_
	);
	LUT2 #(
		.INIT('h8)
	) name26306 (
		_w36141_,
		_w36212_,
		_w36818_
	);
	LUT2 #(
		.INIT('h4)
	) name26307 (
		_w36111_,
		_w36818_,
		_w36819_
	);
	LUT2 #(
		.INIT('h4)
	) name26308 (
		_w36133_,
		_w36600_,
		_w36820_
	);
	LUT2 #(
		.INIT('h8)
	) name26309 (
		_w36144_,
		_w36197_,
		_w36821_
	);
	LUT2 #(
		.INIT('h4)
	) name26310 (
		_w36111_,
		_w36821_,
		_w36822_
	);
	LUT2 #(
		.INIT('h8)
	) name26311 (
		_w36141_,
		_w36197_,
		_w36823_
	);
	LUT2 #(
		.INIT('h4)
	) name26312 (
		_w36111_,
		_w36823_,
		_w36824_
	);
	LUT2 #(
		.INIT('h4)
	) name26313 (
		_w36133_,
		_w36602_,
		_w36825_
	);
	LUT2 #(
		.INIT('h8)
	) name26314 (
		_w36144_,
		_w36202_,
		_w36826_
	);
	LUT2 #(
		.INIT('h4)
	) name26315 (
		_w36111_,
		_w36826_,
		_w36827_
	);
	LUT2 #(
		.INIT('h8)
	) name26316 (
		_w36141_,
		_w36202_,
		_w36828_
	);
	LUT2 #(
		.INIT('h4)
	) name26317 (
		_w36111_,
		_w36828_,
		_w36829_
	);
	LUT2 #(
		.INIT('h4)
	) name26318 (
		_w36133_,
		_w36604_,
		_w36830_
	);
	LUT2 #(
		.INIT('h8)
	) name26319 (
		_w36144_,
		_w36207_,
		_w36831_
	);
	LUT2 #(
		.INIT('h4)
	) name26320 (
		_w36111_,
		_w36831_,
		_w36832_
	);
	LUT2 #(
		.INIT('h8)
	) name26321 (
		_w36141_,
		_w36207_,
		_w36833_
	);
	LUT2 #(
		.INIT('h4)
	) name26322 (
		_w36111_,
		_w36833_,
		_w36834_
	);
	LUT2 #(
		.INIT('h4)
	) name26323 (
		_w36133_,
		_w36606_,
		_w36835_
	);
	LUT2 #(
		.INIT('h8)
	) name26324 (
		_w36149_,
		_w36212_,
		_w36836_
	);
	LUT2 #(
		.INIT('h4)
	) name26325 (
		_w36111_,
		_w36836_,
		_w36837_
	);
	LUT2 #(
		.INIT('h8)
	) name26326 (
		_w36137_,
		_w36212_,
		_w36838_
	);
	LUT2 #(
		.INIT('h4)
	) name26327 (
		_w36111_,
		_w36838_,
		_w36839_
	);
	LUT2 #(
		.INIT('h4)
	) name26328 (
		_w36133_,
		_w36608_,
		_w36840_
	);
	LUT2 #(
		.INIT('h8)
	) name26329 (
		_w36189_,
		_w36278_,
		_w36841_
	);
	LUT2 #(
		.INIT('h4)
	) name26330 (
		_w36111_,
		_w36841_,
		_w36842_
	);
	LUT2 #(
		.INIT('h8)
	) name26331 (
		_w36149_,
		_w36197_,
		_w36843_
	);
	LUT2 #(
		.INIT('h4)
	) name26332 (
		_w36111_,
		_w36843_,
		_w36844_
	);
	LUT2 #(
		.INIT('h8)
	) name26333 (
		_w36137_,
		_w36197_,
		_w36845_
	);
	LUT2 #(
		.INIT('h4)
	) name26334 (
		_w36111_,
		_w36845_,
		_w36846_
	);
	LUT2 #(
		.INIT('h8)
	) name26335 (
		_w36149_,
		_w36202_,
		_w36847_
	);
	LUT2 #(
		.INIT('h4)
	) name26336 (
		_w36111_,
		_w36847_,
		_w36848_
	);
	LUT2 #(
		.INIT('h8)
	) name26337 (
		_w36137_,
		_w36202_,
		_w36849_
	);
	LUT2 #(
		.INIT('h4)
	) name26338 (
		_w36111_,
		_w36849_,
		_w36850_
	);
	LUT2 #(
		.INIT('h4)
	) name26339 (
		_w36101_,
		_w36625_,
		_w36851_
	);
	LUT2 #(
		.INIT('h8)
	) name26340 (
		_w36149_,
		_w36207_,
		_w36852_
	);
	LUT2 #(
		.INIT('h4)
	) name26341 (
		_w36111_,
		_w36852_,
		_w36853_
	);
	LUT2 #(
		.INIT('h4)
	) name26342 (
		_w36133_,
		_w36588_,
		_w36854_
	);
	LUT2 #(
		.INIT('h8)
	) name26343 (
		_w36137_,
		_w36207_,
		_w36855_
	);
	LUT2 #(
		.INIT('h4)
	) name26344 (
		_w36111_,
		_w36855_,
		_w36856_
	);
	LUT2 #(
		.INIT('h8)
	) name26345 (
		_w36135_,
		_w36189_,
		_w36857_
	);
	LUT2 #(
		.INIT('h4)
	) name26346 (
		_w36111_,
		_w36857_,
		_w36858_
	);
	LUT2 #(
		.INIT('h4)
	) name26347 (
		_w36133_,
		_w36611_,
		_w36859_
	);
	LUT2 #(
		.INIT('h8)
	) name26348 (
		_w36189_,
		_w36274_,
		_w36860_
	);
	LUT2 #(
		.INIT('h4)
	) name26349 (
		_w36111_,
		_w36860_,
		_w36861_
	);
	LUT2 #(
		.INIT('h8)
	) name26350 (
		_w36135_,
		_w36158_,
		_w36862_
	);
	LUT2 #(
		.INIT('h4)
	) name26351 (
		_w36111_,
		_w36862_,
		_w36863_
	);
	LUT2 #(
		.INIT('h4)
	) name26352 (
		_w36133_,
		_w36613_,
		_w36864_
	);
	LUT2 #(
		.INIT('h4)
	) name26353 (
		_w36133_,
		_w36617_,
		_w36865_
	);
	LUT2 #(
		.INIT('h8)
	) name26354 (
		_w36186_,
		_w36194_,
		_w36866_
	);
	LUT2 #(
		.INIT('h4)
	) name26355 (
		_w36111_,
		_w36866_,
		_w36867_
	);
	LUT2 #(
		.INIT('h8)
	) name26356 (
		_w36124_,
		_w36158_,
		_w36868_
	);
	LUT2 #(
		.INIT('h4)
	) name26357 (
		_w36111_,
		_w36868_,
		_w36869_
	);
	LUT2 #(
		.INIT('h4)
	) name26358 (
		_w36133_,
		_w36619_,
		_w36870_
	);
	LUT2 #(
		.INIT('h8)
	) name26359 (
		_w36124_,
		_w36162_,
		_w36871_
	);
	LUT2 #(
		.INIT('h4)
	) name26360 (
		_w36111_,
		_w36871_,
		_w36872_
	);
	LUT2 #(
		.INIT('h8)
	) name26361 (
		_w36107_,
		_w36158_,
		_w36873_
	);
	LUT2 #(
		.INIT('h4)
	) name26362 (
		_w36111_,
		_w36873_,
		_w36874_
	);
	LUT2 #(
		.INIT('h8)
	) name26363 (
		_w36107_,
		_w36162_,
		_w36875_
	);
	LUT2 #(
		.INIT('h4)
	) name26364 (
		_w36111_,
		_w36875_,
		_w36876_
	);
	LUT2 #(
		.INIT('h8)
	) name26365 (
		_w36114_,
		_w36158_,
		_w36877_
	);
	LUT2 #(
		.INIT('h4)
	) name26366 (
		_w36111_,
		_w36877_,
		_w36878_
	);
	LUT2 #(
		.INIT('h8)
	) name26367 (
		_w36114_,
		_w36162_,
		_w36879_
	);
	LUT2 #(
		.INIT('h4)
	) name26368 (
		_w36111_,
		_w36879_,
		_w36880_
	);
	LUT2 #(
		.INIT('h4)
	) name26369 (
		_w36133_,
		_w36621_,
		_w36881_
	);
	LUT2 #(
		.INIT('h8)
	) name26370 (
		_w36135_,
		_w36162_,
		_w36882_
	);
	LUT2 #(
		.INIT('h4)
	) name26371 (
		_w36111_,
		_w36882_,
		_w36883_
	);
	LUT2 #(
		.INIT('h8)
	) name26372 (
		_w36124_,
		_w36173_,
		_w36884_
	);
	LUT2 #(
		.INIT('h4)
	) name26373 (
		_w36111_,
		_w36884_,
		_w36885_
	);
	LUT2 #(
		.INIT('h4)
	) name26374 (
		_w36133_,
		_w36623_,
		_w36886_
	);
	LUT2 #(
		.INIT('h8)
	) name26375 (
		_w36124_,
		_w36166_,
		_w36887_
	);
	LUT2 #(
		.INIT('h4)
	) name26376 (
		_w36111_,
		_w36887_,
		_w36888_
	);
	LUT2 #(
		.INIT('h8)
	) name26377 (
		_w36107_,
		_w36173_,
		_w36889_
	);
	LUT2 #(
		.INIT('h4)
	) name26378 (
		_w36111_,
		_w36889_,
		_w36890_
	);
	LUT2 #(
		.INIT('h4)
	) name26379 (
		_w36133_,
		_w36625_,
		_w36891_
	);
	LUT2 #(
		.INIT('h4)
	) name26380 (
		_w36111_,
		_w36615_,
		_w36892_
	);
	LUT2 #(
		.INIT('h4)
	) name26381 (
		_w36133_,
		_w36627_,
		_w36893_
	);
	LUT2 #(
		.INIT('h4)
	) name26382 (
		_w36133_,
		_w36629_,
		_w36894_
	);
	LUT2 #(
		.INIT('h8)
	) name26383 (
		_w36117_,
		_w36166_,
		_w36895_
	);
	LUT2 #(
		.INIT('h4)
	) name26384 (
		_w36111_,
		_w36895_,
		_w36896_
	);
	LUT2 #(
		.INIT('h8)
	) name26385 (
		_w36124_,
		_w36181_,
		_w36897_
	);
	LUT2 #(
		.INIT('h4)
	) name26386 (
		_w36111_,
		_w36897_,
		_w36898_
	);
	LUT2 #(
		.INIT('h4)
	) name26387 (
		_w36133_,
		_w36631_,
		_w36899_
	);
	LUT2 #(
		.INIT('h8)
	) name26388 (
		_w36124_,
		_w36176_,
		_w36900_
	);
	LUT2 #(
		.INIT('h4)
	) name26389 (
		_w36111_,
		_w36900_,
		_w36901_
	);
	LUT2 #(
		.INIT('h8)
	) name26390 (
		_w36158_,
		_w36274_,
		_w36902_
	);
	LUT2 #(
		.INIT('h4)
	) name26391 (
		_w36111_,
		_w36902_,
		_w36903_
	);
	LUT2 #(
		.INIT('h4)
	) name26392 (
		_w36133_,
		_w36633_,
		_w36904_
	);
	LUT2 #(
		.INIT('h8)
	) name26393 (
		_w36107_,
		_w36181_,
		_w36905_
	);
	LUT2 #(
		.INIT('h4)
	) name26394 (
		_w36111_,
		_w36905_,
		_w36906_
	);
	LUT2 #(
		.INIT('h4)
	) name26395 (
		_w36133_,
		_w36635_,
		_w36907_
	);
	LUT2 #(
		.INIT('h8)
	) name26396 (
		_w36114_,
		_w36181_,
		_w36908_
	);
	LUT2 #(
		.INIT('h4)
	) name26397 (
		_w36111_,
		_w36908_,
		_w36909_
	);
	LUT2 #(
		.INIT('h4)
	) name26398 (
		_w36133_,
		_w36637_,
		_w36910_
	);
	LUT2 #(
		.INIT('h8)
	) name26399 (
		_w36117_,
		_w36176_,
		_w36911_
	);
	LUT2 #(
		.INIT('h4)
	) name26400 (
		_w36111_,
		_w36911_,
		_w36912_
	);
	LUT2 #(
		.INIT('h4)
	) name26401 (
		_w36133_,
		_w36639_,
		_w36913_
	);
	LUT2 #(
		.INIT('h8)
	) name26402 (
		_w36124_,
		_w36189_,
		_w36914_
	);
	LUT2 #(
		.INIT('h4)
	) name26403 (
		_w36111_,
		_w36914_,
		_w36915_
	);
	LUT2 #(
		.INIT('h4)
	) name26404 (
		_w36133_,
		_w36641_,
		_w36916_
	);
	LUT2 #(
		.INIT('h8)
	) name26405 (
		_w36107_,
		_w36186_,
		_w36917_
	);
	LUT2 #(
		.INIT('h4)
	) name26406 (
		_w36111_,
		_w36917_,
		_w36918_
	);
	LUT2 #(
		.INIT('h4)
	) name26407 (
		_w36133_,
		_w36643_,
		_w36919_
	);
	LUT2 #(
		.INIT('h8)
	) name26408 (
		_w36162_,
		_w36274_,
		_w36920_
	);
	LUT2 #(
		.INIT('h4)
	) name26409 (
		_w36111_,
		_w36920_,
		_w36921_
	);
	LUT2 #(
		.INIT('h4)
	) name26410 (
		_w36133_,
		_w36645_,
		_w36922_
	);
	LUT2 #(
		.INIT('h8)
	) name26411 (
		_w36114_,
		_w36186_,
		_w36923_
	);
	LUT2 #(
		.INIT('h4)
	) name26412 (
		_w36111_,
		_w36923_,
		_w36924_
	);
	LUT2 #(
		.INIT('h8)
	) name26413 (
		_w36117_,
		_w36189_,
		_w36925_
	);
	LUT2 #(
		.INIT('h4)
	) name26414 (
		_w36111_,
		_w36925_,
		_w36926_
	);
	LUT2 #(
		.INIT('h8)
	) name26415 (
		_w36117_,
		_w36186_,
		_w36927_
	);
	LUT2 #(
		.INIT('h4)
	) name26416 (
		_w36111_,
		_w36927_,
		_w36928_
	);
	LUT2 #(
		.INIT('h4)
	) name26417 (
		_w36111_,
		_w36711_,
		_w36929_
	);
	LUT2 #(
		.INIT('h8)
	) name26418 (
		_w36104_,
		_w36278_,
		_w36930_
	);
	LUT2 #(
		.INIT('h4)
	) name26419 (
		_w36111_,
		_w36930_,
		_w36931_
	);
	LUT2 #(
		.INIT('h4)
	) name26420 (
		_w36133_,
		_w36923_,
		_w36932_
	);
	LUT2 #(
		.INIT('h8)
	) name26421 (
		_w36119_,
		_w36135_,
		_w36933_
	);
	LUT2 #(
		.INIT('h4)
	) name26422 (
		_w36111_,
		_w36933_,
		_w36934_
	);
	LUT2 #(
		.INIT('h8)
	) name26423 (
		_w36104_,
		_w36135_,
		_w36935_
	);
	LUT2 #(
		.INIT('h4)
	) name26424 (
		_w36111_,
		_w36935_,
		_w36936_
	);
	LUT2 #(
		.INIT('h4)
	) name26425 (
		_w36133_,
		_w36647_,
		_w36937_
	);
	LUT2 #(
		.INIT('h8)
	) name26426 (
		_w36119_,
		_w36274_,
		_w36938_
	);
	LUT2 #(
		.INIT('h4)
	) name26427 (
		_w36111_,
		_w36938_,
		_w36939_
	);
	LUT2 #(
		.INIT('h8)
	) name26428 (
		_w36104_,
		_w36274_,
		_w36940_
	);
	LUT2 #(
		.INIT('h4)
	) name26429 (
		_w36111_,
		_w36940_,
		_w36941_
	);
	LUT2 #(
		.INIT('h4)
	) name26430 (
		_w36133_,
		_w36649_,
		_w36942_
	);
	LUT2 #(
		.INIT('h8)
	) name26431 (
		_w36158_,
		_w36194_,
		_w36943_
	);
	LUT2 #(
		.INIT('h4)
	) name26432 (
		_w36111_,
		_w36943_,
		_w36944_
	);
	LUT2 #(
		.INIT('h8)
	) name26433 (
		_w36119_,
		_w36194_,
		_w36945_
	);
	LUT2 #(
		.INIT('h4)
	) name26434 (
		_w36111_,
		_w36945_,
		_w36946_
	);
	LUT2 #(
		.INIT('h4)
	) name26435 (
		_w36133_,
		_w36651_,
		_w36947_
	);
	LUT2 #(
		.INIT('h8)
	) name26436 (
		_w36127_,
		_w36278_,
		_w36948_
	);
	LUT2 #(
		.INIT('h4)
	) name26437 (
		_w36111_,
		_w36948_,
		_w36949_
	);
	LUT2 #(
		.INIT('h8)
	) name26438 (
		_w36127_,
		_w36135_,
		_w36950_
	);
	LUT2 #(
		.INIT('h4)
	) name26439 (
		_w36111_,
		_w36950_,
		_w36951_
	);
	LUT2 #(
		.INIT('h4)
	) name26440 (
		_w36133_,
		_w36653_,
		_w36952_
	);
	LUT2 #(
		.INIT('h8)
	) name26441 (
		_w36127_,
		_w36274_,
		_w36953_
	);
	LUT2 #(
		.INIT('h4)
	) name26442 (
		_w36111_,
		_w36953_,
		_w36954_
	);
	LUT2 #(
		.INIT('h4)
	) name26443 (
		_w36133_,
		_w36655_,
		_w36955_
	);
	LUT2 #(
		.INIT('h8)
	) name26444 (
		_w36123_,
		_w36194_,
		_w36956_
	);
	LUT2 #(
		.INIT('h4)
	) name26445 (
		_w36111_,
		_w36956_,
		_w36957_
	);
	LUT2 #(
		.INIT('h4)
	) name26446 (
		_w36111_,
		_w36816_,
		_w36958_
	);
	LUT2 #(
		.INIT('h8)
	) name26447 (
		_w36144_,
		_w36278_,
		_w36959_
	);
	LUT2 #(
		.INIT('h4)
	) name26448 (
		_w36111_,
		_w36959_,
		_w36960_
	);
	LUT2 #(
		.INIT('h4)
	) name26449 (
		_w36133_,
		_w36657_,
		_w36961_
	);
	LUT2 #(
		.INIT('h4)
	) name26450 (
		_w36111_,
		_w36771_,
		_w36962_
	);
	LUT2 #(
		.INIT('h4)
	) name26451 (
		_w36133_,
		_w36659_,
		_w36963_
	);
	LUT2 #(
		.INIT('h8)
	) name26452 (
		_w36144_,
		_w36274_,
		_w36964_
	);
	LUT2 #(
		.INIT('h4)
	) name26453 (
		_w36111_,
		_w36964_,
		_w36965_
	);
	LUT2 #(
		.INIT('h8)
	) name26454 (
		_w36137_,
		_w36194_,
		_w36966_
	);
	LUT2 #(
		.INIT('h4)
	) name26455 (
		_w36351_,
		_w36966_,
		_w36967_
	);
	LUT2 #(
		.INIT('h4)
	) name26456 (
		_w36133_,
		_w36663_,
		_w36968_
	);
	LUT2 #(
		.INIT('h8)
	) name26457 (
		_w36141_,
		_w36194_,
		_w36969_
	);
	LUT2 #(
		.INIT('h4)
	) name26458 (
		_w36111_,
		_w36969_,
		_w36970_
	);
	LUT2 #(
		.INIT('h4)
	) name26459 (
		_w36133_,
		_w36665_,
		_w36971_
	);
	LUT2 #(
		.INIT('h8)
	) name26460 (
		_w36173_,
		_w36278_,
		_w36972_
	);
	LUT2 #(
		.INIT('h4)
	) name26461 (
		_w36111_,
		_w36972_,
		_w36973_
	);
	LUT2 #(
		.INIT('h4)
	) name26462 (
		_w36133_,
		_w36668_,
		_w36974_
	);
	LUT2 #(
		.INIT('h8)
	) name26463 (
		_w36149_,
		_w36194_,
		_w36975_
	);
	LUT2 #(
		.INIT('h4)
	) name26464 (
		_w36111_,
		_w36975_,
		_w36976_
	);
	LUT2 #(
		.INIT('h4)
	) name26465 (
		_w36133_,
		_w36670_,
		_w36977_
	);
	LUT2 #(
		.INIT('h4)
	) name26466 (
		_w36111_,
		_w36966_,
		_w36978_
	);
	LUT2 #(
		.INIT('h4)
	) name26467 (
		_w36351_,
		_w36975_,
		_w36979_
	);
	LUT2 #(
		.INIT('h8)
	) name26468 (
		_w36119_,
		_w36124_,
		_w36980_
	);
	LUT2 #(
		.INIT('h4)
	) name26469 (
		_w36111_,
		_w36980_,
		_w36981_
	);
	LUT2 #(
		.INIT('h8)
	) name26470 (
		_w36104_,
		_w36124_,
		_w36982_
	);
	LUT2 #(
		.INIT('h4)
	) name26471 (
		_w36111_,
		_w36982_,
		_w36983_
	);
	LUT2 #(
		.INIT('h8)
	) name26472 (
		_w36107_,
		_w36119_,
		_w36984_
	);
	LUT2 #(
		.INIT('h4)
	) name26473 (
		_w36111_,
		_w36984_,
		_w36985_
	);
	LUT2 #(
		.INIT('h4)
	) name26474 (
		_w36133_,
		_w36673_,
		_w36986_
	);
	LUT2 #(
		.INIT('h4)
	) name26475 (
		_w36111_,
		_w36586_,
		_w36987_
	);
	LUT2 #(
		.INIT('h4)
	) name26476 (
		_w36133_,
		_w36675_,
		_w36988_
	);
	LUT2 #(
		.INIT('h4)
	) name26477 (
		_w36351_,
		_w36590_,
		_w36989_
	);
	LUT2 #(
		.INIT('h4)
	) name26478 (
		_w36351_,
		_w36592_,
		_w36990_
	);
	LUT2 #(
		.INIT('h4)
	) name26479 (
		_w36133_,
		_w36920_,
		_w36991_
	);
	LUT2 #(
		.INIT('h4)
	) name26480 (
		_w36351_,
		_w36594_,
		_w36992_
	);
	LUT2 #(
		.INIT('h4)
	) name26481 (
		_w36101_,
		_w36633_,
		_w36993_
	);
	LUT2 #(
		.INIT('h4)
	) name26482 (
		_w36351_,
		_w36596_,
		_w36994_
	);
	LUT2 #(
		.INIT('h4)
	) name26483 (
		_w36133_,
		_w36677_,
		_w36995_
	);
	LUT2 #(
		.INIT('h4)
	) name26484 (
		_w36351_,
		_w36598_,
		_w36996_
	);
	LUT2 #(
		.INIT('h4)
	) name26485 (
		_w36133_,
		_w36679_,
		_w36997_
	);
	LUT2 #(
		.INIT('h4)
	) name26486 (
		_w36351_,
		_w36600_,
		_w36998_
	);
	LUT2 #(
		.INIT('h4)
	) name26487 (
		_w36351_,
		_w36602_,
		_w36999_
	);
	LUT2 #(
		.INIT('h4)
	) name26488 (
		_w36133_,
		_w36681_,
		_w37000_
	);
	LUT2 #(
		.INIT('h4)
	) name26489 (
		_w36351_,
		_w36604_,
		_w37001_
	);
	LUT2 #(
		.INIT('h4)
	) name26490 (
		_w36351_,
		_w36606_,
		_w37002_
	);
	LUT2 #(
		.INIT('h4)
	) name26491 (
		_w36133_,
		_w36684_,
		_w37003_
	);
	LUT2 #(
		.INIT('h4)
	) name26492 (
		_w36351_,
		_w36608_,
		_w37004_
	);
	LUT2 #(
		.INIT('h4)
	) name26493 (
		_w36351_,
		_w36588_,
		_w37005_
	);
	LUT2 #(
		.INIT('h4)
	) name26494 (
		_w36133_,
		_w36686_,
		_w37006_
	);
	LUT2 #(
		.INIT('h4)
	) name26495 (
		_w36351_,
		_w36611_,
		_w37007_
	);
	LUT2 #(
		.INIT('h4)
	) name26496 (
		_w36351_,
		_w36613_,
		_w37008_
	);
	LUT2 #(
		.INIT('h4)
	) name26497 (
		_w36133_,
		_w36688_,
		_w37009_
	);
	LUT2 #(
		.INIT('h4)
	) name26498 (
		_w36351_,
		_w36617_,
		_w37010_
	);
	LUT2 #(
		.INIT('h4)
	) name26499 (
		_w36351_,
		_w36619_,
		_w37011_
	);
	LUT2 #(
		.INIT('h4)
	) name26500 (
		_w36351_,
		_w36621_,
		_w37012_
	);
	LUT2 #(
		.INIT('h4)
	) name26501 (
		_w36351_,
		_w36623_,
		_w37013_
	);
	LUT2 #(
		.INIT('h4)
	) name26502 (
		_w36351_,
		_w36625_,
		_w37014_
	);
	LUT2 #(
		.INIT('h4)
	) name26503 (
		_w36351_,
		_w36627_,
		_w37015_
	);
	LUT2 #(
		.INIT('h4)
	) name26504 (
		_w36351_,
		_w36629_,
		_w37016_
	);
	LUT2 #(
		.INIT('h4)
	) name26505 (
		_w36351_,
		_w36631_,
		_w37017_
	);
	LUT2 #(
		.INIT('h4)
	) name26506 (
		_w36351_,
		_w36633_,
		_w37018_
	);
	LUT2 #(
		.INIT('h4)
	) name26507 (
		_w36351_,
		_w36635_,
		_w37019_
	);
	LUT2 #(
		.INIT('h4)
	) name26508 (
		_w36351_,
		_w36637_,
		_w37020_
	);
	LUT2 #(
		.INIT('h4)
	) name26509 (
		_w36351_,
		_w36639_,
		_w37021_
	);
	LUT2 #(
		.INIT('h4)
	) name26510 (
		_w36133_,
		_w36692_,
		_w37022_
	);
	LUT2 #(
		.INIT('h4)
	) name26511 (
		_w36351_,
		_w36641_,
		_w37023_
	);
	LUT2 #(
		.INIT('h4)
	) name26512 (
		_w36351_,
		_w36643_,
		_w37024_
	);
	LUT2 #(
		.INIT('h4)
	) name26513 (
		_w36351_,
		_w36645_,
		_w37025_
	);
	LUT2 #(
		.INIT('h4)
	) name26514 (
		_w36133_,
		_w36694_,
		_w37026_
	);
	LUT2 #(
		.INIT('h4)
	) name26515 (
		_w36351_,
		_w36647_,
		_w37027_
	);
	LUT2 #(
		.INIT('h4)
	) name26516 (
		_w36351_,
		_w36649_,
		_w37028_
	);
	LUT2 #(
		.INIT('h4)
	) name26517 (
		_w36351_,
		_w36651_,
		_w37029_
	);
	LUT2 #(
		.INIT('h4)
	) name26518 (
		_w36133_,
		_w36917_,
		_w37030_
	);
	LUT2 #(
		.INIT('h4)
	) name26519 (
		_w36133_,
		_w36696_,
		_w37031_
	);
	LUT2 #(
		.INIT('h4)
	) name26520 (
		_w36101_,
		_w36608_,
		_w37032_
	);
	LUT2 #(
		.INIT('h4)
	) name26521 (
		_w36351_,
		_w36653_,
		_w37033_
	);
	LUT2 #(
		.INIT('h4)
	) name26522 (
		_w36351_,
		_w36655_,
		_w37034_
	);
	LUT2 #(
		.INIT('h4)
	) name26523 (
		_w36133_,
		_w36698_,
		_w37035_
	);
	LUT2 #(
		.INIT('h4)
	) name26524 (
		_w36351_,
		_w36657_,
		_w37036_
	);
	LUT2 #(
		.INIT('h4)
	) name26525 (
		_w36351_,
		_w36659_,
		_w37037_
	);
	LUT2 #(
		.INIT('h4)
	) name26526 (
		_w36351_,
		_w36663_,
		_w37038_
	);
	LUT2 #(
		.INIT('h4)
	) name26527 (
		_w36133_,
		_w36701_,
		_w37039_
	);
	LUT2 #(
		.INIT('h4)
	) name26528 (
		_w36351_,
		_w36665_,
		_w37040_
	);
	LUT2 #(
		.INIT('h4)
	) name26529 (
		_w36133_,
		_w36703_,
		_w37041_
	);
	LUT2 #(
		.INIT('h4)
	) name26530 (
		_w36351_,
		_w36668_,
		_w37042_
	);
	LUT2 #(
		.INIT('h4)
	) name26531 (
		_w36351_,
		_w36670_,
		_w37043_
	);
	LUT2 #(
		.INIT('h4)
	) name26532 (
		_w36351_,
		_w36673_,
		_w37044_
	);
	LUT2 #(
		.INIT('h4)
	) name26533 (
		_w36351_,
		_w36675_,
		_w37045_
	);
	LUT2 #(
		.INIT('h4)
	) name26534 (
		_w36133_,
		_w36706_,
		_w37046_
	);
	LUT2 #(
		.INIT('h4)
	) name26535 (
		_w36133_,
		_w36708_,
		_w37047_
	);
	LUT2 #(
		.INIT('h4)
	) name26536 (
		_w36351_,
		_w36677_,
		_w37048_
	);
	LUT2 #(
		.INIT('h4)
	) name26537 (
		_w36351_,
		_w36679_,
		_w37049_
	);
	LUT2 #(
		.INIT('h4)
	) name26538 (
		_w36351_,
		_w36681_,
		_w37050_
	);
	LUT2 #(
		.INIT('h4)
	) name26539 (
		_w36133_,
		_w36713_,
		_w37051_
	);
	LUT2 #(
		.INIT('h4)
	) name26540 (
		_w36351_,
		_w36684_,
		_w37052_
	);
	LUT2 #(
		.INIT('h4)
	) name26541 (
		_w36351_,
		_w36686_,
		_w37053_
	);
	LUT2 #(
		.INIT('h4)
	) name26542 (
		_w36351_,
		_w36688_,
		_w37054_
	);
	LUT2 #(
		.INIT('h4)
	) name26543 (
		_w36133_,
		_w36715_,
		_w37055_
	);
	LUT2 #(
		.INIT('h4)
	) name26544 (
		_w36133_,
		_w36717_,
		_w37056_
	);
	LUT2 #(
		.INIT('h4)
	) name26545 (
		_w36351_,
		_w36692_,
		_w37057_
	);
	LUT2 #(
		.INIT('h4)
	) name26546 (
		_w36133_,
		_w36719_,
		_w37058_
	);
	LUT2 #(
		.INIT('h4)
	) name26547 (
		_w36351_,
		_w36694_,
		_w37059_
	);
	LUT2 #(
		.INIT('h4)
	) name26548 (
		_w36133_,
		_w36721_,
		_w37060_
	);
	LUT2 #(
		.INIT('h4)
	) name26549 (
		_w36351_,
		_w36696_,
		_w37061_
	);
	LUT2 #(
		.INIT('h4)
	) name26550 (
		_w36133_,
		_w36723_,
		_w37062_
	);
	LUT2 #(
		.INIT('h4)
	) name26551 (
		_w36351_,
		_w36698_,
		_w37063_
	);
	LUT2 #(
		.INIT('h4)
	) name26552 (
		_w36133_,
		_w36725_,
		_w37064_
	);
	LUT2 #(
		.INIT('h4)
	) name26553 (
		_w36351_,
		_w36701_,
		_w37065_
	);
	LUT2 #(
		.INIT('h4)
	) name26554 (
		_w36133_,
		_w36728_,
		_w37066_
	);
	LUT2 #(
		.INIT('h4)
	) name26555 (
		_w36351_,
		_w36703_,
		_w37067_
	);
	LUT2 #(
		.INIT('h4)
	) name26556 (
		_w36133_,
		_w36730_,
		_w37068_
	);
	LUT2 #(
		.INIT('h4)
	) name26557 (
		_w36351_,
		_w36706_,
		_w37069_
	);
	LUT2 #(
		.INIT('h4)
	) name26558 (
		_w36133_,
		_w36732_,
		_w37070_
	);
	LUT2 #(
		.INIT('h4)
	) name26559 (
		_w36351_,
		_w36708_,
		_w37071_
	);
	LUT2 #(
		.INIT('h4)
	) name26560 (
		_w36133_,
		_w36734_,
		_w37072_
	);
	LUT2 #(
		.INIT('h4)
	) name26561 (
		_w36351_,
		_w36713_,
		_w37073_
	);
	LUT2 #(
		.INIT('h4)
	) name26562 (
		_w36133_,
		_w36736_,
		_w37074_
	);
	LUT2 #(
		.INIT('h4)
	) name26563 (
		_w36351_,
		_w36715_,
		_w37075_
	);
	LUT2 #(
		.INIT('h4)
	) name26564 (
		_w36133_,
		_w36738_,
		_w37076_
	);
	LUT2 #(
		.INIT('h4)
	) name26565 (
		_w36351_,
		_w36717_,
		_w37077_
	);
	LUT2 #(
		.INIT('h4)
	) name26566 (
		_w36351_,
		_w36719_,
		_w37078_
	);
	LUT2 #(
		.INIT('h4)
	) name26567 (
		_w36351_,
		_w36721_,
		_w37079_
	);
	LUT2 #(
		.INIT('h4)
	) name26568 (
		_w36351_,
		_w36723_,
		_w37080_
	);
	LUT2 #(
		.INIT('h4)
	) name26569 (
		_w36133_,
		_w36740_,
		_w37081_
	);
	LUT2 #(
		.INIT('h4)
	) name26570 (
		_w36351_,
		_w36725_,
		_w37082_
	);
	LUT2 #(
		.INIT('h4)
	) name26571 (
		_w36351_,
		_w36728_,
		_w37083_
	);
	LUT2 #(
		.INIT('h4)
	) name26572 (
		_w36351_,
		_w36730_,
		_w37084_
	);
	LUT2 #(
		.INIT('h4)
	) name26573 (
		_w36351_,
		_w36732_,
		_w37085_
	);
	LUT2 #(
		.INIT('h4)
	) name26574 (
		_w36351_,
		_w36734_,
		_w37086_
	);
	LUT2 #(
		.INIT('h4)
	) name26575 (
		_w36351_,
		_w36736_,
		_w37087_
	);
	LUT2 #(
		.INIT('h4)
	) name26576 (
		_w36133_,
		_w36742_,
		_w37088_
	);
	LUT2 #(
		.INIT('h4)
	) name26577 (
		_w36351_,
		_w36738_,
		_w37089_
	);
	LUT2 #(
		.INIT('h4)
	) name26578 (
		_w36133_,
		_w36744_,
		_w37090_
	);
	LUT2 #(
		.INIT('h4)
	) name26579 (
		_w36351_,
		_w36740_,
		_w37091_
	);
	LUT2 #(
		.INIT('h4)
	) name26580 (
		_w36133_,
		_w36746_,
		_w37092_
	);
	LUT2 #(
		.INIT('h4)
	) name26581 (
		_w36351_,
		_w36742_,
		_w37093_
	);
	LUT2 #(
		.INIT('h4)
	) name26582 (
		_w36133_,
		_w36748_,
		_w37094_
	);
	LUT2 #(
		.INIT('h4)
	) name26583 (
		_w36351_,
		_w36744_,
		_w37095_
	);
	LUT2 #(
		.INIT('h4)
	) name26584 (
		_w36351_,
		_w36746_,
		_w37096_
	);
	LUT2 #(
		.INIT('h4)
	) name26585 (
		_w36351_,
		_w36748_,
		_w37097_
	);
	LUT2 #(
		.INIT('h4)
	) name26586 (
		_w36351_,
		_w36751_,
		_w37098_
	);
	LUT2 #(
		.INIT('h4)
	) name26587 (
		_w36133_,
		_w36751_,
		_w37099_
	);
	LUT2 #(
		.INIT('h4)
	) name26588 (
		_w36351_,
		_w36753_,
		_w37100_
	);
	LUT2 #(
		.INIT('h4)
	) name26589 (
		_w36351_,
		_w36755_,
		_w37101_
	);
	LUT2 #(
		.INIT('h4)
	) name26590 (
		_w36351_,
		_w36757_,
		_w37102_
	);
	LUT2 #(
		.INIT('h4)
	) name26591 (
		_w36351_,
		_w36759_,
		_w37103_
	);
	LUT2 #(
		.INIT('h4)
	) name26592 (
		_w36133_,
		_w36753_,
		_w37104_
	);
	LUT2 #(
		.INIT('h4)
	) name26593 (
		_w36351_,
		_w36956_,
		_w37105_
	);
	LUT2 #(
		.INIT('h4)
	) name26594 (
		_w36351_,
		_w36761_,
		_w37106_
	);
	LUT2 #(
		.INIT('h4)
	) name26595 (
		_w36133_,
		_w36755_,
		_w37107_
	);
	LUT2 #(
		.INIT('h4)
	) name26596 (
		_w36351_,
		_w36763_,
		_w37108_
	);
	LUT2 #(
		.INIT('h4)
	) name26597 (
		_w36133_,
		_w36757_,
		_w37109_
	);
	LUT2 #(
		.INIT('h4)
	) name26598 (
		_w36351_,
		_w36765_,
		_w37110_
	);
	LUT2 #(
		.INIT('h4)
	) name26599 (
		_w36133_,
		_w36759_,
		_w37111_
	);
	LUT2 #(
		.INIT('h4)
	) name26600 (
		_w36351_,
		_w36767_,
		_w37112_
	);
	LUT2 #(
		.INIT('h4)
	) name26601 (
		_w36351_,
		_w36769_,
		_w37113_
	);
	LUT2 #(
		.INIT('h4)
	) name26602 (
		_w36133_,
		_w36911_,
		_w37114_
	);
	LUT2 #(
		.INIT('h4)
	) name26603 (
		_w36133_,
		_w36761_,
		_w37115_
	);
	LUT2 #(
		.INIT('h4)
	) name26604 (
		_w36351_,
		_w36773_,
		_w37116_
	);
	LUT2 #(
		.INIT('h4)
	) name26605 (
		_w36351_,
		_w36775_,
		_w37117_
	);
	LUT2 #(
		.INIT('h4)
	) name26606 (
		_w36351_,
		_w36777_,
		_w37118_
	);
	LUT2 #(
		.INIT('h4)
	) name26607 (
		_w36351_,
		_w36779_,
		_w37119_
	);
	LUT2 #(
		.INIT('h4)
	) name26608 (
		_w36133_,
		_w36763_,
		_w37120_
	);
	LUT2 #(
		.INIT('h4)
	) name26609 (
		_w36351_,
		_w36781_,
		_w37121_
	);
	LUT2 #(
		.INIT('h4)
	) name26610 (
		_w36133_,
		_w36852_,
		_w37122_
	);
	LUT2 #(
		.INIT('h4)
	) name26611 (
		_w36351_,
		_w36784_,
		_w37123_
	);
	LUT2 #(
		.INIT('h4)
	) name26612 (
		_w36351_,
		_w36786_,
		_w37124_
	);
	LUT2 #(
		.INIT('h4)
	) name26613 (
		_w36351_,
		_w36788_,
		_w37125_
	);
	LUT2 #(
		.INIT('h4)
	) name26614 (
		_w36133_,
		_w36765_,
		_w37126_
	);
	LUT2 #(
		.INIT('h4)
	) name26615 (
		_w36351_,
		_w36953_,
		_w37127_
	);
	LUT2 #(
		.INIT('h4)
	) name26616 (
		_w36133_,
		_w36767_,
		_w37128_
	);
	LUT2 #(
		.INIT('h4)
	) name26617 (
		_w36351_,
		_w36791_,
		_w37129_
	);
	LUT2 #(
		.INIT('h4)
	) name26618 (
		_w36133_,
		_w36769_,
		_w37130_
	);
	LUT2 #(
		.INIT('h4)
	) name26619 (
		_w36351_,
		_w36793_,
		_w37131_
	);
	LUT2 #(
		.INIT('h4)
	) name26620 (
		_w36351_,
		_w36795_,
		_w37132_
	);
	LUT2 #(
		.INIT('h4)
	) name26621 (
		_w36351_,
		_w36798_,
		_w37133_
	);
	LUT2 #(
		.INIT('h4)
	) name26622 (
		_w36351_,
		_w36801_,
		_w37134_
	);
	LUT2 #(
		.INIT('h4)
	) name26623 (
		_w36133_,
		_w36773_,
		_w37135_
	);
	LUT2 #(
		.INIT('h4)
	) name26624 (
		_w36351_,
		_w36803_,
		_w37136_
	);
	LUT2 #(
		.INIT('h4)
	) name26625 (
		_w36351_,
		_w36805_,
		_w37137_
	);
	LUT2 #(
		.INIT('h4)
	) name26626 (
		_w36133_,
		_w36775_,
		_w37138_
	);
	LUT2 #(
		.INIT('h4)
	) name26627 (
		_w36351_,
		_w36807_,
		_w37139_
	);
	LUT2 #(
		.INIT('h4)
	) name26628 (
		_w36351_,
		_w36809_,
		_w37140_
	);
	LUT2 #(
		.INIT('h4)
	) name26629 (
		_w36133_,
		_w36777_,
		_w37141_
	);
	LUT2 #(
		.INIT('h4)
	) name26630 (
		_w36351_,
		_w36811_,
		_w37142_
	);
	LUT2 #(
		.INIT('h4)
	) name26631 (
		_w36351_,
		_w36814_,
		_w37143_
	);
	LUT2 #(
		.INIT('h4)
	) name26632 (
		_w36133_,
		_w36779_,
		_w37144_
	);
	LUT2 #(
		.INIT('h4)
	) name26633 (
		_w36133_,
		_w36781_,
		_w37145_
	);
	LUT2 #(
		.INIT('h4)
	) name26634 (
		_w36351_,
		_w36818_,
		_w37146_
	);
	LUT2 #(
		.INIT('h4)
	) name26635 (
		_w36351_,
		_w36821_,
		_w37147_
	);
	LUT2 #(
		.INIT('h4)
	) name26636 (
		_w36133_,
		_w36953_,
		_w37148_
	);
	LUT2 #(
		.INIT('h4)
	) name26637 (
		_w36133_,
		_w36784_,
		_w37149_
	);
	LUT2 #(
		.INIT('h4)
	) name26638 (
		_w36351_,
		_w36823_,
		_w37150_
	);
	LUT2 #(
		.INIT('h4)
	) name26639 (
		_w36351_,
		_w36826_,
		_w37151_
	);
	LUT2 #(
		.INIT('h4)
	) name26640 (
		_w36133_,
		_w36786_,
		_w37152_
	);
	LUT2 #(
		.INIT('h4)
	) name26641 (
		_w36351_,
		_w36828_,
		_w37153_
	);
	LUT2 #(
		.INIT('h4)
	) name26642 (
		_w36351_,
		_w36831_,
		_w37154_
	);
	LUT2 #(
		.INIT('h4)
	) name26643 (
		_w36133_,
		_w36788_,
		_w37155_
	);
	LUT2 #(
		.INIT('h4)
	) name26644 (
		_w36351_,
		_w36833_,
		_w37156_
	);
	LUT2 #(
		.INIT('h4)
	) name26645 (
		_w36351_,
		_w36836_,
		_w37157_
	);
	LUT2 #(
		.INIT('h4)
	) name26646 (
		_w36351_,
		_w36838_,
		_w37158_
	);
	LUT2 #(
		.INIT('h4)
	) name26647 (
		_w36351_,
		_w36841_,
		_w37159_
	);
	LUT2 #(
		.INIT('h4)
	) name26648 (
		_w36351_,
		_w36843_,
		_w37160_
	);
	LUT2 #(
		.INIT('h4)
	) name26649 (
		_w36351_,
		_w36845_,
		_w37161_
	);
	LUT2 #(
		.INIT('h4)
	) name26650 (
		_w36133_,
		_w36791_,
		_w37162_
	);
	LUT2 #(
		.INIT('h4)
	) name26651 (
		_w36351_,
		_w36847_,
		_w37163_
	);
	LUT2 #(
		.INIT('h4)
	) name26652 (
		_w36351_,
		_w36849_,
		_w37164_
	);
	LUT2 #(
		.INIT('h4)
	) name26653 (
		_w36351_,
		_w36852_,
		_w37165_
	);
	LUT2 #(
		.INIT('h4)
	) name26654 (
		_w36351_,
		_w36855_,
		_w37166_
	);
	LUT2 #(
		.INIT('h4)
	) name26655 (
		_w36133_,
		_w36793_,
		_w37167_
	);
	LUT2 #(
		.INIT('h4)
	) name26656 (
		_w36351_,
		_w36857_,
		_w37168_
	);
	LUT2 #(
		.INIT('h4)
	) name26657 (
		_w36133_,
		_w36795_,
		_w37169_
	);
	LUT2 #(
		.INIT('h4)
	) name26658 (
		_w36351_,
		_w36860_,
		_w37170_
	);
	LUT2 #(
		.INIT('h4)
	) name26659 (
		_w36351_,
		_w36862_,
		_w37171_
	);
	LUT2 #(
		.INIT('h4)
	) name26660 (
		_w36133_,
		_w36798_,
		_w37172_
	);
	LUT2 #(
		.INIT('h4)
	) name26661 (
		_w36351_,
		_w36866_,
		_w37173_
	);
	LUT2 #(
		.INIT('h4)
	) name26662 (
		_w36351_,
		_w36868_,
		_w37174_
	);
	LUT2 #(
		.INIT('h4)
	) name26663 (
		_w36351_,
		_w36871_,
		_w37175_
	);
	LUT2 #(
		.INIT('h4)
	) name26664 (
		_w36351_,
		_w36873_,
		_w37176_
	);
	LUT2 #(
		.INIT('h4)
	) name26665 (
		_w36133_,
		_w36801_,
		_w37177_
	);
	LUT2 #(
		.INIT('h4)
	) name26666 (
		_w36351_,
		_w36875_,
		_w37178_
	);
	LUT2 #(
		.INIT('h4)
	) name26667 (
		_w36351_,
		_w36877_,
		_w37179_
	);
	LUT2 #(
		.INIT('h4)
	) name26668 (
		_w36133_,
		_w36803_,
		_w37180_
	);
	LUT2 #(
		.INIT('h4)
	) name26669 (
		_w36351_,
		_w36879_,
		_w37181_
	);
	LUT2 #(
		.INIT('h4)
	) name26670 (
		_w36133_,
		_w36805_,
		_w37182_
	);
	LUT2 #(
		.INIT('h4)
	) name26671 (
		_w36351_,
		_w36882_,
		_w37183_
	);
	LUT2 #(
		.INIT('h4)
	) name26672 (
		_w36133_,
		_w36807_,
		_w37184_
	);
	LUT2 #(
		.INIT('h4)
	) name26673 (
		_w36351_,
		_w36884_,
		_w37185_
	);
	LUT2 #(
		.INIT('h4)
	) name26674 (
		_w36351_,
		_w36887_,
		_w37186_
	);
	LUT2 #(
		.INIT('h4)
	) name26675 (
		_w36133_,
		_w36809_,
		_w37187_
	);
	LUT2 #(
		.INIT('h4)
	) name26676 (
		_w36351_,
		_w36889_,
		_w37188_
	);
	LUT2 #(
		.INIT('h4)
	) name26677 (
		_w36133_,
		_w36811_,
		_w37189_
	);
	LUT2 #(
		.INIT('h4)
	) name26678 (
		_w36351_,
		_w36940_,
		_w37190_
	);
	LUT2 #(
		.INIT('h4)
	) name26679 (
		_w36351_,
		_w36615_,
		_w37191_
	);
	LUT2 #(
		.INIT('h4)
	) name26680 (
		_w36133_,
		_w36814_,
		_w37192_
	);
	LUT2 #(
		.INIT('h4)
	) name26681 (
		_w36351_,
		_w36895_,
		_w37193_
	);
	LUT2 #(
		.INIT('h4)
	) name26682 (
		_w36351_,
		_w36897_,
		_w37194_
	);
	LUT2 #(
		.INIT('h4)
	) name26683 (
		_w36351_,
		_w36938_,
		_w37195_
	);
	LUT2 #(
		.INIT('h4)
	) name26684 (
		_w36351_,
		_w36900_,
		_w37196_
	);
	LUT2 #(
		.INIT('h4)
	) name26685 (
		_w36351_,
		_w36902_,
		_w37197_
	);
	LUT2 #(
		.INIT('h4)
	) name26686 (
		_w36351_,
		_w36905_,
		_w37198_
	);
	LUT2 #(
		.INIT('h4)
	) name26687 (
		_w36133_,
		_w36818_,
		_w37199_
	);
	LUT2 #(
		.INIT('h4)
	) name26688 (
		_w36351_,
		_w36908_,
		_w37200_
	);
	LUT2 #(
		.INIT('h4)
	) name26689 (
		_w36351_,
		_w36935_,
		_w37201_
	);
	LUT2 #(
		.INIT('h4)
	) name26690 (
		_w36133_,
		_w36821_,
		_w37202_
	);
	LUT2 #(
		.INIT('h4)
	) name26691 (
		_w36133_,
		_w36823_,
		_w37203_
	);
	LUT2 #(
		.INIT('h4)
	) name26692 (
		_w36351_,
		_w36911_,
		_w37204_
	);
	LUT2 #(
		.INIT('h4)
	) name26693 (
		_w36351_,
		_w36914_,
		_w37205_
	);
	LUT2 #(
		.INIT('h4)
	) name26694 (
		_w36133_,
		_w36826_,
		_w37206_
	);
	LUT2 #(
		.INIT('h4)
	) name26695 (
		_w36133_,
		_w36828_,
		_w37207_
	);
	LUT2 #(
		.INIT('h4)
	) name26696 (
		_w36351_,
		_w36917_,
		_w37208_
	);
	LUT2 #(
		.INIT('h4)
	) name26697 (
		_w36351_,
		_w36920_,
		_w37209_
	);
	LUT2 #(
		.INIT('h4)
	) name26698 (
		_w36133_,
		_w36831_,
		_w37210_
	);
	LUT2 #(
		.INIT('h4)
	) name26699 (
		_w36351_,
		_w36923_,
		_w37211_
	);
	LUT2 #(
		.INIT('h4)
	) name26700 (
		_w36351_,
		_w36933_,
		_w37212_
	);
	LUT2 #(
		.INIT('h4)
	) name26701 (
		_w36133_,
		_w36833_,
		_w37213_
	);
	LUT2 #(
		.INIT('h4)
	) name26702 (
		_w36351_,
		_w36925_,
		_w37214_
	);
	LUT2 #(
		.INIT('h4)
	) name26703 (
		_w36351_,
		_w36927_,
		_w37215_
	);
	LUT2 #(
		.INIT('h4)
	) name26704 (
		_w36133_,
		_w36836_,
		_w37216_
	);
	LUT2 #(
		.INIT('h4)
	) name26705 (
		_w36351_,
		_w36711_,
		_w37217_
	);
	LUT2 #(
		.INIT('h4)
	) name26706 (
		_w36351_,
		_w36930_,
		_w37218_
	);
	LUT2 #(
		.INIT('h4)
	) name26707 (
		_w36133_,
		_w36838_,
		_w37219_
	);
	LUT2 #(
		.INIT('h4)
	) name26708 (
		_w36133_,
		_w36841_,
		_w37220_
	);
	LUT2 #(
		.INIT('h4)
	) name26709 (
		_w36133_,
		_w36843_,
		_w37221_
	);
	LUT2 #(
		.INIT('h4)
	) name26710 (
		_w36351_,
		_w36943_,
		_w37222_
	);
	LUT2 #(
		.INIT('h4)
	) name26711 (
		_w36351_,
		_w36945_,
		_w37223_
	);
	LUT2 #(
		.INIT('h4)
	) name26712 (
		_w36133_,
		_w36845_,
		_w37224_
	);
	LUT2 #(
		.INIT('h4)
	) name26713 (
		_w36351_,
		_w36948_,
		_w37225_
	);
	LUT2 #(
		.INIT('h4)
	) name26714 (
		_w36133_,
		_w36847_,
		_w37226_
	);
	LUT2 #(
		.INIT('h4)
	) name26715 (
		_w36351_,
		_w36950_,
		_w37227_
	);
	LUT2 #(
		.INIT('h4)
	) name26716 (
		_w36133_,
		_w36849_,
		_w37228_
	);
	LUT2 #(
		.INIT('h4)
	) name26717 (
		_w36133_,
		_w36855_,
		_w37229_
	);
	LUT2 #(
		.INIT('h4)
	) name26718 (
		_w36351_,
		_w36816_,
		_w37230_
	);
	LUT2 #(
		.INIT('h4)
	) name26719 (
		_w36351_,
		_w36959_,
		_w37231_
	);
	LUT2 #(
		.INIT('h4)
	) name26720 (
		_w36133_,
		_w36857_,
		_w37232_
	);
	LUT2 #(
		.INIT('h4)
	) name26721 (
		_w36351_,
		_w36771_,
		_w37233_
	);
	LUT2 #(
		.INIT('h4)
	) name26722 (
		_w36351_,
		_w36964_,
		_w37234_
	);
	LUT2 #(
		.INIT('h4)
	) name26723 (
		_w36133_,
		_w36860_,
		_w37235_
	);
	LUT2 #(
		.INIT('h4)
	) name26724 (
		_w36351_,
		_w36969_,
		_w37236_
	);
	LUT2 #(
		.INIT('h4)
	) name26725 (
		_w36351_,
		_w36972_,
		_w37237_
	);
	LUT2 #(
		.INIT('h4)
	) name26726 (
		_w36133_,
		_w36862_,
		_w37238_
	);
	LUT2 #(
		.INIT('h4)
	) name26727 (
		_w36133_,
		_w36866_,
		_w37239_
	);
	LUT2 #(
		.INIT('h4)
	) name26728 (
		_w36133_,
		_w36868_,
		_w37240_
	);
	LUT2 #(
		.INIT('h4)
	) name26729 (
		_w36351_,
		_w36980_,
		_w37241_
	);
	LUT2 #(
		.INIT('h4)
	) name26730 (
		_w36351_,
		_w36982_,
		_w37242_
	);
	LUT2 #(
		.INIT('h4)
	) name26731 (
		_w36133_,
		_w36871_,
		_w37243_
	);
	LUT2 #(
		.INIT('h4)
	) name26732 (
		_w36351_,
		_w36984_,
		_w37244_
	);
	LUT2 #(
		.INIT('h4)
	) name26733 (
		_w36133_,
		_w36873_,
		_w37245_
	);
	LUT2 #(
		.INIT('h4)
	) name26734 (
		_w36351_,
		_w36586_,
		_w37246_
	);
	LUT2 #(
		.INIT('h4)
	) name26735 (
		_w36133_,
		_w36875_,
		_w37247_
	);
	LUT2 #(
		.INIT('h4)
	) name26736 (
		_w36133_,
		_w36877_,
		_w37248_
	);
	LUT2 #(
		.INIT('h4)
	) name26737 (
		_w36133_,
		_w36972_,
		_w37249_
	);
	LUT2 #(
		.INIT('h4)
	) name26738 (
		_w36101_,
		_w36604_,
		_w37250_
	);
	LUT2 #(
		.INIT('h4)
	) name26739 (
		_w36133_,
		_w36879_,
		_w37251_
	);
	LUT2 #(
		.INIT('h4)
	) name26740 (
		_w36101_,
		_w36602_,
		_w37252_
	);
	LUT2 #(
		.INIT('h4)
	) name26741 (
		_w36101_,
		_w36621_,
		_w37253_
	);
	LUT2 #(
		.INIT('h4)
	) name26742 (
		_w36133_,
		_w36882_,
		_w37254_
	);
	LUT2 #(
		.INIT('h4)
	) name26743 (
		_w36133_,
		_w36884_,
		_w37255_
	);
	LUT2 #(
		.INIT('h4)
	) name26744 (
		_w36101_,
		_w36649_,
		_w37256_
	);
	LUT2 #(
		.INIT('h4)
	) name26745 (
		_w36133_,
		_w36887_,
		_w37257_
	);
	LUT2 #(
		.INIT('h4)
	) name26746 (
		_w36133_,
		_w36889_,
		_w37258_
	);
	LUT2 #(
		.INIT('h4)
	) name26747 (
		_w36133_,
		_w36895_,
		_w37259_
	);
	LUT2 #(
		.INIT('h4)
	) name26748 (
		_w36133_,
		_w36897_,
		_w37260_
	);
	LUT2 #(
		.INIT('h4)
	) name26749 (
		_w36133_,
		_w36900_,
		_w37261_
	);
	LUT2 #(
		.INIT('h4)
	) name26750 (
		_w36133_,
		_w36902_,
		_w37262_
	);
	LUT2 #(
		.INIT('h4)
	) name26751 (
		_w36133_,
		_w36905_,
		_w37263_
	);
	LUT2 #(
		.INIT('h4)
	) name26752 (
		_w36133_,
		_w36908_,
		_w37264_
	);
	LUT2 #(
		.INIT('h4)
	) name26753 (
		_w36133_,
		_w36914_,
		_w37265_
	);
	LUT2 #(
		.INIT('h4)
	) name26754 (
		_w36101_,
		_w36594_,
		_w37266_
	);
	LUT2 #(
		.INIT('h4)
	) name26755 (
		_w36133_,
		_w36925_,
		_w37267_
	);
	LUT2 #(
		.INIT('h4)
	) name26756 (
		_w36133_,
		_w36927_,
		_w37268_
	);
	LUT2 #(
		.INIT('h4)
	) name26757 (
		_w36133_,
		_w36930_,
		_w37269_
	);
	LUT2 #(
		.INIT('h4)
	) name26758 (
		_w36133_,
		_w36933_,
		_w37270_
	);
	LUT2 #(
		.INIT('h4)
	) name26759 (
		_w36133_,
		_w36935_,
		_w37271_
	);
	LUT2 #(
		.INIT('h4)
	) name26760 (
		_w36133_,
		_w36938_,
		_w37272_
	);
	LUT2 #(
		.INIT('h4)
	) name26761 (
		_w36133_,
		_w36940_,
		_w37273_
	);
	LUT2 #(
		.INIT('h4)
	) name26762 (
		_w36133_,
		_w36943_,
		_w37274_
	);
	LUT2 #(
		.INIT('h4)
	) name26763 (
		_w36133_,
		_w36945_,
		_w37275_
	);
	LUT2 #(
		.INIT('h4)
	) name26764 (
		_w36133_,
		_w36948_,
		_w37276_
	);
	LUT2 #(
		.INIT('h4)
	) name26765 (
		_w36133_,
		_w36950_,
		_w37277_
	);
	LUT2 #(
		.INIT('h4)
	) name26766 (
		_w36133_,
		_w36956_,
		_w37278_
	);
	LUT2 #(
		.INIT('h4)
	) name26767 (
		_w36133_,
		_w36959_,
		_w37279_
	);
	LUT2 #(
		.INIT('h4)
	) name26768 (
		_w36133_,
		_w36964_,
		_w37280_
	);
	LUT2 #(
		.INIT('h4)
	) name26769 (
		_w36133_,
		_w36969_,
		_w37281_
	);
	LUT2 #(
		.INIT('h4)
	) name26770 (
		_w36101_,
		_w36613_,
		_w37282_
	);
	LUT2 #(
		.INIT('h4)
	) name26771 (
		_w36133_,
		_w36975_,
		_w37283_
	);
	LUT2 #(
		.INIT('h4)
	) name26772 (
		_w36133_,
		_w36966_,
		_w37284_
	);
	LUT2 #(
		.INIT('h4)
	) name26773 (
		_w36101_,
		_w36611_,
		_w37285_
	);
	LUT2 #(
		.INIT('h4)
	) name26774 (
		_w36133_,
		_w36980_,
		_w37286_
	);
	LUT2 #(
		.INIT('h4)
	) name26775 (
		_w36133_,
		_w36982_,
		_w37287_
	);
	LUT2 #(
		.INIT('h4)
	) name26776 (
		_w36133_,
		_w36984_,
		_w37288_
	);
	LUT2 #(
		.INIT('h4)
	) name26777 (
		_w36133_,
		_w36586_,
		_w37289_
	);
	LUT2 #(
		.INIT('h4)
	) name26778 (
		_w36101_,
		_w36590_,
		_w37290_
	);
	LUT2 #(
		.INIT('h4)
	) name26779 (
		_w36101_,
		_w36596_,
		_w37291_
	);
	LUT2 #(
		.INIT('h4)
	) name26780 (
		_w36101_,
		_w36598_,
		_w37292_
	);
	LUT2 #(
		.INIT('h4)
	) name26781 (
		_w36101_,
		_w36600_,
		_w37293_
	);
	LUT2 #(
		.INIT('h4)
	) name26782 (
		_w36101_,
		_w36606_,
		_w37294_
	);
	LUT2 #(
		.INIT('h4)
	) name26783 (
		_w36101_,
		_w36617_,
		_w37295_
	);
	LUT2 #(
		.INIT('h4)
	) name26784 (
		_w36101_,
		_w36619_,
		_w37296_
	);
	LUT2 #(
		.INIT('h4)
	) name26785 (
		_w36101_,
		_w36623_,
		_w37297_
	);
	LUT2 #(
		.INIT('h4)
	) name26786 (
		_w36101_,
		_w36641_,
		_w37298_
	);
	LUT2 #(
		.INIT('h4)
	) name26787 (
		_w36101_,
		_w36655_,
		_w37299_
	);
	LUT2 #(
		.INIT('h4)
	) name26788 (
		_w36101_,
		_w36657_,
		_w37300_
	);
	LUT2 #(
		.INIT('h4)
	) name26789 (
		_w36101_,
		_w36659_,
		_w37301_
	);
	LUT2 #(
		.INIT('h4)
	) name26790 (
		_w36101_,
		_w36663_,
		_w37302_
	);
	LUT2 #(
		.INIT('h4)
	) name26791 (
		_w36101_,
		_w36665_,
		_w37303_
	);
	LUT2 #(
		.INIT('h4)
	) name26792 (
		_w36101_,
		_w36668_,
		_w37304_
	);
	LUT2 #(
		.INIT('h4)
	) name26793 (
		_w36101_,
		_w36670_,
		_w37305_
	);
	LUT2 #(
		.INIT('h4)
	) name26794 (
		_w36101_,
		_w36673_,
		_w37306_
	);
	LUT2 #(
		.INIT('h4)
	) name26795 (
		_w36101_,
		_w36675_,
		_w37307_
	);
	LUT2 #(
		.INIT('h4)
	) name26796 (
		_w36101_,
		_w36677_,
		_w37308_
	);
	LUT2 #(
		.INIT('h4)
	) name26797 (
		_w36101_,
		_w36679_,
		_w37309_
	);
	LUT2 #(
		.INIT('h4)
	) name26798 (
		_w36101_,
		_w36681_,
		_w37310_
	);
	LUT2 #(
		.INIT('h4)
	) name26799 (
		_w36101_,
		_w36684_,
		_w37311_
	);
	LUT2 #(
		.INIT('h4)
	) name26800 (
		_w36101_,
		_w36686_,
		_w37312_
	);
	LUT2 #(
		.INIT('h4)
	) name26801 (
		_w36101_,
		_w36688_,
		_w37313_
	);
	LUT2 #(
		.INIT('h4)
	) name26802 (
		_w36101_,
		_w36692_,
		_w37314_
	);
	LUT2 #(
		.INIT('h4)
	) name26803 (
		_w36101_,
		_w36694_,
		_w37315_
	);
	LUT2 #(
		.INIT('h4)
	) name26804 (
		_w36101_,
		_w36696_,
		_w37316_
	);
	LUT2 #(
		.INIT('h4)
	) name26805 (
		_w36101_,
		_w36698_,
		_w37317_
	);
	LUT2 #(
		.INIT('h4)
	) name26806 (
		_w36101_,
		_w36701_,
		_w37318_
	);
	LUT2 #(
		.INIT('h4)
	) name26807 (
		_w36101_,
		_w36703_,
		_w37319_
	);
	LUT2 #(
		.INIT('h4)
	) name26808 (
		_w36101_,
		_w36706_,
		_w37320_
	);
	LUT2 #(
		.INIT('h4)
	) name26809 (
		_w36101_,
		_w36708_,
		_w37321_
	);
	LUT2 #(
		.INIT('h4)
	) name26810 (
		_w36101_,
		_w36713_,
		_w37322_
	);
	LUT2 #(
		.INIT('h4)
	) name26811 (
		_w36101_,
		_w36715_,
		_w37323_
	);
	LUT2 #(
		.INIT('h4)
	) name26812 (
		_w36101_,
		_w36717_,
		_w37324_
	);
	LUT2 #(
		.INIT('h4)
	) name26813 (
		_w36101_,
		_w36719_,
		_w37325_
	);
	LUT2 #(
		.INIT('h4)
	) name26814 (
		_w36101_,
		_w36721_,
		_w37326_
	);
	LUT2 #(
		.INIT('h4)
	) name26815 (
		_w36101_,
		_w36723_,
		_w37327_
	);
	LUT2 #(
		.INIT('h4)
	) name26816 (
		_w36101_,
		_w36725_,
		_w37328_
	);
	LUT2 #(
		.INIT('h4)
	) name26817 (
		_w36101_,
		_w36728_,
		_w37329_
	);
	LUT2 #(
		.INIT('h4)
	) name26818 (
		_w36101_,
		_w36730_,
		_w37330_
	);
	LUT2 #(
		.INIT('h4)
	) name26819 (
		_w36101_,
		_w36732_,
		_w37331_
	);
	LUT2 #(
		.INIT('h4)
	) name26820 (
		_w36101_,
		_w36734_,
		_w37332_
	);
	LUT2 #(
		.INIT('h4)
	) name26821 (
		_w36101_,
		_w36736_,
		_w37333_
	);
	LUT2 #(
		.INIT('h4)
	) name26822 (
		_w36101_,
		_w36738_,
		_w37334_
	);
	LUT2 #(
		.INIT('h4)
	) name26823 (
		_w36101_,
		_w36740_,
		_w37335_
	);
	LUT2 #(
		.INIT('h4)
	) name26824 (
		_w36101_,
		_w36742_,
		_w37336_
	);
	LUT2 #(
		.INIT('h4)
	) name26825 (
		_w36101_,
		_w36744_,
		_w37337_
	);
	LUT2 #(
		.INIT('h4)
	) name26826 (
		_w36101_,
		_w36746_,
		_w37338_
	);
	LUT2 #(
		.INIT('h4)
	) name26827 (
		_w36101_,
		_w36748_,
		_w37339_
	);
	LUT2 #(
		.INIT('h4)
	) name26828 (
		_w36101_,
		_w36751_,
		_w37340_
	);
	LUT2 #(
		.INIT('h4)
	) name26829 (
		_w36101_,
		_w36753_,
		_w37341_
	);
	LUT2 #(
		.INIT('h4)
	) name26830 (
		_w36101_,
		_w36755_,
		_w37342_
	);
	LUT2 #(
		.INIT('h4)
	) name26831 (
		_w36101_,
		_w36757_,
		_w37343_
	);
	LUT2 #(
		.INIT('h4)
	) name26832 (
		_w36101_,
		_w36759_,
		_w37344_
	);
	LUT2 #(
		.INIT('h4)
	) name26833 (
		_w36101_,
		_w36761_,
		_w37345_
	);
	LUT2 #(
		.INIT('h4)
	) name26834 (
		_w36101_,
		_w36763_,
		_w37346_
	);
	LUT2 #(
		.INIT('h4)
	) name26835 (
		_w36101_,
		_w36765_,
		_w37347_
	);
	LUT2 #(
		.INIT('h4)
	) name26836 (
		_w36101_,
		_w36767_,
		_w37348_
	);
	LUT2 #(
		.INIT('h4)
	) name26837 (
		_w36101_,
		_w36769_,
		_w37349_
	);
	LUT2 #(
		.INIT('h4)
	) name26838 (
		_w36101_,
		_w36773_,
		_w37350_
	);
	LUT2 #(
		.INIT('h4)
	) name26839 (
		_w36101_,
		_w36775_,
		_w37351_
	);
	LUT2 #(
		.INIT('h4)
	) name26840 (
		_w36101_,
		_w36777_,
		_w37352_
	);
	LUT2 #(
		.INIT('h4)
	) name26841 (
		_w36101_,
		_w36779_,
		_w37353_
	);
	LUT2 #(
		.INIT('h4)
	) name26842 (
		_w36101_,
		_w36781_,
		_w37354_
	);
	LUT2 #(
		.INIT('h4)
	) name26843 (
		_w36101_,
		_w36784_,
		_w37355_
	);
	LUT2 #(
		.INIT('h4)
	) name26844 (
		_w36101_,
		_w36786_,
		_w37356_
	);
	LUT2 #(
		.INIT('h4)
	) name26845 (
		_w36101_,
		_w36788_,
		_w37357_
	);
	LUT2 #(
		.INIT('h4)
	) name26846 (
		_w36101_,
		_w36791_,
		_w37358_
	);
	LUT2 #(
		.INIT('h4)
	) name26847 (
		_w36101_,
		_w36793_,
		_w37359_
	);
	LUT2 #(
		.INIT('h4)
	) name26848 (
		_w36101_,
		_w36795_,
		_w37360_
	);
	LUT2 #(
		.INIT('h4)
	) name26849 (
		_w36101_,
		_w36798_,
		_w37361_
	);
	LUT2 #(
		.INIT('h4)
	) name26850 (
		_w36101_,
		_w36801_,
		_w37362_
	);
	LUT2 #(
		.INIT('h4)
	) name26851 (
		_w36101_,
		_w36803_,
		_w37363_
	);
	LUT2 #(
		.INIT('h4)
	) name26852 (
		_w36101_,
		_w36805_,
		_w37364_
	);
	LUT2 #(
		.INIT('h4)
	) name26853 (
		_w36101_,
		_w36807_,
		_w37365_
	);
	LUT2 #(
		.INIT('h4)
	) name26854 (
		_w36101_,
		_w36809_,
		_w37366_
	);
	LUT2 #(
		.INIT('h4)
	) name26855 (
		_w36101_,
		_w36811_,
		_w37367_
	);
	LUT2 #(
		.INIT('h4)
	) name26856 (
		_w36101_,
		_w36814_,
		_w37368_
	);
	LUT2 #(
		.INIT('h4)
	) name26857 (
		_w36101_,
		_w36818_,
		_w37369_
	);
	LUT2 #(
		.INIT('h4)
	) name26858 (
		_w36101_,
		_w36821_,
		_w37370_
	);
	LUT2 #(
		.INIT('h4)
	) name26859 (
		_w36101_,
		_w36823_,
		_w37371_
	);
	LUT2 #(
		.INIT('h4)
	) name26860 (
		_w36101_,
		_w36826_,
		_w37372_
	);
	LUT2 #(
		.INIT('h4)
	) name26861 (
		_w36101_,
		_w36828_,
		_w37373_
	);
	LUT2 #(
		.INIT('h4)
	) name26862 (
		_w36101_,
		_w36831_,
		_w37374_
	);
	LUT2 #(
		.INIT('h4)
	) name26863 (
		_w36101_,
		_w36833_,
		_w37375_
	);
	LUT2 #(
		.INIT('h4)
	) name26864 (
		_w36101_,
		_w36836_,
		_w37376_
	);
	LUT2 #(
		.INIT('h4)
	) name26865 (
		_w36101_,
		_w36838_,
		_w37377_
	);
	LUT2 #(
		.INIT('h4)
	) name26866 (
		_w36101_,
		_w36841_,
		_w37378_
	);
	LUT2 #(
		.INIT('h4)
	) name26867 (
		_w36101_,
		_w36843_,
		_w37379_
	);
	LUT2 #(
		.INIT('h4)
	) name26868 (
		_w36101_,
		_w36845_,
		_w37380_
	);
	LUT2 #(
		.INIT('h4)
	) name26869 (
		_w36101_,
		_w36847_,
		_w37381_
	);
	LUT2 #(
		.INIT('h4)
	) name26870 (
		_w36101_,
		_w36849_,
		_w37382_
	);
	LUT2 #(
		.INIT('h4)
	) name26871 (
		_w36101_,
		_w36852_,
		_w37383_
	);
	LUT2 #(
		.INIT('h4)
	) name26872 (
		_w36101_,
		_w36855_,
		_w37384_
	);
	LUT2 #(
		.INIT('h4)
	) name26873 (
		_w36101_,
		_w36857_,
		_w37385_
	);
	LUT2 #(
		.INIT('h4)
	) name26874 (
		_w36101_,
		_w36860_,
		_w37386_
	);
	LUT2 #(
		.INIT('h4)
	) name26875 (
		_w36101_,
		_w36862_,
		_w37387_
	);
	LUT2 #(
		.INIT('h4)
	) name26876 (
		_w36101_,
		_w36866_,
		_w37388_
	);
	LUT2 #(
		.INIT('h4)
	) name26877 (
		_w36101_,
		_w36868_,
		_w37389_
	);
	LUT2 #(
		.INIT('h4)
	) name26878 (
		_w36101_,
		_w36871_,
		_w37390_
	);
	LUT2 #(
		.INIT('h4)
	) name26879 (
		_w36101_,
		_w36873_,
		_w37391_
	);
	LUT2 #(
		.INIT('h4)
	) name26880 (
		_w36101_,
		_w36875_,
		_w37392_
	);
	LUT2 #(
		.INIT('h4)
	) name26881 (
		_w36101_,
		_w36877_,
		_w37393_
	);
	LUT2 #(
		.INIT('h4)
	) name26882 (
		_w36101_,
		_w36879_,
		_w37394_
	);
	LUT2 #(
		.INIT('h4)
	) name26883 (
		_w36101_,
		_w36882_,
		_w37395_
	);
	LUT2 #(
		.INIT('h4)
	) name26884 (
		_w36101_,
		_w36884_,
		_w37396_
	);
	LUT2 #(
		.INIT('h4)
	) name26885 (
		_w36101_,
		_w36887_,
		_w37397_
	);
	LUT2 #(
		.INIT('h4)
	) name26886 (
		_w36101_,
		_w36889_,
		_w37398_
	);
	LUT2 #(
		.INIT('h4)
	) name26887 (
		_w36101_,
		_w36615_,
		_w37399_
	);
	LUT2 #(
		.INIT('h4)
	) name26888 (
		_w36101_,
		_w36895_,
		_w37400_
	);
	LUT2 #(
		.INIT('h4)
	) name26889 (
		_w36101_,
		_w36897_,
		_w37401_
	);
	LUT2 #(
		.INIT('h4)
	) name26890 (
		_w36101_,
		_w36900_,
		_w37402_
	);
	LUT2 #(
		.INIT('h4)
	) name26891 (
		_w36101_,
		_w36902_,
		_w37403_
	);
	LUT2 #(
		.INIT('h4)
	) name26892 (
		_w36101_,
		_w36905_,
		_w37404_
	);
	LUT2 #(
		.INIT('h4)
	) name26893 (
		_w36101_,
		_w36908_,
		_w37405_
	);
	LUT2 #(
		.INIT('h4)
	) name26894 (
		_w36101_,
		_w36911_,
		_w37406_
	);
	LUT2 #(
		.INIT('h4)
	) name26895 (
		_w36101_,
		_w36914_,
		_w37407_
	);
	LUT2 #(
		.INIT('h4)
	) name26896 (
		_w36101_,
		_w36917_,
		_w37408_
	);
	LUT2 #(
		.INIT('h4)
	) name26897 (
		_w36101_,
		_w36920_,
		_w37409_
	);
	LUT2 #(
		.INIT('h4)
	) name26898 (
		_w36101_,
		_w36923_,
		_w37410_
	);
	LUT2 #(
		.INIT('h4)
	) name26899 (
		_w36101_,
		_w36925_,
		_w37411_
	);
	LUT2 #(
		.INIT('h4)
	) name26900 (
		_w36101_,
		_w36927_,
		_w37412_
	);
	LUT2 #(
		.INIT('h4)
	) name26901 (
		_w36101_,
		_w36711_,
		_w37413_
	);
	LUT2 #(
		.INIT('h4)
	) name26902 (
		_w36101_,
		_w36930_,
		_w37414_
	);
	LUT2 #(
		.INIT('h4)
	) name26903 (
		_w36101_,
		_w36933_,
		_w37415_
	);
	LUT2 #(
		.INIT('h4)
	) name26904 (
		_w36101_,
		_w36935_,
		_w37416_
	);
	LUT2 #(
		.INIT('h4)
	) name26905 (
		_w36101_,
		_w36938_,
		_w37417_
	);
	LUT2 #(
		.INIT('h4)
	) name26906 (
		_w36101_,
		_w36940_,
		_w37418_
	);
	LUT2 #(
		.INIT('h4)
	) name26907 (
		_w36101_,
		_w36943_,
		_w37419_
	);
	LUT2 #(
		.INIT('h4)
	) name26908 (
		_w36101_,
		_w36945_,
		_w37420_
	);
	LUT2 #(
		.INIT('h4)
	) name26909 (
		_w36101_,
		_w36948_,
		_w37421_
	);
	LUT2 #(
		.INIT('h4)
	) name26910 (
		_w36101_,
		_w36950_,
		_w37422_
	);
	LUT2 #(
		.INIT('h4)
	) name26911 (
		_w36101_,
		_w36953_,
		_w37423_
	);
	LUT2 #(
		.INIT('h4)
	) name26912 (
		_w36101_,
		_w36956_,
		_w37424_
	);
	LUT2 #(
		.INIT('h4)
	) name26913 (
		_w36101_,
		_w36816_,
		_w37425_
	);
	LUT2 #(
		.INIT('h4)
	) name26914 (
		_w36101_,
		_w36959_,
		_w37426_
	);
	LUT2 #(
		.INIT('h4)
	) name26915 (
		_w36101_,
		_w36771_,
		_w37427_
	);
	LUT2 #(
		.INIT('h4)
	) name26916 (
		_w36101_,
		_w36964_,
		_w37428_
	);
	LUT2 #(
		.INIT('h4)
	) name26917 (
		_w36101_,
		_w36969_,
		_w37429_
	);
	LUT2 #(
		.INIT('h4)
	) name26918 (
		_w36101_,
		_w36972_,
		_w37430_
	);
	LUT2 #(
		.INIT('h4)
	) name26919 (
		_w36101_,
		_w36975_,
		_w37431_
	);
	LUT2 #(
		.INIT('h4)
	) name26920 (
		_w36101_,
		_w36966_,
		_w37432_
	);
	LUT2 #(
		.INIT('h4)
	) name26921 (
		_w36101_,
		_w36980_,
		_w37433_
	);
	LUT2 #(
		.INIT('h4)
	) name26922 (
		_w36101_,
		_w36982_,
		_w37434_
	);
	LUT2 #(
		.INIT('h4)
	) name26923 (
		_w36101_,
		_w36984_,
		_w37435_
	);
	LUT2 #(
		.INIT('h4)
	) name26924 (
		\ethreg1_MODER_1_DataOut_reg[4]/NET0131 ,
		_w12484_,
		_w37436_
	);
	LUT2 #(
		.INIT('h8)
	) name26925 (
		\rxethmac1_rxstatem1_StateData0_reg/NET0131 ,
		_w10576_,
		_w37437_
	);
	LUT2 #(
		.INIT('h8)
	) name26926 (
		_w34863_,
		_w37437_,
		_w37438_
	);
	LUT2 #(
		.INIT('h1)
	) name26927 (
		_w37436_,
		_w37438_,
		_w37439_
	);
	LUT2 #(
		.INIT('h8)
	) name26928 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w13499_,
		_w37440_
	);
	LUT2 #(
		.INIT('h8)
	) name26929 (
		_w22959_,
		_w31684_,
		_w37441_
	);
	LUT2 #(
		.INIT('h4)
	) name26930 (
		_w35803_,
		_w35923_,
		_w37442_
	);
	LUT2 #(
		.INIT('h8)
	) name26931 (
		_w23519_,
		_w31684_,
		_w37443_
	);
	LUT2 #(
		.INIT('h8)
	) name26932 (
		_w23519_,
		_w35976_,
		_w37444_
	);
	LUT2 #(
		.INIT('h8)
	) name26933 (
		_w22959_,
		_w35976_,
		_w37445_
	);
	LUT2 #(
		.INIT('h8)
	) name26934 (
		_w23519_,
		_w35705_,
		_w37446_
	);
	LUT2 #(
		.INIT('h8)
	) name26935 (
		_w22966_,
		_w31684_,
		_w37447_
	);
	LUT2 #(
		.INIT('h8)
	) name26936 (
		_w23499_,
		_w31684_,
		_w37448_
	);
	LUT2 #(
		.INIT('h8)
	) name26937 (
		_w22966_,
		_w35976_,
		_w37449_
	);
	LUT2 #(
		.INIT('h8)
	) name26938 (
		_w23499_,
		_w35976_,
		_w37450_
	);
	LUT2 #(
		.INIT('h8)
	) name26939 (
		_w22959_,
		_w35705_,
		_w37451_
	);
	LUT2 #(
		.INIT('h8)
	) name26940 (
		_w22966_,
		_w35705_,
		_w37452_
	);
	LUT2 #(
		.INIT('h8)
	) name26941 (
		_w31683_,
		_w36019_,
		_w37453_
	);
	LUT2 #(
		.INIT('h8)
	) name26942 (
		_w22966_,
		_w37453_,
		_w37454_
	);
	LUT2 #(
		.INIT('h8)
	) name26943 (
		_w22959_,
		_w37453_,
		_w37455_
	);
	LUT2 #(
		.INIT('h8)
	) name26944 (
		_w22952_,
		_w35976_,
		_w37456_
	);
	LUT2 #(
		.INIT('h8)
	) name26945 (
		_w22952_,
		_w35705_,
		_w37457_
	);
	LUT2 #(
		.INIT('h8)
	) name26946 (
		_w22952_,
		_w37453_,
		_w37458_
	);
	LUT2 #(
		.INIT('h8)
	) name26947 (
		_w22952_,
		_w31684_,
		_w37459_
	);
	LUT2 #(
		.INIT('h8)
	) name26948 (
		_w22956_,
		_w31684_,
		_w37460_
	);
	LUT2 #(
		.INIT('h8)
	) name26949 (
		_w22956_,
		_w35976_,
		_w37461_
	);
	LUT2 #(
		.INIT('h8)
	) name26950 (
		_w22956_,
		_w35705_,
		_w37462_
	);
	LUT2 #(
		.INIT('h8)
	) name26951 (
		_w22956_,
		_w37453_,
		_w37463_
	);
	LUT2 #(
		.INIT('h4)
	) name26952 (
		\txethmac1_txcrc_Crc_reg[31]/NET0131 ,
		_w34162_,
		_w37464_
	);
	LUT2 #(
		.INIT('h1)
	) name26953 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w37465_
	);
	LUT2 #(
		.INIT('h2)
	) name26954 (
		_w34164_,
		_w37465_,
		_w37466_
	);
	LUT2 #(
		.INIT('h1)
	) name26955 (
		_w37464_,
		_w37466_,
		_w37467_
	);
	LUT2 #(
		.INIT('h1)
	) name26956 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w37467_,
		_w37468_
	);
	LUT2 #(
		.INIT('h2)
	) name26957 (
		_w11307_,
		_w37468_,
		_w37469_
	);
	LUT2 #(
		.INIT('h8)
	) name26958 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		\txethmac1_random1_x_reg[7]/NET0131 ,
		_w37470_
	);
	LUT2 #(
		.INIT('h2)
	) name26959 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxBDReady_reg/NET0131 ,
		_w37471_
	);
	LUT2 #(
		.INIT('h2)
	) name26960 (
		\wishbone_RxAbortSync3_reg/NET0131 ,
		\wishbone_RxAbortSync4_reg/NET0131 ,
		_w37472_
	);
	LUT2 #(
		.INIT('h2)
	) name26961 (
		_w34202_,
		_w37472_,
		_w37473_
	);
	LUT2 #(
		.INIT('h1)
	) name26962 (
		\wishbone_RxReady_reg/NET0131 ,
		_w37473_,
		_w37474_
	);
	LUT2 #(
		.INIT('h1)
	) name26963 (
		_w37471_,
		_w37474_,
		_w37475_
	);
	LUT2 #(
		.INIT('h2)
	) name26964 (
		\txethmac1_random1_RandomLatched_reg[2]/NET0131 ,
		_w34968_,
		_w37476_
	);
	LUT2 #(
		.INIT('h1)
	) name26965 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w37477_
	);
	LUT2 #(
		.INIT('h4)
	) name26966 (
		_w11273_,
		_w37477_,
		_w37478_
	);
	LUT2 #(
		.INIT('h8)
	) name26967 (
		\txethmac1_random1_x_reg[2]/NET0131 ,
		_w34968_,
		_w37479_
	);
	LUT2 #(
		.INIT('h4)
	) name26968 (
		_w37478_,
		_w37479_,
		_w37480_
	);
	LUT2 #(
		.INIT('h1)
	) name26969 (
		_w37476_,
		_w37480_,
		_w37481_
	);
	LUT2 #(
		.INIT('h1)
	) name26970 (
		\wishbone_RxBDAddress_reg[1]/NET0131 ,
		_w34201_,
		_w37482_
	);
	LUT2 #(
		.INIT('h1)
	) name26971 (
		_w34593_,
		_w37482_,
		_w37483_
	);
	LUT2 #(
		.INIT('h4)
	) name26972 (
		_w34204_,
		_w37483_,
		_w37484_
	);
	LUT2 #(
		.INIT('h8)
	) name26973 (
		\ethreg1_TX_BD_NUM_0_DataOut_reg[0]/NET0131 ,
		_w34204_,
		_w37485_
	);
	LUT2 #(
		.INIT('h1)
	) name26974 (
		_w37484_,
		_w37485_,
		_w37486_
	);
	LUT2 #(
		.INIT('h2)
	) name26975 (
		\wishbone_TxEn_needed_reg/NET0131 ,
		_w17883_,
		_w37487_
	);
	LUT2 #(
		.INIT('h4)
	) name26976 (
		\wishbone_WbEn_q_reg/NET0131 ,
		\wishbone_WbEn_reg/NET0131 ,
		_w37488_
	);
	LUT2 #(
		.INIT('h4)
	) name26977 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w37488_,
		_w37489_
	);
	LUT2 #(
		.INIT('h8)
	) name26978 (
		_w34888_,
		_w37489_,
		_w37490_
	);
	LUT2 #(
		.INIT('h1)
	) name26979 (
		_w37487_,
		_w37490_,
		_w37491_
	);
	LUT2 #(
		.INIT('h8)
	) name26980 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[2]/NET0131 ,
		_w35627_,
		_w37492_
	);
	LUT2 #(
		.INIT('h8)
	) name26981 (
		\ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 ,
		_w35830_,
		_w37493_
	);
	LUT2 #(
		.INIT('h8)
	) name26982 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[2]/NET0131 ,
		_w35625_,
		_w37494_
	);
	LUT2 #(
		.INIT('h8)
	) name26983 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[2]/NET0131 ,
		_w35827_,
		_w37495_
	);
	LUT2 #(
		.INIT('h8)
	) name26984 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		_w34938_,
		_w37496_
	);
	LUT2 #(
		.INIT('h8)
	) name26985 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[2]/NET0131 ,
		_w35622_,
		_w37497_
	);
	LUT2 #(
		.INIT('h8)
	) name26986 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		_w34955_,
		_w37498_
	);
	LUT2 #(
		.INIT('h8)
	) name26987 (
		\ethreg1_TXCTRL_0_DataOut_reg[2]/NET0131 ,
		_w34266_,
		_w37499_
	);
	LUT2 #(
		.INIT('h1)
	) name26988 (
		_w37492_,
		_w37493_,
		_w37500_
	);
	LUT2 #(
		.INIT('h1)
	) name26989 (
		_w37494_,
		_w37495_,
		_w37501_
	);
	LUT2 #(
		.INIT('h1)
	) name26990 (
		_w37496_,
		_w37497_,
		_w37502_
	);
	LUT2 #(
		.INIT('h1)
	) name26991 (
		_w37498_,
		_w37499_,
		_w37503_
	);
	LUT2 #(
		.INIT('h8)
	) name26992 (
		_w37502_,
		_w37503_,
		_w37504_
	);
	LUT2 #(
		.INIT('h8)
	) name26993 (
		_w37500_,
		_w37501_,
		_w37505_
	);
	LUT2 #(
		.INIT('h8)
	) name26994 (
		_w37504_,
		_w37505_,
		_w37506_
	);
	LUT2 #(
		.INIT('h8)
	) name26995 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[4]/NET0131 ,
		_w35627_,
		_w37507_
	);
	LUT2 #(
		.INIT('h8)
	) name26996 (
		\ethreg1_TXCTRL_1_DataOut_reg[4]/NET0131 ,
		_w35830_,
		_w37508_
	);
	LUT2 #(
		.INIT('h8)
	) name26997 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[4]/NET0131 ,
		_w35625_,
		_w37509_
	);
	LUT2 #(
		.INIT('h8)
	) name26998 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[4]/NET0131 ,
		_w35827_,
		_w37510_
	);
	LUT2 #(
		.INIT('h8)
	) name26999 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[4]/NET0131 ,
		_w34938_,
		_w37511_
	);
	LUT2 #(
		.INIT('h8)
	) name27000 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[4]/NET0131 ,
		_w35622_,
		_w37512_
	);
	LUT2 #(
		.INIT('h8)
	) name27001 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[4]/NET0131 ,
		_w34955_,
		_w37513_
	);
	LUT2 #(
		.INIT('h8)
	) name27002 (
		\ethreg1_TXCTRL_0_DataOut_reg[4]/NET0131 ,
		_w34266_,
		_w37514_
	);
	LUT2 #(
		.INIT('h1)
	) name27003 (
		_w37507_,
		_w37508_,
		_w37515_
	);
	LUT2 #(
		.INIT('h1)
	) name27004 (
		_w37509_,
		_w37510_,
		_w37516_
	);
	LUT2 #(
		.INIT('h1)
	) name27005 (
		_w37511_,
		_w37512_,
		_w37517_
	);
	LUT2 #(
		.INIT('h1)
	) name27006 (
		_w37513_,
		_w37514_,
		_w37518_
	);
	LUT2 #(
		.INIT('h8)
	) name27007 (
		_w37517_,
		_w37518_,
		_w37519_
	);
	LUT2 #(
		.INIT('h8)
	) name27008 (
		_w37515_,
		_w37516_,
		_w37520_
	);
	LUT2 #(
		.INIT('h8)
	) name27009 (
		_w37519_,
		_w37520_,
		_w37521_
	);
	LUT2 #(
		.INIT('h8)
	) name27010 (
		\ethreg1_MAC_ADDR0_0_DataOut_reg[5]/NET0131 ,
		_w35627_,
		_w37522_
	);
	LUT2 #(
		.INIT('h8)
	) name27011 (
		\ethreg1_TXCTRL_1_DataOut_reg[5]/NET0131 ,
		_w35830_,
		_w37523_
	);
	LUT2 #(
		.INIT('h8)
	) name27012 (
		\ethreg1_MAC_ADDR0_2_DataOut_reg[5]/NET0131 ,
		_w35625_,
		_w37524_
	);
	LUT2 #(
		.INIT('h8)
	) name27013 (
		\ethreg1_MAC_ADDR0_3_DataOut_reg[5]/NET0131 ,
		_w35827_,
		_w37525_
	);
	LUT2 #(
		.INIT('h8)
	) name27014 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[5]/NET0131 ,
		_w34938_,
		_w37526_
	);
	LUT2 #(
		.INIT('h8)
	) name27015 (
		\ethreg1_MAC_ADDR1_0_DataOut_reg[5]/NET0131 ,
		_w35622_,
		_w37527_
	);
	LUT2 #(
		.INIT('h8)
	) name27016 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[5]/NET0131 ,
		_w34955_,
		_w37528_
	);
	LUT2 #(
		.INIT('h8)
	) name27017 (
		\ethreg1_TXCTRL_0_DataOut_reg[5]/NET0131 ,
		_w34266_,
		_w37529_
	);
	LUT2 #(
		.INIT('h1)
	) name27018 (
		_w37522_,
		_w37523_,
		_w37530_
	);
	LUT2 #(
		.INIT('h1)
	) name27019 (
		_w37524_,
		_w37525_,
		_w37531_
	);
	LUT2 #(
		.INIT('h1)
	) name27020 (
		_w37526_,
		_w37527_,
		_w37532_
	);
	LUT2 #(
		.INIT('h1)
	) name27021 (
		_w37528_,
		_w37529_,
		_w37533_
	);
	LUT2 #(
		.INIT('h8)
	) name27022 (
		_w37532_,
		_w37533_,
		_w37534_
	);
	LUT2 #(
		.INIT('h8)
	) name27023 (
		_w37530_,
		_w37531_,
		_w37535_
	);
	LUT2 #(
		.INIT('h8)
	) name27024 (
		_w37534_,
		_w37535_,
		_w37536_
	);
	LUT2 #(
		.INIT('h1)
	) name27025 (
		\wishbone_TxAbort_wb_reg/NET0131 ,
		\wishbone_TxDone_wb_reg/NET0131 ,
		_w37537_
	);
	LUT2 #(
		.INIT('h1)
	) name27026 (
		\wishbone_BlockingTxStatusWrite_reg/NET0131 ,
		_w34891_,
		_w37538_
	);
	LUT2 #(
		.INIT('h1)
	) name27027 (
		_w37537_,
		_w37538_,
		_w37539_
	);
	LUT2 #(
		.INIT('h2)
	) name27028 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w37540_
	);
	LUT2 #(
		.INIT('h2)
	) name27029 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w37541_
	);
	LUT2 #(
		.INIT('h2)
	) name27030 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w37542_
	);
	LUT2 #(
		.INIT('h2)
	) name27031 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w37543_
	);
	LUT2 #(
		.INIT('h4)
	) name27032 (
		\ethreg1_COLLCONF_0_DataOut_reg[5]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[5]/NET0131 ,
		_w37544_
	);
	LUT2 #(
		.INIT('h4)
	) name27033 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w37545_
	);
	LUT2 #(
		.INIT('h4)
	) name27034 (
		\ethreg1_COLLCONF_0_DataOut_reg[3]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[3]/NET0131 ,
		_w37546_
	);
	LUT2 #(
		.INIT('h4)
	) name27035 (
		\ethreg1_COLLCONF_0_DataOut_reg[0]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[0]/NET0131 ,
		_w37547_
	);
	LUT2 #(
		.INIT('h2)
	) name27036 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w37548_
	);
	LUT2 #(
		.INIT('h4)
	) name27037 (
		\ethreg1_COLLCONF_0_DataOut_reg[2]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[2]/NET0131 ,
		_w37549_
	);
	LUT2 #(
		.INIT('h2)
	) name27038 (
		\ethreg1_COLLCONF_0_DataOut_reg[4]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[4]/NET0131 ,
		_w37550_
	);
	LUT2 #(
		.INIT('h4)
	) name27039 (
		\ethreg1_COLLCONF_0_DataOut_reg[1]/NET0131 ,
		\txethmac1_txcounters1_ByteCnt_reg[1]/NET0131 ,
		_w37551_
	);
	LUT2 #(
		.INIT('h1)
	) name27040 (
		_w10684_,
		_w37540_,
		_w37552_
	);
	LUT2 #(
		.INIT('h1)
	) name27041 (
		_w37541_,
		_w37542_,
		_w37553_
	);
	LUT2 #(
		.INIT('h1)
	) name27042 (
		_w37543_,
		_w37544_,
		_w37554_
	);
	LUT2 #(
		.INIT('h1)
	) name27043 (
		_w37545_,
		_w37546_,
		_w37555_
	);
	LUT2 #(
		.INIT('h1)
	) name27044 (
		_w37547_,
		_w37548_,
		_w37556_
	);
	LUT2 #(
		.INIT('h1)
	) name27045 (
		_w37549_,
		_w37550_,
		_w37557_
	);
	LUT2 #(
		.INIT('h4)
	) name27046 (
		_w37551_,
		_w37557_,
		_w37558_
	);
	LUT2 #(
		.INIT('h8)
	) name27047 (
		_w37555_,
		_w37556_,
		_w37559_
	);
	LUT2 #(
		.INIT('h8)
	) name27048 (
		_w37553_,
		_w37554_,
		_w37560_
	);
	LUT2 #(
		.INIT('h8)
	) name27049 (
		_w37552_,
		_w37560_,
		_w37561_
	);
	LUT2 #(
		.INIT('h8)
	) name27050 (
		_w37558_,
		_w37559_,
		_w37562_
	);
	LUT2 #(
		.INIT('h4)
	) name27051 (
		_w14559_,
		_w37562_,
		_w37563_
	);
	LUT2 #(
		.INIT('h8)
	) name27052 (
		_w37561_,
		_w37563_,
		_w37564_
	);
	LUT2 #(
		.INIT('h1)
	) name27053 (
		\txethmac1_ColWindow_reg/NET0131 ,
		\txethmac1_txstatem1_StateIPG_reg/NET0131 ,
		_w37565_
	);
	LUT2 #(
		.INIT('h4)
	) name27054 (
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w37565_,
		_w37566_
	);
	LUT2 #(
		.INIT('h1)
	) name27055 (
		_w37564_,
		_w37566_,
		_w37567_
	);
	LUT2 #(
		.INIT('h4)
	) name27056 (
		\txethmac1_txcrc_Crc_reg[30]/NET0131 ,
		_w34162_,
		_w37568_
	);
	LUT2 #(
		.INIT('h1)
	) name27057 (
		_w11339_,
		_w37568_,
		_w37569_
	);
	LUT2 #(
		.INIT('h1)
	) name27058 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w37569_,
		_w37570_
	);
	LUT2 #(
		.INIT('h1)
	) name27059 (
		_w11344_,
		_w37570_,
		_w37571_
	);
	LUT2 #(
		.INIT('h1)
	) name27060 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[1]/NET0131 ,
		_w11620_,
		_w37572_
	);
	LUT2 #(
		.INIT('h1)
	) name27061 (
		wb_rst_i_pad,
		_w11621_,
		_w37573_
	);
	LUT2 #(
		.INIT('h4)
	) name27062 (
		_w37572_,
		_w37573_,
		_w37574_
	);
	LUT2 #(
		.INIT('h1)
	) name27063 (
		\wishbone_RxStatusInLatched_reg[0]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[1]/NET0131 ,
		_w37575_
	);
	LUT2 #(
		.INIT('h1)
	) name27064 (
		\wishbone_RxStatusInLatched_reg[3]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[4]/NET0131 ,
		_w37576_
	);
	LUT2 #(
		.INIT('h1)
	) name27065 (
		\wishbone_RxStatusInLatched_reg[5]/NET0131 ,
		\wishbone_RxStatusInLatched_reg[6]/NET0131 ,
		_w37577_
	);
	LUT2 #(
		.INIT('h8)
	) name27066 (
		_w37576_,
		_w37577_,
		_w37578_
	);
	LUT2 #(
		.INIT('h8)
	) name27067 (
		_w37575_,
		_w37578_,
		_w37579_
	);
	LUT2 #(
		.INIT('h2)
	) name27068 (
		\ethreg1_CTRLMODER_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_CTRLMODER_0_DataOut_reg[1]/NET0131 ,
		_w37580_
	);
	LUT2 #(
		.INIT('h2)
	) name27069 (
		\maccontrol1_receivecontrol1_ReceivedPauseFrm_reg/NET0131 ,
		_w37580_,
		_w37581_
	);
	LUT2 #(
		.INIT('h8)
	) name27070 (
		\wishbone_RxStatus_reg[14]/NET0131 ,
		_w34201_,
		_w37582_
	);
	LUT2 #(
		.INIT('h4)
	) name27071 (
		_w37581_,
		_w37582_,
		_w37583_
	);
	LUT2 #(
		.INIT('h4)
	) name27072 (
		\macstatus1_LatchedCrcError_reg/NET0131 ,
		_w37579_,
		_w37584_
	);
	LUT2 #(
		.INIT('h8)
	) name27073 (
		_w37583_,
		_w37584_,
		_w37585_
	);
	LUT2 #(
		.INIT('h4)
	) name27074 (
		_w37579_,
		_w37583_,
		_w37586_
	);
	LUT2 #(
		.INIT('h2)
	) name27075 (
		\miim1_RStat_q2_reg/NET0131 ,
		\miim1_RStat_q3_reg/NET0131 ,
		_w37587_
	);
	LUT2 #(
		.INIT('h1)
	) name27076 (
		\miim1_RStatStart_reg/NET0131 ,
		_w37587_,
		_w37588_
	);
	LUT2 #(
		.INIT('h1)
	) name27077 (
		\miim1_EndBusy_reg/NET0131 ,
		_w37588_,
		_w37589_
	);
	LUT2 #(
		.INIT('h8)
	) name27078 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		_w36005_,
		_w37590_
	);
	LUT2 #(
		.INIT('h1)
	) name27079 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[1]/NET0131 ,
		_w37590_,
		_w37591_
	);
	LUT2 #(
		.INIT('h2)
	) name27080 (
		_w34259_,
		_w36006_,
		_w37592_
	);
	LUT2 #(
		.INIT('h4)
	) name27081 (
		_w37591_,
		_w37592_,
		_w37593_
	);
	LUT2 #(
		.INIT('h1)
	) name27082 (
		\maccontrol1_transmitcontrol1_ControlEnd_q_reg/P0001 ,
		_w34266_,
		_w37594_
	);
	LUT2 #(
		.INIT('h2)
	) name27083 (
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w15175_,
		_w37595_
	);
	LUT2 #(
		.INIT('h2)
	) name27084 (
		\wishbone_ShiftEndedSync3_reg/NET0131 ,
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w37596_
	);
	LUT2 #(
		.INIT('h2)
	) name27085 (
		\wishbone_rx_fifo_cnt_reg[0]/NET0131 ,
		\wishbone_rx_fifo_cnt_reg[1]/NET0131 ,
		_w37597_
	);
	LUT2 #(
		.INIT('h4)
	) name27086 (
		\wishbone_rx_fifo_cnt_reg[2]/NET0131 ,
		_w37597_,
		_w37598_
	);
	LUT2 #(
		.INIT('h8)
	) name27087 (
		_w12553_,
		_w15698_,
		_w37599_
	);
	LUT2 #(
		.INIT('h8)
	) name27088 (
		_w37596_,
		_w37599_,
		_w37600_
	);
	LUT2 #(
		.INIT('h8)
	) name27089 (
		_w37598_,
		_w37600_,
		_w37601_
	);
	LUT2 #(
		.INIT('h1)
	) name27090 (
		_w37595_,
		_w37601_,
		_w37602_
	);
	LUT2 #(
		.INIT('h2)
	) name27091 (
		\txethmac1_random1_RandomLatched_reg[4]/NET0131 ,
		_w34968_,
		_w37603_
	);
	LUT2 #(
		.INIT('h2)
	) name27092 (
		\txethmac1_RetryCnt_reg[2]/NET0131 ,
		_w35740_,
		_w37604_
	);
	LUT2 #(
		.INIT('h1)
	) name27093 (
		\txethmac1_RetryCnt_reg[3]/NET0131 ,
		_w37604_,
		_w37605_
	);
	LUT2 #(
		.INIT('h8)
	) name27094 (
		\txethmac1_random1_x_reg[4]/NET0131 ,
		_w34968_,
		_w37606_
	);
	LUT2 #(
		.INIT('h4)
	) name27095 (
		_w37605_,
		_w37606_,
		_w37607_
	);
	LUT2 #(
		.INIT('h1)
	) name27096 (
		_w37603_,
		_w37607_,
		_w37608_
	);
	LUT2 #(
		.INIT('h1)
	) name27097 (
		\wishbone_RxReady_reg/NET0131 ,
		_w15696_,
		_w37609_
	);
	LUT2 #(
		.INIT('h2)
	) name27098 (
		\wishbone_RxAbortSync2_reg/NET0131 ,
		\wishbone_RxAbortSync3_reg/NET0131 ,
		_w37610_
	);
	LUT2 #(
		.INIT('h2)
	) name27099 (
		\wishbone_r_RxEn_q_reg/NET0131 ,
		_w34199_,
		_w37611_
	);
	LUT2 #(
		.INIT('h1)
	) name27100 (
		\wishbone_ShiftEnded_reg/NET0131 ,
		_w37610_,
		_w37612_
	);
	LUT2 #(
		.INIT('h4)
	) name27101 (
		_w37611_,
		_w37612_,
		_w37613_
	);
	LUT2 #(
		.INIT('h4)
	) name27102 (
		_w37609_,
		_w37613_,
		_w37614_
	);
	LUT2 #(
		.INIT('h8)
	) name27103 (
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		_w11099_,
		_w37615_
	);
	LUT2 #(
		.INIT('h1)
	) name27104 (
		\CarrierSense_Tx2_reg/NET0131 ,
		\ethreg1_MODER_0_DataOut_reg[7]/NET0131 ,
		_w37616_
	);
	LUT2 #(
		.INIT('h1)
	) name27105 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		mcoll_pad_i_pad,
		_w37617_
	);
	LUT2 #(
		.INIT('h8)
	) name27106 (
		_w37616_,
		_w37617_,
		_w37618_
	);
	LUT2 #(
		.INIT('h4)
	) name27107 (
		_w11108_,
		_w37618_,
		_w37619_
	);
	LUT2 #(
		.INIT('h1)
	) name27108 (
		_w37615_,
		_w37619_,
		_w37620_
	);
	LUT2 #(
		.INIT('h1)
	) name27109 (
		\wishbone_Flop_reg/NET0131 ,
		_w12240_,
		_w37621_
	);
	LUT2 #(
		.INIT('h1)
	) name27110 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w37622_
	);
	LUT2 #(
		.INIT('h4)
	) name27111 (
		\maccontrol1_MuxedDone_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		_w37623_
	);
	LUT2 #(
		.INIT('h2)
	) name27112 (
		_w35894_,
		_w37622_,
		_w37624_
	);
	LUT2 #(
		.INIT('h4)
	) name27113 (
		_w37623_,
		_w37624_,
		_w37625_
	);
	LUT2 #(
		.INIT('h1)
	) name27114 (
		_w12246_,
		_w37621_,
		_w37626_
	);
	LUT2 #(
		.INIT('h4)
	) name27115 (
		_w37625_,
		_w37626_,
		_w37627_
	);
	LUT2 #(
		.INIT('h8)
	) name27116 (
		_w36084_,
		_w37627_,
		_w37628_
	);
	LUT2 #(
		.INIT('h4)
	) name27117 (
		\txethmac1_txcrc_Crc_reg[29]/NET0131 ,
		_w34162_,
		_w37629_
	);
	LUT2 #(
		.INIT('h4)
	) name27118 (
		\txethmac1_txstatem1_StateJam_reg/NET0131 ,
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w37630_
	);
	LUT2 #(
		.INIT('h8)
	) name27119 (
		_w34164_,
		_w37630_,
		_w37631_
	);
	LUT2 #(
		.INIT('h1)
	) name27120 (
		_w37629_,
		_w37631_,
		_w37632_
	);
	LUT2 #(
		.INIT('h1)
	) name27121 (
		\txethmac1_txstatem1_StateData_reg[0]/NET0131 ,
		_w37632_,
		_w37633_
	);
	LUT2 #(
		.INIT('h2)
	) name27122 (
		_w11327_,
		_w37633_,
		_w37634_
	);
	LUT2 #(
		.INIT('h8)
	) name27123 (
		\wishbone_TxStatus_reg[14]/NET0131 ,
		_w34892_,
		_w37635_
	);
	LUT2 #(
		.INIT('h1)
	) name27124 (
		\macstatus1_CarrierSenseLost_reg/NET0131 ,
		\macstatus1_LateCollLatched_reg/P0002 ,
		_w37636_
	);
	LUT2 #(
		.INIT('h1)
	) name27125 (
		\macstatus1_RetryLimit_reg/P0002 ,
		\wishbone_TxUnderRun_reg/NET0131 ,
		_w37637_
	);
	LUT2 #(
		.INIT('h8)
	) name27126 (
		_w37636_,
		_w37637_,
		_w37638_
	);
	LUT2 #(
		.INIT('h8)
	) name27127 (
		_w37635_,
		_w37638_,
		_w37639_
	);
	LUT2 #(
		.INIT('h2)
	) name27128 (
		_w37635_,
		_w37638_,
		_w37640_
	);
	LUT2 #(
		.INIT('h1)
	) name27129 (
		\maccontrol1_transmitcontrol1_DlyCrcCnt_reg[0]/NET0131 ,
		_w36005_,
		_w37641_
	);
	LUT2 #(
		.INIT('h2)
	) name27130 (
		_w34259_,
		_w37590_,
		_w37642_
	);
	LUT2 #(
		.INIT('h4)
	) name27131 (
		_w37641_,
		_w37642_,
		_w37643_
	);
	LUT2 #(
		.INIT('h1)
	) name27132 (
		\maccontrol1_receivecontrol1_SlotTimer_reg[0]/NET0131 ,
		_w11619_,
		_w37644_
	);
	LUT2 #(
		.INIT('h1)
	) name27133 (
		wb_rst_i_pad,
		_w11620_,
		_w37645_
	);
	LUT2 #(
		.INIT('h4)
	) name27134 (
		_w37644_,
		_w37645_,
		_w37646_
	);
	LUT2 #(
		.INIT('h2)
	) name27135 (
		\miim1_ScanStat_q2_reg/NET0131 ,
		\miim1_SyncStatMdcEn_reg/NET0131 ,
		_w37647_
	);
	LUT2 #(
		.INIT('h1)
	) name27136 (
		\miim1_Nvalid_reg/NET0131 ,
		_w37647_,
		_w37648_
	);
	LUT2 #(
		.INIT('h4)
	) name27137 (
		\miim1_InProgress_q2_reg/NET0131 ,
		\miim1_InProgress_q3_reg/NET0131 ,
		_w37649_
	);
	LUT2 #(
		.INIT('h1)
	) name27138 (
		_w37648_,
		_w37649_,
		_w37650_
	);
	LUT2 #(
		.INIT('h2)
	) name27139 (
		\TxPauseRq_sync2_reg/NET0131 ,
		\TxPauseRq_sync3_reg/NET0131 ,
		_w37651_
	);
	LUT2 #(
		.INIT('h8)
	) name27140 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_TxUsedDataIn_q_reg/NET0131 ,
		_w37652_
	);
	LUT2 #(
		.INIT('h2)
	) name27141 (
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		_w12240_,
		_w37653_
	);
	LUT2 #(
		.INIT('h8)
	) name27142 (
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		_w34257_,
		_w37654_
	);
	LUT2 #(
		.INIT('h4)
	) name27143 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w37654_,
		_w37655_
	);
	LUT2 #(
		.INIT('h2)
	) name27144 (
		_w37653_,
		_w37655_,
		_w37656_
	);
	LUT2 #(
		.INIT('h1)
	) name27145 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w37656_,
		_w37657_
	);
	LUT2 #(
		.INIT('h1)
	) name27146 (
		_w37652_,
		_w37657_,
		_w37658_
	);
	LUT2 #(
		.INIT('h2)
	) name27147 (
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		\wishbone_BlockingTxStatusWrite_sync3_reg/NET0131 ,
		_w37659_
	);
	LUT2 #(
		.INIT('h2)
	) name27148 (
		\macstatus1_DeferLatched_reg/NET0131 ,
		_w37659_,
		_w37660_
	);
	LUT2 #(
		.INIT('h1)
	) name27149 (
		_w11060_,
		_w37660_,
		_w37661_
	);
	LUT2 #(
		.INIT('h2)
	) name27150 (
		\txethmac1_random1_RandomLatched_reg[3]/NET0131 ,
		_w34968_,
		_w37662_
	);
	LUT2 #(
		.INIT('h8)
	) name27151 (
		\txethmac1_random1_x_reg[3]/NET0131 ,
		_w34968_,
		_w37663_
	);
	LUT2 #(
		.INIT('h4)
	) name27152 (
		_w37477_,
		_w37663_,
		_w37664_
	);
	LUT2 #(
		.INIT('h1)
	) name27153 (
		_w37662_,
		_w37664_,
		_w37665_
	);
	LUT2 #(
		.INIT('h1)
	) name27154 (
		\wishbone_RxStatusWriteLatched_reg/NET0131 ,
		_w34201_,
		_w37666_
	);
	LUT2 #(
		.INIT('h1)
	) name27155 (
		\wishbone_RxStatusWriteLatched_syncb2_reg/NET0131 ,
		_w37666_,
		_w37667_
	);
	LUT2 #(
		.INIT('h2)
	) name27156 (
		\miim1_WCtrlData_q2_reg/NET0131 ,
		\miim1_WCtrlData_q3_reg/NET0131 ,
		_w37668_
	);
	LUT2 #(
		.INIT('h1)
	) name27157 (
		\miim1_WCtrlDataStart_reg/NET0131 ,
		_w37668_,
		_w37669_
	);
	LUT2 #(
		.INIT('h1)
	) name27158 (
		\miim1_EndBusy_reg/NET0131 ,
		_w37669_,
		_w37670_
	);
	LUT2 #(
		.INIT('h2)
	) name27159 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[0]/NET0131 ,
		\ethreg1_MIIADDRESS_1_DataOut_reg[1]/NET0131 ,
		_w37671_
	);
	LUT2 #(
		.INIT('h1)
	) name27160 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		\ethreg1_MIIADDRESS_1_DataOut_reg[3]/NET0131 ,
		_w37672_
	);
	LUT2 #(
		.INIT('h4)
	) name27161 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[4]/NET0131 ,
		_w37672_,
		_w37673_
	);
	LUT2 #(
		.INIT('h8)
	) name27162 (
		_w37671_,
		_w37673_,
		_w37674_
	);
	LUT2 #(
		.INIT('h4)
	) name27163 (
		\miim1_shftrg_ShiftReg_reg[1]/NET0131 ,
		_w37674_,
		_w37675_
	);
	LUT2 #(
		.INIT('h2)
	) name27164 (
		\miim1_shftrg_LinkFail_reg/NET0131 ,
		_w37674_,
		_w37676_
	);
	LUT2 #(
		.INIT('h1)
	) name27165 (
		_w37675_,
		_w37676_,
		_w37677_
	);
	LUT2 #(
		.INIT('h2)
	) name27166 (
		\wishbone_RxEn_needed_reg/NET0131 ,
		_w15696_,
		_w37678_
	);
	LUT2 #(
		.INIT('h4)
	) name27167 (
		\wishbone_RxReady_reg/NET0131 ,
		_w34199_,
		_w37679_
	);
	LUT2 #(
		.INIT('h8)
	) name27168 (
		_w37488_,
		_w37679_,
		_w37680_
	);
	LUT2 #(
		.INIT('h1)
	) name27169 (
		_w37678_,
		_w37680_,
		_w37681_
	);
	LUT2 #(
		.INIT('h4)
	) name27170 (
		wb_err_o_pad,
		_w22937_,
		_w37682_
	);
	LUT2 #(
		.INIT('h4)
	) name27171 (
		_w22941_,
		_w37682_,
		_w37683_
	);
	LUT2 #(
		.INIT('h4)
	) name27172 (
		\maccontrol1_TxDoneInLatched_reg/NET0131 ,
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		_w37684_
	);
	LUT2 #(
		.INIT('h8)
	) name27173 (
		\txethmac1_TxDone_reg/NET0131 ,
		_w37684_,
		_w37685_
	);
	LUT2 #(
		.INIT('h1)
	) name27174 (
		\maccontrol1_MuxedDone_reg/NET0131 ,
		_w37685_,
		_w37686_
	);
	LUT2 #(
		.INIT('h1)
	) name27175 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w37686_,
		_w37687_
	);
	LUT2 #(
		.INIT('h4)
	) name27176 (
		\maccontrol1_TxAbortInLatched_reg/NET0131 ,
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		_w37688_
	);
	LUT2 #(
		.INIT('h8)
	) name27177 (
		\txethmac1_TxAbort_reg/NET0131 ,
		_w37688_,
		_w37689_
	);
	LUT2 #(
		.INIT('h1)
	) name27178 (
		\maccontrol1_MuxedAbort_reg/NET0131 ,
		_w37689_,
		_w37690_
	);
	LUT2 #(
		.INIT('h1)
	) name27179 (
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w37690_,
		_w37691_
	);
	LUT2 #(
		.INIT('h2)
	) name27180 (
		\ethreg1_SetTxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetTxCIrq_sync3_reg/NET0131 ,
		_w37692_
	);
	LUT2 #(
		.INIT('h2)
	) name27181 (
		\ethreg1_SetRxCIrq_sync2_reg/NET0131 ,
		\ethreg1_SetRxCIrq_sync3_reg/NET0131 ,
		_w37693_
	);
	LUT2 #(
		.INIT('h8)
	) name27182 (
		\wishbone_BDRead_reg/NET0131 ,
		_w37488_,
		_w37694_
	);
	LUT2 #(
		.INIT('h1)
	) name27183 (
		\wishbone_BDWrite_reg[0]/NET0131 ,
		\wishbone_BDWrite_reg[1]/NET0131 ,
		_w37695_
	);
	LUT2 #(
		.INIT('h1)
	) name27184 (
		\wishbone_BDWrite_reg[2]/NET0131 ,
		\wishbone_BDWrite_reg[3]/NET0131 ,
		_w37696_
	);
	LUT2 #(
		.INIT('h8)
	) name27185 (
		_w37695_,
		_w37696_,
		_w37697_
	);
	LUT2 #(
		.INIT('h2)
	) name27186 (
		_w36098_,
		_w37697_,
		_w37698_
	);
	LUT2 #(
		.INIT('h1)
	) name27187 (
		_w37694_,
		_w37698_,
		_w37699_
	);
	LUT2 #(
		.INIT('h2)
	) name27188 (
		_w11099_,
		_w37654_,
		_w37700_
	);
	LUT2 #(
		.INIT('h2)
	) name27189 (
		\WillSendControlFrame_sync2_reg/NET0131 ,
		\WillSendControlFrame_sync3_reg/NET0131 ,
		_w37701_
	);
	LUT2 #(
		.INIT('h2)
	) name27190 (
		\txethmac1_random1_RandomLatched_reg[1]/NET0131 ,
		_w34968_,
		_w37702_
	);
	LUT2 #(
		.INIT('h4)
	) name27191 (
		\txethmac1_RetryCnt_reg[1]/NET0131 ,
		_w37477_,
		_w37703_
	);
	LUT2 #(
		.INIT('h8)
	) name27192 (
		\txethmac1_random1_x_reg[1]/NET0131 ,
		_w34968_,
		_w37704_
	);
	LUT2 #(
		.INIT('h4)
	) name27193 (
		_w37703_,
		_w37704_,
		_w37705_
	);
	LUT2 #(
		.INIT('h1)
	) name27194 (
		_w37702_,
		_w37705_,
		_w37706_
	);
	LUT2 #(
		.INIT('h4)
	) name27195 (
		\ethreg1_MODER_2_DataOut_reg[0]/NET0131 ,
		\macstatus1_RxColWindow_reg/NET0131 ,
		_w37707_
	);
	LUT2 #(
		.INIT('h4)
	) name27196 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		mcoll_pad_i_pad,
		_w37708_
	);
	LUT2 #(
		.INIT('h4)
	) name27197 (
		_w37707_,
		_w37708_,
		_w37709_
	);
	LUT2 #(
		.INIT('h1)
	) name27198 (
		\macstatus1_RxLateCollision_reg/NET0131 ,
		_w37709_,
		_w37710_
	);
	LUT2 #(
		.INIT('h1)
	) name27199 (
		\macstatus1_LoadRxStatus_reg/NET0131 ,
		_w37710_,
		_w37711_
	);
	LUT2 #(
		.INIT('h1)
	) name27200 (
		\Collision_Tx1_reg/NET0131 ,
		\Collision_Tx2_reg/NET0131 ,
		_w37712_
	);
	LUT2 #(
		.INIT('h1)
	) name27201 (
		_w11109_,
		_w37712_,
		_w37713_
	);
	LUT2 #(
		.INIT('h2)
	) name27202 (
		\wishbone_RxPointerRead_reg/NET0131 ,
		_w15175_,
		_w37714_
	);
	LUT2 #(
		.INIT('h8)
	) name27203 (
		\wishbone_RxBDRead_reg/NET0131 ,
		\wishbone_RxBDReady_reg/NET0131 ,
		_w37715_
	);
	LUT2 #(
		.INIT('h1)
	) name27204 (
		_w37714_,
		_w37715_,
		_w37716_
	);
	LUT2 #(
		.INIT('h1)
	) name27205 (
		\maccontrol1_TxUsedDataOutDetected_reg/NET0131 ,
		_w12240_,
		_w37717_
	);
	LUT2 #(
		.INIT('h2)
	) name27206 (
		_w34257_,
		_w37717_,
		_w37718_
	);
	LUT2 #(
		.INIT('h2)
	) name27207 (
		\wishbone_ShiftEndedSync1_reg/NET0131 ,
		\wishbone_ShiftEndedSync2_reg/NET0131 ,
		_w37719_
	);
	LUT2 #(
		.INIT('h1)
	) name27208 (
		_w37596_,
		_w37719_,
		_w37720_
	);
	LUT2 #(
		.INIT('h1)
	) name27209 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		\txethmac1_txstatem1_Rule1_reg/NET0131 ,
		_w37721_
	);
	LUT2 #(
		.INIT('h4)
	) name27210 (
		\txethmac1_txstatem1_StatePreamble_reg/NET0131 ,
		_w37721_,
		_w37722_
	);
	LUT2 #(
		.INIT('h1)
	) name27211 (
		\txethmac1_txstatem1_StateBackOff_reg/NET0131 ,
		\txethmac1_txstatem1_StateIdle_reg/NET0131 ,
		_w37723_
	);
	LUT2 #(
		.INIT('h4)
	) name27212 (
		_w37722_,
		_w37723_,
		_w37724_
	);
	LUT2 #(
		.INIT('h1)
	) name27213 (
		\wishbone_TxRetryPacketBlocked_reg/NET0131 ,
		\wishbone_TxRetryPacket_reg/NET0131 ,
		_w37725_
	);
	LUT2 #(
		.INIT('h2)
	) name27214 (
		\wishbone_TxRetry_wb_q_reg/NET0131 ,
		\wishbone_TxRetry_wb_reg/NET0131 ,
		_w37726_
	);
	LUT2 #(
		.INIT('h1)
	) name27215 (
		_w37725_,
		_w37726_,
		_w37727_
	);
	LUT2 #(
		.INIT('h1)
	) name27216 (
		\RxAbort_wb_reg/NET0131 ,
		\wishbone_RxAbortLatched_reg/NET0131 ,
		_w37728_
	);
	LUT2 #(
		.INIT('h1)
	) name27217 (
		\wishbone_RxAbortSyncb2_reg/NET0131 ,
		_w37728_,
		_w37729_
	);
	LUT2 #(
		.INIT('h2)
	) name27218 (
		\maccontrol1_transmitcontrol1_CtrlMux_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w37730_
	);
	LUT2 #(
		.INIT('h1)
	) name27219 (
		_w37653_,
		_w37730_,
		_w37731_
	);
	LUT2 #(
		.INIT('h4)
	) name27220 (
		\wishbone_TxEn_q_reg/NET0131 ,
		\wishbone_TxPointerRead_reg/NET0131 ,
		_w37732_
	);
	LUT2 #(
		.INIT('h8)
	) name27221 (
		\wishbone_TxBDRead_reg/NET0131 ,
		\wishbone_TxBDReady_reg/NET0131 ,
		_w37733_
	);
	LUT2 #(
		.INIT('h1)
	) name27222 (
		_w37732_,
		_w37733_,
		_w37734_
	);
	LUT2 #(
		.INIT('h4)
	) name27223 (
		mrxdv_pad_i_pad,
		_w34199_,
		_w37735_
	);
	LUT2 #(
		.INIT('h1)
	) name27224 (
		_w10584_,
		_w37735_,
		_w37736_
	);
	LUT2 #(
		.INIT('h1)
	) name27225 (
		\wishbone_BlockingIncrementTxPointer_reg/NET0131 ,
		\wishbone_IncrTxPointer_reg/NET0131 ,
		_w37737_
	);
	LUT2 #(
		.INIT('h2)
	) name27226 (
		_w12540_,
		_w37737_,
		_w37738_
	);
	LUT2 #(
		.INIT('h4)
	) name27227 (
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		\wishbone_TxUnderRun_sync1_reg/NET0131 ,
		_w37739_
	);
	LUT2 #(
		.INIT('h1)
	) name27228 (
		\wishbone_TxUnderRun_wb_reg/NET0131 ,
		_w37739_,
		_w37740_
	);
	LUT2 #(
		.INIT('h2)
	) name27229 (
		\miim1_EndBusy_reg/NET0131 ,
		\miim1_WCtrlDataStart_q_reg/NET0131 ,
		_w37741_
	);
	LUT2 #(
		.INIT('h1)
	) name27230 (
		_w28631_,
		_w37741_,
		_w37742_
	);
	LUT2 #(
		.INIT('h2)
	) name27231 (
		\maccontrol1_transmitcontrol1_BlockTxDone_reg/NET0131 ,
		\wishbone_TxStartFrm_reg/NET0131 ,
		_w37743_
	);
	LUT2 #(
		.INIT('h1)
	) name27232 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		_w37743_,
		_w37744_
	);
	LUT2 #(
		.INIT('h1)
	) name27233 (
		\wishbone_TxUnderRun_reg/NET0131 ,
		\wishbone_TxUnderRun_sync1_reg/NET0131 ,
		_w37745_
	);
	LUT2 #(
		.INIT('h1)
	) name27234 (
		\wishbone_BlockingTxStatusWrite_sync2_reg/NET0131 ,
		_w37745_,
		_w37746_
	);
	LUT2 #(
		.INIT('h2)
	) name27235 (
		\maccontrol1_transmitcontrol1_SendingCtrlFrm_reg/NET0131 ,
		\txethmac1_TxDone_reg/NET0131 ,
		_w37747_
	);
	LUT2 #(
		.INIT('h8)
	) name27236 (
		\maccontrol1_transmitcontrol1_TxCtrlStartFrm_reg/NET0131 ,
		\maccontrol1_transmitcontrol1_WillSendControlFrame_reg/NET0131 ,
		_w37748_
	);
	LUT2 #(
		.INIT('h1)
	) name27237 (
		_w37747_,
		_w37748_,
		_w37749_
	);
	LUT2 #(
		.INIT('h1)
	) name27238 (
		\miim1_outctrl_Mdo_2d_reg/NET0131 ,
		\miim1_shftrg_ShiftReg_reg[7]/NET0131 ,
		_w37750_
	);
	LUT2 #(
		.INIT('h8)
	) name27239 (
		\ethreg1_CTRLMODER_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_TXCTRL_2_DataOut_reg[0]/NET0131 ,
		_w37751_
	);
	LUT2 #(
		.INIT('h8)
	) name27240 (
		_w19087_,
		_w20125_,
		_w37752_
	);
	LUT2 #(
		.INIT('h2)
	) name27241 (
		_w18564_,
		_w37752_,
		_w37753_
	);
	LUT2 #(
		.INIT('h1)
	) name27242 (
		_w13475_,
		_w14019_,
		_w37754_
	);
	LUT2 #(
		.INIT('h1)
	) name27243 (
		_w14536_,
		_w15110_,
		_w37755_
	);
	LUT2 #(
		.INIT('h1)
	) name27244 (
		_w16743_,
		_w17287_,
		_w37756_
	);
	LUT2 #(
		.INIT('h1)
	) name27245 (
		_w17810_,
		_w19604_,
		_w37757_
	);
	LUT2 #(
		.INIT('h1)
	) name27246 (
		_w20856_,
		_w21383_,
		_w37758_
	);
	LUT2 #(
		.INIT('h1)
	) name27247 (
		_w21900_,
		_w22415_,
		_w37759_
	);
	LUT2 #(
		.INIT('h4)
	) name27248 (
		_w22932_,
		_w37759_,
		_w37760_
	);
	LUT2 #(
		.INIT('h8)
	) name27249 (
		_w37757_,
		_w37758_,
		_w37761_
	);
	LUT2 #(
		.INIT('h8)
	) name27250 (
		_w37755_,
		_w37756_,
		_w37762_
	);
	LUT2 #(
		.INIT('h4)
	) name27251 (
		_w37753_,
		_w37754_,
		_w37763_
	);
	LUT2 #(
		.INIT('h8)
	) name27252 (
		_w37762_,
		_w37763_,
		_w37764_
	);
	LUT2 #(
		.INIT('h8)
	) name27253 (
		_w37760_,
		_w37761_,
		_w37765_
	);
	LUT2 #(
		.INIT('h8)
	) name27254 (
		_w37764_,
		_w37765_,
		_w37766_
	);
	LUT2 #(
		.INIT('h8)
	) name27255 (
		_w12656_,
		_w15689_,
		_w37767_
	);
	LUT2 #(
		.INIT('h4)
	) name27256 (
		_w37766_,
		_w37767_,
		_w37768_
	);
	LUT2 #(
		.INIT('h2)
	) name27257 (
		\wishbone_TxBDReady_reg/NET0131 ,
		_w12656_,
		_w37769_
	);
	LUT2 #(
		.INIT('h8)
	) name27258 (
		_w34290_,
		_w37769_,
		_w37770_
	);
	LUT2 #(
		.INIT('h1)
	) name27259 (
		_w37768_,
		_w37770_,
		_w37771_
	);
	LUT2 #(
		.INIT('h1)
	) name27260 (
		\wishbone_RxPointerLSB_rst_reg[0]/NET0131 ,
		_w15696_,
		_w37772_
	);
	LUT2 #(
		.INIT('h2)
	) name27261 (
		_w15696_,
		_w24094_,
		_w37773_
	);
	LUT2 #(
		.INIT('h1)
	) name27262 (
		_w15698_,
		_w37772_,
		_w37774_
	);
	LUT2 #(
		.INIT('h4)
	) name27263 (
		_w37773_,
		_w37774_,
		_w37775_
	);
	LUT2 #(
		.INIT('h1)
	) name27264 (
		_w22944_,
		_w31141_,
		_w37776_
	);
	LUT2 #(
		.INIT('h8)
	) name27265 (
		\ethreg1_MAC_ADDR0_1_DataOut_reg[2]/NET0131 ,
		_w22959_,
		_w37777_
	);
	LUT2 #(
		.INIT('h8)
	) name27266 (
		\ethreg1_TXCTRL_1_DataOut_reg[2]/NET0131 ,
		_w23499_,
		_w37778_
	);
	LUT2 #(
		.INIT('h8)
	) name27267 (
		\ethreg1_MAC_ADDR1_1_DataOut_reg[2]/NET0131 ,
		_w23501_,
		_w37779_
	);
	LUT2 #(
		.INIT('h8)
	) name27268 (
		\ethreg1_MIIRX_DATA_DataOut_reg[10]/NET0131 ,
		_w23507_,
		_w37780_
	);
	LUT2 #(
		.INIT('h8)
	) name27269 (
		\ethreg1_RXHASH0_1_DataOut_reg[2]/NET0131 ,
		_w22952_,
		_w37781_
	);
	LUT2 #(
		.INIT('h8)
	) name27270 (
		\ethreg1_RXHASH1_1_DataOut_reg[2]/NET0131 ,
		_w22956_,
		_w37782_
	);
	LUT2 #(
		.INIT('h8)
	) name27271 (
		\ethreg1_MODER_1_DataOut_reg[2]/NET0131 ,
		_w23519_,
		_w37783_
	);
	LUT2 #(
		.INIT('h8)
	) name27272 (
		\ethreg1_PACKETLEN_1_DataOut_reg[2]/NET0131 ,
		_w22966_,
		_w37784_
	);
	LUT2 #(
		.INIT('h8)
	) name27273 (
		\ethreg1_MIIADDRESS_1_DataOut_reg[2]/NET0131 ,
		_w23513_,
		_w37785_
	);
	LUT2 #(
		.INIT('h8)
	) name27274 (
		\ethreg1_MIITX_DATA_1_DataOut_reg[2]/NET0131 ,
		_w23522_,
		_w37786_
	);
	LUT2 #(
		.INIT('h1)
	) name27275 (
		_w37777_,
		_w37778_,
		_w37787_
	);
	LUT2 #(
		.INIT('h1)
	) name27276 (
		_w37779_,
		_w37780_,
		_w37788_
	);
	LUT2 #(
		.INIT('h1)
	) name27277 (
		_w37781_,
		_w37782_,
		_w37789_
	);
	LUT2 #(
		.INIT('h1)
	) name27278 (
		_w37783_,
		_w37785_,
		_w37790_
	);
	LUT2 #(
		.INIT('h4)
	) name27279 (
		_w37786_,
		_w37790_,
		_w37791_
	);
	LUT2 #(
		.INIT('h8)
	) name27280 (
		_w37788_,
		_w37789_,
		_w37792_
	);
	LUT2 #(
		.INIT('h8)
	) name27281 (
		_w22944_,
		_w37787_,
		_w37793_
	);
	LUT2 #(
		.INIT('h8)
	) name27282 (
		_w37792_,
		_w37793_,
		_w37794_
	);
	LUT2 #(
		.INIT('h4)
	) name27283 (
		_w37784_,
		_w37791_,
		_w37795_
	);
	LUT2 #(
		.INIT('h8)
	) name27284 (
		_w37794_,
		_w37795_,
		_w37796_
	);
	LUT2 #(
		.INIT('h1)
	) name27285 (
		_w37776_,
		_w37796_,
		_w37797_
	);
	LUT2 #(
		.INIT('h1)
	) name27286 (
		\wishbone_RxPointerMSB_reg[10]/NET0131 ,
		_w17856_,
		_w37798_
	);
	LUT2 #(
		.INIT('h1)
	) name27287 (
		_w15696_,
		_w17857_,
		_w37799_
	);
	LUT2 #(
		.INIT('h4)
	) name27288 (
		_w37798_,
		_w37799_,
		_w37800_
	);
	LUT2 #(
		.INIT('h8)
	) name27289 (
		_w15696_,
		_w31141_,
		_w37801_
	);
	LUT2 #(
		.INIT('h1)
	) name27290 (
		_w37800_,
		_w37801_,
		_w37802_
	);
	LUT2 #(
		.INIT('h8)
	) name27291 (
		\ethreg1_INT_MASK_0_DataOut_reg[5]/NET0131 ,
		\ethreg1_irq_txc_reg/NET0131 ,
		_w37803_
	);
	LUT2 #(
		.INIT('h8)
	) name27292 (
		\ethreg1_INT_MASK_0_DataOut_reg[4]/NET0131 ,
		\ethreg1_irq_busy_reg/NET0131 ,
		_w37804_
	);
	LUT2 #(
		.INIT('h8)
	) name27293 (
		\ethreg1_INT_MASK_0_DataOut_reg[1]/NET0131 ,
		\ethreg1_irq_txe_reg/NET0131 ,
		_w37805_
	);
	LUT2 #(
		.INIT('h8)
	) name27294 (
		\ethreg1_INT_MASK_0_DataOut_reg[0]/NET0131 ,
		\ethreg1_irq_txb_reg/NET0131 ,
		_w37806_
	);
	LUT2 #(
		.INIT('h8)
	) name27295 (
		\ethreg1_INT_MASK_0_DataOut_reg[2]/NET0131 ,
		\ethreg1_irq_rxb_reg/NET0131 ,
		_w37807_
	);
	LUT2 #(
		.INIT('h8)
	) name27296 (
		\ethreg1_INT_MASK_0_DataOut_reg[6]/NET0131 ,
		\ethreg1_irq_rxc_reg/NET0131 ,
		_w37808_
	);
	LUT2 #(
		.INIT('h8)
	) name27297 (
		\ethreg1_INT_MASK_0_DataOut_reg[3]/NET0131 ,
		\ethreg1_irq_rxe_reg/NET0131 ,
		_w37809_
	);
	LUT2 #(
		.INIT('h1)
	) name27298 (
		_w37803_,
		_w37804_,
		_w37810_
	);
	LUT2 #(
		.INIT('h1)
	) name27299 (
		_w37805_,
		_w37806_,
		_w37811_
	);
	LUT2 #(
		.INIT('h1)
	) name27300 (
		_w37807_,
		_w37808_,
		_w37812_
	);
	LUT2 #(
		.INIT('h4)
	) name27301 (
		_w37809_,
		_w37812_,
		_w37813_
	);
	LUT2 #(
		.INIT('h8)
	) name27302 (
		_w37810_,
		_w37811_,
		_w37814_
	);
	LUT2 #(
		.INIT('h8)
	) name27303 (
		_w37813_,
		_w37814_,
		_w37815_
	);
	LUT2 #(
		.INIT('h2)
	) name27304 (
		\wishbone_tx_fifo_fifo_reg[2][15]/P0001 ,
		_w34464_,
		_w37816_
	);
	LUT2 #(
		.INIT('h8)
	) name27305 (
		\m_wb_dat_i[15]_pad ,
		_w34464_,
		_w37817_
	);
	LUT2 #(
		.INIT('h1)
	) name27306 (
		_w37816_,
		_w37817_,
		_w37818_
	);
	LUT2 #(
		.INIT('h2)
	) name27307 (
		\wishbone_tx_fifo_fifo_reg[2][16]/P0001 ,
		_w34464_,
		_w37819_
	);
	LUT2 #(
		.INIT('h8)
	) name27308 (
		\m_wb_dat_i[16]_pad ,
		_w34464_,
		_w37820_
	);
	LUT2 #(
		.INIT('h1)
	) name27309 (
		_w37819_,
		_w37820_,
		_w37821_
	);
	LUT2 #(
		.INIT('h2)
	) name27310 (
		\wishbone_tx_fifo_fifo_reg[2][17]/P0001 ,
		_w34464_,
		_w37822_
	);
	LUT2 #(
		.INIT('h8)
	) name27311 (
		\m_wb_dat_i[17]_pad ,
		_w34464_,
		_w37823_
	);
	LUT2 #(
		.INIT('h1)
	) name27312 (
		_w37822_,
		_w37823_,
		_w37824_
	);
	LUT2 #(
		.INIT('h2)
	) name27313 (
		\wishbone_tx_fifo_fifo_reg[2][22]/P0001 ,
		_w34464_,
		_w37825_
	);
	LUT2 #(
		.INIT('h8)
	) name27314 (
		\m_wb_dat_i[22]_pad ,
		_w34464_,
		_w37826_
	);
	LUT2 #(
		.INIT('h1)
	) name27315 (
		_w37825_,
		_w37826_,
		_w37827_
	);
	LUT2 #(
		.INIT('h2)
	) name27316 (
		\wishbone_tx_fifo_fifo_reg[2][23]/P0001 ,
		_w34464_,
		_w37828_
	);
	LUT2 #(
		.INIT('h8)
	) name27317 (
		\m_wb_dat_i[23]_pad ,
		_w34464_,
		_w37829_
	);
	LUT2 #(
		.INIT('h1)
	) name27318 (
		_w37828_,
		_w37829_,
		_w37830_
	);
	LUT2 #(
		.INIT('h2)
	) name27319 (
		\wishbone_tx_fifo_fifo_reg[2][25]/P0001 ,
		_w34464_,
		_w37831_
	);
	LUT2 #(
		.INIT('h8)
	) name27320 (
		\m_wb_dat_i[25]_pad ,
		_w34464_,
		_w37832_
	);
	LUT2 #(
		.INIT('h1)
	) name27321 (
		_w37831_,
		_w37832_,
		_w37833_
	);
	LUT2 #(
		.INIT('h2)
	) name27322 (
		\wishbone_tx_fifo_fifo_reg[2][2]/P0001 ,
		_w34464_,
		_w37834_
	);
	LUT2 #(
		.INIT('h8)
	) name27323 (
		\m_wb_dat_i[2]_pad ,
		_w34464_,
		_w37835_
	);
	LUT2 #(
		.INIT('h1)
	) name27324 (
		_w37834_,
		_w37835_,
		_w37836_
	);
	assign \_al_n1  = 1'b0;
	assign \g215539/_0_  = _w10562_ ;
	assign \g215543/_0_  = _w10572_ ;
	assign \g215547/_0_  = _w10581_ ;
	assign \g215551/_0_  = _w10663_ ;
	assign \g215552/_0_  = _w10674_ ;
	assign \g215578/_0_  = _w10678_ ;
	assign \g215587/_1_  = _w11117_ ;
	assign \g215589/_1_  = _w11128_ ;
	assign \g215591/_1_  = _w11132_ ;
	assign \g215593/_1_  = _w11135_ ;
	assign \g215595/_1_  = _w11139_ ;
	assign \g215597/_1_  = _w11143_ ;
	assign \g215599/_1_  = _w11147_ ;
	assign \g215601/_1_  = _w11151_ ;
	assign \g215603/_1_  = _w11155_ ;
	assign \g215605/_1_  = _w11158_ ;
	assign \g215607/_1_  = _w11162_ ;
	assign \g215609/_1_  = _w11165_ ;
	assign \g215611/_1_  = _w11168_ ;
	assign \g215613/_1_  = _w11171_ ;
	assign \g215615/_1_  = _w11174_ ;
	assign \g215617/_1_  = _w11177_ ;
	assign \g215618/_0_  = _w11182_ ;
	assign \g215619/_0_  = _w11183_ ;
	assign \g215620/_0_  = _w11224_ ;
	assign \g215632/_1_  = _w11226_ ;
	assign \g215634/_0_  = _w11240_ ;
	assign \g215635/_0_  = _w11248_ ;
	assign \g215636/_0_  = _w11249_ ;
	assign \g215637/_0_  = _w11252_ ;
	assign \g215638/_0_  = _w11256_ ;
	assign \g215639/_0_  = _w11259_ ;
	assign \g215655/_1_  = _w11272_ ;
	assign \g215657/_1_  = _w11278_ ;
	assign \g215659/_1_  = _w11282_ ;
	assign \g215661/_1_  = _w11285_ ;
	assign \g215662/_0_  = _w11318_ ;
	assign \g215663/_0_  = _w11335_ ;
	assign \g215664/_0_  = _w11353_ ;
	assign \g215665/_0_  = _w11356_ ;
	assign \g215668/_0_  = _w11358_ ;
	assign \g215674/_0_  = _w11372_ ;
	assign \g215677/_0_  = _w11377_ ;
	assign \g215686/_0_  = _w11386_ ;
	assign \g215695/_0_  = _w11389_ ;
	assign \g215696/_0_  = _w11393_ ;
	assign \g215702/_1__syn_2  = _w11386_ ;
	assign \g215705/_0_  = _w11398_ ;
	assign \g215706/_0_  = _w11399_ ;
	assign \g215716/_0_  = _w11404_ ;
	assign \g215717/_0_  = _w11418_ ;
	assign \g215718/_0_  = _w11426_ ;
	assign \g215726/_0_  = _w11431_ ;
	assign \g215727/_0_  = _w11435_ ;
	assign \g215728/_0_  = _w11443_ ;
	assign \g215760/_0_  = _w11447_ ;
	assign \g215764/_0_  = _w11617_ ;
	assign \g215765/_0_  = _w11650_ ;
	assign \g215766/_0_  = _w11655_ ;
	assign \g215767/_3_  = _w11666_ ;
	assign \g215768/_3_  = _w11674_ ;
	assign \g215769/_3_  = _w11679_ ;
	assign \g215770/_3_  = _w11684_ ;
	assign \g215771/_3_  = _w11689_ ;
	assign \g215772/_3_  = _w11694_ ;
	assign \g215773/_3_  = _w11699_ ;
	assign \g215774/_3_  = _w11704_ ;
	assign \g215775/_3_  = _w11710_ ;
	assign \g215776/_3_  = _w11715_ ;
	assign \g215777/_3_  = _w11721_ ;
	assign \g215778/_3_  = _w11726_ ;
	assign \g215779/_3_  = _w11731_ ;
	assign \g215780/_3_  = _w11736_ ;
	assign \g215790/_0_  = _w11747_ ;
	assign \g215791/_0_  = _w11751_ ;
	assign \g215792/_0_  = _w11755_ ;
	assign \g215793/_0_  = _w11756_ ;
	assign \g215801/_0_  = _w11763_ ;
	assign \g215802/_0_  = _w11771_ ;
	assign \g215803/_0_  = _w11775_ ;
	assign \g215804/_0_  = _w11776_ ;
	assign \g215812/_0_  = _w11781_ ;
	assign \g215813/_0_  = _w11785_ ;
	assign \g215821/_0_  = _w11801_ ;
	assign \g215823/_0_  = _w11805_ ;
	assign \g215831/_0_  = _w11809_ ;
	assign \g215832/_0_  = _w11813_ ;
	assign \g215833/_0_  = _w11817_ ;
	assign \g215845/_0_  = _w11822_ ;
	assign \g215846/_0_  = _w11826_ ;
	assign \g215847/_0_  = _w12064_ ;
	assign \g215872/_0_  = _w12068_ ;
	assign \g215873/_0_  = _w12103_ ;
	assign \g215874/_0_  = _w12111_ ;
	assign \g215904/_0_  = _w12119_ ;
	assign \g215905/_0_  = _w12145_ ;
	assign \g215906/_0_  = _w12153_ ;
	assign \g215907/_0_  = _w12157_ ;
	assign \g215908/_0_  = _w12162_ ;
	assign \g215909/_0_  = _w12165_ ;
	assign \g215910/_0_  = _w12169_ ;
	assign \g215911/_0_  = _w12173_ ;
	assign \g215912/_0_  = _w12176_ ;
	assign \g215913/_0_  = _w12181_ ;
	assign \g215914/_0_  = _w12185_ ;
	assign \g215915/_0_  = _w12189_ ;
	assign \g215916/_0_  = _w12193_ ;
	assign \g215917/_0_  = _w12197_ ;
	assign \g215918/_0_  = _w12200_ ;
	assign \g215919/_0_  = _w12203_ ;
	assign \g215920/_0_  = _w12206_ ;
	assign \g215923/_0_  = _w12214_ ;
	assign \g215926/_0_  = _w12217_ ;
	assign \g215941/_0_  = _w12230_ ;
	assign \g215942/_0_  = _w12233_ ;
	assign \g215943/_0_  = _w12236_ ;
	assign \g215944/_0_  = _w12239_ ;
	assign \g215945/_0_  = _w12275_ ;
	assign \g215946/_0_  = _w12298_ ;
	assign \g215947/_0_  = _w12321_ ;
	assign \g215948/_0_  = _w12344_ ;
	assign \g215949/_0_  = _w12367_ ;
	assign \g215950/_0_  = _w12390_ ;
	assign \g215951/_0_  = _w12413_ ;
	assign \g215952/_0_  = _w12436_ ;
	assign \g215953/_0_  = _w12440_ ;
	assign \g215954/_0_  = _w12443_ ;
	assign \g215955/_0_  = _w12445_ ;
	assign \g215956/_0_  = _w12462_ ;
	assign \g215957/_0_  = _w12476_ ;
	assign \g215959/_00_  = _w12494_ ;
	assign \g215960/_0_  = _w12497_ ;
	assign \g215962/_0_  = _w12500_ ;
	assign \g215964/_0_  = _w12529_ ;
	assign \g215966/_0_  = _w12531_ ;
	assign \g215972/_0_  = _w12539_ ;
	assign \g216035/_0_  = _w12640_ ;
	assign \g216037/_0_  = _w12654_ ;
	assign \g216038/_0_  = _w13504_ ;
	assign \g216039/_0_  = _w14024_ ;
	assign \g216040/_0_  = _w14543_ ;
	assign \g216041/_0_  = _w14547_ ;
	assign \g216042/_0_  = _w14551_ ;
	assign \g216046/_0_  = _w14585_ ;
	assign \g216048/_0_  = _w14598_ ;
	assign \g216057/_0_  = _w15121_ ;
	assign \g216263/_0_  = _w15134_ ;
	assign \g216264/_0_  = _w15156_ ;
	assign \g216265/_0_  = _w15159_ ;
	assign \g216266/_0_  = _w15162_ ;
	assign \g216267/_0_  = _w15165_ ;
	assign \g216268/_0_  = _w15168_ ;
	assign \g216269/_0_  = _w15171_ ;
	assign \g216270/_0_  = _w15174_ ;
	assign \g216271/_0_  = _w15692_ ;
	assign \g216272/_0_  = _w15695_ ;
	assign \g216273/_0_  = _w16213_ ;
	assign \g216284/_0_  = _w16217_ ;
	assign \g216289/_0_  = _w16221_ ;
	assign \g216290/_0_  = _w16231_ ;
	assign \g216292/_0_  = _w16775_ ;
	assign \g216296/_0_  = _w17298_ ;
	assign \g216297/_0_  = _w17821_ ;
	assign \g216300/_0_  = _w17826_ ;
	assign \g216301/_0_  = _w17829_ ;
	assign \g216302/_0_  = _w17832_ ;
	assign \g216303/_0_  = _w17835_ ;
	assign \g216304/_0_  = _w17838_ ;
	assign \g216305/_0_  = _w17841_ ;
	assign \g216306/_0_  = _w17844_ ;
	assign \g216307/_0_  = _w17847_ ;
	assign \g216310/_3_  = _w17882_ ;
	assign \g216311/_3_  = _w17920_ ;
	assign \g216314/u3_syn_7  = _w15147_ ;
	assign \g216322/_3_  = _w17926_ ;
	assign \g216323/_3_  = _w17929_ ;
	assign \g216324/_3_  = _w17932_ ;
	assign \g216325/_3_  = _w17935_ ;
	assign \g216326/_3_  = _w17938_ ;
	assign \g216327/_3_  = _w17941_ ;
	assign \g216328/_3_  = _w17944_ ;
	assign \g216329/_3_  = _w17947_ ;
	assign \g216369/_0_  = _w17960_ ;
	assign \g216370/_0_  = _w17973_ ;
	assign \g216371/_0_  = _w17982_ ;
	assign \g216372/_0_  = _w17994_ ;
	assign \g216373/_0_  = _w18005_ ;
	assign \g216374/_0_  = _w18014_ ;
	assign \g216375/_0_  = _w18026_ ;
	assign \g216376/_0_  = _w18039_ ;
	assign \g216379/_0_  = _w18052_ ;
	assign \g216380/_0_  = _w18572_ ;
	assign \g216381/_0_  = _w18573_ ;
	assign \g216385/_0_  = _w19092_ ;
	assign \g216389/_0_  = _w19609_ ;
	assign \g216390/_0_  = _w20130_ ;
	assign \g216402/_0_  = _w20133_ ;
	assign \g216404/_0_  = _w20137_ ;
	assign \g216405/_0_  = _w20149_ ;
	assign \g216406/_0_  = _w20161_ ;
	assign \g216407/_0_  = _w20173_ ;
	assign \g216408/_0_  = _w20185_ ;
	assign \g216409/_0_  = _w20197_ ;
	assign \g216410/_0_  = _w20209_ ;
	assign \g216411/_0_  = _w20218_ ;
	assign \g216412/_0_  = _w20231_ ;
	assign \g216413/_0_  = _w20241_ ;
	assign \g216414/_0_  = _w20253_ ;
	assign \g216415/_0_  = _w20270_ ;
	assign \g216416/_0_  = _w20282_ ;
	assign \g216417/_0_  = _w20294_ ;
	assign \g216418/_0_  = _w20303_ ;
	assign \g216419/_0_  = _w20312_ ;
	assign \g216420/_0_  = _w20321_ ;
	assign \g216421/_0_  = _w20330_ ;
	assign \g216422/_0_  = _w20339_ ;
	assign \g216423/_0_  = _w20341_ ;
	assign \g216424/_0_  = _w20343_ ;
	assign \g216425/_0_  = _w20858_ ;
	assign \g216426/_0_  = _w20860_ ;
	assign \g216427/_0_  = _w20862_ ;
	assign \g216428/_0_  = _w20864_ ;
	assign \g216429/_0_  = _w20866_ ;
	assign \g216430/_0_  = _w20868_ ;
	assign \g216431/_0_  = _w20870_ ;
	assign \g216432/_0_  = _w21385_ ;
	assign \g216433/_0_  = _w21387_ ;
	assign \g216434/_0_  = _w21902_ ;
	assign \g216435/_0_  = _w22417_ ;
	assign \g216436/_0_  = _w22419_ ;
	assign \g216437/_0_  = _w22934_ ;
	assign \g216438/_0_  = _w22936_ ;
	assign \g216439/_3_  = _w22972_ ;
	assign \g216447/_3_  = _w22982_ ;
	assign \g216448/_3_  = _w23534_ ;
	assign \g216452/_0_  = _w23551_ ;
	assign \g216453/_0_  = _w23577_ ;
	assign \g216454/_0_  = _w23580_ ;
	assign \g216455/_0_  = _w24096_ ;
	assign \g216456/_0_  = _w24098_ ;
	assign \g216457/_0_  = _w24100_ ;
	assign \g216458/_3_  = _w24110_ ;
	assign \g216459/_3_  = _w24120_ ;
	assign \g216461/_3_  = _w24130_ ;
	assign \g216462/_3_  = _w24140_ ;
	assign \g216463/_3_  = _w24150_ ;
	assign \g216464/_3_  = _w24160_ ;
	assign \g216465/_3_  = _w24170_ ;
	assign \g216466/_0_  = _w24172_ ;
	assign \g216467/_3_  = _w24182_ ;
	assign \g216468/_3_  = _w24192_ ;
	assign \g216469/_3_  = _w24754_ ;
	assign \g216470/_3_  = _w25304_ ;
	assign \g216471/_3_  = _w25852_ ;
	assign \g216473/_3_  = _w26388_ ;
	assign \g216474/_3_  = _w26924_ ;
	assign \g216475/_3_  = _w27458_ ;
	assign \g216476/_3_  = _w27468_ ;
	assign \g216477/_3_  = _w28002_ ;
	assign \g216478/_0_  = _w28008_ ;
	assign \g216479/_3_  = _w28568_ ;
	assign \g216480/_3_  = _w28612_ ;
	assign \g216481/_3_  = _w28664_ ;
	assign \g216492/_0_  = _w28669_ ;
	assign \g216494/_0_  = _w28690_ ;
	assign \g216495/_3_  = _w28706_ ;
	assign \g216496/_3_  = _w29252_ ;
	assign \g216498/_3_  = _w29264_ ;
	assign \g216499/_3_  = _w29276_ ;
	assign \g216500/_3_  = _w29288_ ;
	assign \g216513/_3_  = _w29296_ ;
	assign \g216514/_3_  = _w29301_ ;
	assign \g216515/_3_  = _w29307_ ;
	assign \g216516/_3_  = _w29312_ ;
	assign \g216517/_3_  = _w29317_ ;
	assign \g216518/_3_  = _w29322_ ;
	assign \g216519/_3_  = _w29327_ ;
	assign \g216520/_3_  = _w29333_ ;
	assign \g216521/_3_  = _w29339_ ;
	assign \g216522/_3_  = _w29344_ ;
	assign \g216523/_3_  = _w29349_ ;
	assign \g216524/_3_  = _w29355_ ;
	assign \g216525/_3_  = _w29361_ ;
	assign \g216526/_3_  = _w29367_ ;
	assign \g216527/_3_  = _w29372_ ;
	assign \g216528/_3_  = _w29378_ ;
	assign \g216529/_3_  = _w29383_ ;
	assign \g216530/_3_  = _w29389_ ;
	assign \g216531/_3_  = _w29394_ ;
	assign \g216532/_3_  = _w29400_ ;
	assign \g216533/_3_  = _w29405_ ;
	assign \g216534/_3_  = _w29411_ ;
	assign \g216535/_3_  = _w29417_ ;
	assign \g216536/_3_  = _w29422_ ;
	assign \g216537/_3_  = _w29430_ ;
	assign \g216538/_3_  = _w29435_ ;
	assign \g216555/_3_  = _w29967_ ;
	assign \g216556/_3_  = _w30499_ ;
	assign \g216557/_3_  = _w30519_ ;
	assign \g216560/_3_  = _w30525_ ;
	assign \g216561/_3_  = _w30530_ ;
	assign \g216562/_3_  = _w30535_ ;
	assign \g216563/_3_  = _w30540_ ;
	assign \g216564/_3_  = _w30545_ ;
	assign \g216565/_3_  = _w30550_ ;
	assign \g216566/_3_  = _w30555_ ;
	assign \g216567/_3_  = _w30561_ ;
	assign \g216568/_3_  = _w30566_ ;
	assign \g216569/_3_  = _w30571_ ;
	assign \g216570/_3_  = _w30576_ ;
	assign \g216571/_3_  = _w30581_ ;
	assign \g216575/_3_  = _w30586_ ;
	assign \g216576/_3_  = _w30591_ ;
	assign \g216577/_3_  = _w30596_ ;
	assign \g216578/_3_  = _w30601_ ;
	assign \g216579/_3_  = _w30606_ ;
	assign \g216580/_3_  = _w30611_ ;
	assign \g216581/_3_  = _w30616_ ;
	assign \g216582/_3_  = _w30621_ ;
	assign \g216583/_3_  = _w30626_ ;
	assign \g216586/_3_  = _w31143_ ;
	assign \g216587/_3_  = _w31148_ ;
	assign \g216588/_3_  = _w31153_ ;
	assign \g216589/_3_  = _w31159_ ;
	assign \g216590/_3_  = _w31164_ ;
	assign \g216591/_3_  = _w31169_ ;
	assign \g216592/_3_  = _w31174_ ;
	assign \g216593/_3_  = _w31179_ ;
	assign \g216594/_3_  = _w31184_ ;
	assign \g216595/_3_  = _w31189_ ;
	assign \g216600/_3_  = _w31211_ ;
	assign \g216683/_0_  = _w31221_ ;
	assign \g216689/_0_  = _w31224_ ;
	assign \g216693/_0_  = _w31237_ ;
	assign \g216694/_0_  = _w31247_ ;
	assign \g216727/_0_  = _w31250_ ;
	assign \g216728/_0_  = _w31253_ ;
	assign \g216729/_0_  = _w31256_ ;
	assign \g216732/_0_  = _w31259_ ;
	assign \g216733/_0_  = _w31263_ ;
	assign \g216734/_0_  = _w31269_ ;
	assign \g216735/_0_  = _w31273_ ;
	assign \g216736/_0_  = _w31276_ ;
	assign \g216737/_0_  = _w31279_ ;
	assign \g216738/_0_  = _w31282_ ;
	assign \g216739/_0_  = _w31286_ ;
	assign \g216740/_0_  = _w31290_ ;
	assign \g216741/_0_  = _w31294_ ;
	assign \g216742/_0_  = _w31298_ ;
	assign \g216743/_0_  = _w31301_ ;
	assign \g216744/_0_  = _w31306_ ;
	assign \g216745/_0_  = _w31310_ ;
	assign \g216746/_0_  = _w31314_ ;
	assign \g216748/_0_  = _w31332_ ;
	assign \g216751/_0_  = _w31342_ ;
	assign \g216754/_0_  = _w31352_ ;
	assign \g216762/_0_  = _w31355_ ;
	assign \g216934/_2_  = _w31357_ ;
	assign \g216952/_0_  = _w31375_ ;
	assign \g216955/_0_  = _w31377_ ;
	assign \g216969/_0_  = _w31385_ ;
	assign \g216979/_0_  = _w31388_ ;
	assign \g216984/_0_  = _w31390_ ;
	assign \g216996/_0_  = _w31393_ ;
	assign \g217002/_0_  = _w31400_ ;
	assign \g217014/_0_  = _w31437_ ;
	assign \g217015/_0_  = _w31449_ ;
	assign \g217016/_0_  = _w31461_ ;
	assign \g217017/_0_  = _w31473_ ;
	assign \g217018/_0_  = _w31485_ ;
	assign \g217019/_0_  = _w31496_ ;
	assign \g217023/_0_  = _w31499_ ;
	assign \g217116/_0_  = _w31681_ ;
	assign \g217146/_3_  = _w31722_ ;
	assign \g217149/_0_  = _w31723_ ;
	assign \g217151/_0_  = _w31727_ ;
	assign \g217160/_0_  = _w31733_ ;
	assign \g217167/_0_  = _w31737_ ;
	assign \g217168/_0_  = _w31742_ ;
	assign \g217169/_0_  = _w31747_ ;
	assign \g217170/_0_  = _w31751_ ;
	assign \g217171/_0_  = _w31755_ ;
	assign \g217172/_0_  = _w31759_ ;
	assign \g217173/_0_  = _w31763_ ;
	assign \g217174/_0_  = _w31767_ ;
	assign \g217175/_0_  = _w31771_ ;
	assign \g217176/_0_  = _w31775_ ;
	assign \g217177/_0_  = _w31779_ ;
	assign \g217178/_0_  = _w31783_ ;
	assign \g217179/_0_  = _w31787_ ;
	assign \g217180/_0_  = _w31791_ ;
	assign \g217181/_0_  = _w31795_ ;
	assign \g217182/_0_  = _w31799_ ;
	assign \g217183/_0_  = _w31803_ ;
	assign \g217187/_0_  = _w31809_ ;
	assign \g217188/_0_  = _w31811_ ;
	assign \g217189/_0_  = _w31816_ ;
	assign \g217193/_0_  = _w31819_ ;
	assign \g217194/_0_  = _w31821_ ;
	assign \g217195/_0_  = _w31848_ ;
	assign \g217196/_0_  = _w31856_ ;
	assign \g217202/_0_  = _w31858_ ;
	assign \g217205/_0_  = _w31863_ ;
	assign \g217206/_0_  = _w31866_ ;
	assign \g217207/_0_  = _w31869_ ;
	assign \g217208/_0_  = _w31872_ ;
	assign \g217209/_0_  = _w31875_ ;
	assign \g217210/_0_  = _w31878_ ;
	assign \g217211/_0_  = _w31881_ ;
	assign \g217212/_0_  = _w31884_ ;
	assign \g217213/_0_  = _w31887_ ;
	assign \g217214/_0_  = _w31890_ ;
	assign \g217215/_0_  = _w31893_ ;
	assign \g217216/_0_  = _w31896_ ;
	assign \g217217/_0_  = _w31899_ ;
	assign \g217218/_0_  = _w31902_ ;
	assign \g217219/_0_  = _w31905_ ;
	assign \g217220/_0_  = _w31908_ ;
	assign \g217223/_0_  = _w31915_ ;
	assign \g217231/_0_  = _w31921_ ;
	assign \g217237/_0_  = _w31931_ ;
	assign \g217238/_0_  = _w31941_ ;
	assign \g217242/_0_  = _w31944_ ;
	assign \g217243/_0_  = _w31949_ ;
	assign \g217250/_3_  = _w32007_ ;
	assign \g217251/_3_  = _w32041_ ;
	assign \g217252/_3_  = _w32073_ ;
	assign \g217253/_3_  = _w32107_ ;
	assign \g217254/_3_  = _w32139_ ;
	assign \g217255/_3_  = _w32173_ ;
	assign \g217256/_3_  = _w32205_ ;
	assign \g217257/_3_  = _w32239_ ;
	assign \g217258/_3_  = _w32271_ ;
	assign \g217259/_3_  = _w32303_ ;
	assign \g217260/_3_  = _w32335_ ;
	assign \g217261/_3_  = _w32369_ ;
	assign \g217262/_3_  = _w32403_ ;
	assign \g217263/_3_  = _w32435_ ;
	assign \g217264/_3_  = _w32467_ ;
	assign \g217265/_3_  = _w32499_ ;
	assign \g217266/_3_  = _w32531_ ;
	assign \g217267/_3_  = _w32563_ ;
	assign \g217268/_3_  = _w32595_ ;
	assign \g217269/_3_  = _w32629_ ;
	assign \g217270/_3_  = _w32663_ ;
	assign \g217271/_3_  = _w32697_ ;
	assign \g217272/_3_  = _w32729_ ;
	assign \g217273/_3_  = _w32761_ ;
	assign \g217274/_3_  = _w32795_ ;
	assign \g217275/_3_  = _w32827_ ;
	assign \g217276/_3_  = _w32861_ ;
	assign \g217277/_3_  = _w32895_ ;
	assign \g217278/_3_  = _w32927_ ;
	assign \g217279/_3_  = _w32961_ ;
	assign \g217280/_3_  = _w32993_ ;
	assign \g217281/_3_  = _w33027_ ;
	assign \g217282/_3_  = _w33085_ ;
	assign \g217283/_3_  = _w33117_ ;
	assign \g217284/_3_  = _w33149_ ;
	assign \g217285/_3_  = _w33181_ ;
	assign \g217286/_3_  = _w33213_ ;
	assign \g217287/_3_  = _w33245_ ;
	assign \g217288/_3_  = _w33277_ ;
	assign \g217289/_3_  = _w33309_ ;
	assign \g217290/_3_  = _w33341_ ;
	assign \g217291/_3_  = _w33373_ ;
	assign \g217292/_3_  = _w33405_ ;
	assign \g217293/_3_  = _w33437_ ;
	assign \g217294/_3_  = _w33469_ ;
	assign \g217295/_3_  = _w33501_ ;
	assign \g217296/_3_  = _w33533_ ;
	assign \g217297/_3_  = _w33565_ ;
	assign \g217298/_3_  = _w33597_ ;
	assign \g217299/_3_  = _w33629_ ;
	assign \g217300/_3_  = _w33661_ ;
	assign \g217301/_3_  = _w33693_ ;
	assign \g217302/_3_  = _w33725_ ;
	assign \g217303/_3_  = _w33757_ ;
	assign \g217304/_3_  = _w33789_ ;
	assign \g217305/_3_  = _w33821_ ;
	assign \g217306/_3_  = _w33853_ ;
	assign \g217307/_3_  = _w33885_ ;
	assign \g217308/_3_  = _w33917_ ;
	assign \g217309/_3_  = _w33949_ ;
	assign \g217310/_3_  = _w33981_ ;
	assign \g217311/_3_  = _w34013_ ;
	assign \g217312/_3_  = _w34045_ ;
	assign \g217313/_3_  = _w34077_ ;
	assign \g217318/_0_  = _w34081_ ;
	assign \g217662/_0_  = _w34101_ ;
	assign \g217663/_0_  = _w34105_ ;
	assign \g217682/_0_  = _w34119_ ;
	assign \g217697/_0_  = _w34130_ ;
	assign \g217698/_0_  = _w34149_ ;
	assign \g217699/_0_  = _w34156_ ;
	assign \g217700/_0_  = _w34159_ ;
	assign \g217701/_0_  = _w34161_ ;
	assign \g217705/_0_  = _w34169_ ;
	assign \g217711/_0_  = _w34173_ ;
	assign \g217747/_0_  = _w34178_ ;
	assign \g217753/_00_  = _w34181_ ;
	assign \g217775/_0_  = _w34198_ ;
	assign \g217781/_0_  = _w34213_ ;
	assign \g217784/_0_  = _w34215_ ;
	assign \g217785/_0_  = _w34220_ ;
	assign \g217786/_0_  = _w34225_ ;
	assign \g217787/_0_  = _w34230_ ;
	assign \g217788/_0_  = _w34235_ ;
	assign \g217790/_0_  = _w34240_ ;
	assign \g217815/_0_  = _w34247_ ;
	assign \g217817/_0_  = _w34250_ ;
	assign \g218145/_0_  = _w34252_ ;
	assign \g218148/_0_  = _w34256_ ;
	assign \g218150/_0_  = _w34282_ ;
	assign \g218167/_0_  = _w34293_ ;
	assign \g218168/_0_  = _w34296_ ;
	assign \g218234/_0_  = _w34297_ ;
	assign \g218235/_0_  = _w34298_ ;
	assign \g218236/_0_  = _w34302_ ;
	assign \g218238/_0_  = _w34308_ ;
	assign \g218242/_0_  = _w34311_ ;
	assign \g218332/_0_  = _w34318_ ;
	assign \g218335/_0_  = _w34327_ ;
	assign \g218336/_0_  = _w34336_ ;
	assign \g218337/_0_  = _w34346_ ;
	assign \g218338/_0_  = _w34350_ ;
	assign \g218339/_0_  = _w34354_ ;
	assign \g218340/_0_  = _w34358_ ;
	assign \g218341/_0_  = _w34362_ ;
	assign \g218342/_0_  = _w34366_ ;
	assign \g218343/_0_  = _w34376_ ;
	assign \g218344/_0_  = _w34380_ ;
	assign \g218345/_0_  = _w34383_ ;
	assign \g218346/_0_  = _w34386_ ;
	assign \g218347/_0_  = _w34389_ ;
	assign \g218348/_0_  = _w34392_ ;
	assign \g218349/_0_  = _w34395_ ;
	assign \g218350/_0_  = _w34398_ ;
	assign \g218351/_0_  = _w34405_ ;
	assign \g218352/_0_  = _w34408_ ;
	assign \g218353/_0_  = _w34411_ ;
	assign \g218354/_0_  = _w34414_ ;
	assign \g218355/_0_  = _w34417_ ;
	assign \g218356/_0_  = _w34420_ ;
	assign \g218357/_0_  = _w34423_ ;
	assign \g218358/_0_  = _w34426_ ;
	assign \g218359/_0_  = _w34429_ ;
	assign \g218360/_0_  = _w34432_ ;
	assign \g218398/_3_  = _w34435_ ;
	assign \g218430/_0_  = _w34439_ ;
	assign \g218440/_0_  = _w34444_ ;
	assign \g218452/u3_syn_4  = _w34451_ ;
	assign \g218495/u3_syn_4  = _w34455_ ;
	assign \g218517/u3_syn_4  = _w34457_ ;
	assign \g218554/u3_syn_4  = _w34462_ ;
	assign \g218575/u3_syn_4  = _w34464_ ;
	assign \g218600/u3_syn_4  = _w34466_ ;
	assign \g218621/u3_syn_4  = _w34467_ ;
	assign \g218638/u3_syn_4  = _w34468_ ;
	assign \g218659/u3_syn_4  = _w34472_ ;
	assign \g218673/u3_syn_4  = _w34476_ ;
	assign \g218707/u3_syn_4  = _w34479_ ;
	assign \g218735/_3_  = _w34482_ ;
	assign \g219186/_0_  = _w34491_ ;
	assign \g219187/_0_  = _w34494_ ;
	assign \g219188/_0_  = _w34497_ ;
	assign \g219189/_0_  = _w34502_ ;
	assign \g219190/_0_  = _w34513_ ;
	assign \g219196/_0_  = _w34518_ ;
	assign \g219198/_0_  = _w34524_ ;
	assign \g219199/_0_  = _w34531_ ;
	assign \g219200/_0_  = _w34535_ ;
	assign \g219308/_0_  = _w34540_ ;
	assign \g219314/_0_  = _w34544_ ;
	assign \g219326/_0_  = _w34546_ ;
	assign \g219328/_0_  = _w34549_ ;
	assign \g219348/_0_  = _w34560_ ;
	assign \g219351/_0_  = _w34562_ ;
	assign \g219363/_0_  = _w34565_ ;
	assign \g219364/_0_  = _w34570_ ;
	assign \g219365/_0_  = _w34573_ ;
	assign \g219366/_0_  = _w34576_ ;
	assign \g219367/_0_  = _w34579_ ;
	assign \g219368/_0_  = _w34582_ ;
	assign \g219369/_0_  = _w34585_ ;
	assign \g219376/_0_  = _w34589_ ;
	assign \g219381/_0_  = _w34592_ ;
	assign \g219382/_0_  = _w34599_ ;
	assign \g219384/_0_  = _w34605_ ;
	assign \g219385/_0_  = _w34614_ ;
	assign \g219391/_0_  = _w34620_ ;
	assign \g219394/_0_  = _w34626_ ;
	assign \g219395/_0_  = _w34629_ ;
	assign \g219396/_0_  = _w34632_ ;
	assign \g219397/_0_  = _w34635_ ;
	assign \g219398/_0_  = _w34638_ ;
	assign \g219399/_0_  = _w34642_ ;
	assign \g219400/_0_  = _w34645_ ;
	assign \g219401/_0_  = _w34648_ ;
	assign \g219402/_0_  = _w34651_ ;
	assign \g219403/_0_  = _w34654_ ;
	assign \g219404/_0_  = _w34657_ ;
	assign \g219405/_0_  = _w34660_ ;
	assign \g219406/_0_  = _w34663_ ;
	assign \g219407/_0_  = _w34666_ ;
	assign \g219408/_0_  = _w34669_ ;
	assign \g219409/_0_  = _w34674_ ;
	assign \g219410/_0_  = _w34677_ ;
	assign \g219411/_0_  = _w34680_ ;
	assign \g219412/_0_  = _w34683_ ;
	assign \g219413/_0_  = _w34686_ ;
	assign \g219414/_0_  = _w34689_ ;
	assign \g219415/_0_  = _w34692_ ;
	assign \g219416/_0_  = _w34695_ ;
	assign \g219417/_0_  = _w34698_ ;
	assign \g219418/_0_  = _w34701_ ;
	assign \g219419/_0_  = _w34704_ ;
	assign \g219420/_0_  = _w34708_ ;
	assign \g219421/_0_  = _w34711_ ;
	assign \g219422/_0_  = _w34714_ ;
	assign \g219423/_0_  = _w34717_ ;
	assign \g219424/_0_  = _w34720_ ;
	assign \g219425/_0_  = _w34723_ ;
	assign \g219426/_0_  = _w34726_ ;
	assign \g219427/_0_  = _w34729_ ;
	assign \g219428/_0_  = _w34732_ ;
	assign \g219429/_0_  = _w34735_ ;
	assign \g219430/_0_  = _w34738_ ;
	assign \g219431/_0_  = _w34743_ ;
	assign \g219432/_0_  = _w34746_ ;
	assign \g219433/_0_  = _w34749_ ;
	assign \g219434/_0_  = _w34752_ ;
	assign \g219435/_0_  = _w34755_ ;
	assign \g219436/_0_  = _w34758_ ;
	assign \g219437/_0_  = _w34761_ ;
	assign \g219438/_0_  = _w34764_ ;
	assign \g219439/_0_  = _w34767_ ;
	assign \g219440/_0_  = _w34770_ ;
	assign \g219441/_0_  = _w34773_ ;
	assign \g219442/_0_  = _w34776_ ;
	assign \g219443/_0_  = _w34779_ ;
	assign \g219444/_0_  = _w34782_ ;
	assign \g219445/_0_  = _w34785_ ;
	assign \g219446/_0_  = _w34788_ ;
	assign \g219447/_0_  = _w34791_ ;
	assign \g219449/_0_  = _w34796_ ;
	assign \g219450/_0_  = _w34799_ ;
	assign \g219451/_0_  = _w34802_ ;
	assign \g219452/_0_  = _w34805_ ;
	assign \g219453/_0_  = _w34808_ ;
	assign \g219454/_0_  = _w34811_ ;
	assign \g219455/_0_  = _w34814_ ;
	assign \g219456/_0_  = _w34817_ ;
	assign \g219457/_0_  = _w34820_ ;
	assign \g219458/_0_  = _w34823_ ;
	assign \g219464/u3_syn_7  = _w34825_ ;
	assign \g219496/u3_syn_4  = _w34826_ ;
	assign \g219512/u3_syn_4  = _w34457_ ;
	assign \g219526/u3_syn_4  = _w34828_ ;
	assign \g219549/u3_syn_4  = _w34829_ ;
	assign \g219571/u3_syn_4  = _w34462_ ;
	assign \g219588/u3_syn_4  = _w34467_ ;
	assign \g219603/u3_syn_4  = _w34476_ ;
	assign \g219621/u3_syn_4  = _w34830_ ;
	assign \g219636/_3_  = _w34834_ ;
	assign \g219652/u3_syn_4  = _w34837_ ;
	assign \g219676/_3_  = _w34841_ ;
	assign \g219686/_0_  = _w34844_ ;
	assign \g219689/_0_  = _w11469_ ;
	assign \g219694/_3_  = _w11484_ ;
	assign \g220062/_0_  = _w34845_ ;
	assign \g220068/_0_  = _w34846_ ;
	assign \g220069/_0_  = _w34847_ ;
	assign \g220072/_0_  = _w34854_ ;
	assign \g220084/_0_  = _w34856_ ;
	assign \g220149/_0_  = _w34868_ ;
	assign \g220162/_0_  = _w34875_ ;
	assign \g220317/_0_  = _w34878_ ;
	assign \g220360/_2_  = _w11759_ ;
	assign \g220368/_2_  = _w34880_ ;
	assign \g220369/_0_  = _w34903_ ;
	assign \g220370/_0_  = _w34910_ ;
	assign \g220371/_0_  = _w34914_ ;
	assign \g220372/_0_  = _w34922_ ;
	assign \g220376/_0_  = _w34933_ ;
	assign \g220390/_0_  = _w34967_ ;
	assign \g220395/_0_  = _w34974_ ;
	assign \g220499/_0_  = _w34997_ ;
	assign \g220500/_0_  = _w35004_ ;
	assign \g220501/_0_  = _w35011_ ;
	assign \g220502/_0_  = _w35018_ ;
	assign \g220503/_0_  = _w35025_ ;
	assign \g220504/_0_  = _w35032_ ;
	assign \g220505/_0_  = _w35039_ ;
	assign \g220506/_0_  = _w35046_ ;
	assign \g220507/_0_  = _w35053_ ;
	assign \g220508/_0_  = _w35060_ ;
	assign \g220509/_0_  = _w35067_ ;
	assign \g220510/_0_  = _w35074_ ;
	assign \g220511/_0_  = _w35081_ ;
	assign \g220512/_0_  = _w35088_ ;
	assign \g220513/_0_  = _w35095_ ;
	assign \g220514/_0_  = _w35102_ ;
	assign \g220515/_0_  = _w35109_ ;
	assign \g220516/_0_  = _w35116_ ;
	assign \g220517/_0_  = _w35123_ ;
	assign \g220518/_0_  = _w35130_ ;
	assign \g220519/_0_  = _w35137_ ;
	assign \g220520/_0_  = _w35144_ ;
	assign \g220521/_0_  = _w35151_ ;
	assign \g220522/_0_  = _w35158_ ;
	assign \g220523/_0_  = _w35165_ ;
	assign \g220524/_0_  = _w35172_ ;
	assign \g220525/_0_  = _w35179_ ;
	assign \g220526/_0_  = _w35186_ ;
	assign \g220527/_0_  = _w35193_ ;
	assign \g220528/_0_  = _w35200_ ;
	assign \g220529/_0_  = _w35207_ ;
	assign \g220530/_0_  = _w35214_ ;
	assign \g220531/_0_  = _w35221_ ;
	assign \g220532/_0_  = _w35228_ ;
	assign \g220533/_0_  = _w35235_ ;
	assign \g220534/_0_  = _w35239_ ;
	assign \g220535/_0_  = _w35243_ ;
	assign \g220557/_0_  = _w35251_ ;
	assign \g220558/_0_  = _w35254_ ;
	assign \g220559/_0_  = _w35257_ ;
	assign \g220560/_0_  = _w35260_ ;
	assign \g220561/_0_  = _w35263_ ;
	assign \g220562/_0_  = _w35266_ ;
	assign \g220563/_0_  = _w35269_ ;
	assign \g220564/_0_  = _w35272_ ;
	assign \g220565/_0_  = _w35275_ ;
	assign \g220566/_0_  = _w35278_ ;
	assign \g220567/_0_  = _w35281_ ;
	assign \g220568/_0_  = _w35284_ ;
	assign \g220569/_0_  = _w35287_ ;
	assign \g220570/_0_  = _w35290_ ;
	assign \g220571/_0_  = _w35296_ ;
	assign \g220572/_0_  = _w35299_ ;
	assign \g220573/_0_  = _w35302_ ;
	assign \g220574/_0_  = _w35305_ ;
	assign \g220575/_0_  = _w35308_ ;
	assign \g220576/_0_  = _w35311_ ;
	assign \g220577/_0_  = _w35314_ ;
	assign \g220578/_0_  = _w35317_ ;
	assign \g220579/_0_  = _w35320_ ;
	assign \g220580/_0_  = _w35323_ ;
	assign \g220581/_0_  = _w35326_ ;
	assign \g220582/_0_  = _w35329_ ;
	assign \g220583/_0_  = _w35332_ ;
	assign \g220584/_0_  = _w35335_ ;
	assign \g220585/_0_  = _w35338_ ;
	assign \g220586/_0_  = _w35341_ ;
	assign \g220587/_0_  = _w35346_ ;
	assign \g220588/_0_  = _w35349_ ;
	assign \g220589/_0_  = _w35352_ ;
	assign \g220590/_0_  = _w35355_ ;
	assign \g220591/_0_  = _w35358_ ;
	assign \g220592/_0_  = _w35361_ ;
	assign \g220593/_0_  = _w35364_ ;
	assign \g220594/_0_  = _w35367_ ;
	assign \g220595/_0_  = _w35370_ ;
	assign \g220596/_0_  = _w35373_ ;
	assign \g220597/_0_  = _w35376_ ;
	assign \g220598/_0_  = _w35379_ ;
	assign \g220599/_0_  = _w35382_ ;
	assign \g220600/_0_  = _w35385_ ;
	assign \g220601/_0_  = _w35388_ ;
	assign \g220602/_0_  = _w35391_ ;
	assign \g220603/_0_  = _w35394_ ;
	assign \g220604/_0_  = _w35398_ ;
	assign \g220605/_0_  = _w35401_ ;
	assign \g220606/_0_  = _w35404_ ;
	assign \g220607/_0_  = _w35407_ ;
	assign \g220608/_0_  = _w35410_ ;
	assign \g220609/_0_  = _w35413_ ;
	assign \g220610/_0_  = _w35416_ ;
	assign \g220611/_0_  = _w35419_ ;
	assign \g220612/_0_  = _w35422_ ;
	assign \g220613/_0_  = _w35425_ ;
	assign \g220614/_0_  = _w35428_ ;
	assign \g220615/_0_  = _w35431_ ;
	assign \g220616/_0_  = _w35434_ ;
	assign \g220617/_0_  = _w35437_ ;
	assign \g220618/_0_  = _w35440_ ;
	assign \g220619/_0_  = _w35443_ ;
	assign \g220620/_0_  = _w35449_ ;
	assign \g220621/_0_  = _w35452_ ;
	assign \g220622/_0_  = _w35455_ ;
	assign \g220623/_0_  = _w35458_ ;
	assign \g220624/_0_  = _w35461_ ;
	assign \g220625/_0_  = _w35464_ ;
	assign \g220626/_0_  = _w35467_ ;
	assign \g220627/_0_  = _w35470_ ;
	assign \g220628/_0_  = _w35473_ ;
	assign \g220629/_0_  = _w35476_ ;
	assign \g220630/_0_  = _w35479_ ;
	assign \g220631/_0_  = _w35482_ ;
	assign \g220632/_0_  = _w35485_ ;
	assign \g220633/_0_  = _w35488_ ;
	assign \g220634/_0_  = _w35491_ ;
	assign \g220635/_0_  = _w35494_ ;
	assign \g220636/_0_  = _w35497_ ;
	assign \g220637/_0_  = _w35500_ ;
	assign \g220638/_0_  = _w35503_ ;
	assign \g220639/_0_  = _w35506_ ;
	assign \g220640/_0_  = _w35509_ ;
	assign \g220641/_0_  = _w35512_ ;
	assign \g220642/_0_  = _w35515_ ;
	assign \g220643/_0_  = _w35522_ ;
	assign \g220644/_0_  = _w35525_ ;
	assign \g220645/_0_  = _w35528_ ;
	assign \g220646/_0_  = _w35531_ ;
	assign \g220647/_0_  = _w35534_ ;
	assign \g220648/_0_  = _w35537_ ;
	assign \g220649/_0_  = _w35540_ ;
	assign \g220650/_0_  = _w35543_ ;
	assign \g220651/_0_  = _w35546_ ;
	assign \g220652/_0_  = _w35549_ ;
	assign \g220653/_0_  = _w35552_ ;
	assign \g220654/_0_  = _w35555_ ;
	assign \g220655/_0_  = _w35558_ ;
	assign \g220656/_0_  = _w35561_ ;
	assign \g220657/_0_  = _w35564_ ;
	assign \g220658/_0_  = _w35567_ ;
	assign \g220659/_0_  = _w35570_ ;
	assign \g220660/_0_  = _w35573_ ;
	assign \g220661/_0_  = _w35576_ ;
	assign \g220662/_0_  = _w35579_ ;
	assign \g220663/_0_  = _w35582_ ;
	assign \g220664/_0_  = _w35585_ ;
	assign \g220665/_0_  = _w35588_ ;
	assign \g220666/_0_  = _w35591_ ;
	assign \g220674/_0_  = _w35595_ ;
	assign \g220679/u3_syn_7  = _w35598_ ;
	assign \g220711/u3_syn_4  = _w35600_ ;
	assign \g220726/u3_syn_4  = _w35601_ ;
	assign \g220739/u3_syn_4  = _w35602_ ;
	assign \g220751/u3_syn_4  = _w35603_ ;
	assign \g220759/u3_syn_4  = _w35605_ ;
	assign \g220773/u3_syn_4  = _w35606_ ;
	assign \g220782/u3_syn_4  = _w35607_ ;
	assign \g220805/u3_syn_4  = _w35608_ ;
	assign \g220828/u3_syn_4  = _w35610_ ;
	assign \g220921/_0_  = _w34306_ ;
	assign \g220930/u3_syn_4  = _w35612_ ;
	assign \g220949/_3_  = _w35616_ ;
	assign \g220994/_3_  = _w11512_ ;
	assign \g221207/_0_  = _w35639_ ;
	assign \g221213/_0_  = _w11380_ ;
	assign \g221223/_0_  = _w35647_ ;
	assign \g221224/_0_  = _w35654_ ;
	assign \g221225/_0_  = _w35659_ ;
	assign \g221226/_0_  = _w35665_ ;
	assign \g221231/_0_  = _w35671_ ;
	assign \g221232/_0_  = _w35675_ ;
	assign \g221234/_0_  = _w35678_ ;
	assign \g221235/_0_  = _w35681_ ;
	assign \g221246/_2_  = _w11382_ ;
	assign \g221249/_2_  = _w11379_ ;
	assign \g221265/_0_  = _w35683_ ;
	assign \g221287/_0_  = _w35685_ ;
	assign \g221325/_0_  = _w35688_ ;
	assign \g221326/_0_  = _w35695_ ;
	assign \g221447/_0_  = _w35698_ ;
	assign \g221449/_0_  = _w35701_ ;
	assign \g221452/_0_  = _w35702_ ;
	assign \g221469/_0_  = _w35703_ ;
	assign \g221473/_0_  = _w35710_ ;
	assign \g221503/_0_  = _w35713_ ;
	assign \g221510/_0_  = _w35720_ ;
	assign \g221512/_0_  = _w35728_ ;
	assign \g221516/_0_  = _w35733_ ;
	assign \g221517/_0_  = _w35738_ ;
	assign \g221524/_0_  = _w35745_ ;
	assign \g221530/_0_  = _w35750_ ;
	assign \g221592/_0_  = _w35753_ ;
	assign \g221593/_0_  = _w35756_ ;
	assign \g221634/u3_syn_4  = _w35248_ ;
	assign \g221669/u3_syn_4  = _w35293_ ;
	assign \g221789/u3_syn_4  = _w35343_ ;
	assign \g221813/u3_syn_4  = _w35395_ ;
	assign \g221829/u3_syn_4  = _w35446_ ;
	assign \g221861/u3_syn_4  = _w35519_ ;
	assign \g221876/_0_  = _w35759_ ;
	assign \g221935/_0_  = _w35762_ ;
	assign \g221944/_3_  = _w11361_ ;
	assign \g230200/_0_  = _w35765_ ;
	assign \g230201/_0_  = _w34545_ ;
	assign \g230205/_0_  = _w35768_ ;
	assign \g230295/_0_  = _w35772_ ;
	assign \g230297/_0_  = _w35778_ ;
	assign \g230298/_0_  = _w35784_ ;
	assign \g230300/_0_  = _w35790_ ;
	assign \g230302/_0_  = _w35799_ ;
	assign \g230303/_0_  = _w35807_ ;
	assign \g230343/_0_  = _w35811_ ;
	assign \g230368/_0_  = _w35813_ ;
	assign \g230511/_0_  = _w35816_ ;
	assign \g230531/_0_  = _w35818_ ;
	assign \g230635/_2_  = _w34527_ ;
	assign \g230661/_0_  = _w35821_ ;
	assign \g230715/_1__syn_2  = _w35822_ ;
	assign \g230731/_0_  = _w35842_ ;
	assign \g230766/_0_  = _w35844_ ;
	assign \g230784/_0_  = _w35848_ ;
	assign \g230785/_0_  = _w35852_ ;
	assign \g230786/_0_  = _w35856_ ;
	assign \g230787/_0_  = _w35860_ ;
	assign \g230797/_0_  = _w35863_ ;
	assign \g230798/_0_  = _w35865_ ;
	assign \g230803/_0_  = _w35867_ ;
	assign \g230804/_00_  = _w35870_ ;
	assign \g230805/_00_  = _w35873_ ;
	assign \g230806/_00_  = _w35876_ ;
	assign \g230807/_00_  = _w35879_ ;
	assign \g230808/_00_  = _w35882_ ;
	assign \g230809/_00_  = _w35885_ ;
	assign \g230815/_0_  = _w35889_ ;
	assign \g230816/_2_  = _w35891_ ;
	assign \g230817/_2_  = _w35893_ ;
	assign \g230829/_0_  = _w35905_ ;
	assign \g230834/_0_  = _w35910_ ;
	assign \g230835/_0_  = _w35914_ ;
	assign \g230836/_0_  = _w35917_ ;
	assign \g230837/_0_  = _w35925_ ;
	assign \g230844/_0_  = _w35928_ ;
	assign \g230863/_3_  = _w35935_ ;
	assign \g230864/_3_  = _w35940_ ;
	assign \g230870/_0_  = _w35945_ ;
	assign \g230988/_3_  = _w35950_ ;
	assign \g231010/_3_  = _w35953_ ;
	assign \g231016/_3_  = _w35956_ ;
	assign \g231042/_3_  = _w35959_ ;
	assign \g231471/_0_  = _w35962_ ;
	assign \g231472/_0_  = _w35965_ ;
	assign \g231476/_3_  = _w11465_ ;
	assign \g231480/_3_  = _w11531_ ;
	assign \g231484/_3_  = _w11506_ ;
	assign \g231504/_0_  = _w35969_ ;
	assign \g231532/_0_  = _w31401_ ;
	assign \g231542/_0_  = _w35972_ ;
	assign \g231560/_1_  = _w35975_ ;
	assign \g231578/_1_  = _w35978_ ;
	assign \g231580/_0_  = _w35981_ ;
	assign \g231590/_1__syn_2  = _w34106_ ;
	assign \g231615/_0_  = _w35984_ ;
	assign \g231623/_1_  = _w35985_ ;
	assign \g231634/_2_  = _w35986_ ;
	assign \g231635/_0_  = _w35988_ ;
	assign \g231638/_2_  = _w35989_ ;
	assign \g231640/_0_  = _w35992_ ;
	assign \g231653/_2_  = _w35993_ ;
	assign \g231787/_0_  = _w35995_ ;
	assign \g231931/_0_  = _w35998_ ;
	assign \g231939/_3_  = _w36000_ ;
	assign \g231940/_0_  = _w36003_ ;
	assign \g231951/_0_  = _w36008_ ;
	assign \g231955/_0_  = _w36009_ ;
	assign \g231956/_0_  = _w36015_ ;
	assign \g231959/_2_  = _w36016_ ;
	assign \g231960/_0_  = _w36017_ ;
	assign \g231964/_0_  = _w36021_ ;
	assign \g231965/_0_  = _w36026_ ;
	assign \g231975/_0_  = _w36031_ ;
	assign \g231986/_1_  = _w36033_ ;
	assign \g231987/_1_  = _w36034_ ;
	assign \g231989/_1_  = _w36036_ ;
	assign \g231990/_1_  = _w36037_ ;
	assign \g231991/_0_  = _w36054_ ;
	assign \g231992/_0_  = _w36070_ ;
	assign \g231995/_0_  = _w36076_ ;
	assign \g231998/_0_  = _w36078_ ;
	assign \g231999/_0_  = _w36082_ ;
	assign \g232002/_3_  = _w36097_ ;
	assign \g232035/u3_syn_4  = _w36109_ ;
	assign \g232038/u3_syn_4  = _w36116_ ;
	assign \g232046/u3_syn_4  = _w36121_ ;
	assign \g232054/u3_syn_4  = _w36126_ ;
	assign \g232062/u3_syn_4  = _w36129_ ;
	assign \g232070/u3_syn_4  = _w36131_ ;
	assign \g232078/u3_syn_4  = _w36139_ ;
	assign \g232079/u3_syn_4  = _w36143_ ;
	assign \g232087/u3_syn_4  = _w36146_ ;
	assign \g232096/u3_syn_4  = _w36148_ ;
	assign \g232104/u3_syn_4  = _w36151_ ;
	assign \g232112/u3_syn_4  = _w36153_ ;
	assign \g232120/u3_syn_4  = _w36160_ ;
	assign \g232128/u3_syn_4  = _w36164_ ;
	assign \g232136/u3_syn_4  = _w36168_ ;
	assign \g232144/u3_syn_4  = _w36172_ ;
	assign \g232152/u3_syn_4  = _w36175_ ;
	assign \g232161/u3_syn_4  = _w36178_ ;
	assign \g232169/u3_syn_4  = _w36180_ ;
	assign \g232177/u3_syn_4  = _w36183_ ;
	assign \g232185/u3_syn_4  = _w36184_ ;
	assign \g232186/u3_syn_4  = _w36188_ ;
	assign \g232194/u3_syn_4  = _w36191_ ;
	assign \g232202/u3_syn_4  = _w36193_ ;
	assign \g232210/u3_syn_4  = _w36196_ ;
	assign \g232218/u3_syn_4  = _w36199_ ;
	assign \g232226/u3_syn_4  = _w36201_ ;
	assign \g232234/u3_syn_4  = _w36204_ ;
	assign \g232242/u3_syn_4  = _w36206_ ;
	assign \g232251/u3_syn_4  = _w36209_ ;
	assign \g232259/u3_syn_4  = _w36211_ ;
	assign \g232267/u3_syn_4  = _w36214_ ;
	assign \g232275/u3_syn_4  = _w36216_ ;
	assign \g232283/u3_syn_4  = _w36218_ ;
	assign \g232291/u3_syn_4  = _w36220_ ;
	assign \g232299/u3_syn_4  = _w36222_ ;
	assign \g232307/u3_syn_4  = _w36224_ ;
	assign \g232315/u3_syn_4  = _w36226_ ;
	assign \g232324/u3_syn_4  = _w36228_ ;
	assign \g232332/u3_syn_4  = _w36230_ ;
	assign \g232341/u3_syn_4  = _w36232_ ;
	assign \g232349/u3_syn_4  = _w36234_ ;
	assign \g232357/u3_syn_4  = _w36236_ ;
	assign \g232366/u3_syn_4  = _w36238_ ;
	assign \g232374/u3_syn_4  = _w36240_ ;
	assign \g232382/u3_syn_4  = _w36242_ ;
	assign \g232390/u3_syn_4  = _w36244_ ;
	assign \g232398/u3_syn_4  = _w36246_ ;
	assign \g232406/u3_syn_4  = _w36248_ ;
	assign \g232414/u3_syn_4  = _w36250_ ;
	assign \g232422/u3_syn_4  = _w36252_ ;
	assign \g232427/u3_syn_4  = _w36253_ ;
	assign \g232431/u3_syn_4  = _w36255_ ;
	assign \g232439/u3_syn_4  = _w36257_ ;
	assign \g232444/u3_syn_4  = _w36258_ ;
	assign \g232452/u3_syn_4  = _w36260_ ;
	assign \g232461/u3_syn_4  = _w36261_ ;
	assign \g232471/u3_syn_4  = _w36263_ ;
	assign \g232479/u3_syn_4  = _w36265_ ;
	assign \g232487/u3_syn_4  = _w36266_ ;
	assign \g232495/u3_syn_4  = _w36267_ ;
	assign \g232503/u3_syn_4  = _w36269_ ;
	assign \g232506/u3_syn_4  = _w36270_ ;
	assign \g232514/u3_syn_4  = _w36272_ ;
	assign \g232527/u3_syn_4  = _w36273_ ;
	assign \g232530/u3_syn_4  = _w36276_ ;
	assign \g232536/u3_syn_4  = _w36277_ ;
	assign \g232544/u3_syn_4  = _w36280_ ;
	assign \g232551/u3_syn_4  = _w36281_ ;
	assign \g232557/u3_syn_4  = _w36283_ ;
	assign \g232568/u3_syn_4  = _w36285_ ;
	assign \g232576/u3_syn_4  = _w36287_ ;
	assign \g232585/u3_syn_4  = _w36288_ ;
	assign \g232593/u3_syn_4  = _w36289_ ;
	assign \g232597/u3_syn_4  = _w36291_ ;
	assign \g232609/u3_syn_4  = _w36293_ ;
	assign \g232617/u3_syn_4  = _w36295_ ;
	assign \g232625/u3_syn_4  = _w36297_ ;
	assign \g232633/u3_syn_4  = _w36299_ ;
	assign \g232641/u3_syn_4  = _w36301_ ;
	assign \g232649/u3_syn_4  = _w36303_ ;
	assign \g232657/u3_syn_4  = _w36305_ ;
	assign \g232665/u3_syn_4  = _w36307_ ;
	assign \g232673/u3_syn_4  = _w36309_ ;
	assign \g232681/u3_syn_4  = _w36311_ ;
	assign \g232689/u3_syn_4  = _w36312_ ;
	assign \g232697/u3_syn_4  = _w36313_ ;
	assign \g232705/u3_syn_4  = _w36315_ ;
	assign \g232713/u3_syn_4  = _w36316_ ;
	assign \g232717/u3_syn_4  = _w36318_ ;
	assign \g232729/u3_syn_4  = _w36320_ ;
	assign \g232737/u3_syn_4  = _w36321_ ;
	assign \g232745/u3_syn_4  = _w36323_ ;
	assign \g232749/u3_syn_4  = _w36324_ ;
	assign \g232761/u3_syn_4  = _w36325_ ;
	assign \g232768/u3_syn_4  = _w36327_ ;
	assign \g232777/u3_syn_4  = _w36329_ ;
	assign \g232785/u3_syn_4  = _w36331_ ;
	assign \g232793/u3_syn_4  = _w36333_ ;
	assign \g232801/u3_syn_4  = _w36335_ ;
	assign \g232809/u3_syn_4  = _w36337_ ;
	assign \g232815/u3_syn_4  = _w36338_ ;
	assign \g232823/u3_syn_4  = _w36340_ ;
	assign \g232833/u3_syn_4  = _w36341_ ;
	assign \g232841/u3_syn_4  = _w36343_ ;
	assign \g232846/u3_syn_4  = _w36344_ ;
	assign \g232851/u3_syn_4  = _w36346_ ;
	assign \g232865/u3_syn_4  = _w36347_ ;
	assign \g232873/u3_syn_4  = _w36348_ ;
	assign \g232881/u3_syn_4  = _w36349_ ;
	assign \g232882/u3_syn_4  = _w36352_ ;
	assign \g232895/u3_syn_4  = _w36353_ ;
	assign \g232904/u3_syn_4  = _w36354_ ;
	assign \g232913/u3_syn_4  = _w36355_ ;
	assign \g232921/u3_syn_4  = _w36356_ ;
	assign \g232928/u3_syn_4  = _w36357_ ;
	assign \g232934/u3_syn_4  = _w36358_ ;
	assign \g232945/u3_syn_4  = _w36359_ ;
	assign \g232953/u3_syn_4  = _w36360_ ;
	assign \g232954/u3_syn_4  = _w36361_ ;
	assign \g232969/u3_syn_4  = _w36362_ ;
	assign \g232977/u3_syn_4  = _w36363_ ;
	assign \g232981/u3_syn_4  = _w36364_ ;
	assign \g232993/u3_syn_4  = _w36365_ ;
	assign \g232995/u3_syn_4  = _w36366_ ;
	assign \g233009/u3_syn_4  = _w36367_ ;
	assign \g233017/u3_syn_4  = _w36368_ ;
	assign \g233025/u3_syn_4  = _w36369_ ;
	assign \g233033/u3_syn_4  = _w36370_ ;
	assign \g233041/u3_syn_4  = _w36371_ ;
	assign \g233047/u3_syn_4  = _w36372_ ;
	assign \g233057/u3_syn_4  = _w36373_ ;
	assign \g233065/u3_syn_4  = _w36374_ ;
	assign \g233073/u3_syn_4  = _w36375_ ;
	assign \g233081/u3_syn_4  = _w36376_ ;
	assign \g233087/u3_syn_4  = _w36377_ ;
	assign \g233097/u3_syn_4  = _w36378_ ;
	assign \g233105/u3_syn_4  = _w36379_ ;
	assign \g233113/u3_syn_4  = _w36380_ ;
	assign \g233121/u3_syn_4  = _w36381_ ;
	assign \g233128/u3_syn_4  = _w36382_ ;
	assign \g233134/u3_syn_4  = _w36383_ ;
	assign \g233144/u3_syn_4  = _w36384_ ;
	assign \g233153/u3_syn_4  = _w36385_ ;
	assign \g233161/u3_syn_4  = _w36386_ ;
	assign \g233169/u3_syn_4  = _w36387_ ;
	assign \g233177/u3_syn_4  = _w36388_ ;
	assign \g233185/u3_syn_4  = _w36389_ ;
	assign \g233193/u3_syn_4  = _w36390_ ;
	assign \g233201/u3_syn_4  = _w36391_ ;
	assign \g233209/u3_syn_4  = _w36392_ ;
	assign \g233217/u3_syn_4  = _w36393_ ;
	assign \g233219/u3_syn_4  = _w36394_ ;
	assign \g233229/u3_syn_4  = _w36395_ ;
	assign \g233241/u3_syn_4  = _w36396_ ;
	assign \g233249/u3_syn_4  = _w36397_ ;
	assign \g233257/u3_syn_4  = _w36398_ ;
	assign \g233265/u3_syn_4  = _w36399_ ;
	assign \g233273/u3_syn_4  = _w36400_ ;
	assign \g233281/u3_syn_4  = _w36401_ ;
	assign \g233289/u3_syn_4  = _w36402_ ;
	assign \g233297/u3_syn_4  = _w36403_ ;
	assign \g233305/u3_syn_4  = _w36404_ ;
	assign \g233313/u3_syn_4  = _w36405_ ;
	assign \g233321/u3_syn_4  = _w36406_ ;
	assign \g233329/u3_syn_4  = _w36407_ ;
	assign \g233337/u3_syn_4  = _w36408_ ;
	assign \g233345/u3_syn_4  = _w36409_ ;
	assign \g233353/u3_syn_4  = _w36410_ ;
	assign \g233361/u3_syn_4  = _w36411_ ;
	assign \g233369/u3_syn_4  = _w36412_ ;
	assign \g233377/u3_syn_4  = _w36413_ ;
	assign \g233382/u3_syn_4  = _w36414_ ;
	assign \g233392/u3_syn_4  = _w36415_ ;
	assign \g233394/u3_syn_4  = _w36416_ ;
	assign \g233409/u3_syn_4  = _w36417_ ;
	assign \g233417/u3_syn_4  = _w36418_ ;
	assign \g233425/u3_syn_4  = _w36419_ ;
	assign \g233433/u3_syn_4  = _w36420_ ;
	assign \g233441/u3_syn_4  = _w36421_ ;
	assign \g233449/u3_syn_4  = _w36422_ ;
	assign \g233453/u3_syn_4  = _w36423_ ;
	assign \g233465/u3_syn_4  = _w36424_ ;
	assign \g233473/u3_syn_4  = _w36425_ ;
	assign \g233481/u3_syn_4  = _w36426_ ;
	assign \g233489/u3_syn_4  = _w36427_ ;
	assign \g233497/u3_syn_4  = _w36428_ ;
	assign \g233505/u3_syn_4  = _w36429_ ;
	assign \g233513/u3_syn_4  = _w36430_ ;
	assign \g233516/u3_syn_4  = _w36431_ ;
	assign \g233529/u3_syn_4  = _w36432_ ;
	assign \g233531/u3_syn_4  = _w36433_ ;
	assign \g233546/u3_syn_4  = _w36434_ ;
	assign \g233554/u3_syn_4  = _w36435_ ;
	assign \g233562/u3_syn_4  = _w36436_ ;
	assign \g233570/u3_syn_4  = _w36437_ ;
	assign \g233578/u3_syn_4  = _w36438_ ;
	assign \g233586/u3_syn_4  = _w36439_ ;
	assign \g233594/u3_syn_4  = _w36440_ ;
	assign \g233602/u3_syn_4  = _w36441_ ;
	assign \g233603/u3_syn_4  = _w36442_ ;
	assign \g233618/u3_syn_4  = _w36443_ ;
	assign \g233626/u3_syn_4  = _w36444_ ;
	assign \g233634/u3_syn_4  = _w36445_ ;
	assign \g233642/u3_syn_4  = _w36446_ ;
	assign \g233650/u3_syn_4  = _w36447_ ;
	assign \g233658/u3_syn_4  = _w36448_ ;
	assign \g233666/u3_syn_4  = _w36449_ ;
	assign \g233674/u3_syn_4  = _w36450_ ;
	assign \g233682/u3_syn_4  = _w36451_ ;
	assign \g233690/u3_syn_4  = _w36452_ ;
	assign \g233698/u3_syn_4  = _w36453_ ;
	assign \g233706/u3_syn_4  = _w36454_ ;
	assign \g233714/u3_syn_4  = _w36455_ ;
	assign \g233722/u3_syn_4  = _w36456_ ;
	assign \g233730/u3_syn_4  = _w36457_ ;
	assign \g233738/u3_syn_4  = _w36458_ ;
	assign \g233746/u3_syn_4  = _w36459_ ;
	assign \g233754/u3_syn_4  = _w36460_ ;
	assign \g233762/u3_syn_4  = _w36461_ ;
	assign \g233770/u3_syn_4  = _w36462_ ;
	assign \g233778/u3_syn_4  = _w36463_ ;
	assign \g233783/u3_syn_4  = _w36464_ ;
	assign \g233794/u3_syn_4  = _w36465_ ;
	assign \g233802/u3_syn_4  = _w36466_ ;
	assign \g233806/u3_syn_4  = _w36467_ ;
	assign \g233818/u3_syn_4  = _w36468_ ;
	assign \g233826/u3_syn_4  = _w36469_ ;
	assign \g233828/u3_syn_4  = _w36470_ ;
	assign \g233838/u3_syn_4  = _w36471_ ;
	assign \g233850/u3_syn_4  = _w36472_ ;
	assign \g233858/u3_syn_4  = _w36473_ ;
	assign \g233860/u3_syn_4  = _w36474_ ;
	assign \g233870/u3_syn_4  = _w36475_ ;
	assign \g233881/u3_syn_4  = _w36476_ ;
	assign \g233890/u3_syn_4  = _w36477_ ;
	assign \g233899/u3_syn_4  = _w36478_ ;
	assign \g233908/u3_syn_4  = _w36479_ ;
	assign \g233917/u3_syn_4  = _w36480_ ;
	assign \g233919/u3_syn_4  = _w36481_ ;
	assign \g233927/u3_syn_4  = _w36482_ ;
	assign \g233935/u3_syn_4  = _w36483_ ;
	assign \g233943/u3_syn_4  = _w36484_ ;
	assign \g233945/u3_syn_4  = _w36485_ ;
	assign \g233953/u3_syn_4  = _w36486_ ;
	assign \g233961/u3_syn_4  = _w36487_ ;
	assign \g233969/u3_syn_4  = _w36488_ ;
	assign \g233977/u3_syn_4  = _w36489_ ;
	assign \g233985/u3_syn_4  = _w36490_ ;
	assign \g233993/u3_syn_4  = _w36491_ ;
	assign \g234001/u3_syn_4  = _w36492_ ;
	assign \g234008/u3_syn_4  = _w36493_ ;
	assign \g234009/u3_syn_4  = _w36494_ ;
	assign \g234024/u3_syn_4  = _w36495_ ;
	assign \g234032/u3_syn_4  = _w36496_ ;
	assign \g234038/u3_syn_4  = _w36497_ ;
	assign \g234056/u3_syn_4  = _w36498_ ;
	assign \g234063/u3_syn_4  = _w36499_ ;
	assign \g234071/u3_syn_4  = _w36500_ ;
	assign \g234079/u3_syn_4  = _w36501_ ;
	assign \g234098/u3_syn_4  = _w36502_ ;
	assign \g234106/u3_syn_4  = _w36503_ ;
	assign \g234114/u3_syn_4  = _w36504_ ;
	assign \g234122/u3_syn_4  = _w36505_ ;
	assign \g234130/u3_syn_4  = _w36506_ ;
	assign \g234138/u3_syn_4  = _w36507_ ;
	assign \g234145/u3_syn_4  = _w36508_ ;
	assign \g234156/u3_syn_4  = _w36509_ ;
	assign \g234162/u3_syn_4  = _w36510_ ;
	assign \g234171/u3_syn_4  = _w36511_ ;
	assign \g234183/u3_syn_4  = _w36512_ ;
	assign \g234248/u3_syn_4  = _w36513_ ;
	assign \g234265/u3_syn_4  = _w36514_ ;
	assign \g234273/u3_syn_4  = _w36515_ ;
	assign \g234281/u3_syn_4  = _w36516_ ;
	assign \g234289/u3_syn_4  = _w36517_ ;
	assign \g234297/u3_syn_4  = _w36518_ ;
	assign \g234306/u3_syn_4  = _w36519_ ;
	assign \g234314/u3_syn_4  = _w36520_ ;
	assign \g234322/u3_syn_4  = _w36521_ ;
	assign \g234331/u3_syn_4  = _w36522_ ;
	assign \g234339/u3_syn_4  = _w36523_ ;
	assign \g234347/u3_syn_4  = _w36524_ ;
	assign \g234355/u3_syn_4  = _w36525_ ;
	assign \g234363/u3_syn_4  = _w36526_ ;
	assign \g234371/u3_syn_4  = _w36527_ ;
	assign \g234379/u3_syn_4  = _w36528_ ;
	assign \g234387/u3_syn_4  = _w36529_ ;
	assign \g234395/u3_syn_4  = _w36530_ ;
	assign \g234403/u3_syn_4  = _w36531_ ;
	assign \g234411/u3_syn_4  = _w36532_ ;
	assign \g234419/u3_syn_4  = _w36533_ ;
	assign \g234427/u3_syn_4  = _w36534_ ;
	assign \g234435/u3_syn_4  = _w36535_ ;
	assign \g234443/u3_syn_4  = _w36536_ ;
	assign \g234451/u3_syn_4  = _w36537_ ;
	assign \g234459/u3_syn_4  = _w36538_ ;
	assign \g234467/u3_syn_4  = _w36539_ ;
	assign \g234475/u3_syn_4  = _w36540_ ;
	assign \g234483/u3_syn_4  = _w36541_ ;
	assign \g234491/u3_syn_4  = _w36542_ ;
	assign \g234499/u3_syn_4  = _w36543_ ;
	assign \g234507/u3_syn_4  = _w36544_ ;
	assign \g234515/u3_syn_4  = _w36545_ ;
	assign \g234523/u3_syn_4  = _w36546_ ;
	assign \g234531/u3_syn_4  = _w36547_ ;
	assign \g234539/u3_syn_4  = _w36548_ ;
	assign \g234547/u3_syn_4  = _w36549_ ;
	assign \g234555/u3_syn_4  = _w36550_ ;
	assign \g234563/u3_syn_4  = _w36551_ ;
	assign \g234571/u3_syn_4  = _w36552_ ;
	assign \g234579/u3_syn_4  = _w36553_ ;
	assign \g234587/u3_syn_4  = _w36554_ ;
	assign \g234595/u3_syn_4  = _w36555_ ;
	assign \g234604/u3_syn_4  = _w36556_ ;
	assign \g234612/u3_syn_4  = _w36557_ ;
	assign \g234620/u3_syn_4  = _w36558_ ;
	assign \g234628/u3_syn_4  = _w36559_ ;
	assign \g234636/u3_syn_4  = _w36560_ ;
	assign \g234644/u3_syn_4  = _w36561_ ;
	assign \g234652/u3_syn_4  = _w36562_ ;
	assign \g234660/u3_syn_4  = _w36563_ ;
	assign \g234668/u3_syn_4  = _w36564_ ;
	assign \g234676/u3_syn_4  = _w36565_ ;
	assign \g234684/u3_syn_4  = _w36566_ ;
	assign \g234692/u3_syn_4  = _w36567_ ;
	assign \g234700/u3_syn_4  = _w36568_ ;
	assign \g234708/u3_syn_4  = _w36569_ ;
	assign \g234716/u3_syn_4  = _w36570_ ;
	assign \g234725/u3_syn_4  = _w36571_ ;
	assign \g234733/u3_syn_4  = _w36572_ ;
	assign \g234741/u3_syn_4  = _w36573_ ;
	assign \g234749/u3_syn_4  = _w36574_ ;
	assign \g234757/u3_syn_4  = _w36575_ ;
	assign \g234765/u3_syn_4  = _w36576_ ;
	assign \g234773/u3_syn_4  = _w36577_ ;
	assign \g234781/u3_syn_4  = _w36578_ ;
	assign \g234789/u3_syn_4  = _w36579_ ;
	assign \g234798/u3_syn_4  = _w36580_ ;
	assign \g234806/u3_syn_4  = _w36581_ ;
	assign \g234814/u3_syn_4  = _w36582_ ;
	assign \g234822/u3_syn_4  = _w36583_ ;
	assign \g234830/u3_syn_4  = _w36584_ ;
	assign \g234838/u3_syn_4  = _w36585_ ;
	assign \g235911/u3_syn_4  = _w36587_ ;
	assign \g235912/u3_syn_4  = _w36589_ ;
	assign \g235920/u3_syn_4  = _w36591_ ;
	assign \g235928/u3_syn_4  = _w36593_ ;
	assign \g235936/u3_syn_4  = _w36595_ ;
	assign \g235944/u3_syn_4  = _w36597_ ;
	assign \g235952/u3_syn_4  = _w36599_ ;
	assign \g235960/u3_syn_4  = _w36601_ ;
	assign \g235968/u3_syn_4  = _w36603_ ;
	assign \g235976/u3_syn_4  = _w36605_ ;
	assign \g235984/u3_syn_4  = _w36607_ ;
	assign \g235992/u3_syn_4  = _w36609_ ;
	assign \g236000/u3_syn_4  = _w36610_ ;
	assign \g236008/u3_syn_4  = _w36612_ ;
	assign \g236016/u3_syn_4  = _w36614_ ;
	assign \g236021/u3_syn_4  = _w36616_ ;
	assign \g236025/u3_syn_4  = _w36618_ ;
	assign \g236033/u3_syn_4  = _w36620_ ;
	assign \g236041/u3_syn_4  = _w36622_ ;
	assign \g236049/u3_syn_4  = _w36624_ ;
	assign \g236057/u3_syn_4  = _w36626_ ;
	assign \g236065/u3_syn_4  = _w36628_ ;
	assign \g236073/u3_syn_4  = _w36630_ ;
	assign \g236081/u3_syn_4  = _w36632_ ;
	assign \g236089/u3_syn_4  = _w36634_ ;
	assign \g236097/u3_syn_4  = _w36636_ ;
	assign \g236105/u3_syn_4  = _w36638_ ;
	assign \g236113/u3_syn_4  = _w36640_ ;
	assign \g236121/u3_syn_4  = _w36642_ ;
	assign \g236129/u3_syn_4  = _w36644_ ;
	assign \g236137/u3_syn_4  = _w36646_ ;
	assign \g236145/u3_syn_4  = _w36648_ ;
	assign \g236153/u3_syn_4  = _w36650_ ;
	assign \g236161/u3_syn_4  = _w36652_ ;
	assign \g236169/u3_syn_4  = _w36654_ ;
	assign \g236177/u3_syn_4  = _w36656_ ;
	assign \g236185/u3_syn_4  = _w36658_ ;
	assign \g236193/u3_syn_4  = _w36660_ ;
	assign \g236196/u3_syn_4  = _w36661_ ;
	assign \g236198/u3_syn_4  = _w36662_ ;
	assign \g236203/u3_syn_4  = _w36664_ ;
	assign \g236211/u3_syn_4  = _w36666_ ;
	assign \g236219/u3_syn_4  = _w36667_ ;
	assign \g236220/u3_syn_4  = _w36669_ ;
	assign \g236229/u3_syn_4  = _w36671_ ;
	assign \g236232/u3_syn_4  = _w36672_ ;
	assign \g236238/u3_syn_4  = _w36674_ ;
	assign \g236246/u3_syn_4  = _w36676_ ;
	assign \g236255/u3_syn_4  = _w36678_ ;
	assign \g236263/u3_syn_4  = _w36680_ ;
	assign \g236271/u3_syn_4  = _w36682_ ;
	assign \g236275/u3_syn_4  = _w36683_ ;
	assign \g236280/u3_syn_4  = _w36685_ ;
	assign \g236288/u3_syn_4  = _w36687_ ;
	assign \g236296/u3_syn_4  = _w36689_ ;
	assign \g236304/u3_syn_4  = _w36690_ ;
	assign \g236305/u3_syn_4  = _w36691_ ;
	assign \g236306/u3_syn_4  = _w36693_ ;
	assign \g236315/u3_syn_4  = _w36695_ ;
	assign \g236323/u3_syn_4  = _w36697_ ;
	assign \g236331/u3_syn_4  = _w36699_ ;
	assign \g236334/u3_syn_4  = _w36700_ ;
	assign \g236340/u3_syn_4  = _w36702_ ;
	assign \g236348/u3_syn_4  = _w36704_ ;
	assign \g236357/u3_syn_4  = _w36705_ ;
	assign \g236359/u3_syn_4  = _w36707_ ;
	assign \g236367/u3_syn_4  = _w36709_ ;
	assign \g236374/u3_syn_4  = _w36710_ ;
	assign \g236376/u3_syn_4  = _w36712_ ;
	assign \g236377/u3_syn_4  = _w36714_ ;
	assign \g236385/u3_syn_4  = _w36716_ ;
	assign \g236393/u3_syn_4  = _w36718_ ;
	assign \g236402/u3_syn_4  = _w36720_ ;
	assign \g236410/u3_syn_4  = _w36722_ ;
	assign \g236419/u3_syn_4  = _w36724_ ;
	assign \g236427/u3_syn_4  = _w36726_ ;
	assign \g236433/u3_syn_4  = _w36727_ ;
	assign \g236436/u3_syn_4  = _w36729_ ;
	assign \g236444/u3_syn_4  = _w36731_ ;
	assign \g236452/u3_syn_4  = _w36733_ ;
	assign \g236460/u3_syn_4  = _w36735_ ;
	assign \g236468/u3_syn_4  = _w36737_ ;
	assign \g236476/u3_syn_4  = _w36739_ ;
	assign \g236484/u3_syn_4  = _w36741_ ;
	assign \g236492/u3_syn_4  = _w36743_ ;
	assign \g236500/u3_syn_4  = _w36745_ ;
	assign \g236508/u3_syn_4  = _w36747_ ;
	assign \g236516/u3_syn_4  = _w36749_ ;
	assign \g236518/u3_syn_4  = _w36750_ ;
	assign \g236525/u3_syn_4  = _w36752_ ;
	assign \g236533/u3_syn_4  = _w36754_ ;
	assign \g236542/u3_syn_4  = _w36756_ ;
	assign \g236550/u3_syn_4  = _w36758_ ;
	assign \g236559/u3_syn_4  = _w36760_ ;
	assign \g236567/u3_syn_4  = _w36762_ ;
	assign \g236575/u3_syn_4  = _w36764_ ;
	assign \g236583/u3_syn_4  = _w36766_ ;
	assign \g236591/u3_syn_4  = _w36768_ ;
	assign \g236599/u3_syn_4  = _w36770_ ;
	assign \g236607/u3_syn_4  = _w36772_ ;
	assign \g236608/u3_syn_4  = _w36774_ ;
	assign \g236616/u3_syn_4  = _w36776_ ;
	assign \g236624/u3_syn_4  = _w36778_ ;
	assign \g236632/u3_syn_4  = _w36780_ ;
	assign \g236640/u3_syn_4  = _w36782_ ;
	assign \g236647/u3_syn_4  = _w36783_ ;
	assign \g236649/u3_syn_4  = _w36785_ ;
	assign \g236659/u3_syn_4  = _w36787_ ;
	assign \g236671/u3_syn_4  = _w36789_ ;
	assign \g236677/u3_syn_4  = _w36790_ ;
	assign \g236688/u3_syn_4  = _w36792_ ;
	assign \g236696/u3_syn_4  = _w36794_ ;
	assign \g236705/u3_syn_4  = _w36796_ ;
	assign \g236712/u3_syn_4  = _w36797_ ;
	assign \g236718/u3_syn_4  = _w36799_ ;
	assign \g236729/u3_syn_4  = _w36800_ ;
	assign \g236732/u3_syn_4  = _w36802_ ;
	assign \g236745/u3_syn_4  = _w36804_ ;
	assign \g236753/u3_syn_4  = _w36806_ ;
	assign \g236761/u3_syn_4  = _w36808_ ;
	assign \g236769/u3_syn_4  = _w36810_ ;
	assign \g236777/u3_syn_4  = _w36812_ ;
	assign \g236779/u3_syn_4  = _w36813_ ;
	assign \g236788/u3_syn_4  = _w36815_ ;
	assign \g236800/u3_syn_4  = _w36817_ ;
	assign \g236802/u3_syn_4  = _w36819_ ;
	assign \g236805/u3_syn_4  = _w36820_ ;
	assign \g236813/u3_syn_4  = _w36822_ ;
	assign \g236825/u3_syn_4  = _w36824_ ;
	assign \g236829/u3_syn_4  = _w36825_ ;
	assign \g236837/u3_syn_4  = _w36827_ ;
	assign \g236849/u3_syn_4  = _w36829_ ;
	assign \g236854/u3_syn_4  = _w36830_ ;
	assign \g236860/u3_syn_4  = _w36832_ ;
	assign \g236872/u3_syn_4  = _w36834_ ;
	assign \g236878/u3_syn_4  = _w36835_ ;
	assign \g236884/u3_syn_4  = _w36837_ ;
	assign \g236896/u3_syn_4  = _w36839_ ;
	assign \g236903/u3_syn_4  = _w36840_ ;
	assign \g236908/u3_syn_4  = _w36842_ ;
	assign \g236920/u3_syn_4  = _w36844_ ;
	assign \g236930/u3_syn_4  = _w36846_ ;
	assign \g236939/u3_syn_4  = _w36848_ ;
	assign \g236947/u3_syn_4  = _w36850_ ;
	assign \g236949/u3_syn_4  = _w36851_ ;
	assign \g236956/u3_syn_4  = _w36853_ ;
	assign \g236962/u3_syn_4  = _w36854_ ;
	assign \g236965/u3_syn_4  = _w36856_ ;
	assign \g236980/u3_syn_4  = _w36858_ ;
	assign \g236988/u3_syn_4  = _w36859_ ;
	assign \g236989/u3_syn_4  = _w36861_ ;
	assign \g237004/u3_syn_4  = _w36863_ ;
	assign \g237005/u3_syn_4  = _w36864_ ;
	assign \g237020/u3_syn_4  = _w36865_ ;
	assign \g237021/u3_syn_4  = _w36867_ ;
	assign \g237033/u3_syn_4  = _w36869_ ;
	assign \g237044/u3_syn_4  = _w36870_ ;
	assign \g237045/u3_syn_4  = _w36872_ ;
	assign \g237056/u3_syn_4  = _w36874_ ;
	assign \g237068/u3_syn_4  = _w36876_ ;
	assign \g237076/u3_syn_4  = _w36878_ ;
	assign \g237084/u3_syn_4  = _w36880_ ;
	assign \g237092/u3_syn_4  = _w36881_ ;
	assign \g237095/u3_syn_4  = _w36883_ ;
	assign \g237107/u3_syn_4  = _w36885_ ;
	assign \g237110/u3_syn_4  = _w36886_ ;
	assign \g237119/u3_syn_4  = _w36888_ ;
	assign \g237131/u3_syn_4  = _w36890_ ;
	assign \g237135/u3_syn_4  = _w36891_ ;
	assign \g237148/u3_syn_4  = _w36892_ ;
	assign \g237152/u3_syn_4  = _w36893_ ;
	assign \g237165/u3_syn_4  = _w36894_ ;
	assign \g237168/u3_syn_4  = _w36896_ ;
	assign \g237180/u3_syn_4  = _w36898_ ;
	assign \g237185/u3_syn_4  = _w36899_ ;
	assign \g237192/u3_syn_4  = _w36901_ ;
	assign \g237204/u3_syn_4  = _w36903_ ;
	assign \g237209/u3_syn_4  = _w36904_ ;
	assign \g237215/u3_syn_4  = _w36906_ ;
	assign \g237229/u3_syn_4  = _w36907_ ;
	assign \g237231/u3_syn_4  = _w36909_ ;
	assign \g237245/u3_syn_4  = _w36910_ ;
	assign \g237251/u3_syn_4  = _w36912_ ;
	assign \g237260/u3_syn_4  = _w36913_ ;
	assign \g237262/u3_syn_4  = _w36915_ ;
	assign \g237277/u3_syn_4  = _w36916_ ;
	assign \g237281/u3_syn_4  = _w36918_ ;
	assign \g237293/u3_syn_4  = _w36919_ ;
	assign \g237294/u3_syn_4  = _w36921_ ;
	assign \g237310/u3_syn_4  = _w36922_ ;
	assign \g237311/u3_syn_4  = _w36924_ ;
	assign \g237323/u3_syn_4  = _w36926_ ;
	assign \g237334/u3_syn_4  = _w36928_ ;
	assign \g237342/u3_syn_4  = _w36929_ ;
	assign \g237350/u3_syn_4  = _w36931_ ;
	assign \g237353/u3_syn_4  = _w36932_ ;
	assign \g237359/u3_syn_4  = _w36934_ ;
	assign \g237367/u3_syn_4  = _w36936_ ;
	assign \g237368/u3_syn_4  = _w36937_ ;
	assign \g237378/u3_syn_4  = _w36939_ ;
	assign \g237391/u3_syn_4  = _w36941_ ;
	assign \g237392/u3_syn_4  = _w36942_ ;
	assign \g237403/u3_syn_4  = _w36944_ ;
	assign \g237415/u3_syn_4  = _w36946_ ;
	assign \g237417/u3_syn_4  = _w36947_ ;
	assign \g237431/u3_syn_4  = _w36949_ ;
	assign \g237439/u3_syn_4  = _w36951_ ;
	assign \g237440/u3_syn_4  = _w36952_ ;
	assign \g237454/u3_syn_4  = _w36954_ ;
	assign \g237457/u3_syn_4  = _w36955_ ;
	assign \g237472/u3_syn_4  = _w36957_ ;
	assign \g237480/u3_syn_4  = _w36958_ ;
	assign \g237488/u3_syn_4  = _w36960_ ;
	assign \g237496/u3_syn_4  = _w36961_ ;
	assign \g237499/u3_syn_4  = _w36962_ ;
	assign \g237512/u3_syn_4  = _w36963_ ;
	assign \g237515/u3_syn_4  = _w36965_ ;
	assign \g237525/u3_syn_4  = _w36967_ ;
	assign \g237529/u3_syn_4  = _w36968_ ;
	assign \g237535/u3_syn_4  = _w36970_ ;
	assign \g237541/u3_syn_4  = _w36971_ ;
	assign \g237553/u3_syn_4  = _w36973_ ;
	assign \g237561/u3_syn_4  = _w36974_ ;
	assign \g237569/u3_syn_4  = _w36976_ ;
	assign \g237575/u3_syn_4  = _w36977_ ;
	assign \g237578/u3_syn_4  = _w36978_ ;
	assign \g237581/u3_syn_4  = _w36979_ ;
	assign \g237591/u3_syn_4  = _w36981_ ;
	assign \g237602/u3_syn_4  = _w36983_ ;
	assign \g237610/u3_syn_4  = _w36985_ ;
	assign \g237617/u3_syn_4  = _w36986_ ;
	assign \g237623/u3_syn_4  = _w36987_ ;
	assign \g237633/u3_syn_4  = _w36988_ ;
	assign \g237635/u3_syn_4  = _w36989_ ;
	assign \g237648/u3_syn_4  = _w36990_ ;
	assign \g237658/u3_syn_4  = _w36991_ ;
	assign \g237659/u3_syn_4  = _w36992_ ;
	assign \g237660/u3_syn_4  = _w36993_ ;
	assign \g237668/u3_syn_4  = _w36994_ ;
	assign \g237675/u3_syn_4  = _w36995_ ;
	assign \g237684/u3_syn_4  = _w36996_ ;
	assign \g237692/u3_syn_4  = _w36997_ ;
	assign \g237693/u3_syn_4  = _w36998_ ;
	assign \g237705/u3_syn_4  = _w36999_ ;
	assign \g237716/u3_syn_4  = _w37000_ ;
	assign \g237717/u3_syn_4  = _w37001_ ;
	assign \g237729/u3_syn_4  = _w37002_ ;
	assign \g237740/u3_syn_4  = _w37003_ ;
	assign \g237741/u3_syn_4  = _w37004_ ;
	assign \g237756/u3_syn_4  = _w37005_ ;
	assign \g237764/u3_syn_4  = _w37006_ ;
	assign \g237768/u3_syn_4  = _w37007_ ;
	assign \g237780/u3_syn_4  = _w37008_ ;
	assign \g237782/u3_syn_4  = _w37009_ ;
	assign \g237792/u3_syn_4  = _w37010_ ;
	assign \g237804/u3_syn_4  = _w37011_ ;
	assign \g237812/u3_syn_4  = _w37012_ ;
	assign \g237820/u3_syn_4  = _w37013_ ;
	assign \g237828/u3_syn_4  = _w37014_ ;
	assign \g237836/u3_syn_4  = _w37015_ ;
	assign \g237844/u3_syn_4  = _w37016_ ;
	assign \g237852/u3_syn_4  = _w37017_ ;
	assign \g237860/u3_syn_4  = _w37018_ ;
	assign \g237868/u3_syn_4  = _w37019_ ;
	assign \g237876/u3_syn_4  = _w37020_ ;
	assign \g237884/u3_syn_4  = _w37021_ ;
	assign \g237888/u3_syn_4  = _w37022_ ;
	assign \g237895/u3_syn_4  = _w37023_ ;
	assign \g237907/u3_syn_4  = _w37024_ ;
	assign \g237916/u3_syn_4  = _w37025_ ;
	assign \g237924/u3_syn_4  = _w37026_ ;
	assign \g237931/u3_syn_4  = _w37027_ ;
	assign \g237940/u3_syn_4  = _w37028_ ;
	assign \g237949/u3_syn_4  = _w37029_ ;
	assign \g237950/u3_syn_4  = _w37030_ ;
	assign \g237955/u3_syn_4  = _w37031_ ;
	assign \g237961/u3_syn_4  = _w37032_ ;
	assign \g237965/u3_syn_4  = _w37033_ ;
	assign \g237975/u3_syn_4  = _w37034_ ;
	assign \g237983/u3_syn_4  = _w37035_ ;
	assign \g237989/u3_syn_4  = _w37036_ ;
	assign \g237999/u3_syn_4  = _w37037_ ;
	assign \g238007/u3_syn_4  = _w37038_ ;
	assign \g238015/u3_syn_4  = _w37039_ ;
	assign \g238017/u3_syn_4  = _w37040_ ;
	assign \g238033/u3_syn_4  = _w37041_ ;
	assign \g238035/u3_syn_4  = _w37042_ ;
	assign \g238049/u3_syn_4  = _w37043_ ;
	assign \g238057/u3_syn_4  = _w37044_ ;
	assign \g238065/u3_syn_4  = _w37045_ ;
	assign \g238072/u3_syn_4  = _w37046_ ;
	assign \g238081/u3_syn_4  = _w37047_ ;
	assign \g238082/u3_syn_4  = _w37048_ ;
	assign \g238097/u3_syn_4  = _w37049_ ;
	assign \g238105/u3_syn_4  = _w37050_ ;
	assign \g238113/u3_syn_4  = _w37051_ ;
	assign \g238114/u3_syn_4  = _w37052_ ;
	assign \g238129/u3_syn_4  = _w37053_ ;
	assign \g238137/u3_syn_4  = _w37054_ ;
	assign \g238145/u3_syn_4  = _w37055_ ;
	assign \g238153/u3_syn_4  = _w37056_ ;
	assign \g238161/u3_syn_4  = _w37057_ ;
	assign \g238163/u3_syn_4  = _w37058_ ;
	assign \g238177/u3_syn_4  = _w37059_ ;
	assign \g238179/u3_syn_4  = _w37060_ ;
	assign \g238194/u3_syn_4  = _w37061_ ;
	assign \g238197/u3_syn_4  = _w37062_ ;
	assign \g238209/u3_syn_4  = _w37063_ ;
	assign \g238213/u3_syn_4  = _w37064_ ;
	assign \g238225/u3_syn_4  = _w37065_ ;
	assign \g238229/u3_syn_4  = _w37066_ ;
	assign \g238237/u3_syn_4  = _w37067_ ;
	assign \g238250/u3_syn_4  = _w37068_ ;
	assign \g238257/u3_syn_4  = _w37069_ ;
	assign \g238263/u3_syn_4  = _w37070_ ;
	assign \g238269/u3_syn_4  = _w37071_ ;
	assign \g238282/u3_syn_4  = _w37072_ ;
	assign \g238285/u3_syn_4  = _w37073_ ;
	assign \g238298/u3_syn_4  = _w37074_ ;
	assign \g238301/u3_syn_4  = _w37075_ ;
	assign \g238314/u3_syn_4  = _w37076_ ;
	assign \g238316/u3_syn_4  = _w37077_ ;
	assign \g238329/u3_syn_4  = _w37078_ ;
	assign \g238338/u3_syn_4  = _w37079_ ;
	assign \g238346/u3_syn_4  = _w37080_ ;
	assign \g238351/u3_syn_4  = _w37081_ ;
	assign \g238356/u3_syn_4  = _w37082_ ;
	assign \g238368/u3_syn_4  = _w37083_ ;
	assign \g238378/u3_syn_4  = _w37084_ ;
	assign \g238386/u3_syn_4  = _w37085_ ;
	assign \g238394/u3_syn_4  = _w37086_ ;
	assign \g238402/u3_syn_4  = _w37087_ ;
	assign \g238409/u3_syn_4  = _w37088_ ;
	assign \g238412/u3_syn_4  = _w37089_ ;
	assign \g238427/u3_syn_4  = _w37090_ ;
	assign \g238429/u3_syn_4  = _w37091_ ;
	assign \g238443/u3_syn_4  = _w37092_ ;
	assign \g238448/u3_syn_4  = _w37093_ ;
	assign \g238457/u3_syn_4  = _w37094_ ;
	assign \g238460/u3_syn_4  = _w37095_ ;
	assign \g238472/u3_syn_4  = _w37096_ ;
	assign \g238484/u3_syn_4  = _w37097_ ;
	assign \g238492/u3_syn_4  = _w37098_ ;
	assign \g238500/u3_syn_4  = _w37099_ ;
	assign \g238505/u3_syn_4  = _w37100_ ;
	assign \g238516/u3_syn_4  = _w37101_ ;
	assign \g238524/u3_syn_4  = _w37102_ ;
	assign \g238532/u3_syn_4  = _w37103_ ;
	assign \g238534/u3_syn_4  = _w37104_ ;
	assign \g238544/u3_syn_4  = _w37105_ ;
	assign \g238549/u3_syn_4  = _w37106_ ;
	assign \g238550/u3_syn_4  = _w37107_ ;
	assign \g238565/u3_syn_4  = _w37108_ ;
	assign \g238566/u3_syn_4  = _w37109_ ;
	assign \g238582/u3_syn_4  = _w37110_ ;
	assign \g238583/u3_syn_4  = _w37111_ ;
	assign \g238594/u3_syn_4  = _w37112_ ;
	assign \g238606/u3_syn_4  = _w37113_ ;
	assign \g238614/u3_syn_4  = _w37114_ ;
	assign \g238615/u3_syn_4  = _w37115_ ;
	assign \g238619/u3_syn_4  = _w37116_ ;
	assign \g238631/u3_syn_4  = _w37117_ ;
	assign \g238639/u3_syn_4  = _w37118_ ;
	assign \g238647/u3_syn_4  = _w37119_ ;
	assign \g238649/u3_syn_4  = _w37120_ ;
	assign \g238659/u3_syn_4  = _w37121_ ;
	assign \g238670/u3_syn_4  = _w37122_ ;
	assign \g238671/u3_syn_4  = _w37123_ ;
	assign \g238680/u3_syn_4  = _w37124_ ;
	assign \g238688/u3_syn_4  = _w37125_ ;
	assign \g238691/u3_syn_4  = _w37126_ ;
	assign \g238696/u3_syn_4  = _w37127_ ;
	assign \g238705/u3_syn_4  = _w37128_ ;
	assign \g238708/u3_syn_4  = _w37129_ ;
	assign \g238721/u3_syn_4  = _w37130_ ;
	assign \g238724/u3_syn_4  = _w37131_ ;
	assign \g238736/u3_syn_4  = _w37132_ ;
	assign \g238745/u3_syn_4  = _w37133_ ;
	assign \g238753/u3_syn_4  = _w37134_ ;
	assign \g238757/u3_syn_4  = _w37135_ ;
	assign \g238764/u3_syn_4  = _w37136_ ;
	assign \g238776/u3_syn_4  = _w37137_ ;
	assign \g238781/u3_syn_4  = _w37138_ ;
	assign \g238787/u3_syn_4  = _w37139_ ;
	assign \g238799/u3_syn_4  = _w37140_ ;
	assign \g238807/u3_syn_4  = _w37141_ ;
	assign \g238811/u3_syn_4  = _w37142_ ;
	assign \g238824/u3_syn_4  = _w37143_ ;
	assign \g238830/u3_syn_4  = _w37144_ ;
	assign \g238841/u3_syn_4  = _w37145_ ;
	assign \g238843/u3_syn_4  = _w37146_ ;
	assign \g238855/u3_syn_4  = _w37147_ ;
	assign \g238859/u3_syn_4  = _w37148_ ;
	assign \g238863/u3_syn_4  = _w37149_ ;
	assign \g238868/u3_syn_4  = _w37150_ ;
	assign \g238880/u3_syn_4  = _w37151_ ;
	assign \g238888/u3_syn_4  = _w37152_ ;
	assign \g238892/u3_syn_4  = _w37153_ ;
	assign \g238903/u3_syn_4  = _w37154_ ;
	assign \g238911/u3_syn_4  = _w37155_ ;
	assign \g238915/u3_syn_4  = _w37156_ ;
	assign \g238927/u3_syn_4  = _w37157_ ;
	assign \g238937/u3_syn_4  = _w37158_ ;
	assign \g238945/u3_syn_4  = _w37159_ ;
	assign \g238953/u3_syn_4  = _w37160_ ;
	assign \g238961/u3_syn_4  = _w37161_ ;
	assign \g238970/u3_syn_4  = _w37162_ ;
	assign \g238971/u3_syn_4  = _w37163_ ;
	assign \g238983/u3_syn_4  = _w37164_ ;
	assign \g238994/u3_syn_4  = _w37165_ ;
	assign \g239002/u3_syn_4  = _w37166_ ;
	assign \g239009/u3_syn_4  = _w37167_ ;
	assign \g239015/u3_syn_4  = _w37168_ ;
	assign \g239025/u3_syn_4  = _w37169_ ;
	assign \g239030/u3_syn_4  = _w37170_ ;
	assign \g239041/u3_syn_4  = _w37171_ ;
	assign \g239048/u3_syn_4  = _w37172_ ;
	assign \g239053/u3_syn_4  = _w37173_ ;
	assign \g239065/u3_syn_4  = _w37174_ ;
	assign \g239073/u3_syn_4  = _w37175_ ;
	assign \g239081/u3_syn_4  = _w37176_ ;
	assign \g239082/u3_syn_4  = _w37177_ ;
	assign \g239093/u3_syn_4  = _w37178_ ;
	assign \g239105/u3_syn_4  = _w37179_ ;
	assign \g239108/u3_syn_4  = _w37180_ ;
	assign \g239117/u3_syn_4  = _w37181_ ;
	assign \g239129/u3_syn_4  = _w37182_ ;
	assign \g239137/u3_syn_4  = _w37183_ ;
	assign \g239139/u3_syn_4  = _w37184_ ;
	assign \g239148/u3_syn_4  = _w37185_ ;
	assign \g239160/u3_syn_4  = _w37186_ ;
	assign \g239162/u3_syn_4  = _w37187_ ;
	assign \g239172/u3_syn_4  = _w37188_ ;
	assign \g239184/u3_syn_4  = _w37189_ ;
	assign \g239187/u3_syn_4  = _w37190_ ;
	assign \g239189/u3_syn_4  = _w37191_ ;
	assign \g239201/u3_syn_4  = _w37192_ ;
	assign \g239208/u3_syn_4  = _w37193_ ;
	assign \g239217/u3_syn_4  = _w37194_ ;
	assign \g239219/u3_syn_4  = _w37195_ ;
	assign \g239226/u3_syn_4  = _w37196_ ;
	assign \g239234/u3_syn_4  = _w37197_ ;
	assign \g239242/u3_syn_4  = _w37198_ ;
	assign \g239246/u3_syn_4  = _w37199_ ;
	assign \g239257/u3_syn_4  = _w37200_ ;
	assign \g239258/u3_syn_4  = _w37201_ ;
	assign \g239263/u3_syn_4  = _w37202_ ;
	assign \g239275/u3_syn_4  = _w37203_ ;
	assign \g239277/u3_syn_4  = _w37204_ ;
	assign \g239291/u3_syn_4  = _w37205_ ;
	assign \g239296/u3_syn_4  = _w37206_ ;
	assign \g239308/u3_syn_4  = _w37207_ ;
	assign \g239311/u3_syn_4  = _w37208_ ;
	assign \g239322/u3_syn_4  = _w37209_ ;
	assign \g239329/u3_syn_4  = _w37210_ ;
	assign \g239338/u3_syn_4  = _w37211_ ;
	assign \g239339/u3_syn_4  = _w37212_ ;
	assign \g239346/u3_syn_4  = _w37213_ ;
	assign \g239351/u3_syn_4  = _w37214_ ;
	assign \g239363/u3_syn_4  = _w37215_ ;
	assign \g239370/u3_syn_4  = _w37216_ ;
	assign \g239375/u3_syn_4  = _w37217_ ;
	assign \g239387/u3_syn_4  = _w37218_ ;
	assign \g239395/u3_syn_4  = _w37219_ ;
	assign \g239418/u3_syn_4  = _w37220_ ;
	assign \g239439/u3_syn_4  = _w37221_ ;
	assign \g239442/u3_syn_4  = _w37222_ ;
	assign \g239454/u3_syn_4  = _w37223_ ;
	assign \g239464/u3_syn_4  = _w37224_ ;
	assign \g239470/u3_syn_4  = _w37225_ ;
	assign \g239481/u3_syn_4  = _w37226_ ;
	assign \g239487/u3_syn_4  = _w37227_ ;
	assign \g239497/u3_syn_4  = _w37228_ ;
	assign \g239520/u3_syn_4  = _w37229_ ;
	assign \g239532/u3_syn_4  = _w37230_ ;
	assign \g239543/u3_syn_4  = _w37231_ ;
	assign \g239551/u3_syn_4  = _w37232_ ;
	assign \g239552/u3_syn_4  = _w37233_ ;
	assign \g239567/u3_syn_4  = _w37234_ ;
	assign \g239575/u3_syn_4  = _w37235_ ;
	assign \g239579/u3_syn_4  = _w37236_ ;
	assign \g239592/u3_syn_4  = _w37237_ ;
	assign \g239594/u3_syn_4  = _w37238_ ;
	assign \g239608/u3_syn_4  = _w37239_ ;
	assign \g239626/u3_syn_4  = _w37240_ ;
	assign \g239634/u3_syn_4  = _w37241_ ;
	assign \g239646/u3_syn_4  = _w37242_ ;
	assign \g239649/u3_syn_4  = _w37243_ ;
	assign \g239657/u3_syn_4  = _w37244_ ;
	assign \g239670/u3_syn_4  = _w37245_ ;
	assign \g239673/u3_syn_4  = _w37246_ ;
	assign \g239686/u3_syn_4  = _w37247_ ;
	assign \g239694/u3_syn_4  = _w37248_ ;
	assign \g239695/u3_syn_4  = _w37249_ ;
	assign \g239701/u3_syn_4  = _w37250_ ;
	assign \g239705/u3_syn_4  = _w37251_ ;
	assign \g239709/u3_syn_4  = _w37252_ ;
	assign \g239715/u3_syn_4  = _w37253_ ;
	assign \g239717/u3_syn_4  = _w37254_ ;
	assign \g239726/u3_syn_4  = _w37255_ ;
	assign \g239734/u3_syn_4  = _w37256_ ;
	assign \g239735/u3_syn_4  = _w37257_ ;
	assign \g239743/u3_syn_4  = _w37258_ ;
	assign \g239760/u3_syn_4  = _w37259_ ;
	assign \g239768/u3_syn_4  = _w37260_ ;
	assign \g239776/u3_syn_4  = _w37261_ ;
	assign \g239784/u3_syn_4  = _w37262_ ;
	assign \g239793/u3_syn_4  = _w37263_ ;
	assign \g239801/u3_syn_4  = _w37264_ ;
	assign \g239817/u3_syn_4  = _w37265_ ;
	assign \g239818/u3_syn_4  = _w37266_ ;
	assign \g239848/u3_syn_4  = _w37267_ ;
	assign \g239856/u3_syn_4  = _w37268_ ;
	assign \g239872/u3_syn_4  = _w37269_ ;
	assign \g239880/u3_syn_4  = _w37270_ ;
	assign \g239888/u3_syn_4  = _w37271_ ;
	assign \g239896/u3_syn_4  = _w37272_ ;
	assign \g239904/u3_syn_4  = _w37273_ ;
	assign \g239912/u3_syn_4  = _w37274_ ;
	assign \g239920/u3_syn_4  = _w37275_ ;
	assign \g239928/u3_syn_4  = _w37276_ ;
	assign \g239936/u3_syn_4  = _w37277_ ;
	assign \g239951/u3_syn_4  = _w37278_ ;
	assign \g239963/u3_syn_4  = _w37279_ ;
	assign \g239979/u3_syn_4  = _w37280_ ;
	assign \g239986/u3_syn_4  = _w37281_ ;
	assign \g239999/u3_syn_4  = _w37282_ ;
	assign \g240000/u3_syn_4  = _w37283_ ;
	assign \g240008/u3_syn_4  = _w37284_ ;
	assign \g240012/u3_syn_4  = _w37285_ ;
	assign \g240018/u3_syn_4  = _w37286_ ;
	assign \g240026/u3_syn_4  = _w37287_ ;
	assign \g240034/u3_syn_4  = _w37288_ ;
	assign \g240042/u3_syn_4  = _w37289_ ;
	assign \g240050/u3_syn_4  = _w37290_ ;
	assign \g240074/u3_syn_4  = _w37291_ ;
	assign \g240091/u3_syn_4  = _w37292_ ;
	assign \g240122/u3_syn_4  = _w37293_ ;
	assign \g240147/u3_syn_4  = _w37294_ ;
	assign \g240209/u3_syn_4  = _w37295_ ;
	assign \g240219/u3_syn_4  = _w37296_ ;
	assign \g240259/u3_syn_4  = _w37297_ ;
	assign \g240334/u3_syn_4  = _w37298_ ;
	assign \g240406/u3_syn_4  = _w37299_ ;
	assign \g240416/u3_syn_4  = _w37300_ ;
	assign \g240424/u3_syn_4  = _w37301_ ;
	assign \g240432/u3_syn_4  = _w37302_ ;
	assign \g240440/u3_syn_4  = _w37303_ ;
	assign \g240448/u3_syn_4  = _w37304_ ;
	assign \g240456/u3_syn_4  = _w37305_ ;
	assign \g240464/u3_syn_4  = _w37306_ ;
	assign \g240472/u3_syn_4  = _w37307_ ;
	assign \g240480/u3_syn_4  = _w37308_ ;
	assign \g240488/u3_syn_4  = _w37309_ ;
	assign \g240496/u3_syn_4  = _w37310_ ;
	assign \g240504/u3_syn_4  = _w37311_ ;
	assign \g240512/u3_syn_4  = _w37312_ ;
	assign \g240520/u3_syn_4  = _w37313_ ;
	assign \g240530/u3_syn_4  = _w37314_ ;
	assign \g240538/u3_syn_4  = _w37315_ ;
	assign \g240547/u3_syn_4  = _w37316_ ;
	assign \g240555/u3_syn_4  = _w37317_ ;
	assign \g240563/u3_syn_4  = _w37318_ ;
	assign \g240571/u3_syn_4  = _w37319_ ;
	assign \g240579/u3_syn_4  = _w37320_ ;
	assign \g240587/u3_syn_4  = _w37321_ ;
	assign \g240595/u3_syn_4  = _w37322_ ;
	assign \g240603/u3_syn_4  = _w37323_ ;
	assign \g240611/u3_syn_4  = _w37324_ ;
	assign \g240619/u3_syn_4  = _w37325_ ;
	assign \g240627/u3_syn_4  = _w37326_ ;
	assign \g240635/u3_syn_4  = _w37327_ ;
	assign \g240643/u3_syn_4  = _w37328_ ;
	assign \g240651/u3_syn_4  = _w37329_ ;
	assign \g240659/u3_syn_4  = _w37330_ ;
	assign \g240667/u3_syn_4  = _w37331_ ;
	assign \g240675/u3_syn_4  = _w37332_ ;
	assign \g240683/u3_syn_4  = _w37333_ ;
	assign \g240691/u3_syn_4  = _w37334_ ;
	assign \g240699/u3_syn_4  = _w37335_ ;
	assign \g240707/u3_syn_4  = _w37336_ ;
	assign \g240715/u3_syn_4  = _w37337_ ;
	assign \g240723/u3_syn_4  = _w37338_ ;
	assign \g240731/u3_syn_4  = _w37339_ ;
	assign \g240739/u3_syn_4  = _w37340_ ;
	assign \g240747/u3_syn_4  = _w37341_ ;
	assign \g240755/u3_syn_4  = _w37342_ ;
	assign \g240763/u3_syn_4  = _w37343_ ;
	assign \g240771/u3_syn_4  = _w37344_ ;
	assign \g240779/u3_syn_4  = _w37345_ ;
	assign \g240787/u3_syn_4  = _w37346_ ;
	assign \g240795/u3_syn_4  = _w37347_ ;
	assign \g240803/u3_syn_4  = _w37348_ ;
	assign \g240811/u3_syn_4  = _w37349_ ;
	assign \g240819/u3_syn_4  = _w37350_ ;
	assign \g240827/u3_syn_4  = _w37351_ ;
	assign \g240835/u3_syn_4  = _w37352_ ;
	assign \g240843/u3_syn_4  = _w37353_ ;
	assign \g240851/u3_syn_4  = _w37354_ ;
	assign \g240859/u3_syn_4  = _w37355_ ;
	assign \g240867/u3_syn_4  = _w37356_ ;
	assign \g240875/u3_syn_4  = _w37357_ ;
	assign \g240883/u3_syn_4  = _w37358_ ;
	assign \g240891/u3_syn_4  = _w37359_ ;
	assign \g240899/u3_syn_4  = _w37360_ ;
	assign \g240907/u3_syn_4  = _w37361_ ;
	assign \g240915/u3_syn_4  = _w37362_ ;
	assign \g240923/u3_syn_4  = _w37363_ ;
	assign \g240931/u3_syn_4  = _w37364_ ;
	assign \g240939/u3_syn_4  = _w37365_ ;
	assign \g240947/u3_syn_4  = _w37366_ ;
	assign \g240955/u3_syn_4  = _w37367_ ;
	assign \g240963/u3_syn_4  = _w37368_ ;
	assign \g240971/u3_syn_4  = _w37369_ ;
	assign \g240979/u3_syn_4  = _w37370_ ;
	assign \g240987/u3_syn_4  = _w37371_ ;
	assign \g240995/u3_syn_4  = _w37372_ ;
	assign \g241003/u3_syn_4  = _w37373_ ;
	assign \g241011/u3_syn_4  = _w37374_ ;
	assign \g241019/u3_syn_4  = _w37375_ ;
	assign \g241027/u3_syn_4  = _w37376_ ;
	assign \g241036/u3_syn_4  = _w37377_ ;
	assign \g241044/u3_syn_4  = _w37378_ ;
	assign \g241052/u3_syn_4  = _w37379_ ;
	assign \g241060/u3_syn_4  = _w37380_ ;
	assign \g241068/u3_syn_4  = _w37381_ ;
	assign \g241076/u3_syn_4  = _w37382_ ;
	assign \g241084/u3_syn_4  = _w37383_ ;
	assign \g241092/u3_syn_4  = _w37384_ ;
	assign \g241100/u3_syn_4  = _w37385_ ;
	assign \g241108/u3_syn_4  = _w37386_ ;
	assign \g241116/u3_syn_4  = _w37387_ ;
	assign \g241124/u3_syn_4  = _w37388_ ;
	assign \g241132/u3_syn_4  = _w37389_ ;
	assign \g241140/u3_syn_4  = _w37390_ ;
	assign \g241148/u3_syn_4  = _w37391_ ;
	assign \g241156/u3_syn_4  = _w37392_ ;
	assign \g241164/u3_syn_4  = _w37393_ ;
	assign \g241172/u3_syn_4  = _w37394_ ;
	assign \g241180/u3_syn_4  = _w37395_ ;
	assign \g241188/u3_syn_4  = _w37396_ ;
	assign \g241196/u3_syn_4  = _w37397_ ;
	assign \g241205/u3_syn_4  = _w37398_ ;
	assign \g241213/u3_syn_4  = _w37399_ ;
	assign \g241221/u3_syn_4  = _w37400_ ;
	assign \g241229/u3_syn_4  = _w37401_ ;
	assign \g241237/u3_syn_4  = _w37402_ ;
	assign \g241245/u3_syn_4  = _w37403_ ;
	assign \g241253/u3_syn_4  = _w37404_ ;
	assign \g241261/u3_syn_4  = _w37405_ ;
	assign \g241269/u3_syn_4  = _w37406_ ;
	assign \g241277/u3_syn_4  = _w37407_ ;
	assign \g241285/u3_syn_4  = _w37408_ ;
	assign \g241293/u3_syn_4  = _w37409_ ;
	assign \g241301/u3_syn_4  = _w37410_ ;
	assign \g241309/u3_syn_4  = _w37411_ ;
	assign \g241317/u3_syn_4  = _w37412_ ;
	assign \g241325/u3_syn_4  = _w37413_ ;
	assign \g241333/u3_syn_4  = _w37414_ ;
	assign \g241341/u3_syn_4  = _w37415_ ;
	assign \g241349/u3_syn_4  = _w37416_ ;
	assign \g241358/u3_syn_4  = _w37417_ ;
	assign \g241366/u3_syn_4  = _w37418_ ;
	assign \g241374/u3_syn_4  = _w37419_ ;
	assign \g241382/u3_syn_4  = _w37420_ ;
	assign \g241390/u3_syn_4  = _w37421_ ;
	assign \g241398/u3_syn_4  = _w37422_ ;
	assign \g241406/u3_syn_4  = _w37423_ ;
	assign \g241415/u3_syn_4  = _w37424_ ;
	assign \g241424/u3_syn_4  = _w37425_ ;
	assign \g241433/u3_syn_4  = _w37426_ ;
	assign \g241441/u3_syn_4  = _w37427_ ;
	assign \g241449/u3_syn_4  = _w37428_ ;
	assign \g241459/u3_syn_4  = _w37429_ ;
	assign \g241470/u3_syn_4  = _w37430_ ;
	assign \g241480/u3_syn_4  = _w37431_ ;
	assign \g241489/u3_syn_4  = _w37432_ ;
	assign \g241497/u3_syn_4  = _w37433_ ;
	assign \g241505/u3_syn_4  = _w37434_ ;
	assign \g241513/u3_syn_4  = _w37435_ ;
	assign \g241545/_3_  = _w11477_ ;
	assign \g241580/_00_  = _w37439_ ;
	assign \g241737/_0_  = _w37440_ ;
	assign \g241752/_0_  = _w37441_ ;
	assign \g241755/_0_  = _w35933_ ;
	assign \g241767/_2__syn_2  = _w37442_ ;
	assign \g241781/_1__syn_2  = _w37443_ ;
	assign \g241782/_0_  = _w35938_ ;
	assign \g241803/_1__syn_2  = _w37444_ ;
	assign \g241805/_0_  = _w37445_ ;
	assign \g241812/_1__syn_2  = _w37446_ ;
	assign \g241814/_1__syn_2  = _w37447_ ;
	assign \g241816/_1__syn_2  = _w37448_ ;
	assign \g241819/_1__syn_2  = _w37449_ ;
	assign \g241822/_1__syn_2  = _w37450_ ;
	assign \g241823/_0_  = _w37451_ ;
	assign \g241833/_1__syn_2  = _w37452_ ;
	assign \g241843/_1__syn_2  = _w37454_ ;
	assign \g241844/_1__syn_2  = _w37455_ ;
	assign \g241848/_1__syn_2  = _w37456_ ;
	assign \g241855/_1__syn_2  = _w37457_ ;
	assign \g241868/_1__syn_2  = _w37458_ ;
	assign \g242013/_1__syn_2  = _w37459_ ;
	assign \g242015/_1__syn_2  = _w37460_ ;
	assign \g242017/_1__syn_2  = _w37461_ ;
	assign \g242021/_1__syn_2  = _w37462_ ;
	assign \g242039/_1__syn_2  = _w37463_ ;
	assign \g242081/_0_  = _w37469_ ;
	assign \g242086/_0_  = _w37470_ ;
	assign \g242101/_3_  = _w11640_ ;
	assign \g242116/_0_  = _w37475_ ;
	assign \g242135/_2_  = _w31852_ ;
	assign \g242147/_0_  = _w37481_ ;
	assign \g242158/_0_  = _w37486_ ;
	assign \g242196/_0_  = _w37491_ ;
	assign \g242202/_0_  = _w37506_ ;
	assign \g242203/_0_  = _w37521_ ;
	assign \g242204/_0_  = _w37536_ ;
	assign \g242212/_0_  = _w37539_ ;
	assign \g242226/_01_  = _w37567_ ;
	assign \g242281/_0_  = _w10568_ ;
	assign \g242407/_0_  = _w37571_ ;
	assign \g242410/_0_  = _w37574_ ;
	assign \g242426/_0_  = _w37585_ ;
	assign \g242438/_2_  = _w37586_ ;
	assign \g242466/_0_  = _w37589_ ;
	assign \g242530/_0_  = _w37593_ ;
	assign \g242532/_0_  = _w37594_ ;
	assign \g243397/_0_  = _w37602_ ;
	assign \g245925/_0_  = _w37608_ ;
	assign \g245932/_0_  = _w37614_ ;
	assign \g245933/_0_  = _w37620_ ;
	assign \g245986/_3_  = _w37628_ ;
	assign \g250157/_3_  = _w11488_ ;
	assign \g250202/_0_  = _w37634_ ;
	assign \g250246/_1_  = _w34888_ ;
	assign \g250248/_0_  = _w37639_ ;
	assign \g250250/_0_  = _w37640_ ;
	assign \g250305/_0_  = _w37643_ ;
	assign \g250323/_0_  = _w37646_ ;
	assign \g250373/_0_  = _w37650_ ;
	assign \g250377/_0_  = _w37651_ ;
	assign \g250412/_0_  = _w37658_ ;
	assign \g250413/_0_  = _w37661_ ;
	assign \g250418/_0_  = _w37665_ ;
	assign \g250419/_0_  = _w37667_ ;
	assign \g250421/_0_  = _w37670_ ;
	assign \g250433/_0_  = _w37677_ ;
	assign \g250448/_3_  = _w37681_ ;
	assign \g250567/_3_  = _w11492_ ;
	assign \g258965/_0_  = _w37683_ ;
	assign \g259006/_0_  = _w37687_ ;
	assign \g259471/_0_  = _w37691_ ;
	assign \g259473/_2_  = _w36080_ ;
	assign \g260557/_0_  = _w37692_ ;
	assign \g261035/_0_  = _w37693_ ;
	assign \g261095/_3_  = _w37699_ ;
	assign \g261207/_2__syn_2  = _w37700_ ;
	assign \g261754/_0_  = _w37701_ ;
	assign \g262017/_0_  = _w37706_ ;
	assign \g262045/_0_  = _w37711_ ;
	assign \g262046/_0_  = _w37713_ ;
	assign \g262100/_3_  = _w37716_ ;
	assign \g263539/_1_  = _w15176_ ;
	assign \g263574/_0_  = _w12656_ ;
	assign \g263858/_0_  = _w11110_ ;
	assign \g264104/_1_  = _w37625_ ;
	assign \g264107/_1_  = _w35898_ ;
	assign \g264117/_0_  = _w37718_ ;
	assign \g264282/_0_  = _w34266_ ;
	assign \g264511/_0_  = _w37720_ ;
	assign \g264541/_0_  = _w37724_ ;
	assign \g264562/_0_  = _w37727_ ;
	assign \g264618/_0_  = _w37729_ ;
	assign \g264660/_0_  = _w37731_ ;
	assign \g264681/_3_  = _w37734_ ;
	assign \g264727/_0_  = _w37736_ ;
	assign \g265013/_0_  = _w37738_ ;
	assign \g265084/_0_  = _w37740_ ;
	assign \g265378/_0_  = _w37742_ ;
	assign \g265413/_0_  = _w37744_ ;
	assign \g265446/_0_  = _w37746_ ;
	assign \g265486/_0_  = _w37749_ ;
	assign \g265524/_3_  = _w10666_ ;
	assign \g265528/_3_  = _w11229_ ;
	assign \g265548/_3_  = _w10655_ ;
	assign \g265579/_0_  = _w11495_ ;
	assign \g265768/_0_  = _w37649_ ;
	assign \g265801/_0_  = _w12240_ ;
	assign \g265819/_1_  = _w34199_ ;
	assign \g265853/_0_  = _w37741_ ;
	assign \g265933/_0_  = _w37750_ ;
	assign \g266022/_0_  = _w37751_ ;
	assign \g266183/_1_  = _w34968_ ;
	assign \g281909/_0_  = _w37771_ ;
	assign \g281965/_1_  = _w30479_ ;
	assign \g282284/_1_  = _w29947_ ;
	assign \g282639/_1_  = _w27980_ ;
	assign \g283047/_0_  = _w37775_ ;
	assign \g283157/_1_  = _w23494_ ;
	assign \g283184/_0_  = _w37797_ ;
	assign \g283334/_3_  = _w37802_ ;
	assign int_o_pad = _w37815_ ;
	assign \m_wb_adr_o[0]_pad  = 1'b0;
	assign \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131_syn_2  = \maccontrol1_transmitcontrol1_ByteCnt_reg[0]/NET0131 ;
	assign \wishbone_tx_fifo_fifo_reg[2][15]/P0001_reg_syn_3  = _w37818_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][16]/P0001_reg_syn_3  = _w37821_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][17]/P0001_reg_syn_3  = _w37824_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][22]/P0001_reg_syn_3  = _w37827_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][23]/P0001_reg_syn_3  = _w37830_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][25]/P0001_reg_syn_3  = _w37833_ ;
	assign \wishbone_tx_fifo_fifo_reg[2][2]/P0001_reg_syn_3  = _w37836_ ;
endmodule;