module top( \FP_R_reg[10]/P0001  , \FP_R_reg[11]/P0001  , \FP_R_reg[12]/P0001  , \FP_R_reg[13]/P0001  , \FP_R_reg[14]/P0001  , \FP_R_reg[15]/P0001  , \FP_R_reg[16]/P0001  , \FP_R_reg[17]/P0001  , \FP_R_reg[18]/P0001  , \FP_R_reg[19]/P0001  , \FP_R_reg[1]/P0001  , \FP_R_reg[20]/P0001  , \FP_R_reg[21]/P0001  , \FP_R_reg[22]/P0001  , \FP_R_reg[23]/P0001  , \FP_R_reg[24]/P0001  , \FP_R_reg[25]/P0001  , \FP_R_reg[26]/P0001  , \FP_R_reg[27]/P0001  , \FP_R_reg[28]/P0001  , \FP_R_reg[29]/P0001  , \FP_R_reg[2]/P0001  , \FP_R_reg[30]/P0001  , \FP_R_reg[31]/P0001  , \FP_R_reg[32]/P0001  , \FP_R_reg[33]/NET0131  , \FP_R_reg[34]/NET0131  , \FP_R_reg[35]/NET0131  , \FP_R_reg[36]/NET0131  , \FP_R_reg[37]/NET0131  , \FP_R_reg[38]/NET0131  , \FP_R_reg[39]/NET0131  , \FP_R_reg[3]/P0001  , \FP_R_reg[40]/NET0131  , \FP_R_reg[41]/NET0131  , \FP_R_reg[42]/NET0131  , \FP_R_reg[43]/NET0131  , \FP_R_reg[44]/NET0131  , \FP_R_reg[45]/NET0131  , \FP_R_reg[46]/NET0131  , \FP_R_reg[47]/NET0131  , \FP_R_reg[48]/NET0131  , \FP_R_reg[49]/NET0131  , \FP_R_reg[4]/P0001  , \FP_R_reg[50]/NET0131  , \FP_R_reg[51]/NET0131  , \FP_R_reg[52]/NET0131  , \FP_R_reg[53]/NET0131  , \FP_R_reg[54]/NET0131  , \FP_R_reg[55]/NET0131  , \FP_R_reg[56]/NET0131  , \FP_R_reg[57]/NET0131  , \FP_R_reg[58]/NET0131  , \FP_R_reg[59]/NET0131  , \FP_R_reg[5]/P0001  , \FP_R_reg[60]/NET0131  , \FP_R_reg[61]/NET0131  , \FP_R_reg[62]/NET0131  , \FP_R_reg[63]/NET0131  , \FP_R_reg[64]/NET0131  , \FP_R_reg[6]/P0001  , \FP_R_reg[7]/P0001  , \FP_R_reg[8]/P0001  , \FP_R_reg[9]/P0001  , decrypt_pad , \desIn[0]_pad  , \desIn[10]_pad  , \desIn[11]_pad  , \desIn[12]_pad  , \desIn[13]_pad  , \desIn[14]_pad  , \desIn[15]_pad  , \desIn[16]_pad  , \desIn[17]_pad  , \desIn[18]_pad  , \desIn[19]_pad  , \desIn[1]_pad  , \desIn[20]_pad  , \desIn[21]_pad  , \desIn[22]_pad  , \desIn[23]_pad  , \desIn[24]_pad  , \desIn[25]_pad  , \desIn[26]_pad  , \desIn[27]_pad  , \desIn[28]_pad  , \desIn[29]_pad  , \desIn[2]_pad  , \desIn[30]_pad  , \desIn[31]_pad  , \desIn[32]_pad  , \desIn[33]_pad  , \desIn[34]_pad  , \desIn[35]_pad  , \desIn[36]_pad  , \desIn[37]_pad  , \desIn[38]_pad  , \desIn[39]_pad  , \desIn[3]_pad  , \desIn[40]_pad  , \desIn[41]_pad  , \desIn[42]_pad  , \desIn[43]_pad  , \desIn[44]_pad  , \desIn[45]_pad  , \desIn[46]_pad  , \desIn[47]_pad  , \desIn[48]_pad  , \desIn[49]_pad  , \desIn[4]_pad  , \desIn[50]_pad  , \desIn[51]_pad  , \desIn[52]_pad  , \desIn[53]_pad  , \desIn[54]_pad  , \desIn[55]_pad  , \desIn[56]_pad  , \desIn[57]_pad  , \desIn[58]_pad  , \desIn[59]_pad  , \desIn[5]_pad  , \desIn[60]_pad  , \desIn[61]_pad  , \desIn[62]_pad  , \desIn[63]_pad  , \desIn[6]_pad  , \desIn[7]_pad  , \desIn[8]_pad  , \desIn[9]_pad  , \key1[0]_pad  , \key1[10]_pad  , \key1[11]_pad  , \key1[12]_pad  , \key1[13]_pad  , \key1[14]_pad  , \key1[15]_pad  , \key1[16]_pad  , \key1[17]_pad  , \key1[18]_pad  , \key1[19]_pad  , \key1[1]_pad  , \key1[20]_pad  , \key1[21]_pad  , \key1[22]_pad  , \key1[23]_pad  , \key1[24]_pad  , \key1[25]_pad  , \key1[26]_pad  , \key1[27]_pad  , \key1[28]_pad  , \key1[29]_pad  , \key1[2]_pad  , \key1[30]_pad  , \key1[31]_pad  , \key1[32]_pad  , \key1[33]_pad  , \key1[34]_pad  , \key1[35]_pad  , \key1[36]_pad  , \key1[37]_pad  , \key1[38]_pad  , \key1[39]_pad  , \key1[3]_pad  , \key1[40]_pad  , \key1[41]_pad  , \key1[42]_pad  , \key1[43]_pad  , \key1[44]_pad  , \key1[45]_pad  , \key1[46]_pad  , \key1[47]_pad  , \key1[48]_pad  , \key1[49]_pad  , \key1[4]_pad  , \key1[50]_pad  , \key1[51]_pad  , \key1[52]_pad  , \key1[53]_pad  , \key1[54]_pad  , \key1[55]_pad  , \key1[5]_pad  , \key1[6]_pad  , \key1[7]_pad  , \key1[8]_pad  , \key1[9]_pad  , \key2[0]_pad  , \key2[10]_pad  , \key2[11]_pad  , \key2[12]_pad  , \key2[13]_pad  , \key2[14]_pad  , \key2[15]_pad  , \key2[16]_pad  , \key2[17]_pad  , \key2[18]_pad  , \key2[19]_pad  , \key2[1]_pad  , \key2[20]_pad  , \key2[21]_pad  , \key2[22]_pad  , \key2[23]_pad  , \key2[24]_pad  , \key2[25]_pad  , \key2[26]_pad  , \key2[27]_pad  , \key2[28]_pad  , \key2[29]_pad  , \key2[2]_pad  , \key2[30]_pad  , \key2[31]_pad  , \key2[32]_pad  , \key2[33]_pad  , \key2[34]_pad  , \key2[35]_pad  , \key2[36]_pad  , \key2[37]_pad  , \key2[38]_pad  , \key2[39]_pad  , \key2[3]_pad  , \key2[40]_pad  , \key2[41]_pad  , \key2[42]_pad  , \key2[43]_pad  , \key2[44]_pad  , \key2[45]_pad  , \key2[46]_pad  , \key2[47]_pad  , \key2[48]_pad  , \key2[49]_pad  , \key2[4]_pad  , \key2[50]_pad  , \key2[51]_pad  , \key2[52]_pad  , \key2[53]_pad  , \key2[54]_pad  , \key2[55]_pad  , \key2[5]_pad  , \key2[6]_pad  , \key2[7]_pad  , \key2[8]_pad  , \key2[9]_pad  , \key3[0]_pad  , \key3[10]_pad  , \key3[11]_pad  , \key3[12]_pad  , \key3[13]_pad  , \key3[14]_pad  , \key3[15]_pad  , \key3[16]_pad  , \key3[17]_pad  , \key3[18]_pad  , \key3[19]_pad  , \key3[1]_pad  , \key3[20]_pad  , \key3[21]_pad  , \key3[22]_pad  , \key3[23]_pad  , \key3[24]_pad  , \key3[25]_pad  , \key3[26]_pad  , \key3[27]_pad  , \key3[28]_pad  , \key3[29]_pad  , \key3[2]_pad  , \key3[30]_pad  , \key3[31]_pad  , \key3[32]_pad  , \key3[33]_pad  , \key3[34]_pad  , \key3[35]_pad  , \key3[36]_pad  , \key3[37]_pad  , \key3[38]_pad  , \key3[39]_pad  , \key3[3]_pad  , \key3[40]_pad  , \key3[41]_pad  , \key3[42]_pad  , \key3[43]_pad  , \key3[44]_pad  , \key3[45]_pad  , \key3[46]_pad  , \key3[47]_pad  , \key3[48]_pad  , \key3[49]_pad  , \key3[4]_pad  , \key3[50]_pad  , \key3[51]_pad  , \key3[52]_pad  , \key3[53]_pad  , \key3[54]_pad  , \key3[55]_pad  , \key3[5]_pad  , \key3[6]_pad  , \key3[7]_pad  , \key3[8]_pad  , \key3[9]_pad  , \roundSel[0]_pad  , \roundSel[1]_pad  , \roundSel[2]_pad  , \roundSel[3]_pad  , \roundSel[4]_pad  , \roundSel[5]_pad  , \_al_n0  , \_al_n1  , \desOut[0]_pad  , \desOut[11]_pad  , \desOut[12]_pad  , \desOut[13]_pad  , \desOut[14]_pad  , \desOut[15]_pad  , \desOut[18]_pad  , \desOut[1]_pad  , \desOut[22]_pad  , \desOut[23]_pad  , \desOut[24]_pad  , \desOut[25]_pad  , \desOut[26]_pad  , \desOut[28]_pad  , \desOut[2]_pad  , \desOut[30]_pad  , \desOut[32]_pad  , \desOut[34]_pad  , \desOut[35]_pad  , \desOut[37]_pad  , \desOut[38]_pad  , \desOut[39]_pad  , \desOut[3]_pad  , \desOut[40]_pad  , \desOut[42]_pad  , \desOut[44]_pad  , \desOut[45]_pad  , \desOut[46]_pad  , \desOut[48]_pad  , \desOut[4]_pad  , \desOut[50]_pad  , \desOut[52]_pad  , \desOut[54]_pad  , \desOut[56]_pad  , \desOut[57]_pad  , \desOut[59]_pad  , \desOut[5]_pad  , \desOut[60]_pad  , \desOut[61]_pad  , \desOut[63]_pad  , \desOut[6]_pad  , \desOut[8]_pad  , \desOut[9]_pad  , \g13525_dup/_0_  , \g13583_dup/_0_  , \g17813/_3_  , \g17816/_3_  , \g17819/_3_  , \g17822/_3_  , \g17836/_3_  , \g17871/_3_  , \g17878/_1_  , \g17881/_3_  , \g17966/_2_  , \g17969/_3_  , \g17996/_2_  , \g19574_dup/_3_  , \g19619_dup/_3_  , \g19756_dup/_3_  , \g20263/_3_  , \g20541/_2_  , \g20691/_1_  , \g20740_dup/_3_  , \g67/_2_  );
  input \FP_R_reg[10]/P0001  ;
  input \FP_R_reg[11]/P0001  ;
  input \FP_R_reg[12]/P0001  ;
  input \FP_R_reg[13]/P0001  ;
  input \FP_R_reg[14]/P0001  ;
  input \FP_R_reg[15]/P0001  ;
  input \FP_R_reg[16]/P0001  ;
  input \FP_R_reg[17]/P0001  ;
  input \FP_R_reg[18]/P0001  ;
  input \FP_R_reg[19]/P0001  ;
  input \FP_R_reg[1]/P0001  ;
  input \FP_R_reg[20]/P0001  ;
  input \FP_R_reg[21]/P0001  ;
  input \FP_R_reg[22]/P0001  ;
  input \FP_R_reg[23]/P0001  ;
  input \FP_R_reg[24]/P0001  ;
  input \FP_R_reg[25]/P0001  ;
  input \FP_R_reg[26]/P0001  ;
  input \FP_R_reg[27]/P0001  ;
  input \FP_R_reg[28]/P0001  ;
  input \FP_R_reg[29]/P0001  ;
  input \FP_R_reg[2]/P0001  ;
  input \FP_R_reg[30]/P0001  ;
  input \FP_R_reg[31]/P0001  ;
  input \FP_R_reg[32]/P0001  ;
  input \FP_R_reg[33]/NET0131  ;
  input \FP_R_reg[34]/NET0131  ;
  input \FP_R_reg[35]/NET0131  ;
  input \FP_R_reg[36]/NET0131  ;
  input \FP_R_reg[37]/NET0131  ;
  input \FP_R_reg[38]/NET0131  ;
  input \FP_R_reg[39]/NET0131  ;
  input \FP_R_reg[3]/P0001  ;
  input \FP_R_reg[40]/NET0131  ;
  input \FP_R_reg[41]/NET0131  ;
  input \FP_R_reg[42]/NET0131  ;
  input \FP_R_reg[43]/NET0131  ;
  input \FP_R_reg[44]/NET0131  ;
  input \FP_R_reg[45]/NET0131  ;
  input \FP_R_reg[46]/NET0131  ;
  input \FP_R_reg[47]/NET0131  ;
  input \FP_R_reg[48]/NET0131  ;
  input \FP_R_reg[49]/NET0131  ;
  input \FP_R_reg[4]/P0001  ;
  input \FP_R_reg[50]/NET0131  ;
  input \FP_R_reg[51]/NET0131  ;
  input \FP_R_reg[52]/NET0131  ;
  input \FP_R_reg[53]/NET0131  ;
  input \FP_R_reg[54]/NET0131  ;
  input \FP_R_reg[55]/NET0131  ;
  input \FP_R_reg[56]/NET0131  ;
  input \FP_R_reg[57]/NET0131  ;
  input \FP_R_reg[58]/NET0131  ;
  input \FP_R_reg[59]/NET0131  ;
  input \FP_R_reg[5]/P0001  ;
  input \FP_R_reg[60]/NET0131  ;
  input \FP_R_reg[61]/NET0131  ;
  input \FP_R_reg[62]/NET0131  ;
  input \FP_R_reg[63]/NET0131  ;
  input \FP_R_reg[64]/NET0131  ;
  input \FP_R_reg[6]/P0001  ;
  input \FP_R_reg[7]/P0001  ;
  input \FP_R_reg[8]/P0001  ;
  input \FP_R_reg[9]/P0001  ;
  input decrypt_pad ;
  input \desIn[0]_pad  ;
  input \desIn[10]_pad  ;
  input \desIn[11]_pad  ;
  input \desIn[12]_pad  ;
  input \desIn[13]_pad  ;
  input \desIn[14]_pad  ;
  input \desIn[15]_pad  ;
  input \desIn[16]_pad  ;
  input \desIn[17]_pad  ;
  input \desIn[18]_pad  ;
  input \desIn[19]_pad  ;
  input \desIn[1]_pad  ;
  input \desIn[20]_pad  ;
  input \desIn[21]_pad  ;
  input \desIn[22]_pad  ;
  input \desIn[23]_pad  ;
  input \desIn[24]_pad  ;
  input \desIn[25]_pad  ;
  input \desIn[26]_pad  ;
  input \desIn[27]_pad  ;
  input \desIn[28]_pad  ;
  input \desIn[29]_pad  ;
  input \desIn[2]_pad  ;
  input \desIn[30]_pad  ;
  input \desIn[31]_pad  ;
  input \desIn[32]_pad  ;
  input \desIn[33]_pad  ;
  input \desIn[34]_pad  ;
  input \desIn[35]_pad  ;
  input \desIn[36]_pad  ;
  input \desIn[37]_pad  ;
  input \desIn[38]_pad  ;
  input \desIn[39]_pad  ;
  input \desIn[3]_pad  ;
  input \desIn[40]_pad  ;
  input \desIn[41]_pad  ;
  input \desIn[42]_pad  ;
  input \desIn[43]_pad  ;
  input \desIn[44]_pad  ;
  input \desIn[45]_pad  ;
  input \desIn[46]_pad  ;
  input \desIn[47]_pad  ;
  input \desIn[48]_pad  ;
  input \desIn[49]_pad  ;
  input \desIn[4]_pad  ;
  input \desIn[50]_pad  ;
  input \desIn[51]_pad  ;
  input \desIn[52]_pad  ;
  input \desIn[53]_pad  ;
  input \desIn[54]_pad  ;
  input \desIn[55]_pad  ;
  input \desIn[56]_pad  ;
  input \desIn[57]_pad  ;
  input \desIn[58]_pad  ;
  input \desIn[59]_pad  ;
  input \desIn[5]_pad  ;
  input \desIn[60]_pad  ;
  input \desIn[61]_pad  ;
  input \desIn[62]_pad  ;
  input \desIn[63]_pad  ;
  input \desIn[6]_pad  ;
  input \desIn[7]_pad  ;
  input \desIn[8]_pad  ;
  input \desIn[9]_pad  ;
  input \key1[0]_pad  ;
  input \key1[10]_pad  ;
  input \key1[11]_pad  ;
  input \key1[12]_pad  ;
  input \key1[13]_pad  ;
  input \key1[14]_pad  ;
  input \key1[15]_pad  ;
  input \key1[16]_pad  ;
  input \key1[17]_pad  ;
  input \key1[18]_pad  ;
  input \key1[19]_pad  ;
  input \key1[1]_pad  ;
  input \key1[20]_pad  ;
  input \key1[21]_pad  ;
  input \key1[22]_pad  ;
  input \key1[23]_pad  ;
  input \key1[24]_pad  ;
  input \key1[25]_pad  ;
  input \key1[26]_pad  ;
  input \key1[27]_pad  ;
  input \key1[28]_pad  ;
  input \key1[29]_pad  ;
  input \key1[2]_pad  ;
  input \key1[30]_pad  ;
  input \key1[31]_pad  ;
  input \key1[32]_pad  ;
  input \key1[33]_pad  ;
  input \key1[34]_pad  ;
  input \key1[35]_pad  ;
  input \key1[36]_pad  ;
  input \key1[37]_pad  ;
  input \key1[38]_pad  ;
  input \key1[39]_pad  ;
  input \key1[3]_pad  ;
  input \key1[40]_pad  ;
  input \key1[41]_pad  ;
  input \key1[42]_pad  ;
  input \key1[43]_pad  ;
  input \key1[44]_pad  ;
  input \key1[45]_pad  ;
  input \key1[46]_pad  ;
  input \key1[47]_pad  ;
  input \key1[48]_pad  ;
  input \key1[49]_pad  ;
  input \key1[4]_pad  ;
  input \key1[50]_pad  ;
  input \key1[51]_pad  ;
  input \key1[52]_pad  ;
  input \key1[53]_pad  ;
  input \key1[54]_pad  ;
  input \key1[55]_pad  ;
  input \key1[5]_pad  ;
  input \key1[6]_pad  ;
  input \key1[7]_pad  ;
  input \key1[8]_pad  ;
  input \key1[9]_pad  ;
  input \key2[0]_pad  ;
  input \key2[10]_pad  ;
  input \key2[11]_pad  ;
  input \key2[12]_pad  ;
  input \key2[13]_pad  ;
  input \key2[14]_pad  ;
  input \key2[15]_pad  ;
  input \key2[16]_pad  ;
  input \key2[17]_pad  ;
  input \key2[18]_pad  ;
  input \key2[19]_pad  ;
  input \key2[1]_pad  ;
  input \key2[20]_pad  ;
  input \key2[21]_pad  ;
  input \key2[22]_pad  ;
  input \key2[23]_pad  ;
  input \key2[24]_pad  ;
  input \key2[25]_pad  ;
  input \key2[26]_pad  ;
  input \key2[27]_pad  ;
  input \key2[28]_pad  ;
  input \key2[29]_pad  ;
  input \key2[2]_pad  ;
  input \key2[30]_pad  ;
  input \key2[31]_pad  ;
  input \key2[32]_pad  ;
  input \key2[33]_pad  ;
  input \key2[34]_pad  ;
  input \key2[35]_pad  ;
  input \key2[36]_pad  ;
  input \key2[37]_pad  ;
  input \key2[38]_pad  ;
  input \key2[39]_pad  ;
  input \key2[3]_pad  ;
  input \key2[40]_pad  ;
  input \key2[41]_pad  ;
  input \key2[42]_pad  ;
  input \key2[43]_pad  ;
  input \key2[44]_pad  ;
  input \key2[45]_pad  ;
  input \key2[46]_pad  ;
  input \key2[47]_pad  ;
  input \key2[48]_pad  ;
  input \key2[49]_pad  ;
  input \key2[4]_pad  ;
  input \key2[50]_pad  ;
  input \key2[51]_pad  ;
  input \key2[52]_pad  ;
  input \key2[53]_pad  ;
  input \key2[54]_pad  ;
  input \key2[55]_pad  ;
  input \key2[5]_pad  ;
  input \key2[6]_pad  ;
  input \key2[7]_pad  ;
  input \key2[8]_pad  ;
  input \key2[9]_pad  ;
  input \key3[0]_pad  ;
  input \key3[10]_pad  ;
  input \key3[11]_pad  ;
  input \key3[12]_pad  ;
  input \key3[13]_pad  ;
  input \key3[14]_pad  ;
  input \key3[15]_pad  ;
  input \key3[16]_pad  ;
  input \key3[17]_pad  ;
  input \key3[18]_pad  ;
  input \key3[19]_pad  ;
  input \key3[1]_pad  ;
  input \key3[20]_pad  ;
  input \key3[21]_pad  ;
  input \key3[22]_pad  ;
  input \key3[23]_pad  ;
  input \key3[24]_pad  ;
  input \key3[25]_pad  ;
  input \key3[26]_pad  ;
  input \key3[27]_pad  ;
  input \key3[28]_pad  ;
  input \key3[29]_pad  ;
  input \key3[2]_pad  ;
  input \key3[30]_pad  ;
  input \key3[31]_pad  ;
  input \key3[32]_pad  ;
  input \key3[33]_pad  ;
  input \key3[34]_pad  ;
  input \key3[35]_pad  ;
  input \key3[36]_pad  ;
  input \key3[37]_pad  ;
  input \key3[38]_pad  ;
  input \key3[39]_pad  ;
  input \key3[3]_pad  ;
  input \key3[40]_pad  ;
  input \key3[41]_pad  ;
  input \key3[42]_pad  ;
  input \key3[43]_pad  ;
  input \key3[44]_pad  ;
  input \key3[45]_pad  ;
  input \key3[46]_pad  ;
  input \key3[47]_pad  ;
  input \key3[48]_pad  ;
  input \key3[49]_pad  ;
  input \key3[4]_pad  ;
  input \key3[50]_pad  ;
  input \key3[51]_pad  ;
  input \key3[52]_pad  ;
  input \key3[53]_pad  ;
  input \key3[54]_pad  ;
  input \key3[55]_pad  ;
  input \key3[5]_pad  ;
  input \key3[6]_pad  ;
  input \key3[7]_pad  ;
  input \key3[8]_pad  ;
  input \key3[9]_pad  ;
  input \roundSel[0]_pad  ;
  input \roundSel[1]_pad  ;
  input \roundSel[2]_pad  ;
  input \roundSel[3]_pad  ;
  input \roundSel[4]_pad  ;
  input \roundSel[5]_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \desOut[0]_pad  ;
  output \desOut[11]_pad  ;
  output \desOut[12]_pad  ;
  output \desOut[13]_pad  ;
  output \desOut[14]_pad  ;
  output \desOut[15]_pad  ;
  output \desOut[18]_pad  ;
  output \desOut[1]_pad  ;
  output \desOut[22]_pad  ;
  output \desOut[23]_pad  ;
  output \desOut[24]_pad  ;
  output \desOut[25]_pad  ;
  output \desOut[26]_pad  ;
  output \desOut[28]_pad  ;
  output \desOut[2]_pad  ;
  output \desOut[30]_pad  ;
  output \desOut[32]_pad  ;
  output \desOut[34]_pad  ;
  output \desOut[35]_pad  ;
  output \desOut[37]_pad  ;
  output \desOut[38]_pad  ;
  output \desOut[39]_pad  ;
  output \desOut[3]_pad  ;
  output \desOut[40]_pad  ;
  output \desOut[42]_pad  ;
  output \desOut[44]_pad  ;
  output \desOut[45]_pad  ;
  output \desOut[46]_pad  ;
  output \desOut[48]_pad  ;
  output \desOut[4]_pad  ;
  output \desOut[50]_pad  ;
  output \desOut[52]_pad  ;
  output \desOut[54]_pad  ;
  output \desOut[56]_pad  ;
  output \desOut[57]_pad  ;
  output \desOut[59]_pad  ;
  output \desOut[5]_pad  ;
  output \desOut[60]_pad  ;
  output \desOut[61]_pad  ;
  output \desOut[63]_pad  ;
  output \desOut[6]_pad  ;
  output \desOut[8]_pad  ;
  output \desOut[9]_pad  ;
  output \g13525_dup/_0_  ;
  output \g13583_dup/_0_  ;
  output \g17813/_3_  ;
  output \g17816/_3_  ;
  output \g17819/_3_  ;
  output \g17822/_3_  ;
  output \g17836/_3_  ;
  output \g17871/_3_  ;
  output \g17878/_1_  ;
  output \g17881/_3_  ;
  output \g17966/_2_  ;
  output \g17969/_3_  ;
  output \g17996/_2_  ;
  output \g19574_dup/_3_  ;
  output \g19619_dup/_3_  ;
  output \g19756_dup/_3_  ;
  output \g20263/_3_  ;
  output \g20541/_2_  ;
  output \g20691/_1_  ;
  output \g20740_dup/_3_  ;
  output \g67/_2_  ;
  wire n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 ;
  assign n304 = ~\roundSel[0]_pad  & ~\roundSel[1]_pad  ;
  assign n305 = ~\roundSel[2]_pad  & ~\roundSel[3]_pad  ;
  assign n306 = n304 & n305 ;
  assign n307 = ~\roundSel[5]_pad  & n306 ;
  assign n308 = ~\roundSel[4]_pad  & n307 ;
  assign n309 = \desIn[27]_pad  & n308 ;
  assign n310 = ~\roundSel[4]_pad  & \roundSel[5]_pad  ;
  assign n311 = n306 & n310 ;
  assign n312 = \roundSel[4]_pad  & n307 ;
  assign n313 = ~n311 & ~n312 ;
  assign n315 = ~\FP_R_reg[20]/P0001  & n313 ;
  assign n314 = ~\FP_R_reg[52]/NET0131  & ~n313 ;
  assign n316 = ~n308 & ~n314 ;
  assign n317 = ~n315 & n316 ;
  assign n318 = ~n309 & ~n317 ;
  assign n343 = \roundSel[0]_pad  & ~\roundSel[1]_pad  ;
  assign n392 = n305 & n343 ;
  assign n319 = \roundSel[4]_pad  & ~\roundSel[5]_pad  ;
  assign n320 = decrypt_pad & ~n319 ;
  assign n321 = ~decrypt_pad & n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n324 = ~decrypt_pad & ~\roundSel[5]_pad  ;
  assign n325 = decrypt_pad & \roundSel[5]_pad  ;
  assign n326 = ~n324 & ~n325 ;
  assign n329 = ~\roundSel[4]_pad  & n326 ;
  assign n395 = \key3[30]_pad  & n329 ;
  assign n393 = \key2[30]_pad  & n319 ;
  assign n327 = ~\roundSel[4]_pad  & ~n326 ;
  assign n394 = \key1[30]_pad  & n327 ;
  assign n396 = ~n393 & ~n394 ;
  assign n397 = ~n395 & n396 ;
  assign n398 = n322 & ~n397 ;
  assign n401 = \key3[9]_pad  & n329 ;
  assign n399 = \key2[9]_pad  & n319 ;
  assign n400 = \key1[9]_pad  & n327 ;
  assign n402 = ~n399 & ~n400 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = ~n322 & ~n403 ;
  assign n405 = ~n398 & ~n404 ;
  assign n406 = n392 & ~n405 ;
  assign n376 = \roundSel[2]_pad  & ~\roundSel[3]_pad  ;
  assign n407 = ~\roundSel[0]_pad  & \roundSel[1]_pad  ;
  assign n408 = n376 & n407 ;
  assign n411 = \key3[49]_pad  & n329 ;
  assign n409 = \key2[49]_pad  & n319 ;
  assign n410 = \key1[49]_pad  & n327 ;
  assign n412 = ~n409 & ~n410 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n322 & ~n413 ;
  assign n417 = \key3[14]_pad  & n329 ;
  assign n415 = \key2[14]_pad  & n319 ;
  assign n416 = \key1[14]_pad  & n327 ;
  assign n418 = ~n415 & ~n416 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = n322 & ~n419 ;
  assign n421 = ~n414 & ~n420 ;
  assign n422 = n408 & ~n421 ;
  assign n495 = ~n406 & ~n422 ;
  assign n423 = n343 & n376 ;
  assign n426 = \key3[8]_pad  & n329 ;
  assign n424 = \key2[8]_pad  & n319 ;
  assign n425 = \key1[8]_pad  & n327 ;
  assign n427 = ~n424 & ~n425 ;
  assign n428 = ~n426 & n427 ;
  assign n429 = ~n322 & ~n428 ;
  assign n432 = \key3[0]_pad  & n329 ;
  assign n430 = \key2[0]_pad  & n319 ;
  assign n431 = \key1[0]_pad  & n327 ;
  assign n433 = ~n430 & ~n431 ;
  assign n434 = ~n432 & n433 ;
  assign n435 = n322 & ~n434 ;
  assign n436 = ~n429 & ~n435 ;
  assign n437 = n423 & ~n436 ;
  assign n438 = n304 & n376 ;
  assign n370 = \key3[45]_pad  & n329 ;
  assign n368 = \key2[45]_pad  & n319 ;
  assign n369 = \key1[45]_pad  & n327 ;
  assign n371 = ~n368 & ~n369 ;
  assign n372 = ~n370 & n371 ;
  assign n439 = n322 & ~n372 ;
  assign n364 = \key3[22]_pad  & n329 ;
  assign n362 = \key2[22]_pad  & n319 ;
  assign n363 = \key1[22]_pad  & n327 ;
  assign n365 = ~n362 & ~n363 ;
  assign n366 = ~n364 & n365 ;
  assign n440 = ~n322 & ~n366 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = n438 & ~n441 ;
  assign n496 = ~n437 & ~n442 ;
  assign n503 = n495 & n496 ;
  assign n330 = \key3[16]_pad  & n329 ;
  assign n323 = \key2[16]_pad  & n319 ;
  assign n328 = \key1[16]_pad  & n327 ;
  assign n331 = ~n323 & ~n328 ;
  assign n332 = ~n330 & n331 ;
  assign n333 = ~n322 & ~n332 ;
  assign n336 = \key3[23]_pad  & n329 ;
  assign n334 = \key2[23]_pad  & n319 ;
  assign n335 = \key1[23]_pad  & n327 ;
  assign n337 = ~n334 & ~n335 ;
  assign n338 = ~n336 & n337 ;
  assign n339 = n322 & ~n338 ;
  assign n340 = ~n333 & ~n339 ;
  assign n341 = n306 & ~n340 ;
  assign n342 = \roundSel[2]_pad  & \roundSel[3]_pad  ;
  assign n344 = n342 & n343 ;
  assign n347 = \key3[44]_pad  & n329 ;
  assign n345 = \key2[44]_pad  & n319 ;
  assign n346 = \key1[44]_pad  & n327 ;
  assign n348 = ~n345 & ~n346 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = ~n322 & ~n349 ;
  assign n353 = \key3[50]_pad  & n329 ;
  assign n351 = \key2[50]_pad  & n319 ;
  assign n352 = \key1[50]_pad  & n327 ;
  assign n354 = ~n351 & ~n352 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n322 & ~n355 ;
  assign n357 = ~n350 & ~n356 ;
  assign n358 = n344 & ~n357 ;
  assign n493 = ~n341 & ~n358 ;
  assign n359 = ~\roundSel[2]_pad  & \roundSel[3]_pad  ;
  assign n360 = \roundSel[0]_pad  & \roundSel[1]_pad  ;
  assign n361 = n359 & n360 ;
  assign n367 = n322 & ~n366 ;
  assign n373 = ~n322 & ~n372 ;
  assign n374 = ~n367 & ~n373 ;
  assign n375 = n361 & ~n374 ;
  assign n377 = n360 & n376 ;
  assign n380 = \key3[35]_pad  & n329 ;
  assign n378 = \key2[35]_pad  & n319 ;
  assign n379 = \key1[35]_pad  & n327 ;
  assign n381 = ~n378 & ~n379 ;
  assign n382 = ~n380 & n381 ;
  assign n383 = ~n322 & ~n382 ;
  assign n386 = \key3[28]_pad  & n329 ;
  assign n384 = \key2[28]_pad  & n319 ;
  assign n385 = \key1[28]_pad  & n327 ;
  assign n387 = ~n384 & ~n385 ;
  assign n388 = ~n386 & n387 ;
  assign n389 = n322 & ~n388 ;
  assign n390 = ~n383 & ~n389 ;
  assign n391 = n377 & ~n390 ;
  assign n494 = ~n375 & ~n391 ;
  assign n504 = n493 & n494 ;
  assign n505 = n503 & n504 ;
  assign n463 = n304 & n342 ;
  assign n466 = \key3[36]_pad  & n329 ;
  assign n464 = \key2[36]_pad  & n319 ;
  assign n465 = \key1[36]_pad  & n327 ;
  assign n467 = ~n464 & ~n465 ;
  assign n468 = ~n466 & n467 ;
  assign n469 = n322 & ~n468 ;
  assign n472 = \key3[31]_pad  & n329 ;
  assign n470 = \key2[31]_pad  & n319 ;
  assign n471 = \key1[31]_pad  & n327 ;
  assign n473 = ~n470 & ~n471 ;
  assign n474 = ~n472 & n473 ;
  assign n475 = ~n322 & ~n474 ;
  assign n476 = ~n469 & ~n475 ;
  assign n477 = n463 & ~n476 ;
  assign n478 = n342 & n407 ;
  assign n479 = ~n322 & ~n397 ;
  assign n480 = n322 & ~n403 ;
  assign n481 = ~n479 & ~n480 ;
  assign n482 = n478 & ~n481 ;
  assign n499 = ~n477 & ~n482 ;
  assign n483 = n342 & n360 ;
  assign n484 = n322 & ~n332 ;
  assign n485 = ~n322 & ~n338 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = n483 & ~n486 ;
  assign n488 = n305 & n360 ;
  assign n489 = n322 & ~n474 ;
  assign n490 = ~n322 & ~n468 ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = n488 & ~n491 ;
  assign n500 = ~n487 & ~n492 ;
  assign n501 = n499 & n500 ;
  assign n443 = n343 & n359 ;
  assign n444 = n322 & ~n413 ;
  assign n445 = ~n322 & ~n419 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n443 & ~n446 ;
  assign n448 = n305 & n407 ;
  assign n449 = n322 & ~n349 ;
  assign n450 = ~n322 & ~n355 ;
  assign n451 = ~n449 & ~n450 ;
  assign n452 = n448 & ~n451 ;
  assign n497 = ~n447 & ~n452 ;
  assign n453 = n304 & n359 ;
  assign n454 = n322 & ~n382 ;
  assign n455 = ~n322 & ~n388 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = n453 & ~n456 ;
  assign n458 = n359 & n407 ;
  assign n459 = n322 & ~n428 ;
  assign n460 = ~n322 & ~n434 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = n458 & ~n461 ;
  assign n498 = ~n457 & ~n462 ;
  assign n502 = n497 & n498 ;
  assign n506 = n501 & n502 ;
  assign n507 = n505 & n506 ;
  assign n508 = ~n318 & n507 ;
  assign n509 = n318 & ~n507 ;
  assign n510 = ~n508 & ~n509 ;
  assign n546 = \key3[51]_pad  & n329 ;
  assign n544 = \key2[51]_pad  & n319 ;
  assign n545 = \key1[51]_pad  & n327 ;
  assign n547 = ~n544 & ~n545 ;
  assign n548 = ~n546 & n547 ;
  assign n549 = n322 & ~n548 ;
  assign n550 = ~n475 & ~n549 ;
  assign n551 = n483 & ~n550 ;
  assign n552 = ~n322 & ~n548 ;
  assign n553 = ~n489 & ~n552 ;
  assign n554 = n306 & ~n553 ;
  assign n608 = ~n551 & ~n554 ;
  assign n530 = \key3[21]_pad  & n329 ;
  assign n528 = \key2[21]_pad  & n319 ;
  assign n529 = \key1[21]_pad  & n327 ;
  assign n531 = ~n528 & ~n529 ;
  assign n532 = ~n530 & n531 ;
  assign n555 = n322 & ~n532 ;
  assign n524 = \key3[2]_pad  & n329 ;
  assign n522 = \key2[2]_pad  & n319 ;
  assign n523 = \key1[2]_pad  & n327 ;
  assign n525 = ~n522 & ~n523 ;
  assign n526 = ~n524 & n525 ;
  assign n556 = ~n322 & ~n526 ;
  assign n557 = ~n555 & ~n556 ;
  assign n558 = n438 & ~n557 ;
  assign n561 = \key3[15]_pad  & n329 ;
  assign n559 = \key2[15]_pad  & n319 ;
  assign n560 = \key1[15]_pad  & n327 ;
  assign n562 = ~n559 & ~n560 ;
  assign n563 = ~n561 & n562 ;
  assign n564 = ~n322 & ~n563 ;
  assign n565 = ~n459 & ~n564 ;
  assign n566 = n377 & ~n565 ;
  assign n609 = ~n558 & ~n566 ;
  assign n616 = n608 & n609 ;
  assign n513 = \key3[29]_pad  & n329 ;
  assign n511 = \key2[29]_pad  & n319 ;
  assign n512 = \key1[29]_pad  & n327 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = ~n513 & n514 ;
  assign n516 = ~n322 & ~n515 ;
  assign n517 = ~n444 & ~n516 ;
  assign n518 = n408 & ~n517 ;
  assign n519 = n322 & ~n515 ;
  assign n520 = ~n414 & ~n519 ;
  assign n521 = n443 & ~n520 ;
  assign n606 = ~n518 & ~n521 ;
  assign n527 = n322 & ~n526 ;
  assign n533 = ~n322 & ~n532 ;
  assign n534 = ~n527 & ~n533 ;
  assign n535 = n361 & ~n534 ;
  assign n538 = \key3[7]_pad  & n329 ;
  assign n536 = \key2[7]_pad  & n319 ;
  assign n537 = \key1[7]_pad  & n327 ;
  assign n539 = ~n536 & ~n537 ;
  assign n540 = ~n538 & n539 ;
  assign n541 = ~n322 & ~n540 ;
  assign n542 = ~n484 & ~n541 ;
  assign n543 = n463 & ~n542 ;
  assign n607 = ~n535 & ~n543 ;
  assign n617 = n606 & n607 ;
  assign n618 = n616 & n617 ;
  assign n591 = \key3[38]_pad  & n329 ;
  assign n589 = \key2[38]_pad  & n319 ;
  assign n590 = \key1[38]_pad  & n327 ;
  assign n592 = ~n589 & ~n590 ;
  assign n593 = ~n591 & n592 ;
  assign n594 = ~n322 & ~n593 ;
  assign n595 = ~n449 & ~n594 ;
  assign n596 = n478 & ~n595 ;
  assign n597 = n322 & ~n593 ;
  assign n598 = ~n350 & ~n597 ;
  assign n599 = n392 & ~n598 ;
  assign n612 = ~n596 & ~n599 ;
  assign n583 = \key3[43]_pad  & n329 ;
  assign n581 = \key2[43]_pad  & n319 ;
  assign n582 = \key1[43]_pad  & n327 ;
  assign n584 = ~n581 & ~n582 ;
  assign n585 = ~n583 & n584 ;
  assign n600 = ~n322 & ~n585 ;
  assign n601 = ~n454 & ~n600 ;
  assign n602 = n423 & ~n601 ;
  assign n603 = n322 & ~n563 ;
  assign n604 = ~n429 & ~n603 ;
  assign n605 = n453 & ~n604 ;
  assign n613 = ~n602 & ~n605 ;
  assign n614 = n612 & n613 ;
  assign n567 = n322 & ~n540 ;
  assign n568 = ~n333 & ~n567 ;
  assign n569 = n488 & ~n568 ;
  assign n572 = \key3[52]_pad  & n329 ;
  assign n570 = \key2[52]_pad  & n319 ;
  assign n571 = \key1[52]_pad  & n327 ;
  assign n573 = ~n570 & ~n571 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = n322 & ~n574 ;
  assign n576 = ~n479 & ~n575 ;
  assign n577 = n448 & ~n576 ;
  assign n610 = ~n569 & ~n577 ;
  assign n578 = ~n322 & ~n574 ;
  assign n579 = ~n398 & ~n578 ;
  assign n580 = n344 & ~n579 ;
  assign n586 = n322 & ~n585 ;
  assign n587 = ~n383 & ~n586 ;
  assign n588 = n458 & ~n587 ;
  assign n611 = ~n580 & ~n588 ;
  assign n615 = n610 & n611 ;
  assign n619 = n614 & n615 ;
  assign n620 = n618 & n619 ;
  assign n621 = \desIn[3]_pad  & n308 ;
  assign n623 = ~\FP_R_reg[17]/P0001  & n313 ;
  assign n622 = ~\FP_R_reg[49]/NET0131  & ~n313 ;
  assign n624 = ~n308 & ~n622 ;
  assign n625 = ~n623 & n624 ;
  assign n626 = ~n621 & ~n625 ;
  assign n627 = n620 & ~n626 ;
  assign n628 = ~n620 & n626 ;
  assign n629 = ~n627 & ~n628 ;
  assign n638 = ~n429 & ~n527 ;
  assign n639 = n448 & ~n638 ;
  assign n640 = ~n373 & ~n575 ;
  assign n641 = n453 & ~n640 ;
  assign n664 = ~n639 & ~n641 ;
  assign n642 = ~n440 & ~n586 ;
  assign n643 = n392 & ~n642 ;
  assign n644 = ~n454 & ~n479 ;
  assign n645 = n361 & ~n644 ;
  assign n665 = ~n643 & ~n645 ;
  assign n672 = n664 & n665 ;
  assign n630 = ~n333 & ~n444 ;
  assign n631 = n463 & ~n630 ;
  assign n632 = ~n439 & ~n578 ;
  assign n633 = n377 & ~n632 ;
  assign n662 = ~n631 & ~n633 ;
  assign n634 = ~n367 & ~n600 ;
  assign n635 = n478 & ~n634 ;
  assign n636 = ~n489 & ~n541 ;
  assign n637 = n408 & ~n636 ;
  assign n663 = ~n635 & ~n637 ;
  assign n673 = n662 & n663 ;
  assign n674 = n672 & n673 ;
  assign n654 = ~n475 & ~n567 ;
  assign n655 = n443 & ~n654 ;
  assign n656 = ~n490 & ~n519 ;
  assign n657 = n483 & ~n656 ;
  assign n668 = ~n655 & ~n657 ;
  assign n658 = ~n350 & ~n555 ;
  assign n659 = n458 & ~n658 ;
  assign n660 = ~n383 & ~n398 ;
  assign n661 = n438 & ~n660 ;
  assign n669 = ~n659 & ~n661 ;
  assign n670 = n668 & n669 ;
  assign n646 = ~n414 & ~n484 ;
  assign n647 = n488 & ~n646 ;
  assign n648 = ~n469 & ~n516 ;
  assign n649 = n306 & ~n648 ;
  assign n666 = ~n647 & ~n649 ;
  assign n650 = ~n459 & ~n556 ;
  assign n651 = n344 & ~n650 ;
  assign n652 = ~n449 & ~n533 ;
  assign n653 = n423 & ~n652 ;
  assign n667 = ~n651 & ~n653 ;
  assign n671 = n666 & n667 ;
  assign n675 = n670 & n671 ;
  assign n676 = n674 & n675 ;
  assign n677 = \desIn[61]_pad  & n308 ;
  assign n679 = ~\FP_R_reg[16]/P0001  & n313 ;
  assign n678 = ~\FP_R_reg[48]/NET0131  & ~n313 ;
  assign n680 = ~n308 & ~n678 ;
  assign n681 = ~n679 & n680 ;
  assign n682 = ~n677 & ~n681 ;
  assign n683 = n676 & ~n682 ;
  assign n684 = ~n676 & n682 ;
  assign n685 = ~n683 & ~n684 ;
  assign n699 = ~n445 & ~n549 ;
  assign n700 = n344 & ~n699 ;
  assign n701 = n306 & ~n640 ;
  assign n737 = ~n700 & ~n701 ;
  assign n702 = ~n450 & ~n603 ;
  assign n703 = n408 & ~n702 ;
  assign n704 = ~n356 & ~n564 ;
  assign n705 = n443 & ~n704 ;
  assign n738 = ~n703 & ~n705 ;
  assign n745 = n737 & n738 ;
  assign n686 = ~n460 & ~n597 ;
  assign n687 = n478 & ~n686 ;
  assign n688 = n453 & ~n648 ;
  assign n735 = ~n687 & ~n688 ;
  assign n691 = \key3[42]_pad  & n329 ;
  assign n689 = \key2[42]_pad  & n319 ;
  assign n690 = \key1[42]_pad  & n327 ;
  assign n692 = ~n689 & ~n690 ;
  assign n693 = ~n691 & n692 ;
  assign n694 = ~n322 & ~n693 ;
  assign n695 = ~n339 & ~n694 ;
  assign n696 = n361 & ~n695 ;
  assign n697 = ~n420 & ~n552 ;
  assign n698 = n448 & ~n697 ;
  assign n736 = ~n696 & ~n698 ;
  assign n746 = n735 & n736 ;
  assign n747 = n745 & n746 ;
  assign n726 = ~n435 & ~n594 ;
  assign n727 = n392 & ~n726 ;
  assign n728 = n377 & ~n656 ;
  assign n741 = ~n727 & ~n728 ;
  assign n708 = \key3[37]_pad  & n329 ;
  assign n706 = \key2[37]_pad  & n319 ;
  assign n707 = \key1[37]_pad  & n327 ;
  assign n709 = ~n706 & ~n707 ;
  assign n710 = ~n708 & n709 ;
  assign n729 = ~n322 & ~n710 ;
  assign n730 = ~n389 & ~n729 ;
  assign n731 = n488 & ~n730 ;
  assign n720 = \key3[1]_pad  & n329 ;
  assign n718 = \key2[1]_pad  & n319 ;
  assign n719 = \key1[1]_pad  & n327 ;
  assign n721 = ~n718 & ~n719 ;
  assign n722 = ~n720 & n721 ;
  assign n732 = n322 & ~n722 ;
  assign n733 = ~n404 & ~n732 ;
  assign n734 = n423 & ~n733 ;
  assign n742 = ~n731 & ~n734 ;
  assign n743 = n741 & n742 ;
  assign n711 = n322 & ~n710 ;
  assign n712 = ~n455 & ~n711 ;
  assign n713 = n463 & ~n712 ;
  assign n714 = n483 & ~n632 ;
  assign n739 = ~n713 & ~n714 ;
  assign n715 = n322 & ~n693 ;
  assign n716 = ~n485 & ~n715 ;
  assign n717 = n438 & ~n716 ;
  assign n723 = ~n322 & ~n722 ;
  assign n724 = ~n480 & ~n723 ;
  assign n725 = n458 & ~n724 ;
  assign n740 = ~n717 & ~n725 ;
  assign n744 = n739 & n740 ;
  assign n748 = n743 & n744 ;
  assign n749 = n747 & n748 ;
  assign n750 = \desIn[35]_pad  & n308 ;
  assign n752 = ~\FP_R_reg[21]/P0001  & n313 ;
  assign n751 = ~\FP_R_reg[53]/NET0131  & ~n313 ;
  assign n753 = ~n308 & ~n751 ;
  assign n754 = ~n752 & n753 ;
  assign n755 = ~n750 & ~n754 ;
  assign n756 = n749 & ~n755 ;
  assign n757 = ~n749 & n755 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = n685 & n758 ;
  assign n760 = n629 & n759 ;
  assign n769 = ~n527 & ~n541 ;
  assign n770 = n438 & ~n769 ;
  assign n771 = ~n350 & ~n549 ;
  assign n772 = n453 & ~n771 ;
  assign n795 = ~n770 & ~n772 ;
  assign n773 = ~n429 & ~n732 ;
  assign n774 = n483 & ~n773 ;
  assign n775 = ~n414 & ~n603 ;
  assign n776 = n392 & ~n775 ;
  assign n796 = ~n774 & ~n776 ;
  assign n803 = n795 & n796 ;
  assign n761 = ~n555 & ~n600 ;
  assign n762 = n463 & ~n761 ;
  assign n763 = ~n459 & ~n723 ;
  assign n764 = n306 & ~n763 ;
  assign n793 = ~n762 & ~n764 ;
  assign n765 = ~n383 & ~n519 ;
  assign n766 = n448 & ~n765 ;
  assign n767 = ~n398 & ~n594 ;
  assign n768 = n408 & ~n767 ;
  assign n794 = ~n766 & ~n768 ;
  assign n804 = n793 & n794 ;
  assign n805 = n803 & n804 ;
  assign n785 = ~n333 & ~n575 ;
  assign n786 = n458 & ~n785 ;
  assign n787 = ~n449 & ~n552 ;
  assign n788 = n377 & ~n787 ;
  assign n799 = ~n786 & ~n788 ;
  assign n789 = ~n454 & ~n516 ;
  assign n790 = n344 & ~n789 ;
  assign n791 = ~n533 & ~n586 ;
  assign n792 = n488 & ~n791 ;
  assign n800 = ~n790 & ~n792 ;
  assign n801 = n799 & n800 ;
  assign n777 = ~n479 & ~n597 ;
  assign n778 = n443 & ~n777 ;
  assign n779 = ~n444 & ~n564 ;
  assign n780 = n478 & ~n779 ;
  assign n797 = ~n778 & ~n780 ;
  assign n781 = ~n484 & ~n578 ;
  assign n782 = n423 & ~n781 ;
  assign n783 = ~n556 & ~n567 ;
  assign n784 = n361 & ~n783 ;
  assign n798 = ~n782 & ~n784 ;
  assign n802 = n797 & n798 ;
  assign n806 = n801 & n802 ;
  assign n807 = n805 & n806 ;
  assign n808 = ~\desIn[19]_pad  & n308 ;
  assign n810 = \FP_R_reg[51]/NET0131  & ~n313 ;
  assign n809 = \FP_R_reg[19]/P0001  & n313 ;
  assign n811 = ~n308 & ~n809 ;
  assign n812 = ~n810 & n811 ;
  assign n813 = ~n808 & ~n812 ;
  assign n814 = n807 & ~n813 ;
  assign n815 = ~n807 & n813 ;
  assign n816 = ~n814 & ~n815 ;
  assign n817 = ~n629 & ~n685 ;
  assign n878 = ~n816 & ~n817 ;
  assign n879 = ~n760 & n878 ;
  assign n826 = ~n339 & ~n600 ;
  assign n827 = n443 & ~n826 ;
  assign n828 = ~n420 & ~n533 ;
  assign n829 = n483 & ~n828 ;
  assign n852 = ~n827 & ~n829 ;
  assign n830 = ~n445 & ~n555 ;
  assign n831 = n306 & ~n830 ;
  assign n832 = ~n485 & ~n586 ;
  assign n833 = n408 & ~n832 ;
  assign n853 = ~n831 & ~n833 ;
  assign n860 = n852 & n853 ;
  assign n818 = ~n519 & ~n729 ;
  assign n819 = n423 & ~n818 ;
  assign n820 = ~n480 & ~n556 ;
  assign n821 = n453 & ~n820 ;
  assign n850 = ~n819 & ~n821 ;
  assign n822 = ~n597 & ~n723 ;
  assign n823 = n463 & ~n822 ;
  assign n824 = ~n455 & ~n567 ;
  assign n825 = n478 & ~n824 ;
  assign n851 = ~n823 & ~n825 ;
  assign n861 = n850 & n851 ;
  assign n862 = n860 & n861 ;
  assign n842 = ~n516 & ~n711 ;
  assign n843 = n458 & ~n842 ;
  assign n844 = ~n404 & ~n527 ;
  assign n845 = n377 & ~n844 ;
  assign n856 = ~n843 & ~n845 ;
  assign n846 = ~n594 & ~n732 ;
  assign n847 = n488 & ~n846 ;
  assign n848 = ~n549 & ~n564 ;
  assign n849 = n361 & ~n848 ;
  assign n857 = ~n847 & ~n849 ;
  assign n858 = n856 & n857 ;
  assign n834 = ~n578 & ~n715 ;
  assign n835 = n448 & ~n834 ;
  assign n836 = ~n389 & ~n541 ;
  assign n837 = n392 & ~n836 ;
  assign n854 = ~n835 & ~n837 ;
  assign n838 = ~n575 & ~n694 ;
  assign n839 = n344 & ~n838 ;
  assign n840 = ~n552 & ~n603 ;
  assign n841 = n438 & ~n840 ;
  assign n855 = ~n839 & ~n841 ;
  assign n859 = n854 & n855 ;
  assign n863 = n858 & n859 ;
  assign n864 = n862 & n863 ;
  assign n865 = \desIn[11]_pad  & n308 ;
  assign n867 = ~\FP_R_reg[18]/P0001  & n313 ;
  assign n866 = ~\FP_R_reg[50]/NET0131  & ~n313 ;
  assign n868 = ~n308 & ~n866 ;
  assign n869 = ~n867 & n868 ;
  assign n870 = ~n865 & ~n869 ;
  assign n871 = ~n864 & n870 ;
  assign n872 = n864 & ~n870 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = ~n685 & ~n758 ;
  assign n875 = n873 & n874 ;
  assign n876 = ~n629 & ~n758 ;
  assign n877 = ~n873 & n876 ;
  assign n880 = ~n875 & ~n877 ;
  assign n881 = n879 & n880 ;
  assign n884 = ~n629 & n759 ;
  assign n882 = n629 & ~n873 ;
  assign n883 = ~n685 & n882 ;
  assign n885 = n816 & ~n883 ;
  assign n886 = ~n884 & n885 ;
  assign n887 = ~n881 & ~n886 ;
  assign n888 = n685 & ~n758 ;
  assign n889 = n629 & n888 ;
  assign n890 = n873 & n889 ;
  assign n891 = n758 & ~n873 ;
  assign n892 = n629 & n891 ;
  assign n893 = ~n890 & ~n892 ;
  assign n894 = ~n887 & n893 ;
  assign n895 = n510 & ~n894 ;
  assign n896 = ~n629 & n875 ;
  assign n897 = ~n890 & ~n896 ;
  assign n898 = ~n685 & n891 ;
  assign n899 = ~n629 & n898 ;
  assign n900 = n897 & ~n899 ;
  assign n901 = ~n816 & ~n900 ;
  assign n916 = n685 & ~n876 ;
  assign n909 = n816 & ~n817 ;
  assign n917 = ~n510 & ~n882 ;
  assign n918 = n909 & n917 ;
  assign n919 = ~n916 & n918 ;
  assign n907 = n629 & ~n758 ;
  assign n908 = ~n816 & ~n907 ;
  assign n910 = ~n510 & ~n873 ;
  assign n911 = ~n908 & n910 ;
  assign n912 = ~n909 & n911 ;
  assign n903 = ~n685 & n758 ;
  assign n904 = n629 & n903 ;
  assign n905 = ~n510 & n873 ;
  assign n906 = n904 & n905 ;
  assign n902 = n759 & n882 ;
  assign n913 = ~n629 & n873 ;
  assign n914 = n685 & n816 ;
  assign n915 = n913 & n914 ;
  assign n920 = ~n902 & ~n915 ;
  assign n921 = ~n906 & n920 ;
  assign n922 = ~n912 & n921 ;
  assign n923 = ~n919 & n922 ;
  assign n924 = ~n901 & n923 ;
  assign n925 = ~n895 & n924 ;
  assign n926 = ~\desIn[0]_pad  & n308 ;
  assign n928 = \FP_R_reg[25]/P0001  & ~n313 ;
  assign n927 = \FP_R_reg[57]/NET0131  & n313 ;
  assign n929 = ~n308 & ~n927 ;
  assign n930 = ~n928 & n929 ;
  assign n931 = ~n926 & ~n930 ;
  assign n932 = n925 & ~n931 ;
  assign n933 = ~n925 & n931 ;
  assign n934 = ~n932 & ~n933 ;
  assign n993 = \key3[4]_pad  & n329 ;
  assign n991 = \key2[4]_pad  & n319 ;
  assign n992 = \key1[4]_pad  & n327 ;
  assign n994 = ~n991 & ~n992 ;
  assign n995 = ~n993 & n994 ;
  assign n996 = n322 & ~n995 ;
  assign n999 = \key3[12]_pad  & n329 ;
  assign n997 = \key2[12]_pad  & n319 ;
  assign n998 = \key1[12]_pad  & n327 ;
  assign n1000 = ~n997 & ~n998 ;
  assign n1001 = ~n999 & n1000 ;
  assign n1002 = ~n322 & ~n1001 ;
  assign n1003 = ~n996 & ~n1002 ;
  assign n1004 = n448 & ~n1003 ;
  assign n1005 = ~n322 & ~n995 ;
  assign n1006 = n322 & ~n1001 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = n344 & ~n1007 ;
  assign n1081 = ~n1004 & ~n1008 ;
  assign n951 = \key3[27]_pad  & n329 ;
  assign n949 = \key2[27]_pad  & n319 ;
  assign n950 = \key1[27]_pad  & n327 ;
  assign n952 = ~n949 & ~n950 ;
  assign n953 = ~n951 & n952 ;
  assign n1009 = ~n322 & ~n953 ;
  assign n957 = \key3[46]_pad  & n329 ;
  assign n955 = \key2[46]_pad  & n319 ;
  assign n956 = \key1[46]_pad  & n327 ;
  assign n958 = ~n955 & ~n956 ;
  assign n959 = ~n957 & n958 ;
  assign n1010 = n322 & ~n959 ;
  assign n1011 = ~n1009 & ~n1010 ;
  assign n1012 = n423 & ~n1011 ;
  assign n1015 = \key3[33]_pad  & n329 ;
  assign n1013 = \key2[33]_pad  & n319 ;
  assign n1014 = \key1[33]_pad  & n327 ;
  assign n1016 = ~n1013 & ~n1014 ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1018 = n322 & ~n1017 ;
  assign n1021 = \key3[40]_pad  & n329 ;
  assign n1019 = \key2[40]_pad  & n319 ;
  assign n1020 = \key1[40]_pad  & n327 ;
  assign n1022 = ~n1019 & ~n1020 ;
  assign n1023 = ~n1021 & n1022 ;
  assign n1024 = ~n322 & ~n1023 ;
  assign n1025 = ~n1018 & ~n1024 ;
  assign n1026 = n483 & ~n1025 ;
  assign n1082 = ~n1012 & ~n1026 ;
  assign n1089 = n1081 & n1082 ;
  assign n937 = \key3[24]_pad  & n329 ;
  assign n935 = \key2[24]_pad  & n319 ;
  assign n936 = \key1[24]_pad  & n327 ;
  assign n938 = ~n935 & ~n936 ;
  assign n939 = ~n937 & n938 ;
  assign n940 = n322 & ~n939 ;
  assign n943 = \key3[17]_pad  & n329 ;
  assign n941 = \key2[17]_pad  & n319 ;
  assign n942 = \key1[17]_pad  & n327 ;
  assign n944 = ~n941 & ~n942 ;
  assign n945 = ~n943 & n944 ;
  assign n946 = ~n322 & ~n945 ;
  assign n947 = ~n940 & ~n946 ;
  assign n948 = n453 & ~n947 ;
  assign n954 = n322 & ~n953 ;
  assign n960 = ~n322 & ~n959 ;
  assign n961 = ~n954 & ~n960 ;
  assign n962 = n458 & ~n961 ;
  assign n1079 = ~n948 & ~n962 ;
  assign n965 = \key3[47]_pad  & n329 ;
  assign n963 = \key2[47]_pad  & n319 ;
  assign n964 = \key1[47]_pad  & n327 ;
  assign n966 = ~n963 & ~n964 ;
  assign n967 = ~n965 & n966 ;
  assign n968 = ~n322 & ~n967 ;
  assign n971 = \key3[26]_pad  & n329 ;
  assign n969 = \key2[26]_pad  & n319 ;
  assign n970 = \key1[26]_pad  & n327 ;
  assign n972 = ~n969 & ~n970 ;
  assign n973 = ~n971 & n972 ;
  assign n974 = n322 & ~n973 ;
  assign n975 = ~n968 & ~n974 ;
  assign n976 = n478 & ~n975 ;
  assign n979 = \key3[32]_pad  & n329 ;
  assign n977 = \key2[32]_pad  & n319 ;
  assign n978 = \key1[32]_pad  & n327 ;
  assign n980 = ~n977 & ~n978 ;
  assign n981 = ~n979 & n980 ;
  assign n982 = ~n322 & ~n981 ;
  assign n985 = \key3[41]_pad  & n329 ;
  assign n983 = \key2[41]_pad  & n319 ;
  assign n984 = \key1[41]_pad  & n327 ;
  assign n986 = ~n983 & ~n984 ;
  assign n987 = ~n985 & n986 ;
  assign n988 = n322 & ~n987 ;
  assign n989 = ~n982 & ~n988 ;
  assign n990 = n361 & ~n989 ;
  assign n1080 = ~n976 & ~n990 ;
  assign n1090 = n1079 & n1080 ;
  assign n1091 = n1089 & n1090 ;
  assign n1063 = ~n322 & ~n939 ;
  assign n1064 = n322 & ~n945 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = n377 & ~n1065 ;
  assign n1043 = \key3[13]_pad  & n329 ;
  assign n1041 = \key2[13]_pad  & n319 ;
  assign n1042 = \key1[13]_pad  & n327 ;
  assign n1044 = ~n1041 & ~n1042 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1067 = n322 & ~n1045 ;
  assign n1049 = \key3[3]_pad  & n329 ;
  assign n1047 = \key2[3]_pad  & n319 ;
  assign n1048 = \key1[3]_pad  & n327 ;
  assign n1050 = ~n1047 & ~n1048 ;
  assign n1051 = ~n1049 & n1050 ;
  assign n1068 = ~n322 & ~n1051 ;
  assign n1069 = ~n1067 & ~n1068 ;
  assign n1070 = n443 & ~n1069 ;
  assign n1085 = ~n1066 & ~n1070 ;
  assign n1071 = ~n322 & ~n1017 ;
  assign n1072 = n322 & ~n1023 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1074 = n306 & ~n1073 ;
  assign n1075 = n322 & ~n967 ;
  assign n1076 = ~n322 & ~n973 ;
  assign n1077 = ~n1075 & ~n1076 ;
  assign n1078 = n392 & ~n1077 ;
  assign n1086 = ~n1074 & ~n1078 ;
  assign n1087 = n1085 & n1086 ;
  assign n1029 = \key3[18]_pad  & n329 ;
  assign n1027 = \key2[18]_pad  & n319 ;
  assign n1028 = \key1[18]_pad  & n327 ;
  assign n1030 = ~n1027 & ~n1028 ;
  assign n1031 = ~n1029 & n1030 ;
  assign n1032 = ~n322 & ~n1031 ;
  assign n1035 = \key3[55]_pad  & n329 ;
  assign n1033 = \key2[55]_pad  & n319 ;
  assign n1034 = \key1[55]_pad  & n327 ;
  assign n1036 = ~n1033 & ~n1034 ;
  assign n1037 = ~n1035 & n1036 ;
  assign n1038 = n322 & ~n1037 ;
  assign n1039 = ~n1032 & ~n1038 ;
  assign n1040 = n463 & ~n1039 ;
  assign n1046 = ~n322 & ~n1045 ;
  assign n1052 = n322 & ~n1051 ;
  assign n1053 = ~n1046 & ~n1052 ;
  assign n1054 = n408 & ~n1053 ;
  assign n1083 = ~n1040 & ~n1054 ;
  assign n1055 = n322 & ~n1031 ;
  assign n1056 = ~n322 & ~n1037 ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = n488 & ~n1057 ;
  assign n1059 = n322 & ~n981 ;
  assign n1060 = ~n322 & ~n987 ;
  assign n1061 = ~n1059 & ~n1060 ;
  assign n1062 = n438 & ~n1061 ;
  assign n1084 = ~n1058 & ~n1062 ;
  assign n1088 = n1083 & n1084 ;
  assign n1092 = n1087 & n1088 ;
  assign n1093 = n1091 & n1092 ;
  assign n1094 = n682 & ~n1093 ;
  assign n1095 = ~n682 & n1093 ;
  assign n1096 = ~n1094 & ~n1095 ;
  assign n1126 = \key3[53]_pad  & n329 ;
  assign n1124 = \key2[53]_pad  & n319 ;
  assign n1125 = \key1[53]_pad  & n327 ;
  assign n1127 = ~n1124 & ~n1125 ;
  assign n1128 = ~n1126 & n1127 ;
  assign n1129 = n322 & ~n1128 ;
  assign n1240 = ~n1032 & ~n1129 ;
  assign n1241 = n443 & ~n1240 ;
  assign n1185 = \key3[39]_pad  & n329 ;
  assign n1183 = \key2[39]_pad  & n319 ;
  assign n1184 = \key1[39]_pad  & n327 ;
  assign n1186 = ~n1183 & ~n1184 ;
  assign n1187 = ~n1185 & n1186 ;
  assign n1202 = ~n322 & ~n1187 ;
  assign n1242 = ~n1059 & ~n1202 ;
  assign n1243 = n377 & ~n1242 ;
  assign n1266 = ~n1241 & ~n1243 ;
  assign n1198 = ~n322 & ~n1128 ;
  assign n1244 = ~n1055 & ~n1198 ;
  assign n1245 = n408 & ~n1244 ;
  assign n1179 = \key3[19]_pad  & n329 ;
  assign n1177 = \key2[19]_pad  & n319 ;
  assign n1178 = \key1[19]_pad  & n327 ;
  assign n1180 = ~n1177 & ~n1178 ;
  assign n1181 = ~n1179 & n1180 ;
  assign n1182 = ~n322 & ~n1181 ;
  assign n1246 = ~n954 & ~n1182 ;
  assign n1247 = n344 & ~n1246 ;
  assign n1267 = ~n1245 & ~n1247 ;
  assign n1274 = n1266 & n1267 ;
  assign n1232 = ~n1063 & ~n1075 ;
  assign n1233 = n438 & ~n1232 ;
  assign n1157 = \key3[48]_pad  & n329 ;
  assign n1155 = \key2[48]_pad  & n319 ;
  assign n1156 = \key1[48]_pad  & n327 ;
  assign n1158 = ~n1155 & ~n1156 ;
  assign n1159 = ~n1157 & n1158 ;
  assign n1160 = ~n322 & ~n1159 ;
  assign n1234 = ~n1038 & ~n1160 ;
  assign n1235 = n306 & ~n1234 ;
  assign n1264 = ~n1233 & ~n1235 ;
  assign n1191 = n322 & ~n1159 ;
  assign n1236 = ~n1056 & ~n1191 ;
  assign n1237 = n483 & ~n1236 ;
  assign n1163 = \key3[10]_pad  & n329 ;
  assign n1161 = \key2[10]_pad  & n319 ;
  assign n1162 = \key1[10]_pad  & n327 ;
  assign n1164 = ~n1161 & ~n1162 ;
  assign n1165 = ~n1163 & n1164 ;
  assign n1166 = n322 & ~n1165 ;
  assign n1238 = ~n1005 & ~n1166 ;
  assign n1239 = n458 & ~n1238 ;
  assign n1265 = ~n1237 & ~n1239 ;
  assign n1275 = n1264 & n1265 ;
  assign n1276 = n1274 & n1275 ;
  assign n1256 = ~n1018 & ~n1046 ;
  assign n1257 = n488 & ~n1256 ;
  assign n1188 = n322 & ~n1187 ;
  assign n1258 = ~n982 & ~n1188 ;
  assign n1259 = n453 & ~n1258 ;
  assign n1270 = ~n1257 & ~n1259 ;
  assign n1132 = \key3[5]_pad  & n329 ;
  assign n1130 = \key2[5]_pad  & n319 ;
  assign n1131 = \key1[5]_pad  & n327 ;
  assign n1133 = ~n1130 & ~n1131 ;
  assign n1134 = ~n1132 & n1133 ;
  assign n1135 = ~n322 & ~n1134 ;
  assign n1260 = ~n988 & ~n1135 ;
  assign n1261 = n478 & ~n1260 ;
  assign n1262 = ~n1067 & ~n1071 ;
  assign n1263 = n463 & ~n1262 ;
  assign n1271 = ~n1261 & ~n1263 ;
  assign n1272 = n1270 & n1271 ;
  assign n1199 = n322 & ~n1134 ;
  assign n1248 = ~n1060 & ~n1199 ;
  assign n1249 = n392 & ~n1248 ;
  assign n1250 = ~n940 & ~n968 ;
  assign n1251 = n361 & ~n1250 ;
  assign n1268 = ~n1249 & ~n1251 ;
  assign n1192 = ~n322 & ~n1165 ;
  assign n1252 = ~n996 & ~n1192 ;
  assign n1253 = n423 & ~n1252 ;
  assign n1203 = n322 & ~n1181 ;
  assign n1254 = ~n1009 & ~n1203 ;
  assign n1255 = n448 & ~n1254 ;
  assign n1269 = ~n1253 & ~n1255 ;
  assign n1273 = n1268 & n1269 ;
  assign n1277 = n1272 & n1273 ;
  assign n1278 = n1276 & n1277 ;
  assign n1279 = \desIn[37]_pad  & n308 ;
  assign n1281 = ~\FP_R_reg[13]/P0001  & n313 ;
  assign n1280 = ~\FP_R_reg[45]/NET0131  & ~n313 ;
  assign n1282 = ~n308 & ~n1280 ;
  assign n1283 = ~n1281 & n1282 ;
  assign n1284 = ~n1279 & ~n1283 ;
  assign n1285 = n1278 & ~n1284 ;
  assign n1286 = ~n1278 & n1284 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1107 = \key3[20]_pad  & n329 ;
  assign n1105 = \key2[20]_pad  & n319 ;
  assign n1106 = \key1[20]_pad  & n327 ;
  assign n1108 = ~n1105 & ~n1106 ;
  assign n1109 = ~n1107 & n1108 ;
  assign n1110 = ~n322 & ~n1109 ;
  assign n1302 = ~n1110 & ~n1129 ;
  assign n1303 = n344 & ~n1302 ;
  assign n1304 = n377 & ~n1025 ;
  assign n1325 = ~n1303 & ~n1304 ;
  assign n1305 = n483 & ~n1065 ;
  assign n1296 = \key3[6]_pad  & n329 ;
  assign n1294 = \key2[6]_pad  & n319 ;
  assign n1295 = \key1[6]_pad  & n327 ;
  assign n1297 = ~n1294 & ~n1295 ;
  assign n1298 = ~n1296 & n1297 ;
  assign n1306 = ~n322 & ~n1298 ;
  assign n1307 = ~n1166 & ~n1306 ;
  assign n1308 = n478 & ~n1307 ;
  assign n1326 = ~n1305 & ~n1308 ;
  assign n1333 = n1325 & n1326 ;
  assign n1171 = \key3[11]_pad  & n329 ;
  assign n1169 = \key2[11]_pad  & n319 ;
  assign n1170 = \key1[11]_pad  & n327 ;
  assign n1172 = ~n1169 & ~n1170 ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1195 = ~n322 & ~n1173 ;
  assign n1288 = ~n1195 & ~n1199 ;
  assign n1289 = n423 & ~n1288 ;
  assign n1143 = \key3[34]_pad  & n329 ;
  assign n1141 = \key2[34]_pad  & n319 ;
  assign n1142 = \key1[34]_pad  & n327 ;
  assign n1144 = ~n1141 & ~n1142 ;
  assign n1145 = ~n1143 & n1144 ;
  assign n1146 = n322 & ~n1145 ;
  assign n1290 = ~n1146 & ~n1202 ;
  assign n1291 = n488 & ~n1290 ;
  assign n1323 = ~n1289 & ~n1291 ;
  assign n1118 = \key3[25]_pad  & n329 ;
  assign n1116 = \key2[25]_pad  & n319 ;
  assign n1117 = \key1[25]_pad  & n327 ;
  assign n1119 = ~n1116 & ~n1117 ;
  assign n1120 = ~n1118 & n1119 ;
  assign n1152 = n322 & ~n1120 ;
  assign n1292 = ~n1152 & ~n1160 ;
  assign n1293 = n361 & ~n1292 ;
  assign n1299 = n322 & ~n1298 ;
  assign n1300 = ~n1192 & ~n1299 ;
  assign n1301 = n392 & ~n1300 ;
  assign n1324 = ~n1293 & ~n1301 ;
  assign n1334 = n1323 & n1324 ;
  assign n1335 = n1333 & n1334 ;
  assign n1316 = n453 & ~n1073 ;
  assign n1099 = \key3[54]_pad  & n329 ;
  assign n1097 = \key2[54]_pad  & n319 ;
  assign n1098 = \key1[54]_pad  & n327 ;
  assign n1100 = ~n1097 & ~n1098 ;
  assign n1101 = ~n1099 & n1100 ;
  assign n1102 = ~n322 & ~n1101 ;
  assign n1317 = ~n1102 & ~n1203 ;
  assign n1318 = n408 & ~n1317 ;
  assign n1329 = ~n1316 & ~n1318 ;
  assign n1174 = n322 & ~n1173 ;
  assign n1319 = ~n1135 & ~n1174 ;
  assign n1320 = n458 & ~n1319 ;
  assign n1113 = n322 & ~n1109 ;
  assign n1321 = ~n1113 & ~n1198 ;
  assign n1322 = n448 & ~n1321 ;
  assign n1330 = ~n1320 & ~n1322 ;
  assign n1331 = n1329 & n1330 ;
  assign n1149 = ~n322 & ~n1145 ;
  assign n1309 = ~n1149 & ~n1188 ;
  assign n1310 = n463 & ~n1309 ;
  assign n1138 = n322 & ~n1101 ;
  assign n1311 = ~n1138 & ~n1182 ;
  assign n1312 = n443 & ~n1311 ;
  assign n1327 = ~n1310 & ~n1312 ;
  assign n1313 = n306 & ~n947 ;
  assign n1121 = ~n322 & ~n1120 ;
  assign n1314 = ~n1121 & ~n1191 ;
  assign n1315 = n438 & ~n1314 ;
  assign n1328 = ~n1313 & ~n1315 ;
  assign n1332 = n1327 & n1328 ;
  assign n1336 = n1331 & n1332 ;
  assign n1337 = n1335 & n1336 ;
  assign n1338 = \desIn[45]_pad  & n308 ;
  assign n1340 = ~\FP_R_reg[14]/P0001  & n313 ;
  assign n1339 = ~\FP_R_reg[46]/NET0131  & ~n313 ;
  assign n1341 = ~n308 & ~n1339 ;
  assign n1342 = ~n1340 & n1341 ;
  assign n1343 = ~n1338 & ~n1342 ;
  assign n1344 = ~n1337 & ~n1343 ;
  assign n1345 = n1337 & n1343 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = n1287 & n1346 ;
  assign n1136 = ~n1129 & ~n1135 ;
  assign n1137 = n438 & ~n1136 ;
  assign n1139 = ~n1005 & ~n1138 ;
  assign n1140 = n483 & ~n1139 ;
  assign n1208 = ~n1137 & ~n1140 ;
  assign n1147 = ~n1063 & ~n1146 ;
  assign n1148 = n443 & ~n1147 ;
  assign n1150 = ~n940 & ~n1149 ;
  assign n1151 = n408 & ~n1150 ;
  assign n1209 = ~n1148 & ~n1151 ;
  assign n1216 = n1208 & n1209 ;
  assign n1103 = ~n996 & ~n1102 ;
  assign n1104 = n306 & ~n1103 ;
  assign n1111 = ~n1067 & ~n1110 ;
  assign n1112 = n377 & ~n1111 ;
  assign n1206 = ~n1104 & ~n1112 ;
  assign n1114 = ~n1046 & ~n1113 ;
  assign n1115 = n453 & ~n1114 ;
  assign n1122 = ~n1018 & ~n1121 ;
  assign n1123 = n344 & ~n1122 ;
  assign n1207 = ~n1115 & ~n1123 ;
  assign n1217 = n1206 & n1207 ;
  assign n1218 = n1216 & n1217 ;
  assign n1193 = ~n1191 & ~n1192 ;
  assign n1194 = n458 & ~n1193 ;
  assign n1196 = ~n1075 & ~n1195 ;
  assign n1197 = n478 & ~n1196 ;
  assign n1212 = ~n1194 & ~n1197 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = n361 & ~n1200 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1205 = n463 & ~n1204 ;
  assign n1213 = ~n1201 & ~n1205 ;
  assign n1214 = n1212 & n1213 ;
  assign n1153 = ~n1071 & ~n1152 ;
  assign n1154 = n448 & ~n1153 ;
  assign n1167 = ~n1160 & ~n1166 ;
  assign n1168 = n423 & ~n1167 ;
  assign n1210 = ~n1154 & ~n1168 ;
  assign n1175 = ~n968 & ~n1174 ;
  assign n1176 = n392 & ~n1175 ;
  assign n1189 = ~n1182 & ~n1188 ;
  assign n1190 = n488 & ~n1189 ;
  assign n1211 = ~n1176 & ~n1190 ;
  assign n1215 = n1210 & n1211 ;
  assign n1219 = n1214 & n1215 ;
  assign n1220 = n1218 & n1219 ;
  assign n1224 = ~\FP_R_reg[44]/NET0131  & n311 ;
  assign n1223 = ~\FP_R_reg[12]/P0001  & ~n311 ;
  assign n1225 = ~n307 & ~n1223 ;
  assign n1226 = ~n1224 & n1225 ;
  assign n1221 = \FP_R_reg[44]/NET0131  & n312 ;
  assign n1222 = \desIn[29]_pad  & n308 ;
  assign n1227 = ~n1221 & ~n1222 ;
  assign n1228 = ~n1226 & n1227 ;
  assign n1229 = ~n1220 & n1228 ;
  assign n1230 = n1220 & ~n1228 ;
  assign n1231 = ~n1229 & ~n1230 ;
  assign n1354 = ~n1052 & ~n1056 ;
  assign n1355 = n463 & ~n1354 ;
  assign n1356 = n453 & ~n1103 ;
  assign n1378 = ~n1355 & ~n1356 ;
  assign n1357 = ~n974 & ~n982 ;
  assign n1358 = n423 & ~n1357 ;
  assign n1359 = ~n1002 & ~n1010 ;
  assign n1360 = n361 & ~n1359 ;
  assign n1379 = ~n1358 & ~n1360 ;
  assign n1386 = n1378 & n1379 ;
  assign n1348 = ~n1032 & ~n1072 ;
  assign n1349 = n408 & ~n1348 ;
  assign n1350 = n377 & ~n1139 ;
  assign n1376 = ~n1349 & ~n1350 ;
  assign n1351 = n306 & ~n1114 ;
  assign n1352 = ~n1024 & ~n1055 ;
  assign n1353 = n443 & ~n1352 ;
  assign n1377 = ~n1351 & ~n1353 ;
  assign n1387 = n1376 & n1377 ;
  assign n1388 = n1386 & n1387 ;
  assign n1369 = ~n1009 & ~n1299 ;
  assign n1370 = n478 & ~n1369 ;
  assign n1371 = n483 & ~n1111 ;
  assign n1382 = ~n1370 & ~n1371 ;
  assign n1372 = ~n946 & ~n988 ;
  assign n1373 = n448 & ~n1372 ;
  assign n1374 = ~n954 & ~n1306 ;
  assign n1375 = n392 & ~n1374 ;
  assign n1383 = ~n1373 & ~n1375 ;
  assign n1384 = n1382 & n1383 ;
  assign n1361 = ~n1038 & ~n1068 ;
  assign n1362 = n488 & ~n1361 ;
  assign n1363 = ~n960 & ~n1006 ;
  assign n1364 = n438 & ~n1363 ;
  assign n1380 = ~n1362 & ~n1364 ;
  assign n1365 = ~n1060 & ~n1064 ;
  assign n1366 = n344 & ~n1365 ;
  assign n1367 = ~n1059 & ~n1076 ;
  assign n1368 = n458 & ~n1367 ;
  assign n1381 = ~n1366 & ~n1368 ;
  assign n1385 = n1380 & n1381 ;
  assign n1389 = n1384 & n1385 ;
  assign n1390 = n1388 & n1389 ;
  assign n1391 = ~n626 & n1390 ;
  assign n1392 = n626 & ~n1390 ;
  assign n1393 = ~n1391 & ~n1392 ;
  assign n1485 = n1231 & ~n1393 ;
  assign n1493 = ~n1347 & ~n1485 ;
  assign n1402 = ~n954 & ~n1135 ;
  assign n1403 = n408 & ~n1402 ;
  assign n1404 = ~n1060 & ~n1191 ;
  assign n1405 = n453 & ~n1404 ;
  assign n1428 = ~n1403 & ~n1405 ;
  assign n1406 = ~n1059 & ~n1121 ;
  assign n1407 = n306 & ~n1406 ;
  assign n1408 = ~n1018 & ~n1063 ;
  assign n1409 = n361 & ~n1408 ;
  assign n1429 = ~n1407 & ~n1409 ;
  assign n1436 = n1428 & n1429 ;
  assign n1394 = ~n968 & ~n1166 ;
  assign n1395 = n488 & ~n1394 ;
  assign n1396 = ~n1055 & ~n1202 ;
  assign n1397 = n478 & ~n1396 ;
  assign n1426 = ~n1395 & ~n1397 ;
  assign n1398 = ~n1075 & ~n1192 ;
  assign n1399 = n463 & ~n1398 ;
  assign n1400 = ~n996 & ~n1198 ;
  assign n1401 = n344 & ~n1400 ;
  assign n1427 = ~n1399 & ~n1401 ;
  assign n1437 = n1426 & n1427 ;
  assign n1438 = n1436 & n1437 ;
  assign n1418 = ~n988 & ~n1160 ;
  assign n1419 = n377 & ~n1418 ;
  assign n1420 = ~n1067 & ~n1182 ;
  assign n1421 = n423 & ~n1420 ;
  assign n1432 = ~n1419 & ~n1421 ;
  assign n1422 = ~n1032 & ~n1188 ;
  assign n1423 = n392 & ~n1422 ;
  assign n1424 = ~n1046 & ~n1203 ;
  assign n1425 = n458 & ~n1424 ;
  assign n1433 = ~n1423 & ~n1425 ;
  assign n1434 = n1432 & n1433 ;
  assign n1410 = ~n940 & ~n1071 ;
  assign n1411 = n438 & ~n1410 ;
  assign n1412 = ~n1005 & ~n1129 ;
  assign n1413 = n448 & ~n1412 ;
  assign n1430 = ~n1411 & ~n1413 ;
  assign n1414 = ~n982 & ~n1152 ;
  assign n1415 = n483 & ~n1414 ;
  assign n1416 = ~n1009 & ~n1199 ;
  assign n1417 = n443 & ~n1416 ;
  assign n1431 = ~n1415 & ~n1417 ;
  assign n1435 = n1430 & n1431 ;
  assign n1439 = n1434 & n1435 ;
  assign n1440 = n1438 & n1439 ;
  assign n1441 = \desIn[53]_pad  & n308 ;
  assign n1443 = ~\FP_R_reg[15]/P0001  & n313 ;
  assign n1442 = ~\FP_R_reg[47]/NET0131  & ~n313 ;
  assign n1444 = ~n308 & ~n1442 ;
  assign n1445 = ~n1443 & n1444 ;
  assign n1446 = ~n1441 & ~n1445 ;
  assign n1447 = ~n1440 & n1446 ;
  assign n1448 = n1440 & ~n1446 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1459 = ~n1231 & n1393 ;
  assign n1492 = n1347 & ~n1459 ;
  assign n1494 = ~n1449 & ~n1492 ;
  assign n1495 = ~n1493 & n1494 ;
  assign n1476 = n1231 & n1393 ;
  assign n1477 = ~n1346 & n1476 ;
  assign n1478 = n1287 & n1477 ;
  assign n1455 = ~n1287 & ~n1346 ;
  assign n1479 = n1455 & n1459 ;
  assign n1480 = ~n1478 & ~n1479 ;
  assign n1462 = ~n1231 & ~n1393 ;
  assign n1484 = n1287 & n1449 ;
  assign n1488 = n1462 & n1484 ;
  assign n1489 = ~n1287 & n1346 ;
  assign n1454 = n1231 & n1449 ;
  assign n1490 = n1393 & n1454 ;
  assign n1491 = n1489 & n1490 ;
  assign n1496 = ~n1488 & ~n1491 ;
  assign n1497 = n1480 & n1496 ;
  assign n1498 = ~n1495 & n1497 ;
  assign n1499 = n1096 & ~n1498 ;
  assign n1460 = n1449 & n1459 ;
  assign n1461 = n1346 & n1460 ;
  assign n1456 = ~n1287 & ~n1393 ;
  assign n1457 = ~n1455 & ~n1456 ;
  assign n1458 = n1454 & ~n1457 ;
  assign n1463 = ~n1287 & ~n1449 ;
  assign n1464 = n1462 & n1463 ;
  assign n1471 = ~n1458 & ~n1464 ;
  assign n1472 = ~n1461 & n1471 ;
  assign n1450 = n1346 & ~n1449 ;
  assign n1451 = n1393 & n1450 ;
  assign n1452 = ~n1347 & ~n1451 ;
  assign n1453 = n1231 & ~n1452 ;
  assign n1465 = ~n1231 & n1287 ;
  assign n1466 = ~n1346 & n1465 ;
  assign n1467 = ~n1393 & n1466 ;
  assign n1468 = n1346 & n1462 ;
  assign n1469 = ~n1287 & n1468 ;
  assign n1470 = ~n1467 & ~n1469 ;
  assign n1473 = ~n1453 & n1470 ;
  assign n1474 = n1472 & n1473 ;
  assign n1475 = ~n1096 & ~n1474 ;
  assign n1481 = ~n1469 & n1480 ;
  assign n1482 = ~n1449 & ~n1481 ;
  assign n1483 = n1449 & n1466 ;
  assign n1486 = n1484 & n1485 ;
  assign n1487 = n1346 & n1486 ;
  assign n1500 = ~n1483 & ~n1487 ;
  assign n1501 = ~n1482 & n1500 ;
  assign n1502 = ~n1475 & n1501 ;
  assign n1503 = ~n1499 & n1502 ;
  assign n1504 = ~\desIn[12]_pad  & n308 ;
  assign n1506 = \FP_R_reg[10]/P0001  & ~n313 ;
  assign n1505 = \FP_R_reg[42]/NET0131  & n313 ;
  assign n1507 = ~n308 & ~n1505 ;
  assign n1508 = ~n1506 & n1507 ;
  assign n1509 = ~n1504 & ~n1508 ;
  assign n1510 = n1503 & ~n1509 ;
  assign n1511 = ~n1503 & n1509 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = \desIn[13]_pad  & n308 ;
  assign n1515 = ~\FP_R_reg[10]/P0001  & n313 ;
  assign n1514 = ~\FP_R_reg[42]/NET0131  & ~n313 ;
  assign n1516 = ~n308 & ~n1514 ;
  assign n1517 = ~n1515 & n1516 ;
  assign n1518 = ~n1513 & ~n1517 ;
  assign n1519 = \desIn[63]_pad  & n308 ;
  assign n1521 = ~\FP_R_reg[8]/P0001  & n313 ;
  assign n1520 = ~\FP_R_reg[40]/NET0131  & ~n313 ;
  assign n1522 = ~n308 & ~n1520 ;
  assign n1523 = ~n1521 & n1522 ;
  assign n1524 = ~n1519 & ~n1523 ;
  assign n1532 = ~n1006 & ~n1149 ;
  assign n1533 = n443 & ~n1532 ;
  assign n1534 = ~n1052 & ~n1195 ;
  assign n1535 = n448 & ~n1534 ;
  assign n1555 = ~n1533 & ~n1535 ;
  assign n1536 = ~n1064 & ~n1102 ;
  assign n1537 = n488 & ~n1536 ;
  assign n1538 = n377 & ~n1236 ;
  assign n1556 = ~n1537 & ~n1538 ;
  assign n1563 = n1555 & n1556 ;
  assign n1525 = n306 & ~n1258 ;
  assign n1526 = ~n946 & ~n1138 ;
  assign n1527 = n463 & ~n1526 ;
  assign n1553 = ~n1525 & ~n1527 ;
  assign n1528 = ~n1072 & ~n1306 ;
  assign n1529 = n361 & ~n1528 ;
  assign n1530 = ~n1024 & ~n1299 ;
  assign n1531 = n438 & ~n1530 ;
  assign n1554 = ~n1529 & ~n1531 ;
  assign n1564 = n1553 & n1554 ;
  assign n1565 = n1563 & n1564 ;
  assign n1547 = n453 & ~n1234 ;
  assign n1548 = ~n1010 & ~n1121 ;
  assign n1549 = n392 & ~n1548 ;
  assign n1559 = ~n1547 & ~n1549 ;
  assign n1550 = n483 & ~n1242 ;
  assign n1551 = ~n974 & ~n1110 ;
  assign n1552 = n458 & ~n1551 ;
  assign n1560 = ~n1550 & ~n1552 ;
  assign n1561 = n1559 & n1560 ;
  assign n1539 = ~n1068 & ~n1174 ;
  assign n1540 = n344 & ~n1539 ;
  assign n1541 = ~n1076 & ~n1113 ;
  assign n1542 = n423 & ~n1541 ;
  assign n1557 = ~n1540 & ~n1542 ;
  assign n1543 = ~n960 & ~n1152 ;
  assign n1544 = n478 & ~n1543 ;
  assign n1545 = ~n1002 & ~n1146 ;
  assign n1546 = n408 & ~n1545 ;
  assign n1558 = ~n1544 & ~n1546 ;
  assign n1562 = n1557 & n1558 ;
  assign n1566 = n1561 & n1562 ;
  assign n1567 = n1565 & n1566 ;
  assign n1568 = n1524 & n1567 ;
  assign n1569 = ~n1524 & ~n1567 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1807 = n453 & ~n1406 ;
  assign n1808 = ~n1002 & ~n1113 ;
  assign n1809 = n344 & ~n1808 ;
  assign n1830 = ~n1807 & ~n1809 ;
  assign n1810 = ~n1056 & ~n1146 ;
  assign n1811 = n478 & ~n1810 ;
  assign n1812 = ~n946 & ~n1072 ;
  assign n1813 = n438 & ~n1812 ;
  assign n1831 = ~n1811 & ~n1813 ;
  assign n1838 = n1830 & n1831 ;
  assign n1800 = n306 & ~n1404 ;
  assign n1801 = ~n1010 & ~n1195 ;
  assign n1802 = n443 & ~n1801 ;
  assign n1828 = ~n1800 & ~n1802 ;
  assign n1803 = ~n1076 & ~n1299 ;
  assign n1804 = n463 & ~n1803 ;
  assign n1805 = ~n1024 & ~n1064 ;
  assign n1806 = n361 & ~n1805 ;
  assign n1829 = ~n1804 & ~n1806 ;
  assign n1839 = n1828 & n1829 ;
  assign n1840 = n1838 & n1839 ;
  assign n1821 = ~n1068 & ~n1138 ;
  assign n1822 = n423 & ~n1821 ;
  assign n1823 = n483 & ~n1418 ;
  assign n1834 = ~n1822 & ~n1823 ;
  assign n1824 = ~n1006 & ~n1110 ;
  assign n1825 = n448 & ~n1824 ;
  assign n1826 = ~n1038 & ~n1149 ;
  assign n1827 = n392 & ~n1826 ;
  assign n1835 = ~n1825 & ~n1827 ;
  assign n1836 = n1834 & n1835 ;
  assign n1814 = ~n974 & ~n1306 ;
  assign n1815 = n488 & ~n1814 ;
  assign n1816 = ~n960 & ~n1174 ;
  assign n1817 = n408 & ~n1816 ;
  assign n1832 = ~n1815 & ~n1817 ;
  assign n1818 = n377 & ~n1414 ;
  assign n1819 = ~n1052 & ~n1102 ;
  assign n1820 = n458 & ~n1819 ;
  assign n1833 = ~n1818 & ~n1820 ;
  assign n1837 = n1832 & n1833 ;
  assign n1841 = n1836 & n1837 ;
  assign n1842 = n1840 & n1841 ;
  assign n1846 = ~\FP_R_reg[39]/NET0131  & n311 ;
  assign n1845 = ~\FP_R_reg[7]/P0001  & ~n311 ;
  assign n1847 = ~n307 & ~n1845 ;
  assign n1848 = ~n1846 & n1847 ;
  assign n1843 = \FP_R_reg[39]/NET0131  & n312 ;
  assign n1844 = \desIn[55]_pad  & n308 ;
  assign n1849 = ~n1843 & ~n1844 ;
  assign n1850 = ~n1848 & n1849 ;
  assign n1851 = ~n1842 & n1850 ;
  assign n1852 = n1842 & ~n1850 ;
  assign n1853 = ~n1851 & ~n1852 ;
  assign n1627 = \desIn[39]_pad  & n308 ;
  assign n1629 = ~\FP_R_reg[5]/P0001  & n313 ;
  assign n1628 = ~\FP_R_reg[37]/NET0131  & ~n313 ;
  assign n1630 = ~n308 & ~n1628 ;
  assign n1631 = ~n1629 & n1630 ;
  assign n1632 = ~n1627 & ~n1631 ;
  assign n1641 = ~n1024 & ~n1075 ;
  assign n1642 = n453 & ~n1641 ;
  assign n1643 = ~n960 & ~n988 ;
  assign n1644 = n488 & ~n1643 ;
  assign n1667 = ~n1642 & ~n1644 ;
  assign n1645 = ~n954 & ~n1068 ;
  assign n1646 = n448 & ~n1645 ;
  assign n1647 = ~n946 & ~n1067 ;
  assign n1648 = n392 & ~n1647 ;
  assign n1668 = ~n1646 & ~n1648 ;
  assign n1675 = n1667 & n1668 ;
  assign n1633 = ~n968 & ~n1072 ;
  assign n1634 = n377 & ~n1633 ;
  assign n1635 = ~n974 & ~n1005 ;
  assign n1636 = n408 & ~n1635 ;
  assign n1665 = ~n1634 & ~n1636 ;
  assign n1637 = ~n1046 & ~n1064 ;
  assign n1638 = n478 & ~n1637 ;
  assign n1639 = ~n1056 & ~n1059 ;
  assign n1640 = n361 & ~n1639 ;
  assign n1666 = ~n1638 & ~n1640 ;
  assign n1676 = n1665 & n1666 ;
  assign n1677 = n1675 & n1676 ;
  assign n1657 = ~n982 & ~n1038 ;
  assign n1658 = n438 & ~n1657 ;
  assign n1659 = ~n940 & ~n1306 ;
  assign n1660 = n483 & ~n1659 ;
  assign n1671 = ~n1658 & ~n1660 ;
  assign n1661 = ~n1010 & ~n1060 ;
  assign n1662 = n463 & ~n1661 ;
  assign n1663 = ~n1002 & ~n1055 ;
  assign n1664 = n458 & ~n1663 ;
  assign n1672 = ~n1662 & ~n1664 ;
  assign n1673 = n1671 & n1672 ;
  assign n1649 = ~n1006 & ~n1032 ;
  assign n1650 = n423 & ~n1649 ;
  assign n1651 = ~n996 & ~n1076 ;
  assign n1652 = n443 & ~n1651 ;
  assign n1669 = ~n1650 & ~n1652 ;
  assign n1653 = ~n1063 & ~n1299 ;
  assign n1654 = n306 & ~n1653 ;
  assign n1655 = ~n1009 & ~n1052 ;
  assign n1656 = n344 & ~n1655 ;
  assign n1670 = ~n1654 & ~n1656 ;
  assign n1674 = n1669 & n1670 ;
  assign n1678 = n1673 & n1674 ;
  assign n1679 = n1677 & n1678 ;
  assign n1680 = n1632 & n1679 ;
  assign n1681 = ~n1632 & ~n1679 ;
  assign n1682 = ~n1680 & ~n1681 ;
  assign n1683 = \desIn[5]_pad  & n308 ;
  assign n1685 = ~\FP_R_reg[9]/P0001  & n313 ;
  assign n1684 = ~\FP_R_reg[41]/NET0131  & ~n313 ;
  assign n1686 = ~n308 & ~n1684 ;
  assign n1687 = ~n1685 & n1686 ;
  assign n1688 = ~n1683 & ~n1687 ;
  assign n1697 = ~n1068 & ~n1129 ;
  assign n1698 = n377 & ~n1697 ;
  assign n1699 = ~n974 & ~n1135 ;
  assign n1700 = n392 & ~n1699 ;
  assign n1723 = ~n1698 & ~n1700 ;
  assign n1701 = ~n946 & ~n1188 ;
  assign n1702 = n408 & ~n1701 ;
  assign n1703 = ~n1152 & ~n1306 ;
  assign n1704 = n423 & ~n1703 ;
  assign n1724 = ~n1702 & ~n1704 ;
  assign n1731 = n1723 & n1724 ;
  assign n1689 = ~n1002 & ~n1203 ;
  assign n1690 = n306 & ~n1689 ;
  assign n1691 = ~n1110 & ~n1174 ;
  assign n1692 = n438 & ~n1691 ;
  assign n1721 = ~n1690 & ~n1692 ;
  assign n1693 = ~n1102 & ~n1146 ;
  assign n1694 = n463 & ~n1693 ;
  assign n1695 = ~n1072 & ~n1160 ;
  assign n1696 = n448 & ~n1695 ;
  assign n1722 = ~n1694 & ~n1696 ;
  assign n1732 = n1721 & n1722 ;
  assign n1733 = n1731 & n1732 ;
  assign n1713 = ~n1121 & ~n1299 ;
  assign n1714 = n458 & ~n1713 ;
  assign n1715 = ~n1052 & ~n1198 ;
  assign n1716 = n453 & ~n1715 ;
  assign n1727 = ~n1714 & ~n1716 ;
  assign n1717 = ~n1113 & ~n1195 ;
  assign n1718 = n361 & ~n1717 ;
  assign n1719 = ~n1076 & ~n1199 ;
  assign n1720 = n478 & ~n1719 ;
  assign n1728 = ~n1718 & ~n1720 ;
  assign n1729 = n1727 & n1728 ;
  assign n1705 = ~n1064 & ~n1202 ;
  assign n1706 = n443 & ~n1705 ;
  assign n1707 = ~n1138 & ~n1149 ;
  assign n1708 = n488 & ~n1707 ;
  assign n1725 = ~n1706 & ~n1708 ;
  assign n1709 = ~n1006 & ~n1182 ;
  assign n1710 = n483 & ~n1709 ;
  assign n1711 = ~n1024 & ~n1191 ;
  assign n1712 = n344 & ~n1711 ;
  assign n1726 = ~n1710 & ~n1712 ;
  assign n1730 = n1725 & n1726 ;
  assign n1734 = n1729 & n1730 ;
  assign n1735 = n1733 & n1734 ;
  assign n1736 = n1688 & n1735 ;
  assign n1737 = ~n1688 & ~n1735 ;
  assign n1738 = ~n1736 & ~n1737 ;
  assign n1740 = \desIn[31]_pad  & n308 ;
  assign n1742 = ~\FP_R_reg[4]/P0001  & n313 ;
  assign n1741 = ~\FP_R_reg[36]/NET0131  & ~n313 ;
  assign n1743 = ~n308 & ~n1741 ;
  assign n1744 = ~n1742 & n1743 ;
  assign n1745 = ~n1740 & ~n1744 ;
  assign n1754 = ~n996 & ~n1195 ;
  assign n1755 = n377 & ~n1754 ;
  assign n1756 = ~n1198 & ~n1203 ;
  assign n1757 = n438 & ~n1756 ;
  assign n1780 = ~n1755 & ~n1757 ;
  assign n1758 = ~n1063 & ~n1191 ;
  assign n1759 = n448 & ~n1758 ;
  assign n1760 = ~n1067 & ~n1149 ;
  assign n1761 = n478 & ~n1760 ;
  assign n1781 = ~n1759 & ~n1761 ;
  assign n1788 = n1780 & n1781 ;
  assign n1746 = ~n954 & ~n1110 ;
  assign n1747 = n306 & ~n1746 ;
  assign n1748 = ~n1018 & ~n1202 ;
  assign n1749 = n423 & ~n1748 ;
  assign n1778 = ~n1747 & ~n1749 ;
  assign n1750 = ~n1129 & ~n1182 ;
  assign n1751 = n361 & ~n1750 ;
  assign n1752 = ~n1135 & ~n1166 ;
  assign n1753 = n463 & ~n1752 ;
  assign n1779 = ~n1751 & ~n1753 ;
  assign n1789 = n1778 & n1779 ;
  assign n1790 = n1788 & n1789 ;
  assign n1770 = ~n1071 & ~n1188 ;
  assign n1771 = n458 & ~n1770 ;
  assign n1772 = ~n1009 & ~n1113 ;
  assign n1773 = n483 & ~n1772 ;
  assign n1784 = ~n1771 & ~n1773 ;
  assign n1774 = ~n968 & ~n1152 ;
  assign n1775 = n443 & ~n1774 ;
  assign n1776 = ~n1075 & ~n1121 ;
  assign n1777 = n408 & ~n1776 ;
  assign n1785 = ~n1775 & ~n1777 ;
  assign n1786 = n1784 & n1785 ;
  assign n1762 = ~n1192 & ~n1199 ;
  assign n1763 = n488 & ~n1762 ;
  assign n1764 = ~n940 & ~n1160 ;
  assign n1765 = n344 & ~n1764 ;
  assign n1782 = ~n1763 & ~n1765 ;
  assign n1766 = ~n1005 & ~n1174 ;
  assign n1767 = n453 & ~n1766 ;
  assign n1768 = ~n1046 & ~n1146 ;
  assign n1769 = n392 & ~n1768 ;
  assign n1783 = ~n1767 & ~n1769 ;
  assign n1787 = n1782 & n1783 ;
  assign n1791 = n1786 & n1787 ;
  assign n1792 = n1790 & n1791 ;
  assign n1793 = n1745 & ~n1792 ;
  assign n1794 = ~n1745 & n1792 ;
  assign n1795 = ~n1793 & ~n1794 ;
  assign n1796 = ~n1738 & ~n1795 ;
  assign n1797 = n1682 & n1796 ;
  assign n1854 = n1682 & ~n1738 ;
  assign n1571 = \desIn[47]_pad  & n308 ;
  assign n1573 = ~\FP_R_reg[6]/P0001  & n313 ;
  assign n1572 = ~\FP_R_reg[38]/NET0131  & ~n313 ;
  assign n1574 = ~n308 & ~n1572 ;
  assign n1575 = ~n1573 & n1574 ;
  assign n1576 = ~n1571 & ~n1575 ;
  assign n1585 = ~n1067 & ~n1306 ;
  assign n1586 = n453 & ~n1585 ;
  assign n1587 = ~n988 & ~n1068 ;
  assign n1588 = n458 & ~n1587 ;
  assign n1611 = ~n1586 & ~n1588 ;
  assign n1589 = ~n1005 & ~n1072 ;
  assign n1590 = n478 & ~n1589 ;
  assign n1591 = ~n974 & ~n1032 ;
  assign n1592 = n344 & ~n1591 ;
  assign n1612 = ~n1590 & ~n1592 ;
  assign n1619 = n1611 & n1612 ;
  assign n1577 = ~n968 & ~n1138 ;
  assign n1578 = n306 & ~n1577 ;
  assign n1579 = ~n1009 & ~n1064 ;
  assign n1580 = n408 & ~n1579 ;
  assign n1609 = ~n1578 & ~n1580 ;
  assign n1581 = ~n1052 & ~n1060 ;
  assign n1582 = n423 & ~n1581 ;
  assign n1583 = ~n996 & ~n1024 ;
  assign n1584 = n392 & ~n1583 ;
  assign n1610 = ~n1582 & ~n1584 ;
  assign n1620 = n1609 & n1610 ;
  assign n1621 = n1619 & n1620 ;
  assign n1601 = ~n982 & ~n1006 ;
  assign n1602 = n463 & ~n1601 ;
  assign n1603 = ~n1046 & ~n1299 ;
  assign n1604 = n377 & ~n1603 ;
  assign n1615 = ~n1602 & ~n1604 ;
  assign n1605 = ~n1055 & ~n1076 ;
  assign n1606 = n448 & ~n1605 ;
  assign n1607 = ~n960 & ~n1038 ;
  assign n1608 = n361 & ~n1607 ;
  assign n1616 = ~n1606 & ~n1608 ;
  assign n1617 = n1615 & n1616 ;
  assign n1593 = ~n1002 & ~n1059 ;
  assign n1594 = n488 & ~n1593 ;
  assign n1595 = ~n946 & ~n954 ;
  assign n1596 = n443 & ~n1595 ;
  assign n1613 = ~n1594 & ~n1596 ;
  assign n1597 = ~n1075 & ~n1102 ;
  assign n1598 = n483 & ~n1597 ;
  assign n1599 = ~n1010 & ~n1056 ;
  assign n1600 = n438 & ~n1599 ;
  assign n1614 = ~n1598 & ~n1600 ;
  assign n1618 = n1613 & n1614 ;
  assign n1622 = n1617 & n1618 ;
  assign n1623 = n1621 & n1622 ;
  assign n1624 = ~n1576 & n1623 ;
  assign n1625 = n1576 & ~n1623 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1855 = n1626 & n1795 ;
  assign n1856 = ~n1854 & n1855 ;
  assign n1857 = ~n1797 & ~n1856 ;
  assign n1858 = ~n1853 & ~n1857 ;
  assign n1739 = ~n1682 & n1738 ;
  assign n1798 = ~n1739 & ~n1797 ;
  assign n1799 = ~n1626 & ~n1798 ;
  assign n1859 = n1626 & n1682 ;
  assign n1860 = ~n1738 & n1795 ;
  assign n1861 = n1859 & n1860 ;
  assign n1862 = n1853 & n1861 ;
  assign n1863 = n1626 & ~n1682 ;
  assign n1864 = n1796 & n1863 ;
  assign n1865 = ~n1626 & n1682 ;
  assign n1866 = ~n1738 & ~n1853 ;
  assign n1867 = n1865 & n1866 ;
  assign n1868 = ~n1864 & ~n1867 ;
  assign n1869 = ~n1862 & n1868 ;
  assign n1870 = ~n1799 & n1869 ;
  assign n1871 = ~n1858 & n1870 ;
  assign n1872 = n1570 & ~n1871 ;
  assign n1873 = ~n1682 & n1795 ;
  assign n1874 = ~n1626 & ~n1682 ;
  assign n1875 = ~n1873 & ~n1874 ;
  assign n1876 = n1853 & ~n1875 ;
  assign n1877 = n1738 & n1795 ;
  assign n1878 = n1682 & n1877 ;
  assign n1879 = ~n1682 & ~n1738 ;
  assign n1880 = n1795 & n1879 ;
  assign n1881 = ~n1878 & ~n1880 ;
  assign n1882 = ~n1626 & ~n1881 ;
  assign n1883 = ~n1876 & ~n1882 ;
  assign n1884 = ~n1570 & ~n1883 ;
  assign n1885 = ~n1795 & n1859 ;
  assign n1886 = n1738 & n1885 ;
  assign n1887 = ~n1626 & n1873 ;
  assign n1888 = n1853 & ~n1887 ;
  assign n1889 = ~n1886 & n1888 ;
  assign n1890 = ~n1626 & n1797 ;
  assign n1891 = ~n1853 & ~n1864 ;
  assign n1892 = ~n1890 & n1891 ;
  assign n1893 = ~n1889 & ~n1892 ;
  assign n1894 = n1738 & ~n1795 ;
  assign n1895 = ~n1861 & ~n1894 ;
  assign n1896 = ~n1570 & ~n1853 ;
  assign n1897 = ~n1874 & n1896 ;
  assign n1898 = ~n1895 & n1897 ;
  assign n1899 = ~n1893 & ~n1898 ;
  assign n1900 = ~n1884 & n1899 ;
  assign n1901 = ~n1872 & n1900 ;
  assign n1902 = ~\desIn[14]_pad  & n308 ;
  assign n1904 = \FP_R_reg[2]/P0001  & ~n313 ;
  assign n1903 = \FP_R_reg[34]/NET0131  & n313 ;
  assign n1905 = ~n308 & ~n1903 ;
  assign n1906 = ~n1904 & n1905 ;
  assign n1907 = ~n1902 & ~n1906 ;
  assign n1908 = n1901 & ~n1907 ;
  assign n1909 = ~n1901 & n1907 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1914 = ~\FP_R_reg[34]/NET0131  & n311 ;
  assign n1913 = ~\FP_R_reg[2]/P0001  & ~n311 ;
  assign n1915 = ~n307 & ~n1913 ;
  assign n1916 = ~n1914 & n1915 ;
  assign n1911 = \FP_R_reg[34]/NET0131  & n312 ;
  assign n1912 = \desIn[15]_pad  & n308 ;
  assign n1917 = ~n1911 & ~n1912 ;
  assign n1918 = ~n1916 & n1917 ;
  assign n2130 = \desIn[51]_pad  & n308 ;
  assign n2132 = ~\FP_R_reg[23]/P0001  & n313 ;
  assign n2131 = ~\FP_R_reg[55]/NET0131  & ~n313 ;
  assign n2133 = ~n308 & ~n2131 ;
  assign n2134 = ~n2132 & n2133 ;
  assign n2135 = ~n2130 & ~n2134 ;
  assign n2142 = ~n414 & ~n439 ;
  assign n2143 = n423 & ~n2142 ;
  assign n2144 = ~n469 & ~n479 ;
  assign n2145 = n344 & ~n2144 ;
  assign n2166 = ~n2143 & ~n2145 ;
  assign n2146 = ~n454 & ~n460 ;
  assign n2147 = n443 & ~n2146 ;
  assign n2148 = ~n333 & ~n356 ;
  assign n2149 = n478 & ~n2148 ;
  assign n2167 = ~n2147 & ~n2149 ;
  assign n2174 = n2166 & n2167 ;
  assign n2136 = n453 & ~n830 ;
  assign n2137 = ~n440 & ~n449 ;
  assign n2138 = n488 & ~n2137 ;
  assign n2164 = ~n2136 & ~n2138 ;
  assign n2139 = ~n398 & ~n490 ;
  assign n2140 = n448 & ~n2139 ;
  assign n2141 = n483 & ~n844 ;
  assign n2165 = ~n2140 & ~n2141 ;
  assign n2175 = n2164 & n2165 ;
  assign n2176 = n2174 & n2175 ;
  assign n2157 = ~n373 & ~n444 ;
  assign n2158 = n458 & ~n2157 ;
  assign n2159 = ~n383 & ~n435 ;
  assign n2160 = n408 & ~n2159 ;
  assign n2170 = ~n2158 & ~n2160 ;
  assign n2161 = n377 & ~n828 ;
  assign n2162 = ~n350 & ~n367 ;
  assign n2163 = n463 & ~n2162 ;
  assign n2171 = ~n2161 & ~n2163 ;
  assign n2172 = n2170 & n2171 ;
  assign n2150 = ~n450 & ~n484 ;
  assign n2151 = n392 & ~n2150 ;
  assign n2152 = n306 & ~n820 ;
  assign n2168 = ~n2151 & ~n2152 ;
  assign n2153 = ~n429 & ~n489 ;
  assign n2154 = n438 & ~n2153 ;
  assign n2155 = ~n459 & ~n475 ;
  assign n2156 = n361 & ~n2155 ;
  assign n2169 = ~n2154 & ~n2156 ;
  assign n2173 = n2168 & n2169 ;
  assign n2177 = n2172 & n2173 ;
  assign n2178 = n2176 & n2177 ;
  assign n2179 = ~n2135 & n2178 ;
  assign n2180 = n2135 & ~n2178 ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2079 = ~n454 & ~n694 ;
  assign n2080 = n377 & ~n2079 ;
  assign n2081 = ~n564 & ~n567 ;
  assign n2082 = n423 & ~n2081 ;
  assign n2105 = ~n2080 & ~n2082 ;
  assign n2083 = ~n555 & ~n723 ;
  assign n2084 = n408 & ~n2083 ;
  assign n2085 = ~n527 & ~n552 ;
  assign n2086 = n344 & ~n2085 ;
  assign n2106 = ~n2084 & ~n2086 ;
  assign n2113 = n2105 & n2106 ;
  assign n2071 = ~n398 & ~n485 ;
  assign n2072 = n306 & ~n2071 ;
  assign n2073 = ~n586 & ~n594 ;
  assign n2074 = n463 & ~n2073 ;
  assign n2103 = ~n2072 & ~n2074 ;
  assign n2075 = ~n533 & ~n732 ;
  assign n2076 = n443 & ~n2075 ;
  assign n2077 = ~n339 & ~n479 ;
  assign n2078 = n483 & ~n2077 ;
  assign n2104 = ~n2076 & ~n2078 ;
  assign n2114 = n2103 & n2104 ;
  assign n2115 = n2113 & n2114 ;
  assign n2095 = ~n383 & ~n715 ;
  assign n2096 = n453 & ~n2095 ;
  assign n2097 = ~n519 & ~n578 ;
  assign n2098 = n361 & ~n2097 ;
  assign n2109 = ~n2096 & ~n2098 ;
  assign n2099 = ~n516 & ~n575 ;
  assign n2100 = n438 & ~n2099 ;
  assign n2101 = ~n541 & ~n603 ;
  assign n2102 = n458 & ~n2101 ;
  assign n2110 = ~n2100 & ~n2102 ;
  assign n2111 = n2109 & n2110 ;
  assign n2087 = ~n597 & ~n600 ;
  assign n2088 = n488 & ~n2087 ;
  assign n2089 = ~n333 & ~n711 ;
  assign n2090 = n392 & ~n2089 ;
  assign n2107 = ~n2088 & ~n2090 ;
  assign n2091 = ~n549 & ~n556 ;
  assign n2092 = n448 & ~n2091 ;
  assign n2093 = ~n484 & ~n729 ;
  assign n2094 = n478 & ~n2093 ;
  assign n2108 = ~n2092 & ~n2094 ;
  assign n2112 = n2107 & n2108 ;
  assign n2116 = n2111 & n2112 ;
  assign n2117 = n2115 & n2116 ;
  assign n2118 = \desIn[1]_pad  & n308 ;
  assign n2120 = ~\FP_R_reg[25]/P0001  & n313 ;
  assign n2119 = ~\FP_R_reg[57]/NET0131  & ~n313 ;
  assign n2121 = ~n308 & ~n2119 ;
  assign n2122 = ~n2120 & n2121 ;
  assign n2123 = ~n2118 & ~n2122 ;
  assign n2124 = ~n2117 & n2123 ;
  assign n2125 = n2117 & ~n2123 ;
  assign n2126 = ~n2124 & ~n2125 ;
  assign n1927 = ~n356 & ~n556 ;
  assign n1928 = n377 & ~n1927 ;
  assign n1929 = ~n350 & ~n459 ;
  assign n1930 = n438 & ~n1929 ;
  assign n1953 = ~n1928 & ~n1930 ;
  assign n1931 = ~n445 & ~n567 ;
  assign n1932 = n483 & ~n1931 ;
  assign n1933 = ~n420 & ~n541 ;
  assign n1934 = n306 & ~n1933 ;
  assign n1954 = ~n1932 & ~n1934 ;
  assign n1961 = n1953 & n1954 ;
  assign n1919 = ~n333 & ~n469 ;
  assign n1920 = n408 & ~n1919 ;
  assign n1921 = ~n383 & ~n439 ;
  assign n1922 = n344 & ~n1921 ;
  assign n1951 = ~n1920 & ~n1922 ;
  assign n1923 = ~n484 & ~n490 ;
  assign n1924 = n443 & ~n1923 ;
  assign n1925 = ~n398 & ~n440 ;
  assign n1926 = n458 & ~n1925 ;
  assign n1952 = ~n1924 & ~n1926 ;
  assign n1962 = n1951 & n1952 ;
  assign n1963 = n1961 & n1962 ;
  assign n1943 = ~n414 & ~n489 ;
  assign n1944 = n463 & ~n1943 ;
  assign n1945 = ~n367 & ~n479 ;
  assign n1946 = n423 & ~n1945 ;
  assign n1957 = ~n1944 & ~n1946 ;
  assign n1947 = ~n450 & ~n527 ;
  assign n1948 = n453 & ~n1947 ;
  assign n1949 = ~n435 & ~n533 ;
  assign n1950 = n478 & ~n1949 ;
  assign n1958 = ~n1948 & ~n1950 ;
  assign n1959 = n1957 & n1958 ;
  assign n1935 = ~n460 & ~n555 ;
  assign n1936 = n392 & ~n1935 ;
  assign n1937 = ~n429 & ~n449 ;
  assign n1938 = n361 & ~n1937 ;
  assign n1955 = ~n1936 & ~n1938 ;
  assign n1939 = ~n444 & ~n475 ;
  assign n1940 = n488 & ~n1939 ;
  assign n1941 = ~n373 & ~n454 ;
  assign n1942 = n448 & ~n1941 ;
  assign n1956 = ~n1940 & ~n1942 ;
  assign n1960 = n1955 & n1956 ;
  assign n1964 = n1959 & n1960 ;
  assign n1965 = n1963 & n1964 ;
  assign n1966 = ~n318 & n1965 ;
  assign n1967 = n318 & ~n1965 ;
  assign n1968 = ~n1966 & ~n1967 ;
  assign n2029 = ~n339 & ~n455 ;
  assign n2030 = n438 & ~n2029 ;
  assign n2031 = ~n420 & ~n729 ;
  assign n2032 = n458 & ~n2031 ;
  assign n2055 = ~n2030 & ~n2032 ;
  assign n2033 = ~n450 & ~n732 ;
  assign n2034 = n344 & ~n2033 ;
  assign n2035 = ~n440 & ~n519 ;
  assign n2036 = n306 & ~n2035 ;
  assign n2056 = ~n2034 & ~n2036 ;
  assign n2063 = n2055 & n2056 ;
  assign n2021 = ~n373 & ~n597 ;
  assign n2022 = n377 & ~n2021 ;
  assign n2023 = ~n367 & ~n516 ;
  assign n2024 = n483 & ~n2023 ;
  assign n2053 = ~n2022 & ~n2024 ;
  assign n2025 = ~n389 & ~n485 ;
  assign n2026 = n361 & ~n2025 ;
  assign n2027 = ~n445 & ~n711 ;
  assign n2028 = n423 & ~n2027 ;
  assign n2054 = ~n2026 & ~n2028 ;
  assign n2064 = n2053 & n2054 ;
  assign n2065 = n2063 & n2064 ;
  assign n2045 = ~n356 & ~n723 ;
  assign n2046 = n448 & ~n2045 ;
  assign n2047 = ~n480 & ~n694 ;
  assign n2048 = n488 & ~n2047 ;
  assign n2059 = ~n2046 & ~n2048 ;
  assign n2049 = ~n404 & ~n715 ;
  assign n2050 = n463 & ~n2049 ;
  assign n2051 = ~n469 & ~n564 ;
  assign n2052 = n392 & ~n2051 ;
  assign n2060 = ~n2050 & ~n2052 ;
  assign n2061 = n2059 & n2060 ;
  assign n2037 = ~n439 & ~n594 ;
  assign n2038 = n453 & ~n2037 ;
  assign n2039 = ~n490 & ~n603 ;
  assign n2040 = n478 & ~n2039 ;
  assign n2057 = ~n2038 & ~n2040 ;
  assign n2041 = ~n435 & ~n552 ;
  assign n2042 = n443 & ~n2041 ;
  assign n2043 = ~n460 & ~n549 ;
  assign n2044 = n408 & ~n2043 ;
  assign n2058 = ~n2042 & ~n2044 ;
  assign n2062 = n2057 & n2058 ;
  assign n2066 = n2061 & n2062 ;
  assign n2067 = n2065 & n2066 ;
  assign n2068 = n755 & ~n2067 ;
  assign n2069 = ~n755 & n2067 ;
  assign n2070 = ~n2068 & ~n2069 ;
  assign n2188 = ~n1968 & n2070 ;
  assign n2189 = n2126 & n2188 ;
  assign n2184 = ~n1968 & ~n2126 ;
  assign n2190 = ~n2070 & n2184 ;
  assign n2191 = ~n2189 & ~n2190 ;
  assign n2192 = ~n2181 & ~n2191 ;
  assign n1976 = ~n389 & ~n490 ;
  assign n1977 = n423 & ~n1976 ;
  assign n1978 = n453 & ~n763 ;
  assign n1999 = ~n1977 & ~n1978 ;
  assign n1979 = ~n439 & ~n485 ;
  assign n1980 = n448 & ~n1979 ;
  assign n1981 = ~n356 & ~n445 ;
  assign n1982 = n361 & ~n1981 ;
  assign n2000 = ~n1980 & ~n1982 ;
  assign n2007 = n1999 & n2000 ;
  assign n1969 = ~n455 & ~n469 ;
  assign n1970 = n458 & ~n1969 ;
  assign n1971 = n483 & ~n787 ;
  assign n1997 = ~n1970 & ~n1971 ;
  assign n1972 = ~n460 & ~n480 ;
  assign n1973 = n463 & ~n1972 ;
  assign n1974 = ~n475 & ~n711 ;
  assign n1975 = n478 & ~n1974 ;
  assign n1998 = ~n1973 & ~n1975 ;
  assign n2008 = n1997 & n1998 ;
  assign n2009 = n2007 & n2008 ;
  assign n1990 = ~n339 & ~n373 ;
  assign n1991 = n344 & ~n1990 ;
  assign n1992 = n377 & ~n773 ;
  assign n2003 = ~n1991 & ~n1992 ;
  assign n1993 = ~n420 & ~n450 ;
  assign n1994 = n438 & ~n1993 ;
  assign n1995 = ~n404 & ~n435 ;
  assign n1996 = n488 & ~n1995 ;
  assign n2004 = ~n1994 & ~n1996 ;
  assign n2005 = n2003 & n2004 ;
  assign n1983 = ~n489 & ~n729 ;
  assign n1984 = n392 & ~n1983 ;
  assign n1985 = n306 & ~n771 ;
  assign n2001 = ~n1984 & ~n1985 ;
  assign n1986 = ~n367 & ~n694 ;
  assign n1987 = n443 & ~n1986 ;
  assign n1988 = ~n440 & ~n715 ;
  assign n1989 = n408 & ~n1988 ;
  assign n2002 = ~n1987 & ~n1989 ;
  assign n2006 = n2001 & n2002 ;
  assign n2010 = n2005 & n2006 ;
  assign n2011 = n2009 & n2010 ;
  assign n2012 = \desIn[43]_pad  & n308 ;
  assign n2014 = ~\FP_R_reg[22]/P0001  & n313 ;
  assign n2013 = ~\FP_R_reg[54]/NET0131  & ~n313 ;
  assign n2015 = ~n308 & ~n2013 ;
  assign n2016 = ~n2014 & n2015 ;
  assign n2017 = ~n2012 & ~n2016 ;
  assign n2018 = ~n2011 & n2017 ;
  assign n2019 = n2011 & ~n2017 ;
  assign n2020 = ~n2018 & ~n2019 ;
  assign n2182 = ~n2020 & n2070 ;
  assign n2183 = n1968 & ~n2182 ;
  assign n2185 = n2070 & n2184 ;
  assign n2186 = ~n2183 & ~n2185 ;
  assign n2187 = n2181 & ~n2186 ;
  assign n2127 = n2070 & n2126 ;
  assign n2128 = n2020 & n2127 ;
  assign n2129 = n1968 & n2128 ;
  assign n2193 = \desIn[59]_pad  & n308 ;
  assign n2195 = ~\FP_R_reg[24]/P0001  & n313 ;
  assign n2194 = ~\FP_R_reg[56]/NET0131  & ~n313 ;
  assign n2196 = ~n308 & ~n2194 ;
  assign n2197 = ~n2195 & n2196 ;
  assign n2198 = ~n2193 & ~n2197 ;
  assign n2206 = n377 & ~n486 ;
  assign n2207 = ~n541 & ~n732 ;
  assign n2208 = n448 & ~n2207 ;
  assign n2229 = ~n2206 & ~n2208 ;
  assign n2209 = ~n556 & ~n711 ;
  assign n2210 = n443 & ~n2209 ;
  assign n2211 = ~n340 & n453 ;
  assign n2230 = ~n2210 & ~n2211 ;
  assign n2237 = n2229 & n2230 ;
  assign n2199 = n306 & ~n456 ;
  assign n2200 = ~n549 & ~n600 ;
  assign n2201 = n458 & ~n2200 ;
  assign n2227 = ~n2199 & ~n2201 ;
  assign n2202 = ~n578 & ~n603 ;
  assign n2203 = n488 & ~n2202 ;
  assign n2204 = ~n555 & ~n694 ;
  assign n2205 = n478 & ~n2204 ;
  assign n2228 = ~n2203 & ~n2205 ;
  assign n2238 = n2227 & n2228 ;
  assign n2239 = n2237 & n2238 ;
  assign n2220 = ~n390 & n483 ;
  assign n2221 = ~n527 & ~n729 ;
  assign n2222 = n408 & ~n2221 ;
  assign n2233 = ~n2220 & ~n2222 ;
  assign n2223 = ~n552 & ~n586 ;
  assign n2224 = n423 & ~n2223 ;
  assign n2225 = ~n519 & ~n594 ;
  assign n2226 = n438 & ~n2225 ;
  assign n2234 = ~n2224 & ~n2226 ;
  assign n2235 = n2233 & n2234 ;
  assign n2212 = ~n516 & ~n597 ;
  assign n2213 = n361 & ~n2212 ;
  assign n2214 = ~n567 & ~n723 ;
  assign n2215 = n344 & ~n2214 ;
  assign n2231 = ~n2213 & ~n2215 ;
  assign n2216 = ~n564 & ~n575 ;
  assign n2217 = n463 & ~n2216 ;
  assign n2218 = ~n533 & ~n715 ;
  assign n2219 = n392 & ~n2218 ;
  assign n2232 = ~n2217 & ~n2219 ;
  assign n2236 = n2231 & n2232 ;
  assign n2240 = n2235 & n2236 ;
  assign n2241 = n2239 & n2240 ;
  assign n2242 = n2198 & ~n2241 ;
  assign n2243 = ~n2198 & n2241 ;
  assign n2244 = ~n2242 & ~n2243 ;
  assign n2245 = ~n2129 & ~n2244 ;
  assign n2246 = ~n2187 & n2245 ;
  assign n2247 = ~n2192 & n2246 ;
  assign n2248 = ~n1968 & ~n2070 ;
  assign n2257 = n2126 & n2248 ;
  assign n2258 = n1968 & n2182 ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = n2181 & ~n2259 ;
  assign n2261 = ~n2126 & n2182 ;
  assign n2253 = n1968 & ~n2070 ;
  assign n2254 = ~n2181 & n2253 ;
  assign n2262 = n2244 & ~n2254 ;
  assign n2263 = ~n2261 & n2262 ;
  assign n2249 = n2020 & ~n2126 ;
  assign n2250 = ~n2020 & n2126 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = n2248 & ~n2251 ;
  assign n2255 = n2020 & n2188 ;
  assign n2256 = n2126 & n2255 ;
  assign n2264 = ~n2252 & ~n2256 ;
  assign n2265 = n2263 & n2264 ;
  assign n2266 = ~n2260 & n2265 ;
  assign n2267 = ~n2247 & ~n2266 ;
  assign n2268 = ~n2020 & n2181 ;
  assign n2269 = n2257 & n2268 ;
  assign n2270 = ~n2020 & ~n2181 ;
  assign n2271 = n1968 & ~n2126 ;
  assign n2272 = n2070 & n2271 ;
  assign n2273 = n1968 & n2126 ;
  assign n2274 = ~n2070 & n2273 ;
  assign n2275 = ~n2272 & ~n2274 ;
  assign n2276 = n2270 & ~n2275 ;
  assign n2277 = ~n2269 & ~n2276 ;
  assign n2278 = ~n2267 & n2277 ;
  assign n2279 = ~\desIn[18]_pad  & n308 ;
  assign n2281 = \FP_R_reg[19]/P0001  & ~n313 ;
  assign n2280 = \FP_R_reg[51]/NET0131  & n313 ;
  assign n2282 = ~n308 & ~n2280 ;
  assign n2283 = ~n2281 & n2282 ;
  assign n2284 = ~n2279 & ~n2283 ;
  assign n2285 = n2278 & ~n2284 ;
  assign n2286 = ~n2278 & n2284 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = ~n889 & ~n898 ;
  assign n2289 = ~n816 & ~n2288 ;
  assign n2290 = ~n816 & ~n913 ;
  assign n2291 = ~n888 & ~n891 ;
  assign n2292 = ~n884 & ~n2291 ;
  assign n2293 = ~n2290 & ~n2292 ;
  assign n2294 = ~n2289 & ~n2293 ;
  assign n2295 = ~n510 & ~n2294 ;
  assign n2306 = n685 & n877 ;
  assign n2307 = ~n816 & n2306 ;
  assign n2308 = ~n816 & n873 ;
  assign n2309 = n758 & n817 ;
  assign n2310 = n2308 & n2309 ;
  assign n2318 = ~n2307 & ~n2310 ;
  assign n2319 = ~n2295 & n2318 ;
  assign n2297 = ~n685 & n907 ;
  assign n2298 = n759 & ~n873 ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = ~n816 & ~n2299 ;
  assign n2301 = n816 & n904 ;
  assign n2296 = n888 & n913 ;
  assign n2302 = ~n902 & ~n2296 ;
  assign n2303 = ~n2301 & n2302 ;
  assign n2304 = ~n2300 & n2303 ;
  assign n2305 = n510 & ~n2304 ;
  assign n2314 = ~n873 & n889 ;
  assign n2311 = n873 & n884 ;
  assign n2312 = ~n758 & n817 ;
  assign n2313 = ~n873 & n2312 ;
  assign n2315 = ~n2311 & ~n2313 ;
  assign n2316 = ~n2314 & n2315 ;
  assign n2317 = n816 & ~n2316 ;
  assign n2320 = ~n2305 & ~n2317 ;
  assign n2321 = n2319 & n2320 ;
  assign n2322 = ~\desIn[22]_pad  & n308 ;
  assign n2324 = \FP_R_reg[3]/P0001  & ~n313 ;
  assign n2323 = \FP_R_reg[35]/NET0131  & n313 ;
  assign n2325 = ~n308 & ~n2323 ;
  assign n2326 = ~n2324 & n2325 ;
  assign n2327 = ~n2322 & ~n2326 ;
  assign n2328 = n2321 & ~n2327 ;
  assign n2329 = ~n2321 & n2327 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = \desIn[23]_pad  & n308 ;
  assign n2333 = ~\FP_R_reg[3]/P0001  & n313 ;
  assign n2332 = ~\FP_R_reg[35]/NET0131  & ~n313 ;
  assign n2334 = ~n308 & ~n2332 ;
  assign n2335 = ~n2333 & n2334 ;
  assign n2336 = ~n2331 & ~n2335 ;
  assign n2337 = ~n1682 & n1894 ;
  assign n2338 = n1626 & n2337 ;
  assign n2339 = n1881 & ~n2338 ;
  assign n2340 = n1853 & ~n2339 ;
  assign n2343 = ~n1626 & n1738 ;
  assign n2344 = ~n1879 & ~n2343 ;
  assign n2345 = ~n1795 & ~n1853 ;
  assign n2346 = ~n2344 & n2345 ;
  assign n2341 = ~n1626 & n1860 ;
  assign n2342 = n1682 & n2341 ;
  assign n2347 = ~n1626 & n1853 ;
  assign n2348 = n1795 & n2347 ;
  assign n2349 = n1796 & n1859 ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = ~n2342 & n2350 ;
  assign n2352 = ~n2346 & n2351 ;
  assign n2353 = ~n2340 & n2352 ;
  assign n2354 = ~n1570 & ~n2353 ;
  assign n2355 = n1682 & ~n1796 ;
  assign n2356 = ~n1877 & n2355 ;
  assign n2357 = n1626 & n2356 ;
  assign n2358 = n1863 & n1877 ;
  assign n2359 = ~n2357 & ~n2358 ;
  assign n2360 = n1570 & ~n2359 ;
  assign n2361 = ~n1626 & n1877 ;
  assign n2362 = ~n1797 & ~n1873 ;
  assign n2363 = ~n2361 & n2362 ;
  assign n2364 = n1570 & ~n1853 ;
  assign n2365 = ~n2363 & n2364 ;
  assign n2366 = ~n1885 & ~n2358 ;
  assign n2367 = ~n1853 & ~n2366 ;
  assign n2368 = n1570 & ~n1795 ;
  assign n2369 = n1853 & n2368 ;
  assign n2370 = ~n2344 & n2369 ;
  assign n2371 = ~n2367 & ~n2370 ;
  assign n2372 = ~n2365 & n2371 ;
  assign n2373 = ~n2360 & n2372 ;
  assign n2374 = ~n2354 & n2373 ;
  assign n2375 = ~\desIn[24]_pad  & n308 ;
  assign n2377 = \FP_R_reg[28]/P0001  & ~n313 ;
  assign n2376 = \FP_R_reg[60]/NET0131  & n313 ;
  assign n2378 = ~n308 & ~n2376 ;
  assign n2379 = ~n2377 & n2378 ;
  assign n2380 = ~n2375 & ~n2379 ;
  assign n2381 = n2374 & ~n2380 ;
  assign n2382 = ~n2374 & n2380 ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = \desIn[25]_pad  & n308 ;
  assign n2386 = ~\FP_R_reg[28]/P0001  & n313 ;
  assign n2385 = ~\FP_R_reg[60]/NET0131  & ~n313 ;
  assign n2387 = ~n308 & ~n2385 ;
  assign n2388 = ~n2386 & n2387 ;
  assign n2389 = ~n2384 & ~n2388 ;
  assign n2407 = n1347 & n1459 ;
  assign n2408 = ~n1478 & ~n2407 ;
  assign n2409 = ~n1287 & n1460 ;
  assign n2414 = ~n1486 & ~n2409 ;
  assign n2410 = ~n1346 & n1464 ;
  assign n2411 = n1231 & ~n1287 ;
  assign n2412 = ~n1465 & ~n2411 ;
  assign n2413 = n1450 & ~n2412 ;
  assign n2415 = ~n2410 & ~n2413 ;
  assign n2416 = n2414 & n2415 ;
  assign n2417 = n2408 & n2416 ;
  assign n2418 = n1096 & ~n2417 ;
  assign n2396 = ~n1484 & ~n1489 ;
  assign n2397 = n1476 & ~n2396 ;
  assign n2394 = ~n1287 & n1449 ;
  assign n2395 = n1462 & n2394 ;
  assign n2398 = ~n1483 & ~n2395 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2390 = ~n1287 & n1393 ;
  assign n2391 = ~n1346 & n1485 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = ~n1449 & ~n2392 ;
  assign n2400 = n1470 & ~n2393 ;
  assign n2401 = n2399 & n2400 ;
  assign n2402 = ~n1096 & ~n2401 ;
  assign n2403 = n1455 & n1485 ;
  assign n2404 = ~n1469 & ~n2403 ;
  assign n2405 = n1449 & ~n2404 ;
  assign n2406 = n1451 & n1465 ;
  assign n2419 = ~n1487 & ~n2406 ;
  assign n2420 = ~n2405 & n2419 ;
  assign n2421 = ~n2402 & n2420 ;
  assign n2422 = ~n2418 & n2421 ;
  assign n2423 = ~\desIn[26]_pad  & n308 ;
  assign n2425 = \FP_R_reg[20]/P0001  & ~n313 ;
  assign n2424 = \FP_R_reg[52]/NET0131  & n313 ;
  assign n2426 = ~n308 & ~n2424 ;
  assign n2427 = ~n2425 & n2426 ;
  assign n2428 = ~n2423 & ~n2427 ;
  assign n2429 = n2422 & ~n2428 ;
  assign n2430 = ~n2422 & n2428 ;
  assign n2431 = ~n2429 & ~n2430 ;
  assign n2432 = \desIn[28]_pad  & n308 ;
  assign n2434 = ~\FP_R_reg[44]/NET0131  & n313 ;
  assign n2433 = ~\FP_R_reg[12]/P0001  & ~n313 ;
  assign n2435 = ~n308 & ~n2433 ;
  assign n2436 = ~n2434 & n2435 ;
  assign n2437 = ~n2432 & ~n2436 ;
  assign n2446 = ~n367 & ~n556 ;
  assign n2447 = n408 & ~n2446 ;
  assign n2448 = ~n490 & ~n586 ;
  assign n2449 = n453 & ~n2448 ;
  assign n2472 = ~n2447 & ~n2449 ;
  assign n2450 = ~n469 & ~n600 ;
  assign n2451 = n377 & ~n2450 ;
  assign n2452 = ~n373 & ~n567 ;
  assign n2453 = n392 & ~n2452 ;
  assign n2473 = ~n2451 & ~n2453 ;
  assign n2480 = n2472 & n2473 ;
  assign n2438 = ~n489 & ~n533 ;
  assign n2439 = n344 & ~n2438 ;
  assign n2440 = ~n435 & ~n578 ;
  assign n2441 = n306 & ~n2440 ;
  assign n2470 = ~n2439 & ~n2441 ;
  assign n2442 = ~n444 & ~n479 ;
  assign n2443 = n438 & ~n2442 ;
  assign n2444 = ~n398 & ~n414 ;
  assign n2445 = n361 & ~n2444 ;
  assign n2471 = ~n2443 & ~n2445 ;
  assign n2481 = n2470 & n2471 ;
  assign n2482 = n2480 & n2481 ;
  assign n2462 = ~n429 & ~n484 ;
  assign n2463 = n458 & ~n2462 ;
  assign n2464 = ~n460 & ~n575 ;
  assign n2465 = n483 & ~n2464 ;
  assign n2476 = ~n2463 & ~n2465 ;
  assign n2466 = ~n440 & ~n527 ;
  assign n2467 = n443 & ~n2466 ;
  assign n2468 = ~n350 & ~n454 ;
  assign n2469 = n488 & ~n2468 ;
  assign n2477 = ~n2467 & ~n2469 ;
  assign n2478 = n2476 & n2477 ;
  assign n2454 = ~n333 & ~n459 ;
  assign n2455 = n423 & ~n2454 ;
  assign n2456 = ~n439 & ~n541 ;
  assign n2457 = n478 & ~n2456 ;
  assign n2474 = ~n2455 & ~n2457 ;
  assign n2458 = ~n475 & ~n555 ;
  assign n2459 = n448 & ~n2458 ;
  assign n2460 = ~n383 & ~n449 ;
  assign n2461 = n463 & ~n2460 ;
  assign n2475 = ~n2459 & ~n2461 ;
  assign n2479 = n2474 & n2475 ;
  assign n2483 = n2478 & n2479 ;
  assign n2484 = n2482 & n2483 ;
  assign n2485 = \desIn[17]_pad  & n308 ;
  assign n2487 = ~\FP_R_reg[27]/P0001  & n313 ;
  assign n2486 = ~\FP_R_reg[59]/NET0131  & ~n313 ;
  assign n2488 = ~n308 & ~n2486 ;
  assign n2489 = ~n2487 & n2488 ;
  assign n2490 = ~n2485 & ~n2489 ;
  assign n2491 = n2484 & ~n2490 ;
  assign n2492 = ~n2484 & n2490 ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2502 = ~n367 & ~n445 ;
  assign n2503 = n458 & ~n2502 ;
  assign n2504 = ~n398 & ~n729 ;
  assign n2505 = n483 & ~n2504 ;
  assign n2528 = ~n2503 & ~n2505 ;
  assign n2506 = ~n455 & ~n459 ;
  assign n2507 = n443 & ~n2506 ;
  assign n2508 = ~n475 & ~n480 ;
  assign n2509 = n344 & ~n2508 ;
  assign n2529 = ~n2507 & ~n2509 ;
  assign n2536 = n2528 & n2529 ;
  assign n2494 = ~n414 & ~n715 ;
  assign n2495 = n377 & ~n2494 ;
  assign n2496 = ~n389 & ~n429 ;
  assign n2497 = n408 & ~n2496 ;
  assign n2526 = ~n2495 & ~n2497 ;
  assign n2498 = ~n435 & ~n490 ;
  assign n2499 = n438 & ~n2498 ;
  assign n2500 = ~n479 & ~n711 ;
  assign n2501 = n306 & ~n2500 ;
  assign n2527 = ~n2499 & ~n2501 ;
  assign n2537 = n2526 & n2527 ;
  assign n2538 = n2536 & n2537 ;
  assign n2518 = ~n460 & ~n469 ;
  assign n2519 = n361 & ~n2518 ;
  assign n2520 = ~n404 & ~n489 ;
  assign n2521 = n448 & ~n2520 ;
  assign n2532 = ~n2519 & ~n2521 ;
  assign n2522 = ~n356 & ~n373 ;
  assign n2523 = n463 & ~n2522 ;
  assign n2524 = ~n449 & ~n485 ;
  assign n2525 = n392 & ~n2524 ;
  assign n2533 = ~n2523 & ~n2525 ;
  assign n2534 = n2532 & n2533 ;
  assign n2510 = ~n339 & ~n350 ;
  assign n2511 = n478 & ~n2510 ;
  assign n2512 = ~n420 & ~n440 ;
  assign n2513 = n423 & ~n2512 ;
  assign n2530 = ~n2511 & ~n2513 ;
  assign n2514 = ~n439 & ~n450 ;
  assign n2515 = n488 & ~n2514 ;
  assign n2516 = ~n444 & ~n694 ;
  assign n2517 = n453 & ~n2516 ;
  assign n2531 = ~n2515 & ~n2517 ;
  assign n2535 = n2530 & n2531 ;
  assign n2539 = n2534 & n2535 ;
  assign n2540 = n2538 & n2539 ;
  assign n2541 = n2123 & ~n2540 ;
  assign n2542 = ~n2123 & n2540 ;
  assign n2543 = ~n2541 & ~n2542 ;
  assign n2550 = ~n552 & ~n732 ;
  assign n2551 = n361 & ~n2550 ;
  assign n2552 = n453 & ~n1933 ;
  assign n2574 = ~n2551 & ~n2552 ;
  assign n2553 = ~n404 & ~n586 ;
  assign n2554 = n478 & ~n2553 ;
  assign n2555 = ~n603 & ~n729 ;
  assign n2556 = n463 & ~n2555 ;
  assign n2575 = ~n2554 & ~n2556 ;
  assign n2582 = n2574 & n2575 ;
  assign n2544 = ~n389 & ~n578 ;
  assign n2545 = n443 & ~n2544 ;
  assign n2546 = n377 & ~n1931 ;
  assign n2572 = ~n2545 & ~n2546 ;
  assign n2547 = n483 & ~n1927 ;
  assign n2548 = ~n480 & ~n600 ;
  assign n2549 = n392 & ~n2548 ;
  assign n2573 = ~n2547 & ~n2549 ;
  assign n2583 = n2572 & n2573 ;
  assign n2584 = n2582 & n2583 ;
  assign n2565 = ~n564 & ~n711 ;
  assign n2566 = n488 & ~n2565 ;
  assign n2567 = n306 & ~n1947 ;
  assign n2578 = ~n2566 & ~n2567 ;
  assign n2568 = ~n485 & ~n519 ;
  assign n2569 = n344 & ~n2568 ;
  assign n2570 = ~n597 & ~n694 ;
  assign n2571 = n423 & ~n2570 ;
  assign n2579 = ~n2569 & ~n2571 ;
  assign n2580 = n2578 & n2579 ;
  assign n2557 = ~n594 & ~n715 ;
  assign n2558 = n458 & ~n2557 ;
  assign n2559 = ~n339 & ~n516 ;
  assign n2560 = n448 & ~n2559 ;
  assign n2576 = ~n2558 & ~n2560 ;
  assign n2561 = ~n455 & ~n575 ;
  assign n2562 = n408 & ~n2561 ;
  assign n2563 = ~n549 & ~n723 ;
  assign n2564 = n438 & ~n2563 ;
  assign n2577 = ~n2562 & ~n2564 ;
  assign n2581 = n2576 & n2577 ;
  assign n2585 = n2580 & n2581 ;
  assign n2586 = n2584 & n2585 ;
  assign n2587 = ~n2198 & ~n2586 ;
  assign n2588 = n2198 & n2586 ;
  assign n2589 = ~n2587 & ~n2588 ;
  assign n2590 = n2543 & ~n2589 ;
  assign n2599 = ~n333 & ~n555 ;
  assign n2600 = n361 & ~n2599 ;
  assign n2601 = ~n475 & ~n597 ;
  assign n2602 = n453 & ~n2601 ;
  assign n2625 = ~n2600 & ~n2602 ;
  assign n2603 = ~n414 & ~n586 ;
  assign n2604 = n448 & ~n2603 ;
  assign n2605 = ~n429 & ~n519 ;
  assign n2606 = n392 & ~n2605 ;
  assign n2626 = ~n2604 & ~n2606 ;
  assign n2633 = n2625 & n2626 ;
  assign n2591 = ~n484 & ~n533 ;
  assign n2592 = n438 & ~n2591 ;
  assign n2593 = ~n440 & ~n603 ;
  assign n2594 = n483 & ~n2593 ;
  assign n2623 = ~n2592 & ~n2594 ;
  assign n2595 = ~n444 & ~n600 ;
  assign n2596 = n344 & ~n2595 ;
  assign n2597 = ~n479 & ~n567 ;
  assign n2598 = n458 & ~n2597 ;
  assign n2624 = ~n2596 & ~n2598 ;
  assign n2634 = n2623 & n2624 ;
  assign n2635 = n2633 & n2634 ;
  assign n2615 = ~n454 & ~n556 ;
  assign n2616 = n463 & ~n2615 ;
  assign n2617 = ~n367 & ~n564 ;
  assign n2618 = n306 & ~n2617 ;
  assign n2629 = ~n2616 & ~n2618 ;
  assign n2619 = ~n459 & ~n516 ;
  assign n2620 = n478 & ~n2619 ;
  assign n2621 = ~n383 & ~n527 ;
  assign n2622 = n488 & ~n2621 ;
  assign n2630 = ~n2620 & ~n2622 ;
  assign n2631 = n2629 & n2630 ;
  assign n2607 = ~n398 & ~n541 ;
  assign n2608 = n423 & ~n2607 ;
  assign n2609 = ~n489 & ~n594 ;
  assign n2610 = n377 & ~n2609 ;
  assign n2627 = ~n2608 & ~n2610 ;
  assign n2611 = ~n350 & ~n575 ;
  assign n2612 = n443 & ~n2611 ;
  assign n2613 = ~n449 & ~n578 ;
  assign n2614 = n408 & ~n2613 ;
  assign n2628 = ~n2612 & ~n2614 ;
  assign n2632 = n2627 & n2628 ;
  assign n2636 = n2631 & n2632 ;
  assign n2637 = n2635 & n2636 ;
  assign n2638 = \desIn[9]_pad  & n308 ;
  assign n2640 = ~\FP_R_reg[26]/P0001  & n313 ;
  assign n2639 = ~\FP_R_reg[58]/NET0131  & ~n313 ;
  assign n2641 = ~n308 & ~n2639 ;
  assign n2642 = ~n2640 & n2641 ;
  assign n2643 = ~n2638 & ~n2642 ;
  assign n2644 = n2637 & n2643 ;
  assign n2645 = ~n2637 & ~n2643 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = ~n2543 & n2646 ;
  assign n2654 = ~n460 & ~n711 ;
  assign n2655 = n344 & ~n2654 ;
  assign n2656 = n377 & ~n2593 ;
  assign n2678 = ~n2655 & ~n2656 ;
  assign n2657 = ~n356 & ~n694 ;
  assign n2658 = n458 & ~n2657 ;
  assign n2659 = ~n469 & ~n723 ;
  assign n2660 = n443 & ~n2659 ;
  assign n2679 = ~n2658 & ~n2660 ;
  assign n2686 = n2678 & n2679 ;
  assign n2648 = ~n450 & ~n715 ;
  assign n2649 = n423 & ~n2648 ;
  assign n2650 = n306 & ~n2601 ;
  assign n2676 = ~n2649 & ~n2650 ;
  assign n2651 = n483 & ~n2609 ;
  assign n2652 = ~n455 & ~n480 ;
  assign n2653 = n361 & ~n2652 ;
  assign n2677 = ~n2651 & ~n2653 ;
  assign n2687 = n2676 & n2677 ;
  assign n2688 = n2686 & n2687 ;
  assign n2669 = ~n435 & ~n729 ;
  assign n2670 = n448 & ~n2669 ;
  assign n2671 = n453 & ~n2617 ;
  assign n2682 = ~n2670 & ~n2671 ;
  assign n2672 = ~n439 & ~n552 ;
  assign n2673 = n392 & ~n2672 ;
  assign n2674 = ~n389 & ~n404 ;
  assign n2675 = n438 & ~n2674 ;
  assign n2683 = ~n2673 & ~n2675 ;
  assign n2684 = n2682 & n2683 ;
  assign n2661 = ~n490 & ~n732 ;
  assign n2662 = n408 & ~n2661 ;
  assign n2663 = ~n373 & ~n549 ;
  assign n2664 = n478 & ~n2663 ;
  assign n2680 = ~n2662 & ~n2664 ;
  assign n2665 = ~n339 & ~n445 ;
  assign n2666 = n463 & ~n2665 ;
  assign n2667 = ~n420 & ~n485 ;
  assign n2668 = n488 & ~n2667 ;
  assign n2681 = ~n2666 & ~n2668 ;
  assign n2685 = n2680 & n2681 ;
  assign n2689 = n2684 & n2685 ;
  assign n2690 = n2688 & n2689 ;
  assign n2691 = \desIn[33]_pad  & n308 ;
  assign n2693 = ~\FP_R_reg[29]/P0001  & n313 ;
  assign n2692 = ~\FP_R_reg[61]/NET0131  & ~n313 ;
  assign n2694 = ~n308 & ~n2692 ;
  assign n2695 = ~n2693 & n2694 ;
  assign n2696 = ~n2691 & ~n2695 ;
  assign n2697 = ~n2690 & ~n2696 ;
  assign n2698 = n2690 & n2696 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n2700 = n2589 & n2699 ;
  assign n2701 = n2647 & n2700 ;
  assign n2702 = ~n2590 & ~n2701 ;
  assign n2703 = n2493 & ~n2702 ;
  assign n2752 = ~n2589 & n2699 ;
  assign n2753 = ~n2543 & ~n2646 ;
  assign n2754 = n2752 & n2753 ;
  assign n2704 = n2543 & ~n2646 ;
  assign n2705 = n2700 & n2704 ;
  assign n2712 = ~n404 & ~n449 ;
  assign n2713 = n443 & ~n2712 ;
  assign n2714 = ~n367 & ~n460 ;
  assign n2715 = n488 & ~n2714 ;
  assign n2736 = ~n2713 & ~n2715 ;
  assign n2716 = ~n445 & ~n459 ;
  assign n2717 = n448 & ~n2716 ;
  assign n2718 = ~n420 & ~n429 ;
  assign n2719 = n344 & ~n2718 ;
  assign n2737 = ~n2717 & ~n2719 ;
  assign n2744 = n2736 & n2737 ;
  assign n2706 = n377 & ~n2077 ;
  assign n2707 = ~n435 & ~n440 ;
  assign n2708 = n463 & ~n2707 ;
  assign n2734 = ~n2706 & ~n2708 ;
  assign n2709 = ~n450 & ~n489 ;
  assign n2710 = n458 & ~n2709 ;
  assign n2711 = n453 & ~n2071 ;
  assign n2735 = ~n2710 & ~n2711 ;
  assign n2745 = n2734 & n2735 ;
  assign n2746 = n2744 & n2745 ;
  assign n2727 = ~n389 & ~n414 ;
  assign n2728 = n478 & ~n2727 ;
  assign n2729 = ~n373 & ~n469 ;
  assign n2730 = n438 & ~n2729 ;
  assign n2740 = ~n2728 & ~n2730 ;
  assign n2731 = n483 & ~n2079 ;
  assign n2732 = ~n439 & ~n490 ;
  assign n2733 = n361 & ~n2732 ;
  assign n2741 = ~n2731 & ~n2733 ;
  assign n2742 = n2740 & n2741 ;
  assign n2720 = ~n350 & ~n480 ;
  assign n2721 = n408 & ~n2720 ;
  assign n2722 = ~n356 & ~n475 ;
  assign n2723 = n423 & ~n2722 ;
  assign n2738 = ~n2721 & ~n2723 ;
  assign n2724 = n306 & ~n2095 ;
  assign n2725 = ~n444 & ~n455 ;
  assign n2726 = n392 & ~n2725 ;
  assign n2739 = ~n2724 & ~n2726 ;
  assign n2743 = n2738 & n2739 ;
  assign n2747 = n2742 & n2743 ;
  assign n2748 = n2746 & n2747 ;
  assign n2749 = ~n2389 & n2748 ;
  assign n2750 = n2389 & ~n2748 ;
  assign n2751 = ~n2749 & ~n2750 ;
  assign n2763 = ~n2705 & n2751 ;
  assign n2764 = ~n2754 & n2763 ;
  assign n2755 = ~n2589 & ~n2699 ;
  assign n2756 = ~n2543 & n2755 ;
  assign n2757 = n2646 & n2756 ;
  assign n2758 = n2493 & ~n2543 ;
  assign n2759 = ~n2704 & ~n2758 ;
  assign n2760 = n2589 & ~n2699 ;
  assign n2761 = ~n2647 & n2760 ;
  assign n2762 = n2759 & n2761 ;
  assign n2765 = ~n2757 & ~n2762 ;
  assign n2766 = n2764 & n2765 ;
  assign n2767 = ~n2703 & n2766 ;
  assign n2778 = ~n2647 & ~n2704 ;
  assign n2777 = ~n2752 & ~n2760 ;
  assign n2779 = ~n2590 & n2777 ;
  assign n2780 = n2778 & n2779 ;
  assign n2768 = ~n2543 & n2699 ;
  assign n2769 = n2646 & ~n2768 ;
  assign n2770 = n2493 & ~n2646 ;
  assign n2771 = ~n2589 & ~n2770 ;
  assign n2772 = ~n2769 & n2771 ;
  assign n2781 = ~n2751 & ~n2772 ;
  assign n2773 = ~n2759 & n2760 ;
  assign n2774 = n2543 & ~n2699 ;
  assign n2775 = ~n2768 & ~n2774 ;
  assign n2776 = ~n2493 & ~n2775 ;
  assign n2782 = ~n2773 & ~n2776 ;
  assign n2783 = n2781 & n2782 ;
  assign n2784 = ~n2780 & n2783 ;
  assign n2785 = ~n2767 & ~n2784 ;
  assign n2786 = n2437 & n2785 ;
  assign n2787 = ~n2437 & ~n2785 ;
  assign n2788 = ~n2786 & ~n2787 ;
  assign n2796 = n483 & ~n1603 ;
  assign n2797 = ~n940 & ~n1110 ;
  assign n2798 = n478 & ~n2797 ;
  assign n2819 = ~n2796 & ~n2798 ;
  assign n2799 = ~n1129 & ~n1160 ;
  assign n2800 = n463 & ~n2799 ;
  assign n2801 = n377 & ~n1597 ;
  assign n2820 = ~n2800 & ~n2801 ;
  assign n2827 = n2819 & n2820 ;
  assign n2789 = n453 & ~n1577 ;
  assign n2790 = ~n1071 & ~n1174 ;
  assign n2791 = n443 & ~n2790 ;
  assign n2817 = ~n2789 & ~n2791 ;
  assign n2792 = ~n1199 & ~n1202 ;
  assign n2793 = n438 & ~n2792 ;
  assign n2794 = ~n1063 & ~n1113 ;
  assign n2795 = n392 & ~n2794 ;
  assign n2818 = ~n2793 & ~n2795 ;
  assign n2828 = n2817 & n2818 ;
  assign n2829 = n2827 & n2828 ;
  assign n2810 = n306 & ~n1585 ;
  assign n2811 = ~n1146 & ~n1192 ;
  assign n2812 = n448 & ~n2811 ;
  assign n2823 = ~n2810 & ~n2812 ;
  assign n2813 = ~n1121 & ~n1203 ;
  assign n2814 = n423 & ~n2813 ;
  assign n2815 = ~n1149 & ~n1166 ;
  assign n2816 = n344 & ~n2815 ;
  assign n2824 = ~n2814 & ~n2816 ;
  assign n2825 = n2823 & n2824 ;
  assign n2802 = ~n1018 & ~n1195 ;
  assign n2803 = n408 & ~n2802 ;
  assign n2804 = ~n1135 & ~n1188 ;
  assign n2805 = n361 & ~n2804 ;
  assign n2821 = ~n2803 & ~n2805 ;
  assign n2806 = ~n1191 & ~n1198 ;
  assign n2807 = n488 & ~n2806 ;
  assign n2808 = ~n1152 & ~n1182 ;
  assign n2809 = n458 & ~n2808 ;
  assign n2822 = ~n2807 & ~n2809 ;
  assign n2826 = n2821 & n2822 ;
  assign n2830 = n2825 & n2826 ;
  assign n2831 = n2829 & n2830 ;
  assign n2832 = ~n1745 & ~n2831 ;
  assign n2833 = n1745 & n2831 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2842 = n306 & ~n1715 ;
  assign n2843 = ~n954 & ~n1005 ;
  assign n2844 = n438 & ~n2843 ;
  assign n2865 = ~n2842 & ~n2844 ;
  assign n2845 = ~n1010 & ~n1192 ;
  assign n2846 = n478 & ~n2845 ;
  assign n2847 = ~n960 & ~n1166 ;
  assign n2848 = n392 & ~n2847 ;
  assign n2866 = ~n2846 & ~n2848 ;
  assign n2873 = n2865 & n2866 ;
  assign n2835 = n453 & ~n1689 ;
  assign n2836 = ~n1059 & ~n1063 ;
  assign n2837 = n344 & ~n2836 ;
  assign n2863 = ~n2835 & ~n2837 ;
  assign n2838 = ~n1060 & ~n1075 ;
  assign n2839 = n458 & ~n2838 ;
  assign n2840 = ~n940 & ~n982 ;
  assign n2841 = n448 & ~n2840 ;
  assign n2864 = ~n2839 & ~n2841 ;
  assign n2874 = n2863 & n2864 ;
  assign n2875 = n2873 & n2874 ;
  assign n2856 = ~n968 & ~n988 ;
  assign n2857 = n423 & ~n2856 ;
  assign n2858 = n483 & ~n1697 ;
  assign n2869 = ~n2857 & ~n2858 ;
  assign n2859 = ~n996 & ~n1009 ;
  assign n2860 = n361 & ~n2859 ;
  assign n2861 = ~n1046 & ~n1055 ;
  assign n2862 = n463 & ~n2861 ;
  assign n2870 = ~n2860 & ~n2862 ;
  assign n2871 = n2869 & n2870 ;
  assign n2849 = ~n1032 & ~n1067 ;
  assign n2850 = n488 & ~n2849 ;
  assign n2851 = ~n1038 & ~n1071 ;
  assign n2852 = n408 & ~n2851 ;
  assign n2867 = ~n2850 & ~n2852 ;
  assign n2853 = n377 & ~n1709 ;
  assign n2854 = ~n1018 & ~n1056 ;
  assign n2855 = n443 & ~n2854 ;
  assign n2868 = ~n2853 & ~n2855 ;
  assign n2872 = n2867 & n2868 ;
  assign n2876 = n2871 & n2872 ;
  assign n2877 = n2875 & n2876 ;
  assign n2878 = n2336 & ~n2877 ;
  assign n2879 = ~n2336 & n2877 ;
  assign n2880 = ~n2878 & ~n2879 ;
  assign n2887 = ~n1195 & ~n1203 ;
  assign n2888 = n344 & ~n2887 ;
  assign n2889 = n377 & ~n1659 ;
  assign n2911 = ~n2888 & ~n2889 ;
  assign n2890 = ~n1160 & ~n1188 ;
  assign n2891 = n438 & ~n2890 ;
  assign n2892 = ~n1146 & ~n1198 ;
  assign n2893 = n458 & ~n2892 ;
  assign n2912 = ~n2891 & ~n2893 ;
  assign n2919 = n2911 & n2912 ;
  assign n2881 = ~n1113 & ~n1192 ;
  assign n2882 = n443 & ~n2881 ;
  assign n2883 = n306 & ~n1641 ;
  assign n2909 = ~n2882 & ~n2883 ;
  assign n2884 = n483 & ~n1633 ;
  assign n2885 = ~n1110 & ~n1166 ;
  assign n2886 = n408 & ~n2885 ;
  assign n2910 = ~n2884 & ~n2886 ;
  assign n2920 = n2909 & n2910 ;
  assign n2921 = n2919 & n2920 ;
  assign n2902 = ~n1018 & ~n1102 ;
  assign n2903 = n478 & ~n2902 ;
  assign n2904 = n453 & ~n1653 ;
  assign n2915 = ~n2903 & ~n2904 ;
  assign n2905 = ~n1174 & ~n1182 ;
  assign n2906 = n448 & ~n2905 ;
  assign n2907 = ~n1071 & ~n1138 ;
  assign n2908 = n392 & ~n2907 ;
  assign n2916 = ~n2906 & ~n2908 ;
  assign n2917 = n2915 & n2916 ;
  assign n2894 = ~n1135 & ~n1152 ;
  assign n2895 = n488 & ~n2894 ;
  assign n2896 = ~n1191 & ~n1202 ;
  assign n2897 = n361 & ~n2896 ;
  assign n2913 = ~n2895 & ~n2897 ;
  assign n2898 = ~n1129 & ~n1149 ;
  assign n2899 = n423 & ~n2898 ;
  assign n2900 = ~n1121 & ~n1199 ;
  assign n2901 = n463 & ~n2900 ;
  assign n2914 = ~n2899 & ~n2901 ;
  assign n2918 = n2913 & n2914 ;
  assign n2922 = n2917 & n2918 ;
  assign n2923 = n2921 & n2922 ;
  assign n2924 = \desIn[57]_pad  & n308 ;
  assign n2926 = ~\FP_R_reg[32]/P0001  & n313 ;
  assign n2925 = ~\FP_R_reg[64]/NET0131  & ~n313 ;
  assign n2927 = ~n308 & ~n2925 ;
  assign n2928 = ~n2926 & n2927 ;
  assign n2929 = ~n2924 & ~n2928 ;
  assign n2930 = ~n2923 & n2929 ;
  assign n2931 = n2923 & ~n2929 ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2940 = ~n1002 & ~n1052 ;
  assign n2941 = n438 & ~n2940 ;
  assign n2942 = n377 & ~n1772 ;
  assign n2963 = ~n2941 & ~n2942 ;
  assign n2943 = n483 & ~n1754 ;
  assign n2944 = ~n1060 & ~n1299 ;
  assign n2945 = n408 & ~n2944 ;
  assign n2964 = ~n2943 & ~n2945 ;
  assign n2971 = n2963 & n2964 ;
  assign n2933 = ~n1055 & ~n1102 ;
  assign n2934 = n392 & ~n2933 ;
  assign n2935 = n453 & ~n1746 ;
  assign n2961 = ~n2934 & ~n2935 ;
  assign n2936 = ~n1056 & ~n1064 ;
  assign n2937 = n423 & ~n2936 ;
  assign n2938 = ~n960 & ~n974 ;
  assign n2939 = n463 & ~n2938 ;
  assign n2962 = ~n2937 & ~n2939 ;
  assign n2972 = n2961 & n2962 ;
  assign n2973 = n2971 & n2972 ;
  assign n2954 = ~n982 & ~n1072 ;
  assign n2955 = n344 & ~n2954 ;
  assign n2956 = n306 & ~n1766 ;
  assign n2967 = ~n2955 & ~n2956 ;
  assign n2957 = ~n988 & ~n1306 ;
  assign n2958 = n443 & ~n2957 ;
  assign n2959 = ~n946 & ~n1038 ;
  assign n2960 = n458 & ~n2959 ;
  assign n2968 = ~n2958 & ~n2960 ;
  assign n2969 = n2967 & n2968 ;
  assign n2946 = ~n1032 & ~n1138 ;
  assign n2947 = n478 & ~n2946 ;
  assign n2948 = ~n1010 & ~n1076 ;
  assign n2949 = n488 & ~n2948 ;
  assign n2965 = ~n2947 & ~n2949 ;
  assign n2950 = ~n1024 & ~n1059 ;
  assign n2951 = n448 & ~n2950 ;
  assign n2952 = ~n1006 & ~n1068 ;
  assign n2953 = n361 & ~n2952 ;
  assign n2966 = ~n2951 & ~n2953 ;
  assign n2970 = n2965 & n2966 ;
  assign n2974 = n2969 & n2970 ;
  assign n2975 = n2973 & n2974 ;
  assign n2979 = ~\FP_R_reg[33]/NET0131  & n311 ;
  assign n2978 = ~\FP_R_reg[1]/P0001  & ~n311 ;
  assign n2980 = ~n307 & ~n2978 ;
  assign n2981 = ~n2979 & n2980 ;
  assign n2976 = \FP_R_reg[33]/NET0131  & n312 ;
  assign n2977 = \desIn[7]_pad  & n308 ;
  assign n2982 = ~n2976 & ~n2977 ;
  assign n2983 = ~n2981 & n2982 ;
  assign n2984 = ~n2975 & n2983 ;
  assign n2985 = n2975 & ~n2983 ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n3051 = ~n1010 & ~n1063 ;
  assign n3052 = n408 & ~n3051 ;
  assign n3053 = ~n1076 & ~n1203 ;
  assign n3054 = n483 & ~n3053 ;
  assign n3077 = ~n3052 & ~n3054 ;
  assign n3055 = ~n1009 & ~n1055 ;
  assign n3056 = n438 & ~n3055 ;
  assign n3057 = ~n968 & ~n1038 ;
  assign n3058 = n344 & ~n3057 ;
  assign n3078 = ~n3056 & ~n3058 ;
  assign n3085 = n3077 & n3078 ;
  assign n3043 = ~n954 & ~n1032 ;
  assign n3044 = n361 & ~n3043 ;
  assign n3045 = ~n1002 & ~n1018 ;
  assign n3046 = n392 & ~n3045 ;
  assign n3075 = ~n3044 & ~n3046 ;
  assign n3047 = ~n996 & ~n1060 ;
  assign n3048 = n488 & ~n3047 ;
  assign n3049 = ~n1056 & ~n1075 ;
  assign n3050 = n448 & ~n3049 ;
  assign n3076 = ~n3048 & ~n3050 ;
  assign n3086 = n3075 & n3076 ;
  assign n3087 = n3085 & n3086 ;
  assign n3067 = ~n974 & ~n1182 ;
  assign n3068 = n306 & ~n3067 ;
  assign n3069 = ~n982 & ~n1067 ;
  assign n3070 = n458 & ~n3069 ;
  assign n3081 = ~n3068 & ~n3070 ;
  assign n3071 = ~n940 & ~n960 ;
  assign n3072 = n443 & ~n3071 ;
  assign n3073 = ~n1052 & ~n1192 ;
  assign n3074 = n377 & ~n3073 ;
  assign n3082 = ~n3072 & ~n3074 ;
  assign n3083 = n3081 & n3082 ;
  assign n3059 = ~n988 & ~n1005 ;
  assign n3060 = n463 & ~n3059 ;
  assign n3061 = ~n1006 & ~n1071 ;
  assign n3062 = n478 & ~n3061 ;
  assign n3079 = ~n3060 & ~n3062 ;
  assign n3063 = ~n1046 & ~n1059 ;
  assign n3064 = n423 & ~n3063 ;
  assign n3065 = ~n1068 & ~n1166 ;
  assign n3066 = n453 & ~n3065 ;
  assign n3080 = ~n3064 & ~n3066 ;
  assign n3084 = n3079 & n3080 ;
  assign n3088 = n3083 & n3084 ;
  assign n3089 = n3087 & n3088 ;
  assign n3090 = ~n1918 & ~n3089 ;
  assign n3091 = n1918 & n3089 ;
  assign n3092 = ~n3090 & ~n3091 ;
  assign n3118 = ~n2986 & n3092 ;
  assign n3119 = ~n2932 & ~n3118 ;
  assign n2995 = ~n1005 & ~n1188 ;
  assign n2996 = n443 & ~n2995 ;
  assign n2997 = ~n1055 & ~n1121 ;
  assign n2998 = n377 & ~n2997 ;
  assign n3021 = ~n2996 & ~n2998 ;
  assign n2999 = ~n1018 & ~n1192 ;
  assign n3000 = n438 & ~n2999 ;
  assign n3001 = ~n996 & ~n1202 ;
  assign n3002 = n408 & ~n3001 ;
  assign n3022 = ~n3000 & ~n3002 ;
  assign n3029 = n3021 & n3022 ;
  assign n2987 = ~n968 & ~n1129 ;
  assign n2988 = n458 & ~n2987 ;
  assign n2989 = ~n1060 & ~n1146 ;
  assign n2990 = n483 & ~n2989 ;
  assign n3019 = ~n2988 & ~n2990 ;
  assign n2991 = ~n988 & ~n1149 ;
  assign n2992 = n306 & ~n2991 ;
  assign n2993 = ~n1067 & ~n1135 ;
  assign n2994 = n344 & ~n2993 ;
  assign n3020 = ~n2992 & ~n2994 ;
  assign n3030 = n3019 & n3020 ;
  assign n3031 = n3029 & n3030 ;
  assign n3011 = ~n940 & ~n1182 ;
  assign n3012 = n463 & ~n3011 ;
  assign n3013 = ~n1032 & ~n1152 ;
  assign n3014 = n453 & ~n3013 ;
  assign n3025 = ~n3012 & ~n3014 ;
  assign n3015 = ~n954 & ~n1160 ;
  assign n3016 = n478 & ~n3015 ;
  assign n3017 = ~n1009 & ~n1191 ;
  assign n3018 = n392 & ~n3017 ;
  assign n3026 = ~n3016 & ~n3018 ;
  assign n3027 = n3025 & n3026 ;
  assign n3003 = ~n1071 & ~n1166 ;
  assign n3004 = n361 & ~n3003 ;
  assign n3005 = ~n1046 & ~n1199 ;
  assign n3006 = n448 & ~n3005 ;
  assign n3023 = ~n3004 & ~n3006 ;
  assign n3007 = ~n1063 & ~n1203 ;
  assign n3008 = n488 & ~n3007 ;
  assign n3009 = ~n1075 & ~n1198 ;
  assign n3010 = n423 & ~n3009 ;
  assign n3024 = ~n3008 & ~n3010 ;
  assign n3028 = n3023 & n3024 ;
  assign n3032 = n3027 & n3028 ;
  assign n3033 = n3031 & n3032 ;
  assign n3034 = n1632 & ~n3033 ;
  assign n3035 = ~n1632 & n3033 ;
  assign n3036 = ~n3034 & ~n3035 ;
  assign n3039 = n2932 & n3036 ;
  assign n3120 = n3039 & n3118 ;
  assign n3121 = ~n3119 & ~n3120 ;
  assign n3122 = n2880 & ~n3121 ;
  assign n3123 = n2932 & n3092 ;
  assign n3124 = ~n2880 & ~n3123 ;
  assign n3125 = ~n3119 & n3124 ;
  assign n3109 = n2986 & ~n3092 ;
  assign n3116 = n3036 & n3109 ;
  assign n3093 = n2932 & n2986 ;
  assign n3094 = ~n3036 & n3093 ;
  assign n3117 = n3092 & n3094 ;
  assign n3126 = ~n3116 & ~n3117 ;
  assign n3127 = ~n3125 & n3126 ;
  assign n3128 = ~n3122 & n3127 ;
  assign n3129 = ~n2834 & ~n3128 ;
  assign n3037 = ~n2986 & ~n3036 ;
  assign n3038 = n2932 & n3037 ;
  assign n3040 = n2986 & n3039 ;
  assign n3041 = ~n3038 & ~n3040 ;
  assign n3042 = n2880 & ~n3041 ;
  assign n3095 = ~n2932 & n3036 ;
  assign n3096 = ~n2986 & n3095 ;
  assign n3097 = ~n3094 & ~n3096 ;
  assign n3098 = ~n3092 & ~n3097 ;
  assign n3099 = ~n3042 & ~n3098 ;
  assign n3100 = n2834 & ~n3099 ;
  assign n3101 = n2834 & ~n2880 ;
  assign n3102 = ~n2932 & ~n3036 ;
  assign n3103 = ~n3039 & ~n3102 ;
  assign n3104 = ~n2986 & ~n3103 ;
  assign n3105 = ~n2932 & n3092 ;
  assign n3106 = ~n3036 & n3105 ;
  assign n3107 = ~n3104 & ~n3106 ;
  assign n3108 = n3101 & ~n3107 ;
  assign n3110 = ~n3036 & n3109 ;
  assign n3111 = n2986 & n3092 ;
  assign n3112 = n3036 & n3111 ;
  assign n3113 = ~n3110 & ~n3112 ;
  assign n3114 = n2880 & ~n2932 ;
  assign n3115 = ~n3113 & n3114 ;
  assign n3130 = ~n3108 & ~n3115 ;
  assign n3131 = ~n3100 & n3130 ;
  assign n3132 = ~n3129 & n3131 ;
  assign n3133 = ~\desIn[2]_pad  & n308 ;
  assign n3135 = \FP_R_reg[17]/P0001  & ~n313 ;
  assign n3134 = \FP_R_reg[49]/NET0131  & n313 ;
  assign n3136 = ~n308 & ~n3134 ;
  assign n3137 = ~n3135 & n3136 ;
  assign n3138 = ~n3133 & ~n3137 ;
  assign n3139 = n3132 & ~n3138 ;
  assign n3140 = ~n3132 & n3138 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3148 = n2020 & n2273 ;
  assign n3149 = ~n2070 & n3148 ;
  assign n3150 = ~n1968 & n2250 ;
  assign n3151 = ~n2272 & ~n3150 ;
  assign n3152 = ~n3149 & n3151 ;
  assign n3153 = n2181 & ~n3152 ;
  assign n3142 = n2020 & n2257 ;
  assign n3143 = ~n2185 & ~n3142 ;
  assign n3144 = ~n2181 & ~n3143 ;
  assign n3145 = n2270 & n2273 ;
  assign n3146 = ~n2020 & ~n2070 ;
  assign n3147 = n2271 & n3146 ;
  assign n3154 = ~n3145 & ~n3147 ;
  assign n3155 = ~n3144 & n3154 ;
  assign n3156 = ~n3153 & n3155 ;
  assign n3157 = ~n2244 & ~n3156 ;
  assign n3159 = ~n1968 & ~n2020 ;
  assign n3160 = ~n2261 & ~n3159 ;
  assign n3161 = ~n2181 & ~n3160 ;
  assign n3158 = ~n1968 & n2261 ;
  assign n3162 = n2268 & n2273 ;
  assign n3163 = ~n2128 & ~n3162 ;
  assign n3164 = ~n3158 & n3163 ;
  assign n3165 = ~n3161 & n3164 ;
  assign n3166 = n2244 & ~n3165 ;
  assign n3167 = n2020 & n2181 ;
  assign n3168 = n2191 & ~n2272 ;
  assign n3169 = n3167 & ~n3168 ;
  assign n3171 = ~n2070 & n2271 ;
  assign n3172 = n2070 & n2273 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = n2020 & n3173 ;
  assign n3170 = ~n2020 & ~n2184 ;
  assign n3175 = ~n2181 & ~n3170 ;
  assign n3176 = ~n3174 & n3175 ;
  assign n3177 = ~n3169 & ~n3176 ;
  assign n3178 = ~n3166 & n3177 ;
  assign n3179 = ~n3157 & n3178 ;
  assign n3180 = ~\desIn[30]_pad  & n308 ;
  assign n3182 = \FP_R_reg[4]/P0001  & ~n313 ;
  assign n3181 = \FP_R_reg[36]/NET0131  & n313 ;
  assign n3183 = ~n308 & ~n3181 ;
  assign n3184 = ~n3182 & n3183 ;
  assign n3185 = ~n3180 & ~n3184 ;
  assign n3186 = n3179 & ~n3185 ;
  assign n3187 = ~n3179 & n3185 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3193 = n2020 & n2272 ;
  assign n3202 = n2188 & ~n2249 ;
  assign n3203 = ~n3193 & ~n3202 ;
  assign n3204 = n2181 & ~n3203 ;
  assign n3207 = ~n2182 & n2184 ;
  assign n3208 = ~n3148 & ~n3207 ;
  assign n3209 = ~n2181 & ~n3208 ;
  assign n3205 = n2270 & n2271 ;
  assign n3206 = ~n3149 & ~n3205 ;
  assign n3210 = ~n2252 & n3206 ;
  assign n3211 = ~n3209 & n3210 ;
  assign n3212 = ~n3204 & n3211 ;
  assign n3213 = n2244 & ~n3212 ;
  assign n3189 = ~n2255 & ~n3146 ;
  assign n3190 = ~n2126 & ~n3189 ;
  assign n3191 = n3173 & ~n3190 ;
  assign n3192 = n2181 & ~n3191 ;
  assign n3194 = ~n2020 & ~n2248 ;
  assign n3195 = ~n2271 & n3194 ;
  assign n3196 = ~n3193 & ~n3195 ;
  assign n3197 = ~n2181 & ~n3196 ;
  assign n3198 = ~n3142 & ~n3197 ;
  assign n3199 = ~n3192 & n3198 ;
  assign n3200 = ~n2244 & ~n3199 ;
  assign n3201 = n2127 & n2268 ;
  assign n3214 = ~n3147 & ~n3201 ;
  assign n3215 = ~n3200 & n3214 ;
  assign n3216 = ~n3213 & n3215 ;
  assign n3217 = ~\desIn[32]_pad  & n308 ;
  assign n3219 = \FP_R_reg[29]/P0001  & ~n313 ;
  assign n3218 = \FP_R_reg[61]/NET0131  & n313 ;
  assign n3220 = ~n308 & ~n3218 ;
  assign n3221 = ~n3219 & n3220 ;
  assign n3222 = ~n3217 & ~n3221 ;
  assign n3223 = n3216 & ~n3222 ;
  assign n3224 = ~n3216 & n3222 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3234 = ~n356 & ~n600 ;
  assign n3235 = n453 & ~n3234 ;
  assign n3236 = ~n450 & ~n586 ;
  assign n3237 = n377 & ~n3236 ;
  assign n3260 = ~n3235 & ~n3237 ;
  assign n3238 = ~n485 & ~n603 ;
  assign n3239 = n423 & ~n3238 ;
  assign n3240 = ~n480 & ~n516 ;
  assign n3241 = n443 & ~n3240 ;
  assign n3261 = ~n3239 & ~n3241 ;
  assign n3268 = n3260 & n3261 ;
  assign n3226 = ~n404 & ~n519 ;
  assign n3227 = n408 & ~n3226 ;
  assign n3228 = ~n455 & ~n597 ;
  assign n3229 = n344 & ~n3228 ;
  assign n3258 = ~n3227 & ~n3229 ;
  assign n3230 = ~n445 & ~n575 ;
  assign n3231 = n478 & ~n3230 ;
  assign n3232 = ~n339 & ~n564 ;
  assign n3233 = n458 & ~n3232 ;
  assign n3259 = ~n3231 & ~n3233 ;
  assign n3269 = n3258 & n3259 ;
  assign n3270 = n3268 & n3269 ;
  assign n3250 = ~n389 & ~n594 ;
  assign n3251 = n448 & ~n3250 ;
  assign n3252 = ~n729 & ~n732 ;
  assign n3253 = n438 & ~n3252 ;
  assign n3264 = ~n3251 & ~n3253 ;
  assign n3254 = ~n711 & ~n723 ;
  assign n3255 = n361 & ~n3254 ;
  assign n3256 = ~n549 & ~n694 ;
  assign n3257 = n463 & ~n3256 ;
  assign n3265 = ~n3255 & ~n3257 ;
  assign n3266 = n3264 & n3265 ;
  assign n3242 = ~n460 & ~n567 ;
  assign n3243 = n306 & ~n3242 ;
  assign n3244 = ~n435 & ~n541 ;
  assign n3245 = n483 & ~n3244 ;
  assign n3262 = ~n3243 & ~n3245 ;
  assign n3246 = ~n552 & ~n715 ;
  assign n3247 = n488 & ~n3246 ;
  assign n3248 = ~n420 & ~n578 ;
  assign n3249 = n392 & ~n3248 ;
  assign n3263 = ~n3247 & ~n3249 ;
  assign n3267 = n3262 & n3263 ;
  assign n3271 = n3266 & n3267 ;
  assign n3272 = n3270 & n3271 ;
  assign n3273 = ~n2929 & n3272 ;
  assign n3274 = n2929 & ~n3272 ;
  assign n3275 = ~n3273 & ~n3274 ;
  assign n3284 = ~n356 & ~n460 ;
  assign n3285 = n438 & ~n3284 ;
  assign n3286 = ~n414 & ~n732 ;
  assign n3287 = n306 & ~n3286 ;
  assign n3310 = ~n3285 & ~n3287 ;
  assign n3288 = ~n339 & ~n475 ;
  assign n3289 = n408 & ~n3288 ;
  assign n3290 = ~n485 & ~n489 ;
  assign n3291 = n443 & ~n3290 ;
  assign n3311 = ~n3289 & ~n3291 ;
  assign n3318 = n3310 & n3311 ;
  assign n3276 = ~n389 & ~n440 ;
  assign n3277 = n344 & ~n3276 ;
  assign n3278 = ~n350 & ~n711 ;
  assign n3279 = n377 & ~n3278 ;
  assign n3308 = ~n3277 & ~n3279 ;
  assign n3280 = ~n444 & ~n723 ;
  assign n3281 = n483 & ~n3280 ;
  assign n3282 = ~n404 & ~n439 ;
  assign n3283 = n458 & ~n3282 ;
  assign n3309 = ~n3281 & ~n3283 ;
  assign n3319 = n3308 & n3309 ;
  assign n3320 = n3318 & n3319 ;
  assign n3300 = ~n429 & ~n715 ;
  assign n3301 = n478 & ~n3300 ;
  assign n3302 = ~n449 & ~n729 ;
  assign n3303 = n453 & ~n3302 ;
  assign n3314 = ~n3301 & ~n3303 ;
  assign n3304 = ~n445 & ~n469 ;
  assign n3305 = n488 & ~n3304 ;
  assign n3306 = ~n420 & ~n490 ;
  assign n3307 = n463 & ~n3306 ;
  assign n3315 = ~n3305 & ~n3307 ;
  assign n3316 = n3314 & n3315 ;
  assign n3292 = ~n435 & ~n450 ;
  assign n3293 = n361 & ~n3292 ;
  assign n3294 = ~n459 & ~n694 ;
  assign n3295 = n392 & ~n3294 ;
  assign n3312 = ~n3293 & ~n3295 ;
  assign n3296 = ~n373 & ~n480 ;
  assign n3297 = n423 & ~n3296 ;
  assign n3298 = ~n367 & ~n455 ;
  assign n3299 = n448 & ~n3298 ;
  assign n3313 = ~n3297 & ~n3299 ;
  assign n3317 = n3312 & n3313 ;
  assign n3321 = n3316 & n3317 ;
  assign n3322 = n3320 & n3321 ;
  assign n3323 = \desIn[49]_pad  & n308 ;
  assign n3325 = ~\FP_R_reg[31]/P0001  & n313 ;
  assign n3324 = ~\FP_R_reg[63]/NET0131  & ~n313 ;
  assign n3326 = ~n308 & ~n3324 ;
  assign n3327 = ~n3325 & n3326 ;
  assign n3328 = ~n3323 & ~n3327 ;
  assign n3329 = n3322 & ~n3328 ;
  assign n3330 = ~n3322 & n3328 ;
  assign n3331 = ~n3329 & ~n3330 ;
  assign n3439 = ~n383 & ~n420 ;
  assign n3440 = n478 & ~n3439 ;
  assign n3441 = ~n389 & ~n533 ;
  assign n3442 = n306 & ~n3441 ;
  assign n3465 = ~n3440 & ~n3442 ;
  assign n3443 = ~n445 & ~n454 ;
  assign n3444 = n392 & ~n3443 ;
  assign n3445 = ~n449 & ~n490 ;
  assign n3446 = n458 & ~n3445 ;
  assign n3466 = ~n3444 & ~n3446 ;
  assign n3473 = n3465 & n3466 ;
  assign n3431 = ~n356 & ~n479 ;
  assign n3432 = n408 & ~n3431 ;
  assign n3433 = ~n455 & ~n555 ;
  assign n3434 = n483 & ~n3433 ;
  assign n3463 = ~n3432 & ~n3434 ;
  assign n3435 = ~n404 & ~n484 ;
  assign n3436 = n453 & ~n3435 ;
  assign n3437 = ~n440 & ~n489 ;
  assign n3438 = n361 & ~n3437 ;
  assign n3464 = ~n3436 & ~n3438 ;
  assign n3474 = n3463 & n3464 ;
  assign n3475 = n3473 & n3474 ;
  assign n3455 = ~n414 & ~n435 ;
  assign n3456 = n344 & ~n3455 ;
  assign n3457 = ~n333 & ~n480 ;
  assign n3458 = n377 & ~n3457 ;
  assign n3469 = ~n3456 & ~n3458 ;
  assign n3459 = ~n444 & ~n460 ;
  assign n3460 = n448 & ~n3459 ;
  assign n3461 = ~n350 & ~n469 ;
  assign n3462 = n423 & ~n3461 ;
  assign n3470 = ~n3460 & ~n3462 ;
  assign n3471 = n3469 & n3470 ;
  assign n3447 = ~n367 & ~n475 ;
  assign n3448 = n438 & ~n3447 ;
  assign n3449 = ~n429 & ~n439 ;
  assign n3450 = n463 & ~n3449 ;
  assign n3467 = ~n3448 & ~n3450 ;
  assign n3451 = ~n373 & ~n459 ;
  assign n3452 = n488 & ~n3451 ;
  assign n3453 = ~n398 & ~n450 ;
  assign n3454 = n443 & ~n3453 ;
  assign n3468 = ~n3452 & ~n3454 ;
  assign n3472 = n3467 & n3468 ;
  assign n3476 = n3471 & n3472 ;
  assign n3477 = n3475 & n3476 ;
  assign n3478 = ~n2983 & ~n3477 ;
  assign n3479 = n2983 & n3477 ;
  assign n3480 = ~n3478 & ~n3479 ;
  assign n3338 = ~n454 & ~n564 ;
  assign n3339 = n408 & ~n3338 ;
  assign n3340 = n377 & ~n3280 ;
  assign n3362 = ~n3339 & ~n3340 ;
  assign n3341 = ~n567 & ~n600 ;
  assign n3342 = n438 & ~n3341 ;
  assign n3343 = ~n519 & ~n533 ;
  assign n3344 = n458 & ~n3343 ;
  assign n3363 = ~n3342 & ~n3344 ;
  assign n3370 = n3362 & n3363 ;
  assign n3332 = ~n383 & ~n603 ;
  assign n3333 = n443 & ~n3332 ;
  assign n3334 = n306 & ~n3302 ;
  assign n3360 = ~n3333 & ~n3334 ;
  assign n3335 = n483 & ~n3278 ;
  assign n3336 = ~n484 & ~n594 ;
  assign n3337 = n344 & ~n3336 ;
  assign n3361 = ~n3335 & ~n3337 ;
  assign n3371 = n3360 & n3361 ;
  assign n3372 = n3370 & n3371 ;
  assign n3353 = ~n516 & ~n555 ;
  assign n3354 = n423 & ~n3353 ;
  assign n3355 = n453 & ~n3286 ;
  assign n3366 = ~n3354 & ~n3355 ;
  assign n3356 = ~n527 & ~n578 ;
  assign n3357 = n463 & ~n3356 ;
  assign n3358 = ~n398 & ~n552 ;
  assign n3359 = n478 & ~n3358 ;
  assign n3367 = ~n3357 & ~n3359 ;
  assign n3368 = n3366 & n3367 ;
  assign n3345 = ~n541 & ~n586 ;
  assign n3346 = n361 & ~n3345 ;
  assign n3347 = ~n479 & ~n549 ;
  assign n3348 = n392 & ~n3347 ;
  assign n3364 = ~n3346 & ~n3348 ;
  assign n3349 = ~n556 & ~n575 ;
  assign n3350 = n488 & ~n3349 ;
  assign n3351 = ~n333 & ~n597 ;
  assign n3352 = n448 & ~n3351 ;
  assign n3365 = ~n3350 & ~n3352 ;
  assign n3369 = n3364 & n3365 ;
  assign n3373 = n3368 & n3369 ;
  assign n3374 = n3372 & n3373 ;
  assign n3375 = \desIn[41]_pad  & n308 ;
  assign n3377 = ~\FP_R_reg[30]/P0001  & n313 ;
  assign n3376 = ~\FP_R_reg[62]/NET0131  & ~n313 ;
  assign n3378 = ~n308 & ~n3376 ;
  assign n3379 = ~n3377 & n3378 ;
  assign n3380 = ~n3375 & ~n3379 ;
  assign n3381 = n3374 & ~n3380 ;
  assign n3382 = ~n3374 & n3380 ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3391 = ~n455 & ~n549 ;
  assign n3392 = n423 & ~n3391 ;
  assign n3393 = n453 & ~n2440 ;
  assign n3414 = ~n3392 & ~n3393 ;
  assign n3394 = ~n715 & ~n729 ;
  assign n3395 = n361 & ~n3394 ;
  assign n3396 = ~n450 & ~n519 ;
  assign n3397 = n478 & ~n3396 ;
  assign n3415 = ~n3395 & ~n3397 ;
  assign n3422 = n3414 & n3415 ;
  assign n3384 = ~n356 & ~n516 ;
  assign n3385 = n392 & ~n3384 ;
  assign n3386 = n306 & ~n2448 ;
  assign n3412 = ~n3385 & ~n3386 ;
  assign n3387 = ~n404 & ~n603 ;
  assign n3388 = n344 & ~n3387 ;
  assign n3389 = ~n339 & ~n723 ;
  assign n3390 = n488 & ~n3389 ;
  assign n3413 = ~n3388 & ~n3390 ;
  assign n3423 = n3412 & n3413 ;
  assign n3424 = n3422 & n3423 ;
  assign n3405 = ~n480 & ~n564 ;
  assign n3406 = n448 & ~n3405 ;
  assign n3407 = n483 & ~n2450 ;
  assign n3418 = ~n3406 & ~n3407 ;
  assign n3408 = ~n389 & ~n552 ;
  assign n3409 = n458 & ~n3408 ;
  assign n3410 = ~n445 & ~n597 ;
  assign n3411 = n408 & ~n3410 ;
  assign n3419 = ~n3409 & ~n3411 ;
  assign n3420 = n3418 & n3419 ;
  assign n3398 = ~n420 & ~n594 ;
  assign n3399 = n443 & ~n3398 ;
  assign n3400 = n377 & ~n2464 ;
  assign n3416 = ~n3399 & ~n3400 ;
  assign n3401 = ~n694 & ~n711 ;
  assign n3402 = n438 & ~n3401 ;
  assign n3403 = ~n485 & ~n732 ;
  assign n3404 = n463 & ~n3403 ;
  assign n3417 = ~n3402 & ~n3404 ;
  assign n3421 = n3416 & n3417 ;
  assign n3425 = n3420 & n3421 ;
  assign n3426 = n3424 & n3425 ;
  assign n3427 = ~n2696 & n3426 ;
  assign n3428 = n2696 & ~n3426 ;
  assign n3429 = ~n3427 & ~n3428 ;
  assign n3533 = ~n3383 & ~n3429 ;
  assign n3534 = ~n3480 & n3533 ;
  assign n3488 = ~n594 & ~n603 ;
  assign n3489 = n361 & ~n3488 ;
  assign n3490 = n453 & ~n3441 ;
  assign n3511 = ~n3489 & ~n3490 ;
  assign n3491 = ~n485 & ~n527 ;
  assign n3492 = n478 & ~n3491 ;
  assign n3493 = ~n339 & ~n556 ;
  assign n3494 = n392 & ~n3493 ;
  assign n3512 = ~n3492 & ~n3494 ;
  assign n3519 = n3511 & n3512 ;
  assign n3481 = ~n564 & ~n597 ;
  assign n3482 = n438 & ~n3481 ;
  assign n3483 = n483 & ~n3457 ;
  assign n3509 = ~n3482 & ~n3483 ;
  assign n3484 = ~n516 & ~n549 ;
  assign n3485 = n488 & ~n3484 ;
  assign n3486 = ~n575 & ~n723 ;
  assign n3487 = n423 & ~n3486 ;
  assign n3510 = ~n3485 & ~n3487 ;
  assign n3520 = n3509 & n3510 ;
  assign n3521 = n3519 & n3520 ;
  assign n3502 = ~n586 & ~n729 ;
  assign n3503 = n344 & ~n3502 ;
  assign n3504 = n377 & ~n3433 ;
  assign n3515 = ~n3503 & ~n3504 ;
  assign n3505 = ~n541 & ~n715 ;
  assign n3506 = n443 & ~n3505 ;
  assign n3507 = ~n578 & ~n732 ;
  assign n3508 = n458 & ~n3507 ;
  assign n3516 = ~n3506 & ~n3508 ;
  assign n3517 = n3515 & n3516 ;
  assign n3495 = ~n567 & ~n694 ;
  assign n3496 = n408 & ~n3495 ;
  assign n3497 = n306 & ~n3435 ;
  assign n3513 = ~n3496 & ~n3497 ;
  assign n3498 = ~n519 & ~n552 ;
  assign n3499 = n463 & ~n3498 ;
  assign n3500 = ~n600 & ~n711 ;
  assign n3501 = n448 & ~n3500 ;
  assign n3514 = ~n3499 & ~n3501 ;
  assign n3518 = n3513 & n3514 ;
  assign n3522 = n3517 & n3518 ;
  assign n3523 = n3521 & n3522 ;
  assign n3524 = ~n2389 & n3523 ;
  assign n3525 = n2389 & ~n3523 ;
  assign n3526 = ~n3524 & ~n3525 ;
  assign n3535 = n3480 & ~n3526 ;
  assign n3529 = ~n3383 & n3526 ;
  assign n3536 = n3429 & ~n3529 ;
  assign n3537 = ~n3535 & n3536 ;
  assign n3538 = ~n3534 & ~n3537 ;
  assign n3539 = n3331 & ~n3538 ;
  assign n3540 = ~n3429 & n3535 ;
  assign n3541 = n3480 & n3526 ;
  assign n3542 = n3429 & n3541 ;
  assign n3543 = ~n3540 & ~n3542 ;
  assign n3544 = n3383 & ~n3543 ;
  assign n3430 = n3383 & ~n3429 ;
  assign n3527 = ~n3480 & n3526 ;
  assign n3528 = n3430 & n3527 ;
  assign n3530 = n3480 & n3529 ;
  assign n3531 = ~n3528 & ~n3530 ;
  assign n3532 = ~n3331 & ~n3531 ;
  assign n3545 = ~n3526 & n3534 ;
  assign n3546 = ~n3532 & ~n3545 ;
  assign n3547 = ~n3544 & n3546 ;
  assign n3548 = ~n3539 & n3547 ;
  assign n3549 = n3275 & ~n3548 ;
  assign n3550 = n3430 & n3526 ;
  assign n3551 = ~n3542 & ~n3550 ;
  assign n3552 = n3331 & ~n3551 ;
  assign n3553 = n3383 & ~n3526 ;
  assign n3554 = n3429 & n3553 ;
  assign n3555 = n3429 & n3480 ;
  assign n3556 = ~n3331 & ~n3526 ;
  assign n3557 = n3555 & n3556 ;
  assign n3567 = ~n3554 & ~n3557 ;
  assign n3563 = n3533 & n3535 ;
  assign n3564 = ~n3480 & ~n3526 ;
  assign n3565 = ~n3331 & n3383 ;
  assign n3566 = n3564 & n3565 ;
  assign n3568 = ~n3563 & ~n3566 ;
  assign n3569 = n3567 & n3568 ;
  assign n3558 = n3480 & n3550 ;
  assign n3559 = ~n3331 & ~n3383 ;
  assign n3560 = ~n3383 & n3429 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = n3527 & ~n3561 ;
  assign n3570 = ~n3558 & ~n3562 ;
  assign n3571 = n3569 & n3570 ;
  assign n3572 = ~n3552 & n3571 ;
  assign n3573 = ~n3275 & ~n3572 ;
  assign n3574 = ~n3526 & n3533 ;
  assign n3575 = n3331 & n3574 ;
  assign n3576 = n3429 & n3527 ;
  assign n3577 = n3559 & n3576 ;
  assign n3578 = ~n3575 & ~n3577 ;
  assign n3579 = ~n3573 & n3578 ;
  assign n3580 = ~n3549 & n3579 ;
  assign n3581 = ~\desIn[34]_pad  & n308 ;
  assign n3583 = \FP_R_reg[21]/P0001  & ~n313 ;
  assign n3582 = \FP_R_reg[53]/NET0131  & n313 ;
  assign n3584 = ~n308 & ~n3582 ;
  assign n3585 = ~n3583 & n3584 ;
  assign n3586 = ~n3581 & ~n3585 ;
  assign n3587 = n3580 & ~n3586 ;
  assign n3588 = ~n3580 & n3586 ;
  assign n3589 = ~n3587 & ~n3588 ;
  assign n3590 = ~n3529 & ~n3555 ;
  assign n3591 = n3429 & n3530 ;
  assign n3592 = ~n3590 & ~n3591 ;
  assign n3593 = n3331 & ~n3592 ;
  assign n3594 = ~n3331 & ~n3550 ;
  assign n3595 = ~n3574 & n3594 ;
  assign n3596 = ~n3593 & ~n3595 ;
  assign n3597 = n3429 & n3564 ;
  assign n3598 = n3383 & n3597 ;
  assign n3599 = ~n3596 & ~n3598 ;
  assign n3600 = n3275 & ~n3599 ;
  assign n3601 = ~n3429 & ~n3480 ;
  assign n3602 = ~n3526 & n3601 ;
  assign n3603 = ~n3558 & ~n3602 ;
  assign n3604 = ~n3275 & ~n3603 ;
  assign n3605 = ~n3541 & ~n3560 ;
  assign n3606 = ~n3590 & n3605 ;
  assign n3607 = n3553 & n3601 ;
  assign n3608 = ~n3563 & ~n3607 ;
  assign n3609 = ~n3606 & n3608 ;
  assign n3610 = ~n3604 & n3609 ;
  assign n3611 = n3331 & ~n3610 ;
  assign n3615 = n3480 & ~n3553 ;
  assign n3616 = ~n3331 & ~n3601 ;
  assign n3617 = ~n3615 & n3616 ;
  assign n3612 = n3331 & ~n3555 ;
  assign n3613 = n3529 & ~n3612 ;
  assign n3614 = n3383 & n3576 ;
  assign n3618 = ~n3613 & ~n3614 ;
  assign n3619 = ~n3617 & n3618 ;
  assign n3620 = ~n3275 & ~n3619 ;
  assign n3621 = n3542 & n3559 ;
  assign n3622 = ~n3620 & ~n3621 ;
  assign n3623 = ~n3611 & n3622 ;
  assign n3624 = ~n3600 & n3623 ;
  assign n3625 = ~\desIn[38]_pad  & n308 ;
  assign n3627 = \FP_R_reg[5]/P0001  & ~n313 ;
  assign n3626 = \FP_R_reg[37]/NET0131  & n313 ;
  assign n3628 = ~n308 & ~n3626 ;
  assign n3629 = ~n3627 & n3628 ;
  assign n3630 = ~n3625 & ~n3629 ;
  assign n3631 = n3624 & ~n3630 ;
  assign n3632 = ~n3624 & n3630 ;
  assign n3633 = ~n3631 & ~n3632 ;
  assign n3641 = ~n960 & ~n1138 ;
  assign n3642 = n344 & ~n3641 ;
  assign n3643 = n453 & ~n2991 ;
  assign n3664 = ~n3642 & ~n3643 ;
  assign n3644 = n483 & ~n2997 ;
  assign n3645 = ~n1064 & ~n1076 ;
  assign n3646 = n438 & ~n3645 ;
  assign n3665 = ~n3644 & ~n3646 ;
  assign n3672 = n3664 & n3665 ;
  assign n3634 = ~n1056 & ~n1113 ;
  assign n3635 = n408 & ~n3634 ;
  assign n3636 = n306 & ~n3013 ;
  assign n3662 = ~n3635 & ~n3636 ;
  assign n3637 = ~n982 & ~n1174 ;
  assign n3638 = n478 & ~n3637 ;
  assign n3639 = ~n1038 & ~n1110 ;
  assign n3640 = n443 & ~n3639 ;
  assign n3663 = ~n3638 & ~n3640 ;
  assign n3673 = n3662 & n3663 ;
  assign n3674 = n3672 & n3673 ;
  assign n3655 = ~n1024 & ~n1052 ;
  assign n3656 = n488 & ~n3655 ;
  assign n3657 = n377 & ~n2989 ;
  assign n3668 = ~n3656 & ~n3657 ;
  assign n3658 = ~n1059 & ~n1195 ;
  assign n3659 = n392 & ~n3658 ;
  assign n3660 = ~n1010 & ~n1102 ;
  assign n3661 = n448 & ~n3660 ;
  assign n3669 = ~n3659 & ~n3661 ;
  assign n3670 = n3668 & n3669 ;
  assign n3647 = ~n1006 & ~n1306 ;
  assign n3648 = n458 & ~n3647 ;
  assign n3649 = ~n946 & ~n974 ;
  assign n3650 = n361 & ~n3649 ;
  assign n3666 = ~n3648 & ~n3650 ;
  assign n3651 = ~n1068 & ~n1072 ;
  assign n3652 = n463 & ~n3651 ;
  assign n3653 = ~n1002 & ~n1299 ;
  assign n3654 = n423 & ~n3653 ;
  assign n3667 = ~n3652 & ~n3654 ;
  assign n3671 = n3666 & n3667 ;
  assign n3675 = n3670 & n3671 ;
  assign n3676 = n3674 & n3675 ;
  assign n3677 = n1688 & n3676 ;
  assign n3678 = ~n1688 & ~n3676 ;
  assign n3679 = ~n3677 & ~n3678 ;
  assign n3688 = ~n1056 & ~n1199 ;
  assign n3689 = n306 & ~n3688 ;
  assign n3690 = ~n1138 & ~n1306 ;
  assign n3691 = n438 & ~n3690 ;
  assign n3714 = ~n3689 & ~n3691 ;
  assign n3692 = ~n1038 & ~n1135 ;
  assign n3693 = n483 & ~n3692 ;
  assign n3694 = ~n1052 & ~n1121 ;
  assign n3695 = n443 & ~n3694 ;
  assign n3715 = ~n3693 & ~n3695 ;
  assign n3722 = n3714 & n3715 ;
  assign n3680 = ~n960 & ~n1188 ;
  assign n3681 = n377 & ~n3680 ;
  assign n3682 = ~n1068 & ~n1152 ;
  assign n3683 = n408 & ~n3682 ;
  assign n3712 = ~n3681 & ~n3683 ;
  assign n3684 = ~n1076 & ~n1146 ;
  assign n3685 = n344 & ~n3684 ;
  assign n3686 = ~n1064 & ~n1195 ;
  assign n3687 = n458 & ~n3686 ;
  assign n3713 = ~n3685 & ~n3687 ;
  assign n3723 = n3712 & n3713 ;
  assign n3724 = n3722 & n3723 ;
  assign n3704 = ~n1072 & ~n1110 ;
  assign n3705 = n488 & ~n3704 ;
  assign n3706 = ~n1010 & ~n1202 ;
  assign n3707 = n453 & ~n3706 ;
  assign n3718 = ~n3705 & ~n3707 ;
  assign n3708 = ~n974 & ~n1149 ;
  assign n3709 = n448 & ~n3708 ;
  assign n3710 = ~n946 & ~n1174 ;
  assign n3711 = n423 & ~n3710 ;
  assign n3719 = ~n3709 & ~n3711 ;
  assign n3720 = n3718 & n3719 ;
  assign n3696 = ~n1002 & ~n1191 ;
  assign n3697 = n478 & ~n3696 ;
  assign n3698 = ~n1024 & ~n1113 ;
  assign n3699 = n463 & ~n3698 ;
  assign n3716 = ~n3697 & ~n3699 ;
  assign n3700 = ~n1102 & ~n1299 ;
  assign n3701 = n361 & ~n3700 ;
  assign n3702 = ~n1006 & ~n1160 ;
  assign n3703 = n392 & ~n3702 ;
  assign n3717 = ~n3701 & ~n3703 ;
  assign n3721 = n3716 & n3717 ;
  assign n3725 = n3720 & n3721 ;
  assign n3726 = n3724 & n3725 ;
  assign n3727 = n1284 & n3726 ;
  assign n3728 = ~n1284 & ~n3726 ;
  assign n3729 = ~n3727 & ~n3728 ;
  assign n3730 = ~n3679 & n3729 ;
  assign n3739 = ~n1102 & ~n1199 ;
  assign n3740 = n344 & ~n3739 ;
  assign n3741 = ~n974 & ~n1071 ;
  assign n3742 = n483 & ~n3741 ;
  assign n3765 = ~n3740 & ~n3742 ;
  assign n3743 = ~n1129 & ~n1306 ;
  assign n3744 = n408 & ~n3743 ;
  assign n3745 = ~n1113 & ~n1202 ;
  assign n3746 = n458 & ~n3745 ;
  assign n3766 = ~n3744 & ~n3746 ;
  assign n3773 = n3765 & n3766 ;
  assign n3731 = ~n1135 & ~n1138 ;
  assign n3732 = n448 & ~n3731 ;
  assign n3733 = ~n946 & ~n1166 ;
  assign n3734 = n377 & ~n3733 ;
  assign n3763 = ~n3732 & ~n3734 ;
  assign n3735 = ~n1018 & ~n1076 ;
  assign n3736 = n306 & ~n3735 ;
  assign n3737 = ~n1024 & ~n1203 ;
  assign n3738 = n478 & ~n3737 ;
  assign n3764 = ~n3736 & ~n3738 ;
  assign n3774 = n3763 & n3764 ;
  assign n3775 = n3773 & n3774 ;
  assign n3755 = ~n1198 & ~n1299 ;
  assign n3756 = n443 & ~n3755 ;
  assign n3757 = ~n1064 & ~n1192 ;
  assign n3758 = n453 & ~n3757 ;
  assign n3769 = ~n3756 & ~n3758 ;
  assign n3759 = ~n1121 & ~n1146 ;
  assign n3760 = n361 & ~n3759 ;
  assign n3761 = ~n1072 & ~n1182 ;
  assign n3762 = n392 & ~n3761 ;
  assign n3770 = ~n3760 & ~n3762 ;
  assign n3771 = n3769 & n3770 ;
  assign n3747 = ~n1160 & ~n1174 ;
  assign n3748 = n488 & ~n3747 ;
  assign n3749 = ~n1110 & ~n1188 ;
  assign n3750 = n423 & ~n3749 ;
  assign n3767 = ~n3748 & ~n3750 ;
  assign n3751 = ~n1191 & ~n1195 ;
  assign n3752 = n463 & ~n3751 ;
  assign n3753 = ~n1149 & ~n1152 ;
  assign n3754 = n438 & ~n3753 ;
  assign n3768 = ~n3752 & ~n3754 ;
  assign n3772 = n3767 & n3768 ;
  assign n3776 = n3771 & n3772 ;
  assign n3777 = n3775 & n3776 ;
  assign n3778 = ~n1518 & n3777 ;
  assign n3779 = n1518 & ~n3777 ;
  assign n3780 = ~n3778 & ~n3779 ;
  assign n3889 = n3730 & n3780 ;
  assign n3789 = ~n1102 & ~n1113 ;
  assign n3790 = n438 & ~n3789 ;
  assign n3791 = ~n960 & ~n1129 ;
  assign n3792 = n306 & ~n3791 ;
  assign n3815 = ~n3790 & ~n3792 ;
  assign n3793 = ~n1010 & ~n1198 ;
  assign n3794 = n483 & ~n3793 ;
  assign n3795 = ~n1076 & ~n1191 ;
  assign n3796 = n408 & ~n3795 ;
  assign n3816 = ~n3794 & ~n3796 ;
  assign n3823 = n3815 & n3816 ;
  assign n3781 = ~n1195 & ~n1299 ;
  assign n3782 = n488 & ~n3781 ;
  assign n3783 = ~n1006 & ~n1135 ;
  assign n3784 = n453 & ~n3783 ;
  assign n3813 = ~n3782 & ~n3784 ;
  assign n3785 = ~n1174 & ~n1306 ;
  assign n3786 = n463 & ~n3785 ;
  assign n3787 = ~n1064 & ~n1121 ;
  assign n3788 = n448 & ~n3787 ;
  assign n3814 = ~n3786 & ~n3788 ;
  assign n3824 = n3813 & n3814 ;
  assign n3825 = n3823 & n3824 ;
  assign n3805 = ~n1110 & ~n1138 ;
  assign n3806 = n361 & ~n3805 ;
  assign n3807 = ~n1052 & ~n1202 ;
  assign n3808 = n392 & ~n3807 ;
  assign n3819 = ~n3806 & ~n3808 ;
  assign n3809 = ~n1024 & ~n1146 ;
  assign n3810 = n423 & ~n3809 ;
  assign n3811 = ~n1068 & ~n1188 ;
  assign n3812 = n478 & ~n3811 ;
  assign n3820 = ~n3810 & ~n3812 ;
  assign n3821 = n3819 & n3820 ;
  assign n3797 = ~n946 & ~n1152 ;
  assign n3798 = n344 & ~n3797 ;
  assign n3799 = ~n974 & ~n1160 ;
  assign n3800 = n443 & ~n3799 ;
  assign n3817 = ~n3798 & ~n3800 ;
  assign n3801 = ~n1072 & ~n1149 ;
  assign n3802 = n458 & ~n3801 ;
  assign n3803 = ~n1002 & ~n1199 ;
  assign n3804 = n377 & ~n3803 ;
  assign n3818 = ~n3802 & ~n3804 ;
  assign n3822 = n3817 & n3818 ;
  assign n3826 = n3821 & n3822 ;
  assign n3827 = n3825 & n3826 ;
  assign n3828 = n1524 & n3827 ;
  assign n3829 = ~n1524 & ~n3827 ;
  assign n3830 = ~n3828 & ~n3829 ;
  assign n3831 = n3780 & ~n3830 ;
  assign n3832 = ~n3730 & ~n3831 ;
  assign n3841 = ~n946 & ~n1006 ;
  assign n3842 = n488 & ~n3841 ;
  assign n3843 = ~n1002 & ~n1064 ;
  assign n3844 = n463 & ~n3843 ;
  assign n3867 = ~n3842 & ~n3844 ;
  assign n3845 = ~n974 & ~n1068 ;
  assign n3846 = n438 & ~n3845 ;
  assign n3847 = ~n1038 & ~n1306 ;
  assign n3848 = n448 & ~n3847 ;
  assign n3868 = ~n3846 & ~n3848 ;
  assign n3875 = n3867 & n3868 ;
  assign n3833 = ~n954 & ~n1149 ;
  assign n3834 = n483 & ~n3833 ;
  assign n3835 = ~n1060 & ~n1113 ;
  assign n3836 = n478 & ~n3835 ;
  assign n3865 = ~n3834 & ~n3836 ;
  assign n3837 = ~n960 & ~n1072 ;
  assign n3838 = n423 & ~n3837 ;
  assign n3839 = ~n1059 & ~n1102 ;
  assign n3840 = n443 & ~n3839 ;
  assign n3866 = ~n3838 & ~n3840 ;
  assign n3876 = n3865 & n3866 ;
  assign n3877 = n3875 & n3876 ;
  assign n3857 = ~n1032 & ~n1174 ;
  assign n3858 = n377 & ~n3857 ;
  assign n3859 = ~n1052 & ~n1076 ;
  assign n3860 = n361 & ~n3859 ;
  assign n3871 = ~n3858 & ~n3860 ;
  assign n3861 = ~n1056 & ~n1299 ;
  assign n3862 = n344 & ~n3861 ;
  assign n3863 = ~n982 & ~n1138 ;
  assign n3864 = n408 & ~n3863 ;
  assign n3872 = ~n3862 & ~n3864 ;
  assign n3873 = n3871 & n3872 ;
  assign n3849 = ~n1055 & ~n1195 ;
  assign n3850 = n453 & ~n3849 ;
  assign n3851 = ~n1010 & ~n1024 ;
  assign n3852 = n458 & ~n3851 ;
  assign n3869 = ~n3850 & ~n3852 ;
  assign n3853 = ~n988 & ~n1110 ;
  assign n3854 = n392 & ~n3853 ;
  assign n3855 = ~n1009 & ~n1146 ;
  assign n3856 = n306 & ~n3855 ;
  assign n3870 = ~n3854 & ~n3856 ;
  assign n3874 = n3869 & n3870 ;
  assign n3878 = n3873 & n3874 ;
  assign n3879 = n3877 & n3878 ;
  assign n3880 = \desIn[21]_pad  & n308 ;
  assign n3882 = ~\FP_R_reg[11]/P0001  & n313 ;
  assign n3881 = ~\FP_R_reg[43]/NET0131  & ~n313 ;
  assign n3883 = ~n308 & ~n3881 ;
  assign n3884 = ~n3882 & n3883 ;
  assign n3885 = ~n3880 & ~n3884 ;
  assign n3886 = n3879 & ~n3885 ;
  assign n3887 = ~n3879 & n3885 ;
  assign n3888 = ~n3886 & ~n3887 ;
  assign n3890 = ~n3832 & n3888 ;
  assign n3891 = ~n3889 & n3890 ;
  assign n3892 = ~n3831 & ~n3888 ;
  assign n3893 = n3679 & n3830 ;
  assign n3894 = ~n3730 & ~n3893 ;
  assign n3895 = n3892 & n3894 ;
  assign n3907 = ~n954 & ~n982 ;
  assign n3908 = n488 & ~n3907 ;
  assign n3909 = ~n1010 & ~n1046 ;
  assign n3910 = n344 & ~n3909 ;
  assign n3931 = ~n3908 & ~n3910 ;
  assign n3911 = ~n968 & ~n1006 ;
  assign n3912 = n408 & ~n3911 ;
  assign n3913 = ~n960 & ~n1067 ;
  assign n3914 = n448 & ~n3913 ;
  assign n3932 = ~n3912 & ~n3914 ;
  assign n3939 = n3931 & n3932 ;
  assign n3901 = n453 & ~n3735 ;
  assign n3902 = ~n1009 & ~n1059 ;
  assign n3903 = n463 & ~n3902 ;
  assign n3929 = ~n3901 & ~n3903 ;
  assign n3904 = ~n1002 & ~n1075 ;
  assign n3905 = n443 & ~n3904 ;
  assign n3906 = n483 & ~n3733 ;
  assign n3930 = ~n3905 & ~n3906 ;
  assign n3940 = n3929 & n3930 ;
  assign n3941 = n3939 & n3940 ;
  assign n3922 = ~n988 & ~n1032 ;
  assign n3923 = n438 & ~n3922 ;
  assign n3924 = ~n1055 & ~n1060 ;
  assign n3925 = n361 & ~n3924 ;
  assign n3935 = ~n3923 & ~n3925 ;
  assign n3926 = n377 & ~n3741 ;
  assign n3927 = ~n996 & ~n1056 ;
  assign n3928 = n458 & ~n3927 ;
  assign n3936 = ~n3926 & ~n3928 ;
  assign n3937 = n3935 & n3936 ;
  assign n3915 = ~n940 & ~n1068 ;
  assign n3916 = n392 & ~n3915 ;
  assign n3917 = ~n1052 & ~n1063 ;
  assign n3918 = n478 & ~n3917 ;
  assign n3933 = ~n3916 & ~n3918 ;
  assign n3919 = n306 & ~n3757 ;
  assign n3920 = ~n1005 & ~n1038 ;
  assign n3921 = n423 & ~n3920 ;
  assign n3934 = ~n3919 & ~n3921 ;
  assign n3938 = n3933 & n3934 ;
  assign n3942 = n3937 & n3938 ;
  assign n3943 = n3941 & n3942 ;
  assign n3944 = ~n1228 & n3943 ;
  assign n3945 = n1228 & ~n3943 ;
  assign n3946 = ~n3944 & ~n3945 ;
  assign n3950 = ~n3895 & ~n3946 ;
  assign n3896 = n3679 & ~n3780 ;
  assign n3897 = n3729 & n3830 ;
  assign n3898 = ~n3729 & ~n3830 ;
  assign n3899 = ~n3897 & ~n3898 ;
  assign n3900 = n3896 & ~n3899 ;
  assign n3947 = n3679 & ~n3729 ;
  assign n3948 = n3830 & n3947 ;
  assign n3949 = n3780 & n3948 ;
  assign n3951 = ~n3900 & ~n3949 ;
  assign n3952 = n3950 & n3951 ;
  assign n3953 = ~n3891 & n3952 ;
  assign n3956 = ~n3729 & n3830 ;
  assign n3957 = ~n3780 & n3956 ;
  assign n3958 = n3780 & n3897 ;
  assign n3959 = ~n3957 & ~n3958 ;
  assign n3960 = n3888 & n3959 ;
  assign n3961 = ~n3679 & n3897 ;
  assign n3962 = n3892 & ~n3961 ;
  assign n3963 = ~n3960 & ~n3962 ;
  assign n3964 = ~n3780 & n3888 ;
  assign n3965 = n3729 & ~n3830 ;
  assign n3966 = n3679 & n3965 ;
  assign n3967 = n3964 & n3966 ;
  assign n3954 = ~n3679 & n3780 ;
  assign n3955 = ~n3898 & n3954 ;
  assign n3968 = n3946 & ~n3955 ;
  assign n3969 = ~n3967 & n3968 ;
  assign n3970 = ~n3963 & n3969 ;
  assign n3971 = ~n3953 & ~n3970 ;
  assign n3972 = ~n3888 & n3889 ;
  assign n3973 = n3780 & n3947 ;
  assign n3974 = ~n3830 & n3888 ;
  assign n3975 = n3973 & n3974 ;
  assign n3976 = ~n3972 & ~n3975 ;
  assign n3977 = ~n3971 & n3976 ;
  assign n3978 = ~\desIn[40]_pad  & n308 ;
  assign n3980 = \FP_R_reg[30]/P0001  & ~n313 ;
  assign n3979 = \FP_R_reg[62]/NET0131  & n313 ;
  assign n3981 = ~n308 & ~n3979 ;
  assign n3982 = ~n3980 & n3981 ;
  assign n3983 = ~n3978 & ~n3982 ;
  assign n3984 = n3977 & ~n3983 ;
  assign n3985 = ~n3977 & n3983 ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n4015 = n2589 & n2774 ;
  assign n4016 = ~n2757 & ~n4015 ;
  assign n4017 = ~n2493 & ~n4016 ;
  assign n3993 = n2493 & ~n2589 ;
  assign n4018 = n2646 & n2774 ;
  assign n4019 = ~n2753 & ~n4018 ;
  assign n4020 = n3993 & ~n4019 ;
  assign n4005 = n2753 & n2760 ;
  assign n4021 = ~n2701 & ~n4005 ;
  assign n4022 = ~n4020 & n4021 ;
  assign n4023 = ~n4017 & n4022 ;
  assign n4024 = n2751 & ~n4023 ;
  assign n3989 = n2590 & n2699 ;
  assign n3987 = n2700 & n2753 ;
  assign n3988 = ~n2646 & n2755 ;
  assign n3990 = ~n3987 & ~n3988 ;
  assign n3991 = ~n3989 & n3990 ;
  assign n3992 = ~n2493 & ~n3991 ;
  assign n3998 = n2646 & ~n2758 ;
  assign n3999 = n2760 & n3998 ;
  assign n3994 = ~n2752 & ~n3993 ;
  assign n3995 = n2647 & ~n3994 ;
  assign n3996 = ~n2589 & n2704 ;
  assign n3997 = ~n2699 & n3996 ;
  assign n4000 = ~n3995 & ~n3997 ;
  assign n4001 = ~n3999 & n4000 ;
  assign n4002 = ~n3992 & n4001 ;
  assign n4003 = ~n2751 & ~n4002 ;
  assign n4006 = ~n2705 & ~n4005 ;
  assign n4007 = ~n2543 & n2752 ;
  assign n4008 = n4006 & ~n4007 ;
  assign n4009 = n2493 & ~n4008 ;
  assign n4004 = ~n2493 & n3996 ;
  assign n4012 = n2493 & ~n2768 ;
  assign n4010 = n2543 & n2589 ;
  assign n4011 = ~n2493 & ~n4010 ;
  assign n4013 = n2646 & ~n4011 ;
  assign n4014 = ~n4012 & n4013 ;
  assign n4025 = ~n4004 & ~n4014 ;
  assign n4026 = ~n4009 & n4025 ;
  assign n4027 = ~n4003 & n4026 ;
  assign n4028 = ~n4024 & n4027 ;
  assign n4029 = ~\desIn[42]_pad  & n308 ;
  assign n4031 = \FP_R_reg[22]/P0001  & ~n313 ;
  assign n4030 = \FP_R_reg[54]/NET0131  & n313 ;
  assign n4032 = ~n308 & ~n4030 ;
  assign n4033 = ~n4031 & n4032 ;
  assign n4034 = ~n4029 & ~n4033 ;
  assign n4035 = n4028 & ~n4034 ;
  assign n4036 = ~n4028 & n4034 ;
  assign n4037 = ~n4035 & ~n4036 ;
  assign n4043 = n873 & n907 ;
  assign n4044 = ~n902 & ~n2309 ;
  assign n4045 = ~n4043 & n4044 ;
  assign n4046 = ~n2306 & n4045 ;
  assign n4047 = n816 & ~n4046 ;
  assign n4038 = n759 & n873 ;
  assign n4039 = ~n883 & ~n2312 ;
  assign n4040 = ~n4038 & n4039 ;
  assign n4041 = ~n816 & ~n4040 ;
  assign n4042 = ~n758 & n883 ;
  assign n4048 = ~n2311 & ~n4042 ;
  assign n4049 = ~n4041 & n4048 ;
  assign n4050 = ~n4047 & n4049 ;
  assign n4051 = ~n510 & ~n4050 ;
  assign n4052 = ~n882 & n903 ;
  assign n4053 = ~n889 & ~n2298 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4055 = ~n816 & ~n4054 ;
  assign n4056 = n816 & ~n873 ;
  assign n4057 = ~n904 & ~n2312 ;
  assign n4058 = n4056 & ~n4057 ;
  assign n4059 = ~n882 & ~n913 ;
  assign n4060 = n759 & ~n2308 ;
  assign n4061 = n4059 & n4060 ;
  assign n4062 = n888 & ~n4059 ;
  assign n4063 = ~n4061 & ~n4062 ;
  assign n4064 = ~n4058 & n4063 ;
  assign n4065 = ~n4055 & n4064 ;
  assign n4066 = n510 & ~n4065 ;
  assign n4067 = ~n2297 & ~n2309 ;
  assign n4068 = n873 & ~n4067 ;
  assign n4069 = n816 & ~n4068 ;
  assign n4070 = ~n816 & ~n896 ;
  assign n4071 = ~n2314 & n4070 ;
  assign n4072 = ~n4069 & ~n4071 ;
  assign n4073 = ~n4066 & ~n4072 ;
  assign n4074 = ~n4051 & n4073 ;
  assign n4075 = ~\desIn[44]_pad  & n308 ;
  assign n4077 = \FP_R_reg[14]/P0001  & ~n313 ;
  assign n4076 = \FP_R_reg[46]/NET0131  & n313 ;
  assign n4078 = ~n308 & ~n4076 ;
  assign n4079 = ~n4077 & n4078 ;
  assign n4080 = ~n4075 & ~n4079 ;
  assign n4081 = n4074 & ~n4080 ;
  assign n4082 = ~n4074 & n4080 ;
  assign n4083 = ~n4081 & ~n4082 ;
  assign n4106 = ~n3896 & ~n3899 ;
  assign n4107 = ~n3954 & n4106 ;
  assign n4101 = ~n3896 & ~n3954 ;
  assign n4102 = n3830 & n3888 ;
  assign n4103 = n3899 & ~n4102 ;
  assign n4104 = ~n4101 & n4103 ;
  assign n4093 = ~n3679 & ~n3780 ;
  assign n4105 = n4093 & n4102 ;
  assign n4108 = ~n4104 & ~n4105 ;
  assign n4109 = ~n4107 & n4108 ;
  assign n4110 = ~n3946 & ~n4109 ;
  assign n4084 = n3780 & n3956 ;
  assign n4085 = n3730 & ~n3830 ;
  assign n4086 = ~n4084 & ~n4085 ;
  assign n4087 = ~n3947 & n4086 ;
  assign n4088 = n3946 & ~n4087 ;
  assign n4089 = n3896 & n3897 ;
  assign n4090 = ~n3973 & ~n4089 ;
  assign n4091 = ~n4088 & n4090 ;
  assign n4092 = n3888 & ~n4091 ;
  assign n4094 = n3830 & ~n4093 ;
  assign n4095 = ~n3888 & n3946 ;
  assign n4096 = ~n3730 & n4095 ;
  assign n4097 = ~n3947 & n4096 ;
  assign n4098 = ~n4094 & n4097 ;
  assign n4099 = ~n3679 & n3946 ;
  assign n4100 = n3958 & n4099 ;
  assign n4111 = ~n4098 & ~n4100 ;
  assign n4112 = ~n4092 & n4111 ;
  assign n4113 = ~n4110 & n4112 ;
  assign n4114 = ~\desIn[46]_pad  & n308 ;
  assign n4116 = \FP_R_reg[6]/P0001  & ~n313 ;
  assign n4115 = \FP_R_reg[38]/NET0131  & n313 ;
  assign n4117 = ~n308 & ~n4115 ;
  assign n4118 = ~n4116 & n4117 ;
  assign n4119 = ~n4114 & ~n4118 ;
  assign n4120 = n4113 & ~n4119 ;
  assign n4121 = ~n4113 & n4119 ;
  assign n4122 = ~n4120 & ~n4121 ;
  assign n4123 = ~n2986 & n3036 ;
  assign n4124 = ~n3092 & n3102 ;
  assign n4125 = ~n4123 & ~n4124 ;
  assign n4126 = n2880 & ~n4125 ;
  assign n4130 = n2880 & n3092 ;
  assign n4131 = n3095 & n4130 ;
  assign n4127 = ~n2880 & n3093 ;
  assign n4128 = ~n2932 & ~n2986 ;
  assign n4129 = ~n3092 & n4128 ;
  assign n4134 = ~n4127 & ~n4129 ;
  assign n4135 = ~n4131 & n4134 ;
  assign n4132 = n3038 & n3092 ;
  assign n4133 = ~n2834 & ~n3096 ;
  assign n4136 = ~n4132 & n4133 ;
  assign n4137 = n4135 & n4136 ;
  assign n4138 = ~n4126 & n4137 ;
  assign n4139 = n2880 & ~n3092 ;
  assign n4146 = n3094 & n4139 ;
  assign n4147 = ~n3120 & ~n4146 ;
  assign n4142 = n2986 & n3102 ;
  assign n4143 = n2880 & n3039 ;
  assign n4144 = ~n4142 & ~n4143 ;
  assign n4145 = n3092 & ~n4144 ;
  assign n4140 = n2986 & n3095 ;
  assign n4141 = n4139 & n4140 ;
  assign n4148 = n2834 & ~n4141 ;
  assign n4149 = ~n4145 & n4148 ;
  assign n4150 = n4147 & n4149 ;
  assign n4151 = ~n4138 & ~n4150 ;
  assign n4160 = n3036 & n4129 ;
  assign n4158 = ~n3036 & n3111 ;
  assign n4159 = n3039 & n3109 ;
  assign n4161 = ~n4158 & ~n4159 ;
  assign n4162 = ~n4160 & n4161 ;
  assign n4163 = ~n2880 & ~n4162 ;
  assign n4152 = n3038 & ~n3092 ;
  assign n4153 = n3105 & ~n4123 ;
  assign n4154 = ~n4152 & ~n4153 ;
  assign n4155 = n3101 & ~n4154 ;
  assign n4156 = ~n3036 & n4128 ;
  assign n4157 = n4139 & n4156 ;
  assign n4164 = n2880 & n2932 ;
  assign n4165 = n3118 & n4164 ;
  assign n4166 = ~n4157 & ~n4165 ;
  assign n4167 = ~n4155 & n4166 ;
  assign n4168 = ~n4163 & n4167 ;
  assign n4169 = ~n4151 & n4168 ;
  assign n4170 = ~\desIn[48]_pad  & n308 ;
  assign n4172 = \FP_R_reg[31]/P0001  & ~n313 ;
  assign n4171 = \FP_R_reg[63]/NET0131  & n313 ;
  assign n4173 = ~n308 & ~n4171 ;
  assign n4174 = ~n4172 & n4173 ;
  assign n4175 = ~n4170 & ~n4174 ;
  assign n4176 = n4169 & ~n4175 ;
  assign n4177 = ~n4169 & n4175 ;
  assign n4178 = ~n4176 & ~n4177 ;
  assign n4194 = ~n3096 & ~n4142 ;
  assign n4195 = n3041 & n4194 ;
  assign n4196 = ~n3092 & ~n4195 ;
  assign n4179 = ~n3037 & ~n4140 ;
  assign n4193 = n4130 & ~n4179 ;
  assign n4197 = ~n3117 & ~n4193 ;
  assign n4198 = ~n4196 & n4197 ;
  assign n4199 = ~n2834 & ~n4198 ;
  assign n4180 = ~n2880 & n4179 ;
  assign n4181 = n2880 & ~n4123 ;
  assign n4182 = ~n3110 & n4181 ;
  assign n4183 = ~n4142 & n4182 ;
  assign n4184 = ~n4180 & ~n4183 ;
  assign n4185 = ~n3092 & n3104 ;
  assign n4186 = n2932 & n3112 ;
  assign n4187 = ~n4185 & ~n4186 ;
  assign n4188 = ~n4184 & n4187 ;
  assign n4189 = n2834 & ~n4188 ;
  assign n4190 = ~n2932 & n3116 ;
  assign n4191 = ~n4186 & ~n4190 ;
  assign n4192 = ~n2880 & ~n4191 ;
  assign n4200 = ~n4189 & ~n4192 ;
  assign n4201 = ~n4199 & n4200 ;
  assign n4202 = ~\desIn[4]_pad  & n308 ;
  assign n4204 = \FP_R_reg[9]/P0001  & ~n313 ;
  assign n4203 = \FP_R_reg[41]/NET0131  & n313 ;
  assign n4205 = ~n308 & ~n4203 ;
  assign n4206 = ~n4204 & n4205 ;
  assign n4207 = ~n4202 & ~n4206 ;
  assign n4208 = n4201 & ~n4207 ;
  assign n4209 = ~n4201 & n4207 ;
  assign n4210 = ~n4208 & ~n4209 ;
  assign n4211 = n3039 & ~n3092 ;
  assign n4212 = ~n3093 & ~n4211 ;
  assign n4213 = ~n2880 & ~n4212 ;
  assign n4215 = n2880 & n4142 ;
  assign n4216 = n3095 & n4139 ;
  assign n4214 = n3037 & n3092 ;
  assign n4217 = ~n3116 & ~n4214 ;
  assign n4218 = ~n4216 & n4217 ;
  assign n4219 = ~n4215 & n4218 ;
  assign n4220 = ~n4213 & n4219 ;
  assign n4221 = n2834 & ~n4220 ;
  assign n4222 = n2880 & n4140 ;
  assign n4223 = ~n4157 & ~n4222 ;
  assign n4224 = n4147 & n4223 ;
  assign n4225 = ~n2834 & ~n4224 ;
  assign n4230 = ~n4152 & n4194 ;
  assign n4231 = ~n2834 & ~n2880 ;
  assign n4232 = ~n4230 & n4231 ;
  assign n4229 = n3092 & n4215 ;
  assign n4226 = ~n2880 & n3092 ;
  assign n4227 = ~n3097 & n4226 ;
  assign n4228 = ~n2880 & n4159 ;
  assign n4233 = ~n4165 & ~n4228 ;
  assign n4234 = ~n4227 & n4233 ;
  assign n4235 = ~n4229 & n4234 ;
  assign n4236 = ~n4232 & n4235 ;
  assign n4237 = ~n4225 & n4236 ;
  assign n4238 = ~n4221 & n4237 ;
  assign n4239 = ~\desIn[50]_pad  & n308 ;
  assign n4241 = \FP_R_reg[23]/P0001  & ~n313 ;
  assign n4240 = \FP_R_reg[55]/NET0131  & n313 ;
  assign n4242 = ~n308 & ~n4240 ;
  assign n4243 = ~n4241 & n4242 ;
  assign n4244 = ~n4239 & ~n4243 ;
  assign n4245 = n4238 & ~n4244 ;
  assign n4246 = ~n4238 & n4244 ;
  assign n4247 = ~n4245 & ~n4246 ;
  assign n4249 = ~n3383 & n3555 ;
  assign n4248 = n3429 & n3526 ;
  assign n4250 = ~n3602 & ~n4248 ;
  assign n4251 = ~n4249 & n4250 ;
  assign n4252 = n3331 & ~n4251 ;
  assign n4253 = n3533 & n3541 ;
  assign n4254 = ~n4252 & ~n4253 ;
  assign n4255 = ~n3275 & ~n4254 ;
  assign n4258 = n3565 & n3601 ;
  assign n4256 = n3526 & n3560 ;
  assign n4260 = ~n3528 & ~n4256 ;
  assign n4261 = ~n4258 & n4260 ;
  assign n4257 = n3331 & n3540 ;
  assign n4259 = n3480 & n3554 ;
  assign n4262 = ~n4257 & ~n4259 ;
  assign n4263 = n4261 & n4262 ;
  assign n4264 = n3275 & ~n4263 ;
  assign n4265 = ~n3275 & ~n3429 ;
  assign n4266 = n3526 & n4265 ;
  assign n4268 = ~n3563 & ~n4266 ;
  assign n4269 = n3594 & n4268 ;
  assign n4267 = ~n3383 & n3597 ;
  assign n4270 = ~n4259 & ~n4267 ;
  assign n4271 = n4269 & n4270 ;
  assign n4272 = n3331 & ~n3545 ;
  assign n4273 = ~n3598 & n4272 ;
  assign n4274 = ~n4271 & ~n4273 ;
  assign n4275 = ~n4264 & ~n4274 ;
  assign n4276 = ~n4255 & n4275 ;
  assign n4277 = ~\desIn[52]_pad  & n308 ;
  assign n4279 = \FP_R_reg[15]/P0001  & ~n313 ;
  assign n4278 = \FP_R_reg[47]/NET0131  & n313 ;
  assign n4280 = ~n308 & ~n4278 ;
  assign n4281 = ~n4279 & n4280 ;
  assign n4282 = ~n4277 & ~n4281 ;
  assign n4283 = n4276 & ~n4282 ;
  assign n4284 = ~n4276 & n4282 ;
  assign n4285 = ~n4283 & ~n4284 ;
  assign n4286 = ~\desIn[54]_pad  & n308 ;
  assign n4288 = \FP_R_reg[7]/P0001  & ~n313 ;
  assign n4287 = \FP_R_reg[39]/NET0131  & n313 ;
  assign n4289 = ~n308 & ~n4287 ;
  assign n4290 = ~n4288 & n4289 ;
  assign n4291 = ~n4286 & ~n4290 ;
  assign n4292 = n2753 & n2755 ;
  assign n4295 = ~n2704 & ~n2777 ;
  assign n4296 = ~n2769 & n2777 ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4293 = ~n2493 & n2751 ;
  assign n4294 = n2493 & ~n2751 ;
  assign n4298 = ~n4293 & ~n4294 ;
  assign n4299 = ~n3987 & n4298 ;
  assign n4300 = ~n4297 & n4299 ;
  assign n4303 = n2589 & ~n2778 ;
  assign n4302 = n2543 & ~n2777 ;
  assign n4301 = ~n2646 & n2752 ;
  assign n4304 = n4293 & ~n4301 ;
  assign n4305 = ~n4302 & n4304 ;
  assign n4306 = ~n4303 & n4305 ;
  assign n4307 = ~n4300 & ~n4306 ;
  assign n4308 = ~n4292 & ~n4307 ;
  assign n4309 = ~n2646 & n2700 ;
  assign n4310 = n4294 & ~n4309 ;
  assign n4311 = ~n3997 & n4310 ;
  assign n4312 = ~n4295 & n4311 ;
  assign n4313 = ~n4308 & ~n4312 ;
  assign n4314 = ~n4291 & ~n4313 ;
  assign n4315 = n4291 & n4313 ;
  assign n4316 = ~n4314 & ~n4315 ;
  assign n4323 = n2589 & n2768 ;
  assign n4324 = ~n4018 & ~n4301 ;
  assign n4325 = ~n4323 & n4324 ;
  assign n4326 = n2493 & ~n4325 ;
  assign n4317 = n2699 & n3996 ;
  assign n4318 = n2647 & ~n2777 ;
  assign n4319 = n2543 & n2700 ;
  assign n4320 = ~n4292 & ~n4319 ;
  assign n4321 = ~n4318 & n4320 ;
  assign n4322 = ~n2493 & ~n4321 ;
  assign n4327 = ~n4317 & ~n4322 ;
  assign n4328 = ~n4326 & n4327 ;
  assign n4329 = n2751 & ~n4328 ;
  assign n4330 = n2646 & n2752 ;
  assign n4334 = n2543 & n4330 ;
  assign n4335 = ~n3997 & n4006 ;
  assign n4336 = ~n4334 & n4335 ;
  assign n4331 = ~n2756 & ~n4330 ;
  assign n4332 = n2493 & ~n4331 ;
  assign n4333 = n2776 & ~n4330 ;
  assign n4337 = ~n4332 & ~n4333 ;
  assign n4338 = n4336 & n4337 ;
  assign n4339 = ~n2751 & ~n4338 ;
  assign n4340 = n2493 & n4005 ;
  assign n4341 = ~n2589 & n4018 ;
  assign n4342 = ~n2646 & n4010 ;
  assign n4343 = ~n4341 & ~n4342 ;
  assign n4344 = ~n2493 & ~n4343 ;
  assign n4345 = ~n4340 & ~n4344 ;
  assign n4346 = ~n4339 & n4345 ;
  assign n4347 = ~n4329 & n4346 ;
  assign n4348 = ~\desIn[56]_pad  & n308 ;
  assign n4350 = \FP_R_reg[32]/P0001  & ~n313 ;
  assign n4349 = \FP_R_reg[64]/NET0131  & n313 ;
  assign n4351 = ~n308 & ~n4349 ;
  assign n4352 = ~n4350 & n4351 ;
  assign n4353 = ~n4348 & ~n4352 ;
  assign n4354 = n4347 & ~n4353 ;
  assign n4355 = ~n4347 & n4353 ;
  assign n4356 = ~n4354 & ~n4355 ;
  assign n4357 = ~n3679 & n3898 ;
  assign n4358 = ~n3948 & ~n4357 ;
  assign n4366 = ~n3780 & n3897 ;
  assign n4367 = n4358 & ~n4366 ;
  assign n4368 = ~n3946 & ~n4367 ;
  assign n4369 = n3679 & n3831 ;
  assign n4370 = ~n3780 & n3965 ;
  assign n4371 = ~n3958 & ~n4370 ;
  assign n4372 = n3946 & ~n4371 ;
  assign n4373 = ~n4369 & ~n4372 ;
  assign n4374 = ~n4368 & n4373 ;
  assign n4375 = ~n3888 & ~n4374 ;
  assign n4359 = n3730 & n4102 ;
  assign n4360 = ~n3966 & ~n4359 ;
  assign n4361 = n4358 & n4360 ;
  assign n4362 = ~n3780 & ~n4361 ;
  assign n4363 = ~n3679 & n4084 ;
  assign n4364 = ~n4362 & ~n4363 ;
  assign n4365 = n3946 & ~n4364 ;
  assign n4376 = n3679 & ~n3898 ;
  assign n4377 = n3888 & ~n3897 ;
  assign n4378 = ~n4357 & n4377 ;
  assign n4379 = ~n4376 & n4378 ;
  assign n4380 = ~n4089 & ~n4379 ;
  assign n4381 = ~n3946 & ~n4380 ;
  assign n4382 = n3729 & n3893 ;
  assign n4383 = ~n4085 & ~n4382 ;
  assign n4384 = n3780 & n3888 ;
  assign n4385 = ~n4383 & n4384 ;
  assign n4386 = ~n4381 & ~n4385 ;
  assign n4387 = ~n4365 & n4386 ;
  assign n4388 = ~n4375 & n4387 ;
  assign n4389 = ~\desIn[60]_pad  & n308 ;
  assign n4391 = \FP_R_reg[16]/P0001  & ~n313 ;
  assign n4390 = \FP_R_reg[48]/NET0131  & n313 ;
  assign n4392 = ~n308 & ~n4390 ;
  assign n4393 = ~n4391 & n4392 ;
  assign n4394 = ~n4389 & ~n4393 ;
  assign n4395 = n4388 & ~n4394 ;
  assign n4396 = ~n4388 & n4394 ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4414 = n1449 & ~n1468 ;
  assign n4415 = ~n2403 & n4414 ;
  assign n4417 = n1393 & n2411 ;
  assign n4416 = n1346 & n1485 ;
  assign n4418 = ~n1449 & ~n4416 ;
  assign n4419 = ~n4417 & n4418 ;
  assign n4420 = ~n4415 & ~n4419 ;
  assign n4421 = n1287 & n4416 ;
  assign n4422 = n2408 & ~n4421 ;
  assign n4423 = ~n4420 & n4422 ;
  assign n4424 = ~n1096 & ~n4423 ;
  assign n4408 = ~n1346 & ~n1459 ;
  assign n4407 = ~n1449 & ~n1485 ;
  assign n4409 = n1287 & n4407 ;
  assign n4410 = ~n4408 & n4409 ;
  assign n4400 = n1287 & n2391 ;
  assign n4406 = ~n1231 & n1455 ;
  assign n4411 = ~n4400 & ~n4406 ;
  assign n4412 = ~n4410 & n4411 ;
  assign n4413 = n1096 & ~n4412 ;
  assign n4398 = ~n1467 & n1480 ;
  assign n4399 = n1449 & ~n4398 ;
  assign n4402 = n1346 & n2411 ;
  assign n4403 = ~n2390 & ~n4402 ;
  assign n4404 = n1096 & n1449 ;
  assign n4405 = ~n4403 & n4404 ;
  assign n4401 = ~n1449 & n4400 ;
  assign n4425 = ~n2410 & ~n4401 ;
  assign n4426 = ~n4405 & n4425 ;
  assign n4427 = ~n4399 & n4426 ;
  assign n4428 = ~n4413 & n4427 ;
  assign n4429 = ~n4424 & n4428 ;
  assign n4430 = ~\desIn[6]_pad  & n308 ;
  assign n4432 = \FP_R_reg[1]/P0001  & ~n313 ;
  assign n4431 = \FP_R_reg[33]/NET0131  & n313 ;
  assign n4433 = ~n308 & ~n4431 ;
  assign n4434 = ~n4432 & n4433 ;
  assign n4435 = ~n4430 & ~n4434 ;
  assign n4436 = n4429 & ~n4435 ;
  assign n4437 = ~n4429 & n4435 ;
  assign n4438 = ~n4436 & ~n4437 ;
  assign n4439 = ~\desIn[8]_pad  & n308 ;
  assign n4441 = \FP_R_reg[26]/P0001  & ~n313 ;
  assign n4440 = \FP_R_reg[58]/NET0131  & n313 ;
  assign n4442 = ~n308 & ~n4440 ;
  assign n4443 = ~n4441 & n4442 ;
  assign n4444 = ~n4439 & ~n4443 ;
  assign n4446 = n1459 & n1489 ;
  assign n4447 = ~n1477 & ~n4446 ;
  assign n4448 = ~n1449 & ~n4447 ;
  assign n4451 = ~n1347 & ~n2394 ;
  assign n4452 = n1462 & ~n4451 ;
  assign n4449 = ~n1346 & n1459 ;
  assign n4450 = ~n1463 & n4449 ;
  assign n4453 = ~n4400 & ~n4450 ;
  assign n4454 = ~n4452 & n4453 ;
  assign n4455 = ~n4448 & n4454 ;
  assign n4456 = n1096 & ~n4455 ;
  assign n4457 = n1484 & n4408 ;
  assign n4458 = ~n1486 & ~n2407 ;
  assign n4459 = ~n4402 & n4458 ;
  assign n4460 = ~n4457 & n4459 ;
  assign n4461 = ~n1096 & ~n4460 ;
  assign n4462 = ~n1456 & ~n4406 ;
  assign n4463 = ~n1096 & ~n1449 ;
  assign n4464 = ~n4462 & n4463 ;
  assign n4445 = n1347 & n1460 ;
  assign n4467 = ~n1491 & ~n4445 ;
  assign n4465 = n1463 & n4416 ;
  assign n4466 = n1492 & n4407 ;
  assign n4468 = ~n4465 & ~n4466 ;
  assign n4469 = n4467 & n4468 ;
  assign n4470 = ~n4464 & n4469 ;
  assign n4471 = ~n4461 & n4470 ;
  assign n4472 = ~n4456 & n4471 ;
  assign n4473 = ~n4444 & n4472 ;
  assign n4474 = n4444 & ~n4472 ;
  assign n4475 = ~n4473 & ~n4474 ;
  assign n4476 = ~n1682 & n2341 ;
  assign n4477 = ~n2358 & ~n4476 ;
  assign n4479 = ~n1853 & ~n2337 ;
  assign n4478 = n1865 & n1877 ;
  assign n4480 = ~n2349 & ~n4478 ;
  assign n4481 = n4479 & n4480 ;
  assign n4482 = n4477 & n4481 ;
  assign n4483 = ~n1739 & n1855 ;
  assign n4484 = n1853 & ~n4483 ;
  assign n4485 = ~n2356 & n4484 ;
  assign n4486 = ~n4482 & ~n4485 ;
  assign n4488 = ~n1874 & ~n2347 ;
  assign n4489 = n1796 & ~n4488 ;
  assign n4487 = n1739 & n2348 ;
  assign n4490 = n1570 & ~n4487 ;
  assign n4491 = ~n4489 & n4490 ;
  assign n4492 = ~n4486 & n4491 ;
  assign n4494 = ~n2343 & n2355 ;
  assign n4495 = ~n1853 & ~n4494 ;
  assign n4497 = n1626 & n1796 ;
  assign n4496 = n1738 & n1865 ;
  assign n4498 = n1853 & ~n4496 ;
  assign n4499 = ~n4497 & n4498 ;
  assign n4500 = ~n4495 & ~n4499 ;
  assign n4493 = ~n1626 & n2337 ;
  assign n4501 = ~n1570 & n1868 ;
  assign n4502 = ~n4493 & n4501 ;
  assign n4503 = n4477 & n4502 ;
  assign n4504 = ~n4500 & n4503 ;
  assign n4505 = ~n4492 & ~n4504 ;
  assign n4506 = ~\desIn[36]_pad  & n308 ;
  assign n4508 = \FP_R_reg[13]/P0001  & ~n313 ;
  assign n4507 = \FP_R_reg[45]/NET0131  & n313 ;
  assign n4509 = ~n308 & ~n4507 ;
  assign n4510 = ~n4508 & n4509 ;
  assign n4511 = ~n4506 & ~n4510 ;
  assign n4512 = ~n4505 & ~n4511 ;
  assign n4513 = n4505 & n4511 ;
  assign n4514 = ~n4512 & ~n4513 ;
  assign n4529 = ~n1798 & n1853 ;
  assign n4527 = ~n1878 & ~n2341 ;
  assign n4528 = ~n1853 & ~n4527 ;
  assign n4530 = ~n1886 & ~n4528 ;
  assign n4531 = ~n4529 & n4530 ;
  assign n4532 = ~n1570 & ~n4531 ;
  assign n4516 = n1853 & n1880 ;
  assign n4518 = ~n1861 & ~n2358 ;
  assign n4515 = n1863 & n2345 ;
  assign n4517 = ~n1860 & n1865 ;
  assign n4519 = ~n4515 & ~n4517 ;
  assign n4520 = n4518 & n4519 ;
  assign n4521 = ~n4516 & n4520 ;
  assign n4522 = n1570 & ~n4521 ;
  assign n4523 = n1626 & n1860 ;
  assign n4524 = ~n4493 & ~n4523 ;
  assign n4525 = n1853 & ~n4524 ;
  assign n4526 = n1879 & n2345 ;
  assign n4533 = ~n4525 & ~n4526 ;
  assign n4534 = ~n4522 & n4533 ;
  assign n4535 = ~n4532 & n4534 ;
  assign n4536 = ~\desIn[10]_pad  & n308 ;
  assign n4538 = \FP_R_reg[18]/P0001  & ~n313 ;
  assign n4537 = \FP_R_reg[50]/NET0131  & n313 ;
  assign n4539 = ~n308 & ~n4537 ;
  assign n4540 = ~n4538 & n4539 ;
  assign n4541 = ~n4536 & ~n4540 ;
  assign n4542 = n4535 & ~n4541 ;
  assign n4543 = ~n4535 & n4541 ;
  assign n4544 = ~n4542 & ~n4543 ;
  assign n4559 = ~n2070 & n3167 ;
  assign n4560 = ~n2261 & ~n4559 ;
  assign n4561 = n1968 & ~n4560 ;
  assign n4566 = n3206 & ~n4561 ;
  assign n4562 = ~n2255 & ~n2258 ;
  assign n4563 = ~n2181 & ~n4562 ;
  assign n4564 = ~n2257 & ~n3159 ;
  assign n4565 = n2181 & ~n4564 ;
  assign n4567 = ~n4563 & ~n4565 ;
  assign n4568 = n4566 & n4567 ;
  assign n4569 = ~n2244 & ~n4568 ;
  assign n4545 = ~n2020 & ~n2189 ;
  assign n4546 = ~n2274 & n4545 ;
  assign n4547 = ~n2181 & ~n2255 ;
  assign n4548 = ~n3148 & n4547 ;
  assign n4549 = ~n4546 & n4548 ;
  assign n4550 = ~n2255 & ~n3147 ;
  assign n4551 = ~n3172 & n4550 ;
  assign n4552 = n2181 & ~n4551 ;
  assign n4553 = ~n4549 & ~n4552 ;
  assign n4554 = n2244 & ~n4553 ;
  assign n4557 = ~n3148 & ~n3158 ;
  assign n4558 = n2181 & ~n4557 ;
  assign n4555 = ~n2190 & ~n2272 ;
  assign n4556 = n2270 & ~n4555 ;
  assign n4570 = ~n2269 & ~n4556 ;
  assign n4571 = ~n4558 & n4570 ;
  assign n4572 = ~n4554 & n4571 ;
  assign n4573 = ~n4569 & n4572 ;
  assign n4574 = ~\desIn[20]_pad  & n308 ;
  assign n4576 = \FP_R_reg[11]/P0001  & ~n313 ;
  assign n4575 = \FP_R_reg[43]/NET0131  & n313 ;
  assign n4577 = ~n308 & ~n4575 ;
  assign n4578 = ~n4576 & n4577 ;
  assign n4579 = ~n4574 & ~n4578 ;
  assign n4580 = n4573 & ~n4579 ;
  assign n4581 = ~n4573 & n4579 ;
  assign n4582 = ~n4580 & ~n4581 ;
  assign n4586 = ~n3542 & ~n3574 ;
  assign n4587 = ~n3597 & n4586 ;
  assign n4588 = ~n3331 & ~n4587 ;
  assign n4583 = ~n3526 & n4249 ;
  assign n4584 = ~n3576 & ~n4583 ;
  assign n4585 = n3331 & ~n4584 ;
  assign n4589 = ~n3534 & ~n3558 ;
  assign n4590 = ~n3598 & n4589 ;
  assign n4591 = ~n4585 & n4590 ;
  assign n4592 = ~n4588 & n4591 ;
  assign n4593 = n3275 & ~n4592 ;
  assign n4595 = n3331 & ~n3554 ;
  assign n4594 = ~n3480 & ~n3560 ;
  assign n4596 = ~n4249 & ~n4594 ;
  assign n4597 = n4595 & n4596 ;
  assign n4598 = n3527 & n3565 ;
  assign n4599 = ~n3557 & ~n3607 ;
  assign n4600 = ~n4598 & n4599 ;
  assign n4601 = ~n4597 & n4600 ;
  assign n4602 = ~n3275 & ~n4601 ;
  assign n4605 = ~n3331 & n3606 ;
  assign n4603 = n3331 & n3480 ;
  assign n4604 = n3430 & n4603 ;
  assign n4606 = ~n3621 & ~n4604 ;
  assign n4607 = ~n4605 & n4606 ;
  assign n4608 = ~n4602 & n4607 ;
  assign n4609 = ~n4593 & n4608 ;
  assign n4610 = ~\desIn[16]_pad  & n308 ;
  assign n4612 = \FP_R_reg[27]/P0001  & ~n313 ;
  assign n4611 = \FP_R_reg[59]/NET0131  & n313 ;
  assign n4613 = ~n308 & ~n4611 ;
  assign n4614 = ~n4612 & n4613 ;
  assign n4615 = ~n4610 & ~n4614 ;
  assign n4616 = n4609 & ~n4615 ;
  assign n4617 = ~n4609 & n4615 ;
  assign n4618 = ~n4616 & ~n4617 ;
  assign n4632 = ~n884 & ~n2313 ;
  assign n4633 = ~n816 & ~n4632 ;
  assign n4634 = n685 & n4056 ;
  assign n4635 = ~n4068 & ~n4634 ;
  assign n4636 = ~n4633 & n4635 ;
  assign n4637 = n510 & ~n4636 ;
  assign n4622 = n760 & ~n816 ;
  assign n4623 = ~n883 & ~n4622 ;
  assign n4624 = n897 & n4623 ;
  assign n4619 = n903 & ~n913 ;
  assign n4620 = ~n884 & ~n4619 ;
  assign n4621 = n816 & ~n4620 ;
  assign n4625 = ~n2307 & ~n4621 ;
  assign n4626 = n4624 & n4625 ;
  assign n4627 = ~n510 & ~n4626 ;
  assign n4629 = n758 & n883 ;
  assign n4630 = ~n4043 & ~n4629 ;
  assign n4631 = ~n816 & ~n4630 ;
  assign n4628 = n816 & n2296 ;
  assign n4638 = ~n2310 & ~n4628 ;
  assign n4639 = ~n4631 & n4638 ;
  assign n4640 = ~n4627 & n4639 ;
  assign n4641 = ~n4637 & n4640 ;
  assign n4642 = ~\desIn[62]_pad  & n308 ;
  assign n4644 = \FP_R_reg[8]/P0001  & ~n313 ;
  assign n4643 = \FP_R_reg[40]/NET0131  & n313 ;
  assign n4645 = ~n308 & ~n4643 ;
  assign n4646 = ~n4644 & n4645 ;
  assign n4647 = ~n4642 & ~n4646 ;
  assign n4648 = n4641 & ~n4647 ;
  assign n4649 = ~n4641 & n4647 ;
  assign n4650 = ~n4648 & ~n4649 ;
  assign n4662 = ~n3961 & ~n4369 ;
  assign n4663 = n3959 & n4662 ;
  assign n4664 = n3888 & ~n4663 ;
  assign n4665 = n3729 & n4369 ;
  assign n4666 = ~n4664 & ~n4665 ;
  assign n4667 = ~n3946 & ~n4666 ;
  assign n4651 = ~n3888 & n4106 ;
  assign n4656 = n3679 & ~n3956 ;
  assign n4657 = n3964 & n4656 ;
  assign n4658 = ~n4651 & ~n4657 ;
  assign n4652 = ~n3679 & n3831 ;
  assign n4653 = ~n4084 & ~n4652 ;
  assign n4654 = n3888 & ~n4653 ;
  assign n4655 = n3896 & n4103 ;
  assign n4659 = ~n4654 & ~n4655 ;
  assign n4660 = n4658 & n4659 ;
  assign n4661 = n3946 & ~n4660 ;
  assign n4671 = ~n3900 & n4086 ;
  assign n4672 = ~n3888 & ~n3946 ;
  assign n4673 = ~n4671 & n4672 ;
  assign n4669 = n3780 & ~n3888 ;
  assign n4670 = n4357 & n4669 ;
  assign n4668 = ~n3729 & n4105 ;
  assign n4674 = ~n3967 & ~n4668 ;
  assign n4675 = ~n4670 & n4674 ;
  assign n4676 = ~n4673 & n4675 ;
  assign n4677 = ~n4661 & n4676 ;
  assign n4678 = ~n4667 & n4677 ;
  assign n4679 = ~\desIn[58]_pad  & n308 ;
  assign n4681 = \FP_R_reg[24]/P0001  & ~n313 ;
  assign n4680 = \FP_R_reg[56]/NET0131  & n313 ;
  assign n4682 = ~n308 & ~n4680 ;
  assign n4683 = ~n4681 & n4682 ;
  assign n4684 = ~n4679 & ~n4683 ;
  assign n4685 = n4678 & ~n4684 ;
  assign n4686 = ~n4678 & n4684 ;
  assign n4687 = ~n4685 & ~n4686 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \desOut[0]_pad  = n934 ;
  assign \desOut[11]_pad  = ~n870 ;
  assign \desOut[12]_pad  = n1512 ;
  assign \desOut[13]_pad  = ~n1518 ;
  assign \desOut[14]_pad  = n1910 ;
  assign \desOut[15]_pad  = ~n1918 ;
  assign \desOut[18]_pad  = n2287 ;
  assign \desOut[1]_pad  = ~n2123 ;
  assign \desOut[22]_pad  = n2330 ;
  assign \desOut[23]_pad  = ~n2336 ;
  assign \desOut[24]_pad  = n2383 ;
  assign \desOut[25]_pad  = ~n2389 ;
  assign \desOut[26]_pad  = n2431 ;
  assign \desOut[28]_pad  = ~n2788 ;
  assign \desOut[2]_pad  = n3141 ;
  assign \desOut[30]_pad  = n3188 ;
  assign \desOut[32]_pad  = ~n3225 ;
  assign \desOut[34]_pad  = n3589 ;
  assign \desOut[35]_pad  = ~n755 ;
  assign \desOut[37]_pad  = ~n1284 ;
  assign \desOut[38]_pad  = ~n3633 ;
  assign \desOut[39]_pad  = ~n1632 ;
  assign \desOut[3]_pad  = ~n626 ;
  assign \desOut[40]_pad  = ~n3986 ;
  assign \desOut[42]_pad  = n4037 ;
  assign \desOut[44]_pad  = n4083 ;
  assign \desOut[45]_pad  = ~n1343 ;
  assign \desOut[46]_pad  = n4122 ;
  assign \desOut[48]_pad  = n4178 ;
  assign \desOut[4]_pad  = n4210 ;
  assign \desOut[50]_pad  = ~n4247 ;
  assign \desOut[52]_pad  = n4285 ;
  assign \desOut[54]_pad  = n4316 ;
  assign \desOut[56]_pad  = n4356 ;
  assign \desOut[57]_pad  = ~n2929 ;
  assign \desOut[59]_pad  = ~n2198 ;
  assign \desOut[5]_pad  = ~n1688 ;
  assign \desOut[60]_pad  = n4397 ;
  assign \desOut[61]_pad  = ~n682 ;
  assign \desOut[63]_pad  = ~n1524 ;
  assign \desOut[6]_pad  = n4438 ;
  assign \desOut[8]_pad  = n4475 ;
  assign \desOut[9]_pad  = ~n2643 ;
  assign \g13525_dup/_0_  = ~n4514 ;
  assign \g13583_dup/_0_  = n4544 ;
  assign \g17813/_3_  = ~n1745 ;
  assign \g17816/_3_  = ~n3380 ;
  assign \g17819/_3_  = ~n1446 ;
  assign \g17822/_3_  = ~n2135 ;
  assign \g17836/_3_  = ~n2490 ;
  assign \g17871/_3_  = ~n1576 ;
  assign \g17878/_1_  = ~n318 ;
  assign \g17881/_3_  = ~n3885 ;
  assign \g17966/_2_  = ~n3328 ;
  assign \g17969/_3_  = ~n2017 ;
  assign \g17996/_2_  = ~n1228 ;
  assign \g19574_dup/_3_  = ~n4582 ;
  assign \g19619_dup/_3_  = n4618 ;
  assign \g19756_dup/_3_  = n4650 ;
  assign \g20263/_3_  = ~n2696 ;
  assign \g20541/_2_  = ~n2983 ;
  assign \g20691/_1_  = n813 ;
  assign \g20740_dup/_3_  = n4687 ;
  assign \g67/_2_  = ~n1850 ;
endmodule
