module top( a_pad , b_pad , c_pad , d_pad , e_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , \a0_pad  , \b0_pad  , \c0_pad  , \d0_pad  , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  output \a0_pad  ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \d0_pad  ;
  output r_pad ;
  output s_pad ;
  output t_pad ;
  output u_pad ;
  output v_pad ;
  output w_pad ;
  output x_pad ;
  output y_pad ;
  output z_pad ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n17 = a_pad & ~l_pad ;
  assign n18 = m_pad & n_pad ;
  assign n19 = ~m_pad & ~n_pad ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = n17 & ~n20 ;
  assign n22 = c_pad & d_pad ;
  assign n23 = e_pad & n22 ;
  assign n24 = k_pad & n_pad ;
  assign n25 = ~n23 & n24 ;
  assign n26 = m_pad & n17 ;
  assign n27 = n25 & n26 ;
  assign n28 = b_pad & ~n24 ;
  assign n29 = b_pad & e_pad ;
  assign n30 = n22 & n29 ;
  assign n31 = ~n28 & ~n30 ;
  assign n32 = ~b_pad & n_pad ;
  assign n33 = n26 & ~n32 ;
  assign n34 = n31 & n33 ;
  assign n35 = ~k_pad & n17 ;
  assign n36 = n18 & n35 ;
  assign n37 = ~b_pad & ~m_pad ;
  assign n38 = ~n_pad & n37 ;
  assign n39 = ~m_pad & n_pad ;
  assign n40 = m_pad & n24 ;
  assign n41 = g_pad & h_pad ;
  assign n42 = i_pad & j_pad ;
  assign n43 = n41 & n42 ;
  assign n44 = n40 & n43 ;
  assign n45 = n40 & ~n43 ;
  assign n46 = n23 & ~n39 ;
  assign n47 = b_pad & k_pad ;
  assign n48 = ~n46 & n47 ;
  assign n49 = n23 & n24 ;
  assign n50 = n26 & ~n49 ;
  assign \a0_pad  = n21 ;
  assign \b0_pad  = n27 ;
  assign \c0_pad  = n34 ;
  assign \d0_pad  = n36 ;
  assign r_pad = ~n38 ;
  assign s_pad = ~n39 ;
  assign t_pad = ~n44 ;
  assign u_pad = ~n45 ;
  assign v_pad = ~p_pad ;
  assign w_pad = ~o_pad ;
  assign x_pad = n48 ;
  assign y_pad = ~q_pad ;
  assign z_pad = ~n50 ;
endmodule
