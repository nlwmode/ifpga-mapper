module top( \inA0_pad  , \inA10_pad  , \inA11_pad  , \inA12_pad  , \inA13_pad  , \inA14_pad  , \inA15_pad  , \inA1_pad  , \inA2_pad  , \inA3_pad  , \inA4_pad  , \inA5_pad  , \inA6_pad  , \inA7_pad  , \inA8_pad  , \inA9_pad  , \inB0_pad  , \inB10_pad  , \inB11_pad  , \inB12_pad  , \inB13_pad  , \inB14_pad  , \inB15_pad  , \inB1_pad  , \inB2_pad  , \inB3_pad  , \inB4_pad  , \inB5_pad  , \inB6_pad  , \inB7_pad  , \inB8_pad  , \inB9_pad  , \inC0_pad  , \inC10_pad  , \inC11_pad  , \inC12_pad  , \inC13_pad  , \inC14_pad  , \inC15_pad  , \inC1_pad  , \inC2_pad  , \inC3_pad  , \inC4_pad  , \inC5_pad  , \inC6_pad  , \inC7_pad  , \inC8_pad  , \inC9_pad  , \inD0_pad  , \inD10_pad  , \inD11_pad  , \inD12_pad  , \inD13_pad  , \inD14_pad  , \inD15_pad  , \inD1_pad  , \inD2_pad  , \inD3_pad  , \inD4_pad  , \inD5_pad  , \inD6_pad  , \inD7_pad  , \inD8_pad  , \inD9_pad  , \musel1_pad  , \musel2_pad  , \musel3_pad  , \musel4_pad  , \opsel0_pad  , \opsel1_pad  , \opsel2_pad  , \opsel3_pad  , \sh0_pad  , \sh1_pad  , \sh2_pad  , \O0_pad  , \O10_pad  , \O11_pad  , \O12_pad  , \O13_pad  , \O14_pad  , \O15_pad  , \O1_pad  , \O2_pad  , \O3_pad  , \O4_pad  , \O5_pad  , \O6_pad  , \O7_pad  , \O8_pad  , \O9_pad  );
  input \inA0_pad  ;
  input \inA10_pad  ;
  input \inA11_pad  ;
  input \inA12_pad  ;
  input \inA13_pad  ;
  input \inA14_pad  ;
  input \inA15_pad  ;
  input \inA1_pad  ;
  input \inA2_pad  ;
  input \inA3_pad  ;
  input \inA4_pad  ;
  input \inA5_pad  ;
  input \inA6_pad  ;
  input \inA7_pad  ;
  input \inA8_pad  ;
  input \inA9_pad  ;
  input \inB0_pad  ;
  input \inB10_pad  ;
  input \inB11_pad  ;
  input \inB12_pad  ;
  input \inB13_pad  ;
  input \inB14_pad  ;
  input \inB15_pad  ;
  input \inB1_pad  ;
  input \inB2_pad  ;
  input \inB3_pad  ;
  input \inB4_pad  ;
  input \inB5_pad  ;
  input \inB6_pad  ;
  input \inB7_pad  ;
  input \inB8_pad  ;
  input \inB9_pad  ;
  input \inC0_pad  ;
  input \inC10_pad  ;
  input \inC11_pad  ;
  input \inC12_pad  ;
  input \inC13_pad  ;
  input \inC14_pad  ;
  input \inC15_pad  ;
  input \inC1_pad  ;
  input \inC2_pad  ;
  input \inC3_pad  ;
  input \inC4_pad  ;
  input \inC5_pad  ;
  input \inC6_pad  ;
  input \inC7_pad  ;
  input \inC8_pad  ;
  input \inC9_pad  ;
  input \inD0_pad  ;
  input \inD10_pad  ;
  input \inD11_pad  ;
  input \inD12_pad  ;
  input \inD13_pad  ;
  input \inD14_pad  ;
  input \inD15_pad  ;
  input \inD1_pad  ;
  input \inD2_pad  ;
  input \inD3_pad  ;
  input \inD4_pad  ;
  input \inD5_pad  ;
  input \inD6_pad  ;
  input \inD7_pad  ;
  input \inD8_pad  ;
  input \inD9_pad  ;
  input \musel1_pad  ;
  input \musel2_pad  ;
  input \musel3_pad  ;
  input \musel4_pad  ;
  input \opsel0_pad  ;
  input \opsel1_pad  ;
  input \opsel2_pad  ;
  input \opsel3_pad  ;
  input \sh0_pad  ;
  input \sh1_pad  ;
  input \sh2_pad  ;
  output \O0_pad  ;
  output \O10_pad  ;
  output \O11_pad  ;
  output \O12_pad  ;
  output \O13_pad  ;
  output \O14_pad  ;
  output \O15_pad  ;
  output \O1_pad  ;
  output \O2_pad  ;
  output \O3_pad  ;
  output \O4_pad  ;
  output \O5_pad  ;
  output \O6_pad  ;
  output \O7_pad  ;
  output \O8_pad  ;
  output \O9_pad  ;
  wire n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 ;
  assign n76 = ~\opsel2_pad  & \opsel3_pad  ;
  assign n77 = ~\musel3_pad  & \musel4_pad  ;
  assign n78 = ~\musel1_pad  & ~\musel2_pad  ;
  assign n79 = n77 & n78 ;
  assign n80 = \inD3_pad  & n79 ;
  assign n81 = \musel3_pad  & ~\musel4_pad  ;
  assign n82 = \musel1_pad  & \musel2_pad  ;
  assign n83 = ~n78 & ~n82 ;
  assign n84 = \inB3_pad  & n83 ;
  assign n85 = \inD3_pad  & n82 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = n81 & ~n86 ;
  assign n88 = ~n80 & ~n87 ;
  assign n89 = ~\sh2_pad  & ~n88 ;
  assign n90 = \inD0_pad  & n79 ;
  assign n91 = \inB0_pad  & n83 ;
  assign n92 = \inD0_pad  & n82 ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = n81 & ~n93 ;
  assign n95 = ~n90 & ~n94 ;
  assign n96 = \sh2_pad  & ~n95 ;
  assign n97 = ~n89 & ~n96 ;
  assign n98 = \sh1_pad  & ~n97 ;
  assign n99 = \inD5_pad  & n79 ;
  assign n100 = \inB5_pad  & n83 ;
  assign n101 = \inD5_pad  & n82 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = n81 & ~n102 ;
  assign n104 = ~n99 & ~n103 ;
  assign n105 = \sh2_pad  & ~n104 ;
  assign n106 = \inD1_pad  & n79 ;
  assign n107 = \inB1_pad  & n83 ;
  assign n108 = \inD1_pad  & n82 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = n81 & ~n109 ;
  assign n111 = ~n106 & ~n110 ;
  assign n112 = ~\sh2_pad  & ~n111 ;
  assign n113 = ~n105 & ~n112 ;
  assign n114 = ~\sh1_pad  & ~n113 ;
  assign n115 = ~n98 & ~n114 ;
  assign n116 = \sh0_pad  & ~n115 ;
  assign n134 = \inD4_pad  & n79 ;
  assign n135 = \inB4_pad  & n83 ;
  assign n136 = \inD4_pad  & n82 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = n81 & ~n137 ;
  assign n139 = ~n134 & ~n138 ;
  assign n140 = \sh2_pad  & ~n139 ;
  assign n133 = ~\sh2_pad  & ~n95 ;
  assign n141 = ~\sh1_pad  & ~n133 ;
  assign n142 = ~n140 & n141 ;
  assign n124 = \inD2_pad  & n79 ;
  assign n125 = \inB2_pad  & n83 ;
  assign n126 = \inD2_pad  & n82 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = n81 & ~n127 ;
  assign n129 = ~n124 & ~n128 ;
  assign n130 = ~\sh2_pad  & ~n129 ;
  assign n117 = \inD8_pad  & n79 ;
  assign n118 = \inB8_pad  & n83 ;
  assign n119 = \inD8_pad  & n82 ;
  assign n120 = ~n118 & ~n119 ;
  assign n121 = n81 & ~n120 ;
  assign n122 = ~n117 & ~n121 ;
  assign n123 = \sh2_pad  & ~n122 ;
  assign n131 = \sh1_pad  & ~n123 ;
  assign n132 = ~n130 & n131 ;
  assign n143 = ~\sh0_pad  & ~n132 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = ~n116 & ~n144 ;
  assign n146 = ~\opsel0_pad  & ~\opsel1_pad  ;
  assign n147 = ~n145 & n146 ;
  assign n148 = \opsel0_pad  & \opsel1_pad  ;
  assign n149 = ~n146 & ~n148 ;
  assign n150 = ~\musel2_pad  & \musel3_pad  ;
  assign n151 = \inD0_pad  & n150 ;
  assign n152 = \musel2_pad  & ~\musel3_pad  ;
  assign n153 = \inB0_pad  & n152 ;
  assign n154 = ~n151 & ~n153 ;
  assign n155 = ~\musel1_pad  & ~n154 ;
  assign n156 = \musel1_pad  & ~\musel3_pad  ;
  assign n157 = \inA0_pad  & ~\musel2_pad  ;
  assign n158 = \inC0_pad  & \musel2_pad  ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = n156 & ~n159 ;
  assign n161 = ~n155 & ~n160 ;
  assign n162 = ~\musel4_pad  & ~n161 ;
  assign n163 = \inC0_pad  & n79 ;
  assign n164 = \inA0_pad  & n83 ;
  assign n165 = \musel1_pad  & n158 ;
  assign n166 = ~n164 & ~n165 ;
  assign n167 = n81 & ~n166 ;
  assign n168 = ~n163 & ~n167 ;
  assign n169 = ~n162 & ~n168 ;
  assign n170 = n162 & n168 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = n149 & ~n171 ;
  assign n173 = ~n147 & ~n172 ;
  assign n174 = n76 & ~n173 ;
  assign n175 = \opsel2_pad  & ~n146 ;
  assign n181 = n145 & n175 ;
  assign n176 = \inC0_pad  & ~\musel1_pad  ;
  assign n177 = ~n157 & ~n176 ;
  assign n178 = n77 & ~n78 ;
  assign n179 = ~n177 & n178 ;
  assign n180 = ~n175 & ~n179 ;
  assign n182 = ~\opsel2_pad  & n146 ;
  assign n183 = ~\opsel3_pad  & ~n182 ;
  assign n184 = ~n180 & n183 ;
  assign n185 = ~n181 & n184 ;
  assign n186 = ~n174 & ~n185 ;
  assign n187 = \inD14_pad  & n79 ;
  assign n188 = \inB14_pad  & n83 ;
  assign n189 = \inD14_pad  & n82 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n81 & ~n190 ;
  assign n192 = ~n187 & ~n191 ;
  assign n193 = \sh2_pad  & ~n192 ;
  assign n194 = \inD10_pad  & n79 ;
  assign n195 = \inB10_pad  & n83 ;
  assign n196 = \inD10_pad  & n82 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = n81 & ~n197 ;
  assign n199 = ~n194 & ~n198 ;
  assign n200 = ~\sh2_pad  & ~n199 ;
  assign n201 = ~n193 & ~n200 ;
  assign n202 = ~\sh1_pad  & ~n201 ;
  assign n203 = \inD12_pad  & n79 ;
  assign n204 = \inB12_pad  & n83 ;
  assign n205 = \inD12_pad  & n82 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = n81 & ~n206 ;
  assign n208 = ~n203 & ~n207 ;
  assign n209 = ~\sh2_pad  & ~n208 ;
  assign n210 = \inD15_pad  & n79 ;
  assign n211 = \inB15_pad  & n83 ;
  assign n212 = \inD15_pad  & n82 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = n81 & ~n213 ;
  assign n215 = ~n210 & ~n214 ;
  assign n216 = \sh2_pad  & ~n215 ;
  assign n217 = ~n209 & ~n216 ;
  assign n218 = \sh1_pad  & ~n217 ;
  assign n219 = ~n202 & ~n218 ;
  assign n220 = ~\sh0_pad  & ~n219 ;
  assign n231 = \inD11_pad  & n79 ;
  assign n232 = \inB11_pad  & n83 ;
  assign n233 = \inD11_pad  & n82 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = n81 & ~n234 ;
  assign n236 = ~n231 & ~n235 ;
  assign n237 = ~\sh2_pad  & ~n236 ;
  assign n238 = ~n216 & ~n237 ;
  assign n239 = ~\sh1_pad  & n238 ;
  assign n222 = \inD13_pad  & n79 ;
  assign n223 = \inB13_pad  & n83 ;
  assign n224 = \inD13_pad  & n82 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = n81 & ~n225 ;
  assign n227 = ~n222 & ~n226 ;
  assign n228 = ~\sh2_pad  & ~n227 ;
  assign n221 = \sh2_pad  & ~n199 ;
  assign n229 = \sh1_pad  & ~n221 ;
  assign n230 = ~n228 & n229 ;
  assign n240 = \sh0_pad  & ~n230 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = ~n220 & ~n241 ;
  assign n243 = n146 & ~n242 ;
  assign n252 = \opsel2_pad  & ~\opsel3_pad  ;
  assign n253 = \opsel1_pad  & ~n252 ;
  assign n251 = ~\opsel1_pad  & ~n76 ;
  assign n254 = ~\opsel0_pad  & ~n251 ;
  assign n255 = ~n253 & n254 ;
  assign n465 = \inC10_pad  & n79 ;
  assign n466 = \inA10_pad  & n83 ;
  assign n467 = \inC10_pad  & \musel2_pad  ;
  assign n468 = \musel1_pad  & n467 ;
  assign n469 = ~n466 & ~n468 ;
  assign n470 = n81 & ~n469 ;
  assign n471 = ~n465 & ~n470 ;
  assign n472 = ~n255 & ~n471 ;
  assign n473 = n255 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = \inD10_pad  & n150 ;
  assign n476 = \inB10_pad  & n152 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~\musel1_pad  & ~n477 ;
  assign n479 = \inA10_pad  & ~\musel2_pad  ;
  assign n480 = ~n467 & ~n479 ;
  assign n481 = n156 & ~n480 ;
  assign n482 = ~n478 & ~n481 ;
  assign n483 = ~\musel4_pad  & ~n482 ;
  assign n484 = ~n474 & n483 ;
  assign n244 = \inC9_pad  & n79 ;
  assign n245 = \inA9_pad  & n83 ;
  assign n246 = \inC9_pad  & \musel2_pad  ;
  assign n247 = \musel1_pad  & n246 ;
  assign n248 = ~n245 & ~n247 ;
  assign n249 = n81 & ~n248 ;
  assign n250 = ~n244 & ~n249 ;
  assign n256 = ~n250 & ~n255 ;
  assign n257 = n250 & n255 ;
  assign n258 = ~n256 & ~n257 ;
  assign n259 = \inD9_pad  & n150 ;
  assign n260 = \inB9_pad  & n152 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = ~\musel1_pad  & ~n261 ;
  assign n263 = \inA9_pad  & ~\musel2_pad  ;
  assign n264 = ~n246 & ~n263 ;
  assign n265 = n156 & ~n264 ;
  assign n266 = ~n262 & ~n265 ;
  assign n267 = ~\musel4_pad  & ~n266 ;
  assign n268 = n258 & ~n267 ;
  assign n269 = ~n258 & n267 ;
  assign n270 = \inC8_pad  & n79 ;
  assign n271 = \inA8_pad  & n83 ;
  assign n272 = \inC8_pad  & \musel2_pad  ;
  assign n273 = \musel1_pad  & n272 ;
  assign n274 = ~n271 & ~n273 ;
  assign n275 = n81 & ~n274 ;
  assign n276 = ~n270 & ~n275 ;
  assign n277 = ~n255 & ~n276 ;
  assign n278 = n255 & n276 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = \inD8_pad  & n150 ;
  assign n281 = \inB8_pad  & n152 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = ~\musel1_pad  & ~n282 ;
  assign n284 = \inA8_pad  & ~\musel2_pad  ;
  assign n285 = ~n272 & ~n284 ;
  assign n286 = n156 & ~n285 ;
  assign n287 = ~n283 & ~n286 ;
  assign n288 = ~\musel4_pad  & ~n287 ;
  assign n289 = n279 & ~n288 ;
  assign n290 = ~n279 & n288 ;
  assign n291 = \inC4_pad  & n79 ;
  assign n293 = \inC4_pad  & \musel2_pad  ;
  assign n294 = ~n83 & ~n293 ;
  assign n292 = ~\inA4_pad  & n83 ;
  assign n295 = n81 & ~n292 ;
  assign n296 = ~n294 & n295 ;
  assign n297 = ~n291 & ~n296 ;
  assign n298 = ~n255 & ~n297 ;
  assign n299 = n255 & n297 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = \inD4_pad  & n150 ;
  assign n302 = \inB4_pad  & n152 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~\musel1_pad  & ~n303 ;
  assign n305 = \inA4_pad  & ~\musel2_pad  ;
  assign n306 = ~n293 & ~n305 ;
  assign n307 = n156 & ~n306 ;
  assign n308 = ~n304 & ~n307 ;
  assign n309 = ~\musel4_pad  & ~n308 ;
  assign n310 = n300 & ~n309 ;
  assign n331 = \inC2_pad  & n79 ;
  assign n332 = \inA2_pad  & n83 ;
  assign n333 = \inC2_pad  & \musel2_pad  ;
  assign n334 = \musel1_pad  & n333 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = n81 & ~n335 ;
  assign n337 = ~n331 & ~n336 ;
  assign n338 = ~n255 & ~n337 ;
  assign n339 = n255 & n337 ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = \inD2_pad  & n150 ;
  assign n342 = \inB2_pad  & n152 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = ~\musel1_pad  & ~n343 ;
  assign n345 = \inA2_pad  & ~\musel2_pad  ;
  assign n346 = ~n333 & ~n345 ;
  assign n347 = n156 & ~n346 ;
  assign n348 = ~n344 & ~n347 ;
  assign n349 = ~\musel4_pad  & ~n348 ;
  assign n350 = n340 & ~n349 ;
  assign n311 = \inC3_pad  & n79 ;
  assign n312 = \inA3_pad  & n83 ;
  assign n313 = \inC3_pad  & \musel2_pad  ;
  assign n314 = \musel1_pad  & n313 ;
  assign n315 = ~n312 & ~n314 ;
  assign n316 = n81 & ~n315 ;
  assign n317 = ~n311 & ~n316 ;
  assign n318 = ~n255 & ~n317 ;
  assign n319 = n255 & n317 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = \inD3_pad  & n150 ;
  assign n322 = \inB3_pad  & n152 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = ~\musel1_pad  & ~n323 ;
  assign n325 = \inA3_pad  & ~\musel2_pad  ;
  assign n326 = ~n313 & ~n325 ;
  assign n327 = n156 & ~n326 ;
  assign n328 = ~n324 & ~n327 ;
  assign n329 = ~\musel4_pad  & ~n328 ;
  assign n351 = n320 & ~n329 ;
  assign n352 = ~n350 & ~n351 ;
  assign n379 = n168 & ~n255 ;
  assign n378 = ~n168 & n255 ;
  assign n380 = n162 & ~n378 ;
  assign n381 = ~n379 & n380 ;
  assign n376 = ~n340 & n349 ;
  assign n353 = \inC1_pad  & n79 ;
  assign n354 = \inA1_pad  & n83 ;
  assign n355 = \inC1_pad  & \musel2_pad  ;
  assign n356 = \musel1_pad  & n355 ;
  assign n357 = ~n354 & ~n356 ;
  assign n358 = n81 & ~n357 ;
  assign n359 = ~n353 & ~n358 ;
  assign n360 = ~n255 & ~n359 ;
  assign n361 = n255 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = \inD1_pad  & n150 ;
  assign n364 = \inB1_pad  & n152 ;
  assign n365 = ~n363 & ~n364 ;
  assign n366 = ~\musel1_pad  & ~n365 ;
  assign n367 = \inA1_pad  & ~\musel2_pad  ;
  assign n368 = ~n355 & ~n367 ;
  assign n369 = n156 & ~n368 ;
  assign n370 = ~n366 & ~n369 ;
  assign n371 = ~\musel4_pad  & ~n370 ;
  assign n377 = ~n362 & n371 ;
  assign n382 = ~n376 & ~n377 ;
  assign n383 = ~n381 & n382 ;
  assign n384 = n352 & ~n383 ;
  assign n330 = ~n320 & n329 ;
  assign n372 = n362 & ~n371 ;
  assign n373 = ~n169 & n255 ;
  assign n374 = ~n372 & n373 ;
  assign n375 = n352 & n374 ;
  assign n385 = ~n330 & ~n375 ;
  assign n386 = ~n384 & n385 ;
  assign n387 = ~n310 & ~n386 ;
  assign n388 = \inC6_pad  & n79 ;
  assign n390 = \inC6_pad  & \musel2_pad  ;
  assign n391 = ~n83 & ~n390 ;
  assign n389 = ~\inA6_pad  & n83 ;
  assign n392 = n81 & ~n389 ;
  assign n393 = ~n391 & n392 ;
  assign n394 = ~n388 & ~n393 ;
  assign n395 = ~n255 & ~n394 ;
  assign n396 = n255 & n394 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = \inD6_pad  & n150 ;
  assign n399 = \inB6_pad  & n152 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = ~\musel1_pad  & ~n400 ;
  assign n402 = \inA6_pad  & ~\musel2_pad  ;
  assign n403 = ~n390 & ~n402 ;
  assign n404 = n156 & ~n403 ;
  assign n405 = ~n401 & ~n404 ;
  assign n406 = ~\musel4_pad  & ~n405 ;
  assign n407 = n397 & ~n406 ;
  assign n408 = \inC7_pad  & n79 ;
  assign n410 = \inC7_pad  & \musel2_pad  ;
  assign n411 = ~n83 & ~n410 ;
  assign n409 = ~\inA7_pad  & n83 ;
  assign n412 = n81 & ~n409 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n408 & ~n413 ;
  assign n415 = ~n255 & ~n414 ;
  assign n416 = n255 & n414 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = \inD7_pad  & n150 ;
  assign n419 = \inB7_pad  & n152 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~\musel1_pad  & ~n420 ;
  assign n422 = \inA7_pad  & ~\musel2_pad  ;
  assign n423 = ~n410 & ~n422 ;
  assign n424 = n156 & ~n423 ;
  assign n425 = ~n421 & ~n424 ;
  assign n426 = ~\musel4_pad  & ~n425 ;
  assign n427 = n417 & ~n426 ;
  assign n428 = ~n407 & ~n427 ;
  assign n429 = \inC5_pad  & n79 ;
  assign n431 = \inC5_pad  & \musel2_pad  ;
  assign n432 = ~n83 & ~n431 ;
  assign n430 = ~\inA5_pad  & n83 ;
  assign n433 = n81 & ~n430 ;
  assign n434 = ~n432 & n433 ;
  assign n435 = ~n429 & ~n434 ;
  assign n436 = ~n255 & ~n435 ;
  assign n437 = n255 & n435 ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = \inD5_pad  & n150 ;
  assign n440 = \inB5_pad  & n152 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~\musel1_pad  & ~n441 ;
  assign n443 = \inA5_pad  & ~\musel2_pad  ;
  assign n444 = ~n431 & ~n443 ;
  assign n445 = n156 & ~n444 ;
  assign n446 = ~n442 & ~n445 ;
  assign n447 = ~\musel4_pad  & ~n446 ;
  assign n448 = n438 & ~n447 ;
  assign n449 = n428 & ~n448 ;
  assign n450 = n387 & n449 ;
  assign n451 = ~n417 & n426 ;
  assign n452 = ~n300 & n309 ;
  assign n453 = ~n448 & n452 ;
  assign n454 = ~n438 & n447 ;
  assign n455 = ~n397 & n406 ;
  assign n456 = ~n454 & ~n455 ;
  assign n457 = ~n453 & n456 ;
  assign n458 = n428 & ~n457 ;
  assign n459 = ~n451 & ~n458 ;
  assign n460 = ~n450 & n459 ;
  assign n461 = ~n290 & n460 ;
  assign n462 = ~n289 & ~n461 ;
  assign n463 = ~n269 & ~n462 ;
  assign n464 = ~n268 & ~n463 ;
  assign n485 = n474 & ~n483 ;
  assign n488 = n464 & ~n485 ;
  assign n489 = ~n484 & n488 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~n464 & ~n486 ;
  assign n490 = n149 & ~n487 ;
  assign n491 = ~n489 & n490 ;
  assign n492 = ~n243 & ~n491 ;
  assign n493 = n76 & ~n492 ;
  assign n552 = n175 & n242 ;
  assign n494 = \inA15_pad  & ~\musel2_pad  ;
  assign n495 = \inC15_pad  & ~\musel1_pad  ;
  assign n496 = ~n494 & ~n495 ;
  assign n497 = ~n78 & n496 ;
  assign n498 = \inC10_pad  & ~\musel1_pad  ;
  assign n499 = ~n479 & ~n498 ;
  assign n500 = n497 & ~n499 ;
  assign n501 = ~n78 & ~n496 ;
  assign n502 = n499 & n501 ;
  assign n503 = ~n500 & ~n502 ;
  assign n514 = \inC2_pad  & ~\musel1_pad  ;
  assign n515 = ~n345 & ~n514 ;
  assign n517 = n496 & n515 ;
  assign n516 = ~n496 & ~n515 ;
  assign n518 = n178 & ~n516 ;
  assign n519 = ~n517 & n518 ;
  assign n520 = \inC3_pad  & ~\musel1_pad  ;
  assign n521 = ~n325 & ~n520 ;
  assign n522 = n497 & ~n521 ;
  assign n523 = n501 & n521 ;
  assign n524 = ~n522 & ~n523 ;
  assign n534 = n519 & ~n524 ;
  assign n525 = n178 & ~n496 ;
  assign n526 = n177 & n525 ;
  assign n527 = n179 & ~n521 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = \inC1_pad  & ~\musel1_pad  ;
  assign n530 = ~n367 & ~n529 ;
  assign n531 = n501 & n530 ;
  assign n532 = n497 & ~n530 ;
  assign n533 = ~n531 & ~n532 ;
  assign n535 = ~n528 & ~n533 ;
  assign n536 = n534 & n535 ;
  assign n504 = \inC9_pad  & ~\musel1_pad  ;
  assign n505 = ~n263 & ~n504 ;
  assign n506 = n497 & ~n505 ;
  assign n507 = n501 & n505 ;
  assign n508 = ~n506 & ~n507 ;
  assign n544 = ~n503 & ~n508 ;
  assign n509 = \inC8_pad  & ~\musel1_pad  ;
  assign n510 = ~n284 & ~n509 ;
  assign n511 = n497 & ~n510 ;
  assign n512 = n501 & n510 ;
  assign n513 = ~n511 & ~n512 ;
  assign n537 = \inA11_pad  & ~\musel2_pad  ;
  assign n538 = \inC11_pad  & ~\musel1_pad  ;
  assign n539 = ~n537 & ~n538 ;
  assign n541 = n501 & ~n539 ;
  assign n540 = n496 & n539 ;
  assign n542 = n178 & ~n540 ;
  assign n543 = ~n541 & n542 ;
  assign n545 = ~n513 & n543 ;
  assign n546 = n544 & n545 ;
  assign n547 = n536 & n546 ;
  assign n548 = n501 & n547 ;
  assign n549 = n77 & ~n548 ;
  assign n550 = ~n503 & n549 ;
  assign n551 = ~n175 & ~n550 ;
  assign n553 = n183 & ~n551 ;
  assign n554 = ~n552 & n553 ;
  assign n555 = ~n493 & ~n554 ;
  assign n556 = \sh0_pad  & \sh1_pad  ;
  assign n557 = n215 & ~n556 ;
  assign n558 = n236 & n556 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = \sh2_pad  & ~n559 ;
  assign n565 = ~\sh1_pad  & ~n236 ;
  assign n566 = \sh1_pad  & ~n227 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~\sh0_pad  & ~n567 ;
  assign n561 = \sh1_pad  & ~n192 ;
  assign n562 = ~\sh1_pad  & ~n208 ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = \sh0_pad  & ~n563 ;
  assign n569 = ~\sh2_pad  & ~n564 ;
  assign n570 = ~n568 & n569 ;
  assign n571 = ~n560 & ~n570 ;
  assign n572 = n146 & n571 ;
  assign n573 = \inC11_pad  & n79 ;
  assign n574 = \inA11_pad  & n83 ;
  assign n575 = \inC11_pad  & \musel2_pad  ;
  assign n576 = \musel1_pad  & n575 ;
  assign n577 = ~n574 & ~n576 ;
  assign n578 = n81 & ~n577 ;
  assign n579 = ~n573 & ~n578 ;
  assign n580 = ~n255 & ~n579 ;
  assign n581 = n255 & n579 ;
  assign n582 = ~n580 & ~n581 ;
  assign n583 = \inD11_pad  & n150 ;
  assign n584 = \inB11_pad  & n152 ;
  assign n585 = ~n583 & ~n584 ;
  assign n586 = ~\musel1_pad  & ~n585 ;
  assign n587 = ~n537 & ~n575 ;
  assign n588 = n156 & ~n587 ;
  assign n589 = ~n586 & ~n588 ;
  assign n590 = ~\musel4_pad  & ~n589 ;
  assign n591 = n582 & ~n590 ;
  assign n592 = ~n582 & n590 ;
  assign n593 = ~n591 & ~n592 ;
  assign n595 = ~n484 & ~n593 ;
  assign n596 = ~n488 & n595 ;
  assign n594 = n488 & n593 ;
  assign n597 = n149 & ~n594 ;
  assign n598 = ~n596 & n597 ;
  assign n599 = ~n572 & ~n598 ;
  assign n600 = n76 & ~n599 ;
  assign n603 = n175 & ~n571 ;
  assign n601 = n543 & ~n548 ;
  assign n602 = ~n175 & ~n601 ;
  assign n604 = n183 & ~n602 ;
  assign n605 = ~n603 & n604 ;
  assign n606 = ~n600 & ~n605 ;
  assign n608 = ~\sh0_pad  & ~n563 ;
  assign n607 = ~n215 & n556 ;
  assign n609 = \sh0_pad  & ~\sh1_pad  ;
  assign n610 = ~n227 & n609 ;
  assign n611 = ~n607 & ~n610 ;
  assign n612 = ~n608 & n611 ;
  assign n613 = ~\sh2_pad  & ~n612 ;
  assign n614 = n208 & n556 ;
  assign n615 = \sh2_pad  & ~n557 ;
  assign n616 = ~n614 & n615 ;
  assign n617 = ~n613 & ~n616 ;
  assign n618 = n146 & ~n617 ;
  assign n619 = \inC12_pad  & n79 ;
  assign n620 = \inA12_pad  & n83 ;
  assign n621 = \inC12_pad  & \musel2_pad  ;
  assign n622 = \musel1_pad  & n621 ;
  assign n623 = ~n620 & ~n622 ;
  assign n624 = n81 & ~n623 ;
  assign n625 = ~n619 & ~n624 ;
  assign n626 = ~n255 & ~n625 ;
  assign n627 = n255 & n625 ;
  assign n628 = ~n626 & ~n627 ;
  assign n629 = \inD12_pad  & n150 ;
  assign n630 = \inB12_pad  & n152 ;
  assign n631 = ~n629 & ~n630 ;
  assign n632 = ~\musel1_pad  & ~n631 ;
  assign n633 = \inA12_pad  & ~\musel2_pad  ;
  assign n634 = ~n621 & ~n633 ;
  assign n635 = n156 & ~n634 ;
  assign n636 = ~n632 & ~n635 ;
  assign n637 = ~\musel4_pad  & ~n636 ;
  assign n638 = n628 & ~n637 ;
  assign n639 = ~n628 & n637 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = ~n268 & ~n289 ;
  assign n642 = ~n485 & ~n591 ;
  assign n643 = n641 & n642 ;
  assign n644 = ~n460 & n643 ;
  assign n646 = n640 & n644 ;
  assign n645 = ~n640 & ~n644 ;
  assign n647 = n149 & ~n645 ;
  assign n648 = ~n646 & n647 ;
  assign n649 = ~n618 & ~n648 ;
  assign n650 = n76 & ~n649 ;
  assign n682 = n175 & n617 ;
  assign n659 = \inC5_pad  & ~\musel1_pad  ;
  assign n660 = ~n443 & ~n659 ;
  assign n662 = n501 & ~n660 ;
  assign n661 = n496 & n660 ;
  assign n663 = n178 & ~n661 ;
  assign n664 = ~n662 & n663 ;
  assign n651 = \inC4_pad  & ~\musel1_pad  ;
  assign n652 = ~n305 & ~n651 ;
  assign n653 = n497 & ~n652 ;
  assign n654 = n501 & n652 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = \inC6_pad  & ~\musel1_pad  ;
  assign n657 = ~n402 & ~n656 ;
  assign n658 = ~n78 & ~n657 ;
  assign n665 = \inC7_pad  & ~\musel1_pad  ;
  assign n666 = ~n422 & ~n665 ;
  assign n667 = n525 & n666 ;
  assign n668 = ~n658 & n667 ;
  assign n669 = ~n655 & n668 ;
  assign n670 = n664 & n669 ;
  assign n671 = n547 & n670 ;
  assign n672 = \inC12_pad  & ~\musel1_pad  ;
  assign n673 = ~n633 & ~n672 ;
  assign n675 = n501 & ~n673 ;
  assign n674 = n496 & n673 ;
  assign n676 = n178 & ~n674 ;
  assign n677 = ~n675 & n676 ;
  assign n678 = n671 & n677 ;
  assign n679 = ~n671 & ~n677 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = ~n175 & ~n680 ;
  assign n683 = n183 & ~n681 ;
  assign n684 = ~n682 & n683 ;
  assign n685 = ~n650 & ~n684 ;
  assign n692 = \sh0_pad  & n192 ;
  assign n688 = ~\sh1_pad  & ~\sh2_pad  ;
  assign n691 = ~\sh0_pad  & n227 ;
  assign n693 = n688 & ~n691 ;
  assign n694 = ~n692 & n693 ;
  assign n686 = \sh2_pad  & n556 ;
  assign n687 = ~n227 & n686 ;
  assign n689 = ~n686 & ~n688 ;
  assign n690 = ~n215 & n689 ;
  assign n695 = ~n687 & ~n690 ;
  assign n696 = ~n694 & n695 ;
  assign n697 = n146 & ~n696 ;
  assign n698 = \inC13_pad  & n79 ;
  assign n699 = \inA13_pad  & n83 ;
  assign n700 = \inC13_pad  & \musel2_pad  ;
  assign n701 = \musel1_pad  & n700 ;
  assign n702 = ~n699 & ~n701 ;
  assign n703 = n81 & ~n702 ;
  assign n704 = ~n698 & ~n703 ;
  assign n705 = ~n255 & ~n704 ;
  assign n706 = n255 & n704 ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = \inD13_pad  & n150 ;
  assign n709 = \inB13_pad  & n152 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = ~\musel1_pad  & ~n710 ;
  assign n712 = \inA13_pad  & ~\musel2_pad  ;
  assign n713 = ~n700 & ~n712 ;
  assign n714 = n156 & ~n713 ;
  assign n715 = ~n711 & ~n714 ;
  assign n716 = ~\musel4_pad  & ~n715 ;
  assign n717 = n707 & ~n716 ;
  assign n718 = ~n707 & n716 ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = ~n638 & n644 ;
  assign n721 = ~n639 & ~n720 ;
  assign n722 = ~n719 & n721 ;
  assign n723 = n719 & n720 ;
  assign n724 = n149 & ~n723 ;
  assign n725 = ~n722 & n724 ;
  assign n726 = ~n697 & ~n725 ;
  assign n727 = n76 & ~n726 ;
  assign n729 = \inC13_pad  & ~\musel1_pad  ;
  assign n730 = ~n712 & ~n729 ;
  assign n731 = n497 & ~n730 ;
  assign n732 = n501 & n730 ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = n77 & ~n733 ;
  assign n735 = ~n678 & ~n734 ;
  assign n736 = n678 & ~n733 ;
  assign n737 = ~n735 & ~n736 ;
  assign n738 = ~n175 & ~n737 ;
  assign n728 = n175 & n696 ;
  assign n739 = n183 & ~n728 ;
  assign n740 = ~n738 & n739 ;
  assign n741 = ~n727 & ~n740 ;
  assign n742 = ~n717 & n720 ;
  assign n743 = \inC14_pad  & n79 ;
  assign n744 = \inA14_pad  & n83 ;
  assign n745 = \inC14_pad  & \musel2_pad  ;
  assign n746 = \musel1_pad  & n745 ;
  assign n747 = ~n744 & ~n746 ;
  assign n748 = n81 & ~n747 ;
  assign n749 = ~n743 & ~n748 ;
  assign n750 = ~n255 & ~n749 ;
  assign n751 = n255 & n749 ;
  assign n752 = ~n750 & ~n751 ;
  assign n753 = \inD14_pad  & n150 ;
  assign n754 = \inB14_pad  & n152 ;
  assign n755 = ~n753 & ~n754 ;
  assign n756 = ~\musel1_pad  & ~n755 ;
  assign n757 = \inA14_pad  & ~\musel2_pad  ;
  assign n758 = ~n745 & ~n757 ;
  assign n759 = n156 & ~n758 ;
  assign n760 = ~n756 & ~n759 ;
  assign n761 = ~\musel4_pad  & ~n760 ;
  assign n762 = n752 & ~n761 ;
  assign n763 = ~n752 & n761 ;
  assign n764 = ~n762 & ~n763 ;
  assign n765 = ~n718 & n764 ;
  assign n766 = ~n742 & n765 ;
  assign n767 = ~n718 & n721 ;
  assign n768 = ~n717 & ~n764 ;
  assign n769 = ~n767 & n768 ;
  assign n770 = ~n766 & ~n769 ;
  assign n771 = n149 & ~n770 ;
  assign n772 = \sh0_pad  & \sh2_pad  ;
  assign n773 = ~n688 & ~n772 ;
  assign n774 = ~n609 & ~n773 ;
  assign n775 = ~n192 & n774 ;
  assign n776 = ~n215 & ~n774 ;
  assign n777 = ~n775 & ~n776 ;
  assign n778 = n146 & ~n777 ;
  assign n779 = ~n771 & ~n778 ;
  assign n780 = n76 & ~n779 ;
  assign n782 = \inC14_pad  & ~\musel1_pad  ;
  assign n783 = ~n757 & ~n782 ;
  assign n785 = n501 & ~n783 ;
  assign n784 = n496 & n783 ;
  assign n786 = n178 & ~n784 ;
  assign n787 = ~n785 & n786 ;
  assign n788 = n736 & n787 ;
  assign n789 = ~n736 & ~n787 ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = ~n175 & ~n790 ;
  assign n781 = n175 & n777 ;
  assign n792 = n183 & ~n781 ;
  assign n793 = ~n791 & n792 ;
  assign n794 = ~n780 & ~n793 ;
  assign n795 = n146 & ~n215 ;
  assign n796 = ~n762 & ~n766 ;
  assign n797 = \inC15_pad  & n79 ;
  assign n798 = \inA15_pad  & n83 ;
  assign n799 = \inC15_pad  & \musel2_pad  ;
  assign n800 = \musel1_pad  & n799 ;
  assign n801 = ~n798 & ~n800 ;
  assign n802 = n81 & ~n801 ;
  assign n803 = ~n797 & ~n802 ;
  assign n804 = \inD15_pad  & n150 ;
  assign n805 = \inB15_pad  & n152 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = ~\musel1_pad  & ~n806 ;
  assign n808 = ~n494 & ~n799 ;
  assign n809 = n156 & ~n808 ;
  assign n810 = ~n807 & ~n809 ;
  assign n811 = ~\musel4_pad  & ~n810 ;
  assign n812 = n803 & ~n811 ;
  assign n813 = ~n803 & n811 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = n255 & n814 ;
  assign n816 = ~n255 & ~n814 ;
  assign n817 = ~n815 & ~n816 ;
  assign n820 = n796 & n817 ;
  assign n818 = ~n763 & ~n817 ;
  assign n819 = ~n796 & n818 ;
  assign n821 = n149 & ~n819 ;
  assign n822 = ~n820 & n821 ;
  assign n823 = ~n795 & ~n822 ;
  assign n824 = n76 & ~n823 ;
  assign n826 = ~n175 & ~n788 ;
  assign n825 = n175 & n215 ;
  assign n827 = n183 & ~n825 ;
  assign n828 = ~n826 & n827 ;
  assign n829 = ~n824 & ~n828 ;
  assign n830 = \inD9_pad  & n79 ;
  assign n831 = \inB9_pad  & n83 ;
  assign n832 = \inD9_pad  & n82 ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = n81 & ~n833 ;
  assign n835 = ~n830 & ~n834 ;
  assign n836 = \sh2_pad  & ~n835 ;
  assign n837 = ~n89 & ~n836 ;
  assign n838 = \sh1_pad  & ~n837 ;
  assign n839 = ~n114 & ~n838 ;
  assign n840 = ~\sh0_pad  & ~n839 ;
  assign n841 = \inD6_pad  & n79 ;
  assign n842 = \inB6_pad  & n83 ;
  assign n843 = \inD6_pad  & n82 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = n81 & ~n844 ;
  assign n846 = ~n841 & ~n845 ;
  assign n847 = \sh2_pad  & ~n846 ;
  assign n848 = ~n130 & ~n847 ;
  assign n849 = ~\sh1_pad  & ~n848 ;
  assign n850 = ~\sh2_pad  & ~n139 ;
  assign n851 = \sh2_pad  & ~n111 ;
  assign n852 = ~n850 & ~n851 ;
  assign n853 = \sh1_pad  & ~n852 ;
  assign n854 = ~n849 & ~n853 ;
  assign n855 = \sh0_pad  & ~n854 ;
  assign n856 = ~n840 & ~n855 ;
  assign n857 = n146 & ~n856 ;
  assign n858 = ~n372 & ~n377 ;
  assign n859 = ~n169 & ~n379 ;
  assign n861 = n858 & n859 ;
  assign n860 = ~n858 & ~n859 ;
  assign n862 = n149 & ~n860 ;
  assign n863 = ~n861 & n862 ;
  assign n864 = ~n857 & ~n863 ;
  assign n865 = n76 & ~n864 ;
  assign n866 = n175 & ~n856 ;
  assign n867 = n77 & ~n533 ;
  assign n868 = ~n526 & ~n867 ;
  assign n869 = ~n78 & ~n530 ;
  assign n870 = n526 & ~n869 ;
  assign n871 = ~n175 & ~n870 ;
  assign n872 = ~n868 & n871 ;
  assign n873 = ~n866 & ~n872 ;
  assign n874 = n183 & ~n873 ;
  assign n875 = ~n865 & ~n874 ;
  assign n876 = ~n221 & ~n850 ;
  assign n877 = \sh1_pad  & ~n876 ;
  assign n878 = ~n849 & ~n877 ;
  assign n879 = ~\sh0_pad  & ~n878 ;
  assign n880 = \inD7_pad  & n79 ;
  assign n881 = \inB7_pad  & n83 ;
  assign n882 = \inD7_pad  & n82 ;
  assign n883 = ~n881 & ~n882 ;
  assign n884 = n81 & ~n883 ;
  assign n885 = ~n880 & ~n884 ;
  assign n886 = \sh2_pad  & ~n885 ;
  assign n887 = ~n89 & ~n886 ;
  assign n888 = ~\sh1_pad  & ~n887 ;
  assign n889 = ~\sh2_pad  & ~n104 ;
  assign n890 = \sh2_pad  & ~n129 ;
  assign n891 = ~n889 & ~n890 ;
  assign n892 = \sh1_pad  & ~n891 ;
  assign n893 = ~n888 & ~n892 ;
  assign n894 = \sh0_pad  & ~n893 ;
  assign n895 = ~n879 & ~n894 ;
  assign n896 = n146 & ~n895 ;
  assign n897 = ~n350 & ~n376 ;
  assign n898 = ~n372 & n859 ;
  assign n900 = ~n377 & ~n898 ;
  assign n901 = ~n897 & n900 ;
  assign n899 = n897 & n898 ;
  assign n902 = n149 & ~n899 ;
  assign n903 = ~n901 & n902 ;
  assign n904 = ~n896 & ~n903 ;
  assign n905 = n76 & ~n904 ;
  assign n906 = n175 & ~n895 ;
  assign n908 = n519 & n870 ;
  assign n907 = ~n519 & ~n870 ;
  assign n909 = ~n175 & ~n907 ;
  assign n910 = ~n908 & n909 ;
  assign n911 = ~n906 & ~n910 ;
  assign n912 = n183 & ~n911 ;
  assign n913 = ~n905 & ~n912 ;
  assign n914 = \sh2_pad  & ~n236 ;
  assign n915 = ~n889 & ~n914 ;
  assign n916 = \sh1_pad  & ~n915 ;
  assign n917 = ~n888 & ~n916 ;
  assign n918 = ~\sh0_pad  & ~n917 ;
  assign n919 = ~n123 & ~n850 ;
  assign n920 = ~\sh1_pad  & ~n919 ;
  assign n921 = ~\sh2_pad  & ~n846 ;
  assign n922 = \sh2_pad  & ~n88 ;
  assign n923 = ~n921 & ~n922 ;
  assign n924 = \sh1_pad  & ~n923 ;
  assign n925 = ~n920 & ~n924 ;
  assign n926 = \sh0_pad  & ~n925 ;
  assign n927 = ~n918 & ~n926 ;
  assign n928 = n146 & ~n927 ;
  assign n929 = ~n350 & ~n900 ;
  assign n930 = ~n330 & ~n351 ;
  assign n932 = ~n376 & ~n930 ;
  assign n933 = ~n929 & n932 ;
  assign n931 = n929 & n930 ;
  assign n934 = n149 & ~n931 ;
  assign n935 = ~n933 & n934 ;
  assign n936 = ~n928 & ~n935 ;
  assign n937 = n76 & ~n936 ;
  assign n943 = n175 & n927 ;
  assign n940 = n524 & n908 ;
  assign n938 = n77 & ~n524 ;
  assign n939 = ~n908 & n938 ;
  assign n941 = ~n175 & ~n939 ;
  assign n942 = ~n940 & n941 ;
  assign n944 = n183 & ~n942 ;
  assign n945 = ~n943 & n944 ;
  assign n946 = ~n937 & ~n945 ;
  assign n947 = \sh2_pad  & ~n208 ;
  assign n948 = ~n921 & ~n947 ;
  assign n949 = \sh1_pad  & ~n948 ;
  assign n950 = ~n920 & ~n949 ;
  assign n951 = ~\sh0_pad  & ~n950 ;
  assign n952 = ~n836 & ~n889 ;
  assign n953 = ~\sh1_pad  & ~n952 ;
  assign n954 = ~\sh2_pad  & ~n885 ;
  assign n955 = ~n140 & ~n954 ;
  assign n956 = \sh1_pad  & ~n955 ;
  assign n957 = ~n953 & ~n956 ;
  assign n958 = \sh0_pad  & ~n957 ;
  assign n959 = ~n951 & ~n958 ;
  assign n960 = n146 & ~n959 ;
  assign n961 = ~n310 & ~n452 ;
  assign n963 = n386 & ~n961 ;
  assign n962 = ~n386 & n961 ;
  assign n964 = n149 & ~n962 ;
  assign n965 = ~n963 & n964 ;
  assign n966 = ~n960 & ~n965 ;
  assign n967 = n76 & ~n966 ;
  assign n974 = n175 & n959 ;
  assign n968 = n501 & n536 ;
  assign n969 = n77 & ~n655 ;
  assign n970 = n968 & n969 ;
  assign n971 = ~n968 & ~n969 ;
  assign n972 = ~n970 & ~n971 ;
  assign n973 = ~n175 & ~n972 ;
  assign n975 = n183 & ~n973 ;
  assign n976 = ~n974 & n975 ;
  assign n977 = ~n967 & ~n976 ;
  assign n978 = \sh2_pad  & ~n227 ;
  assign n979 = ~n954 & ~n978 ;
  assign n980 = \sh1_pad  & ~n979 ;
  assign n981 = ~n953 & ~n980 ;
  assign n982 = ~\sh0_pad  & ~n981 ;
  assign n983 = ~n221 & ~n921 ;
  assign n984 = ~\sh1_pad  & ~n983 ;
  assign n985 = ~\sh2_pad  & ~n122 ;
  assign n986 = ~n105 & ~n985 ;
  assign n987 = \sh1_pad  & ~n986 ;
  assign n988 = ~n984 & ~n987 ;
  assign n989 = \sh0_pad  & ~n988 ;
  assign n990 = ~n982 & ~n989 ;
  assign n991 = n146 & ~n990 ;
  assign n992 = ~n448 & ~n454 ;
  assign n995 = n387 & n992 ;
  assign n993 = ~n452 & ~n992 ;
  assign n994 = ~n387 & n993 ;
  assign n996 = n149 & ~n994 ;
  assign n997 = ~n995 & n996 ;
  assign n998 = ~n991 & ~n997 ;
  assign n999 = n76 & ~n998 ;
  assign n1005 = n175 & n990 ;
  assign n1000 = ~n664 & ~n970 ;
  assign n1001 = ~n78 & ~n660 ;
  assign n1002 = n970 & ~n1001 ;
  assign n1003 = ~n1000 & ~n1002 ;
  assign n1004 = ~n175 & ~n1003 ;
  assign n1006 = n183 & ~n1004 ;
  assign n1007 = ~n1005 & n1006 ;
  assign n1008 = ~n999 & ~n1007 ;
  assign n1009 = ~n193 & ~n985 ;
  assign n1010 = \sh1_pad  & ~n1009 ;
  assign n1011 = ~n984 & ~n1010 ;
  assign n1012 = ~\sh0_pad  & ~n1011 ;
  assign n1013 = ~n914 & ~n954 ;
  assign n1014 = ~\sh1_pad  & ~n1013 ;
  assign n1015 = ~\sh2_pad  & ~n835 ;
  assign n1016 = ~n847 & ~n1015 ;
  assign n1017 = \sh1_pad  & ~n1016 ;
  assign n1018 = ~n1014 & ~n1017 ;
  assign n1019 = \sh0_pad  & ~n1018 ;
  assign n1020 = ~n1012 & ~n1019 ;
  assign n1021 = n146 & ~n1020 ;
  assign n1023 = ~n387 & ~n454 ;
  assign n1024 = ~n448 & ~n1023 ;
  assign n1027 = ~n407 & n1024 ;
  assign n1028 = ~n455 & n1027 ;
  assign n1022 = ~n407 & ~n455 ;
  assign n1025 = ~n453 & ~n1022 ;
  assign n1026 = ~n1024 & n1025 ;
  assign n1029 = n149 & ~n1026 ;
  assign n1030 = ~n1028 & n1029 ;
  assign n1031 = ~n1021 & ~n1030 ;
  assign n1032 = n76 & ~n1031 ;
  assign n1035 = n501 & ~n657 ;
  assign n1034 = n496 & n657 ;
  assign n1036 = n178 & ~n1034 ;
  assign n1037 = ~n1035 & n1036 ;
  assign n1038 = n1002 & n1037 ;
  assign n1039 = ~n1002 & ~n1037 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1041 = ~n175 & ~n1040 ;
  assign n1033 = n175 & n1020 ;
  assign n1042 = n183 & ~n1033 ;
  assign n1043 = ~n1041 & n1042 ;
  assign n1044 = ~n1032 & ~n1043 ;
  assign n1045 = ~n216 & ~n1015 ;
  assign n1046 = \sh1_pad  & ~n1045 ;
  assign n1047 = ~n1014 & ~n1046 ;
  assign n1048 = ~\sh0_pad  & ~n1047 ;
  assign n1049 = ~n947 & ~n985 ;
  assign n1050 = ~\sh1_pad  & ~n1049 ;
  assign n1051 = ~n200 & ~n886 ;
  assign n1052 = \sh1_pad  & ~n1051 ;
  assign n1053 = ~n1050 & ~n1052 ;
  assign n1054 = \sh0_pad  & ~n1053 ;
  assign n1055 = ~n1048 & ~n1054 ;
  assign n1056 = n146 & ~n1055 ;
  assign n1057 = ~n427 & ~n451 ;
  assign n1059 = ~n455 & ~n1057 ;
  assign n1060 = ~n1027 & n1059 ;
  assign n1058 = n1027 & n1057 ;
  assign n1061 = n149 & ~n1058 ;
  assign n1062 = ~n1060 & n1061 ;
  assign n1063 = ~n1056 & ~n1062 ;
  assign n1064 = n76 & ~n1063 ;
  assign n1065 = n77 & ~n666 ;
  assign n1066 = n497 & n1065 ;
  assign n1067 = ~n667 & ~n1066 ;
  assign n1068 = n1038 & ~n1067 ;
  assign n1069 = ~n1038 & n1067 ;
  assign n1070 = ~n1068 & ~n1069 ;
  assign n1071 = ~n175 & ~n1070 ;
  assign n1072 = n175 & n1055 ;
  assign n1073 = n183 & ~n1072 ;
  assign n1074 = ~n1071 & n1073 ;
  assign n1075 = ~n1064 & ~n1074 ;
  assign n1076 = ~n200 & ~n216 ;
  assign n1077 = \sh1_pad  & ~n1076 ;
  assign n1078 = ~n1050 & ~n1077 ;
  assign n1079 = ~\sh0_pad  & ~n1078 ;
  assign n1080 = ~n978 & ~n1015 ;
  assign n1081 = ~\sh1_pad  & ~n1080 ;
  assign n1082 = ~n123 & ~n237 ;
  assign n1083 = \sh1_pad  & ~n1082 ;
  assign n1084 = ~n1081 & ~n1083 ;
  assign n1085 = \sh0_pad  & ~n1084 ;
  assign n1086 = ~n1079 & ~n1085 ;
  assign n1087 = n146 & ~n1086 ;
  assign n1088 = ~n289 & ~n290 ;
  assign n1090 = n460 & ~n1088 ;
  assign n1089 = ~n460 & n1088 ;
  assign n1091 = n149 & ~n1089 ;
  assign n1092 = ~n1090 & n1091 ;
  assign n1093 = ~n1087 & ~n1092 ;
  assign n1094 = n76 & ~n1093 ;
  assign n1095 = n175 & ~n1086 ;
  assign n1096 = ~n175 & n549 ;
  assign n1097 = ~n513 & n1096 ;
  assign n1098 = ~n1095 & ~n1097 ;
  assign n1099 = n183 & ~n1098 ;
  assign n1100 = ~n1094 & ~n1099 ;
  assign n1101 = \sh1_pad  & ~n238 ;
  assign n1102 = ~n1081 & ~n1101 ;
  assign n1103 = ~\sh0_pad  & ~n1102 ;
  assign n1104 = ~n209 & ~n836 ;
  assign n1105 = \sh1_pad  & ~n1104 ;
  assign n1106 = ~n202 & ~n1105 ;
  assign n1107 = \sh0_pad  & ~n1106 ;
  assign n1108 = ~n1103 & ~n1107 ;
  assign n1109 = n146 & ~n1108 ;
  assign n1110 = ~n268 & ~n269 ;
  assign n1112 = n462 & n1110 ;
  assign n1111 = ~n462 & ~n1110 ;
  assign n1113 = n149 & ~n1111 ;
  assign n1114 = ~n1112 & n1113 ;
  assign n1115 = ~n1109 & ~n1114 ;
  assign n1116 = n76 & ~n1115 ;
  assign n1117 = n175 & ~n1108 ;
  assign n1118 = ~n508 & n1096 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n183 & ~n1119 ;
  assign n1121 = ~n1116 & ~n1120 ;
  assign \O0_pad  = ~n186 ;
  assign \O10_pad  = ~n555 ;
  assign \O11_pad  = ~n606 ;
  assign \O12_pad  = ~n685 ;
  assign \O13_pad  = ~n741 ;
  assign \O14_pad  = ~n794 ;
  assign \O15_pad  = ~n829 ;
  assign \O1_pad  = ~n875 ;
  assign \O2_pad  = ~n913 ;
  assign \O3_pad  = ~n946 ;
  assign \O4_pad  = ~n977 ;
  assign \O5_pad  = ~n1008 ;
  assign \O6_pad  = ~n1044 ;
  assign \O7_pad  = ~n1075 ;
  assign \O8_pad  = ~n1100 ;
  assign \O9_pad  = ~n1121 ;
endmodule
