module top (\B_reg/NET0131 , \IR_reg[0]/NET0131 , \IR_reg[10]/NET0131 , \IR_reg[11]/NET0131 , \IR_reg[12]/NET0131 , \IR_reg[13]/NET0131 , \IR_reg[14]/NET0131 , \IR_reg[15]/NET0131 , \IR_reg[16]/NET0131 , \IR_reg[17]/NET0131 , \IR_reg[18]/NET0131 , \IR_reg[19]/NET0131 , \IR_reg[1]/NET0131 , \IR_reg[20]/NET0131 , \IR_reg[21]/NET0131 , \IR_reg[22]/NET0131 , \IR_reg[23]/NET0131 , \IR_reg[24]/NET0131 , \IR_reg[25]/NET0131 , \IR_reg[26]/NET0131 , \IR_reg[27]/NET0131 , \IR_reg[28]/NET0131 , \IR_reg[29]/NET0131 , \IR_reg[2]/NET0131 , \IR_reg[30]/NET0131 , \IR_reg[31]/NET0131 , \IR_reg[3]/NET0131 , \IR_reg[4]/NET0131 , \IR_reg[5]/NET0131 , \IR_reg[6]/NET0131 , \IR_reg[7]/NET0131 , \IR_reg[8]/NET0131 , \IR_reg[9]/NET0131 , \addr[0]_pad , \addr[10]_pad , \addr[11]_pad , \addr[12]_pad , \addr[13]_pad , \addr[14]_pad , \addr[15]_pad , \addr[16]_pad , \addr[17]_pad , \addr[18]_pad , \addr[19]_pad , \addr[1]_pad , \addr[2]_pad , \addr[3]_pad , \addr[4]_pad , \addr[5]_pad , \addr[6]_pad , \addr[7]_pad , \addr[8]_pad , \addr[9]_pad , \d_reg[0]/NET0131 , \d_reg[1]/NET0131 , \datai[0]_pad , \datai[10]_pad , \datai[11]_pad , \datai[12]_pad , \datai[13]_pad , \datai[14]_pad , \datai[15]_pad , \datai[16]_pad , \datai[17]_pad , \datai[18]_pad , \datai[19]_pad , \datai[1]_pad , \datai[20]_pad , \datai[21]_pad , \datai[22]_pad , \datai[23]_pad , \datai[24]_pad , \datai[25]_pad , \datai[26]_pad , \datai[27]_pad , \datai[28]_pad , \datai[29]_pad , \datai[2]_pad , \datai[30]_pad , \datai[31]_pad , \datai[3]_pad , \datai[4]_pad , \datai[5]_pad , \datai[6]_pad , \datai[7]_pad , \datai[8]_pad , \datai[9]_pad , \reg0_reg[0]/NET0131 , \reg0_reg[10]/NET0131 , \reg0_reg[11]/NET0131 , \reg0_reg[12]/NET0131 , \reg0_reg[13]/NET0131 , \reg0_reg[14]/NET0131 , \reg0_reg[15]/NET0131 , \reg0_reg[16]/NET0131 , \reg0_reg[17]/NET0131 , \reg0_reg[18]/NET0131 , \reg0_reg[19]/NET0131 , \reg0_reg[1]/NET0131 , \reg0_reg[20]/NET0131 , \reg0_reg[21]/NET0131 , \reg0_reg[22]/NET0131 , \reg0_reg[23]/NET0131 , \reg0_reg[24]/NET0131 , \reg0_reg[25]/NET0131 , \reg0_reg[26]/NET0131 , \reg0_reg[27]/NET0131 , \reg0_reg[28]/NET0131 , \reg0_reg[29]/NET0131 , \reg0_reg[2]/NET0131 , \reg0_reg[30]/NET0131 , \reg0_reg[31]/NET0131 , \reg0_reg[3]/NET0131 , \reg0_reg[4]/NET0131 , \reg0_reg[5]/NET0131 , \reg0_reg[6]/NET0131 , \reg0_reg[7]/NET0131 , \reg0_reg[8]/NET0131 , \reg0_reg[9]/NET0131 , \reg1_reg[0]/NET0131 , \reg1_reg[10]/NET0131 , \reg1_reg[11]/NET0131 , \reg1_reg[12]/NET0131 , \reg1_reg[13]/NET0131 , \reg1_reg[14]/NET0131 , \reg1_reg[15]/NET0131 , \reg1_reg[16]/NET0131 , \reg1_reg[17]/NET0131 , \reg1_reg[18]/NET0131 , \reg1_reg[19]/NET0131 , \reg1_reg[1]/NET0131 , \reg1_reg[20]/NET0131 , \reg1_reg[21]/NET0131 , \reg1_reg[22]/NET0131 , \reg1_reg[23]/NET0131 , \reg1_reg[24]/NET0131 , \reg1_reg[25]/NET0131 , \reg1_reg[26]/NET0131 , \reg1_reg[27]/NET0131 , \reg1_reg[28]/NET0131 , \reg1_reg[29]/NET0131 , \reg1_reg[2]/NET0131 , \reg1_reg[30]/NET0131 , \reg1_reg[31]/NET0131 , \reg1_reg[3]/NET0131 , \reg1_reg[4]/NET0131 , \reg1_reg[5]/NET0131 , \reg1_reg[6]/NET0131 , \reg1_reg[7]/NET0131 , \reg1_reg[8]/NET0131 , \reg1_reg[9]/NET0131 , \reg2_reg[0]/NET0131 , \reg2_reg[10]/NET0131 , \reg2_reg[11]/NET0131 , \reg2_reg[12]/NET0131 , \reg2_reg[13]/NET0131 , \reg2_reg[14]/NET0131 , \reg2_reg[15]/NET0131 , \reg2_reg[16]/NET0131 , \reg2_reg[17]/NET0131 , \reg2_reg[18]/NET0131 , \reg2_reg[19]/NET0131 , \reg2_reg[1]/NET0131 , \reg2_reg[20]/NET0131 , \reg2_reg[21]/NET0131 , \reg2_reg[22]/NET0131 , \reg2_reg[23]/NET0131 , \reg2_reg[24]/NET0131 , \reg2_reg[25]/NET0131 , \reg2_reg[26]/NET0131 , \reg2_reg[27]/NET0131 , \reg2_reg[28]/NET0131 , \reg2_reg[29]/NET0131 , \reg2_reg[2]/NET0131 , \reg2_reg[30]/NET0131 , \reg2_reg[31]/NET0131 , \reg2_reg[3]/NET0131 , \reg2_reg[4]/NET0131 , \reg2_reg[5]/NET0131 , \reg2_reg[6]/NET0131 , \reg2_reg[7]/NET0131 , \reg2_reg[8]/NET0131 , \reg2_reg[9]/NET0131 , \reg3_reg[0]/NET0131 , \reg3_reg[10]/NET0131 , \reg3_reg[11]/NET0131 , \reg3_reg[12]/NET0131 , \reg3_reg[13]/NET0131 , \reg3_reg[14]/NET0131 , \reg3_reg[15]/NET0131 , \reg3_reg[16]/NET0131 , \reg3_reg[17]/NET0131 , \reg3_reg[18]/NET0131 , \reg3_reg[19]/NET0131 , \reg3_reg[1]/NET0131 , \reg3_reg[20]/NET0131 , \reg3_reg[21]/NET0131 , \reg3_reg[22]/NET0131 , \reg3_reg[23]/NET0131 , \reg3_reg[24]/NET0131 , \reg3_reg[25]/NET0131 , \reg3_reg[26]/NET0131 , \reg3_reg[27]/NET0131 , \reg3_reg[28]/NET0131 , \reg3_reg[2]/NET0131 , \reg3_reg[3]/NET0131 , \reg3_reg[4]/NET0131 , \reg3_reg[5]/NET0131 , \reg3_reg[6]/NET0131 , \reg3_reg[7]/NET0131 , \reg3_reg[8]/NET0131 , \reg3_reg[9]/NET0131 , \state_reg[0]/NET0131 , \_al_n0 , \_al_n1 , \g29_dup/_0_ , \g33_dup47063/_0_ , \g36117/_0_ , \g36132/_0_ , \g36133/_0_ , \g36134/_0_ , \g36135/_0_ , \g36136/_0_ , \g36153/_0_ , \g36154/_0_ , \g36155/_0_ , \g36156/_0_ , \g36157/_0_ , \g36158/_0_ , \g36186/_0_ , \g36187/_0_ , \g36193/_0_ , \g36197/_0_ , \g36198/_0_ , \g36199/_0_ , \g36200/_0_ , \g36201/_0_ , \g36202/_0_ , \g36203/_0_ , \g36204/_0_ , \g36239/_0_ , \g36240/_0_ , \g36242/_0_ , \g36246/_0_ , \g36255/_0_ , \g36259/_0_ , \g36260/_0_ , \g36261/_0_ , \g36262/_0_ , \g36263/_0_ , \g36264/_0_ , \g36265/_0_ , \g36266/_0_ , \g36267/_0_ , \g36268/_0_ , \g36269/_0_ , \g36270/_0_ , \g36271/_0_ , \g36272/_0_ , \g36273/_0_ , \g36274/_0_ , \g36321/_0_ , \g36322/_0_ , \g36323/_0_ , \g36324/_0_ , \g36325/_0_ , \g36341/_0_ , \g36343/_0_ , \g36344/_0_ , \g36345/_0_ , \g36346/_0_ , \g36347/_0_ , \g36348/_0_ , \g36349/_0_ , \g36350/_0_ , \g36351/_0_ , \g36352/_0_ , \g36353/_0_ , \g36354/_0_ , \g36355/_0_ , \g36356/_0_ , \g36357/_0_ , \g36358/_0_ , \g36359/_0_ , \g36360/_0_ , \g36361/_0_ , \g36362/_0_ , \g36363/_0_ , \g36410/_0_ , \g36413/_0_ , \g36414/_0_ , \g36415/_0_ , \g36416/_0_ , \g36424/_0_ , \g36425/_0_ , \g36452/_0_ , \g36455/_0_ , \g36456/_0_ , \g36457/_0_ , \g36458/_0_ , \g36459/_0_ , \g36460/_0_ , \g36461/_0_ , \g36462/_0_ , \g36463/_0_ , \g36464/_0_ , \g36465/_0_ , \g36466/_0_ , \g36467/_0_ , \g36468/_0_ , \g36469/_0_ , \g36470/_0_ , \g36471/_0_ , \g36472/_0_ , \g36473/_0_ , \g36557/_0_ , \g36558/_0_ , \g36559/_0_ , \g36560/_0_ , \g36561/_0_ , \g36562/_0_ , \g36563/_0_ , \g36564/_0_ , \g36565/_0_ , \g36566/_0_ , \g36567/_0_ , \g36568/_0_ , \g36569/_0_ , \g36570/_0_ , \g36571/_0_ , \g36572/_0_ , \g36573/_0_ , \g36574/_0_ , \g36575/_0_ , \g36576/_0_ , \g36577/_0_ , \g36672/_0_ , \g36673/_0_ , \g36674/_0_ , \g38/_0_ , \g38_dup47616/_1_ , \g39789/u3_syn_4 , \g40089/_0_ , \g40090/_0_ , \g40092/_0_ , \g40093/_0_ , \g40095/_0_ , \g40096/_0_ , \g40097/_0_ , \g40098/_0_ , \g40099/_0_ , \g40100/_0_ , \g40105/_0_ , \g40106/_0_ , \g40108/_0_ , \g40109/_0_ , \g40219/_0_ , \g40220/_0_ , \g40221/_0_ , \g40222/_0_ , \g40223/_0_ , \g40228/_0_ , \g40434/_0_ , \g40495/_0_ , \g40760/_0_ , \g41149/u3_syn_4 , \g42397/_0_ , \g42487/_0_ , \g42553/_0_ , \g43089/_0_ , \g43163/_0_ , \g43169/_0_ , \g43180/_0_ , \g43189_dup/_0_ , \g43196/_0_ , \g43217/_0_ , \g43236/_0_ , \g43251/_0_ , \g43256/_0_ , \g43272/_0_ , \g43277/_0_ , \g43324/_0_ , \g43341/_0_ , \g43350/_0_ , \g43360/_0_ , \g44419/_3_ , \g44452/_3_ , \g44514/_3_ , \g44515/_3_ , \g44516/_3_ , \g44583/_3_ , \g44586/_3_ , \g44587/_3_ , \g44588/_3_ , \g44589/_3_ , \g44590/_3_ , \g44591/_3_ , \g44679/_0_ , \g44680/_3_ , \g44681/_3_ , \g44682/_3_ , \g44686/_3_ , \g44687/_3_ , \g44688/_3_ , \g44689/_3_ , \g44771/_3_ , \g44785/_3_ , \g44795/_3_ , \g44796/_3_ , \g44906/_3_ , \g44968/_3_ , \g44984/_3_ , \g45042/_3_ , \g45044/_3_ , \g45115/_3_ , \g45116/_3_ , \g46478/_1_ , \g46505/_0_ , \g46519/_0_ , \g46696/_0_ , \g47017/_2_ , \g47072_dup/_0_ , \g47395/_0_ , \g47397/_0_ , \g47401/_0_ , \g47404/_0_ , \g47458/_0_ , \g47540/_0_ , \g47791/_0_ , \state_reg[0]/NET0131_syn_2 );
	input \B_reg/NET0131  ;
	input \IR_reg[0]/NET0131  ;
	input \IR_reg[10]/NET0131  ;
	input \IR_reg[11]/NET0131  ;
	input \IR_reg[12]/NET0131  ;
	input \IR_reg[13]/NET0131  ;
	input \IR_reg[14]/NET0131  ;
	input \IR_reg[15]/NET0131  ;
	input \IR_reg[16]/NET0131  ;
	input \IR_reg[17]/NET0131  ;
	input \IR_reg[18]/NET0131  ;
	input \IR_reg[19]/NET0131  ;
	input \IR_reg[1]/NET0131  ;
	input \IR_reg[20]/NET0131  ;
	input \IR_reg[21]/NET0131  ;
	input \IR_reg[22]/NET0131  ;
	input \IR_reg[23]/NET0131  ;
	input \IR_reg[24]/NET0131  ;
	input \IR_reg[25]/NET0131  ;
	input \IR_reg[26]/NET0131  ;
	input \IR_reg[27]/NET0131  ;
	input \IR_reg[28]/NET0131  ;
	input \IR_reg[29]/NET0131  ;
	input \IR_reg[2]/NET0131  ;
	input \IR_reg[30]/NET0131  ;
	input \IR_reg[31]/NET0131  ;
	input \IR_reg[3]/NET0131  ;
	input \IR_reg[4]/NET0131  ;
	input \IR_reg[5]/NET0131  ;
	input \IR_reg[6]/NET0131  ;
	input \IR_reg[7]/NET0131  ;
	input \IR_reg[8]/NET0131  ;
	input \IR_reg[9]/NET0131  ;
	input \addr[0]_pad  ;
	input \addr[10]_pad  ;
	input \addr[11]_pad  ;
	input \addr[12]_pad  ;
	input \addr[13]_pad  ;
	input \addr[14]_pad  ;
	input \addr[15]_pad  ;
	input \addr[16]_pad  ;
	input \addr[17]_pad  ;
	input \addr[18]_pad  ;
	input \addr[19]_pad  ;
	input \addr[1]_pad  ;
	input \addr[2]_pad  ;
	input \addr[3]_pad  ;
	input \addr[4]_pad  ;
	input \addr[5]_pad  ;
	input \addr[6]_pad  ;
	input \addr[7]_pad  ;
	input \addr[8]_pad  ;
	input \addr[9]_pad  ;
	input \d_reg[0]/NET0131  ;
	input \d_reg[1]/NET0131  ;
	input \datai[0]_pad  ;
	input \datai[10]_pad  ;
	input \datai[11]_pad  ;
	input \datai[12]_pad  ;
	input \datai[13]_pad  ;
	input \datai[14]_pad  ;
	input \datai[15]_pad  ;
	input \datai[16]_pad  ;
	input \datai[17]_pad  ;
	input \datai[18]_pad  ;
	input \datai[19]_pad  ;
	input \datai[1]_pad  ;
	input \datai[20]_pad  ;
	input \datai[21]_pad  ;
	input \datai[22]_pad  ;
	input \datai[23]_pad  ;
	input \datai[24]_pad  ;
	input \datai[25]_pad  ;
	input \datai[26]_pad  ;
	input \datai[27]_pad  ;
	input \datai[28]_pad  ;
	input \datai[29]_pad  ;
	input \datai[2]_pad  ;
	input \datai[30]_pad  ;
	input \datai[31]_pad  ;
	input \datai[3]_pad  ;
	input \datai[4]_pad  ;
	input \datai[5]_pad  ;
	input \datai[6]_pad  ;
	input \datai[7]_pad  ;
	input \datai[8]_pad  ;
	input \datai[9]_pad  ;
	input \reg0_reg[0]/NET0131  ;
	input \reg0_reg[10]/NET0131  ;
	input \reg0_reg[11]/NET0131  ;
	input \reg0_reg[12]/NET0131  ;
	input \reg0_reg[13]/NET0131  ;
	input \reg0_reg[14]/NET0131  ;
	input \reg0_reg[15]/NET0131  ;
	input \reg0_reg[16]/NET0131  ;
	input \reg0_reg[17]/NET0131  ;
	input \reg0_reg[18]/NET0131  ;
	input \reg0_reg[19]/NET0131  ;
	input \reg0_reg[1]/NET0131  ;
	input \reg0_reg[20]/NET0131  ;
	input \reg0_reg[21]/NET0131  ;
	input \reg0_reg[22]/NET0131  ;
	input \reg0_reg[23]/NET0131  ;
	input \reg0_reg[24]/NET0131  ;
	input \reg0_reg[25]/NET0131  ;
	input \reg0_reg[26]/NET0131  ;
	input \reg0_reg[27]/NET0131  ;
	input \reg0_reg[28]/NET0131  ;
	input \reg0_reg[29]/NET0131  ;
	input \reg0_reg[2]/NET0131  ;
	input \reg0_reg[30]/NET0131  ;
	input \reg0_reg[31]/NET0131  ;
	input \reg0_reg[3]/NET0131  ;
	input \reg0_reg[4]/NET0131  ;
	input \reg0_reg[5]/NET0131  ;
	input \reg0_reg[6]/NET0131  ;
	input \reg0_reg[7]/NET0131  ;
	input \reg0_reg[8]/NET0131  ;
	input \reg0_reg[9]/NET0131  ;
	input \reg1_reg[0]/NET0131  ;
	input \reg1_reg[10]/NET0131  ;
	input \reg1_reg[11]/NET0131  ;
	input \reg1_reg[12]/NET0131  ;
	input \reg1_reg[13]/NET0131  ;
	input \reg1_reg[14]/NET0131  ;
	input \reg1_reg[15]/NET0131  ;
	input \reg1_reg[16]/NET0131  ;
	input \reg1_reg[17]/NET0131  ;
	input \reg1_reg[18]/NET0131  ;
	input \reg1_reg[19]/NET0131  ;
	input \reg1_reg[1]/NET0131  ;
	input \reg1_reg[20]/NET0131  ;
	input \reg1_reg[21]/NET0131  ;
	input \reg1_reg[22]/NET0131  ;
	input \reg1_reg[23]/NET0131  ;
	input \reg1_reg[24]/NET0131  ;
	input \reg1_reg[25]/NET0131  ;
	input \reg1_reg[26]/NET0131  ;
	input \reg1_reg[27]/NET0131  ;
	input \reg1_reg[28]/NET0131  ;
	input \reg1_reg[29]/NET0131  ;
	input \reg1_reg[2]/NET0131  ;
	input \reg1_reg[30]/NET0131  ;
	input \reg1_reg[31]/NET0131  ;
	input \reg1_reg[3]/NET0131  ;
	input \reg1_reg[4]/NET0131  ;
	input \reg1_reg[5]/NET0131  ;
	input \reg1_reg[6]/NET0131  ;
	input \reg1_reg[7]/NET0131  ;
	input \reg1_reg[8]/NET0131  ;
	input \reg1_reg[9]/NET0131  ;
	input \reg2_reg[0]/NET0131  ;
	input \reg2_reg[10]/NET0131  ;
	input \reg2_reg[11]/NET0131  ;
	input \reg2_reg[12]/NET0131  ;
	input \reg2_reg[13]/NET0131  ;
	input \reg2_reg[14]/NET0131  ;
	input \reg2_reg[15]/NET0131  ;
	input \reg2_reg[16]/NET0131  ;
	input \reg2_reg[17]/NET0131  ;
	input \reg2_reg[18]/NET0131  ;
	input \reg2_reg[19]/NET0131  ;
	input \reg2_reg[1]/NET0131  ;
	input \reg2_reg[20]/NET0131  ;
	input \reg2_reg[21]/NET0131  ;
	input \reg2_reg[22]/NET0131  ;
	input \reg2_reg[23]/NET0131  ;
	input \reg2_reg[24]/NET0131  ;
	input \reg2_reg[25]/NET0131  ;
	input \reg2_reg[26]/NET0131  ;
	input \reg2_reg[27]/NET0131  ;
	input \reg2_reg[28]/NET0131  ;
	input \reg2_reg[29]/NET0131  ;
	input \reg2_reg[2]/NET0131  ;
	input \reg2_reg[30]/NET0131  ;
	input \reg2_reg[31]/NET0131  ;
	input \reg2_reg[3]/NET0131  ;
	input \reg2_reg[4]/NET0131  ;
	input \reg2_reg[5]/NET0131  ;
	input \reg2_reg[6]/NET0131  ;
	input \reg2_reg[7]/NET0131  ;
	input \reg2_reg[8]/NET0131  ;
	input \reg2_reg[9]/NET0131  ;
	input \reg3_reg[0]/NET0131  ;
	input \reg3_reg[10]/NET0131  ;
	input \reg3_reg[11]/NET0131  ;
	input \reg3_reg[12]/NET0131  ;
	input \reg3_reg[13]/NET0131  ;
	input \reg3_reg[14]/NET0131  ;
	input \reg3_reg[15]/NET0131  ;
	input \reg3_reg[16]/NET0131  ;
	input \reg3_reg[17]/NET0131  ;
	input \reg3_reg[18]/NET0131  ;
	input \reg3_reg[19]/NET0131  ;
	input \reg3_reg[1]/NET0131  ;
	input \reg3_reg[20]/NET0131  ;
	input \reg3_reg[21]/NET0131  ;
	input \reg3_reg[22]/NET0131  ;
	input \reg3_reg[23]/NET0131  ;
	input \reg3_reg[24]/NET0131  ;
	input \reg3_reg[25]/NET0131  ;
	input \reg3_reg[26]/NET0131  ;
	input \reg3_reg[27]/NET0131  ;
	input \reg3_reg[28]/NET0131  ;
	input \reg3_reg[2]/NET0131  ;
	input \reg3_reg[3]/NET0131  ;
	input \reg3_reg[4]/NET0131  ;
	input \reg3_reg[5]/NET0131  ;
	input \reg3_reg[6]/NET0131  ;
	input \reg3_reg[7]/NET0131  ;
	input \reg3_reg[8]/NET0131  ;
	input \reg3_reg[9]/NET0131  ;
	input \state_reg[0]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g29_dup/_0_  ;
	output \g33_dup47063/_0_  ;
	output \g36117/_0_  ;
	output \g36132/_0_  ;
	output \g36133/_0_  ;
	output \g36134/_0_  ;
	output \g36135/_0_  ;
	output \g36136/_0_  ;
	output \g36153/_0_  ;
	output \g36154/_0_  ;
	output \g36155/_0_  ;
	output \g36156/_0_  ;
	output \g36157/_0_  ;
	output \g36158/_0_  ;
	output \g36186/_0_  ;
	output \g36187/_0_  ;
	output \g36193/_0_  ;
	output \g36197/_0_  ;
	output \g36198/_0_  ;
	output \g36199/_0_  ;
	output \g36200/_0_  ;
	output \g36201/_0_  ;
	output \g36202/_0_  ;
	output \g36203/_0_  ;
	output \g36204/_0_  ;
	output \g36239/_0_  ;
	output \g36240/_0_  ;
	output \g36242/_0_  ;
	output \g36246/_0_  ;
	output \g36255/_0_  ;
	output \g36259/_0_  ;
	output \g36260/_0_  ;
	output \g36261/_0_  ;
	output \g36262/_0_  ;
	output \g36263/_0_  ;
	output \g36264/_0_  ;
	output \g36265/_0_  ;
	output \g36266/_0_  ;
	output \g36267/_0_  ;
	output \g36268/_0_  ;
	output \g36269/_0_  ;
	output \g36270/_0_  ;
	output \g36271/_0_  ;
	output \g36272/_0_  ;
	output \g36273/_0_  ;
	output \g36274/_0_  ;
	output \g36321/_0_  ;
	output \g36322/_0_  ;
	output \g36323/_0_  ;
	output \g36324/_0_  ;
	output \g36325/_0_  ;
	output \g36341/_0_  ;
	output \g36343/_0_  ;
	output \g36344/_0_  ;
	output \g36345/_0_  ;
	output \g36346/_0_  ;
	output \g36347/_0_  ;
	output \g36348/_0_  ;
	output \g36349/_0_  ;
	output \g36350/_0_  ;
	output \g36351/_0_  ;
	output \g36352/_0_  ;
	output \g36353/_0_  ;
	output \g36354/_0_  ;
	output \g36355/_0_  ;
	output \g36356/_0_  ;
	output \g36357/_0_  ;
	output \g36358/_0_  ;
	output \g36359/_0_  ;
	output \g36360/_0_  ;
	output \g36361/_0_  ;
	output \g36362/_0_  ;
	output \g36363/_0_  ;
	output \g36410/_0_  ;
	output \g36413/_0_  ;
	output \g36414/_0_  ;
	output \g36415/_0_  ;
	output \g36416/_0_  ;
	output \g36424/_0_  ;
	output \g36425/_0_  ;
	output \g36452/_0_  ;
	output \g36455/_0_  ;
	output \g36456/_0_  ;
	output \g36457/_0_  ;
	output \g36458/_0_  ;
	output \g36459/_0_  ;
	output \g36460/_0_  ;
	output \g36461/_0_  ;
	output \g36462/_0_  ;
	output \g36463/_0_  ;
	output \g36464/_0_  ;
	output \g36465/_0_  ;
	output \g36466/_0_  ;
	output \g36467/_0_  ;
	output \g36468/_0_  ;
	output \g36469/_0_  ;
	output \g36470/_0_  ;
	output \g36471/_0_  ;
	output \g36472/_0_  ;
	output \g36473/_0_  ;
	output \g36557/_0_  ;
	output \g36558/_0_  ;
	output \g36559/_0_  ;
	output \g36560/_0_  ;
	output \g36561/_0_  ;
	output \g36562/_0_  ;
	output \g36563/_0_  ;
	output \g36564/_0_  ;
	output \g36565/_0_  ;
	output \g36566/_0_  ;
	output \g36567/_0_  ;
	output \g36568/_0_  ;
	output \g36569/_0_  ;
	output \g36570/_0_  ;
	output \g36571/_0_  ;
	output \g36572/_0_  ;
	output \g36573/_0_  ;
	output \g36574/_0_  ;
	output \g36575/_0_  ;
	output \g36576/_0_  ;
	output \g36577/_0_  ;
	output \g36672/_0_  ;
	output \g36673/_0_  ;
	output \g36674/_0_  ;
	output \g38/_0_  ;
	output \g38_dup47616/_1_  ;
	output \g39789/u3_syn_4  ;
	output \g40089/_0_  ;
	output \g40090/_0_  ;
	output \g40092/_0_  ;
	output \g40093/_0_  ;
	output \g40095/_0_  ;
	output \g40096/_0_  ;
	output \g40097/_0_  ;
	output \g40098/_0_  ;
	output \g40099/_0_  ;
	output \g40100/_0_  ;
	output \g40105/_0_  ;
	output \g40106/_0_  ;
	output \g40108/_0_  ;
	output \g40109/_0_  ;
	output \g40219/_0_  ;
	output \g40220/_0_  ;
	output \g40221/_0_  ;
	output \g40222/_0_  ;
	output \g40223/_0_  ;
	output \g40228/_0_  ;
	output \g40434/_0_  ;
	output \g40495/_0_  ;
	output \g40760/_0_  ;
	output \g41149/u3_syn_4  ;
	output \g42397/_0_  ;
	output \g42487/_0_  ;
	output \g42553/_0_  ;
	output \g43089/_0_  ;
	output \g43163/_0_  ;
	output \g43169/_0_  ;
	output \g43180/_0_  ;
	output \g43189_dup/_0_  ;
	output \g43196/_0_  ;
	output \g43217/_0_  ;
	output \g43236/_0_  ;
	output \g43251/_0_  ;
	output \g43256/_0_  ;
	output \g43272/_0_  ;
	output \g43277/_0_  ;
	output \g43324/_0_  ;
	output \g43341/_0_  ;
	output \g43350/_0_  ;
	output \g43360/_0_  ;
	output \g44419/_3_  ;
	output \g44452/_3_  ;
	output \g44514/_3_  ;
	output \g44515/_3_  ;
	output \g44516/_3_  ;
	output \g44583/_3_  ;
	output \g44586/_3_  ;
	output \g44587/_3_  ;
	output \g44588/_3_  ;
	output \g44589/_3_  ;
	output \g44590/_3_  ;
	output \g44591/_3_  ;
	output \g44679/_0_  ;
	output \g44680/_3_  ;
	output \g44681/_3_  ;
	output \g44682/_3_  ;
	output \g44686/_3_  ;
	output \g44687/_3_  ;
	output \g44688/_3_  ;
	output \g44689/_3_  ;
	output \g44771/_3_  ;
	output \g44785/_3_  ;
	output \g44795/_3_  ;
	output \g44796/_3_  ;
	output \g44906/_3_  ;
	output \g44968/_3_  ;
	output \g44984/_3_  ;
	output \g45042/_3_  ;
	output \g45044/_3_  ;
	output \g45115/_3_  ;
	output \g45116/_3_  ;
	output \g46478/_1_  ;
	output \g46505/_0_  ;
	output \g46519/_0_  ;
	output \g46696/_0_  ;
	output \g47017/_2_  ;
	output \g47072_dup/_0_  ;
	output \g47395/_0_  ;
	output \g47397/_0_  ;
	output \g47401/_0_  ;
	output \g47404/_0_  ;
	output \g47458/_0_  ;
	output \g47540/_0_  ;
	output \g47791/_0_  ;
	output \state_reg[0]/NET0131_syn_2  ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\state_reg[0]/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\IR_reg[6]/NET0131 ,
		\IR_reg[7]/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('h0001)
	) name2 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[3]/NET0131 ,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\IR_reg[4]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		_w218_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		_w216_,
		_w217_,
		_w218_,
		_w219_
	);
	LUT3 #(
		.INIT('h01)
	) name5 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[8]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w220_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[12]/NET0131 ,
		\IR_reg[13]/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w220_,
		_w221_,
		_w222_
	);
	LUT3 #(
		.INIT('h2a)
	) name8 (
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		_w224_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[18]/NET0131 ,
		\IR_reg[19]/NET0131 ,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT3 #(
		.INIT('h01)
	) name12 (
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		\IR_reg[23]/NET0131 ,
		_w227_
	);
	LUT4 #(
		.INIT('h0001)
	) name13 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		\IR_reg[23]/NET0131 ,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		_w229_
	);
	LUT4 #(
		.INIT('h8000)
	) name15 (
		_w224_,
		_w225_,
		_w228_,
		_w229_,
		_w230_
	);
	LUT3 #(
		.INIT('h01)
	) name16 (
		\IR_reg[27]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		\IR_reg[29]/NET0131 ,
		_w231_
	);
	LUT4 #(
		.INIT('h0001)
	) name17 (
		\IR_reg[26]/NET0131 ,
		\IR_reg[27]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		\IR_reg[29]/NET0131 ,
		_w232_
	);
	LUT3 #(
		.INIT('h2a)
	) name18 (
		\IR_reg[31]/NET0131 ,
		_w230_,
		_w232_,
		_w233_
	);
	LUT3 #(
		.INIT('h56)
	) name19 (
		\IR_reg[30]/NET0131 ,
		_w223_,
		_w233_,
		_w234_
	);
	LUT3 #(
		.INIT('h01)
	) name20 (
		\IR_reg[6]/NET0131 ,
		\IR_reg[7]/NET0131 ,
		\IR_reg[8]/NET0131 ,
		_w235_
	);
	LUT4 #(
		.INIT('h0001)
	) name21 (
		\IR_reg[10]/NET0131 ,
		\IR_reg[11]/NET0131 ,
		\IR_reg[12]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w236_
	);
	LUT4 #(
		.INIT('h8000)
	) name22 (
		_w217_,
		_w218_,
		_w235_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		\IR_reg[20]/NET0131 ,
		_w238_
	);
	LUT3 #(
		.INIT('h01)
	) name24 (
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		_w239_
	);
	LUT4 #(
		.INIT('h0001)
	) name25 (
		\IR_reg[24]/NET0131 ,
		\IR_reg[25]/NET0131 ,
		\IR_reg[26]/NET0131 ,
		\IR_reg[27]/NET0131 ,
		_w240_
	);
	LUT4 #(
		.INIT('h0001)
	) name26 (
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		\IR_reg[23]/NET0131 ,
		\IR_reg[28]/NET0131 ,
		_w241_
	);
	LUT4 #(
		.INIT('h8000)
	) name27 (
		_w225_,
		_w238_,
		_w240_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('ha666)
	) name28 (
		\IR_reg[29]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w237_,
		_w242_,
		_w243_
	);
	LUT4 #(
		.INIT('h0056)
	) name29 (
		\IR_reg[30]/NET0131 ,
		_w223_,
		_w233_,
		_w243_,
		_w244_
	);
	LUT4 #(
		.INIT('ha900)
	) name30 (
		\IR_reg[30]/NET0131 ,
		_w223_,
		_w233_,
		_w243_,
		_w245_
	);
	LUT4 #(
		.INIT('hf53f)
	) name31 (
		\reg1_reg[5]/NET0131 ,
		\reg2_reg[5]/NET0131 ,
		_w234_,
		_w243_,
		_w246_
	);
	LUT4 #(
		.INIT('h5600)
	) name32 (
		\IR_reg[30]/NET0131 ,
		_w223_,
		_w233_,
		_w243_,
		_w247_
	);
	LUT3 #(
		.INIT('h78)
	) name33 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		_w248_
	);
	LUT4 #(
		.INIT('h00a9)
	) name34 (
		\IR_reg[30]/NET0131 ,
		_w223_,
		_w233_,
		_w243_,
		_w249_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name35 (
		\reg0_reg[5]/NET0131 ,
		_w234_,
		_w243_,
		_w248_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w246_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h7)
	) name37 (
		_w246_,
		_w250_,
		_w252_
	);
	LUT4 #(
		.INIT('h8000)
	) name38 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		\reg3_reg[6]/NET0131 ,
		_w253_
	);
	LUT4 #(
		.INIT('h8000)
	) name39 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		\reg3_reg[9]/NET0131 ,
		_w253_,
		_w254_
	);
	LUT3 #(
		.INIT('h80)
	) name40 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h8000)
	) name41 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		\reg3_reg[12]/NET0131 ,
		_w254_,
		_w256_
	);
	LUT2 #(
		.INIT('h6)
	) name42 (
		\reg3_reg[13]/NET0131 ,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name43 (
		\reg0_reg[13]/NET0131 ,
		_w234_,
		_w243_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('hf53f)
	) name44 (
		\reg1_reg[13]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w234_,
		_w243_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w258_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h7)
	) name46 (
		_w258_,
		_w259_,
		_w261_
	);
	LUT3 #(
		.INIT('h40)
	) name47 (
		\IR_reg[14]/NET0131 ,
		_w220_,
		_w221_,
		_w262_
	);
	LUT4 #(
		.INIT('h0001)
	) name48 (
		\IR_reg[15]/NET0131 ,
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[18]/NET0131 ,
		_w263_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name49 (
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w262_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\IR_reg[19]/NET0131 ,
		\IR_reg[20]/NET0131 ,
		_w265_
	);
	LUT4 #(
		.INIT('h0001)
	) name51 (
		\IR_reg[19]/NET0131 ,
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\IR_reg[31]/NET0131 ,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h56)
	) name53 (
		\IR_reg[23]/NET0131 ,
		_w264_,
		_w267_,
		_w268_
	);
	LUT4 #(
		.INIT('h4448)
	) name54 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w264_,
		_w267_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\B_reg/NET0131 ,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name56 (
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w222_,
		_w226_,
		_w271_
	);
	LUT2 #(
		.INIT('h9)
	) name57 (
		\IR_reg[20]/NET0131 ,
		_w271_,
		_w272_
	);
	LUT3 #(
		.INIT('h80)
	) name58 (
		_w227_,
		_w239_,
		_w265_,
		_w273_
	);
	LUT4 #(
		.INIT('h8000)
	) name59 (
		_w219_,
		_w262_,
		_w263_,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('ha6)
	) name60 (
		\IR_reg[27]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w274_,
		_w275_
	);
	LUT3 #(
		.INIT('h2a)
	) name61 (
		\IR_reg[31]/NET0131 ,
		_w228_,
		_w240_,
		_w276_
	);
	LUT3 #(
		.INIT('h56)
	) name62 (
		\IR_reg[28]/NET0131 ,
		_w271_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w275_,
		_w277_,
		_w278_
	);
	LUT3 #(
		.INIT('ha8)
	) name64 (
		\datai[31]_pad ,
		_w275_,
		_w277_,
		_w279_
	);
	LUT3 #(
		.INIT('h80)
	) name65 (
		\reg3_reg[12]/NET0131 ,
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		_w280_
	);
	LUT4 #(
		.INIT('h8000)
	) name66 (
		\reg3_reg[12]/NET0131 ,
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		\reg3_reg[15]/NET0131 ,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\reg3_reg[16]/NET0131 ,
		_w281_,
		_w282_
	);
	LUT4 #(
		.INIT('h8000)
	) name68 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		_w254_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w284_
	);
	LUT3 #(
		.INIT('h80)
	) name70 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		\reg3_reg[22]/NET0131 ,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\reg3_reg[17]/NET0131 ,
		\reg3_reg[18]/NET0131 ,
		_w286_
	);
	LUT3 #(
		.INIT('h80)
	) name72 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[23]/NET0131 ,
		\reg3_reg[24]/NET0131 ,
		_w287_
	);
	LUT3 #(
		.INIT('h80)
	) name73 (
		_w285_,
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w283_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		\reg3_reg[27]/NET0131 ,
		\reg3_reg[28]/NET0131 ,
		_w290_
	);
	LUT3 #(
		.INIT('h80)
	) name76 (
		_w283_,
		_w288_,
		_w290_,
		_w291_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name77 (
		\reg0_reg[31]/NET0131 ,
		_w234_,
		_w243_,
		_w291_,
		_w292_
	);
	LUT4 #(
		.INIT('hf53f)
	) name78 (
		\reg1_reg[31]/NET0131 ,
		\reg2_reg[31]/NET0131 ,
		_w234_,
		_w243_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h7)
	) name80 (
		_w292_,
		_w293_,
		_w295_
	);
	LUT3 #(
		.INIT('ha8)
	) name81 (
		\datai[30]_pad ,
		_w275_,
		_w277_,
		_w296_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name82 (
		\reg0_reg[30]/NET0131 ,
		_w234_,
		_w243_,
		_w291_,
		_w297_
	);
	LUT4 #(
		.INIT('hf53f)
	) name83 (
		\reg1_reg[30]/NET0131 ,
		\reg2_reg[30]/NET0131 ,
		_w234_,
		_w243_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h7)
	) name85 (
		_w297_,
		_w298_,
		_w300_
	);
	LUT3 #(
		.INIT('h15)
	) name86 (
		_w296_,
		_w297_,
		_w298_,
		_w301_
	);
	LUT3 #(
		.INIT('ha8)
	) name87 (
		_w279_,
		_w294_,
		_w301_,
		_w302_
	);
	LUT3 #(
		.INIT('ha8)
	) name88 (
		\datai[29]_pad ,
		_w275_,
		_w277_,
		_w303_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name89 (
		\reg1_reg[29]/NET0131 ,
		_w234_,
		_w243_,
		_w291_,
		_w304_
	);
	LUT4 #(
		.INIT('hff35)
	) name90 (
		\reg0_reg[29]/NET0131 ,
		\reg2_reg[29]/NET0131 ,
		_w234_,
		_w243_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w304_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h7)
	) name92 (
		_w304_,
		_w305_,
		_w307_
	);
	LUT3 #(
		.INIT('h15)
	) name93 (
		_w303_,
		_w304_,
		_w305_,
		_w308_
	);
	LUT3 #(
		.INIT('h80)
	) name94 (
		_w303_,
		_w304_,
		_w305_,
		_w309_
	);
	LUT3 #(
		.INIT('ha8)
	) name95 (
		\datai[28]_pad ,
		_w275_,
		_w277_,
		_w310_
	);
	LUT4 #(
		.INIT('h8000)
	) name96 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		_w283_,
		_w288_,
		_w311_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name97 (
		\reg3_reg[27]/NET0131 ,
		\reg3_reg[28]/NET0131 ,
		_w291_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\reg2_reg[28]/NET0131 ,
		_w244_,
		_w313_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name99 (
		\reg0_reg[28]/NET0131 ,
		\reg1_reg[28]/NET0131 ,
		_w234_,
		_w243_,
		_w314_
	);
	LUT4 #(
		.INIT('h1300)
	) name100 (
		_w247_,
		_w313_,
		_w312_,
		_w314_,
		_w315_
	);
	LUT4 #(
		.INIT('hecff)
	) name101 (
		_w247_,
		_w313_,
		_w312_,
		_w314_,
		_w316_
	);
	LUT4 #(
		.INIT('h5554)
	) name102 (
		_w308_,
		_w309_,
		_w310_,
		_w315_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w310_,
		_w315_,
		_w318_
	);
	LUT3 #(
		.INIT('h15)
	) name104 (
		_w309_,
		_w310_,
		_w315_,
		_w319_
	);
	LUT3 #(
		.INIT('ha8)
	) name105 (
		\datai[27]_pad ,
		_w275_,
		_w277_,
		_w320_
	);
	LUT2 #(
		.INIT('h6)
	) name106 (
		\reg3_reg[27]/NET0131 ,
		_w311_,
		_w321_
	);
	LUT3 #(
		.INIT('h48)
	) name107 (
		\reg3_reg[27]/NET0131 ,
		_w247_,
		_w311_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\reg0_reg[27]/NET0131 ,
		_w249_,
		_w323_
	);
	LUT4 #(
		.INIT('hf53f)
	) name109 (
		\reg1_reg[27]/NET0131 ,
		\reg2_reg[27]/NET0131 ,
		_w234_,
		_w243_,
		_w324_
	);
	LUT3 #(
		.INIT('h10)
	) name110 (
		_w323_,
		_w322_,
		_w324_,
		_w325_
	);
	LUT3 #(
		.INIT('hef)
	) name111 (
		_w323_,
		_w322_,
		_w324_,
		_w326_
	);
	LUT4 #(
		.INIT('h0200)
	) name112 (
		_w320_,
		_w323_,
		_w322_,
		_w324_,
		_w327_
	);
	LUT3 #(
		.INIT('ha8)
	) name113 (
		\datai[26]_pad ,
		_w275_,
		_w277_,
		_w328_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name114 (
		\reg3_reg[25]/NET0131 ,
		\reg3_reg[26]/NET0131 ,
		_w283_,
		_w288_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w247_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\reg1_reg[26]/NET0131 ,
		_w245_,
		_w331_
	);
	LUT4 #(
		.INIT('hff35)
	) name117 (
		\reg0_reg[26]/NET0131 ,
		\reg2_reg[26]/NET0131 ,
		_w234_,
		_w243_,
		_w332_
	);
	LUT3 #(
		.INIT('h10)
	) name118 (
		_w331_,
		_w330_,
		_w332_,
		_w333_
	);
	LUT3 #(
		.INIT('hef)
	) name119 (
		_w331_,
		_w330_,
		_w332_,
		_w334_
	);
	LUT4 #(
		.INIT('h0200)
	) name120 (
		_w328_,
		_w331_,
		_w330_,
		_w332_,
		_w335_
	);
	LUT3 #(
		.INIT('ha8)
	) name121 (
		\datai[25]_pad ,
		_w275_,
		_w277_,
		_w336_
	);
	LUT3 #(
		.INIT('h6a)
	) name122 (
		\reg3_reg[25]/NET0131 ,
		_w283_,
		_w288_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w247_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\reg2_reg[25]/NET0131 ,
		_w244_,
		_w339_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name125 (
		\reg0_reg[25]/NET0131 ,
		\reg1_reg[25]/NET0131 ,
		_w234_,
		_w243_,
		_w340_
	);
	LUT3 #(
		.INIT('h10)
	) name126 (
		_w339_,
		_w338_,
		_w340_,
		_w341_
	);
	LUT3 #(
		.INIT('hef)
	) name127 (
		_w339_,
		_w338_,
		_w340_,
		_w342_
	);
	LUT4 #(
		.INIT('h0200)
	) name128 (
		_w336_,
		_w339_,
		_w338_,
		_w340_,
		_w343_
	);
	LUT4 #(
		.INIT('h5455)
	) name129 (
		_w336_,
		_w339_,
		_w338_,
		_w340_,
		_w344_
	);
	LUT3 #(
		.INIT('ha8)
	) name130 (
		\datai[24]_pad ,
		_w275_,
		_w277_,
		_w345_
	);
	LUT3 #(
		.INIT('h80)
	) name131 (
		\reg3_reg[19]/NET0131 ,
		_w283_,
		_w286_,
		_w346_
	);
	LUT4 #(
		.INIT('h8000)
	) name132 (
		\reg3_reg[19]/NET0131 ,
		_w283_,
		_w285_,
		_w286_,
		_w347_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name133 (
		\reg3_reg[23]/NET0131 ,
		\reg3_reg[24]/NET0131 ,
		_w289_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\reg2_reg[24]/NET0131 ,
		_w244_,
		_w349_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name135 (
		\reg0_reg[24]/NET0131 ,
		\reg1_reg[24]/NET0131 ,
		_w234_,
		_w243_,
		_w350_
	);
	LUT4 #(
		.INIT('h1300)
	) name136 (
		_w247_,
		_w349_,
		_w348_,
		_w350_,
		_w351_
	);
	LUT4 #(
		.INIT('hecff)
	) name137 (
		_w247_,
		_w349_,
		_w348_,
		_w350_,
		_w352_
	);
	LUT3 #(
		.INIT('h0e)
	) name138 (
		_w345_,
		_w351_,
		_w344_,
		_w353_
	);
	LUT4 #(
		.INIT('h5501)
	) name139 (
		_w343_,
		_w345_,
		_w351_,
		_w344_,
		_w354_
	);
	LUT4 #(
		.INIT('h5455)
	) name140 (
		_w320_,
		_w323_,
		_w322_,
		_w324_,
		_w355_
	);
	LUT4 #(
		.INIT('h5455)
	) name141 (
		_w328_,
		_w331_,
		_w330_,
		_w332_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT4 #(
		.INIT('h1055)
	) name143 (
		_w327_,
		_w335_,
		_w354_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w345_,
		_w351_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w343_,
		_w335_,
		_w360_
	);
	LUT3 #(
		.INIT('h01)
	) name146 (
		_w343_,
		_w327_,
		_w335_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w359_,
		_w361_,
		_w362_
	);
	LUT3 #(
		.INIT('ha8)
	) name148 (
		\datai[22]_pad ,
		_w275_,
		_w277_,
		_w363_
	);
	LUT4 #(
		.INIT('h8000)
	) name149 (
		\reg3_reg[19]/NET0131 ,
		_w283_,
		_w284_,
		_w286_,
		_w364_
	);
	LUT3 #(
		.INIT('h32)
	) name150 (
		\reg3_reg[22]/NET0131 ,
		_w347_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('h4888)
	) name151 (
		\reg3_reg[22]/NET0131 ,
		_w247_,
		_w284_,
		_w346_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\reg0_reg[22]/NET0131 ,
		_w249_,
		_w367_
	);
	LUT4 #(
		.INIT('hf53f)
	) name153 (
		\reg1_reg[22]/NET0131 ,
		\reg2_reg[22]/NET0131 ,
		_w234_,
		_w243_,
		_w368_
	);
	LUT3 #(
		.INIT('h10)
	) name154 (
		_w367_,
		_w366_,
		_w368_,
		_w369_
	);
	LUT3 #(
		.INIT('hef)
	) name155 (
		_w367_,
		_w366_,
		_w368_,
		_w370_
	);
	LUT4 #(
		.INIT('h0200)
	) name156 (
		_w363_,
		_w367_,
		_w366_,
		_w368_,
		_w371_
	);
	LUT3 #(
		.INIT('ha8)
	) name157 (
		\datai[23]_pad ,
		_w275_,
		_w277_,
		_w372_
	);
	LUT2 #(
		.INIT('h6)
	) name158 (
		\reg3_reg[23]/NET0131 ,
		_w347_,
		_w373_
	);
	LUT3 #(
		.INIT('h48)
	) name159 (
		\reg3_reg[23]/NET0131 ,
		_w247_,
		_w347_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\reg1_reg[23]/NET0131 ,
		_w245_,
		_w375_
	);
	LUT4 #(
		.INIT('hff35)
	) name161 (
		\reg0_reg[23]/NET0131 ,
		\reg2_reg[23]/NET0131 ,
		_w234_,
		_w243_,
		_w376_
	);
	LUT3 #(
		.INIT('h10)
	) name162 (
		_w375_,
		_w374_,
		_w376_,
		_w377_
	);
	LUT3 #(
		.INIT('hef)
	) name163 (
		_w375_,
		_w374_,
		_w376_,
		_w378_
	);
	LUT4 #(
		.INIT('h0200)
	) name164 (
		_w372_,
		_w375_,
		_w374_,
		_w376_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w371_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('ha8)
	) name166 (
		\datai[21]_pad ,
		_w275_,
		_w277_,
		_w381_
	);
	LUT3 #(
		.INIT('h6c)
	) name167 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w346_,
		_w382_
	);
	LUT4 #(
		.INIT('h60c0)
	) name168 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w247_,
		_w346_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\reg2_reg[21]/NET0131 ,
		_w244_,
		_w384_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name170 (
		\reg0_reg[21]/NET0131 ,
		\reg1_reg[21]/NET0131 ,
		_w234_,
		_w243_,
		_w385_
	);
	LUT3 #(
		.INIT('h10)
	) name171 (
		_w384_,
		_w383_,
		_w385_,
		_w386_
	);
	LUT3 #(
		.INIT('hef)
	) name172 (
		_w384_,
		_w383_,
		_w385_,
		_w387_
	);
	LUT4 #(
		.INIT('h5455)
	) name173 (
		_w381_,
		_w384_,
		_w383_,
		_w385_,
		_w388_
	);
	LUT3 #(
		.INIT('ha8)
	) name174 (
		\datai[20]_pad ,
		_w275_,
		_w277_,
		_w389_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name175 (
		\reg3_reg[19]/NET0131 ,
		\reg3_reg[20]/NET0131 ,
		_w283_,
		_w286_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w247_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\reg2_reg[20]/NET0131 ,
		_w244_,
		_w392_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name178 (
		\reg0_reg[20]/NET0131 ,
		\reg1_reg[20]/NET0131 ,
		_w234_,
		_w243_,
		_w393_
	);
	LUT3 #(
		.INIT('h10)
	) name179 (
		_w392_,
		_w391_,
		_w393_,
		_w394_
	);
	LUT3 #(
		.INIT('hef)
	) name180 (
		_w392_,
		_w391_,
		_w393_,
		_w395_
	);
	LUT4 #(
		.INIT('h5455)
	) name181 (
		_w389_,
		_w392_,
		_w391_,
		_w393_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w388_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h0200)
	) name183 (
		_w381_,
		_w384_,
		_w383_,
		_w385_,
		_w398_
	);
	LUT3 #(
		.INIT('h71)
	) name184 (
		_w381_,
		_w386_,
		_w396_,
		_w399_
	);
	LUT4 #(
		.INIT('h5455)
	) name185 (
		_w372_,
		_w375_,
		_w374_,
		_w376_,
		_w400_
	);
	LUT4 #(
		.INIT('h5455)
	) name186 (
		_w363_,
		_w367_,
		_w366_,
		_w368_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w400_,
		_w401_,
		_w402_
	);
	LUT3 #(
		.INIT('h71)
	) name188 (
		_w372_,
		_w377_,
		_w401_,
		_w403_
	);
	LUT3 #(
		.INIT('h07)
	) name189 (
		_w380_,
		_w399_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h6)
	) name190 (
		\IR_reg[19]/NET0131 ,
		_w264_,
		_w405_
	);
	LUT4 #(
		.INIT('h5457)
	) name191 (
		\datai[19]_pad ,
		_w275_,
		_w277_,
		_w405_,
		_w406_
	);
	LUT3 #(
		.INIT('h6a)
	) name192 (
		\reg3_reg[19]/NET0131 ,
		_w283_,
		_w286_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w247_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\reg1_reg[19]/NET0131 ,
		_w245_,
		_w409_
	);
	LUT4 #(
		.INIT('hff35)
	) name195 (
		\reg0_reg[19]/NET0131 ,
		\reg2_reg[19]/NET0131 ,
		_w234_,
		_w243_,
		_w410_
	);
	LUT3 #(
		.INIT('h10)
	) name196 (
		_w409_,
		_w408_,
		_w410_,
		_w411_
	);
	LUT3 #(
		.INIT('hef)
	) name197 (
		_w409_,
		_w408_,
		_w410_,
		_w412_
	);
	LUT4 #(
		.INIT('h0100)
	) name198 (
		_w406_,
		_w409_,
		_w408_,
		_w410_,
		_w413_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name199 (
		\IR_reg[15]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w262_,
		_w414_
	);
	LUT3 #(
		.INIT('he0)
	) name200 (
		\IR_reg[16]/NET0131 ,
		\IR_reg[17]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w415_
	);
	LUT3 #(
		.INIT('h56)
	) name201 (
		\IR_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w416_
	);
	LUT4 #(
		.INIT('haba8)
	) name202 (
		\datai[18]_pad ,
		_w275_,
		_w277_,
		_w416_,
		_w417_
	);
	LUT3 #(
		.INIT('h6c)
	) name203 (
		\reg3_reg[17]/NET0131 ,
		\reg3_reg[18]/NET0131 ,
		_w283_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w247_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\reg2_reg[18]/NET0131 ,
		_w244_,
		_w420_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name206 (
		\reg0_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w234_,
		_w243_,
		_w421_
	);
	LUT3 #(
		.INIT('h10)
	) name207 (
		_w420_,
		_w419_,
		_w421_,
		_w422_
	);
	LUT3 #(
		.INIT('hef)
	) name208 (
		_w420_,
		_w419_,
		_w421_,
		_w423_
	);
	LUT4 #(
		.INIT('h0200)
	) name209 (
		_w417_,
		_w420_,
		_w419_,
		_w421_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w413_,
		_w424_,
		_w425_
	);
	LUT4 #(
		.INIT('hf53f)
	) name211 (
		\reg1_reg[17]/NET0131 ,
		\reg2_reg[17]/NET0131 ,
		_w234_,
		_w243_,
		_w426_
	);
	LUT2 #(
		.INIT('h6)
	) name212 (
		\reg3_reg[17]/NET0131 ,
		_w283_,
		_w427_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name213 (
		\reg0_reg[17]/NET0131 ,
		_w234_,
		_w243_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w426_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h7)
	) name215 (
		_w426_,
		_w428_,
		_w430_
	);
	LUT4 #(
		.INIT('h0001)
	) name216 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[14]/NET0131 ,
		\IR_reg[15]/NET0131 ,
		\IR_reg[16]/NET0131 ,
		_w431_
	);
	LUT4 #(
		.INIT('ha666)
	) name217 (
		\IR_reg[17]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w237_,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('haba8)
	) name218 (
		\datai[17]_pad ,
		_w275_,
		_w277_,
		_w432_,
		_w433_
	);
	LUT3 #(
		.INIT('h07)
	) name219 (
		_w426_,
		_w428_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h6)
	) name220 (
		\IR_reg[16]/NET0131 ,
		_w414_,
		_w435_
	);
	LUT4 #(
		.INIT('haba8)
	) name221 (
		\datai[16]_pad ,
		_w275_,
		_w277_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h8000)
	) name222 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		_w254_,
		_w281_,
		_w437_
	);
	LUT3 #(
		.INIT('h32)
	) name223 (
		\reg3_reg[16]/NET0131 ,
		_w283_,
		_w437_,
		_w438_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name224 (
		\reg0_reg[16]/NET0131 ,
		_w234_,
		_w243_,
		_w438_,
		_w439_
	);
	LUT4 #(
		.INIT('hf53f)
	) name225 (
		\reg1_reg[16]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w234_,
		_w243_,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h7)
	) name227 (
		_w439_,
		_w440_,
		_w442_
	);
	LUT3 #(
		.INIT('h15)
	) name228 (
		_w436_,
		_w439_,
		_w440_,
		_w443_
	);
	LUT3 #(
		.INIT('h80)
	) name229 (
		_w426_,
		_w428_,
		_w433_,
		_w444_
	);
	LUT3 #(
		.INIT('h71)
	) name230 (
		_w429_,
		_w433_,
		_w443_,
		_w445_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name231 (
		_w406_,
		_w409_,
		_w408_,
		_w410_,
		_w446_
	);
	LUT4 #(
		.INIT('h5455)
	) name232 (
		_w417_,
		_w420_,
		_w419_,
		_w421_,
		_w447_
	);
	LUT3 #(
		.INIT('hb2)
	) name233 (
		_w406_,
		_w411_,
		_w447_,
		_w448_
	);
	LUT3 #(
		.INIT('h07)
	) name234 (
		_w425_,
		_w445_,
		_w448_,
		_w449_
	);
	LUT4 #(
		.INIT('h0200)
	) name235 (
		_w389_,
		_w392_,
		_w391_,
		_w393_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w398_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('h0001)
	) name237 (
		_w371_,
		_w379_,
		_w398_,
		_w450_,
		_w452_
	);
	LUT4 #(
		.INIT('hf800)
	) name238 (
		_w425_,
		_w445_,
		_w448_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w404_,
		_w453_,
		_w454_
	);
	LUT4 #(
		.INIT('h78f0)
	) name240 (
		\reg3_reg[12]/NET0131 ,
		\reg3_reg[13]/NET0131 ,
		\reg3_reg[14]/NET0131 ,
		_w255_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w247_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		\reg1_reg[14]/NET0131 ,
		_w245_,
		_w457_
	);
	LUT4 #(
		.INIT('hff35)
	) name243 (
		\reg0_reg[14]/NET0131 ,
		\reg2_reg[14]/NET0131 ,
		_w234_,
		_w243_,
		_w458_
	);
	LUT3 #(
		.INIT('h10)
	) name244 (
		_w456_,
		_w457_,
		_w458_,
		_w459_
	);
	LUT3 #(
		.INIT('hef)
	) name245 (
		_w456_,
		_w457_,
		_w458_,
		_w460_
	);
	LUT4 #(
		.INIT('ha666)
	) name246 (
		\IR_reg[14]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w222_,
		_w461_
	);
	LUT4 #(
		.INIT('h5457)
	) name247 (
		\datai[14]_pad ,
		_w275_,
		_w277_,
		_w461_,
		_w462_
	);
	LUT4 #(
		.INIT('h0010)
	) name248 (
		_w456_,
		_w457_,
		_w458_,
		_w462_,
		_w463_
	);
	LUT3 #(
		.INIT('h6a)
	) name249 (
		\reg3_reg[15]/NET0131 ,
		_w255_,
		_w280_,
		_w464_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name250 (
		\reg0_reg[15]/NET0131 ,
		_w234_,
		_w243_,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('hf53f)
	) name251 (
		\reg1_reg[15]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		_w234_,
		_w243_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h7)
	) name253 (
		_w465_,
		_w466_,
		_w468_
	);
	LUT4 #(
		.INIT('ha666)
	) name254 (
		\IR_reg[15]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w262_,
		_w469_
	);
	LUT4 #(
		.INIT('haba8)
	) name255 (
		\datai[15]_pad ,
		_w275_,
		_w277_,
		_w469_,
		_w470_
	);
	LUT3 #(
		.INIT('h80)
	) name256 (
		_w465_,
		_w466_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w463_,
		_w471_,
		_w472_
	);
	LUT3 #(
		.INIT('ha6)
	) name258 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w237_,
		_w473_
	);
	LUT4 #(
		.INIT('h5457)
	) name259 (
		\datai[13]_pad ,
		_w275_,
		_w277_,
		_w473_,
		_w474_
	);
	LUT3 #(
		.INIT('h08)
	) name260 (
		_w258_,
		_w259_,
		_w474_,
		_w475_
	);
	LUT3 #(
		.INIT('h70)
	) name261 (
		_w258_,
		_w259_,
		_w474_,
		_w476_
	);
	LUT4 #(
		.INIT('hff35)
	) name262 (
		\reg0_reg[12]/NET0131 ,
		\reg2_reg[12]/NET0131 ,
		_w234_,
		_w243_,
		_w477_
	);
	LUT4 #(
		.INIT('h78f0)
	) name263 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		\reg3_reg[12]/NET0131 ,
		_w254_,
		_w478_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name264 (
		\reg1_reg[12]/NET0131 ,
		_w234_,
		_w243_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		_w477_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h7)
	) name266 (
		_w477_,
		_w479_,
		_w481_
	);
	LUT4 #(
		.INIT('h8000)
	) name267 (
		_w216_,
		_w217_,
		_w218_,
		_w220_,
		_w482_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name268 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[12]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w482_,
		_w483_
	);
	LUT4 #(
		.INIT('haba8)
	) name269 (
		\datai[12]_pad ,
		_w275_,
		_w277_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h07)
	) name270 (
		_w477_,
		_w479_,
		_w484_,
		_w485_
	);
	LUT3 #(
		.INIT('h54)
	) name271 (
		_w475_,
		_w476_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('hef00)
	) name272 (
		_w456_,
		_w457_,
		_w458_,
		_w462_,
		_w487_
	);
	LUT3 #(
		.INIT('h07)
	) name273 (
		_w465_,
		_w466_,
		_w470_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('h54)
	) name275 (
		_w471_,
		_w487_,
		_w488_,
		_w490_
	);
	LUT3 #(
		.INIT('h07)
	) name276 (
		_w472_,
		_w486_,
		_w490_,
		_w491_
	);
	LUT3 #(
		.INIT('h59)
	) name277 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w482_,
		_w492_
	);
	LUT4 #(
		.INIT('h5754)
	) name278 (
		\datai[11]_pad ,
		_w275_,
		_w277_,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h6c)
	) name279 (
		\reg3_reg[10]/NET0131 ,
		\reg3_reg[11]/NET0131 ,
		_w254_,
		_w494_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name280 (
		\reg1_reg[11]/NET0131 ,
		_w234_,
		_w243_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('hff35)
	) name281 (
		\reg0_reg[11]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w234_,
		_w243_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h7)
	) name283 (
		_w495_,
		_w496_,
		_w498_
	);
	LUT3 #(
		.INIT('h40)
	) name284 (
		_w493_,
		_w495_,
		_w496_,
		_w499_
	);
	LUT2 #(
		.INIT('h6)
	) name285 (
		\reg3_reg[10]/NET0131 ,
		_w254_,
		_w500_
	);
	LUT4 #(
		.INIT('h37f7)
	) name286 (
		\reg2_reg[10]/NET0131 ,
		_w234_,
		_w243_,
		_w500_,
		_w501_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name287 (
		\reg0_reg[10]/NET0131 ,
		\reg1_reg[10]/NET0131 ,
		_w234_,
		_w243_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h7)
	) name289 (
		_w501_,
		_w502_,
		_w504_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name290 (
		\IR_reg[31]/NET0131 ,
		_w217_,
		_w218_,
		_w235_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[9]/NET0131 ,
		_w506_
	);
	LUT3 #(
		.INIT('h56)
	) name292 (
		\IR_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w507_
	);
	LUT4 #(
		.INIT('haba8)
	) name293 (
		\datai[10]_pad ,
		_w275_,
		_w277_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('h80)
	) name294 (
		_w501_,
		_w502_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w499_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h9)
	) name296 (
		\IR_reg[9]/NET0131 ,
		_w505_,
		_w511_
	);
	LUT4 #(
		.INIT('h5754)
	) name297 (
		\datai[9]_pad ,
		_w275_,
		_w277_,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h78f0)
	) name298 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		\reg3_reg[9]/NET0131 ,
		_w253_,
		_w513_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name299 (
		\reg1_reg[9]/NET0131 ,
		_w234_,
		_w243_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('hff35)
	) name300 (
		\reg0_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w234_,
		_w243_,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h7)
	) name302 (
		_w514_,
		_w515_,
		_w517_
	);
	LUT3 #(
		.INIT('h2a)
	) name303 (
		_w512_,
		_w514_,
		_w515_,
		_w518_
	);
	LUT3 #(
		.INIT('h40)
	) name304 (
		_w512_,
		_w514_,
		_w515_,
		_w519_
	);
	LUT3 #(
		.INIT('h6c)
	) name305 (
		\reg3_reg[7]/NET0131 ,
		\reg3_reg[8]/NET0131 ,
		_w253_,
		_w520_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name306 (
		\reg1_reg[8]/NET0131 ,
		_w234_,
		_w243_,
		_w520_,
		_w521_
	);
	LUT4 #(
		.INIT('hff35)
	) name307 (
		\reg0_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w234_,
		_w243_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w521_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h7)
	) name309 (
		_w521_,
		_w522_,
		_w524_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name310 (
		\IR_reg[31]/NET0131 ,
		_w216_,
		_w217_,
		_w218_,
		_w525_
	);
	LUT2 #(
		.INIT('h6)
	) name311 (
		\IR_reg[8]/NET0131 ,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('haba8)
	) name312 (
		\datai[8]_pad ,
		_w275_,
		_w277_,
		_w526_,
		_w527_
	);
	LUT3 #(
		.INIT('h07)
	) name313 (
		_w521_,
		_w522_,
		_w527_,
		_w528_
	);
	LUT3 #(
		.INIT('h23)
	) name314 (
		_w519_,
		_w518_,
		_w528_,
		_w529_
	);
	LUT3 #(
		.INIT('h2a)
	) name315 (
		_w493_,
		_w495_,
		_w496_,
		_w530_
	);
	LUT3 #(
		.INIT('h07)
	) name316 (
		_w501_,
		_w502_,
		_w508_,
		_w531_
	);
	LUT3 #(
		.INIT('h32)
	) name317 (
		_w530_,
		_w499_,
		_w531_,
		_w532_
	);
	LUT3 #(
		.INIT('h0d)
	) name318 (
		_w510_,
		_w529_,
		_w532_,
		_w533_
	);
	LUT3 #(
		.INIT('h80)
	) name319 (
		_w477_,
		_w479_,
		_w484_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w475_,
		_w534_,
		_w535_
	);
	LUT4 #(
		.INIT('h0001)
	) name321 (
		_w463_,
		_w471_,
		_w475_,
		_w534_,
		_w536_
	);
	LUT4 #(
		.INIT('hf200)
	) name322 (
		_w510_,
		_w529_,
		_w532_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		_w491_,
		_w537_,
		_w538_
	);
	LUT4 #(
		.INIT('h3999)
	) name324 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[6]/NET0131 ,
		_w217_,
		_w218_,
		_w539_
	);
	LUT4 #(
		.INIT('h5754)
	) name325 (
		\datai[6]_pad ,
		_w275_,
		_w277_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('hf53f)
	) name326 (
		\reg1_reg[6]/NET0131 ,
		\reg2_reg[6]/NET0131 ,
		_w234_,
		_w243_,
		_w541_
	);
	LUT4 #(
		.INIT('h7f80)
	) name327 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		\reg3_reg[5]/NET0131 ,
		\reg3_reg[6]/NET0131 ,
		_w542_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name328 (
		\reg0_reg[6]/NET0131 ,
		_w234_,
		_w243_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w541_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h7)
	) name330 (
		_w541_,
		_w543_,
		_w545_
	);
	LUT3 #(
		.INIT('h40)
	) name331 (
		_w540_,
		_w541_,
		_w543_,
		_w546_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name332 (
		\reg0_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w234_,
		_w243_,
		_w547_
	);
	LUT2 #(
		.INIT('h6)
	) name333 (
		\reg3_reg[7]/NET0131 ,
		_w253_,
		_w548_
	);
	LUT4 #(
		.INIT('h37f7)
	) name334 (
		\reg2_reg[7]/NET0131 ,
		_w234_,
		_w243_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w547_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h7)
	) name336 (
		_w547_,
		_w549_,
		_w551_
	);
	LUT4 #(
		.INIT('h7555)
	) name337 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[6]/NET0131 ,
		_w217_,
		_w218_,
		_w552_
	);
	LUT2 #(
		.INIT('h9)
	) name338 (
		\IR_reg[7]/NET0131 ,
		_w552_,
		_w553_
	);
	LUT4 #(
		.INIT('haba8)
	) name339 (
		\datai[7]_pad ,
		_w275_,
		_w277_,
		_w553_,
		_w554_
	);
	LUT3 #(
		.INIT('h80)
	) name340 (
		_w547_,
		_w549_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w546_,
		_w555_,
		_w556_
	);
	LUT3 #(
		.INIT('h39)
	) name342 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		_w217_,
		_w557_
	);
	LUT4 #(
		.INIT('h5754)
	) name343 (
		\datai[4]_pad ,
		_w275_,
		_w277_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h6)
	) name344 (
		\reg3_reg[3]/NET0131 ,
		\reg3_reg[4]/NET0131 ,
		_w559_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name345 (
		\reg1_reg[4]/NET0131 ,
		_w234_,
		_w243_,
		_w559_,
		_w560_
	);
	LUT4 #(
		.INIT('hff35)
	) name346 (
		\reg0_reg[4]/NET0131 ,
		\reg2_reg[4]/NET0131 ,
		_w234_,
		_w243_,
		_w561_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		_w560_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h7)
	) name348 (
		_w560_,
		_w561_,
		_w563_
	);
	LUT3 #(
		.INIT('h40)
	) name349 (
		_w558_,
		_w560_,
		_w561_,
		_w564_
	);
	LUT4 #(
		.INIT('h785a)
	) name350 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\IR_reg[5]/NET0131 ,
		_w217_,
		_w565_
	);
	LUT4 #(
		.INIT('haba8)
	) name351 (
		\datai[5]_pad ,
		_w275_,
		_w277_,
		_w565_,
		_w566_
	);
	LUT3 #(
		.INIT('h80)
	) name352 (
		_w246_,
		_w250_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w564_,
		_w567_,
		_w568_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name354 (
		\reg0_reg[2]/NET0131 ,
		\reg1_reg[2]/NET0131 ,
		_w234_,
		_w243_,
		_w569_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name355 (
		\reg2_reg[2]/NET0131 ,
		\reg3_reg[2]/NET0131 ,
		_w234_,
		_w243_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h7)
	) name357 (
		_w569_,
		_w570_,
		_w572_
	);
	LUT4 #(
		.INIT('he10f)
	) name358 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w573_
	);
	LUT4 #(
		.INIT('h5754)
	) name359 (
		\datai[2]_pad ,
		_w275_,
		_w277_,
		_w573_,
		_w574_
	);
	LUT3 #(
		.INIT('h08)
	) name360 (
		_w569_,
		_w570_,
		_w574_,
		_w575_
	);
	LUT4 #(
		.INIT('hc5ff)
	) name361 (
		\reg1_reg[3]/NET0131 ,
		\reg3_reg[3]/NET0131 ,
		_w234_,
		_w243_,
		_w576_
	);
	LUT4 #(
		.INIT('hff35)
	) name362 (
		\reg0_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w234_,
		_w243_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		_w576_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h7)
	) name364 (
		_w576_,
		_w577_,
		_w579_
	);
	LUT4 #(
		.INIT('hfe00)
	) name365 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[2]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w580_
	);
	LUT2 #(
		.INIT('h6)
	) name366 (
		\IR_reg[3]/NET0131 ,
		_w580_,
		_w581_
	);
	LUT4 #(
		.INIT('h5457)
	) name367 (
		\datai[3]_pad ,
		_w275_,
		_w277_,
		_w581_,
		_w582_
	);
	LUT3 #(
		.INIT('h08)
	) name368 (
		_w576_,
		_w577_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w575_,
		_w583_,
		_w584_
	);
	LUT4 #(
		.INIT('h35ff)
	) name370 (
		\reg1_reg[1]/NET0131 ,
		\reg3_reg[1]/NET0131 ,
		_w234_,
		_w243_,
		_w585_
	);
	LUT4 #(
		.INIT('hff35)
	) name371 (
		\reg0_reg[1]/NET0131 ,
		\reg2_reg[1]/NET0131 ,
		_w234_,
		_w243_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w585_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h7)
	) name373 (
		_w585_,
		_w586_,
		_w588_
	);
	LUT3 #(
		.INIT('h93)
	) name374 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w589_
	);
	LUT4 #(
		.INIT('h5754)
	) name375 (
		\datai[1]_pad ,
		_w275_,
		_w277_,
		_w589_,
		_w590_
	);
	LUT3 #(
		.INIT('h08)
	) name376 (
		_w585_,
		_w586_,
		_w590_,
		_w591_
	);
	LUT3 #(
		.INIT('h70)
	) name377 (
		_w585_,
		_w586_,
		_w590_,
		_w592_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name378 (
		\reg0_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w234_,
		_w243_,
		_w593_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name379 (
		\reg2_reg[0]/NET0131 ,
		\reg3_reg[0]/NET0131 ,
		_w234_,
		_w243_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h7)
	) name381 (
		_w593_,
		_w594_,
		_w596_
	);
	LUT4 #(
		.INIT('h3335)
	) name382 (
		\IR_reg[0]/NET0131 ,
		\datai[0]_pad ,
		_w275_,
		_w277_,
		_w597_
	);
	LUT3 #(
		.INIT('h08)
	) name383 (
		_w593_,
		_w594_,
		_w597_,
		_w598_
	);
	LUT3 #(
		.INIT('h23)
	) name384 (
		_w592_,
		_w591_,
		_w598_,
		_w599_
	);
	LUT3 #(
		.INIT('h70)
	) name385 (
		_w576_,
		_w577_,
		_w582_,
		_w600_
	);
	LUT3 #(
		.INIT('h70)
	) name386 (
		_w569_,
		_w570_,
		_w574_,
		_w601_
	);
	LUT3 #(
		.INIT('h32)
	) name387 (
		_w600_,
		_w583_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('haa80)
	) name388 (
		_w568_,
		_w584_,
		_w599_,
		_w602_,
		_w603_
	);
	LUT3 #(
		.INIT('h07)
	) name389 (
		_w246_,
		_w250_,
		_w566_,
		_w604_
	);
	LUT3 #(
		.INIT('h2a)
	) name390 (
		_w558_,
		_w560_,
		_w561_,
		_w605_
	);
	LUT3 #(
		.INIT('h45)
	) name391 (
		_w604_,
		_w567_,
		_w605_,
		_w606_
	);
	LUT3 #(
		.INIT('h2a)
	) name392 (
		_w540_,
		_w541_,
		_w543_,
		_w607_
	);
	LUT3 #(
		.INIT('h07)
	) name393 (
		_w547_,
		_w549_,
		_w554_,
		_w608_
	);
	LUT3 #(
		.INIT('h54)
	) name394 (
		_w555_,
		_w607_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('h0075)
	) name395 (
		_w556_,
		_w603_,
		_w606_,
		_w609_,
		_w610_
	);
	LUT4 #(
		.INIT('h0b02)
	) name396 (
		_w260_,
		_w474_,
		_w487_,
		_w534_,
		_w611_
	);
	LUT3 #(
		.INIT('h31)
	) name397 (
		_w472_,
		_w488_,
		_w611_,
		_w612_
	);
	LUT3 #(
		.INIT('h80)
	) name398 (
		_w521_,
		_w522_,
		_w527_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w519_,
		_w613_,
		_w614_
	);
	LUT4 #(
		.INIT('h00d4)
	) name400 (
		_w512_,
		_w516_,
		_w613_,
		_w531_,
		_w615_
	);
	LUT3 #(
		.INIT('h51)
	) name401 (
		_w530_,
		_w510_,
		_w615_,
		_w616_
	);
	LUT3 #(
		.INIT('ha8)
	) name402 (
		_w491_,
		_w612_,
		_w616_,
		_w617_
	);
	LUT3 #(
		.INIT('h80)
	) name403 (
		_w436_,
		_w439_,
		_w440_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w444_,
		_w618_,
		_w619_
	);
	LUT4 #(
		.INIT('h0001)
	) name405 (
		_w413_,
		_w424_,
		_w444_,
		_w618_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w452_,
		_w620_,
		_w621_
	);
	LUT4 #(
		.INIT('h5700)
	) name407 (
		_w491_,
		_w612_,
		_w616_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h80aa)
	) name408 (
		_w454_,
		_w538_,
		_w610_,
		_w622_,
		_w623_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name409 (
		_w319_,
		_w362_,
		_w358_,
		_w623_,
		_w624_
	);
	LUT3 #(
		.INIT('h15)
	) name410 (
		_w279_,
		_w292_,
		_w293_,
		_w625_
	);
	LUT4 #(
		.INIT('h0777)
	) name411 (
		_w292_,
		_w293_,
		_w297_,
		_w298_,
		_w626_
	);
	LUT3 #(
		.INIT('h51)
	) name412 (
		_w625_,
		_w296_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('h0233)
	) name413 (
		_w317_,
		_w302_,
		_w624_,
		_w627_,
		_w628_
	);
	LUT3 #(
		.INIT('h2a)
	) name414 (
		\IR_reg[31]/NET0131 ,
		_w225_,
		_w238_,
		_w629_
	);
	LUT4 #(
		.INIT('h55a6)
	) name415 (
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w237_,
		_w629_,
		_w630_
	);
	LUT3 #(
		.INIT('he0)
	) name416 (
		\IR_reg[20]/NET0131 ,
		\IR_reg[21]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w631_
	);
	LUT3 #(
		.INIT('h56)
	) name417 (
		\IR_reg[22]/NET0131 ,
		_w271_,
		_w631_,
		_w632_
	);
	LUT4 #(
		.INIT('h4448)
	) name418 (
		\IR_reg[22]/NET0131 ,
		_w630_,
		_w271_,
		_w631_,
		_w633_
	);
	LUT3 #(
		.INIT('h84)
	) name419 (
		_w272_,
		_w633_,
		_w628_,
		_w634_
	);
	LUT3 #(
		.INIT('h80)
	) name420 (
		_w279_,
		_w292_,
		_w293_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w635_,
		_w301_,
		_w636_
	);
	LUT3 #(
		.INIT('h80)
	) name422 (
		_w296_,
		_w297_,
		_w298_,
		_w637_
	);
	LUT4 #(
		.INIT('h0515)
	) name423 (
		_w625_,
		_w637_,
		_w636_,
		_w317_,
		_w638_
	);
	LUT4 #(
		.INIT('h0001)
	) name424 (
		_w499_,
		_w509_,
		_w519_,
		_w613_,
		_w639_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name425 (
		_w536_,
		_w538_,
		_w610_,
		_w639_,
		_w640_
	);
	LUT4 #(
		.INIT('h5d00)
	) name426 (
		_w454_,
		_w621_,
		_w640_,
		_w362_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w625_,
		_w637_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w642_,
		_w319_,
		_w643_
	);
	LUT4 #(
		.INIT('h0155)
	) name429 (
		_w638_,
		_w641_,
		_w358_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h2221)
	) name430 (
		\IR_reg[22]/NET0131 ,
		_w630_,
		_w271_,
		_w631_,
		_w645_
	);
	LUT3 #(
		.INIT('h84)
	) name431 (
		_w272_,
		_w645_,
		_w644_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w604_,
		_w607_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w600_,
		_w605_,
		_w648_
	);
	LUT3 #(
		.INIT('h70)
	) name434 (
		_w593_,
		_w594_,
		_w597_,
		_w649_
	);
	LUT4 #(
		.INIT('h002b)
	) name435 (
		_w587_,
		_w590_,
		_w649_,
		_w601_,
		_w650_
	);
	LUT4 #(
		.INIT('h22a2)
	) name436 (
		_w568_,
		_w648_,
		_w584_,
		_w650_,
		_w651_
	);
	LUT3 #(
		.INIT('h01)
	) name437 (
		_w476_,
		_w518_,
		_w531_,
		_w652_
	);
	LUT4 #(
		.INIT('h0001)
	) name438 (
		_w485_,
		_w530_,
		_w528_,
		_w608_,
		_w653_
	);
	LUT3 #(
		.INIT('h80)
	) name439 (
		_w489_,
		_w652_,
		_w653_,
		_w654_
	);
	LUT4 #(
		.INIT('h5d00)
	) name440 (
		_w556_,
		_w647_,
		_w651_,
		_w654_,
		_w655_
	);
	LUT4 #(
		.INIT('h0001)
	) name441 (
		_w446_,
		_w447_,
		_w434_,
		_w443_,
		_w656_
	);
	LUT3 #(
		.INIT('h80)
	) name442 (
		_w402_,
		_w397_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w371_,
		_w398_,
		_w658_
	);
	LUT3 #(
		.INIT('h01)
	) name444 (
		_w371_,
		_w398_,
		_w450_,
		_w659_
	);
	LUT4 #(
		.INIT('h4054)
	) name445 (
		_w400_,
		_w363_,
		_w369_,
		_w388_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('h5440)
	) name447 (
		_w447_,
		_w429_,
		_w433_,
		_w618_,
		_w662_
	);
	LUT4 #(
		.INIT('h2232)
	) name448 (
		_w446_,
		_w379_,
		_w425_,
		_w662_,
		_w663_
	);
	LUT3 #(
		.INIT('h8a)
	) name449 (
		_w404_,
		_w661_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h001f)
	) name450 (
		_w617_,
		_w655_,
		_w657_,
		_w664_,
		_w665_
	);
	LUT3 #(
		.INIT('h0e)
	) name451 (
		_w310_,
		_w315_,
		_w355_,
		_w666_
	);
	LUT3 #(
		.INIT('h01)
	) name452 (
		_w635_,
		_w308_,
		_w301_,
		_w667_
	);
	LUT4 #(
		.INIT('h0001)
	) name453 (
		_w635_,
		_w308_,
		_w301_,
		_w356_,
		_w668_
	);
	LUT3 #(
		.INIT('h80)
	) name454 (
		_w666_,
		_w353_,
		_w668_,
		_w669_
	);
	LUT3 #(
		.INIT('h54)
	) name455 (
		_w635_,
		_w625_,
		_w637_,
		_w670_
	);
	LUT3 #(
		.INIT('h15)
	) name456 (
		_w343_,
		_w345_,
		_w351_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w344_,
		_w356_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w327_,
		_w335_,
		_w673_
	);
	LUT4 #(
		.INIT('h20aa)
	) name459 (
		_w666_,
		_w671_,
		_w672_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h1151)
	) name460 (
		_w670_,
		_w667_,
		_w319_,
		_w674_,
		_w675_
	);
	LUT3 #(
		.INIT('hb0)
	) name461 (
		_w665_,
		_w669_,
		_w675_,
		_w676_
	);
	LUT4 #(
		.INIT('h2228)
	) name462 (
		\B_reg/NET0131 ,
		\IR_reg[23]/NET0131 ,
		_w264_,
		_w267_,
		_w677_
	);
	LUT4 #(
		.INIT('h1112)
	) name463 (
		\IR_reg[22]/NET0131 ,
		_w630_,
		_w271_,
		_w631_,
		_w678_
	);
	LUT4 #(
		.INIT('hf600)
	) name464 (
		_w676_,
		_w272_,
		_w677_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h0100)
	) name465 (
		_w336_,
		_w339_,
		_w338_,
		_w340_,
		_w680_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name466 (
		_w336_,
		_w339_,
		_w338_,
		_w340_,
		_w681_
	);
	LUT4 #(
		.INIT('h5655)
	) name467 (
		_w336_,
		_w339_,
		_w338_,
		_w340_,
		_w682_
	);
	LUT4 #(
		.INIT('h5655)
	) name468 (
		_w406_,
		_w409_,
		_w408_,
		_w410_,
		_w683_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name469 (
		_w389_,
		_w392_,
		_w391_,
		_w393_,
		_w684_
	);
	LUT4 #(
		.INIT('h0100)
	) name470 (
		_w389_,
		_w392_,
		_w391_,
		_w393_,
		_w685_
	);
	LUT4 #(
		.INIT('h5655)
	) name471 (
		_w389_,
		_w392_,
		_w391_,
		_w393_,
		_w686_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name472 (
		_w417_,
		_w420_,
		_w419_,
		_w421_,
		_w687_
	);
	LUT4 #(
		.INIT('h0100)
	) name473 (
		_w417_,
		_w420_,
		_w419_,
		_w421_,
		_w688_
	);
	LUT4 #(
		.INIT('h5655)
	) name474 (
		_w417_,
		_w420_,
		_w419_,
		_w421_,
		_w689_
	);
	LUT4 #(
		.INIT('h0004)
	) name475 (
		_w682_,
		_w683_,
		_w686_,
		_w689_,
		_w690_
	);
	LUT4 #(
		.INIT('h0006)
	) name476 (
		_w279_,
		_w294_,
		_w637_,
		_w301_,
		_w691_
	);
	LUT3 #(
		.INIT('h08)
	) name477 (
		_w477_,
		_w479_,
		_w484_,
		_w692_
	);
	LUT3 #(
		.INIT('h70)
	) name478 (
		_w477_,
		_w479_,
		_w484_,
		_w693_
	);
	LUT3 #(
		.INIT('h87)
	) name479 (
		_w477_,
		_w479_,
		_w484_,
		_w694_
	);
	LUT3 #(
		.INIT('h95)
	) name480 (
		_w540_,
		_w541_,
		_w543_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT4 #(
		.INIT('h10ef)
	) name482 (
		_w456_,
		_w457_,
		_w458_,
		_w462_,
		_w697_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name483 (
		_w328_,
		_w331_,
		_w330_,
		_w332_,
		_w698_
	);
	LUT4 #(
		.INIT('h0100)
	) name484 (
		_w328_,
		_w331_,
		_w330_,
		_w332_,
		_w699_
	);
	LUT4 #(
		.INIT('h5655)
	) name485 (
		_w328_,
		_w331_,
		_w330_,
		_w332_,
		_w700_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		_w697_,
		_w700_,
		_w701_
	);
	LUT4 #(
		.INIT('h8000)
	) name487 (
		_w691_,
		_w696_,
		_w701_,
		_w690_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w345_,
		_w351_,
		_w703_
	);
	LUT2 #(
		.INIT('h9)
	) name489 (
		_w345_,
		_w351_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w310_,
		_w315_,
		_w705_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		_w310_,
		_w315_,
		_w706_
	);
	LUT2 #(
		.INIT('h9)
	) name492 (
		_w310_,
		_w315_,
		_w707_
	);
	LUT4 #(
		.INIT('h0660)
	) name493 (
		_w310_,
		_w315_,
		_w345_,
		_w351_,
		_w708_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name494 (
		_w381_,
		_w384_,
		_w383_,
		_w385_,
		_w709_
	);
	LUT4 #(
		.INIT('h0100)
	) name495 (
		_w381_,
		_w384_,
		_w383_,
		_w385_,
		_w710_
	);
	LUT4 #(
		.INIT('h5655)
	) name496 (
		_w381_,
		_w384_,
		_w383_,
		_w385_,
		_w711_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name497 (
		_w372_,
		_w375_,
		_w374_,
		_w376_,
		_w712_
	);
	LUT4 #(
		.INIT('h0100)
	) name498 (
		_w372_,
		_w375_,
		_w374_,
		_w376_,
		_w713_
	);
	LUT4 #(
		.INIT('h5655)
	) name499 (
		_w372_,
		_w375_,
		_w374_,
		_w376_,
		_w714_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name500 (
		_w363_,
		_w367_,
		_w366_,
		_w368_,
		_w715_
	);
	LUT4 #(
		.INIT('h0100)
	) name501 (
		_w363_,
		_w367_,
		_w366_,
		_w368_,
		_w716_
	);
	LUT4 #(
		.INIT('h5655)
	) name502 (
		_w363_,
		_w367_,
		_w366_,
		_w368_,
		_w717_
	);
	LUT4 #(
		.INIT('h0100)
	) name503 (
		_w320_,
		_w323_,
		_w322_,
		_w324_,
		_w718_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name504 (
		_w320_,
		_w323_,
		_w322_,
		_w324_,
		_w719_
	);
	LUT4 #(
		.INIT('h5655)
	) name505 (
		_w320_,
		_w323_,
		_w322_,
		_w324_,
		_w720_
	);
	LUT4 #(
		.INIT('h0001)
	) name506 (
		_w711_,
		_w714_,
		_w717_,
		_w720_,
		_w721_
	);
	LUT3 #(
		.INIT('h95)
	) name507 (
		_w493_,
		_w495_,
		_w496_,
		_w722_
	);
	LUT3 #(
		.INIT('h08)
	) name508 (
		_w246_,
		_w250_,
		_w566_,
		_w723_
	);
	LUT3 #(
		.INIT('h70)
	) name509 (
		_w246_,
		_w250_,
		_w566_,
		_w724_
	);
	LUT3 #(
		.INIT('h87)
	) name510 (
		_w246_,
		_w250_,
		_w566_,
		_w725_
	);
	LUT3 #(
		.INIT('h08)
	) name511 (
		_w426_,
		_w428_,
		_w433_,
		_w726_
	);
	LUT3 #(
		.INIT('h70)
	) name512 (
		_w426_,
		_w428_,
		_w433_,
		_w727_
	);
	LUT3 #(
		.INIT('h87)
	) name513 (
		_w426_,
		_w428_,
		_w433_,
		_w728_
	);
	LUT3 #(
		.INIT('h6a)
	) name514 (
		_w303_,
		_w304_,
		_w305_,
		_w729_
	);
	LUT4 #(
		.INIT('h0200)
	) name515 (
		_w722_,
		_w725_,
		_w728_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('h08)
	) name516 (
		_w547_,
		_w549_,
		_w554_,
		_w731_
	);
	LUT3 #(
		.INIT('h70)
	) name517 (
		_w547_,
		_w549_,
		_w554_,
		_w732_
	);
	LUT3 #(
		.INIT('h87)
	) name518 (
		_w547_,
		_w549_,
		_w554_,
		_w733_
	);
	LUT3 #(
		.INIT('h95)
	) name519 (
		_w558_,
		_w560_,
		_w561_,
		_w734_
	);
	LUT3 #(
		.INIT('h87)
	) name520 (
		_w593_,
		_w594_,
		_w597_,
		_w735_
	);
	LUT3 #(
		.INIT('h70)
	) name521 (
		_w521_,
		_w522_,
		_w527_,
		_w736_
	);
	LUT3 #(
		.INIT('h08)
	) name522 (
		_w521_,
		_w522_,
		_w527_,
		_w737_
	);
	LUT3 #(
		.INIT('h87)
	) name523 (
		_w521_,
		_w522_,
		_w527_,
		_w738_
	);
	LUT4 #(
		.INIT('h0040)
	) name524 (
		_w733_,
		_w734_,
		_w735_,
		_w738_,
		_w739_
	);
	LUT3 #(
		.INIT('h80)
	) name525 (
		_w576_,
		_w577_,
		_w582_,
		_w740_
	);
	LUT3 #(
		.INIT('h07)
	) name526 (
		_w576_,
		_w577_,
		_w582_,
		_w741_
	);
	LUT3 #(
		.INIT('h78)
	) name527 (
		_w576_,
		_w577_,
		_w582_,
		_w742_
	);
	LUT3 #(
		.INIT('h87)
	) name528 (
		_w258_,
		_w259_,
		_w474_,
		_w743_
	);
	LUT3 #(
		.INIT('h08)
	) name529 (
		_w465_,
		_w466_,
		_w470_,
		_w744_
	);
	LUT3 #(
		.INIT('h70)
	) name530 (
		_w465_,
		_w466_,
		_w470_,
		_w745_
	);
	LUT3 #(
		.INIT('h87)
	) name531 (
		_w465_,
		_w466_,
		_w470_,
		_w746_
	);
	LUT3 #(
		.INIT('h87)
	) name532 (
		_w569_,
		_w570_,
		_w574_,
		_w747_
	);
	LUT4 #(
		.INIT('h0400)
	) name533 (
		_w742_,
		_w743_,
		_w746_,
		_w747_,
		_w748_
	);
	LUT3 #(
		.INIT('h40)
	) name534 (
		_w436_,
		_w439_,
		_w440_,
		_w749_
	);
	LUT3 #(
		.INIT('h2a)
	) name535 (
		_w436_,
		_w439_,
		_w440_,
		_w750_
	);
	LUT3 #(
		.INIT('h95)
	) name536 (
		_w436_,
		_w439_,
		_w440_,
		_w751_
	);
	LUT3 #(
		.INIT('h70)
	) name537 (
		_w501_,
		_w502_,
		_w508_,
		_w752_
	);
	LUT3 #(
		.INIT('h08)
	) name538 (
		_w501_,
		_w502_,
		_w508_,
		_w753_
	);
	LUT3 #(
		.INIT('h87)
	) name539 (
		_w501_,
		_w502_,
		_w508_,
		_w754_
	);
	LUT3 #(
		.INIT('h95)
	) name540 (
		_w512_,
		_w514_,
		_w515_,
		_w755_
	);
	LUT3 #(
		.INIT('h87)
	) name541 (
		_w585_,
		_w586_,
		_w590_,
		_w756_
	);
	LUT4 #(
		.INIT('h1000)
	) name542 (
		_w751_,
		_w754_,
		_w755_,
		_w756_,
		_w757_
	);
	LUT4 #(
		.INIT('h8000)
	) name543 (
		_w748_,
		_w757_,
		_w730_,
		_w739_,
		_w758_
	);
	LUT4 #(
		.INIT('h8000)
	) name544 (
		_w721_,
		_w758_,
		_w702_,
		_w708_,
		_w759_
	);
	LUT4 #(
		.INIT('h171d)
	) name545 (
		_w630_,
		_w272_,
		_w677_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('h9996)
	) name546 (
		\IR_reg[22]/NET0131 ,
		_w630_,
		_w271_,
		_w631_,
		_w761_
	);
	LUT3 #(
		.INIT('h21)
	) name547 (
		\IR_reg[20]/NET0131 ,
		_w630_,
		_w271_,
		_w762_
	);
	LUT3 #(
		.INIT('h02)
	) name548 (
		_w677_,
		_w761_,
		_w762_,
		_w763_
	);
	LUT3 #(
		.INIT('h0e)
	) name549 (
		_w632_,
		_w760_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w679_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name551 (
		_w269_,
		_w646_,
		_w634_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('he)
	) name552 (
		_w270_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		\IR_reg[31]/NET0131 ,
		_w228_,
		_w768_
	);
	LUT3 #(
		.INIT('h56)
	) name554 (
		\IR_reg[24]/NET0131 ,
		_w271_,
		_w768_,
		_w769_
	);
	LUT4 #(
		.INIT('hd555)
	) name555 (
		\IR_reg[31]/NET0131 ,
		_w219_,
		_w222_,
		_w230_,
		_w770_
	);
	LUT2 #(
		.INIT('h9)
	) name556 (
		\IR_reg[26]/NET0131 ,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w769_,
		_w771_,
		_w772_
	);
	LUT4 #(
		.INIT('h0001)
	) name558 (
		\IR_reg[21]/NET0131 ,
		\IR_reg[22]/NET0131 ,
		\IR_reg[23]/NET0131 ,
		\IR_reg[24]/NET0131 ,
		_w773_
	);
	LUT4 #(
		.INIT('h0d05)
	) name559 (
		\IR_reg[31]/NET0131 ,
		_w237_,
		_w629_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h9)
	) name560 (
		\IR_reg[25]/NET0131 ,
		_w774_,
		_w775_
	);
	LUT4 #(
		.INIT('h6669)
	) name561 (
		\B_reg/NET0131 ,
		\IR_reg[24]/NET0131 ,
		_w271_,
		_w768_,
		_w776_
	);
	LUT3 #(
		.INIT('h21)
	) name562 (
		\IR_reg[26]/NET0131 ,
		\d_reg[0]/NET0131 ,
		_w770_,
		_w777_
	);
	LUT3 #(
		.INIT('he0)
	) name563 (
		_w775_,
		_w776_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w772_,
		_w778_,
		_w779_
	);
	LUT4 #(
		.INIT('hb8bc)
	) name565 (
		\d_reg[1]/NET0131 ,
		_w771_,
		_w775_,
		_w776_,
		_w780_
	);
	LUT3 #(
		.INIT('h10)
	) name566 (
		_w772_,
		_w778_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name567 (
		_w312_,
		_w772_,
		_w778_,
		_w780_,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w620_,
		_w536_,
		_w783_
	);
	LUT4 #(
		.INIT('h7500)
	) name569 (
		_w533_,
		_w610_,
		_w639_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('hf800)
	) name570 (
		_w472_,
		_w486_,
		_w490_,
		_w620_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w449_,
		_w785_,
		_w786_
	);
	LUT3 #(
		.INIT('h40)
	) name572 (
		_w359_,
		_w452_,
		_w361_,
		_w787_
	);
	LUT3 #(
		.INIT('h0b)
	) name573 (
		_w404_,
		_w362_,
		_w358_,
		_w788_
	);
	LUT4 #(
		.INIT('h4f00)
	) name574 (
		_w784_,
		_w786_,
		_w787_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('h0b07)
	) name575 (
		_w707_,
		_w781_,
		_w782_,
		_w789_,
		_w790_
	);
	LUT4 #(
		.INIT('h404a)
	) name576 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w791_
	);
	LUT3 #(
		.INIT('h80)
	) name577 (
		_w258_,
		_w259_,
		_w474_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w692_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h1000)
	) name579 (
		_w456_,
		_w457_,
		_w458_,
		_w462_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w744_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h0001)
	) name581 (
		_w692_,
		_w744_,
		_w792_,
		_w794_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w726_,
		_w749_,
		_w797_
	);
	LUT4 #(
		.INIT('h0200)
	) name583 (
		_w406_,
		_w409_,
		_w408_,
		_w410_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w688_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h0001)
	) name585 (
		_w726_,
		_w749_,
		_w688_,
		_w798_,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		_w796_,
		_w800_,
		_w801_
	);
	LUT3 #(
		.INIT('h80)
	) name587 (
		_w493_,
		_w495_,
		_w496_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w753_,
		_w802_,
		_w803_
	);
	LUT3 #(
		.INIT('h15)
	) name589 (
		_w512_,
		_w514_,
		_w515_,
		_w804_
	);
	LUT3 #(
		.INIT('h80)
	) name590 (
		_w512_,
		_w514_,
		_w515_,
		_w805_
	);
	LUT3 #(
		.INIT('h31)
	) name591 (
		_w736_,
		_w804_,
		_w805_,
		_w806_
	);
	LUT3 #(
		.INIT('h15)
	) name592 (
		_w493_,
		_w495_,
		_w496_,
		_w807_
	);
	LUT3 #(
		.INIT('h32)
	) name593 (
		_w752_,
		_w802_,
		_w807_,
		_w808_
	);
	LUT3 #(
		.INIT('h0d)
	) name594 (
		_w803_,
		_w806_,
		_w808_,
		_w809_
	);
	LUT3 #(
		.INIT('h80)
	) name595 (
		_w540_,
		_w541_,
		_w543_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w731_,
		_w810_,
		_w811_
	);
	LUT3 #(
		.INIT('h80)
	) name597 (
		_w558_,
		_w560_,
		_w561_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w723_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h07)
	) name599 (
		_w585_,
		_w586_,
		_w590_,
		_w814_
	);
	LUT3 #(
		.INIT('h07)
	) name600 (
		_w593_,
		_w594_,
		_w597_,
		_w815_
	);
	LUT3 #(
		.INIT('h80)
	) name601 (
		_w585_,
		_w586_,
		_w590_,
		_w816_
	);
	LUT3 #(
		.INIT('h51)
	) name602 (
		_w814_,
		_w815_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h80)
	) name603 (
		_w569_,
		_w570_,
		_w574_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w740_,
		_w818_,
		_w819_
	);
	LUT3 #(
		.INIT('h07)
	) name605 (
		_w569_,
		_w570_,
		_w574_,
		_w820_
	);
	LUT3 #(
		.INIT('h54)
	) name606 (
		_w740_,
		_w741_,
		_w820_,
		_w821_
	);
	LUT4 #(
		.INIT('haa20)
	) name607 (
		_w813_,
		_w817_,
		_w819_,
		_w821_,
		_w822_
	);
	LUT3 #(
		.INIT('h15)
	) name608 (
		_w558_,
		_w560_,
		_w561_,
		_w823_
	);
	LUT3 #(
		.INIT('h23)
	) name609 (
		_w723_,
		_w724_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('h15)
	) name610 (
		_w540_,
		_w541_,
		_w543_,
		_w825_
	);
	LUT3 #(
		.INIT('h23)
	) name611 (
		_w731_,
		_w732_,
		_w825_,
		_w826_
	);
	LUT3 #(
		.INIT('hd0)
	) name612 (
		_w811_,
		_w824_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w737_,
		_w805_,
		_w828_
	);
	LUT4 #(
		.INIT('h0001)
	) name614 (
		_w737_,
		_w753_,
		_w802_,
		_w805_,
		_w829_
	);
	LUT4 #(
		.INIT('h8f00)
	) name615 (
		_w811_,
		_w822_,
		_w827_,
		_w829_,
		_w830_
	);
	LUT3 #(
		.INIT('h07)
	) name616 (
		_w258_,
		_w259_,
		_w474_,
		_w831_
	);
	LUT3 #(
		.INIT('h0d)
	) name617 (
		_w693_,
		_w792_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h00ef)
	) name618 (
		_w456_,
		_w457_,
		_w458_,
		_w462_,
		_w833_
	);
	LUT3 #(
		.INIT('h23)
	) name619 (
		_w744_,
		_w745_,
		_w833_,
		_w834_
	);
	LUT3 #(
		.INIT('hd0)
	) name620 (
		_w795_,
		_w832_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h08cc)
	) name621 (
		_w795_,
		_w800_,
		_w832_,
		_w834_,
		_w836_
	);
	LUT3 #(
		.INIT('h54)
	) name622 (
		_w726_,
		_w727_,
		_w750_,
		_w837_
	);
	LUT4 #(
		.INIT('h5455)
	) name623 (
		_w406_,
		_w409_,
		_w408_,
		_w410_,
		_w838_
	);
	LUT3 #(
		.INIT('h0d)
	) name624 (
		_w687_,
		_w798_,
		_w838_,
		_w839_
	);
	LUT3 #(
		.INIT('h70)
	) name625 (
		_w799_,
		_w837_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w836_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('h5d00)
	) name627 (
		_w801_,
		_w809_,
		_w830_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w699_,
		_w718_,
		_w843_
	);
	LUT3 #(
		.INIT('h01)
	) name629 (
		_w699_,
		_w718_,
		_w680_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w703_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w710_,
		_w716_,
		_w846_
	);
	LUT3 #(
		.INIT('h01)
	) name632 (
		_w710_,
		_w716_,
		_w685_,
		_w847_
	);
	LUT4 #(
		.INIT('h0001)
	) name633 (
		_w710_,
		_w713_,
		_w716_,
		_w685_,
		_w848_
	);
	LUT3 #(
		.INIT('h40)
	) name634 (
		_w703_,
		_w844_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w712_,
		_w715_,
		_w850_
	);
	LUT3 #(
		.INIT('h45)
	) name636 (
		_w709_,
		_w710_,
		_w684_,
		_w851_
	);
	LUT4 #(
		.INIT('h0b02)
	) name637 (
		_w381_,
		_w386_,
		_w716_,
		_w684_,
		_w852_
	);
	LUT3 #(
		.INIT('h51)
	) name638 (
		_w713_,
		_w850_,
		_w852_,
		_w853_
	);
	LUT4 #(
		.INIT('h00fd)
	) name639 (
		_w345_,
		_w351_,
		_w680_,
		_w681_,
		_w854_
	);
	LUT4 #(
		.INIT('h1303)
	) name640 (
		_w698_,
		_w719_,
		_w843_,
		_w854_,
		_w855_
	);
	LUT3 #(
		.INIT('h70)
	) name641 (
		_w845_,
		_w853_,
		_w855_,
		_w856_
	);
	LUT4 #(
		.INIT('h65aa)
	) name642 (
		_w707_,
		_w842_,
		_w849_,
		_w856_,
		_w857_
	);
	LUT4 #(
		.INIT('h1a10)
	) name643 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w858_
	);
	LUT4 #(
		.INIT('h2e00)
	) name644 (
		_w312_,
		_w781_,
		_w857_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h8000)
	) name645 (
		_w582_,
		_w574_,
		_w590_,
		_w597_,
		_w860_
	);
	LUT3 #(
		.INIT('h40)
	) name646 (
		_w566_,
		_w558_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		_w540_,
		_w554_,
		_w862_
	);
	LUT4 #(
		.INIT('h4000)
	) name648 (
		_w566_,
		_w558_,
		_w860_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		_w512_,
		_w527_,
		_w864_
	);
	LUT4 #(
		.INIT('h0020)
	) name650 (
		_w474_,
		_w484_,
		_w493_,
		_w508_,
		_w865_
	);
	LUT3 #(
		.INIT('h80)
	) name651 (
		_w863_,
		_w864_,
		_w865_,
		_w866_
	);
	LUT3 #(
		.INIT('h02)
	) name652 (
		_w462_,
		_w470_,
		_w436_,
		_w867_
	);
	LUT4 #(
		.INIT('h0002)
	) name653 (
		_w462_,
		_w470_,
		_w433_,
		_w436_,
		_w868_
	);
	LUT4 #(
		.INIT('h8000)
	) name654 (
		_w863_,
		_w864_,
		_w865_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h02)
	) name655 (
		_w406_,
		_w417_,
		_w389_,
		_w870_
	);
	LUT4 #(
		.INIT('h111f)
	) name656 (
		\datai[23]_pad ,
		\datai[24]_pad ,
		_w275_,
		_w277_,
		_w871_
	);
	LUT4 #(
		.INIT('h111f)
	) name657 (
		\datai[21]_pad ,
		\datai[22]_pad ,
		_w275_,
		_w277_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w871_,
		_w872_,
		_w873_
	);
	LUT3 #(
		.INIT('h80)
	) name659 (
		_w869_,
		_w870_,
		_w873_,
		_w874_
	);
	LUT4 #(
		.INIT('h111f)
	) name660 (
		\datai[25]_pad ,
		\datai[26]_pad ,
		_w275_,
		_w277_,
		_w875_
	);
	LUT4 #(
		.INIT('h8000)
	) name661 (
		_w869_,
		_w870_,
		_w873_,
		_w875_,
		_w876_
	);
	LUT4 #(
		.INIT('h6050)
	) name662 (
		_w310_,
		_w320_,
		_w781_,
		_w876_,
		_w877_
	);
	LUT3 #(
		.INIT('h10)
	) name663 (
		_w268_,
		_w632_,
		_w762_,
		_w878_
	);
	LUT3 #(
		.INIT('he0)
	) name664 (
		_w782_,
		_w877_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h0777)
	) name665 (
		_w292_,
		_w293_,
		_w593_,
		_w594_,
		_w880_
	);
	LUT4 #(
		.INIT('h0100)
	) name666 (
		_w578_,
		_w571_,
		_w587_,
		_w880_,
		_w881_
	);
	LUT4 #(
		.INIT('h0777)
	) name667 (
		_w246_,
		_w250_,
		_w560_,
		_w561_,
		_w882_
	);
	LUT4 #(
		.INIT('h0777)
	) name668 (
		_w541_,
		_w543_,
		_w547_,
		_w549_,
		_w883_
	);
	LUT4 #(
		.INIT('h0777)
	) name669 (
		_w495_,
		_w496_,
		_w501_,
		_w502_,
		_w884_
	);
	LUT4 #(
		.INIT('h0777)
	) name670 (
		_w514_,
		_w515_,
		_w521_,
		_w522_,
		_w885_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w884_,
		_w885_,
		_w886_
	);
	LUT4 #(
		.INIT('h8000)
	) name672 (
		_w881_,
		_w882_,
		_w883_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h0777)
	) name673 (
		_w258_,
		_w259_,
		_w465_,
		_w466_,
		_w888_
	);
	LUT3 #(
		.INIT('h10)
	) name674 (
		_w459_,
		_w480_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		_w887_,
		_w889_,
		_w890_
	);
	LUT4 #(
		.INIT('h0777)
	) name676 (
		_w426_,
		_w428_,
		_w439_,
		_w440_,
		_w891_
	);
	LUT3 #(
		.INIT('h10)
	) name677 (
		_w411_,
		_w422_,
		_w891_,
		_w892_
	);
	LUT3 #(
		.INIT('h80)
	) name678 (
		_w887_,
		_w889_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w369_,
		_w386_,
		_w894_
	);
	LUT4 #(
		.INIT('h0001)
	) name680 (
		_w377_,
		_w369_,
		_w386_,
		_w394_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w341_,
		_w351_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w325_,
		_w333_,
		_w898_
	);
	LUT3 #(
		.INIT('h01)
	) name684 (
		_w315_,
		_w325_,
		_w333_,
		_w899_
	);
	LUT3 #(
		.INIT('h80)
	) name685 (
		_w895_,
		_w896_,
		_w899_,
		_w900_
	);
	LUT4 #(
		.INIT('h8000)
	) name686 (
		_w887_,
		_w889_,
		_w892_,
		_w900_,
		_w901_
	);
	LUT4 #(
		.INIT('h0200)
	) name687 (
		_w277_,
		_w323_,
		_w322_,
		_w324_,
		_w902_
	);
	LUT4 #(
		.INIT('h00eb)
	) name688 (
		_w277_,
		_w306_,
		_w901_,
		_w902_,
		_w903_
	);
	LUT3 #(
		.INIT('h80)
	) name689 (
		_w268_,
		_w632_,
		_w762_,
		_w904_
	);
	LUT3 #(
		.INIT('h04)
	) name690 (
		_w268_,
		_w630_,
		_w632_,
		_w905_
	);
	LUT4 #(
		.INIT('h1000)
	) name691 (
		_w772_,
		_w778_,
		_w780_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h10)
	) name692 (
		_w268_,
		_w272_,
		_w645_,
		_w907_
	);
	LUT3 #(
		.INIT('ha8)
	) name693 (
		_w310_,
		_w906_,
		_w907_,
		_w908_
	);
	LUT3 #(
		.INIT('h08)
	) name694 (
		_w268_,
		_w632_,
		_w762_,
		_w909_
	);
	LUT4 #(
		.INIT('hef00)
	) name695 (
		_w772_,
		_w778_,
		_w780_,
		_w905_,
		_w910_
	);
	LUT4 #(
		.INIT('hef00)
	) name696 (
		_w772_,
		_w778_,
		_w780_,
		_w904_,
		_w911_
	);
	LUT4 #(
		.INIT('haaa8)
	) name697 (
		_w312_,
		_w909_,
		_w910_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w908_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('h7f00)
	) name699 (
		_w781_,
		_w903_,
		_w904_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w879_,
		_w914_,
		_w915_
	);
	LUT4 #(
		.INIT('h0b00)
	) name701 (
		_w790_,
		_w791_,
		_w859_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('h80)
	) name702 (
		_w769_,
		_w771_,
		_w775_,
		_w917_
	);
	LUT4 #(
		.INIT('h1555)
	) name703 (
		_w268_,
		_w769_,
		_w771_,
		_w775_,
		_w918_
	);
	LUT4 #(
		.INIT('h4000)
	) name704 (
		_w268_,
		_w769_,
		_w771_,
		_w775_,
		_w919_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		_w312_,
		_w919_,
		_w920_
	);
	LUT4 #(
		.INIT('haa20)
	) name706 (
		\state_reg[0]/NET0131 ,
		_w916_,
		_w918_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h2)
	) name707 (
		\reg3_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w922_
	);
	LUT3 #(
		.INIT('h07)
	) name708 (
		_w269_,
		_w312_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('hb)
	) name709 (
		_w921_,
		_w923_,
		_w924_
	);
	LUT3 #(
		.INIT('he0)
	) name710 (
		_w772_,
		_w778_,
		_w780_,
		_w925_
	);
	LUT4 #(
		.INIT('h02aa)
	) name711 (
		\reg2_reg[28]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w926_
	);
	LUT4 #(
		.INIT('hc355)
	) name712 (
		\reg2_reg[28]/NET0131 ,
		_w707_,
		_w789_,
		_w925_,
		_w927_
	);
	LUT4 #(
		.INIT('h30a0)
	) name713 (
		\reg2_reg[28]/NET0131 ,
		_w857_,
		_w858_,
		_w925_,
		_w928_
	);
	LUT4 #(
		.INIT('h6500)
	) name714 (
		_w310_,
		_w320_,
		_w876_,
		_w925_,
		_w929_
	);
	LUT3 #(
		.INIT('ha8)
	) name715 (
		_w878_,
		_w926_,
		_w929_,
		_w930_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name716 (
		\reg2_reg[28]/NET0131 ,
		_w903_,
		_w904_,
		_w925_,
		_w931_
	);
	LUT4 #(
		.INIT('h1f00)
	) name717 (
		_w772_,
		_w778_,
		_w780_,
		_w905_,
		_w932_
	);
	LUT3 #(
		.INIT('ha8)
	) name718 (
		\reg2_reg[28]/NET0131 ,
		_w909_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name719 (
		_w312_,
		_w907_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		_w310_,
		_w905_,
		_w935_
	);
	LUT3 #(
		.INIT('h13)
	) name721 (
		_w925_,
		_w934_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name722 (
		_w933_,
		_w936_,
		_w937_
	);
	LUT3 #(
		.INIT('h10)
	) name723 (
		_w930_,
		_w931_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('h0d00)
	) name724 (
		_w791_,
		_w927_,
		_w928_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		\reg2_reg[28]/NET0131 ,
		_w919_,
		_w940_
	);
	LUT4 #(
		.INIT('haa08)
	) name726 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w939_,
		_w940_,
		_w941_
	);
	LUT4 #(
		.INIT('h8884)
	) name727 (
		\IR_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w264_,
		_w267_,
		_w942_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		\reg2_reg[28]/NET0131 ,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('he)
	) name729 (
		_w941_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		\reg2_reg[29]/NET0131 ,
		_w942_,
		_w945_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		\reg2_reg[29]/NET0131 ,
		_w919_,
		_w946_
	);
	LUT4 #(
		.INIT('h0100)
	) name732 (
		_w303_,
		_w310_,
		_w320_,
		_w876_,
		_w947_
	);
	LUT4 #(
		.INIT('h5655)
	) name733 (
		_w303_,
		_w310_,
		_w320_,
		_w876_,
		_w948_
	);
	LUT4 #(
		.INIT('hc808)
	) name734 (
		\reg2_reg[29]/NET0131 ,
		_w878_,
		_w925_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		_w277_,
		_w315_,
		_w950_
	);
	LUT4 #(
		.INIT('h8828)
	) name736 (
		\B_reg/NET0131 ,
		\IR_reg[27]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		_w274_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w277_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('hef00)
	) name738 (
		_w299_,
		_w306_,
		_w901_,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('h6500)
	) name739 (
		_w299_,
		_w306_,
		_w901_,
		_w952_,
		_w954_
	);
	LUT4 #(
		.INIT('h111d)
	) name740 (
		\reg2_reg[29]/NET0131 ,
		_w925_,
		_w950_,
		_w954_,
		_w955_
	);
	LUT3 #(
		.INIT('ha8)
	) name741 (
		\reg2_reg[29]/NET0131 ,
		_w909_,
		_w932_,
		_w956_
	);
	LUT4 #(
		.INIT('h0400)
	) name742 (
		_w268_,
		_w291_,
		_w272_,
		_w645_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		_w303_,
		_w905_,
		_w958_
	);
	LUT3 #(
		.INIT('h13)
	) name744 (
		_w925_,
		_w957_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h4)
	) name745 (
		_w956_,
		_w959_,
		_w960_
	);
	LUT4 #(
		.INIT('h3100)
	) name746 (
		_w904_,
		_w949_,
		_w955_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w792_,
		_w794_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w749_,
		_w744_,
		_w963_
	);
	LUT4 #(
		.INIT('h0001)
	) name749 (
		_w749_,
		_w744_,
		_w792_,
		_w794_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w726_,
		_w688_,
		_w965_
	);
	LUT4 #(
		.INIT('h0001)
	) name751 (
		_w726_,
		_w685_,
		_w688_,
		_w798_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		_w964_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w692_,
		_w802_,
		_w968_
	);
	LUT3 #(
		.INIT('h45)
	) name754 (
		_w752_,
		_w753_,
		_w804_,
		_w969_
	);
	LUT3 #(
		.INIT('h23)
	) name755 (
		_w692_,
		_w693_,
		_w807_,
		_w970_
	);
	LUT3 #(
		.INIT('hd0)
	) name756 (
		_w968_,
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w731_,
		_w737_,
		_w972_
	);
	LUT4 #(
		.INIT('h008e)
	) name758 (
		_w587_,
		_w590_,
		_w815_,
		_w820_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w741_,
		_w823_,
		_w974_
	);
	LUT3 #(
		.INIT('h01)
	) name760 (
		_w723_,
		_w810_,
		_w812_,
		_w975_
	);
	LUT4 #(
		.INIT('h2f00)
	) name761 (
		_w819_,
		_w973_,
		_w974_,
		_w975_,
		_w976_
	);
	LUT3 #(
		.INIT('h0d)
	) name762 (
		_w724_,
		_w810_,
		_w825_,
		_w977_
	);
	LUT3 #(
		.INIT('h31)
	) name763 (
		_w732_,
		_w736_,
		_w737_,
		_w978_
	);
	LUT3 #(
		.INIT('hd0)
	) name764 (
		_w972_,
		_w977_,
		_w978_,
		_w979_
	);
	LUT3 #(
		.INIT('h70)
	) name765 (
		_w972_,
		_w976_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w753_,
		_w805_,
		_w981_
	);
	LUT4 #(
		.INIT('h0001)
	) name767 (
		_w692_,
		_w753_,
		_w802_,
		_w805_,
		_w982_
	);
	LUT4 #(
		.INIT('h8f00)
	) name768 (
		_w972_,
		_w976_,
		_w979_,
		_w982_,
		_w983_
	);
	LUT3 #(
		.INIT('h0b)
	) name769 (
		_w794_,
		_w831_,
		_w833_,
		_w984_
	);
	LUT3 #(
		.INIT('h54)
	) name770 (
		_w749_,
		_w750_,
		_w745_,
		_w985_
	);
	LUT3 #(
		.INIT('h0d)
	) name771 (
		_w963_,
		_w984_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('hcc08)
	) name772 (
		_w963_,
		_w966_,
		_w984_,
		_w985_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w684_,
		_w838_,
		_w988_
	);
	LUT3 #(
		.INIT('h31)
	) name774 (
		_w727_,
		_w687_,
		_w688_,
		_w989_
	);
	LUT4 #(
		.INIT('h00b2)
	) name775 (
		_w417_,
		_w422_,
		_w727_,
		_w798_,
		_w990_
	);
	LUT3 #(
		.INIT('h51)
	) name776 (
		_w685_,
		_w988_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w987_,
		_w991_,
		_w992_
	);
	LUT4 #(
		.INIT('h5d00)
	) name778 (
		_w967_,
		_w971_,
		_w983_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		_w705_,
		_w844_,
		_w994_
	);
	LUT3 #(
		.INIT('h0b)
	) name780 (
		_w345_,
		_w351_,
		_w713_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		_w846_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h4000)
	) name782 (
		_w705_,
		_w844_,
		_w846_,
		_w995_,
		_w997_
	);
	LUT3 #(
		.INIT('h31)
	) name783 (
		_w709_,
		_w715_,
		_w716_,
		_w998_
	);
	LUT3 #(
		.INIT('h4d)
	) name784 (
		_w345_,
		_w351_,
		_w712_,
		_w999_
	);
	LUT3 #(
		.INIT('hd0)
	) name785 (
		_w995_,
		_w998_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		_w698_,
		_w681_,
		_w1001_
	);
	LUT4 #(
		.INIT('h0b02)
	) name787 (
		_w328_,
		_w333_,
		_w718_,
		_w681_,
		_w1002_
	);
	LUT4 #(
		.INIT('h2223)
	) name788 (
		_w705_,
		_w706_,
		_w719_,
		_w1002_,
		_w1003_
	);
	LUT3 #(
		.INIT('hd0)
	) name789 (
		_w994_,
		_w1000_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('h9a55)
	) name790 (
		_w729_,
		_w993_,
		_w997_,
		_w1004_,
		_w1005_
	);
	LUT4 #(
		.INIT('h08c8)
	) name791 (
		\reg2_reg[29]/NET0131 ,
		_w858_,
		_w925_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w509_,
		_w519_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w534_,
		_w499_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0001)
	) name794 (
		_w534_,
		_w499_,
		_w509_,
		_w519_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w613_,
		_w555_,
		_w1010_
	);
	LUT4 #(
		.INIT('h0b02)
	) name796 (
		_w587_,
		_w590_,
		_w601_,
		_w598_,
		_w1011_
	);
	LUT3 #(
		.INIT('h01)
	) name797 (
		_w564_,
		_w575_,
		_w583_,
		_w1012_
	);
	LUT3 #(
		.INIT('h54)
	) name798 (
		_w564_,
		_w600_,
		_w605_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w546_,
		_w567_,
		_w1014_
	);
	LUT4 #(
		.INIT('hf400)
	) name800 (
		_w1011_,
		_w1012_,
		_w1013_,
		_w1014_,
		_w1015_
	);
	LUT3 #(
		.INIT('h80)
	) name801 (
		_w1009_,
		_w1010_,
		_w1015_,
		_w1016_
	);
	LUT3 #(
		.INIT('h54)
	) name802 (
		_w546_,
		_w604_,
		_w607_,
		_w1017_
	);
	LUT3 #(
		.INIT('h54)
	) name803 (
		_w613_,
		_w528_,
		_w608_,
		_w1018_
	);
	LUT3 #(
		.INIT('h07)
	) name804 (
		_w1010_,
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('haa80)
	) name805 (
		_w1009_,
		_w1010_,
		_w1017_,
		_w1018_,
		_w1020_
	);
	LUT3 #(
		.INIT('h54)
	) name806 (
		_w509_,
		_w518_,
		_w531_,
		_w1021_
	);
	LUT3 #(
		.INIT('h32)
	) name807 (
		_w485_,
		_w534_,
		_w530_,
		_w1022_
	);
	LUT3 #(
		.INIT('h07)
	) name808 (
		_w1008_,
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		_w1020_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w424_,
		_w444_,
		_w1025_
	);
	LUT4 #(
		.INIT('h0001)
	) name811 (
		_w413_,
		_w424_,
		_w444_,
		_w450_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w463_,
		_w475_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w471_,
		_w618_,
		_w1028_
	);
	LUT4 #(
		.INIT('h0001)
	) name814 (
		_w463_,
		_w471_,
		_w475_,
		_w618_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		_w1026_,
		_w1029_,
		_w1030_
	);
	LUT3 #(
		.INIT('h54)
	) name816 (
		_w463_,
		_w476_,
		_w487_,
		_w1031_
	);
	LUT3 #(
		.INIT('h31)
	) name817 (
		_w488_,
		_w443_,
		_w618_,
		_w1032_
	);
	LUT3 #(
		.INIT('h70)
	) name818 (
		_w1028_,
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h80aa)
	) name819 (
		_w1026_,
		_w1028_,
		_w1031_,
		_w1032_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w446_,
		_w396_,
		_w1035_
	);
	LUT3 #(
		.INIT('h0e)
	) name821 (
		_w447_,
		_w434_,
		_w424_,
		_w1036_
	);
	LUT4 #(
		.INIT('h0071)
	) name822 (
		_w417_,
		_w422_,
		_w434_,
		_w413_,
		_w1037_
	);
	LUT3 #(
		.INIT('h51)
	) name823 (
		_w450_,
		_w1035_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1034_,
		_w1038_,
		_w1039_
	);
	LUT4 #(
		.INIT('h4f00)
	) name825 (
		_w1016_,
		_w1024_,
		_w1030_,
		_w1039_,
		_w1040_
	);
	LUT3 #(
		.INIT('h07)
	) name826 (
		_w345_,
		_w351_,
		_w379_,
		_w1041_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w658_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h4000)
	) name828 (
		_w318_,
		_w658_,
		_w361_,
		_w1041_,
		_w1043_
	);
	LUT3 #(
		.INIT('h51)
	) name829 (
		_w401_,
		_w388_,
		_w371_,
		_w1044_
	);
	LUT3 #(
		.INIT('h8e)
	) name830 (
		_w345_,
		_w351_,
		_w400_,
		_w1045_
	);
	LUT3 #(
		.INIT('hd0)
	) name831 (
		_w1041_,
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT4 #(
		.INIT('h08aa)
	) name832 (
		_w361_,
		_w1041_,
		_w1044_,
		_w1045_,
		_w1047_
	);
	LUT3 #(
		.INIT('h2b)
	) name833 (
		_w344_,
		_w328_,
		_w333_,
		_w1048_
	);
	LUT4 #(
		.INIT('h000e)
	) name834 (
		_w344_,
		_w356_,
		_w327_,
		_w335_,
		_w1049_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		_w666_,
		_w1049_,
		_w1050_
	);
	LUT3 #(
		.INIT('h45)
	) name836 (
		_w318_,
		_w1047_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('h559a)
	) name837 (
		_w729_,
		_w1040_,
		_w1043_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('hc808)
	) name838 (
		\reg2_reg[29]/NET0131 ,
		_w791_,
		_w925_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name839 (
		_w918_,
		_w1006_,
		_w1053_,
		_w961_,
		_w1054_
	);
	LUT4 #(
		.INIT('heeec)
	) name840 (
		\state_reg[0]/NET0131 ,
		_w945_,
		_w946_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		\reg0_reg[28]/NET0131 ,
		_w942_,
		_w1056_
	);
	LUT3 #(
		.INIT('h0e)
	) name842 (
		_w772_,
		_w778_,
		_w780_,
		_w1057_
	);
	LUT4 #(
		.INIT('hc355)
	) name843 (
		\reg0_reg[28]/NET0131 ,
		_w707_,
		_w789_,
		_w1057_,
		_w1058_
	);
	LUT4 #(
		.INIT('h30a0)
	) name844 (
		\reg0_reg[28]/NET0131 ,
		_w857_,
		_w858_,
		_w1057_,
		_w1059_
	);
	LUT4 #(
		.INIT('h6500)
	) name845 (
		_w310_,
		_w320_,
		_w876_,
		_w878_,
		_w1060_
	);
	LUT4 #(
		.INIT('h0007)
	) name846 (
		_w903_,
		_w904_,
		_w935_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('hf100)
	) name847 (
		_w772_,
		_w778_,
		_w780_,
		_w904_,
		_w1062_
	);
	LUT4 #(
		.INIT('h7f5e)
	) name848 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w1063_
	);
	LUT4 #(
		.INIT('hfafb)
	) name849 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w1064_
	);
	LUT4 #(
		.INIT('h00f1)
	) name850 (
		_w772_,
		_w778_,
		_w780_,
		_w1064_,
		_w1065_
	);
	LUT3 #(
		.INIT('h04)
	) name851 (
		_w1062_,
		_w1063_,
		_w1065_,
		_w1066_
	);
	LUT4 #(
		.INIT('haa8a)
	) name852 (
		\reg0_reg[28]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w1067_
	);
	LUT3 #(
		.INIT('h0d)
	) name853 (
		_w1057_,
		_w1061_,
		_w1067_,
		_w1068_
	);
	LUT4 #(
		.INIT('h0d00)
	) name854 (
		_w791_,
		_w1058_,
		_w1059_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		\reg0_reg[28]/NET0131 ,
		_w919_,
		_w1070_
	);
	LUT4 #(
		.INIT('haa08)
	) name856 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1069_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('he)
	) name857 (
		_w1056_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		\reg1_reg[28]/NET0131 ,
		_w942_,
		_w1073_
	);
	LUT3 #(
		.INIT('h01)
	) name859 (
		_w772_,
		_w778_,
		_w780_,
		_w1074_
	);
	LUT4 #(
		.INIT('hc355)
	) name860 (
		\reg1_reg[28]/NET0131 ,
		_w707_,
		_w789_,
		_w1074_,
		_w1075_
	);
	LUT4 #(
		.INIT('h30a0)
	) name861 (
		\reg1_reg[28]/NET0131 ,
		_w857_,
		_w858_,
		_w1074_,
		_w1076_
	);
	LUT4 #(
		.INIT('hfe00)
	) name862 (
		_w772_,
		_w778_,
		_w780_,
		_w904_,
		_w1077_
	);
	LUT4 #(
		.INIT('h00fe)
	) name863 (
		_w772_,
		_w778_,
		_w780_,
		_w1064_,
		_w1078_
	);
	LUT4 #(
		.INIT('haaa2)
	) name864 (
		\reg1_reg[28]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w1079_
	);
	LUT3 #(
		.INIT('h0b)
	) name865 (
		_w1061_,
		_w1074_,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('h0d00)
	) name866 (
		_w791_,
		_w1075_,
		_w1076_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		\reg1_reg[28]/NET0131 ,
		_w919_,
		_w1082_
	);
	LUT4 #(
		.INIT('haa08)
	) name868 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1081_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('he)
	) name869 (
		_w1073_,
		_w1083_,
		_w1084_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name870 (
		_w464_,
		_w772_,
		_w778_,
		_w780_,
		_w1085_
	);
	LUT3 #(
		.INIT('h07)
	) name871 (
		_w1022_,
		_w1027_,
		_w1031_,
		_w1086_
	);
	LUT4 #(
		.INIT('h0001)
	) name872 (
		_w463_,
		_w475_,
		_w534_,
		_w499_,
		_w1087_
	);
	LUT4 #(
		.INIT('h0001)
	) name873 (
		_w509_,
		_w519_,
		_w613_,
		_w555_,
		_w1088_
	);
	LUT3 #(
		.INIT('h07)
	) name874 (
		_w1007_,
		_w1018_,
		_w1021_,
		_w1089_
	);
	LUT4 #(
		.INIT('h1f00)
	) name875 (
		_w1015_,
		_w1017_,
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT4 #(
		.INIT('h66a6)
	) name876 (
		_w746_,
		_w1086_,
		_w1087_,
		_w1090_,
		_w1091_
	);
	LUT4 #(
		.INIT('he020)
	) name877 (
		_w464_,
		_w781_,
		_w791_,
		_w1091_,
		_w1092_
	);
	LUT4 #(
		.INIT('h0001)
	) name878 (
		_w731_,
		_w737_,
		_w753_,
		_w805_,
		_w1093_
	);
	LUT3 #(
		.INIT('h8a)
	) name879 (
		_w969_,
		_w978_,
		_w981_,
		_w1094_
	);
	LUT4 #(
		.INIT('h4f00)
	) name880 (
		_w976_,
		_w977_,
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h0001)
	) name881 (
		_w692_,
		_w792_,
		_w794_,
		_w802_,
		_w1096_
	);
	LUT3 #(
		.INIT('hd0)
	) name882 (
		_w962_,
		_w970_,
		_w984_,
		_w1097_
	);
	LUT4 #(
		.INIT('h65aa)
	) name883 (
		_w746_,
		_w1095_,
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h20e0)
	) name884 (
		_w464_,
		_w781_,
		_w858_,
		_w1098_,
		_w1099_
	);
	LUT4 #(
		.INIT('h1444)
	) name885 (
		_w277_,
		_w441_,
		_w887_,
		_w889_,
		_w1100_
	);
	LUT4 #(
		.INIT('h0200)
	) name886 (
		_w277_,
		_w456_,
		_w457_,
		_w458_,
		_w1101_
	);
	LUT4 #(
		.INIT('h3331)
	) name887 (
		_w781_,
		_w1085_,
		_w1100_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('h8000)
	) name888 (
		_w462_,
		_w863_,
		_w864_,
		_w865_,
		_w1103_
	);
	LUT4 #(
		.INIT('h070b)
	) name889 (
		_w470_,
		_w781_,
		_w1085_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('ha8)
	) name890 (
		_w470_,
		_w906_,
		_w907_,
		_w1105_
	);
	LUT3 #(
		.INIT('ha8)
	) name891 (
		_w464_,
		_w909_,
		_w910_,
		_w1106_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1105_,
		_w1106_,
		_w1107_
	);
	LUT3 #(
		.INIT('hd0)
	) name893 (
		_w878_,
		_w1104_,
		_w1107_,
		_w1108_
	);
	LUT3 #(
		.INIT('hd0)
	) name894 (
		_w904_,
		_w1102_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1110_
	);
	LUT4 #(
		.INIT('hef00)
	) name896 (
		_w1092_,
		_w1099_,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT4 #(
		.INIT('hdd1d)
	) name897 (
		\reg3_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w464_,
		_w918_,
		_w1112_
	);
	LUT2 #(
		.INIT('hb)
	) name898 (
		_w1111_,
		_w1112_,
		_w1113_
	);
	LUT4 #(
		.INIT('h02aa)
	) name899 (
		\reg2_reg[27]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1114_
	);
	LUT3 #(
		.INIT('hd0)
	) name900 (
		_w847_,
		_w988_,
		_w998_,
		_w1115_
	);
	LUT4 #(
		.INIT('h20f0)
	) name901 (
		_w847_,
		_w988_,
		_w995_,
		_w998_,
		_w1116_
	);
	LUT4 #(
		.INIT('h88c8)
	) name902 (
		_w680_,
		_w1001_,
		_w999_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w699_,
		_w1117_,
		_w1118_
	);
	LUT4 #(
		.INIT('h0001)
	) name904 (
		_w726_,
		_w749_,
		_w744_,
		_w688_,
		_w1119_
	);
	LUT4 #(
		.INIT('h4f00)
	) name905 (
		_w1095_,
		_w1096_,
		_w1097_,
		_w1119_,
		_w1120_
	);
	LUT3 #(
		.INIT('h70)
	) name906 (
		_w965_,
		_w985_,
		_w989_,
		_w1121_
	);
	LUT4 #(
		.INIT('h000b)
	) name907 (
		_w345_,
		_w351_,
		_w713_,
		_w680_,
		_w1122_
	);
	LUT4 #(
		.INIT('h0001)
	) name908 (
		_w710_,
		_w716_,
		_w685_,
		_w798_,
		_w1123_
	);
	LUT3 #(
		.INIT('h40)
	) name909 (
		_w699_,
		_w1123_,
		_w1122_,
		_w1124_
	);
	LUT4 #(
		.INIT('h1055)
	) name910 (
		_w1118_,
		_w1120_,
		_w1121_,
		_w1124_,
		_w1125_
	);
	LUT4 #(
		.INIT('h35c5)
	) name911 (
		\reg2_reg[27]/NET0131 ,
		_w720_,
		_w925_,
		_w1125_,
		_w1126_
	);
	LUT4 #(
		.INIT('h0001)
	) name912 (
		_w471_,
		_w424_,
		_w444_,
		_w618_,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w1087_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('hf800)
	) name914 (
		_w1022_,
		_w1027_,
		_w1031_,
		_w1127_,
		_w1129_
	);
	LUT3 #(
		.INIT('h0d)
	) name915 (
		_w1025_,
		_w1032_,
		_w1036_,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name916 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT4 #(
		.INIT('h0001)
	) name917 (
		_w343_,
		_w335_,
		_w413_,
		_w450_,
		_w1132_
	);
	LUT3 #(
		.INIT('h80)
	) name918 (
		_w658_,
		_w1041_,
		_w1132_,
		_w1133_
	);
	LUT4 #(
		.INIT('h4f00)
	) name919 (
		_w1090_,
		_w1128_,
		_w1131_,
		_w1133_,
		_w1134_
	);
	LUT3 #(
		.INIT('hd0)
	) name920 (
		_w659_,
		_w1035_,
		_w1044_,
		_w1135_
	);
	LUT4 #(
		.INIT('h20f0)
	) name921 (
		_w659_,
		_w1035_,
		_w1041_,
		_w1044_,
		_w1136_
	);
	LUT4 #(
		.INIT('h050d)
	) name922 (
		_w360_,
		_w1045_,
		_w1048_,
		_w1136_,
		_w1137_
	);
	LUT4 #(
		.INIT('h8488)
	) name923 (
		_w720_,
		_w925_,
		_w1134_,
		_w1137_,
		_w1138_
	);
	LUT3 #(
		.INIT('ha8)
	) name924 (
		_w791_,
		_w1114_,
		_w1138_,
		_w1139_
	);
	LUT4 #(
		.INIT('h8000)
	) name925 (
		_w887_,
		_w889_,
		_w892_,
		_w897_,
		_w1140_
	);
	LUT4 #(
		.INIT('h0d05)
	) name926 (
		_w315_,
		_w898_,
		_w901_,
		_w1140_,
		_w1141_
	);
	LUT4 #(
		.INIT('h7020)
	) name927 (
		_w277_,
		_w333_,
		_w925_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h3c55)
	) name928 (
		\reg2_reg[27]/NET0131 ,
		_w320_,
		_w876_,
		_w925_,
		_w1143_
	);
	LUT3 #(
		.INIT('ha8)
	) name929 (
		\reg2_reg[27]/NET0131 ,
		_w909_,
		_w932_,
		_w1144_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w321_,
		_w907_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		_w320_,
		_w905_,
		_w1146_
	);
	LUT3 #(
		.INIT('h13)
	) name932 (
		_w925_,
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		_w1144_,
		_w1147_,
		_w1148_
	);
	LUT3 #(
		.INIT('hd0)
	) name934 (
		_w878_,
		_w1143_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h5700)
	) name935 (
		_w904_,
		_w1114_,
		_w1142_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h0d00)
	) name936 (
		_w858_,
		_w1126_,
		_w1139_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		\reg2_reg[27]/NET0131 ,
		_w919_,
		_w1152_
	);
	LUT4 #(
		.INIT('haa08)
	) name938 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\reg2_reg[27]/NET0131 ,
		_w942_,
		_w1154_
	);
	LUT2 #(
		.INIT('he)
	) name940 (
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		\reg0_reg[27]/NET0131 ,
		_w942_,
		_w1156_
	);
	LUT4 #(
		.INIT('haa02)
	) name942 (
		\reg0_reg[27]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1157_
	);
	LUT4 #(
		.INIT('h35c5)
	) name943 (
		\reg0_reg[27]/NET0131 ,
		_w720_,
		_w1057_,
		_w1125_,
		_w1158_
	);
	LUT4 #(
		.INIT('h8488)
	) name944 (
		_w720_,
		_w1057_,
		_w1134_,
		_w1137_,
		_w1159_
	);
	LUT3 #(
		.INIT('ha8)
	) name945 (
		_w791_,
		_w1157_,
		_w1159_,
		_w1160_
	);
	LUT4 #(
		.INIT('h7020)
	) name946 (
		_w277_,
		_w333_,
		_w904_,
		_w1141_,
		_w1161_
	);
	LUT4 #(
		.INIT('h006f)
	) name947 (
		_w320_,
		_w876_,
		_w878_,
		_w1146_,
		_w1162_
	);
	LUT4 #(
		.INIT('haa8a)
	) name948 (
		\reg0_reg[27]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w1163_
	);
	LUT4 #(
		.INIT('h0075)
	) name949 (
		_w1057_,
		_w1161_,
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('h0d00)
	) name950 (
		_w858_,
		_w1158_,
		_w1160_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		\reg0_reg[27]/NET0131 ,
		_w919_,
		_w1166_
	);
	LUT4 #(
		.INIT('haa08)
	) name952 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1165_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('he)
	) name953 (
		_w1156_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\reg0_reg[29]/NET0131 ,
		_w942_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		\reg0_reg[29]/NET0131 ,
		_w919_,
		_w1170_
	);
	LUT4 #(
		.INIT('hf800)
	) name956 (
		_w878_,
		_w948_,
		_w958_,
		_w1057_,
		_w1171_
	);
	LUT4 #(
		.INIT('h0355)
	) name957 (
		\reg0_reg[29]/NET0131 ,
		_w950_,
		_w954_,
		_w1057_,
		_w1172_
	);
	LUT3 #(
		.INIT('ha2)
	) name958 (
		\reg0_reg[29]/NET0131 ,
		_w1063_,
		_w1065_,
		_w1173_
	);
	LUT4 #(
		.INIT('h0031)
	) name959 (
		_w904_,
		_w1171_,
		_w1172_,
		_w1173_,
		_w1174_
	);
	LUT4 #(
		.INIT('h0c88)
	) name960 (
		\reg0_reg[29]/NET0131 ,
		_w858_,
		_w1005_,
		_w1057_,
		_w1175_
	);
	LUT4 #(
		.INIT('hc088)
	) name961 (
		\reg0_reg[29]/NET0131 ,
		_w791_,
		_w1052_,
		_w1057_,
		_w1176_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name962 (
		_w918_,
		_w1175_,
		_w1176_,
		_w1174_,
		_w1177_
	);
	LUT4 #(
		.INIT('heeec)
	) name963 (
		\state_reg[0]/NET0131 ,
		_w1169_,
		_w1170_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h2)
	) name964 (
		\reg1_reg[27]/NET0131 ,
		_w942_,
		_w1179_
	);
	LUT4 #(
		.INIT('haaa8)
	) name965 (
		\reg1_reg[27]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1180_
	);
	LUT4 #(
		.INIT('h35c5)
	) name966 (
		\reg1_reg[27]/NET0131 ,
		_w720_,
		_w1074_,
		_w1125_,
		_w1181_
	);
	LUT4 #(
		.INIT('h8488)
	) name967 (
		_w720_,
		_w1074_,
		_w1134_,
		_w1137_,
		_w1182_
	);
	LUT3 #(
		.INIT('ha8)
	) name968 (
		_w791_,
		_w1180_,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('haaa2)
	) name969 (
		\reg1_reg[27]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w1184_
	);
	LUT4 #(
		.INIT('h0075)
	) name970 (
		_w1074_,
		_w1161_,
		_w1162_,
		_w1184_,
		_w1185_
	);
	LUT4 #(
		.INIT('h0d00)
	) name971 (
		_w858_,
		_w1181_,
		_w1183_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		\reg1_reg[27]/NET0131 ,
		_w919_,
		_w1187_
	);
	LUT4 #(
		.INIT('haa08)
	) name973 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('he)
	) name974 (
		_w1179_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		\reg1_reg[29]/NET0131 ,
		_w942_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name976 (
		\reg1_reg[29]/NET0131 ,
		_w919_,
		_w1191_
	);
	LUT4 #(
		.INIT('hf800)
	) name977 (
		_w878_,
		_w948_,
		_w958_,
		_w1074_,
		_w1192_
	);
	LUT4 #(
		.INIT('h0355)
	) name978 (
		\reg1_reg[29]/NET0131 ,
		_w950_,
		_w954_,
		_w1074_,
		_w1193_
	);
	LUT3 #(
		.INIT('ha2)
	) name979 (
		\reg1_reg[29]/NET0131 ,
		_w1063_,
		_w1078_,
		_w1194_
	);
	LUT4 #(
		.INIT('h0031)
	) name980 (
		_w904_,
		_w1192_,
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT4 #(
		.INIT('h0c88)
	) name981 (
		\reg1_reg[29]/NET0131 ,
		_w858_,
		_w1005_,
		_w1074_,
		_w1196_
	);
	LUT4 #(
		.INIT('hc088)
	) name982 (
		\reg1_reg[29]/NET0131 ,
		_w791_,
		_w1052_,
		_w1074_,
		_w1197_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name983 (
		_w918_,
		_w1196_,
		_w1197_,
		_w1195_,
		_w1198_
	);
	LUT4 #(
		.INIT('heeec)
	) name984 (
		\state_reg[0]/NET0131 ,
		_w1190_,
		_w1191_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		_w494_,
		_w919_,
		_w1200_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name986 (
		_w494_,
		_w772_,
		_w778_,
		_w780_,
		_w1201_
	);
	LUT4 #(
		.INIT('h007b)
	) name987 (
		_w722_,
		_w781_,
		_w1090_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		_w791_,
		_w1202_,
		_w1203_
	);
	LUT3 #(
		.INIT('h80)
	) name989 (
		_w277_,
		_w501_,
		_w502_,
		_w1204_
	);
	LUT4 #(
		.INIT('h00eb)
	) name990 (
		_w277_,
		_w480_,
		_w887_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('he020)
	) name991 (
		_w494_,
		_w781_,
		_w904_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h00b7)
	) name992 (
		_w722_,
		_w781_,
		_w1095_,
		_w1201_,
		_w1207_
	);
	LUT4 #(
		.INIT('h2000)
	) name993 (
		_w493_,
		_w508_,
		_w863_,
		_w864_,
		_w1208_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name994 (
		_w493_,
		_w508_,
		_w863_,
		_w864_,
		_w1209_
	);
	LUT4 #(
		.INIT('he020)
	) name995 (
		_w494_,
		_w781_,
		_w878_,
		_w1209_,
		_w1210_
	);
	LUT3 #(
		.INIT('h54)
	) name996 (
		_w493_,
		_w906_,
		_w907_,
		_w1211_
	);
	LUT3 #(
		.INIT('ha8)
	) name997 (
		_w494_,
		_w909_,
		_w910_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w1211_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name999 (
		_w1210_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1000 (
		_w858_,
		_w1207_,
		_w1206_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('h1311)
	) name1001 (
		_w918_,
		_w1200_,
		_w1203_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		\reg3_reg[11]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1217_
	);
	LUT3 #(
		.INIT('h07)
	) name1003 (
		_w269_,
		_w494_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('h2f)
	) name1004 (
		\state_reg[0]/NET0131 ,
		_w1216_,
		_w1218_,
		_w1219_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w478_,
		_w919_,
		_w1220_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1006 (
		_w478_,
		_w772_,
		_w778_,
		_w780_,
		_w1221_
	);
	LUT4 #(
		.INIT('h758a)
	) name1007 (
		_w533_,
		_w610_,
		_w639_,
		_w694_,
		_w1222_
	);
	LUT4 #(
		.INIT('he020)
	) name1008 (
		_w478_,
		_w781_,
		_w791_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('h4484)
	) name1009 (
		_w694_,
		_w781_,
		_w809_,
		_w830_,
		_w1224_
	);
	LUT3 #(
		.INIT('ha8)
	) name1010 (
		_w858_,
		_w1221_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('h2122)
	) name1011 (
		_w260_,
		_w277_,
		_w480_,
		_w887_,
		_w1226_
	);
	LUT3 #(
		.INIT('h80)
	) name1012 (
		_w277_,
		_w495_,
		_w496_,
		_w1227_
	);
	LUT4 #(
		.INIT('h3331)
	) name1013 (
		_w781_,
		_w1221_,
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('h007b)
	) name1014 (
		_w484_,
		_w781_,
		_w1208_,
		_w1221_,
		_w1229_
	);
	LUT3 #(
		.INIT('ha8)
	) name1015 (
		_w484_,
		_w906_,
		_w907_,
		_w1230_
	);
	LUT3 #(
		.INIT('ha8)
	) name1016 (
		_w478_,
		_w909_,
		_w910_,
		_w1231_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1230_,
		_w1231_,
		_w1232_
	);
	LUT3 #(
		.INIT('hd0)
	) name1018 (
		_w878_,
		_w1229_,
		_w1232_,
		_w1233_
	);
	LUT3 #(
		.INIT('hd0)
	) name1019 (
		_w904_,
		_w1228_,
		_w1233_,
		_w1234_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1020 (
		_w918_,
		_w1223_,
		_w1225_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h2)
	) name1021 (
		\reg3_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1236_
	);
	LUT3 #(
		.INIT('h07)
	) name1022 (
		_w269_,
		_w478_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1023 (
		\state_reg[0]/NET0131 ,
		_w1220_,
		_w1235_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h8)
	) name1024 (
		_w348_,
		_w919_,
		_w1239_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1025 (
		_w348_,
		_w772_,
		_w778_,
		_w780_,
		_w1240_
	);
	LUT4 #(
		.INIT('h0800)
	) name1026 (
		_w621_,
		_w536_,
		_w610_,
		_w639_,
		_w1241_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1027 (
		_w491_,
		_w449_,
		_w620_,
		_w537_,
		_w1242_
	);
	LUT3 #(
		.INIT('ha2)
	) name1028 (
		_w404_,
		_w452_,
		_w1242_,
		_w1243_
	);
	LUT4 #(
		.INIT('h8488)
	) name1029 (
		_w704_,
		_w781_,
		_w1241_,
		_w1243_,
		_w1244_
	);
	LUT3 #(
		.INIT('ha8)
	) name1030 (
		_w791_,
		_w1240_,
		_w1244_,
		_w1245_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1031 (
		_w277_,
		_w375_,
		_w374_,
		_w376_,
		_w1246_
	);
	LUT4 #(
		.INIT('h8000)
	) name1032 (
		_w887_,
		_w889_,
		_w892_,
		_w895_,
		_w1247_
	);
	LUT3 #(
		.INIT('h8a)
	) name1033 (
		_w341_,
		_w351_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w277_,
		_w1140_,
		_w1249_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1035 (
		_w781_,
		_w1246_,
		_w1248_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('ha8)
	) name1036 (
		_w345_,
		_w906_,
		_w907_,
		_w1251_
	);
	LUT3 #(
		.INIT('ha8)
	) name1037 (
		_w348_,
		_w909_,
		_w910_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h5700)
	) name1039 (
		_w904_,
		_w1240_,
		_w1250_,
		_w1253_,
		_w1254_
	);
	LUT3 #(
		.INIT('h40)
	) name1040 (
		_w381_,
		_w869_,
		_w870_,
		_w1255_
	);
	LUT4 #(
		.INIT('h1000)
	) name1041 (
		_w363_,
		_w381_,
		_w869_,
		_w870_,
		_w1256_
	);
	LUT4 #(
		.INIT('h0705)
	) name1042 (
		_w345_,
		_w372_,
		_w874_,
		_w1256_,
		_w1257_
	);
	LUT4 #(
		.INIT('he020)
	) name1043 (
		_w348_,
		_w781_,
		_w878_,
		_w1257_,
		_w1258_
	);
	LUT4 #(
		.INIT('haa08)
	) name1044 (
		_w796_,
		_w803_,
		_w806_,
		_w808_,
		_w1259_
	);
	LUT4 #(
		.INIT('h50d0)
	) name1045 (
		_w800_,
		_w835_,
		_w840_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h80f0)
	) name1046 (
		_w801_,
		_w830_,
		_w848_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('h4448)
	) name1047 (
		_w704_,
		_w781_,
		_w853_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h0507)
	) name1048 (
		_w858_,
		_w1240_,
		_w1258_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1049 (
		_w918_,
		_w1245_,
		_w1254_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\reg3_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1265_
	);
	LUT3 #(
		.INIT('h07)
	) name1051 (
		_w269_,
		_w348_,
		_w1265_,
		_w1266_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1052 (
		\state_reg[0]/NET0131 ,
		_w1239_,
		_w1264_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		_w373_,
		_w919_,
		_w1268_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1054 (
		_w373_,
		_w772_,
		_w778_,
		_w780_,
		_w1269_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1055 (
		_w1115_,
		_w1120_,
		_w1121_,
		_w1123_,
		_w1270_
	);
	LUT4 #(
		.INIT('h070b)
	) name1056 (
		_w714_,
		_w781_,
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT4 #(
		.INIT('h0001)
	) name1057 (
		_w371_,
		_w398_,
		_w413_,
		_w450_,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		_w1127_,
		_w1272_,
		_w1273_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1059 (
		_w1086_,
		_w1087_,
		_w1090_,
		_w1273_,
		_w1274_
	);
	LUT4 #(
		.INIT('hf200)
	) name1060 (
		_w1025_,
		_w1032_,
		_w1036_,
		_w1272_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		_w1135_,
		_w1275_,
		_w1276_
	);
	LUT4 #(
		.INIT('h8488)
	) name1062 (
		_w714_,
		_w781_,
		_w1274_,
		_w1276_,
		_w1277_
	);
	LUT3 #(
		.INIT('ha8)
	) name1063 (
		_w791_,
		_w1269_,
		_w1277_,
		_w1278_
	);
	LUT4 #(
		.INIT('h007b)
	) name1064 (
		_w372_,
		_w781_,
		_w1256_,
		_w1269_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name1065 (
		_w878_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h0200)
	) name1066 (
		_w277_,
		_w367_,
		_w366_,
		_w368_,
		_w1281_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1067 (
		_w277_,
		_w351_,
		_w1247_,
		_w1281_,
		_w1282_
	);
	LUT4 #(
		.INIT('he020)
	) name1068 (
		_w373_,
		_w781_,
		_w904_,
		_w1282_,
		_w1283_
	);
	LUT3 #(
		.INIT('ha8)
	) name1069 (
		_w373_,
		_w909_,
		_w910_,
		_w1284_
	);
	LUT3 #(
		.INIT('ha8)
	) name1070 (
		_w372_,
		_w906_,
		_w907_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT3 #(
		.INIT('h10)
	) name1072 (
		_w1283_,
		_w1280_,
		_w1286_,
		_w1287_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1073 (
		_w858_,
		_w1271_,
		_w1278_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1074 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1268_,
		_w1288_,
		_w1289_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name1075 (
		\reg3_reg[23]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w268_,
		_w347_,
		_w1290_
	);
	LUT2 #(
		.INIT('hb)
	) name1076 (
		_w1289_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h2)
	) name1077 (
		\reg0_reg[15]/NET0131 ,
		_w942_,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		\reg0_reg[15]/NET0131 ,
		_w919_,
		_w1293_
	);
	LUT4 #(
		.INIT('hc808)
	) name1079 (
		\reg0_reg[15]/NET0131 ,
		_w791_,
		_w1057_,
		_w1091_,
		_w1294_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1080 (
		\reg0_reg[15]/NET0131 ,
		_w858_,
		_w1057_,
		_w1098_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		_w470_,
		_w905_,
		_w1296_
	);
	LUT4 #(
		.INIT('h007b)
	) name1082 (
		_w470_,
		_w878_,
		_w1103_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1083 (
		_w904_,
		_w1100_,
		_w1101_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1084 (
		\reg0_reg[15]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w1299_
	);
	LUT3 #(
		.INIT('h0d)
	) name1085 (
		_w1057_,
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1086 (
		_w918_,
		_w1294_,
		_w1295_,
		_w1300_,
		_w1301_
	);
	LUT4 #(
		.INIT('heeec)
	) name1087 (
		\state_reg[0]/NET0131 ,
		_w1292_,
		_w1293_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		\reg0_reg[23]/NET0131 ,
		_w942_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name1089 (
		\reg0_reg[23]/NET0131 ,
		_w919_,
		_w1304_
	);
	LUT4 #(
		.INIT('haa02)
	) name1090 (
		\reg0_reg[23]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1305_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1091 (
		\reg0_reg[23]/NET0131 ,
		_w714_,
		_w1057_,
		_w1270_,
		_w1306_
	);
	LUT4 #(
		.INIT('h8488)
	) name1092 (
		_w714_,
		_w1057_,
		_w1274_,
		_w1276_,
		_w1307_
	);
	LUT3 #(
		.INIT('ha8)
	) name1093 (
		_w791_,
		_w1305_,
		_w1307_,
		_w1308_
	);
	LUT3 #(
		.INIT('h84)
	) name1094 (
		_w372_,
		_w878_,
		_w1256_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name1095 (
		_w372_,
		_w905_,
		_w1310_
	);
	LUT4 #(
		.INIT('h0007)
	) name1096 (
		_w904_,
		_w1282_,
		_w1310_,
		_w1309_,
		_w1311_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1097 (
		\reg0_reg[23]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w1312_
	);
	LUT3 #(
		.INIT('h0d)
	) name1098 (
		_w1057_,
		_w1311_,
		_w1312_,
		_w1313_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1099 (
		_w858_,
		_w1306_,
		_w1308_,
		_w1313_,
		_w1314_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1100 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1304_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('he)
	) name1101 (
		_w1303_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h2)
	) name1102 (
		\reg0_reg[24]/NET0131 ,
		_w942_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		\reg0_reg[24]/NET0131 ,
		_w919_,
		_w1318_
	);
	LUT4 #(
		.INIT('haa02)
	) name1104 (
		\reg0_reg[24]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1319_
	);
	LUT4 #(
		.INIT('h8488)
	) name1105 (
		_w704_,
		_w1057_,
		_w1241_,
		_w1243_,
		_w1320_
	);
	LUT3 #(
		.INIT('ha8)
	) name1106 (
		_w791_,
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1107 (
		_w1057_,
		_w1246_,
		_w1248_,
		_w1249_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name1108 (
		_w345_,
		_w905_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w1057_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('hf100)
	) name1110 (
		_w772_,
		_w778_,
		_w780_,
		_w905_,
		_w1325_
	);
	LUT3 #(
		.INIT('ha2)
	) name1111 (
		\reg0_reg[24]/NET0131 ,
		_w1063_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('h5700)
	) name1113 (
		_w904_,
		_w1319_,
		_w1322_,
		_w1327_,
		_w1328_
	);
	LUT4 #(
		.INIT('hc808)
	) name1114 (
		\reg0_reg[24]/NET0131 ,
		_w878_,
		_w1057_,
		_w1257_,
		_w1329_
	);
	LUT4 #(
		.INIT('h5060)
	) name1115 (
		_w704_,
		_w853_,
		_w1057_,
		_w1261_,
		_w1330_
	);
	LUT4 #(
		.INIT('h0507)
	) name1116 (
		_w858_,
		_w1319_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1117 (
		_w918_,
		_w1321_,
		_w1328_,
		_w1331_,
		_w1332_
	);
	LUT4 #(
		.INIT('heeec)
	) name1118 (
		\state_reg[0]/NET0131 ,
		_w1317_,
		_w1318_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h2)
	) name1119 (
		\reg1_reg[15]/NET0131 ,
		_w942_,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		\reg1_reg[15]/NET0131 ,
		_w919_,
		_w1335_
	);
	LUT4 #(
		.INIT('hc808)
	) name1121 (
		\reg1_reg[15]/NET0131 ,
		_w791_,
		_w1074_,
		_w1091_,
		_w1336_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1122 (
		\reg1_reg[15]/NET0131 ,
		_w858_,
		_w1074_,
		_w1098_,
		_w1337_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1123 (
		\reg1_reg[15]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w1338_
	);
	LUT3 #(
		.INIT('h0d)
	) name1124 (
		_w1074_,
		_w1298_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1125 (
		_w918_,
		_w1336_,
		_w1337_,
		_w1339_,
		_w1340_
	);
	LUT4 #(
		.INIT('heeec)
	) name1126 (
		\state_reg[0]/NET0131 ,
		_w1334_,
		_w1335_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		\reg1_reg[23]/NET0131 ,
		_w942_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		\reg1_reg[23]/NET0131 ,
		_w919_,
		_w1343_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1129 (
		\reg1_reg[23]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1344_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1130 (
		\reg1_reg[23]/NET0131 ,
		_w714_,
		_w1074_,
		_w1270_,
		_w1345_
	);
	LUT4 #(
		.INIT('h8488)
	) name1131 (
		_w714_,
		_w1074_,
		_w1274_,
		_w1276_,
		_w1346_
	);
	LUT3 #(
		.INIT('ha8)
	) name1132 (
		_w791_,
		_w1344_,
		_w1346_,
		_w1347_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1133 (
		\reg1_reg[23]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w1348_
	);
	LUT3 #(
		.INIT('h0d)
	) name1134 (
		_w1074_,
		_w1311_,
		_w1348_,
		_w1349_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1135 (
		_w858_,
		_w1345_,
		_w1347_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1136 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1343_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('he)
	) name1137 (
		_w1342_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name1138 (
		\reg2_reg[15]/NET0131 ,
		_w942_,
		_w1353_
	);
	LUT2 #(
		.INIT('h8)
	) name1139 (
		\reg2_reg[15]/NET0131 ,
		_w919_,
		_w1354_
	);
	LUT4 #(
		.INIT('hc808)
	) name1140 (
		\reg2_reg[15]/NET0131 ,
		_w791_,
		_w925_,
		_w1091_,
		_w1355_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1141 (
		\reg2_reg[15]/NET0131 ,
		_w858_,
		_w925_,
		_w1098_,
		_w1356_
	);
	LUT4 #(
		.INIT('h0400)
	) name1142 (
		_w268_,
		_w464_,
		_w272_,
		_w645_,
		_w1357_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1143 (
		_w772_,
		_w778_,
		_w780_,
		_w904_,
		_w1358_
	);
	LUT4 #(
		.INIT('h001f)
	) name1144 (
		_w772_,
		_w778_,
		_w780_,
		_w1064_,
		_w1359_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1145 (
		\reg2_reg[15]/NET0131 ,
		_w909_,
		_w1358_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1357_,
		_w1360_,
		_w1361_
	);
	LUT3 #(
		.INIT('hd0)
	) name1147 (
		_w925_,
		_w1298_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1148 (
		_w918_,
		_w1355_,
		_w1356_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('heeec)
	) name1149 (
		\state_reg[0]/NET0131 ,
		_w1353_,
		_w1354_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h2)
	) name1150 (
		\reg2_reg[23]/NET0131 ,
		_w942_,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\reg2_reg[23]/NET0131 ,
		_w919_,
		_w1366_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1152 (
		\reg2_reg[23]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1367_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1153 (
		\reg2_reg[23]/NET0131 ,
		_w714_,
		_w925_,
		_w1270_,
		_w1368_
	);
	LUT4 #(
		.INIT('h8488)
	) name1154 (
		_w714_,
		_w925_,
		_w1274_,
		_w1276_,
		_w1369_
	);
	LUT3 #(
		.INIT('ha8)
	) name1155 (
		_w791_,
		_w1367_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		_w373_,
		_w907_,
		_w1371_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1157 (
		\reg2_reg[23]/NET0131 ,
		_w909_,
		_w1358_,
		_w1359_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT3 #(
		.INIT('hd0)
	) name1159 (
		_w925_,
		_w1311_,
		_w1373_,
		_w1374_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1160 (
		_w858_,
		_w1368_,
		_w1370_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1161 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1366_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('he)
	) name1162 (
		_w1365_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		_w455_,
		_w919_,
		_w1378_
	);
	LUT4 #(
		.INIT('h8088)
	) name1164 (
		_w614_,
		_w556_,
		_w603_,
		_w606_,
		_w1379_
	);
	LUT3 #(
		.INIT('h4c)
	) name1165 (
		_w614_,
		_w529_,
		_w609_,
		_w1380_
	);
	LUT4 #(
		.INIT('h0001)
	) name1166 (
		_w475_,
		_w534_,
		_w499_,
		_w509_,
		_w1381_
	);
	LUT3 #(
		.INIT('h15)
	) name1167 (
		_w486_,
		_w535_,
		_w532_,
		_w1382_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1168 (
		_w1379_,
		_w1380_,
		_w1381_,
		_w1382_,
		_w1383_
	);
	LUT3 #(
		.INIT('h84)
	) name1169 (
		_w697_,
		_w791_,
		_w1383_,
		_w1384_
	);
	LUT3 #(
		.INIT('h70)
	) name1170 (
		_w793_,
		_w808_,
		_w832_,
		_w1385_
	);
	LUT4 #(
		.INIT('h0001)
	) name1171 (
		_w731_,
		_w737_,
		_w805_,
		_w810_,
		_w1386_
	);
	LUT3 #(
		.INIT('h8a)
	) name1172 (
		_w806_,
		_w826_,
		_w828_,
		_w1387_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1173 (
		_w822_,
		_w824_,
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h0001)
	) name1174 (
		_w692_,
		_w753_,
		_w792_,
		_w802_,
		_w1389_
	);
	LUT4 #(
		.INIT('h1511)
	) name1175 (
		_w697_,
		_w1385_,
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT4 #(
		.INIT('h8088)
	) name1176 (
		_w697_,
		_w1385_,
		_w1388_,
		_w1389_,
		_w1391_
	);
	LUT3 #(
		.INIT('h02)
	) name1177 (
		_w858_,
		_w1391_,
		_w1390_,
		_w1392_
	);
	LUT3 #(
		.INIT('h15)
	) name1178 (
		_w277_,
		_w465_,
		_w466_,
		_w1393_
	);
	LUT4 #(
		.INIT('h0100)
	) name1179 (
		_w260_,
		_w459_,
		_w480_,
		_w887_,
		_w1394_
	);
	LUT3 #(
		.INIT('h70)
	) name1180 (
		_w258_,
		_w259_,
		_w277_,
		_w1395_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1181 (
		_w890_,
		_w1393_,
		_w1394_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h1555)
	) name1182 (
		_w462_,
		_w863_,
		_w864_,
		_w865_,
		_w1397_
	);
	LUT3 #(
		.INIT('h02)
	) name1183 (
		_w878_,
		_w1103_,
		_w1397_,
		_w1398_
	);
	LUT3 #(
		.INIT('h0d)
	) name1184 (
		_w904_,
		_w1396_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1185 (
		_w781_,
		_w1392_,
		_w1384_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('h54)
	) name1186 (
		_w462_,
		_w906_,
		_w907_,
		_w1401_
	);
	LUT3 #(
		.INIT('h09)
	) name1187 (
		_w268_,
		_w632_,
		_w762_,
		_w1402_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1188 (
		_w772_,
		_w778_,
		_w780_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1189 (
		_w455_,
		_w909_,
		_w910_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w1401_,
		_w1404_,
		_w1405_
	);
	LUT4 #(
		.INIT('h1311)
	) name1191 (
		_w918_,
		_w1378_,
		_w1400_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		\reg3_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1407_
	);
	LUT3 #(
		.INIT('h07)
	) name1193 (
		_w269_,
		_w455_,
		_w1407_,
		_w1408_
	);
	LUT3 #(
		.INIT('h2f)
	) name1194 (
		\state_reg[0]/NET0131 ,
		_w1406_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		_w438_,
		_w919_,
		_w1410_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1196 (
		_w438_,
		_w772_,
		_w778_,
		_w780_,
		_w1411_
	);
	LUT4 #(
		.INIT('h009f)
	) name1197 (
		_w640_,
		_w751_,
		_w781_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name1198 (
		_w791_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1199 (
		_w796_,
		_w809_,
		_w830_,
		_w835_,
		_w1414_
	);
	LUT4 #(
		.INIT('h070b)
	) name1200 (
		_w751_,
		_w781_,
		_w1411_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('h1000)
	) name1201 (
		_w429_,
		_w441_,
		_w887_,
		_w889_,
		_w1416_
	);
	LUT4 #(
		.INIT('h6555)
	) name1202 (
		_w429_,
		_w441_,
		_w887_,
		_w889_,
		_w1417_
	);
	LUT4 #(
		.INIT('h7020)
	) name1203 (
		_w277_,
		_w467_,
		_w781_,
		_w1417_,
		_w1418_
	);
	LUT3 #(
		.INIT('ha8)
	) name1204 (
		_w904_,
		_w1411_,
		_w1418_,
		_w1419_
	);
	LUT4 #(
		.INIT('h2d0f)
	) name1205 (
		_w462_,
		_w470_,
		_w436_,
		_w866_,
		_w1420_
	);
	LUT4 #(
		.INIT('he020)
	) name1206 (
		_w438_,
		_w781_,
		_w878_,
		_w1420_,
		_w1421_
	);
	LUT3 #(
		.INIT('ha8)
	) name1207 (
		_w436_,
		_w906_,
		_w907_,
		_w1422_
	);
	LUT3 #(
		.INIT('ha8)
	) name1208 (
		_w438_,
		_w909_,
		_w910_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h4)
	) name1210 (
		_w1421_,
		_w1424_,
		_w1425_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1211 (
		_w858_,
		_w1415_,
		_w1419_,
		_w1425_,
		_w1426_
	);
	LUT4 #(
		.INIT('h1311)
	) name1212 (
		_w918_,
		_w1410_,
		_w1413_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\reg3_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1428_
	);
	LUT3 #(
		.INIT('h07)
	) name1214 (
		_w269_,
		_w438_,
		_w1428_,
		_w1429_
	);
	LUT3 #(
		.INIT('h2f)
	) name1215 (
		\state_reg[0]/NET0131 ,
		_w1427_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w548_,
		_w919_,
		_w1431_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1217 (
		_w548_,
		_w772_,
		_w778_,
		_w780_,
		_w1432_
	);
	LUT4 #(
		.INIT('h4000)
	) name1218 (
		_w523_,
		_w881_,
		_w882_,
		_w883_,
		_w1433_
	);
	LUT4 #(
		.INIT('h9555)
	) name1219 (
		_w523_,
		_w881_,
		_w882_,
		_w883_,
		_w1434_
	);
	LUT4 #(
		.INIT('h7020)
	) name1220 (
		_w277_,
		_w544_,
		_w781_,
		_w1434_,
		_w1435_
	);
	LUT3 #(
		.INIT('ha8)
	) name1221 (
		_w904_,
		_w1432_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('h8884)
	) name1222 (
		_w733_,
		_w781_,
		_w1015_,
		_w1017_,
		_w1437_
	);
	LUT3 #(
		.INIT('ha8)
	) name1223 (
		_w791_,
		_w1432_,
		_w1437_,
		_w1438_
	);
	LUT4 #(
		.INIT('h4844)
	) name1224 (
		_w733_,
		_w781_,
		_w976_,
		_w977_,
		_w1439_
	);
	LUT4 #(
		.INIT('h9300)
	) name1225 (
		_w540_,
		_w554_,
		_w861_,
		_w878_,
		_w1440_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1226 (
		_w772_,
		_w778_,
		_w780_,
		_w1064_,
		_w1441_
	);
	LUT3 #(
		.INIT('ha8)
	) name1227 (
		_w548_,
		_w909_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('ha8)
	) name1228 (
		_w554_,
		_w906_,
		_w907_,
		_w1443_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1442_,
		_w1443_,
		_w1444_
	);
	LUT3 #(
		.INIT('h70)
	) name1230 (
		_w781_,
		_w1440_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('h5700)
	) name1231 (
		_w858_,
		_w1432_,
		_w1439_,
		_w1445_,
		_w1446_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1232 (
		_w918_,
		_w1438_,
		_w1436_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name1233 (
		\reg3_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1448_
	);
	LUT3 #(
		.INIT('h07)
	) name1234 (
		_w269_,
		_w548_,
		_w1448_,
		_w1449_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1235 (
		\state_reg[0]/NET0131 ,
		_w1431_,
		_w1447_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\reg3_reg[19]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1451_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1237 (
		_w407_,
		_w772_,
		_w778_,
		_w780_,
		_w1452_
	);
	LUT4 #(
		.INIT('h8488)
	) name1238 (
		_w683_,
		_w781_,
		_w1120_,
		_w1121_,
		_w1453_
	);
	LUT3 #(
		.INIT('ha8)
	) name1239 (
		_w858_,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h65aa)
	) name1240 (
		_w683_,
		_w1090_,
		_w1128_,
		_w1131_,
		_w1455_
	);
	LUT4 #(
		.INIT('h20e0)
	) name1241 (
		_w407_,
		_w781_,
		_w791_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h4000)
	) name1242 (
		_w394_,
		_w887_,
		_w889_,
		_w892_,
		_w1457_
	);
	LUT4 #(
		.INIT('h9555)
	) name1243 (
		_w394_,
		_w887_,
		_w889_,
		_w892_,
		_w1458_
	);
	LUT4 #(
		.INIT('h7020)
	) name1244 (
		_w277_,
		_w422_,
		_w781_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h90a0)
	) name1245 (
		_w406_,
		_w417_,
		_w781_,
		_w869_,
		_w1460_
	);
	LUT3 #(
		.INIT('h54)
	) name1246 (
		_w406_,
		_w906_,
		_w907_,
		_w1461_
	);
	LUT4 #(
		.INIT('h5700)
	) name1247 (
		_w407_,
		_w909_,
		_w910_,
		_w918_,
		_w1462_
	);
	LUT2 #(
		.INIT('h4)
	) name1248 (
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h5700)
	) name1249 (
		_w878_,
		_w1452_,
		_w1460_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('h5700)
	) name1250 (
		_w904_,
		_w1452_,
		_w1459_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name1251 (
		_w1456_,
		_w1465_,
		_w1466_
	);
	LUT3 #(
		.INIT('ha8)
	) name1252 (
		\state_reg[0]/NET0131 ,
		_w407_,
		_w918_,
		_w1467_
	);
	LUT4 #(
		.INIT('hefaa)
	) name1253 (
		_w1451_,
		_w1454_,
		_w1466_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		_w390_,
		_w919_,
		_w1469_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1255 (
		_w390_,
		_w772_,
		_w778_,
		_w780_,
		_w1470_
	);
	LUT4 #(
		.INIT('h8488)
	) name1256 (
		_w686_,
		_w781_,
		_w784_,
		_w786_,
		_w1471_
	);
	LUT3 #(
		.INIT('ha8)
	) name1257 (
		_w791_,
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT4 #(
		.INIT('h007b)
	) name1258 (
		_w686_,
		_w781_,
		_w842_,
		_w1470_,
		_w1473_
	);
	LUT4 #(
		.INIT('h0200)
	) name1259 (
		_w277_,
		_w409_,
		_w408_,
		_w410_,
		_w1474_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1260 (
		_w277_,
		_w386_,
		_w1457_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('he020)
	) name1261 (
		_w390_,
		_w781_,
		_w904_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h2d0f)
	) name1262 (
		_w406_,
		_w417_,
		_w389_,
		_w869_,
		_w1477_
	);
	LUT4 #(
		.INIT('he020)
	) name1263 (
		_w390_,
		_w781_,
		_w878_,
		_w1477_,
		_w1478_
	);
	LUT3 #(
		.INIT('ha8)
	) name1264 (
		_w389_,
		_w906_,
		_w907_,
		_w1479_
	);
	LUT3 #(
		.INIT('ha8)
	) name1265 (
		_w390_,
		_w909_,
		_w910_,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w1478_,
		_w1481_,
		_w1482_
	);
	LUT4 #(
		.INIT('h3100)
	) name1268 (
		_w858_,
		_w1476_,
		_w1473_,
		_w1482_,
		_w1483_
	);
	LUT4 #(
		.INIT('h1311)
	) name1269 (
		_w918_,
		_w1469_,
		_w1472_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h2)
	) name1270 (
		\reg3_reg[20]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1485_
	);
	LUT3 #(
		.INIT('h07)
	) name1271 (
		_w269_,
		_w390_,
		_w1485_,
		_w1486_
	);
	LUT3 #(
		.INIT('h2f)
	) name1272 (
		\state_reg[0]/NET0131 ,
		_w1484_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h07)
	) name1273 (
		_w490_,
		_w619_,
		_w445_,
		_w1488_
	);
	LUT4 #(
		.INIT('h0001)
	) name1274 (
		_w463_,
		_w471_,
		_w444_,
		_w618_,
		_w1489_
	);
	LUT4 #(
		.INIT('h0001)
	) name1275 (
		_w398_,
		_w413_,
		_w424_,
		_w450_,
		_w1490_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		_w671_,
		_w380_,
		_w1491_
	);
	LUT3 #(
		.INIT('h80)
	) name1277 (
		_w671_,
		_w380_,
		_w1490_,
		_w1492_
	);
	LUT4 #(
		.INIT('h7300)
	) name1278 (
		_w1383_,
		_w1488_,
		_w1489_,
		_w1492_,
		_w1493_
	);
	LUT3 #(
		.INIT('h15)
	) name1279 (
		_w399_,
		_w448_,
		_w451_,
		_w1494_
	);
	LUT3 #(
		.INIT('h07)
	) name1280 (
		_w671_,
		_w403_,
		_w354_,
		_w1495_
	);
	LUT3 #(
		.INIT('hd0)
	) name1281 (
		_w1491_,
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT4 #(
		.INIT('h4844)
	) name1282 (
		_w700_,
		_w781_,
		_w1493_,
		_w1496_,
		_w1497_
	);
	LUT4 #(
		.INIT('h5455)
	) name1283 (
		_w329_,
		_w772_,
		_w778_,
		_w780_,
		_w1498_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		_w791_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w710_,
		_w685_,
		_w1500_
	);
	LUT4 #(
		.INIT('h0001)
	) name1286 (
		_w710_,
		_w685_,
		_w688_,
		_w798_,
		_w1501_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		_w716_,
		_w1122_,
		_w1502_
	);
	LUT3 #(
		.INIT('h40)
	) name1288 (
		_w716_,
		_w1122_,
		_w1501_,
		_w1503_
	);
	LUT4 #(
		.INIT('h0001)
	) name1289 (
		_w726_,
		_w749_,
		_w744_,
		_w794_,
		_w1504_
	);
	LUT4 #(
		.INIT('h4000)
	) name1290 (
		_w716_,
		_w1122_,
		_w1501_,
		_w1504_,
		_w1505_
	);
	LUT3 #(
		.INIT('h40)
	) name1291 (
		_w1388_,
		_w1389_,
		_w1505_,
		_w1506_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1292 (
		_w793_,
		_w808_,
		_w832_,
		_w1504_,
		_w1507_
	);
	LUT3 #(
		.INIT('h0d)
	) name1293 (
		_w797_,
		_w834_,
		_w837_,
		_w1508_
	);
	LUT3 #(
		.INIT('h8a)
	) name1294 (
		_w1503_,
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT3 #(
		.INIT('h8c)
	) name1295 (
		_w839_,
		_w851_,
		_w1500_,
		_w1510_
	);
	LUT3 #(
		.INIT('h8a)
	) name1296 (
		_w854_,
		_w850_,
		_w1122_,
		_w1511_
	);
	LUT3 #(
		.INIT('hd0)
	) name1297 (
		_w1502_,
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name1298 (
		_w1509_,
		_w1512_,
		_w1513_
	);
	LUT4 #(
		.INIT('h4844)
	) name1299 (
		_w700_,
		_w858_,
		_w1506_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1300 (
		_w277_,
		_w339_,
		_w338_,
		_w340_,
		_w1515_
	);
	LUT4 #(
		.INIT('h1c11)
	) name1301 (
		_w277_,
		_w325_,
		_w333_,
		_w1140_,
		_w1516_
	);
	LUT4 #(
		.INIT('h6300)
	) name1302 (
		_w336_,
		_w328_,
		_w874_,
		_w878_,
		_w1517_
	);
	LUT4 #(
		.INIT('h0057)
	) name1303 (
		_w904_,
		_w1515_,
		_w1516_,
		_w1517_,
		_w1518_
	);
	LUT3 #(
		.INIT('ha8)
	) name1304 (
		_w328_,
		_w906_,
		_w907_,
		_w1519_
	);
	LUT4 #(
		.INIT('he4ef)
	) name1305 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w1520_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1306 (
		_w772_,
		_w778_,
		_w780_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h0001)
	) name1307 (
		_w909_,
		_w910_,
		_w911_,
		_w1521_,
		_w1522_
	);
	LUT3 #(
		.INIT('h31)
	) name1308 (
		_w329_,
		_w1519_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h7500)
	) name1309 (
		_w781_,
		_w1514_,
		_w1518_,
		_w1523_,
		_w1524_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1310 (
		_w918_,
		_w1497_,
		_w1499_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h8)
	) name1311 (
		_w329_,
		_w919_,
		_w1526_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		\reg3_reg[26]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1527_
	);
	LUT3 #(
		.INIT('h07)
	) name1313 (
		_w269_,
		_w329_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1314 (
		\state_reg[0]/NET0131 ,
		_w1525_,
		_w1526_,
		_w1528_,
		_w1529_
	);
	LUT4 #(
		.INIT('h6050)
	) name1315 (
		_w279_,
		_w296_,
		_w878_,
		_w947_,
		_w1530_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w279_,
		_w905_,
		_w1531_
	);
	LUT3 #(
		.INIT('h70)
	) name1317 (
		_w292_,
		_w293_,
		_w904_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w953_,
		_w1532_,
		_w1533_
	);
	LUT3 #(
		.INIT('h13)
	) name1319 (
		_w953_,
		_w1531_,
		_w1532_,
		_w1534_
	);
	LUT4 #(
		.INIT('h1311)
	) name1320 (
		_w925_,
		_w957_,
		_w1530_,
		_w1534_,
		_w1535_
	);
	LUT4 #(
		.INIT('h001f)
	) name1321 (
		_w772_,
		_w778_,
		_w780_,
		_w907_,
		_w1536_
	);
	LUT3 #(
		.INIT('h20)
	) name1322 (
		\state_reg[0]/NET0131 ,
		_w909_,
		_w918_,
		_w1537_
	);
	LUT3 #(
		.INIT('h8a)
	) name1323 (
		\reg2_reg[31]/NET0131 ,
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('hf2)
	) name1324 (
		_w1110_,
		_w1535_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		\reg2_reg[26]/NET0131 ,
		_w942_,
		_w1540_
	);
	LUT4 #(
		.INIT('h4844)
	) name1326 (
		_w700_,
		_w925_,
		_w1493_,
		_w1496_,
		_w1541_
	);
	LUT4 #(
		.INIT('h0155)
	) name1327 (
		\reg2_reg[26]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1542_
	);
	LUT2 #(
		.INIT('h2)
	) name1328 (
		_w791_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		_w328_,
		_w905_,
		_w1544_
	);
	LUT3 #(
		.INIT('h04)
	) name1330 (
		_w1514_,
		_w1518_,
		_w1544_,
		_w1545_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1331 (
		_w925_,
		_w1514_,
		_w1518_,
		_w1544_,
		_w1546_
	);
	LUT4 #(
		.INIT('h0400)
	) name1332 (
		_w268_,
		_w329_,
		_w272_,
		_w645_,
		_w1547_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1333 (
		_w772_,
		_w778_,
		_w780_,
		_w858_,
		_w1548_
	);
	LUT3 #(
		.INIT('h01)
	) name1334 (
		_w909_,
		_w1359_,
		_w1548_,
		_w1549_
	);
	LUT4 #(
		.INIT('h0001)
	) name1335 (
		_w909_,
		_w1358_,
		_w1359_,
		_w1548_,
		_w1550_
	);
	LUT3 #(
		.INIT('h31)
	) name1336 (
		\reg2_reg[26]/NET0131 ,
		_w1547_,
		_w1550_,
		_w1551_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1337 (
		_w1541_,
		_w1543_,
		_w1546_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		\reg2_reg[26]/NET0131 ,
		_w919_,
		_w1553_
	);
	LUT4 #(
		.INIT('haa08)
	) name1339 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('he)
	) name1340 (
		_w1540_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\reg0_reg[20]/NET0131 ,
		_w942_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name1342 (
		\reg0_reg[20]/NET0131 ,
		_w919_,
		_w1557_
	);
	LUT4 #(
		.INIT('haa02)
	) name1343 (
		\reg0_reg[20]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1558_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1344 (
		_w686_,
		_w784_,
		_w786_,
		_w1057_,
		_w1559_
	);
	LUT3 #(
		.INIT('ha8)
	) name1345 (
		_w791_,
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1346 (
		\reg0_reg[20]/NET0131 ,
		_w686_,
		_w842_,
		_w1057_,
		_w1561_
	);
	LUT4 #(
		.INIT('hc808)
	) name1347 (
		\reg0_reg[20]/NET0131 ,
		_w904_,
		_w1057_,
		_w1475_,
		_w1562_
	);
	LUT4 #(
		.INIT('hc808)
	) name1348 (
		\reg0_reg[20]/NET0131 ,
		_w878_,
		_w1057_,
		_w1477_,
		_w1563_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w389_,
		_w905_,
		_w1564_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		_w1057_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('ha2)
	) name1351 (
		\reg0_reg[20]/NET0131 ,
		_w1063_,
		_w1325_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		_w1565_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h4)
	) name1353 (
		_w1563_,
		_w1567_,
		_w1568_
	);
	LUT4 #(
		.INIT('h3100)
	) name1354 (
		_w858_,
		_w1562_,
		_w1561_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('h1311)
	) name1355 (
		_w918_,
		_w1557_,
		_w1560_,
		_w1569_,
		_w1570_
	);
	LUT3 #(
		.INIT('hce)
	) name1356 (
		\state_reg[0]/NET0131 ,
		_w1556_,
		_w1570_,
		_w1571_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1357 (
		_w772_,
		_w778_,
		_w780_,
		_w1520_,
		_w1572_
	);
	LUT3 #(
		.INIT('h02)
	) name1358 (
		_w1063_,
		_w1325_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('hf100)
	) name1359 (
		_w772_,
		_w778_,
		_w780_,
		_w791_,
		_w1574_
	);
	LUT2 #(
		.INIT('h2)
	) name1360 (
		_w1110_,
		_w1574_,
		_w1575_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1361 (
		\reg0_reg[26]/NET0131 ,
		_w1062_,
		_w1573_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h8488)
	) name1362 (
		_w700_,
		_w791_,
		_w1493_,
		_w1496_,
		_w1577_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w1057_,
		_w1110_,
		_w1578_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name1364 (
		_w1545_,
		_w1576_,
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		\reg1_reg[11]/NET0131 ,
		_w942_,
		_w1580_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\reg1_reg[11]/NET0131 ,
		_w919_,
		_w1581_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1367 (
		\reg1_reg[11]/NET0131 ,
		_w722_,
		_w1074_,
		_w1090_,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		_w791_,
		_w1582_,
		_w1583_
	);
	LUT4 #(
		.INIT('hc808)
	) name1369 (
		\reg1_reg[11]/NET0131 ,
		_w904_,
		_w1074_,
		_w1205_,
		_w1584_
	);
	LUT4 #(
		.INIT('hc535)
	) name1370 (
		\reg1_reg[11]/NET0131 ,
		_w722_,
		_w1074_,
		_w1095_,
		_w1585_
	);
	LUT3 #(
		.INIT('ha2)
	) name1371 (
		\reg1_reg[11]/NET0131 ,
		_w1063_,
		_w1078_,
		_w1586_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w493_,
		_w905_,
		_w1587_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1373 (
		_w878_,
		_w1074_,
		_w1209_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w1586_,
		_w1588_,
		_w1589_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1375 (
		_w858_,
		_w1585_,
		_w1584_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('h1311)
	) name1376 (
		_w918_,
		_w1581_,
		_w1583_,
		_w1590_,
		_w1591_
	);
	LUT3 #(
		.INIT('hce)
	) name1377 (
		\state_reg[0]/NET0131 ,
		_w1580_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		\reg1_reg[12]/NET0131 ,
		_w942_,
		_w1593_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		\reg1_reg[12]/NET0131 ,
		_w919_,
		_w1594_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1380 (
		\reg1_reg[12]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1595_
	);
	LUT4 #(
		.INIT('hc808)
	) name1381 (
		\reg1_reg[12]/NET0131 ,
		_w791_,
		_w1074_,
		_w1222_,
		_w1596_
	);
	LUT4 #(
		.INIT('h5900)
	) name1382 (
		_w694_,
		_w809_,
		_w830_,
		_w1074_,
		_w1597_
	);
	LUT3 #(
		.INIT('ha8)
	) name1383 (
		_w858_,
		_w1595_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1384 (
		\reg1_reg[12]/NET0131 ,
		_w1074_,
		_w1226_,
		_w1227_,
		_w1599_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1385 (
		\reg1_reg[12]/NET0131 ,
		_w484_,
		_w1074_,
		_w1208_,
		_w1600_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		_w484_,
		_w905_,
		_w1601_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w1074_,
		_w1601_,
		_w1602_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1388 (
		_w772_,
		_w778_,
		_w780_,
		_w905_,
		_w1603_
	);
	LUT3 #(
		.INIT('ha2)
	) name1389 (
		\reg1_reg[12]/NET0131 ,
		_w1063_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w1602_,
		_w1604_,
		_w1605_
	);
	LUT3 #(
		.INIT('hd0)
	) name1391 (
		_w878_,
		_w1600_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('hd0)
	) name1392 (
		_w904_,
		_w1599_,
		_w1606_,
		_w1607_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1393 (
		_w918_,
		_w1596_,
		_w1598_,
		_w1607_,
		_w1608_
	);
	LUT4 #(
		.INIT('heeec)
	) name1394 (
		\state_reg[0]/NET0131 ,
		_w1593_,
		_w1594_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h2)
	) name1395 (
		\reg1_reg[20]/NET0131 ,
		_w942_,
		_w1610_
	);
	LUT2 #(
		.INIT('h8)
	) name1396 (
		\reg1_reg[20]/NET0131 ,
		_w919_,
		_w1611_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1397 (
		\reg1_reg[20]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1612_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1398 (
		_w686_,
		_w784_,
		_w786_,
		_w1074_,
		_w1613_
	);
	LUT3 #(
		.INIT('ha8)
	) name1399 (
		_w791_,
		_w1612_,
		_w1613_,
		_w1614_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1400 (
		\reg1_reg[20]/NET0131 ,
		_w686_,
		_w842_,
		_w1074_,
		_w1615_
	);
	LUT4 #(
		.INIT('hc808)
	) name1401 (
		\reg1_reg[20]/NET0131 ,
		_w904_,
		_w1074_,
		_w1475_,
		_w1616_
	);
	LUT4 #(
		.INIT('hc808)
	) name1402 (
		\reg1_reg[20]/NET0131 ,
		_w878_,
		_w1074_,
		_w1477_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		_w1074_,
		_w1564_,
		_w1618_
	);
	LUT3 #(
		.INIT('ha2)
	) name1404 (
		\reg1_reg[20]/NET0131 ,
		_w1063_,
		_w1603_,
		_w1619_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		_w1618_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h4)
	) name1406 (
		_w1617_,
		_w1620_,
		_w1621_
	);
	LUT4 #(
		.INIT('h3100)
	) name1407 (
		_w858_,
		_w1616_,
		_w1615_,
		_w1621_,
		_w1622_
	);
	LUT4 #(
		.INIT('h1311)
	) name1408 (
		_w918_,
		_w1611_,
		_w1614_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('hce)
	) name1409 (
		\state_reg[0]/NET0131 ,
		_w1610_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h2)
	) name1410 (
		\reg1_reg[24]/NET0131 ,
		_w942_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		\reg1_reg[24]/NET0131 ,
		_w919_,
		_w1626_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1412 (
		\reg1_reg[24]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1627_
	);
	LUT4 #(
		.INIT('h8488)
	) name1413 (
		_w704_,
		_w1074_,
		_w1241_,
		_w1243_,
		_w1628_
	);
	LUT3 #(
		.INIT('ha8)
	) name1414 (
		_w791_,
		_w1627_,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1415 (
		_w1074_,
		_w1246_,
		_w1248_,
		_w1249_,
		_w1630_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		_w1074_,
		_w1323_,
		_w1631_
	);
	LUT3 #(
		.INIT('ha2)
	) name1417 (
		\reg1_reg[24]/NET0131 ,
		_w1063_,
		_w1603_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT4 #(
		.INIT('h5700)
	) name1419 (
		_w904_,
		_w1627_,
		_w1630_,
		_w1633_,
		_w1634_
	);
	LUT4 #(
		.INIT('hc808)
	) name1420 (
		\reg1_reg[24]/NET0131 ,
		_w878_,
		_w1074_,
		_w1257_,
		_w1635_
	);
	LUT4 #(
		.INIT('h5060)
	) name1421 (
		_w704_,
		_w853_,
		_w1074_,
		_w1261_,
		_w1636_
	);
	LUT4 #(
		.INIT('h0507)
	) name1422 (
		_w858_,
		_w1627_,
		_w1635_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1423 (
		_w918_,
		_w1629_,
		_w1634_,
		_w1637_,
		_w1638_
	);
	LUT4 #(
		.INIT('heeec)
	) name1424 (
		\state_reg[0]/NET0131 ,
		_w1625_,
		_w1626_,
		_w1638_,
		_w1639_
	);
	LUT2 #(
		.INIT('h2)
	) name1425 (
		\reg1_reg[25]/NET0131 ,
		_w942_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		\reg1_reg[25]/NET0131 ,
		_w919_,
		_w1641_
	);
	LUT4 #(
		.INIT('h8899)
	) name1427 (
		_w268_,
		_w632_,
		_w272_,
		_w633_,
		_w1642_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1428 (
		_w772_,
		_w778_,
		_w780_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h0002)
	) name1429 (
		_w1063_,
		_w1077_,
		_w1078_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		\reg1_reg[25]/NET0131 ,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1431 (
		_w1009_,
		_w1010_,
		_w1015_,
		_w1019_,
		_w1646_
	);
	LUT4 #(
		.INIT('hf800)
	) name1432 (
		_w1008_,
		_w1021_,
		_w1022_,
		_w1029_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name1433 (
		_w1033_,
		_w1647_,
		_w1648_
	);
	LUT4 #(
		.INIT('h050d)
	) name1434 (
		_w1026_,
		_w1033_,
		_w1038_,
		_w1647_,
		_w1649_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1435 (
		_w1030_,
		_w1042_,
		_w1646_,
		_w1649_,
		_w1650_
	);
	LUT4 #(
		.INIT('h8848)
	) name1436 (
		_w682_,
		_w791_,
		_w1046_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1437 (
		_w964_,
		_w968_,
		_w969_,
		_w970_,
		_w1652_
	);
	LUT4 #(
		.INIT('h050d)
	) name1438 (
		_w966_,
		_w986_,
		_w991_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('h80f0)
	) name1439 (
		_w967_,
		_w983_,
		_w996_,
		_w1653_,
		_w1654_
	);
	LUT4 #(
		.INIT('h4484)
	) name1440 (
		_w682_,
		_w858_,
		_w1000_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		_w277_,
		_w351_,
		_w1656_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1442 (
		_w277_,
		_w333_,
		_w1140_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1443 (
		_w336_,
		_w905_,
		_w1658_
	);
	LUT4 #(
		.INIT('h9555)
	) name1444 (
		_w336_,
		_w869_,
		_w870_,
		_w873_,
		_w1659_
	);
	LUT3 #(
		.INIT('h13)
	) name1445 (
		_w878_,
		_w1658_,
		_w1659_,
		_w1660_
	);
	LUT3 #(
		.INIT('h70)
	) name1446 (
		_w904_,
		_w1657_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1447 (
		_w1074_,
		_w1651_,
		_w1655_,
		_w1661_,
		_w1662_
	);
	LUT4 #(
		.INIT('h1113)
	) name1448 (
		_w918_,
		_w1641_,
		_w1645_,
		_w1662_,
		_w1663_
	);
	LUT3 #(
		.INIT('hce)
	) name1449 (
		\state_reg[0]/NET0131 ,
		_w1640_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		\reg2_reg[12]/NET0131 ,
		_w942_,
		_w1665_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		\reg2_reg[12]/NET0131 ,
		_w919_,
		_w1666_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1452 (
		\reg2_reg[12]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1667_
	);
	LUT4 #(
		.INIT('hc808)
	) name1453 (
		\reg2_reg[12]/NET0131 ,
		_w791_,
		_w925_,
		_w1222_,
		_w1668_
	);
	LUT4 #(
		.INIT('h5900)
	) name1454 (
		_w694_,
		_w809_,
		_w830_,
		_w925_,
		_w1669_
	);
	LUT3 #(
		.INIT('ha8)
	) name1455 (
		_w858_,
		_w1667_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1456 (
		\reg2_reg[12]/NET0131 ,
		_w925_,
		_w1226_,
		_w1227_,
		_w1671_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1457 (
		\reg2_reg[12]/NET0131 ,
		_w484_,
		_w925_,
		_w1208_,
		_w1672_
	);
	LUT3 #(
		.INIT('ha8)
	) name1458 (
		\reg2_reg[12]/NET0131 ,
		_w909_,
		_w932_,
		_w1673_
	);
	LUT4 #(
		.INIT('h0400)
	) name1459 (
		_w268_,
		_w478_,
		_w272_,
		_w645_,
		_w1674_
	);
	LUT3 #(
		.INIT('h07)
	) name1460 (
		_w925_,
		_w1601_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h4)
	) name1461 (
		_w1673_,
		_w1675_,
		_w1676_
	);
	LUT3 #(
		.INIT('hd0)
	) name1462 (
		_w878_,
		_w1672_,
		_w1676_,
		_w1677_
	);
	LUT3 #(
		.INIT('hd0)
	) name1463 (
		_w904_,
		_w1671_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1464 (
		_w918_,
		_w1668_,
		_w1670_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('heeec)
	) name1465 (
		\state_reg[0]/NET0131 ,
		_w1665_,
		_w1666_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\reg2_reg[11]/NET0131 ,
		_w942_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		\reg2_reg[11]/NET0131 ,
		_w919_,
		_w1682_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1468 (
		\reg2_reg[11]/NET0131 ,
		_w722_,
		_w925_,
		_w1090_,
		_w1683_
	);
	LUT2 #(
		.INIT('h2)
	) name1469 (
		_w791_,
		_w1683_,
		_w1684_
	);
	LUT4 #(
		.INIT('hc808)
	) name1470 (
		\reg2_reg[11]/NET0131 ,
		_w904_,
		_w925_,
		_w1205_,
		_w1685_
	);
	LUT4 #(
		.INIT('hc535)
	) name1471 (
		\reg2_reg[11]/NET0131 ,
		_w722_,
		_w925_,
		_w1095_,
		_w1686_
	);
	LUT4 #(
		.INIT('hc808)
	) name1472 (
		\reg2_reg[11]/NET0131 ,
		_w878_,
		_w925_,
		_w1209_,
		_w1687_
	);
	LUT3 #(
		.INIT('ha8)
	) name1473 (
		\reg2_reg[11]/NET0131 ,
		_w909_,
		_w932_,
		_w1688_
	);
	LUT4 #(
		.INIT('h0400)
	) name1474 (
		_w268_,
		_w494_,
		_w272_,
		_w645_,
		_w1689_
	);
	LUT3 #(
		.INIT('h07)
	) name1475 (
		_w925_,
		_w1587_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h4)
	) name1477 (
		_w1687_,
		_w1691_,
		_w1692_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1478 (
		_w858_,
		_w1686_,
		_w1685_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h1311)
	) name1479 (
		_w918_,
		_w1682_,
		_w1684_,
		_w1693_,
		_w1694_
	);
	LUT3 #(
		.INIT('hce)
	) name1480 (
		\state_reg[0]/NET0131 ,
		_w1681_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h2)
	) name1481 (
		\reg0_reg[11]/NET0131 ,
		_w942_,
		_w1696_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		\reg0_reg[11]/NET0131 ,
		_w919_,
		_w1697_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1483 (
		\reg0_reg[11]/NET0131 ,
		_w722_,
		_w1057_,
		_w1090_,
		_w1698_
	);
	LUT2 #(
		.INIT('h2)
	) name1484 (
		_w791_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('hc808)
	) name1485 (
		\reg0_reg[11]/NET0131 ,
		_w904_,
		_w1057_,
		_w1205_,
		_w1700_
	);
	LUT4 #(
		.INIT('hc535)
	) name1486 (
		\reg0_reg[11]/NET0131 ,
		_w722_,
		_w1057_,
		_w1095_,
		_w1701_
	);
	LUT3 #(
		.INIT('ha2)
	) name1487 (
		\reg0_reg[11]/NET0131 ,
		_w1063_,
		_w1065_,
		_w1702_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1488 (
		_w878_,
		_w1057_,
		_w1209_,
		_w1587_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1490 (
		_w858_,
		_w1701_,
		_w1700_,
		_w1704_,
		_w1705_
	);
	LUT4 #(
		.INIT('h1311)
	) name1491 (
		_w918_,
		_w1697_,
		_w1699_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('hce)
	) name1492 (
		\state_reg[0]/NET0131 ,
		_w1696_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		\reg2_reg[20]/NET0131 ,
		_w942_,
		_w1708_
	);
	LUT2 #(
		.INIT('h8)
	) name1494 (
		\reg2_reg[20]/NET0131 ,
		_w919_,
		_w1709_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1495 (
		\reg2_reg[20]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1710_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1496 (
		_w686_,
		_w784_,
		_w786_,
		_w925_,
		_w1711_
	);
	LUT3 #(
		.INIT('ha8)
	) name1497 (
		_w791_,
		_w1710_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h3c55)
	) name1498 (
		\reg2_reg[20]/NET0131 ,
		_w686_,
		_w842_,
		_w925_,
		_w1713_
	);
	LUT4 #(
		.INIT('hc808)
	) name1499 (
		\reg2_reg[20]/NET0131 ,
		_w904_,
		_w925_,
		_w1475_,
		_w1714_
	);
	LUT4 #(
		.INIT('hc808)
	) name1500 (
		\reg2_reg[20]/NET0131 ,
		_w878_,
		_w925_,
		_w1477_,
		_w1715_
	);
	LUT3 #(
		.INIT('ha8)
	) name1501 (
		\reg2_reg[20]/NET0131 ,
		_w909_,
		_w932_,
		_w1716_
	);
	LUT4 #(
		.INIT('h0400)
	) name1502 (
		_w268_,
		_w390_,
		_w272_,
		_w645_,
		_w1717_
	);
	LUT3 #(
		.INIT('h07)
	) name1503 (
		_w925_,
		_w1564_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w1716_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h4)
	) name1505 (
		_w1715_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('h3100)
	) name1506 (
		_w858_,
		_w1714_,
		_w1713_,
		_w1720_,
		_w1721_
	);
	LUT4 #(
		.INIT('h1311)
	) name1507 (
		_w918_,
		_w1709_,
		_w1712_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('hce)
	) name1508 (
		\state_reg[0]/NET0131 ,
		_w1708_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1509 (
		\reg0_reg[12]/NET0131 ,
		_w942_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\reg0_reg[12]/NET0131 ,
		_w919_,
		_w1725_
	);
	LUT4 #(
		.INIT('haa02)
	) name1511 (
		\reg0_reg[12]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1726_
	);
	LUT4 #(
		.INIT('hc808)
	) name1512 (
		\reg0_reg[12]/NET0131 ,
		_w791_,
		_w1057_,
		_w1222_,
		_w1727_
	);
	LUT4 #(
		.INIT('h5900)
	) name1513 (
		_w694_,
		_w809_,
		_w830_,
		_w1057_,
		_w1728_
	);
	LUT3 #(
		.INIT('ha8)
	) name1514 (
		_w858_,
		_w1726_,
		_w1728_,
		_w1729_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1515 (
		\reg0_reg[12]/NET0131 ,
		_w1057_,
		_w1226_,
		_w1227_,
		_w1730_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1516 (
		\reg0_reg[12]/NET0131 ,
		_w484_,
		_w1057_,
		_w1208_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name1517 (
		_w1057_,
		_w1601_,
		_w1732_
	);
	LUT3 #(
		.INIT('ha2)
	) name1518 (
		\reg0_reg[12]/NET0131 ,
		_w1063_,
		_w1325_,
		_w1733_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT3 #(
		.INIT('hd0)
	) name1520 (
		_w878_,
		_w1731_,
		_w1734_,
		_w1735_
	);
	LUT3 #(
		.INIT('hd0)
	) name1521 (
		_w904_,
		_w1730_,
		_w1735_,
		_w1736_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1522 (
		_w918_,
		_w1727_,
		_w1729_,
		_w1736_,
		_w1737_
	);
	LUT4 #(
		.INIT('heeec)
	) name1523 (
		\state_reg[0]/NET0131 ,
		_w1724_,
		_w1725_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h2)
	) name1524 (
		\reg2_reg[24]/NET0131 ,
		_w942_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		\reg2_reg[24]/NET0131 ,
		_w919_,
		_w1740_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1526 (
		\reg2_reg[24]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1741_
	);
	LUT4 #(
		.INIT('h8488)
	) name1527 (
		_w704_,
		_w925_,
		_w1241_,
		_w1243_,
		_w1742_
	);
	LUT3 #(
		.INIT('ha8)
	) name1528 (
		_w791_,
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1529 (
		_w925_,
		_w1246_,
		_w1248_,
		_w1249_,
		_w1744_
	);
	LUT3 #(
		.INIT('ha8)
	) name1530 (
		\reg2_reg[24]/NET0131 ,
		_w909_,
		_w932_,
		_w1745_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		_w348_,
		_w907_,
		_w1746_
	);
	LUT3 #(
		.INIT('h07)
	) name1532 (
		_w925_,
		_w1323_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h4)
	) name1533 (
		_w1745_,
		_w1747_,
		_w1748_
	);
	LUT4 #(
		.INIT('h5700)
	) name1534 (
		_w904_,
		_w1741_,
		_w1744_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('hc808)
	) name1535 (
		\reg2_reg[24]/NET0131 ,
		_w878_,
		_w925_,
		_w1257_,
		_w1750_
	);
	LUT4 #(
		.INIT('h5060)
	) name1536 (
		_w704_,
		_w853_,
		_w925_,
		_w1261_,
		_w1751_
	);
	LUT4 #(
		.INIT('h0507)
	) name1537 (
		_w858_,
		_w1741_,
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1538 (
		_w918_,
		_w1743_,
		_w1749_,
		_w1752_,
		_w1753_
	);
	LUT4 #(
		.INIT('heeec)
	) name1539 (
		\state_reg[0]/NET0131 ,
		_w1739_,
		_w1740_,
		_w1753_,
		_w1754_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w257_,
		_w919_,
		_w1755_
	);
	LUT4 #(
		.INIT('h4844)
	) name1541 (
		_w743_,
		_w791_,
		_w1016_,
		_w1024_,
		_w1756_
	);
	LUT4 #(
		.INIT('h90a0)
	) name1542 (
		_w474_,
		_w484_,
		_w878_,
		_w1208_,
		_w1757_
	);
	LUT4 #(
		.INIT('h8848)
	) name1543 (
		_w743_,
		_w858_,
		_w971_,
		_w983_,
		_w1758_
	);
	LUT3 #(
		.INIT('h01)
	) name1544 (
		_w1757_,
		_w1758_,
		_w1756_,
		_w1759_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1545 (
		_w781_,
		_w1757_,
		_w1758_,
		_w1756_,
		_w1760_
	);
	LUT4 #(
		.INIT('h3633)
	) name1546 (
		_w260_,
		_w459_,
		_w480_,
		_w887_,
		_w1761_
	);
	LUT4 #(
		.INIT('h80d0)
	) name1547 (
		_w277_,
		_w480_,
		_w781_,
		_w1761_,
		_w1762_
	);
	LUT4 #(
		.INIT('h5455)
	) name1548 (
		_w257_,
		_w772_,
		_w778_,
		_w780_,
		_w1763_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		_w904_,
		_w1763_,
		_w1764_
	);
	LUT3 #(
		.INIT('h54)
	) name1550 (
		_w474_,
		_w906_,
		_w907_,
		_w1765_
	);
	LUT4 #(
		.INIT('ha4a5)
	) name1551 (
		_w268_,
		_w630_,
		_w632_,
		_w272_,
		_w1766_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1552 (
		_w772_,
		_w778_,
		_w780_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1553 (
		_w257_,
		_w909_,
		_w910_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w1765_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('hb0)
	) name1555 (
		_w1762_,
		_w1764_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h1311)
	) name1556 (
		_w918_,
		_w1755_,
		_w1760_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		\reg3_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1772_
	);
	LUT3 #(
		.INIT('h07)
	) name1558 (
		_w257_,
		_w269_,
		_w1772_,
		_w1773_
	);
	LUT3 #(
		.INIT('h2f)
	) name1559 (
		\state_reg[0]/NET0131 ,
		_w1771_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h8)
	) name1560 (
		_w427_,
		_w919_,
		_w1775_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1561 (
		_w427_,
		_w772_,
		_w778_,
		_w780_,
		_w1776_
	);
	LUT3 #(
		.INIT('h80)
	) name1562 (
		_w277_,
		_w439_,
		_w440_,
		_w1777_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1563 (
		_w277_,
		_w422_,
		_w1416_,
		_w1777_,
		_w1778_
	);
	LUT4 #(
		.INIT('he020)
	) name1564 (
		_w427_,
		_w781_,
		_w904_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('h8444)
	) name1565 (
		_w433_,
		_w781_,
		_w866_,
		_w867_,
		_w1780_
	);
	LUT3 #(
		.INIT('ha8)
	) name1566 (
		_w433_,
		_w906_,
		_w907_,
		_w1781_
	);
	LUT3 #(
		.INIT('ha8)
	) name1567 (
		_w427_,
		_w909_,
		_w910_,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT4 #(
		.INIT('h5700)
	) name1569 (
		_w878_,
		_w1776_,
		_w1780_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h4)
	) name1570 (
		_w1779_,
		_w1784_,
		_w1785_
	);
	LUT4 #(
		.INIT('h65a5)
	) name1571 (
		_w728_,
		_w1029_,
		_w1648_,
		_w1646_,
		_w1786_
	);
	LUT4 #(
		.INIT('h20e0)
	) name1572 (
		_w427_,
		_w781_,
		_w791_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1573 (
		_w964_,
		_w971_,
		_w983_,
		_w986_,
		_w1788_
	);
	LUT4 #(
		.INIT('h070b)
	) name1574 (
		_w728_,
		_w781_,
		_w1776_,
		_w1788_,
		_w1789_
	);
	LUT3 #(
		.INIT('h31)
	) name1575 (
		_w858_,
		_w1787_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h3111)
	) name1576 (
		_w918_,
		_w1775_,
		_w1785_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h2)
	) name1577 (
		\reg3_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1792_
	);
	LUT3 #(
		.INIT('h07)
	) name1578 (
		_w269_,
		_w427_,
		_w1792_,
		_w1793_
	);
	LUT3 #(
		.INIT('h2f)
	) name1579 (
		\state_reg[0]/NET0131 ,
		_w1791_,
		_w1793_,
		_w1794_
	);
	LUT3 #(
		.INIT('h54)
	) name1580 (
		_w582_,
		_w906_,
		_w907_,
		_w1795_
	);
	LUT4 #(
		.INIT('h3060)
	) name1581 (
		_w575_,
		_w742_,
		_w791_,
		_w1011_,
		_w1796_
	);
	LUT3 #(
		.INIT('h04)
	) name1582 (
		_w741_,
		_w819_,
		_w973_,
		_w1797_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name1583 (
		_w742_,
		_w818_,
		_w858_,
		_w973_,
		_w1798_
	);
	LUT4 #(
		.INIT('h1555)
	) name1584 (
		_w582_,
		_w574_,
		_w590_,
		_w597_,
		_w1799_
	);
	LUT3 #(
		.INIT('h04)
	) name1585 (
		_w860_,
		_w878_,
		_w1799_,
		_w1800_
	);
	LUT4 #(
		.INIT('h0045)
	) name1586 (
		_w1796_,
		_w1797_,
		_w1798_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1587 (
		_w277_,
		_w569_,
		_w570_,
		_w904_,
		_w1802_
	);
	LUT4 #(
		.INIT('heb00)
	) name1588 (
		_w277_,
		_w562_,
		_w881_,
		_w1802_,
		_w1803_
	);
	LUT4 #(
		.INIT('h1131)
	) name1589 (
		_w781_,
		_w1795_,
		_w1801_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1590 (
		_w772_,
		_w778_,
		_w780_,
		_w1642_,
		_w1805_
	);
	LUT4 #(
		.INIT('h0001)
	) name1591 (
		_w909_,
		_w917_,
		_w1441_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		\reg3_reg[3]/NET0131 ,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('hcc04)
	) name1593 (
		_w917_,
		_w942_,
		_w1804_,
		_w1807_,
		_w1808_
	);
	LUT3 #(
		.INIT('h9d)
	) name1594 (
		\reg3_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w268_,
		_w1809_
	);
	LUT2 #(
		.INIT('hb)
	) name1595 (
		_w1808_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w248_,
		_w919_,
		_w1811_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1597 (
		_w248_,
		_w772_,
		_w778_,
		_w780_,
		_w1812_
	);
	LUT4 #(
		.INIT('h1444)
	) name1598 (
		_w277_,
		_w544_,
		_w881_,
		_w882_,
		_w1813_
	);
	LUT3 #(
		.INIT('h80)
	) name1599 (
		_w277_,
		_w560_,
		_w561_,
		_w1814_
	);
	LUT4 #(
		.INIT('h3331)
	) name1600 (
		_w781_,
		_w1812_,
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		_w904_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h0455)
	) name1602 (
		_w812_,
		_w819_,
		_w973_,
		_w974_,
		_w1817_
	);
	LUT4 #(
		.INIT('h0b07)
	) name1603 (
		_w725_,
		_w781_,
		_w1812_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('haa65)
	) name1604 (
		_w725_,
		_w1011_,
		_w1012_,
		_w1013_,
		_w1819_
	);
	LUT4 #(
		.INIT('he020)
	) name1605 (
		_w248_,
		_w781_,
		_w791_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h9050)
	) name1606 (
		_w566_,
		_w558_,
		_w781_,
		_w860_,
		_w1821_
	);
	LUT3 #(
		.INIT('ha8)
	) name1607 (
		_w878_,
		_w1812_,
		_w1821_,
		_w1822_
	);
	LUT3 #(
		.INIT('ha8)
	) name1608 (
		_w566_,
		_w906_,
		_w907_,
		_w1823_
	);
	LUT3 #(
		.INIT('ha8)
	) name1609 (
		_w248_,
		_w909_,
		_w910_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w1823_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w1822_,
		_w1825_,
		_w1826_
	);
	LUT4 #(
		.INIT('h3100)
	) name1612 (
		_w858_,
		_w1820_,
		_w1818_,
		_w1826_,
		_w1827_
	);
	LUT4 #(
		.INIT('h1311)
	) name1613 (
		_w918_,
		_w1811_,
		_w1816_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1614 (
		\reg3_reg[5]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1829_
	);
	LUT3 #(
		.INIT('h07)
	) name1615 (
		_w248_,
		_w269_,
		_w1829_,
		_w1830_
	);
	LUT3 #(
		.INIT('h2f)
	) name1616 (
		\state_reg[0]/NET0131 ,
		_w1828_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		_w513_,
		_w919_,
		_w1832_
	);
	LUT4 #(
		.INIT('h4144)
	) name1618 (
		_w277_,
		_w503_,
		_w516_,
		_w1433_,
		_w1833_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1619 (
		_w277_,
		_w521_,
		_w522_,
		_w904_,
		_w1834_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1621 (
		_w512_,
		_w527_,
		_w863_,
		_w878_,
		_w1836_
	);
	LUT4 #(
		.INIT('h00b7)
	) name1622 (
		_w755_,
		_w858_,
		_w980_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1623 (
		_w755_,
		_w1010_,
		_w1015_,
		_w1019_,
		_w1838_
	);
	LUT4 #(
		.INIT('h1500)
	) name1624 (
		_w755_,
		_w1010_,
		_w1015_,
		_w1019_,
		_w1839_
	);
	LUT3 #(
		.INIT('h02)
	) name1625 (
		_w791_,
		_w1839_,
		_w1838_,
		_w1840_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1626 (
		_w781_,
		_w1837_,
		_w1840_,
		_w1835_,
		_w1841_
	);
	LUT3 #(
		.INIT('h54)
	) name1627 (
		_w512_,
		_w906_,
		_w907_,
		_w1842_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1628 (
		_w513_,
		_w909_,
		_w910_,
		_w1403_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('h1311)
	) name1630 (
		_w918_,
		_w1832_,
		_w1841_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		\reg3_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1846_
	);
	LUT3 #(
		.INIT('h07)
	) name1632 (
		_w269_,
		_w513_,
		_w1846_,
		_w1847_
	);
	LUT3 #(
		.INIT('h2f)
	) name1633 (
		\state_reg[0]/NET0131 ,
		_w1845_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		_w365_,
		_w919_,
		_w1849_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1635 (
		_w365_,
		_w772_,
		_w778_,
		_w780_,
		_w1850_
	);
	LUT4 #(
		.INIT('h7500)
	) name1636 (
		_w1385_,
		_w1388_,
		_w1389_,
		_w1504_,
		_w1851_
	);
	LUT4 #(
		.INIT('h50d0)
	) name1637 (
		_w1501_,
		_w1508_,
		_w1510_,
		_w1851_,
		_w1852_
	);
	LUT4 #(
		.INIT('h070b)
	) name1638 (
		_w717_,
		_w781_,
		_w1850_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		_w1489_,
		_w1490_,
		_w1854_
	);
	LUT4 #(
		.INIT('hf800)
	) name1640 (
		_w490_,
		_w619_,
		_w445_,
		_w1490_,
		_w1855_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		_w1494_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('h65aa)
	) name1642 (
		_w717_,
		_w1383_,
		_w1854_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('he020)
	) name1643 (
		_w365_,
		_w781_,
		_w791_,
		_w1857_,
		_w1858_
	);
	LUT4 #(
		.INIT('h0d05)
	) name1644 (
		_w377_,
		_w894_,
		_w1247_,
		_w1457_,
		_w1859_
	);
	LUT4 #(
		.INIT('h7020)
	) name1645 (
		_w277_,
		_w386_,
		_w781_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('h8040)
	) name1646 (
		_w363_,
		_w781_,
		_w878_,
		_w1255_,
		_w1861_
	);
	LUT3 #(
		.INIT('ha8)
	) name1647 (
		_w365_,
		_w909_,
		_w1441_,
		_w1862_
	);
	LUT3 #(
		.INIT('ha8)
	) name1648 (
		_w363_,
		_w906_,
		_w907_,
		_w1863_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w1862_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h4)
	) name1650 (
		_w1861_,
		_w1864_,
		_w1865_
	);
	LUT4 #(
		.INIT('h5700)
	) name1651 (
		_w904_,
		_w1850_,
		_w1860_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1652 (
		_w858_,
		_w1853_,
		_w1858_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1653 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w1849_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h2)
	) name1654 (
		\reg3_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w1869_
	);
	LUT4 #(
		.INIT('h4888)
	) name1655 (
		\reg3_reg[22]/NET0131 ,
		_w269_,
		_w284_,
		_w346_,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		_w1869_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('hb)
	) name1657 (
		_w1868_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('h8a)
	) name1658 (
		\reg2_reg[30]/NET0131 ,
		_w1536_,
		_w1537_,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		_w296_,
		_w905_,
		_w1874_
	);
	LUT4 #(
		.INIT('h007b)
	) name1660 (
		_w296_,
		_w878_,
		_w947_,
		_w1874_,
		_w1875_
	);
	LUT4 #(
		.INIT('h1311)
	) name1661 (
		_w925_,
		_w957_,
		_w1533_,
		_w1875_,
		_w1876_
	);
	LUT3 #(
		.INIT('hce)
	) name1662 (
		_w1110_,
		_w1873_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h2)
	) name1663 (
		\reg2_reg[7]/NET0131 ,
		_w942_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		\reg2_reg[7]/NET0131 ,
		_w919_,
		_w1879_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1665 (
		\reg2_reg[7]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1880_
	);
	LUT4 #(
		.INIT('h8884)
	) name1666 (
		_w733_,
		_w925_,
		_w1015_,
		_w1017_,
		_w1881_
	);
	LUT3 #(
		.INIT('ha8)
	) name1667 (
		_w791_,
		_w1880_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h7020)
	) name1668 (
		_w277_,
		_w544_,
		_w925_,
		_w1434_,
		_w1883_
	);
	LUT3 #(
		.INIT('ha8)
	) name1669 (
		_w904_,
		_w1880_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('h4844)
	) name1670 (
		_w733_,
		_w925_,
		_w976_,
		_w977_,
		_w1885_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		_w554_,
		_w905_,
		_w1886_
	);
	LUT4 #(
		.INIT('h0400)
	) name1672 (
		_w268_,
		_w548_,
		_w272_,
		_w645_,
		_w1887_
	);
	LUT4 #(
		.INIT('h0057)
	) name1673 (
		\reg2_reg[7]/NET0131 ,
		_w909_,
		_w1359_,
		_w1887_,
		_w1888_
	);
	LUT4 #(
		.INIT('h5700)
	) name1674 (
		_w925_,
		_w1440_,
		_w1886_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h5700)
	) name1675 (
		_w858_,
		_w1880_,
		_w1885_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1676 (
		_w918_,
		_w1884_,
		_w1882_,
		_w1890_,
		_w1891_
	);
	LUT4 #(
		.INIT('heeec)
	) name1677 (
		\state_reg[0]/NET0131 ,
		_w1878_,
		_w1879_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h19)
	) name1678 (
		_w268_,
		_w632_,
		_w762_,
		_w1893_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1679 (
		_w772_,
		_w778_,
		_w780_,
		_w1893_,
		_w1894_
	);
	LUT4 #(
		.INIT('h0020)
	) name1680 (
		_w1063_,
		_w1065_,
		_w1110_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h2)
	) name1681 (
		\reg0_reg[14]/NET0131 ,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h4)
	) name1682 (
		_w462_,
		_w905_,
		_w1897_
	);
	LUT4 #(
		.INIT('h0010)
	) name1683 (
		_w1392_,
		_w1384_,
		_w1399_,
		_w1897_,
		_w1898_
	);
	LUT3 #(
		.INIT('hce)
	) name1684 (
		_w1578_,
		_w1896_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		\reg0_reg[16]/NET0131 ,
		_w942_,
		_w1900_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		\reg0_reg[16]/NET0131 ,
		_w919_,
		_w1901_
	);
	LUT4 #(
		.INIT('haa02)
	) name1687 (
		\reg0_reg[16]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1902_
	);
	LUT4 #(
		.INIT('hc355)
	) name1688 (
		\reg0_reg[16]/NET0131 ,
		_w640_,
		_w751_,
		_w1057_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name1689 (
		_w791_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1690 (
		\reg0_reg[16]/NET0131 ,
		_w751_,
		_w1057_,
		_w1414_,
		_w1905_
	);
	LUT4 #(
		.INIT('h7020)
	) name1691 (
		_w277_,
		_w467_,
		_w1057_,
		_w1417_,
		_w1906_
	);
	LUT3 #(
		.INIT('ha8)
	) name1692 (
		_w904_,
		_w1902_,
		_w1906_,
		_w1907_
	);
	LUT3 #(
		.INIT('ha2)
	) name1693 (
		\reg0_reg[16]/NET0131 ,
		_w1063_,
		_w1065_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		_w436_,
		_w905_,
		_w1909_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1695 (
		_w878_,
		_w1057_,
		_w1420_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w1908_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1697 (
		_w858_,
		_w1905_,
		_w1907_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('h1311)
	) name1698 (
		_w918_,
		_w1901_,
		_w1904_,
		_w1912_,
		_w1913_
	);
	LUT3 #(
		.INIT('hce)
	) name1699 (
		\state_reg[0]/NET0131 ,
		_w1900_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('haa02)
	) name1700 (
		\reg0_reg[19]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1915_
	);
	LUT4 #(
		.INIT('h8488)
	) name1701 (
		_w683_,
		_w1057_,
		_w1120_,
		_w1121_,
		_w1916_
	);
	LUT3 #(
		.INIT('ha8)
	) name1702 (
		_w858_,
		_w1915_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1703 (
		\reg0_reg[19]/NET0131 ,
		_w791_,
		_w1057_,
		_w1455_,
		_w1918_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1704 (
		\reg0_reg[19]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w1919_
	);
	LUT4 #(
		.INIT('h7020)
	) name1705 (
		_w277_,
		_w422_,
		_w904_,
		_w1458_,
		_w1920_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1706 (
		_w406_,
		_w417_,
		_w869_,
		_w878_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w406_,
		_w905_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT4 #(
		.INIT('h1311)
	) name1709 (
		_w1057_,
		_w1919_,
		_w1920_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		_w1918_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		\reg0_reg[19]/NET0131 ,
		_w919_,
		_w1926_
	);
	LUT4 #(
		.INIT('h0075)
	) name1712 (
		_w918_,
		_w1917_,
		_w1925_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h2)
	) name1713 (
		\reg0_reg[19]/NET0131 ,
		_w942_,
		_w1928_
	);
	LUT3 #(
		.INIT('hf2)
	) name1714 (
		\state_reg[0]/NET0131 ,
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('haa02)
	) name1715 (
		\reg0_reg[25]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1930_
	);
	LUT4 #(
		.INIT('ha060)
	) name1716 (
		_w682_,
		_w1046_,
		_w1578_,
		_w1650_,
		_w1931_
	);
	LUT3 #(
		.INIT('ha8)
	) name1717 (
		_w791_,
		_w1930_,
		_w1931_,
		_w1932_
	);
	LUT4 #(
		.INIT('hf100)
	) name1718 (
		_w772_,
		_w778_,
		_w780_,
		_w858_,
		_w1933_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		_w1110_,
		_w1933_,
		_w1934_
	);
	LUT3 #(
		.INIT('h2a)
	) name1720 (
		\reg0_reg[25]/NET0131 ,
		_w1066_,
		_w1934_,
		_w1935_
	);
	LUT4 #(
		.INIT('h0075)
	) name1721 (
		_w1578_,
		_w1655_,
		_w1661_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('hb)
	) name1722 (
		_w1932_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		\reg0_reg[30]/NET0131 ,
		_w1895_,
		_w1938_
	);
	LUT3 #(
		.INIT('hf2)
	) name1724 (
		_w1578_,
		_w1875_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h2)
	) name1725 (
		\reg0_reg[31]/NET0131 ,
		_w1895_,
		_w1940_
	);
	LUT4 #(
		.INIT('hffb0)
	) name1726 (
		_w1530_,
		_w1534_,
		_w1578_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		\reg0_reg[7]/NET0131 ,
		_w942_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1728 (
		\reg0_reg[7]/NET0131 ,
		_w919_,
		_w1943_
	);
	LUT4 #(
		.INIT('haa02)
	) name1729 (
		\reg0_reg[7]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1944_
	);
	LUT4 #(
		.INIT('h7020)
	) name1730 (
		_w277_,
		_w544_,
		_w1057_,
		_w1434_,
		_w1945_
	);
	LUT3 #(
		.INIT('ha8)
	) name1731 (
		_w904_,
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('ha900)
	) name1732 (
		_w733_,
		_w1015_,
		_w1017_,
		_w1057_,
		_w1947_
	);
	LUT3 #(
		.INIT('ha8)
	) name1733 (
		_w791_,
		_w1944_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h6500)
	) name1734 (
		_w733_,
		_w976_,
		_w977_,
		_w1057_,
		_w1949_
	);
	LUT3 #(
		.INIT('ha2)
	) name1735 (
		\reg0_reg[7]/NET0131 ,
		_w1063_,
		_w1065_,
		_w1950_
	);
	LUT4 #(
		.INIT('h0057)
	) name1736 (
		_w1057_,
		_w1440_,
		_w1886_,
		_w1950_,
		_w1951_
	);
	LUT4 #(
		.INIT('h5700)
	) name1737 (
		_w858_,
		_w1944_,
		_w1949_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1738 (
		_w918_,
		_w1948_,
		_w1946_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('heeec)
	) name1739 (
		\state_reg[0]/NET0131 ,
		_w1942_,
		_w1943_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('h2)
	) name1740 (
		\reg0_reg[8]/NET0131 ,
		_w942_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		\reg0_reg[8]/NET0131 ,
		_w919_,
		_w1956_
	);
	LUT4 #(
		.INIT('hc355)
	) name1742 (
		\reg0_reg[8]/NET0131 ,
		_w610_,
		_w738_,
		_w1057_,
		_w1957_
	);
	LUT2 #(
		.INIT('h2)
	) name1743 (
		_w791_,
		_w1957_,
		_w1958_
	);
	LUT3 #(
		.INIT('h80)
	) name1744 (
		_w277_,
		_w547_,
		_w549_,
		_w1959_
	);
	LUT4 #(
		.INIT('h00eb)
	) name1745 (
		_w277_,
		_w516_,
		_w1433_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('hc808)
	) name1746 (
		\reg0_reg[8]/NET0131 ,
		_w904_,
		_w1057_,
		_w1960_,
		_w1961_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1747 (
		_w738_,
		_w811_,
		_w822_,
		_w827_,
		_w1962_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1748 (
		\reg0_reg[8]/NET0131 ,
		_w858_,
		_w1057_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('ha2)
	) name1749 (
		\reg0_reg[8]/NET0131 ,
		_w1063_,
		_w1065_,
		_w1964_
	);
	LUT2 #(
		.INIT('h8)
	) name1750 (
		_w527_,
		_w905_,
		_w1965_
	);
	LUT4 #(
		.INIT('h006f)
	) name1751 (
		_w527_,
		_w863_,
		_w878_,
		_w1965_,
		_w1966_
	);
	LUT3 #(
		.INIT('h31)
	) name1752 (
		_w1057_,
		_w1964_,
		_w1966_,
		_w1967_
	);
	LUT3 #(
		.INIT('h10)
	) name1753 (
		_w1961_,
		_w1963_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h1311)
	) name1754 (
		_w918_,
		_w1956_,
		_w1958_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('hce)
	) name1755 (
		\state_reg[0]/NET0131 ,
		_w1955_,
		_w1969_,
		_w1970_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1756 (
		_w772_,
		_w778_,
		_w780_,
		_w1893_,
		_w1971_
	);
	LUT4 #(
		.INIT('h0020)
	) name1757 (
		_w1063_,
		_w1078_,
		_w1110_,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		\reg1_reg[14]/NET0131 ,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		_w1074_,
		_w1110_,
		_w1974_
	);
	LUT3 #(
		.INIT('hdc)
	) name1760 (
		_w1898_,
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h2)
	) name1761 (
		\reg1_reg[16]/NET0131 ,
		_w942_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		\reg1_reg[16]/NET0131 ,
		_w919_,
		_w1977_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1763 (
		\reg1_reg[16]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1978_
	);
	LUT4 #(
		.INIT('hc355)
	) name1764 (
		\reg1_reg[16]/NET0131 ,
		_w640_,
		_w751_,
		_w1074_,
		_w1979_
	);
	LUT2 #(
		.INIT('h2)
	) name1765 (
		_w791_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1766 (
		\reg1_reg[16]/NET0131 ,
		_w751_,
		_w1074_,
		_w1414_,
		_w1981_
	);
	LUT4 #(
		.INIT('h7020)
	) name1767 (
		_w277_,
		_w467_,
		_w1074_,
		_w1417_,
		_w1982_
	);
	LUT3 #(
		.INIT('ha8)
	) name1768 (
		_w904_,
		_w1978_,
		_w1982_,
		_w1983_
	);
	LUT3 #(
		.INIT('ha2)
	) name1769 (
		\reg1_reg[16]/NET0131 ,
		_w1063_,
		_w1078_,
		_w1984_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1770 (
		_w878_,
		_w1074_,
		_w1420_,
		_w1909_,
		_w1985_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w1984_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1772 (
		_w858_,
		_w1981_,
		_w1983_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h1311)
	) name1773 (
		_w918_,
		_w1977_,
		_w1980_,
		_w1987_,
		_w1988_
	);
	LUT3 #(
		.INIT('hce)
	) name1774 (
		\state_reg[0]/NET0131 ,
		_w1976_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		\reg1_reg[19]/NET0131 ,
		_w942_,
		_w1990_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1776 (
		\reg1_reg[19]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w1991_
	);
	LUT4 #(
		.INIT('h8488)
	) name1777 (
		_w683_,
		_w1074_,
		_w1120_,
		_w1121_,
		_w1992_
	);
	LUT3 #(
		.INIT('ha8)
	) name1778 (
		_w858_,
		_w1991_,
		_w1992_,
		_w1993_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1779 (
		\reg1_reg[19]/NET0131 ,
		_w791_,
		_w1074_,
		_w1455_,
		_w1994_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1780 (
		\reg1_reg[19]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w1995_
	);
	LUT4 #(
		.INIT('h0075)
	) name1781 (
		_w1074_,
		_w1920_,
		_w1923_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w1994_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		\reg1_reg[19]/NET0131 ,
		_w919_,
		_w1998_
	);
	LUT4 #(
		.INIT('h0075)
	) name1784 (
		_w918_,
		_w1993_,
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT3 #(
		.INIT('hce)
	) name1785 (
		\state_reg[0]/NET0131 ,
		_w1990_,
		_w1999_,
		_w2000_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1786 (
		_w772_,
		_w778_,
		_w780_,
		_w1520_,
		_w2001_
	);
	LUT3 #(
		.INIT('h02)
	) name1787 (
		_w1063_,
		_w1603_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1788 (
		_w772_,
		_w778_,
		_w780_,
		_w791_,
		_w2003_
	);
	LUT2 #(
		.INIT('h2)
	) name1789 (
		_w1110_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('h2a)
	) name1790 (
		\reg1_reg[26]/NET0131 ,
		_w2002_,
		_w2004_,
		_w2005_
	);
	LUT4 #(
		.INIT('hffd0)
	) name1791 (
		_w1545_,
		_w1577_,
		_w1974_,
		_w2005_,
		_w2006_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1792 (
		\reg1_reg[30]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2007_
	);
	LUT4 #(
		.INIT('h006f)
	) name1793 (
		_w296_,
		_w947_,
		_w1974_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h0008)
	) name1794 (
		_w1063_,
		_w1110_,
		_w1603_,
		_w1971_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		\reg1_reg[30]/NET0131 ,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('hf800)
	) name1796 (
		_w953_,
		_w1532_,
		_w1874_,
		_w1974_,
		_w2011_
	);
	LUT4 #(
		.INIT('hffce)
	) name1797 (
		_w878_,
		_w2010_,
		_w2008_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		\reg1_reg[31]/NET0131 ,
		_w1972_,
		_w2013_
	);
	LUT4 #(
		.INIT('hffb0)
	) name1799 (
		_w1530_,
		_w1534_,
		_w1974_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h2)
	) name1800 (
		\reg1_reg[7]/NET0131 ,
		_w942_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		\reg1_reg[7]/NET0131 ,
		_w919_,
		_w2016_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1802 (
		\reg1_reg[7]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2017_
	);
	LUT4 #(
		.INIT('h7020)
	) name1803 (
		_w277_,
		_w544_,
		_w1074_,
		_w1434_,
		_w2018_
	);
	LUT3 #(
		.INIT('ha8)
	) name1804 (
		_w904_,
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('ha900)
	) name1805 (
		_w733_,
		_w1015_,
		_w1017_,
		_w1074_,
		_w2020_
	);
	LUT3 #(
		.INIT('ha8)
	) name1806 (
		_w791_,
		_w2017_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h6500)
	) name1807 (
		_w733_,
		_w976_,
		_w977_,
		_w1074_,
		_w2022_
	);
	LUT3 #(
		.INIT('ha2)
	) name1808 (
		\reg1_reg[7]/NET0131 ,
		_w1063_,
		_w1078_,
		_w2023_
	);
	LUT4 #(
		.INIT('h0057)
	) name1809 (
		_w1074_,
		_w1440_,
		_w1886_,
		_w2023_,
		_w2024_
	);
	LUT4 #(
		.INIT('h5700)
	) name1810 (
		_w858_,
		_w2017_,
		_w2022_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1811 (
		_w918_,
		_w2021_,
		_w2019_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('heeec)
	) name1812 (
		\state_reg[0]/NET0131 ,
		_w2015_,
		_w2016_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1813 (
		_w772_,
		_w778_,
		_w780_,
		_w791_,
		_w2028_
	);
	LUT2 #(
		.INIT('h2)
	) name1814 (
		_w1110_,
		_w2028_,
		_w2029_
	);
	LUT3 #(
		.INIT('ha2)
	) name1815 (
		\reg2_reg[14]/NET0131 ,
		_w1110_,
		_w2028_,
		_w2030_
	);
	LUT4 #(
		.INIT('h0400)
	) name1816 (
		_w268_,
		_w455_,
		_w272_,
		_w645_,
		_w2031_
	);
	LUT3 #(
		.INIT('h90)
	) name1817 (
		_w268_,
		_w632_,
		_w762_,
		_w2032_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1818 (
		_w772_,
		_w778_,
		_w780_,
		_w2032_,
		_w2033_
	);
	LUT4 #(
		.INIT('h0001)
	) name1819 (
		_w909_,
		_w932_,
		_w1548_,
		_w2033_,
		_w2034_
	);
	LUT3 #(
		.INIT('h31)
	) name1820 (
		\reg2_reg[14]/NET0131 ,
		_w2031_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1821 (
		_w925_,
		_w1110_,
		_w1898_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('he)
	) name1822 (
		_w2030_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h2)
	) name1823 (
		\reg2_reg[16]/NET0131 ,
		_w942_,
		_w2038_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		\reg2_reg[16]/NET0131 ,
		_w919_,
		_w2039_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1825 (
		\reg2_reg[16]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2040_
	);
	LUT4 #(
		.INIT('hc355)
	) name1826 (
		\reg2_reg[16]/NET0131 ,
		_w640_,
		_w751_,
		_w925_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		_w791_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1828 (
		\reg2_reg[16]/NET0131 ,
		_w751_,
		_w925_,
		_w1414_,
		_w2043_
	);
	LUT4 #(
		.INIT('h7020)
	) name1829 (
		_w277_,
		_w467_,
		_w925_,
		_w1417_,
		_w2044_
	);
	LUT3 #(
		.INIT('ha8)
	) name1830 (
		_w904_,
		_w2040_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1831 (
		_w878_,
		_w925_,
		_w1420_,
		_w1909_,
		_w2046_
	);
	LUT4 #(
		.INIT('h0400)
	) name1832 (
		_w268_,
		_w438_,
		_w272_,
		_w645_,
		_w2047_
	);
	LUT4 #(
		.INIT('h0057)
	) name1833 (
		\reg2_reg[16]/NET0131 ,
		_w909_,
		_w1359_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w2046_,
		_w2048_,
		_w2049_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1835 (
		_w858_,
		_w2043_,
		_w2045_,
		_w2049_,
		_w2050_
	);
	LUT4 #(
		.INIT('h1311)
	) name1836 (
		_w918_,
		_w2039_,
		_w2042_,
		_w2050_,
		_w2051_
	);
	LUT3 #(
		.INIT('hce)
	) name1837 (
		\state_reg[0]/NET0131 ,
		_w2038_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		\reg2_reg[19]/NET0131 ,
		_w942_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name1839 (
		\reg2_reg[19]/NET0131 ,
		_w919_,
		_w2054_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1840 (
		\reg2_reg[19]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2055_
	);
	LUT4 #(
		.INIT('h8488)
	) name1841 (
		_w683_,
		_w925_,
		_w1120_,
		_w1121_,
		_w2056_
	);
	LUT3 #(
		.INIT('ha8)
	) name1842 (
		_w858_,
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1843 (
		\reg2_reg[19]/NET0131 ,
		_w791_,
		_w925_,
		_w1455_,
		_w2058_
	);
	LUT4 #(
		.INIT('h0400)
	) name1844 (
		_w268_,
		_w407_,
		_w272_,
		_w645_,
		_w2059_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1845 (
		\reg2_reg[19]/NET0131 ,
		_w909_,
		_w932_,
		_w2033_,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h7500)
	) name1847 (
		_w925_,
		_w1920_,
		_w1923_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		_w2058_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h1311)
	) name1849 (
		_w918_,
		_w2054_,
		_w2057_,
		_w2063_,
		_w2064_
	);
	LUT3 #(
		.INIT('hce)
	) name1850 (
		\state_reg[0]/NET0131 ,
		_w2053_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		\reg2_reg[25]/NET0131 ,
		_w942_,
		_w2066_
	);
	LUT2 #(
		.INIT('h8)
	) name1852 (
		\reg2_reg[25]/NET0131 ,
		_w919_,
		_w2067_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1853 (
		\reg2_reg[25]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2068_
	);
	LUT4 #(
		.INIT('h8848)
	) name1854 (
		_w682_,
		_w925_,
		_w1046_,
		_w1650_,
		_w2069_
	);
	LUT3 #(
		.INIT('ha8)
	) name1855 (
		_w791_,
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT4 #(
		.INIT('h4484)
	) name1856 (
		_w682_,
		_w925_,
		_w1000_,
		_w1654_,
		_w2071_
	);
	LUT3 #(
		.INIT('ha8)
	) name1857 (
		_w858_,
		_w2068_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('hc808)
	) name1858 (
		\reg2_reg[25]/NET0131 ,
		_w904_,
		_w925_,
		_w1657_,
		_w2073_
	);
	LUT4 #(
		.INIT('hc808)
	) name1859 (
		\reg2_reg[25]/NET0131 ,
		_w878_,
		_w925_,
		_w1659_,
		_w2074_
	);
	LUT3 #(
		.INIT('ha8)
	) name1860 (
		\reg2_reg[25]/NET0131 ,
		_w909_,
		_w932_,
		_w2075_
	);
	LUT4 #(
		.INIT('h0400)
	) name1861 (
		_w268_,
		_w337_,
		_w272_,
		_w645_,
		_w2076_
	);
	LUT3 #(
		.INIT('h07)
	) name1862 (
		_w925_,
		_w1658_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w2075_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		_w2074_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name1865 (
		_w2073_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1866 (
		_w918_,
		_w2070_,
		_w2072_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('heeec)
	) name1867 (
		\state_reg[0]/NET0131 ,
		_w2066_,
		_w2067_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		\reg3_reg[1]/NET0131 ,
		_w942_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		\reg3_reg[1]/NET0131 ,
		_w919_,
		_w2084_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1870 (
		\reg3_reg[1]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2085_
	);
	LUT4 #(
		.INIT('h2d00)
	) name1871 (
		_w595_,
		_w597_,
		_w756_,
		_w781_,
		_w2086_
	);
	LUT3 #(
		.INIT('ha8)
	) name1872 (
		_w791_,
		_w2085_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('h4144)
	) name1873 (
		_w277_,
		_w571_,
		_w587_,
		_w880_,
		_w2088_
	);
	LUT3 #(
		.INIT('h80)
	) name1874 (
		_w277_,
		_w593_,
		_w594_,
		_w2089_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1875 (
		\reg3_reg[1]/NET0131 ,
		_w781_,
		_w2088_,
		_w2089_,
		_w2090_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1876 (
		\reg3_reg[1]/NET0131 ,
		_w756_,
		_w781_,
		_w815_,
		_w2091_
	);
	LUT2 #(
		.INIT('h6)
	) name1877 (
		_w590_,
		_w597_,
		_w2092_
	);
	LUT4 #(
		.INIT('he020)
	) name1878 (
		\reg3_reg[1]/NET0131 ,
		_w781_,
		_w878_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h0100)
	) name1879 (
		_w590_,
		_w772_,
		_w778_,
		_w780_,
		_w2094_
	);
	LUT4 #(
		.INIT('h0080)
	) name1880 (
		\reg3_reg[1]/NET0131 ,
		_w268_,
		_w632_,
		_w762_,
		_w2095_
	);
	LUT3 #(
		.INIT('h0b)
	) name1881 (
		_w590_,
		_w907_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('h5700)
	) name1882 (
		_w905_,
		_w2085_,
		_w2094_,
		_w2096_,
		_w2097_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1883 (
		_w858_,
		_w2091_,
		_w2093_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1884 (
		_w904_,
		_w2090_,
		_w2087_,
		_w2098_,
		_w2099_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1885 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2084_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('he)
	) name1886 (
		_w2083_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		\reg3_reg[2]/NET0131 ,
		_w942_,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name1888 (
		\reg3_reg[2]/NET0131 ,
		_w919_,
		_w2103_
	);
	LUT4 #(
		.INIT('h5655)
	) name1889 (
		_w578_,
		_w571_,
		_w587_,
		_w880_,
		_w2104_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1890 (
		_w277_,
		_w585_,
		_w586_,
		_w904_,
		_w2105_
	);
	LUT3 #(
		.INIT('he0)
	) name1891 (
		_w277_,
		_w2104_,
		_w2105_,
		_w2106_
	);
	LUT4 #(
		.INIT('h0701)
	) name1892 (
		_w587_,
		_w590_,
		_w747_,
		_w815_,
		_w2107_
	);
	LUT4 #(
		.INIT('h80e0)
	) name1893 (
		_w587_,
		_w590_,
		_w747_,
		_w815_,
		_w2108_
	);
	LUT3 #(
		.INIT('h02)
	) name1894 (
		_w858_,
		_w2108_,
		_w2107_,
		_w2109_
	);
	LUT4 #(
		.INIT('h4d00)
	) name1895 (
		_w587_,
		_w590_,
		_w598_,
		_w747_,
		_w2110_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1896 (
		_w587_,
		_w590_,
		_w598_,
		_w747_,
		_w2111_
	);
	LUT3 #(
		.INIT('h02)
	) name1897 (
		_w791_,
		_w2111_,
		_w2110_,
		_w2112_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1898 (
		_w781_,
		_w2109_,
		_w2106_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w574_,
		_w907_,
		_w2114_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1900 (
		\reg3_reg[2]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2115_
	);
	LUT3 #(
		.INIT('h6a)
	) name1901 (
		_w574_,
		_w590_,
		_w597_,
		_w2116_
	);
	LUT4 #(
		.INIT('he020)
	) name1902 (
		\reg3_reg[2]/NET0131 ,
		_w781_,
		_w878_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1903 (
		_w772_,
		_w778_,
		_w780_,
		_w1893_,
		_w2118_
	);
	LUT3 #(
		.INIT('ha8)
	) name1904 (
		\reg3_reg[2]/NET0131 ,
		_w909_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h0100)
	) name1905 (
		_w574_,
		_w772_,
		_w778_,
		_w780_,
		_w2120_
	);
	LUT3 #(
		.INIT('ha8)
	) name1906 (
		_w905_,
		_w2115_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h0001)
	) name1907 (
		_w2114_,
		_w2117_,
		_w2119_,
		_w2121_,
		_w2122_
	);
	LUT4 #(
		.INIT('h1311)
	) name1908 (
		_w918_,
		_w2103_,
		_w2113_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('hce)
	) name1909 (
		\state_reg[0]/NET0131 ,
		_w2102_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h8)
	) name1910 (
		_w559_,
		_w919_,
		_w2125_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1911 (
		_w559_,
		_w772_,
		_w778_,
		_w780_,
		_w2126_
	);
	LUT3 #(
		.INIT('h2a)
	) name1912 (
		_w277_,
		_w576_,
		_w577_,
		_w2127_
	);
	LUT4 #(
		.INIT('h1211)
	) name1913 (
		_w251_,
		_w277_,
		_w562_,
		_w881_,
		_w2128_
	);
	LUT4 #(
		.INIT('h1113)
	) name1914 (
		_w781_,
		_w2126_,
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h2)
	) name1915 (
		_w904_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1916 (
		_w584_,
		_w599_,
		_w602_,
		_w734_,
		_w2131_
	);
	LUT4 #(
		.INIT('he020)
	) name1917 (
		_w559_,
		_w781_,
		_w791_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h559a)
	) name1918 (
		_w734_,
		_w817_,
		_w819_,
		_w821_,
		_w2133_
	);
	LUT4 #(
		.INIT('h20e0)
	) name1919 (
		_w559_,
		_w781_,
		_w858_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('h00b7)
	) name1920 (
		_w558_,
		_w781_,
		_w860_,
		_w2126_,
		_w2135_
	);
	LUT3 #(
		.INIT('h54)
	) name1921 (
		_w558_,
		_w906_,
		_w907_,
		_w2136_
	);
	LUT3 #(
		.INIT('ha8)
	) name1922 (
		_w559_,
		_w909_,
		_w910_,
		_w2137_
	);
	LUT4 #(
		.INIT('h0031)
	) name1923 (
		_w878_,
		_w2136_,
		_w2135_,
		_w2137_,
		_w2138_
	);
	LUT3 #(
		.INIT('h10)
	) name1924 (
		_w2134_,
		_w2132_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h1311)
	) name1925 (
		_w918_,
		_w2125_,
		_w2130_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name1926 (
		\reg3_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2141_
	);
	LUT3 #(
		.INIT('h07)
	) name1927 (
		_w269_,
		_w559_,
		_w2141_,
		_w2142_
	);
	LUT3 #(
		.INIT('h2f)
	) name1928 (
		\state_reg[0]/NET0131 ,
		_w2140_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		_w542_,
		_w919_,
		_w2144_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1930 (
		_w542_,
		_w772_,
		_w778_,
		_w780_,
		_w2145_
	);
	LUT4 #(
		.INIT('h4b00)
	) name1931 (
		_w603_,
		_w606_,
		_w695_,
		_w781_,
		_w2146_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name1932 (
		_w540_,
		_w566_,
		_w558_,
		_w860_,
		_w2147_
	);
	LUT4 #(
		.INIT('he020)
	) name1933 (
		_w542_,
		_w781_,
		_w878_,
		_w2147_,
		_w2148_
	);
	LUT3 #(
		.INIT('h54)
	) name1934 (
		_w540_,
		_w906_,
		_w907_,
		_w2149_
	);
	LUT3 #(
		.INIT('ha8)
	) name1935 (
		_w542_,
		_w909_,
		_w910_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w2149_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name1937 (
		_w2148_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h5700)
	) name1938 (
		_w791_,
		_w2145_,
		_w2146_,
		_w2152_,
		_w2153_
	);
	LUT3 #(
		.INIT('h70)
	) name1939 (
		_w246_,
		_w250_,
		_w277_,
		_w2154_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1940 (
		_w544_,
		_w550_,
		_w881_,
		_w882_,
		_w2155_
	);
	LUT4 #(
		.INIT('h1555)
	) name1941 (
		_w277_,
		_w881_,
		_w882_,
		_w883_,
		_w2156_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1942 (
		_w781_,
		_w2154_,
		_w2155_,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('ha8)
	) name1943 (
		_w904_,
		_w2145_,
		_w2157_,
		_w2158_
	);
	LUT4 #(
		.INIT('h8488)
	) name1944 (
		_w695_,
		_w781_,
		_w822_,
		_w824_,
		_w2159_
	);
	LUT3 #(
		.INIT('ha8)
	) name1945 (
		_w858_,
		_w2145_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1946 (
		_w918_,
		_w2158_,
		_w2160_,
		_w2153_,
		_w2161_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		\reg3_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2162_
	);
	LUT3 #(
		.INIT('h07)
	) name1948 (
		_w269_,
		_w542_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1949 (
		\state_reg[0]/NET0131 ,
		_w2144_,
		_w2161_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name1950 (
		_w520_,
		_w919_,
		_w2165_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1951 (
		_w520_,
		_w772_,
		_w778_,
		_w780_,
		_w2166_
	);
	LUT4 #(
		.INIT('he020)
	) name1952 (
		_w520_,
		_w781_,
		_w904_,
		_w1960_,
		_w2167_
	);
	LUT4 #(
		.INIT('h009f)
	) name1953 (
		_w610_,
		_w738_,
		_w781_,
		_w2166_,
		_w2168_
	);
	LUT4 #(
		.INIT('h20e0)
	) name1954 (
		_w520_,
		_w781_,
		_w858_,
		_w1962_,
		_w2169_
	);
	LUT4 #(
		.INIT('h8400)
	) name1955 (
		_w527_,
		_w781_,
		_w863_,
		_w878_,
		_w2170_
	);
	LUT3 #(
		.INIT('ha8)
	) name1956 (
		_w520_,
		_w909_,
		_w1441_,
		_w2171_
	);
	LUT3 #(
		.INIT('ha8)
	) name1957 (
		_w527_,
		_w906_,
		_w907_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name1958 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name1959 (
		_w2170_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1960 (
		_w791_,
		_w2168_,
		_w2169_,
		_w2174_,
		_w2175_
	);
	LUT4 #(
		.INIT('h1311)
	) name1961 (
		_w918_,
		_w2165_,
		_w2167_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		\reg3_reg[8]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2177_
	);
	LUT3 #(
		.INIT('h07)
	) name1963 (
		_w269_,
		_w520_,
		_w2177_,
		_w2178_
	);
	LUT3 #(
		.INIT('h2f)
	) name1964 (
		\state_reg[0]/NET0131 ,
		_w2176_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		\reg3_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2180_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1966 (
		_w500_,
		_w772_,
		_w778_,
		_w780_,
		_w2181_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1967 (
		_w497_,
		_w503_,
		_w516_,
		_w1433_,
		_w2182_
	);
	LUT3 #(
		.INIT('h80)
	) name1968 (
		_w277_,
		_w514_,
		_w515_,
		_w2183_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1969 (
		_w277_,
		_w887_,
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT4 #(
		.INIT('he020)
	) name1970 (
		_w500_,
		_w781_,
		_w904_,
		_w2184_,
		_w2185_
	);
	LUT4 #(
		.INIT('h8488)
	) name1971 (
		_w754_,
		_w781_,
		_w1379_,
		_w1380_,
		_w2186_
	);
	LUT3 #(
		.INIT('ha8)
	) name1972 (
		_w791_,
		_w2181_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('h007b)
	) name1973 (
		_w754_,
		_w781_,
		_w1388_,
		_w2181_,
		_w2188_
	);
	LUT4 #(
		.INIT('h9500)
	) name1974 (
		_w508_,
		_w863_,
		_w864_,
		_w878_,
		_w2189_
	);
	LUT3 #(
		.INIT('ha8)
	) name1975 (
		_w508_,
		_w906_,
		_w907_,
		_w2190_
	);
	LUT4 #(
		.INIT('h5070)
	) name1976 (
		_w500_,
		_w909_,
		_w918_,
		_w1441_,
		_w2191_
	);
	LUT2 #(
		.INIT('h4)
	) name1977 (
		_w2190_,
		_w2191_,
		_w2192_
	);
	LUT3 #(
		.INIT('h70)
	) name1978 (
		_w781_,
		_w2189_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('hd0)
	) name1979 (
		_w858_,
		_w2188_,
		_w2193_,
		_w2194_
	);
	LUT3 #(
		.INIT('ha8)
	) name1980 (
		\state_reg[0]/NET0131 ,
		_w500_,
		_w918_,
		_w2195_
	);
	LUT4 #(
		.INIT('hef00)
	) name1981 (
		_w2185_,
		_w2187_,
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('he)
	) name1982 (
		_w2180_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		\reg3_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2198_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1984 (
		_w418_,
		_w772_,
		_w778_,
		_w780_,
		_w2199_
	);
	LUT4 #(
		.INIT('h6a5a)
	) name1985 (
		_w689_,
		_w1383_,
		_w1488_,
		_w1489_,
		_w2200_
	);
	LUT4 #(
		.INIT('he020)
	) name1986 (
		_w418_,
		_w781_,
		_w791_,
		_w2200_,
		_w2201_
	);
	LUT4 #(
		.INIT('h0705)
	) name1987 (
		_w411_,
		_w422_,
		_w893_,
		_w1416_,
		_w2202_
	);
	LUT4 #(
		.INIT('h7020)
	) name1988 (
		_w277_,
		_w429_,
		_w781_,
		_w2202_,
		_w2203_
	);
	LUT3 #(
		.INIT('ha8)
	) name1989 (
		_w904_,
		_w2199_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('h4484)
	) name1990 (
		_w689_,
		_w781_,
		_w1508_,
		_w1851_,
		_w2205_
	);
	LUT4 #(
		.INIT('h8400)
	) name1991 (
		_w417_,
		_w781_,
		_w869_,
		_w878_,
		_w2206_
	);
	LUT3 #(
		.INIT('ha8)
	) name1992 (
		_w417_,
		_w906_,
		_w907_,
		_w2207_
	);
	LUT4 #(
		.INIT('h5070)
	) name1993 (
		_w418_,
		_w909_,
		_w918_,
		_w1441_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w2207_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		_w2206_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('h5700)
	) name1996 (
		_w858_,
		_w2199_,
		_w2205_,
		_w2210_,
		_w2211_
	);
	LUT3 #(
		.INIT('ha8)
	) name1997 (
		\state_reg[0]/NET0131 ,
		_w418_,
		_w918_,
		_w2212_
	);
	LUT4 #(
		.INIT('hef00)
	) name1998 (
		_w2201_,
		_w2204_,
		_w2211_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('he)
	) name1999 (
		_w2198_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w382_,
		_w919_,
		_w2215_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2001 (
		_w382_,
		_w772_,
		_w778_,
		_w780_,
		_w2216_
	);
	LUT4 #(
		.INIT('h4144)
	) name2002 (
		_w277_,
		_w369_,
		_w386_,
		_w1457_,
		_w2217_
	);
	LUT4 #(
		.INIT('h0200)
	) name2003 (
		_w277_,
		_w392_,
		_w391_,
		_w393_,
		_w2218_
	);
	LUT4 #(
		.INIT('h3331)
	) name2004 (
		_w781_,
		_w2216_,
		_w2217_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		_w904_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h007b)
	) name2006 (
		_w711_,
		_w781_,
		_w993_,
		_w2216_,
		_w2221_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		_w858_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h00b7)
	) name2008 (
		_w711_,
		_w781_,
		_w1040_,
		_w2216_,
		_w2223_
	);
	LUT4 #(
		.INIT('h8444)
	) name2009 (
		_w381_,
		_w781_,
		_w869_,
		_w870_,
		_w2224_
	);
	LUT3 #(
		.INIT('ha8)
	) name2010 (
		_w381_,
		_w906_,
		_w907_,
		_w2225_
	);
	LUT3 #(
		.INIT('ha8)
	) name2011 (
		_w382_,
		_w909_,
		_w910_,
		_w2226_
	);
	LUT2 #(
		.INIT('h1)
	) name2012 (
		_w2225_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('h5700)
	) name2013 (
		_w878_,
		_w2216_,
		_w2224_,
		_w2227_,
		_w2228_
	);
	LUT3 #(
		.INIT('hd0)
	) name2014 (
		_w791_,
		_w2223_,
		_w2228_,
		_w2229_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2015 (
		_w918_,
		_w2220_,
		_w2222_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name2016 (
		\reg3_reg[21]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2231_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2017 (
		\reg3_reg[20]/NET0131 ,
		\reg3_reg[21]/NET0131 ,
		_w269_,
		_w346_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name2018 (
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2019 (
		\state_reg[0]/NET0131 ,
		_w2215_,
		_w2230_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name2020 (
		\reg2_reg[5]/NET0131 ,
		_w942_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		\reg2_reg[5]/NET0131 ,
		_w919_,
		_w2236_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2022 (
		\reg2_reg[5]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2237_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2023 (
		\reg2_reg[5]/NET0131 ,
		_w925_,
		_w1813_,
		_w1814_,
		_w2238_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		_w904_,
		_w2238_,
		_w2239_
	);
	LUT4 #(
		.INIT('hc535)
	) name2025 (
		\reg2_reg[5]/NET0131 ,
		_w725_,
		_w925_,
		_w1817_,
		_w2240_
	);
	LUT4 #(
		.INIT('hc808)
	) name2026 (
		\reg2_reg[5]/NET0131 ,
		_w791_,
		_w925_,
		_w1819_,
		_w2241_
	);
	LUT4 #(
		.INIT('h9500)
	) name2027 (
		_w566_,
		_w558_,
		_w860_,
		_w925_,
		_w2242_
	);
	LUT3 #(
		.INIT('ha8)
	) name2028 (
		_w878_,
		_w2237_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('ha8)
	) name2029 (
		\reg2_reg[5]/NET0131 ,
		_w909_,
		_w932_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		_w566_,
		_w905_,
		_w2245_
	);
	LUT4 #(
		.INIT('h0200)
	) name2031 (
		_w248_,
		_w268_,
		_w272_,
		_w645_,
		_w2246_
	);
	LUT3 #(
		.INIT('h07)
	) name2032 (
		_w925_,
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		_w2244_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name2034 (
		_w2243_,
		_w2248_,
		_w2249_
	);
	LUT4 #(
		.INIT('h3100)
	) name2035 (
		_w858_,
		_w2241_,
		_w2240_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h1311)
	) name2036 (
		_w918_,
		_w2236_,
		_w2239_,
		_w2250_,
		_w2251_
	);
	LUT3 #(
		.INIT('hce)
	) name2037 (
		\state_reg[0]/NET0131 ,
		_w2235_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		\reg0_reg[17]/NET0131 ,
		_w942_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		\reg0_reg[17]/NET0131 ,
		_w919_,
		_w2254_
	);
	LUT4 #(
		.INIT('hc808)
	) name2040 (
		\reg0_reg[17]/NET0131 ,
		_w904_,
		_w1057_,
		_w1778_,
		_w2255_
	);
	LUT3 #(
		.INIT('ha2)
	) name2041 (
		\reg0_reg[17]/NET0131 ,
		_w1063_,
		_w1065_,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w433_,
		_w905_,
		_w2257_
	);
	LUT4 #(
		.INIT('h9500)
	) name2043 (
		_w433_,
		_w866_,
		_w867_,
		_w878_,
		_w2258_
	);
	LUT4 #(
		.INIT('h1113)
	) name2044 (
		_w1057_,
		_w2256_,
		_w2257_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w2255_,
		_w2259_,
		_w2260_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2046 (
		\reg0_reg[17]/NET0131 ,
		_w791_,
		_w1057_,
		_w1786_,
		_w2261_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2047 (
		\reg0_reg[17]/NET0131 ,
		_w728_,
		_w1057_,
		_w1788_,
		_w2262_
	);
	LUT3 #(
		.INIT('h31)
	) name2048 (
		_w858_,
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h3111)
	) name2049 (
		_w918_,
		_w2254_,
		_w2260_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('hce)
	) name2050 (
		\state_reg[0]/NET0131 ,
		_w2253_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\reg0_reg[1]/NET0131 ,
		_w942_,
		_w2266_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		\reg0_reg[1]/NET0131 ,
		_w919_,
		_w2267_
	);
	LUT4 #(
		.INIT('haa02)
	) name2053 (
		\reg0_reg[1]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2268_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2054 (
		_w595_,
		_w597_,
		_w756_,
		_w1057_,
		_w2269_
	);
	LUT3 #(
		.INIT('ha8)
	) name2055 (
		_w791_,
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2056 (
		\reg0_reg[1]/NET0131 ,
		_w1057_,
		_w2088_,
		_w2089_,
		_w2271_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2057 (
		\reg0_reg[1]/NET0131 ,
		_w756_,
		_w815_,
		_w1057_,
		_w2272_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		_w858_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h0054)
	) name2059 (
		_w590_,
		_w772_,
		_w778_,
		_w780_,
		_w2274_
	);
	LUT3 #(
		.INIT('ha8)
	) name2060 (
		_w905_,
		_w2268_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		\reg0_reg[1]/NET0131 ,
		_w1063_,
		_w2276_
	);
	LUT4 #(
		.INIT('hc808)
	) name2062 (
		\reg0_reg[1]/NET0131 ,
		_w878_,
		_w1057_,
		_w2092_,
		_w2277_
	);
	LUT3 #(
		.INIT('h01)
	) name2063 (
		_w2276_,
		_w2277_,
		_w2275_,
		_w2278_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2064 (
		_w904_,
		_w2271_,
		_w2273_,
		_w2278_,
		_w2279_
	);
	LUT4 #(
		.INIT('h1311)
	) name2065 (
		_w918_,
		_w2267_,
		_w2270_,
		_w2279_,
		_w2280_
	);
	LUT3 #(
		.INIT('hce)
	) name2066 (
		\state_reg[0]/NET0131 ,
		_w2266_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('haa02)
	) name2067 (
		\reg0_reg[21]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2282_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2068 (
		_w1578_,
		_w2217_,
		_w2218_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name2069 (
		_w904_,
		_w2283_,
		_w2284_
	);
	LUT3 #(
		.INIT('h2a)
	) name2070 (
		\reg0_reg[21]/NET0131 ,
		_w1573_,
		_w1575_,
		_w2285_
	);
	LUT3 #(
		.INIT('h48)
	) name2071 (
		_w711_,
		_w791_,
		_w1040_,
		_w2286_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w381_,
		_w905_,
		_w2287_
	);
	LUT4 #(
		.INIT('h9500)
	) name2073 (
		_w381_,
		_w869_,
		_w870_,
		_w878_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2075 (
		_w711_,
		_w858_,
		_w993_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h1311)
	) name2076 (
		_w1578_,
		_w2285_,
		_w2286_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('hb)
	) name2077 (
		_w2284_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		\reg0_reg[22]/NET0131 ,
		_w942_,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		\reg0_reg[22]/NET0131 ,
		_w919_,
		_w2294_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2080 (
		\reg0_reg[22]/NET0131 ,
		_w717_,
		_w1057_,
		_w1852_,
		_w2295_
	);
	LUT4 #(
		.INIT('hc808)
	) name2081 (
		\reg0_reg[22]/NET0131 ,
		_w791_,
		_w1057_,
		_w1857_,
		_w2296_
	);
	LUT4 #(
		.INIT('h7020)
	) name2082 (
		_w277_,
		_w386_,
		_w904_,
		_w1859_,
		_w2297_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		_w363_,
		_w905_,
		_w2298_
	);
	LUT4 #(
		.INIT('h007b)
	) name2084 (
		_w363_,
		_w878_,
		_w1255_,
		_w2298_,
		_w2299_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2085 (
		\reg0_reg[22]/NET0131 ,
		_w1062_,
		_w1063_,
		_w1065_,
		_w2300_
	);
	LUT4 #(
		.INIT('h0075)
	) name2086 (
		_w1057_,
		_w2297_,
		_w2299_,
		_w2300_,
		_w2301_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2087 (
		_w858_,
		_w2295_,
		_w2296_,
		_w2301_,
		_w2302_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2088 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2294_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('he)
	) name2089 (
		_w2293_,
		_w2303_,
		_w2304_
	);
	LUT4 #(
		.INIT('h04cc)
	) name2090 (
		_w277_,
		_w1895_,
		_w2104_,
		_w2105_,
		_w2305_
	);
	LUT2 #(
		.INIT('h2)
	) name2091 (
		\reg0_reg[2]/NET0131 ,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2092 (
		_w574_,
		_w590_,
		_w597_,
		_w878_,
		_w2307_
	);
	LUT2 #(
		.INIT('h4)
	) name2093 (
		_w574_,
		_w905_,
		_w2308_
	);
	LUT2 #(
		.INIT('h1)
	) name2094 (
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('h0100)
	) name2095 (
		_w2109_,
		_w2106_,
		_w2112_,
		_w2309_,
		_w2310_
	);
	LUT3 #(
		.INIT('hce)
	) name2096 (
		_w1578_,
		_w2306_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h4)
	) name2097 (
		_w582_,
		_w905_,
		_w2312_
	);
	LUT3 #(
		.INIT('h2a)
	) name2098 (
		\reg0_reg[3]/NET0131 ,
		_w1573_,
		_w1575_,
		_w2313_
	);
	LUT4 #(
		.INIT('hffa2)
	) name2099 (
		_w1578_,
		_w1801_,
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		\reg0_reg[5]/NET0131 ,
		_w942_,
		_w2315_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		\reg0_reg[5]/NET0131 ,
		_w919_,
		_w2316_
	);
	LUT4 #(
		.INIT('haa02)
	) name2102 (
		\reg0_reg[5]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2317_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2103 (
		\reg0_reg[5]/NET0131 ,
		_w1057_,
		_w1813_,
		_w1814_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name2104 (
		_w904_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('hc535)
	) name2105 (
		\reg0_reg[5]/NET0131 ,
		_w725_,
		_w1057_,
		_w1817_,
		_w2320_
	);
	LUT4 #(
		.INIT('hc808)
	) name2106 (
		\reg0_reg[5]/NET0131 ,
		_w791_,
		_w1057_,
		_w1819_,
		_w2321_
	);
	LUT4 #(
		.INIT('h9500)
	) name2107 (
		_w566_,
		_w558_,
		_w860_,
		_w1057_,
		_w2322_
	);
	LUT3 #(
		.INIT('ha8)
	) name2108 (
		_w878_,
		_w2317_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('ha2)
	) name2109 (
		\reg0_reg[5]/NET0131 ,
		_w1063_,
		_w1325_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name2110 (
		_w1057_,
		_w2245_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h4)
	) name2112 (
		_w2323_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h3100)
	) name2113 (
		_w858_,
		_w2321_,
		_w2320_,
		_w2327_,
		_w2328_
	);
	LUT4 #(
		.INIT('h1311)
	) name2114 (
		_w918_,
		_w2316_,
		_w2319_,
		_w2328_,
		_w2329_
	);
	LUT3 #(
		.INIT('hce)
	) name2115 (
		\state_reg[0]/NET0131 ,
		_w2315_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h7020)
	) name2116 (
		_w277_,
		_w480_,
		_w904_,
		_w1761_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name2117 (
		_w474_,
		_w905_,
		_w2332_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT4 #(
		.INIT('h6050)
	) name2119 (
		_w474_,
		_w484_,
		_w1074_,
		_w1208_,
		_w2334_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2120 (
		\reg1_reg[13]/NET0131 ,
		_w878_,
		_w2009_,
		_w2334_,
		_w2335_
	);
	LUT4 #(
		.INIT('hff4c)
	) name2121 (
		_w1759_,
		_w1974_,
		_w2333_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		\reg1_reg[17]/NET0131 ,
		_w942_,
		_w2337_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		\reg1_reg[17]/NET0131 ,
		_w919_,
		_w2338_
	);
	LUT4 #(
		.INIT('hc808)
	) name2124 (
		\reg1_reg[17]/NET0131 ,
		_w904_,
		_w1074_,
		_w1778_,
		_w2339_
	);
	LUT3 #(
		.INIT('ha2)
	) name2125 (
		\reg1_reg[17]/NET0131 ,
		_w1063_,
		_w1078_,
		_w2340_
	);
	LUT4 #(
		.INIT('h0057)
	) name2126 (
		_w1074_,
		_w2257_,
		_w2258_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h4)
	) name2127 (
		_w2339_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2128 (
		\reg1_reg[17]/NET0131 ,
		_w791_,
		_w1074_,
		_w1786_,
		_w2343_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2129 (
		\reg1_reg[17]/NET0131 ,
		_w728_,
		_w1074_,
		_w1788_,
		_w2344_
	);
	LUT3 #(
		.INIT('h31)
	) name2130 (
		_w858_,
		_w2343_,
		_w2344_,
		_w2345_
	);
	LUT4 #(
		.INIT('h3111)
	) name2131 (
		_w918_,
		_w2338_,
		_w2342_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('hce)
	) name2132 (
		\state_reg[0]/NET0131 ,
		_w2337_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		\reg1_reg[1]/NET0131 ,
		_w942_,
		_w2348_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		\reg1_reg[1]/NET0131 ,
		_w919_,
		_w2349_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2135 (
		\reg1_reg[1]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2350_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2136 (
		_w595_,
		_w597_,
		_w756_,
		_w1074_,
		_w2351_
	);
	LUT3 #(
		.INIT('ha8)
	) name2137 (
		_w791_,
		_w2350_,
		_w2351_,
		_w2352_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2138 (
		\reg1_reg[1]/NET0131 ,
		_w1074_,
		_w2088_,
		_w2089_,
		_w2353_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2139 (
		\reg1_reg[1]/NET0131 ,
		_w756_,
		_w815_,
		_w1074_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		_w858_,
		_w2354_,
		_w2355_
	);
	LUT4 #(
		.INIT('h0001)
	) name2141 (
		_w590_,
		_w772_,
		_w778_,
		_w780_,
		_w2356_
	);
	LUT3 #(
		.INIT('ha8)
	) name2142 (
		_w905_,
		_w2350_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		\reg1_reg[1]/NET0131 ,
		_w1063_,
		_w2358_
	);
	LUT4 #(
		.INIT('hc808)
	) name2144 (
		\reg1_reg[1]/NET0131 ,
		_w878_,
		_w1074_,
		_w2092_,
		_w2359_
	);
	LUT3 #(
		.INIT('h01)
	) name2145 (
		_w2358_,
		_w2359_,
		_w2357_,
		_w2360_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2146 (
		_w904_,
		_w2353_,
		_w2355_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h1311)
	) name2147 (
		_w918_,
		_w2349_,
		_w2352_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('hce)
	) name2148 (
		\state_reg[0]/NET0131 ,
		_w2348_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		\reg1_reg[22]/NET0131 ,
		_w942_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		\reg1_reg[22]/NET0131 ,
		_w919_,
		_w2365_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2151 (
		\reg1_reg[22]/NET0131 ,
		_w717_,
		_w1074_,
		_w1852_,
		_w2366_
	);
	LUT4 #(
		.INIT('hc808)
	) name2152 (
		\reg1_reg[22]/NET0131 ,
		_w791_,
		_w1074_,
		_w1857_,
		_w2367_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2153 (
		\reg1_reg[22]/NET0131 ,
		_w1063_,
		_w1077_,
		_w1078_,
		_w2368_
	);
	LUT4 #(
		.INIT('h0075)
	) name2154 (
		_w1074_,
		_w2297_,
		_w2299_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2155 (
		_w858_,
		_w2366_,
		_w2367_,
		_w2369_,
		_w2370_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2156 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2365_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('he)
	) name2157 (
		_w2364_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h2)
	) name2158 (
		\reg1_reg[2]/NET0131 ,
		_w1972_,
		_w2373_
	);
	LUT3 #(
		.INIT('hf2)
	) name2159 (
		_w1974_,
		_w2310_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h2)
	) name2160 (
		\reg0_reg[10]/NET0131 ,
		_w942_,
		_w2375_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		\reg0_reg[10]/NET0131 ,
		_w919_,
		_w2376_
	);
	LUT4 #(
		.INIT('haa02)
	) name2162 (
		\reg0_reg[10]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2377_
	);
	LUT4 #(
		.INIT('hc808)
	) name2163 (
		\reg0_reg[10]/NET0131 ,
		_w904_,
		_w1057_,
		_w2184_,
		_w2378_
	);
	LUT4 #(
		.INIT('h8488)
	) name2164 (
		_w754_,
		_w1057_,
		_w1379_,
		_w1380_,
		_w2379_
	);
	LUT3 #(
		.INIT('ha8)
	) name2165 (
		_w791_,
		_w2377_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2166 (
		\reg0_reg[10]/NET0131 ,
		_w1063_,
		_w1325_,
		_w1572_,
		_w2381_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		_w508_,
		_w905_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w2189_,
		_w2382_,
		_w2383_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2169 (
		_w754_,
		_w858_,
		_w1388_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h31)
	) name2170 (
		_w1057_,
		_w2381_,
		_w2384_,
		_w2385_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2171 (
		_w918_,
		_w2378_,
		_w2380_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('heeec)
	) name2172 (
		\state_reg[0]/NET0131 ,
		_w2375_,
		_w2376_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('h2a)
	) name2173 (
		\reg1_reg[3]/NET0131 ,
		_w2002_,
		_w2004_,
		_w2388_
	);
	LUT4 #(
		.INIT('hffc4)
	) name2174 (
		_w1801_,
		_w1974_,
		_w2312_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name2175 (
		\reg1_reg[5]/NET0131 ,
		_w942_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		\reg1_reg[5]/NET0131 ,
		_w919_,
		_w2391_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2177 (
		\reg1_reg[5]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2392_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2178 (
		\reg1_reg[5]/NET0131 ,
		_w1074_,
		_w1813_,
		_w1814_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name2179 (
		_w904_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('hc535)
	) name2180 (
		\reg1_reg[5]/NET0131 ,
		_w725_,
		_w1074_,
		_w1817_,
		_w2395_
	);
	LUT4 #(
		.INIT('hc808)
	) name2181 (
		\reg1_reg[5]/NET0131 ,
		_w791_,
		_w1074_,
		_w1819_,
		_w2396_
	);
	LUT4 #(
		.INIT('h9500)
	) name2182 (
		_w566_,
		_w558_,
		_w860_,
		_w1074_,
		_w2397_
	);
	LUT3 #(
		.INIT('ha8)
	) name2183 (
		_w878_,
		_w2392_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('ha2)
	) name2184 (
		\reg1_reg[5]/NET0131 ,
		_w1063_,
		_w1603_,
		_w2399_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		_w1074_,
		_w2245_,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name2186 (
		_w2399_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h4)
	) name2187 (
		_w2398_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('h3100)
	) name2188 (
		_w858_,
		_w2396_,
		_w2395_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h1311)
	) name2189 (
		_w918_,
		_w2391_,
		_w2394_,
		_w2403_,
		_w2404_
	);
	LUT3 #(
		.INIT('hce)
	) name2190 (
		\state_reg[0]/NET0131 ,
		_w2390_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('h0200)
	) name2191 (
		_w257_,
		_w268_,
		_w272_,
		_w645_,
		_w2406_
	);
	LUT4 #(
		.INIT('h00d5)
	) name2192 (
		_w925_,
		_w1759_,
		_w2333_,
		_w2406_,
		_w2407_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2193 (
		_w632_,
		_w772_,
		_w778_,
		_w780_,
		_w2408_
	);
	LUT4 #(
		.INIT('h0004)
	) name2194 (
		_w909_,
		_w1110_,
		_w1359_,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		\reg2_reg[13]/NET0131 ,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('hf2)
	) name2196 (
		_w1110_,
		_w2407_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name2197 (
		\reg2_reg[17]/NET0131 ,
		_w942_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		\reg2_reg[17]/NET0131 ,
		_w919_,
		_w2413_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2199 (
		\reg2_reg[17]/NET0131 ,
		_w791_,
		_w925_,
		_w1786_,
		_w2414_
	);
	LUT4 #(
		.INIT('h0400)
	) name2200 (
		_w268_,
		_w427_,
		_w272_,
		_w645_,
		_w2415_
	);
	LUT4 #(
		.INIT('h0057)
	) name2201 (
		\reg2_reg[17]/NET0131 ,
		_w909_,
		_w1359_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h5700)
	) name2202 (
		_w925_,
		_w2257_,
		_w2258_,
		_w2416_,
		_w2417_
	);
	LUT2 #(
		.INIT('h4)
	) name2203 (
		_w2414_,
		_w2417_,
		_w2418_
	);
	LUT4 #(
		.INIT('hc808)
	) name2204 (
		\reg2_reg[17]/NET0131 ,
		_w904_,
		_w925_,
		_w1778_,
		_w2419_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2205 (
		\reg2_reg[17]/NET0131 ,
		_w728_,
		_w925_,
		_w1788_,
		_w2420_
	);
	LUT3 #(
		.INIT('h31)
	) name2206 (
		_w858_,
		_w2419_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('h3111)
	) name2207 (
		_w918_,
		_w2413_,
		_w2418_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('hce)
	) name2208 (
		\state_reg[0]/NET0131 ,
		_w2412_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name2209 (
		\reg2_reg[22]/NET0131 ,
		_w942_,
		_w2424_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		\reg2_reg[22]/NET0131 ,
		_w919_,
		_w2425_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2211 (
		\reg2_reg[22]/NET0131 ,
		_w717_,
		_w925_,
		_w1852_,
		_w2426_
	);
	LUT4 #(
		.INIT('hc808)
	) name2212 (
		\reg2_reg[22]/NET0131 ,
		_w791_,
		_w925_,
		_w1857_,
		_w2427_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2213 (
		\reg2_reg[22]/NET0131 ,
		_w909_,
		_w1358_,
		_w1359_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w365_,
		_w907_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT4 #(
		.INIT('h7500)
	) name2216 (
		_w925_,
		_w2297_,
		_w2299_,
		_w2430_,
		_w2431_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2217 (
		_w858_,
		_w2426_,
		_w2427_,
		_w2431_,
		_w2432_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2218 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2425_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('he)
	) name2219 (
		_w2424_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('h0200)
	) name2220 (
		\reg3_reg[2]/NET0131 ,
		_w268_,
		_w272_,
		_w645_,
		_w2435_
	);
	LUT4 #(
		.INIT('hcc08)
	) name2221 (
		_w925_,
		_w1110_,
		_w2310_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h2a)
	) name2222 (
		\reg2_reg[2]/NET0131 ,
		_w1549_,
		_w2029_,
		_w2437_
	);
	LUT2 #(
		.INIT('he)
	) name2223 (
		_w2436_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2224 (
		_w772_,
		_w778_,
		_w780_,
		_w1402_,
		_w2439_
	);
	LUT4 #(
		.INIT('h0008)
	) name2225 (
		_w1063_,
		_w1110_,
		_w1325_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		\reg0_reg[13]/NET0131 ,
		_w2440_,
		_w2441_
	);
	LUT4 #(
		.INIT('hff2a)
	) name2227 (
		_w1578_,
		_w1759_,
		_w2333_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		\reg2_reg[4]/NET0131 ,
		_w942_,
		_w2443_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		\reg2_reg[4]/NET0131 ,
		_w919_,
		_w2444_
	);
	LUT4 #(
		.INIT('h111d)
	) name2230 (
		\reg2_reg[4]/NET0131 ,
		_w925_,
		_w2127_,
		_w2128_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		_w904_,
		_w2445_,
		_w2446_
	);
	LUT4 #(
		.INIT('hc808)
	) name2232 (
		\reg2_reg[4]/NET0131 ,
		_w791_,
		_w925_,
		_w2131_,
		_w2447_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2233 (
		\reg2_reg[4]/NET0131 ,
		_w858_,
		_w925_,
		_w2133_,
		_w2448_
	);
	LUT4 #(
		.INIT('hc355)
	) name2234 (
		\reg2_reg[4]/NET0131 ,
		_w558_,
		_w860_,
		_w925_,
		_w2449_
	);
	LUT3 #(
		.INIT('ha8)
	) name2235 (
		\reg2_reg[4]/NET0131 ,
		_w909_,
		_w932_,
		_w2450_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w558_,
		_w905_,
		_w2451_
	);
	LUT4 #(
		.INIT('h0400)
	) name2237 (
		_w268_,
		_w559_,
		_w272_,
		_w645_,
		_w2452_
	);
	LUT3 #(
		.INIT('h07)
	) name2238 (
		_w925_,
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2239 (
		_w878_,
		_w2449_,
		_w2450_,
		_w2453_,
		_w2454_
	);
	LUT3 #(
		.INIT('h10)
	) name2240 (
		_w2448_,
		_w2447_,
		_w2454_,
		_w2455_
	);
	LUT4 #(
		.INIT('h1311)
	) name2241 (
		_w918_,
		_w2444_,
		_w2446_,
		_w2455_,
		_w2456_
	);
	LUT3 #(
		.INIT('hce)
	) name2242 (
		\state_reg[0]/NET0131 ,
		_w2443_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		\reg2_reg[6]/NET0131 ,
		_w942_,
		_w2458_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		\reg2_reg[6]/NET0131 ,
		_w919_,
		_w2459_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2245 (
		\reg2_reg[6]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2460_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2246 (
		_w925_,
		_w2154_,
		_w2155_,
		_w2156_,
		_w2461_
	);
	LUT4 #(
		.INIT('hc808)
	) name2247 (
		\reg2_reg[6]/NET0131 ,
		_w878_,
		_w925_,
		_w2147_,
		_w2462_
	);
	LUT3 #(
		.INIT('ha8)
	) name2248 (
		\reg2_reg[6]/NET0131 ,
		_w909_,
		_w932_,
		_w2463_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w540_,
		_w905_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0400)
	) name2250 (
		_w268_,
		_w542_,
		_w272_,
		_w645_,
		_w2465_
	);
	LUT3 #(
		.INIT('h07)
	) name2251 (
		_w925_,
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name2252 (
		_w2463_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h4)
	) name2253 (
		_w2462_,
		_w2467_,
		_w2468_
	);
	LUT4 #(
		.INIT('h5700)
	) name2254 (
		_w904_,
		_w2460_,
		_w2461_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2255 (
		_w695_,
		_w822_,
		_w824_,
		_w925_,
		_w2470_
	);
	LUT3 #(
		.INIT('ha8)
	) name2256 (
		_w858_,
		_w2460_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('h4b00)
	) name2257 (
		_w603_,
		_w606_,
		_w695_,
		_w925_,
		_w2472_
	);
	LUT3 #(
		.INIT('ha8)
	) name2258 (
		_w791_,
		_w2460_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2259 (
		_w918_,
		_w2471_,
		_w2473_,
		_w2469_,
		_w2474_
	);
	LUT4 #(
		.INIT('heeec)
	) name2260 (
		\state_reg[0]/NET0131 ,
		_w2458_,
		_w2459_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h2)
	) name2261 (
		\reg2_reg[8]/NET0131 ,
		_w942_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name2262 (
		\reg2_reg[8]/NET0131 ,
		_w919_,
		_w2477_
	);
	LUT4 #(
		.INIT('hc355)
	) name2263 (
		\reg2_reg[8]/NET0131 ,
		_w610_,
		_w738_,
		_w925_,
		_w2478_
	);
	LUT2 #(
		.INIT('h2)
	) name2264 (
		_w791_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('hc808)
	) name2265 (
		\reg2_reg[8]/NET0131 ,
		_w904_,
		_w925_,
		_w1960_,
		_w2480_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2266 (
		\reg2_reg[8]/NET0131 ,
		_w858_,
		_w925_,
		_w1962_,
		_w2481_
	);
	LUT4 #(
		.INIT('h0400)
	) name2267 (
		_w268_,
		_w520_,
		_w272_,
		_w645_,
		_w2482_
	);
	LUT4 #(
		.INIT('h0057)
	) name2268 (
		\reg2_reg[8]/NET0131 ,
		_w909_,
		_w1359_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('hd0)
	) name2269 (
		_w925_,
		_w1966_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h10)
	) name2270 (
		_w2480_,
		_w2481_,
		_w2484_,
		_w2485_
	);
	LUT4 #(
		.INIT('h1311)
	) name2271 (
		_w918_,
		_w2477_,
		_w2479_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('hce)
	) name2272 (
		\state_reg[0]/NET0131 ,
		_w2476_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name2273 (
		_w512_,
		_w905_,
		_w2488_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2274 (
		_w925_,
		_w1837_,
		_w1840_,
		_w2488_,
		_w2489_
	);
	LUT4 #(
		.INIT('h0400)
	) name2275 (
		_w268_,
		_w513_,
		_w272_,
		_w645_,
		_w2490_
	);
	LUT3 #(
		.INIT('h2a)
	) name2276 (
		\reg2_reg[9]/NET0131 ,
		_w1549_,
		_w2029_,
		_w2491_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2277 (
		_w1110_,
		_w2489_,
		_w2490_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name2278 (
		\reg0_reg[18]/NET0131 ,
		_w1066_,
		_w1574_,
		_w1934_,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w791_,
		_w2200_,
		_w2494_
	);
	LUT4 #(
		.INIT('h4484)
	) name2280 (
		_w689_,
		_w858_,
		_w1508_,
		_w1851_,
		_w2495_
	);
	LUT4 #(
		.INIT('h7020)
	) name2281 (
		_w277_,
		_w429_,
		_w904_,
		_w2202_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name2282 (
		_w417_,
		_w905_,
		_w2497_
	);
	LUT4 #(
		.INIT('h006f)
	) name2283 (
		_w417_,
		_w869_,
		_w878_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h10)
	) name2284 (
		_w2496_,
		_w2495_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('hecee)
	) name2285 (
		_w1578_,
		_w2493_,
		_w2494_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name2286 (
		\reg0_reg[4]/NET0131 ,
		_w942_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		\reg0_reg[4]/NET0131 ,
		_w919_,
		_w2502_
	);
	LUT4 #(
		.INIT('h111d)
	) name2288 (
		\reg0_reg[4]/NET0131 ,
		_w1057_,
		_w2127_,
		_w2128_,
		_w2503_
	);
	LUT2 #(
		.INIT('h2)
	) name2289 (
		_w904_,
		_w2503_,
		_w2504_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2290 (
		\reg0_reg[4]/NET0131 ,
		_w858_,
		_w1057_,
		_w2133_,
		_w2505_
	);
	LUT4 #(
		.INIT('hc808)
	) name2291 (
		\reg0_reg[4]/NET0131 ,
		_w791_,
		_w1057_,
		_w2131_,
		_w2506_
	);
	LUT4 #(
		.INIT('hc355)
	) name2292 (
		\reg0_reg[4]/NET0131 ,
		_w558_,
		_w860_,
		_w1057_,
		_w2507_
	);
	LUT3 #(
		.INIT('ha2)
	) name2293 (
		\reg0_reg[4]/NET0131 ,
		_w1063_,
		_w1325_,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		_w1057_,
		_w2451_,
		_w2509_
	);
	LUT4 #(
		.INIT('h0031)
	) name2295 (
		_w878_,
		_w2508_,
		_w2507_,
		_w2509_,
		_w2510_
	);
	LUT3 #(
		.INIT('h10)
	) name2296 (
		_w2506_,
		_w2505_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('h1311)
	) name2297 (
		_w918_,
		_w2502_,
		_w2504_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('hce)
	) name2298 (
		\state_reg[0]/NET0131 ,
		_w2501_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h2)
	) name2299 (
		\reg0_reg[6]/NET0131 ,
		_w942_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		\reg0_reg[6]/NET0131 ,
		_w919_,
		_w2515_
	);
	LUT4 #(
		.INIT('haa02)
	) name2301 (
		\reg0_reg[6]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2516_
	);
	LUT4 #(
		.INIT('h4b00)
	) name2302 (
		_w603_,
		_w606_,
		_w695_,
		_w1057_,
		_w2517_
	);
	LUT4 #(
		.INIT('hc808)
	) name2303 (
		\reg0_reg[6]/NET0131 ,
		_w878_,
		_w1057_,
		_w2147_,
		_w2518_
	);
	LUT3 #(
		.INIT('ha2)
	) name2304 (
		\reg0_reg[6]/NET0131 ,
		_w1063_,
		_w1325_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		_w1057_,
		_w2464_,
		_w2520_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w2519_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w2518_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('h5700)
	) name2308 (
		_w791_,
		_w2516_,
		_w2517_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2309 (
		_w1057_,
		_w2154_,
		_w2155_,
		_w2156_,
		_w2524_
	);
	LUT3 #(
		.INIT('ha8)
	) name2310 (
		_w904_,
		_w2516_,
		_w2524_,
		_w2525_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2311 (
		_w695_,
		_w822_,
		_w824_,
		_w1057_,
		_w2526_
	);
	LUT3 #(
		.INIT('ha8)
	) name2312 (
		_w858_,
		_w2516_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2313 (
		_w918_,
		_w2525_,
		_w2527_,
		_w2523_,
		_w2528_
	);
	LUT4 #(
		.INIT('heeec)
	) name2314 (
		\state_reg[0]/NET0131 ,
		_w2514_,
		_w2515_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2315 (
		_w1578_,
		_w1837_,
		_w1840_,
		_w2488_,
		_w2530_
	);
	LUT3 #(
		.INIT('h2a)
	) name2316 (
		\reg0_reg[9]/NET0131 ,
		_w1573_,
		_w1575_,
		_w2531_
	);
	LUT2 #(
		.INIT('he)
	) name2317 (
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h2)
	) name2318 (
		\reg1_reg[10]/NET0131 ,
		_w942_,
		_w2533_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		\reg1_reg[10]/NET0131 ,
		_w919_,
		_w2534_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2320 (
		\reg1_reg[10]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2535_
	);
	LUT4 #(
		.INIT('hc808)
	) name2321 (
		\reg1_reg[10]/NET0131 ,
		_w904_,
		_w1074_,
		_w2184_,
		_w2536_
	);
	LUT4 #(
		.INIT('h8488)
	) name2322 (
		_w754_,
		_w1074_,
		_w1379_,
		_w1380_,
		_w2537_
	);
	LUT3 #(
		.INIT('ha8)
	) name2323 (
		_w791_,
		_w2535_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2324 (
		\reg1_reg[10]/NET0131 ,
		_w1063_,
		_w1603_,
		_w2001_,
		_w2539_
	);
	LUT3 #(
		.INIT('h0d)
	) name2325 (
		_w1074_,
		_w2384_,
		_w2539_,
		_w2540_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2326 (
		_w918_,
		_w2536_,
		_w2538_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('heeec)
	) name2327 (
		\state_reg[0]/NET0131 ,
		_w2533_,
		_w2534_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		\reg1_reg[18]/NET0131 ,
		_w942_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		\reg1_reg[18]/NET0131 ,
		_w919_,
		_w2544_
	);
	LUT2 #(
		.INIT('h2)
	) name2330 (
		\reg1_reg[18]/NET0131 ,
		_w1644_,
		_w2545_
	);
	LUT4 #(
		.INIT('h0075)
	) name2331 (
		_w1074_,
		_w2494_,
		_w2499_,
		_w2545_,
		_w2546_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2332 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2544_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('he)
	) name2333 (
		_w2543_,
		_w2547_,
		_w2548_
	);
	LUT3 #(
		.INIT('h2a)
	) name2334 (
		\reg1_reg[21]/NET0131 ,
		_w2002_,
		_w2004_,
		_w2549_
	);
	LUT4 #(
		.INIT('hff8a)
	) name2335 (
		_w1974_,
		_w2286_,
		_w2290_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h2)
	) name2336 (
		\reg1_reg[4]/NET0131 ,
		_w942_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		\reg1_reg[4]/NET0131 ,
		_w919_,
		_w2552_
	);
	LUT4 #(
		.INIT('h111d)
	) name2338 (
		\reg1_reg[4]/NET0131 ,
		_w1074_,
		_w2127_,
		_w2128_,
		_w2553_
	);
	LUT2 #(
		.INIT('h2)
	) name2339 (
		_w904_,
		_w2553_,
		_w2554_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2340 (
		\reg1_reg[4]/NET0131 ,
		_w858_,
		_w1074_,
		_w2133_,
		_w2555_
	);
	LUT4 #(
		.INIT('hc808)
	) name2341 (
		\reg1_reg[4]/NET0131 ,
		_w791_,
		_w1074_,
		_w2131_,
		_w2556_
	);
	LUT4 #(
		.INIT('hc355)
	) name2342 (
		\reg1_reg[4]/NET0131 ,
		_w558_,
		_w860_,
		_w1074_,
		_w2557_
	);
	LUT3 #(
		.INIT('ha2)
	) name2343 (
		\reg1_reg[4]/NET0131 ,
		_w1063_,
		_w1603_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		_w1074_,
		_w2451_,
		_w2559_
	);
	LUT4 #(
		.INIT('h0031)
	) name2345 (
		_w878_,
		_w2558_,
		_w2557_,
		_w2559_,
		_w2560_
	);
	LUT3 #(
		.INIT('h10)
	) name2346 (
		_w2556_,
		_w2555_,
		_w2560_,
		_w2561_
	);
	LUT4 #(
		.INIT('h1311)
	) name2347 (
		_w918_,
		_w2552_,
		_w2554_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('hce)
	) name2348 (
		\state_reg[0]/NET0131 ,
		_w2551_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name2349 (
		\reg1_reg[6]/NET0131 ,
		_w942_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		\reg1_reg[6]/NET0131 ,
		_w919_,
		_w2565_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2351 (
		\reg1_reg[6]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2566_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2352 (
		_w1074_,
		_w2154_,
		_w2155_,
		_w2156_,
		_w2567_
	);
	LUT4 #(
		.INIT('hc808)
	) name2353 (
		\reg1_reg[6]/NET0131 ,
		_w878_,
		_w1074_,
		_w2147_,
		_w2568_
	);
	LUT3 #(
		.INIT('ha2)
	) name2354 (
		\reg1_reg[6]/NET0131 ,
		_w1063_,
		_w1603_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		_w1074_,
		_w2464_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h4)
	) name2357 (
		_w2568_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('h5700)
	) name2358 (
		_w904_,
		_w2566_,
		_w2567_,
		_w2572_,
		_w2573_
	);
	LUT4 #(
		.INIT('h4b00)
	) name2359 (
		_w603_,
		_w606_,
		_w695_,
		_w1074_,
		_w2574_
	);
	LUT3 #(
		.INIT('ha8)
	) name2360 (
		_w791_,
		_w2566_,
		_w2574_,
		_w2575_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2361 (
		_w695_,
		_w822_,
		_w824_,
		_w1074_,
		_w2576_
	);
	LUT3 #(
		.INIT('ha8)
	) name2362 (
		_w858_,
		_w2566_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2363 (
		_w918_,
		_w2575_,
		_w2577_,
		_w2573_,
		_w2578_
	);
	LUT4 #(
		.INIT('heeec)
	) name2364 (
		\state_reg[0]/NET0131 ,
		_w2564_,
		_w2565_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2365 (
		\reg1_reg[8]/NET0131 ,
		_w942_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		\reg1_reg[8]/NET0131 ,
		_w919_,
		_w2581_
	);
	LUT4 #(
		.INIT('hc355)
	) name2367 (
		\reg1_reg[8]/NET0131 ,
		_w610_,
		_w738_,
		_w1074_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2368 (
		_w791_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('hc808)
	) name2369 (
		\reg1_reg[8]/NET0131 ,
		_w904_,
		_w1074_,
		_w1960_,
		_w2584_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2370 (
		\reg1_reg[8]/NET0131 ,
		_w858_,
		_w1074_,
		_w1962_,
		_w2585_
	);
	LUT3 #(
		.INIT('ha2)
	) name2371 (
		\reg1_reg[8]/NET0131 ,
		_w1063_,
		_w1078_,
		_w2586_
	);
	LUT3 #(
		.INIT('h0d)
	) name2372 (
		_w1074_,
		_w1966_,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('h10)
	) name2373 (
		_w2584_,
		_w2585_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('h1311)
	) name2374 (
		_w918_,
		_w2581_,
		_w2583_,
		_w2588_,
		_w2589_
	);
	LUT3 #(
		.INIT('hce)
	) name2375 (
		\state_reg[0]/NET0131 ,
		_w2580_,
		_w2589_,
		_w2590_
	);
	LUT3 #(
		.INIT('h2a)
	) name2376 (
		\reg1_reg[9]/NET0131 ,
		_w2002_,
		_w2004_,
		_w2591_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name2377 (
		_w1837_,
		_w1840_,
		_w1974_,
		_w2488_,
		_w2592_
	);
	LUT2 #(
		.INIT('he)
	) name2378 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h2)
	) name2379 (
		\reg2_reg[10]/NET0131 ,
		_w942_,
		_w2594_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		\reg2_reg[10]/NET0131 ,
		_w919_,
		_w2595_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2381 (
		\reg2_reg[10]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2596_
	);
	LUT4 #(
		.INIT('hc808)
	) name2382 (
		\reg2_reg[10]/NET0131 ,
		_w904_,
		_w925_,
		_w2184_,
		_w2597_
	);
	LUT4 #(
		.INIT('h8488)
	) name2383 (
		_w754_,
		_w925_,
		_w1379_,
		_w1380_,
		_w2598_
	);
	LUT3 #(
		.INIT('ha8)
	) name2384 (
		_w791_,
		_w2596_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h0400)
	) name2385 (
		_w268_,
		_w500_,
		_w272_,
		_w645_,
		_w2600_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2386 (
		\reg2_reg[10]/NET0131 ,
		_w909_,
		_w1359_,
		_w1548_,
		_w2601_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT3 #(
		.INIT('hd0)
	) name2388 (
		_w925_,
		_w2384_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2389 (
		_w918_,
		_w2597_,
		_w2599_,
		_w2603_,
		_w2604_
	);
	LUT4 #(
		.INIT('heeec)
	) name2390 (
		\state_reg[0]/NET0131 ,
		_w2594_,
		_w2595_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name2391 (
		\reg2_reg[18]/NET0131 ,
		_w942_,
		_w2606_
	);
	LUT2 #(
		.INIT('h8)
	) name2392 (
		\reg2_reg[18]/NET0131 ,
		_w919_,
		_w2607_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2393 (
		_w925_,
		_w2496_,
		_w2495_,
		_w2498_,
		_w2608_
	);
	LUT4 #(
		.INIT('h0155)
	) name2394 (
		\reg2_reg[18]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2609_
	);
	LUT2 #(
		.INIT('h2)
	) name2395 (
		_w791_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h0400)
	) name2396 (
		_w268_,
		_w418_,
		_w272_,
		_w645_,
		_w2611_
	);
	LUT3 #(
		.INIT('h0d)
	) name2397 (
		\reg2_reg[18]/NET0131 ,
		_w1550_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2398 (
		_w925_,
		_w2200_,
		_w2610_,
		_w2612_,
		_w2613_
	);
	LUT4 #(
		.INIT('h1311)
	) name2399 (
		_w918_,
		_w2607_,
		_w2608_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('hce)
	) name2400 (
		\state_reg[0]/NET0131 ,
		_w2606_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h2)
	) name2401 (
		\reg2_reg[1]/NET0131 ,
		_w942_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		\reg2_reg[1]/NET0131 ,
		_w919_,
		_w2617_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2403 (
		\reg2_reg[1]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2618_
	);
	LUT4 #(
		.INIT('h2d00)
	) name2404 (
		_w595_,
		_w597_,
		_w756_,
		_w925_,
		_w2619_
	);
	LUT3 #(
		.INIT('ha8)
	) name2405 (
		_w791_,
		_w2618_,
		_w2619_,
		_w2620_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2406 (
		\reg2_reg[1]/NET0131 ,
		_w925_,
		_w2088_,
		_w2089_,
		_w2621_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2407 (
		\reg2_reg[1]/NET0131 ,
		_w756_,
		_w815_,
		_w925_,
		_w2622_
	);
	LUT4 #(
		.INIT('hc808)
	) name2408 (
		\reg2_reg[1]/NET0131 ,
		_w878_,
		_w925_,
		_w2092_,
		_w2623_
	);
	LUT4 #(
		.INIT('h5400)
	) name2409 (
		_w590_,
		_w772_,
		_w778_,
		_w780_,
		_w2624_
	);
	LUT4 #(
		.INIT('h0200)
	) name2410 (
		\reg3_reg[1]/NET0131 ,
		_w268_,
		_w272_,
		_w645_,
		_w2625_
	);
	LUT4 #(
		.INIT('h0080)
	) name2411 (
		\reg2_reg[1]/NET0131 ,
		_w268_,
		_w632_,
		_w762_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		_w2625_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('h5700)
	) name2413 (
		_w905_,
		_w2618_,
		_w2624_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2414 (
		_w858_,
		_w2622_,
		_w2623_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2415 (
		_w904_,
		_w2621_,
		_w2620_,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2416 (
		\state_reg[0]/NET0131 ,
		_w918_,
		_w2617_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('he)
	) name2417 (
		_w2616_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name2418 (
		\reg2_reg[21]/NET0131 ,
		_w942_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		\reg2_reg[21]/NET0131 ,
		_w919_,
		_w2634_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2420 (
		\reg2_reg[21]/NET0131 ,
		_w925_,
		_w2217_,
		_w2218_,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name2421 (
		_w904_,
		_w2635_,
		_w2636_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2422 (
		\reg2_reg[21]/NET0131 ,
		_w711_,
		_w925_,
		_w993_,
		_w2637_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		_w858_,
		_w2637_,
		_w2638_
	);
	LUT4 #(
		.INIT('hc535)
	) name2424 (
		\reg2_reg[21]/NET0131 ,
		_w711_,
		_w925_,
		_w1040_,
		_w2639_
	);
	LUT2 #(
		.INIT('h8)
	) name2425 (
		_w382_,
		_w907_,
		_w2640_
	);
	LUT4 #(
		.INIT('h0057)
	) name2426 (
		\reg2_reg[21]/NET0131 ,
		_w909_,
		_w1359_,
		_w2640_,
		_w2641_
	);
	LUT4 #(
		.INIT('h5700)
	) name2427 (
		_w925_,
		_w2287_,
		_w2288_,
		_w2641_,
		_w2642_
	);
	LUT3 #(
		.INIT('hd0)
	) name2428 (
		_w791_,
		_w2639_,
		_w2642_,
		_w2643_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2429 (
		_w918_,
		_w2636_,
		_w2638_,
		_w2643_,
		_w2644_
	);
	LUT4 #(
		.INIT('heeec)
	) name2430 (
		\state_reg[0]/NET0131 ,
		_w2633_,
		_w2634_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		\reg1_reg[0]/NET0131 ,
		_w942_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		\reg1_reg[0]/NET0131 ,
		_w919_,
		_w2647_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2433 (
		\reg1_reg[0]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2648_
	);
	LUT4 #(
		.INIT('h4100)
	) name2434 (
		_w277_,
		_w587_,
		_w880_,
		_w1074_,
		_w2649_
	);
	LUT3 #(
		.INIT('ha8)
	) name2435 (
		_w904_,
		_w2648_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('h003a)
	) name2436 (
		\reg1_reg[0]/NET0131 ,
		_w735_,
		_w1074_,
		_w1642_,
		_w2651_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		\reg1_reg[0]/NET0131 ,
		_w1063_,
		_w2652_
	);
	LUT4 #(
		.INIT('h0001)
	) name2438 (
		_w597_,
		_w772_,
		_w778_,
		_w780_,
		_w2653_
	);
	LUT4 #(
		.INIT('h2223)
	) name2439 (
		_w1064_,
		_w2652_,
		_w2648_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h4)
	) name2440 (
		_w2651_,
		_w2654_,
		_w2655_
	);
	LUT4 #(
		.INIT('h1311)
	) name2441 (
		_w918_,
		_w2647_,
		_w2650_,
		_w2655_,
		_w2656_
	);
	LUT3 #(
		.INIT('hce)
	) name2442 (
		\state_reg[0]/NET0131 ,
		_w2646_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name2443 (
		\reg2_reg[0]/NET0131 ,
		_w942_,
		_w2658_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		\reg2_reg[0]/NET0131 ,
		_w919_,
		_w2659_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2445 (
		\reg2_reg[0]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2660_
	);
	LUT4 #(
		.INIT('h4100)
	) name2446 (
		_w277_,
		_w587_,
		_w880_,
		_w925_,
		_w2661_
	);
	LUT3 #(
		.INIT('ha8)
	) name2447 (
		_w904_,
		_w2660_,
		_w2661_,
		_w2662_
	);
	LUT4 #(
		.INIT('h003a)
	) name2448 (
		\reg2_reg[0]/NET0131 ,
		_w735_,
		_w925_,
		_w1642_,
		_w2663_
	);
	LUT4 #(
		.INIT('h5400)
	) name2449 (
		_w597_,
		_w772_,
		_w778_,
		_w780_,
		_w2664_
	);
	LUT4 #(
		.INIT('h0200)
	) name2450 (
		\reg3_reg[0]/NET0131 ,
		_w268_,
		_w272_,
		_w645_,
		_w2665_
	);
	LUT4 #(
		.INIT('h0080)
	) name2451 (
		\reg2_reg[0]/NET0131 ,
		_w268_,
		_w632_,
		_w762_,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('hab00)
	) name2453 (
		_w1064_,
		_w2660_,
		_w2664_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h4)
	) name2454 (
		_w2663_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h1311)
	) name2455 (
		_w918_,
		_w2659_,
		_w2662_,
		_w2669_,
		_w2670_
	);
	LUT3 #(
		.INIT('hce)
	) name2456 (
		\state_reg[0]/NET0131 ,
		_w2658_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		\reg0_reg[0]/NET0131 ,
		_w942_,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		\reg0_reg[0]/NET0131 ,
		_w919_,
		_w2673_
	);
	LUT4 #(
		.INIT('haa02)
	) name2459 (
		\reg0_reg[0]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w2674_
	);
	LUT4 #(
		.INIT('h4100)
	) name2460 (
		_w277_,
		_w587_,
		_w880_,
		_w1057_,
		_w2675_
	);
	LUT3 #(
		.INIT('ha8)
	) name2461 (
		_w904_,
		_w2674_,
		_w2675_,
		_w2676_
	);
	LUT4 #(
		.INIT('h0054)
	) name2462 (
		_w597_,
		_w772_,
		_w778_,
		_w780_,
		_w2677_
	);
	LUT3 #(
		.INIT('h54)
	) name2463 (
		_w1064_,
		_w2674_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\reg0_reg[0]/NET0131 ,
		_w1063_,
		_w2679_
	);
	LUT4 #(
		.INIT('h003a)
	) name2465 (
		\reg0_reg[0]/NET0131 ,
		_w735_,
		_w1057_,
		_w1642_,
		_w2680_
	);
	LUT3 #(
		.INIT('h01)
	) name2466 (
		_w2679_,
		_w2680_,
		_w2678_,
		_w2681_
	);
	LUT4 #(
		.INIT('h1311)
	) name2467 (
		_w918_,
		_w2673_,
		_w2676_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('hce)
	) name2468 (
		\state_reg[0]/NET0131 ,
		_w2672_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('ha060)
	) name2469 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w482_,
		_w2684_
	);
	LUT4 #(
		.INIT('h0509)
	) name2470 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w482_,
		_w2685_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2471 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[11]/NET0131 ,
		_w482_,
		_w2686_
	);
	LUT3 #(
		.INIT('h12)
	) name2472 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w552_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		\reg2_reg[6]/NET0131 ,
		_w539_,
		_w2688_
	);
	LUT2 #(
		.INIT('h4)
	) name2474 (
		\reg2_reg[6]/NET0131 ,
		_w539_,
		_w2689_
	);
	LUT3 #(
		.INIT('h48)
	) name2475 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w580_,
		_w2690_
	);
	LUT3 #(
		.INIT('h21)
	) name2476 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w580_,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w2692_
	);
	LUT3 #(
		.INIT('h4d)
	) name2478 (
		\reg2_reg[1]/NET0131 ,
		_w589_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h020b)
	) name2479 (
		\reg2_reg[2]/NET0131 ,
		_w573_,
		_w2691_,
		_w2693_,
		_w2694_
	);
	LUT4 #(
		.INIT('h444d)
	) name2480 (
		\reg2_reg[4]/NET0131 ,
		_w557_,
		_w2690_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h080e)
	) name2481 (
		\reg2_reg[5]/NET0131 ,
		_w565_,
		_w2689_,
		_w2695_,
		_w2696_
	);
	LUT3 #(
		.INIT('h84)
	) name2482 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w552_,
		_w2697_
	);
	LUT3 #(
		.INIT('h48)
	) name2483 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w525_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name2484 (
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT4 #(
		.INIT('hab00)
	) name2485 (
		_w2687_,
		_w2688_,
		_w2696_,
		_w2699_,
		_w2700_
	);
	LUT3 #(
		.INIT('h21)
	) name2486 (
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w505_,
		_w2701_
	);
	LUT3 #(
		.INIT('h21)
	) name2487 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w525_,
		_w2702_
	);
	LUT2 #(
		.INIT('h1)
	) name2488 (
		_w2701_,
		_w2702_,
		_w2703_
	);
	LUT3 #(
		.INIT('h48)
	) name2489 (
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w505_,
		_w2704_
	);
	LUT4 #(
		.INIT('h4448)
	) name2490 (
		\IR_reg[10]/NET0131 ,
		\reg2_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w2704_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h2221)
	) name2492 (
		\IR_reg[10]/NET0131 ,
		\reg2_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2707_
	);
	LUT4 #(
		.INIT('h004f)
	) name2493 (
		_w2700_,
		_w2703_,
		_w2706_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h8)
	) name2494 (
		_w275_,
		_w277_,
		_w2709_
	);
	LUT3 #(
		.INIT('h28)
	) name2495 (
		_w2709_,
		_w2686_,
		_w2708_,
		_w2710_
	);
	LUT4 #(
		.INIT('ha060)
	) name2496 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[11]/NET0131 ,
		_w482_,
		_w2711_
	);
	LUT4 #(
		.INIT('h2221)
	) name2497 (
		\IR_reg[10]/NET0131 ,
		\reg1_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2712_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		\reg1_reg[6]/NET0131 ,
		_w539_,
		_w2713_
	);
	LUT3 #(
		.INIT('h48)
	) name2499 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w580_,
		_w2714_
	);
	LUT3 #(
		.INIT('h21)
	) name2500 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w580_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w2716_
	);
	LUT3 #(
		.INIT('h4d)
	) name2502 (
		\reg1_reg[1]/NET0131 ,
		_w589_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('h020b)
	) name2503 (
		\reg1_reg[2]/NET0131 ,
		_w573_,
		_w2715_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h444d)
	) name2504 (
		\reg1_reg[4]/NET0131 ,
		_w557_,
		_w2714_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h0701)
	) name2505 (
		\reg1_reg[5]/NET0131 ,
		_w565_,
		_w2713_,
		_w2719_,
		_w2720_
	);
	LUT3 #(
		.INIT('h12)
	) name2506 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w552_,
		_w2721_
	);
	LUT2 #(
		.INIT('h4)
	) name2507 (
		\reg1_reg[6]/NET0131 ,
		_w539_,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		_w2721_,
		_w2722_,
		_w2723_
	);
	LUT3 #(
		.INIT('h48)
	) name2509 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w525_,
		_w2724_
	);
	LUT3 #(
		.INIT('h84)
	) name2510 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w552_,
		_w2725_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT3 #(
		.INIT('h21)
	) name2512 (
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w505_,
		_w2727_
	);
	LUT3 #(
		.INIT('h21)
	) name2513 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w525_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2515 (
		_w2720_,
		_w2723_,
		_w2726_,
		_w2729_,
		_w2730_
	);
	LUT3 #(
		.INIT('h48)
	) name2516 (
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w505_,
		_w2731_
	);
	LUT4 #(
		.INIT('h4448)
	) name2517 (
		\IR_reg[10]/NET0131 ,
		\reg1_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w2731_,
		_w2732_,
		_w2733_
	);
	LUT3 #(
		.INIT('h45)
	) name2519 (
		_w2712_,
		_w2730_,
		_w2733_,
		_w2734_
	);
	LUT4 #(
		.INIT('h0509)
	) name2520 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[11]/NET0131 ,
		_w482_,
		_w2735_
	);
	LUT4 #(
		.INIT('h0045)
	) name2521 (
		_w2712_,
		_w2730_,
		_w2733_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h4)
	) name2522 (
		_w275_,
		_w277_,
		_w2737_
	);
	LUT4 #(
		.INIT('h6900)
	) name2523 (
		\reg1_reg[11]/NET0131 ,
		_w492_,
		_w2734_,
		_w2737_,
		_w2738_
	);
	LUT3 #(
		.INIT('hc8)
	) name2524 (
		_w275_,
		_w492_,
		_w919_,
		_w2739_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name2525 (
		\addr[11]_pad ,
		_w275_,
		_w277_,
		_w919_,
		_w2740_
	);
	LUT2 #(
		.INIT('h4)
	) name2526 (
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2527 (
		\state_reg[0]/NET0131 ,
		_w2738_,
		_w2741_,
		_w2710_,
		_w2742_
	);
	LUT2 #(
		.INIT('he)
	) name2528 (
		_w1217_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		\reg2_reg[12]/NET0131 ,
		_w483_,
		_w2744_
	);
	LUT2 #(
		.INIT('h6)
	) name2530 (
		\reg2_reg[12]/NET0131 ,
		_w483_,
		_w2745_
	);
	LUT4 #(
		.INIT('h1117)
	) name2531 (
		\reg2_reg[7]/NET0131 ,
		_w553_,
		_w2688_,
		_w2696_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w2698_,
		_w2704_,
		_w2747_
	);
	LUT4 #(
		.INIT('h0155)
	) name2533 (
		_w2701_,
		_w2702_,
		_w2746_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w2684_,
		_w2705_,
		_w2749_
	);
	LUT4 #(
		.INIT('h1055)
	) name2535 (
		_w2685_,
		_w2707_,
		_w2748_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('h28)
	) name2536 (
		_w2709_,
		_w2745_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		\reg1_reg[12]/NET0131 ,
		_w483_,
		_w2752_
	);
	LUT2 #(
		.INIT('h6)
	) name2538 (
		\reg1_reg[12]/NET0131 ,
		_w483_,
		_w2753_
	);
	LUT4 #(
		.INIT('h888e)
	) name2539 (
		\reg1_reg[7]/NET0131 ,
		_w553_,
		_w2720_,
		_w2722_,
		_w2754_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w2724_,
		_w2731_,
		_w2755_
	);
	LUT4 #(
		.INIT('h1055)
	) name2541 (
		_w2727_,
		_w2728_,
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name2542 (
		_w2732_,
		_w2711_,
		_w2757_
	);
	LUT4 #(
		.INIT('h1033)
	) name2543 (
		_w2712_,
		_w2735_,
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT3 #(
		.INIT('h01)
	) name2544 (
		\addr[12]_pad ,
		_w275_,
		_w919_,
		_w2759_
	);
	LUT4 #(
		.INIT('h3031)
	) name2545 (
		_w275_,
		_w277_,
		_w483_,
		_w919_,
		_w2760_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h00d7)
	) name2547 (
		_w2737_,
		_w2753_,
		_w2758_,
		_w2761_,
		_w2762_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2548 (
		\reg3_reg[12]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2751_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		\reg1_reg[15]/NET0131 ,
		_w469_,
		_w2764_
	);
	LUT4 #(
		.INIT('h0509)
	) name2550 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[13]/NET0131 ,
		_w237_,
		_w2765_
	);
	LUT3 #(
		.INIT('h0e)
	) name2551 (
		\reg1_reg[12]/NET0131 ,
		_w483_,
		_w2765_,
		_w2766_
	);
	LUT3 #(
		.INIT('h07)
	) name2552 (
		\reg1_reg[12]/NET0131 ,
		_w483_,
		_w2711_,
		_w2767_
	);
	LUT4 #(
		.INIT('ha060)
	) name2553 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[13]/NET0131 ,
		_w237_,
		_w2768_
	);
	LUT3 #(
		.INIT('h07)
	) name2554 (
		\reg1_reg[14]/NET0131 ,
		_w461_,
		_w2768_,
		_w2769_
	);
	LUT4 #(
		.INIT('h7300)
	) name2555 (
		_w2736_,
		_w2766_,
		_w2767_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		\reg1_reg[14]/NET0131 ,
		_w461_,
		_w2771_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2557 (
		\reg1_reg[14]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w461_,
		_w469_,
		_w2772_
	);
	LUT3 #(
		.INIT('h10)
	) name2558 (
		_w2764_,
		_w2770_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h6)
	) name2559 (
		\reg1_reg[15]/NET0131 ,
		_w469_,
		_w2774_
	);
	LUT4 #(
		.INIT('h888a)
	) name2560 (
		_w2737_,
		_w2774_,
		_w2770_,
		_w2771_,
		_w2775_
	);
	LUT2 #(
		.INIT('h1)
	) name2561 (
		\reg2_reg[15]/NET0131 ,
		_w469_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name2562 (
		\reg2_reg[15]/NET0131 ,
		_w469_,
		_w2777_
	);
	LUT2 #(
		.INIT('h6)
	) name2563 (
		\reg2_reg[15]/NET0131 ,
		_w469_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		\reg2_reg[14]/NET0131 ,
		_w461_,
		_w2779_
	);
	LUT4 #(
		.INIT('h0509)
	) name2565 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w237_,
		_w2780_
	);
	LUT3 #(
		.INIT('h0e)
	) name2566 (
		\reg2_reg[12]/NET0131 ,
		_w483_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w2685_,
		_w2707_,
		_w2782_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2568 (
		_w2700_,
		_w2703_,
		_w2706_,
		_w2782_,
		_w2783_
	);
	LUT3 #(
		.INIT('h07)
	) name2569 (
		\reg2_reg[12]/NET0131 ,
		_w483_,
		_w2684_,
		_w2784_
	);
	LUT4 #(
		.INIT('ha060)
	) name2570 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w237_,
		_w2785_
	);
	LUT3 #(
		.INIT('h07)
	) name2571 (
		\reg2_reg[14]/NET0131 ,
		_w461_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h7500)
	) name2572 (
		_w2781_,
		_w2783_,
		_w2784_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h8882)
	) name2573 (
		_w2709_,
		_w2778_,
		_w2779_,
		_w2787_,
		_w2788_
	);
	LUT3 #(
		.INIT('h01)
	) name2574 (
		\addr[15]_pad ,
		_w275_,
		_w919_,
		_w2789_
	);
	LUT4 #(
		.INIT('h3031)
	) name2575 (
		_w275_,
		_w277_,
		_w469_,
		_w919_,
		_w2790_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w2789_,
		_w2790_,
		_w2791_
	);
	LUT4 #(
		.INIT('h1011)
	) name2577 (
		_w2788_,
		_w2791_,
		_w2773_,
		_w2775_,
		_w2792_
	);
	LUT3 #(
		.INIT('h2e)
	) name2578 (
		\reg3_reg[15]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		\reg2_reg[17]/NET0131 ,
		_w432_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		\reg2_reg[17]/NET0131 ,
		_w432_,
		_w2795_
	);
	LUT2 #(
		.INIT('h6)
	) name2581 (
		\reg2_reg[17]/NET0131 ,
		_w432_,
		_w2796_
	);
	LUT3 #(
		.INIT('h48)
	) name2582 (
		\IR_reg[16]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w414_,
		_w2797_
	);
	LUT3 #(
		.INIT('h21)
	) name2583 (
		\IR_reg[16]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w414_,
		_w2798_
	);
	LUT2 #(
		.INIT('h1)
	) name2584 (
		_w2776_,
		_w2798_,
		_w2799_
	);
	LUT4 #(
		.INIT('hab00)
	) name2585 (
		_w2777_,
		_w2779_,
		_w2787_,
		_w2799_,
		_w2800_
	);
	LUT4 #(
		.INIT('h2228)
	) name2586 (
		_w2709_,
		_w2796_,
		_w2797_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name2587 (
		\reg1_reg[17]/NET0131 ,
		_w432_,
		_w2802_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		\reg1_reg[17]/NET0131 ,
		_w432_,
		_w2803_
	);
	LUT2 #(
		.INIT('h6)
	) name2589 (
		\reg1_reg[17]/NET0131 ,
		_w432_,
		_w2804_
	);
	LUT3 #(
		.INIT('h21)
	) name2590 (
		\IR_reg[16]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w414_,
		_w2805_
	);
	LUT3 #(
		.INIT('h48)
	) name2591 (
		\IR_reg[16]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w414_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w2764_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h040f)
	) name2593 (
		_w2770_,
		_w2772_,
		_w2805_,
		_w2807_,
		_w2808_
	);
	LUT3 #(
		.INIT('h01)
	) name2594 (
		\addr[17]_pad ,
		_w275_,
		_w919_,
		_w2809_
	);
	LUT4 #(
		.INIT('h3031)
	) name2595 (
		_w275_,
		_w277_,
		_w432_,
		_w919_,
		_w2810_
	);
	LUT2 #(
		.INIT('h4)
	) name2596 (
		_w2809_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h00d7)
	) name2597 (
		_w2737_,
		_w2804_,
		_w2808_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2598 (
		\reg3_reg[17]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2801_,
		_w2812_,
		_w2813_
	);
	LUT3 #(
		.INIT('h01)
	) name2599 (
		\addr[5]_pad ,
		_w275_,
		_w919_,
		_w2814_
	);
	LUT4 #(
		.INIT('h3031)
	) name2600 (
		_w275_,
		_w277_,
		_w565_,
		_w919_,
		_w2815_
	);
	LUT2 #(
		.INIT('h6)
	) name2601 (
		\reg2_reg[5]/NET0131 ,
		_w565_,
		_w2816_
	);
	LUT4 #(
		.INIT('h8008)
	) name2602 (
		_w275_,
		_w277_,
		_w2695_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h6)
	) name2603 (
		\reg1_reg[5]/NET0131 ,
		_w565_,
		_w2818_
	);
	LUT4 #(
		.INIT('h4004)
	) name2604 (
		_w275_,
		_w277_,
		_w2719_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w2817_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2606 (
		\state_reg[0]/NET0131 ,
		_w2814_,
		_w2815_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('he)
	) name2607 (
		_w1829_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h9)
	) name2608 (
		\reg2_reg[6]/NET0131 ,
		_w539_,
		_w2823_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2609 (
		\reg2_reg[5]/NET0131 ,
		_w565_,
		_w2695_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('h0071)
	) name2610 (
		\reg2_reg[5]/NET0131 ,
		_w565_,
		_w2695_,
		_w2823_,
		_w2825_
	);
	LUT3 #(
		.INIT('h02)
	) name2611 (
		_w2709_,
		_w2825_,
		_w2824_,
		_w2826_
	);
	LUT2 #(
		.INIT('h9)
	) name2612 (
		\reg1_reg[6]/NET0131 ,
		_w539_,
		_w2827_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2613 (
		\reg1_reg[5]/NET0131 ,
		_w565_,
		_w2719_,
		_w2827_,
		_w2828_
	);
	LUT4 #(
		.INIT('h0071)
	) name2614 (
		\reg1_reg[5]/NET0131 ,
		_w565_,
		_w2719_,
		_w2827_,
		_w2829_
	);
	LUT3 #(
		.INIT('h02)
	) name2615 (
		_w2737_,
		_w2829_,
		_w2828_,
		_w2830_
	);
	LUT3 #(
		.INIT('hc8)
	) name2616 (
		_w275_,
		_w539_,
		_w919_,
		_w2831_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name2617 (
		\addr[6]_pad ,
		_w275_,
		_w277_,
		_w919_,
		_w2832_
	);
	LUT4 #(
		.INIT('h0045)
	) name2618 (
		_w2830_,
		_w2831_,
		_w2832_,
		_w2826_,
		_w2833_
	);
	LUT3 #(
		.INIT('h2e)
	) name2619 (
		\reg3_reg[6]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h69)
	) name2620 (
		\IR_reg[7]/NET0131 ,
		\reg2_reg[7]/NET0131 ,
		_w552_,
		_w2835_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2621 (
		_w2709_,
		_w2688_,
		_w2696_,
		_w2835_,
		_w2836_
	);
	LUT3 #(
		.INIT('h69)
	) name2622 (
		\IR_reg[7]/NET0131 ,
		\reg1_reg[7]/NET0131 ,
		_w552_,
		_w2837_
	);
	LUT4 #(
		.INIT('he010)
	) name2623 (
		_w2720_,
		_w2722_,
		_w2737_,
		_w2837_,
		_w2838_
	);
	LUT3 #(
		.INIT('h01)
	) name2624 (
		\addr[7]_pad ,
		_w275_,
		_w919_,
		_w2839_
	);
	LUT4 #(
		.INIT('h3031)
	) name2625 (
		_w275_,
		_w277_,
		_w553_,
		_w919_,
		_w2840_
	);
	LUT4 #(
		.INIT('h0045)
	) name2626 (
		_w2838_,
		_w2839_,
		_w2840_,
		_w2836_,
		_w2841_
	);
	LUT3 #(
		.INIT('h2e)
	) name2627 (
		\reg3_reg[7]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2841_,
		_w2842_
	);
	LUT3 #(
		.INIT('h96)
	) name2628 (
		\IR_reg[8]/NET0131 ,
		\reg2_reg[8]/NET0131 ,
		_w525_,
		_w2843_
	);
	LUT3 #(
		.INIT('h82)
	) name2629 (
		_w2709_,
		_w2746_,
		_w2843_,
		_w2844_
	);
	LUT3 #(
		.INIT('h01)
	) name2630 (
		\addr[8]_pad ,
		_w275_,
		_w919_,
		_w2845_
	);
	LUT4 #(
		.INIT('h3031)
	) name2631 (
		_w275_,
		_w277_,
		_w526_,
		_w919_,
		_w2846_
	);
	LUT2 #(
		.INIT('h4)
	) name2632 (
		_w2845_,
		_w2846_,
		_w2847_
	);
	LUT3 #(
		.INIT('h96)
	) name2633 (
		\IR_reg[8]/NET0131 ,
		\reg1_reg[8]/NET0131 ,
		_w525_,
		_w2848_
	);
	LUT3 #(
		.INIT('h28)
	) name2634 (
		_w2737_,
		_w2754_,
		_w2848_,
		_w2849_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2635 (
		\state_reg[0]/NET0131 ,
		_w2847_,
		_w2849_,
		_w2844_,
		_w2850_
	);
	LUT2 #(
		.INIT('he)
	) name2636 (
		_w2177_,
		_w2850_,
		_w2851_
	);
	LUT3 #(
		.INIT('h96)
	) name2637 (
		\IR_reg[9]/NET0131 ,
		\reg2_reg[9]/NET0131 ,
		_w505_,
		_w2852_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w2698_,
		_w2852_,
		_w2853_
	);
	LUT3 #(
		.INIT('he0)
	) name2639 (
		_w2702_,
		_w2746_,
		_w2853_,
		_w2854_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2640 (
		_w2709_,
		_w2700_,
		_w2703_,
		_w2704_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name2641 (
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name2642 (
		_w2730_,
		_w2731_,
		_w2857_
	);
	LUT3 #(
		.INIT('h96)
	) name2643 (
		\IR_reg[9]/NET0131 ,
		\reg1_reg[9]/NET0131 ,
		_w505_,
		_w2858_
	);
	LUT4 #(
		.INIT('h004f)
	) name2644 (
		_w2720_,
		_w2723_,
		_w2726_,
		_w2728_,
		_w2859_
	);
	LUT3 #(
		.INIT('ha8)
	) name2645 (
		_w2737_,
		_w2858_,
		_w2859_,
		_w2860_
	);
	LUT3 #(
		.INIT('hc8)
	) name2646 (
		_w275_,
		_w511_,
		_w919_,
		_w2861_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name2647 (
		\addr[9]_pad ,
		_w275_,
		_w277_,
		_w919_,
		_w2862_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w2861_,
		_w2862_,
		_w2863_
	);
	LUT3 #(
		.INIT('h0b)
	) name2649 (
		_w2857_,
		_w2860_,
		_w2863_,
		_w2864_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2650 (
		\reg3_reg[9]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2856_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h6)
	) name2651 (
		\reg2_reg[14]/NET0131 ,
		_w461_,
		_w2866_
	);
	LUT4 #(
		.INIT('h173f)
	) name2652 (
		\reg2_reg[12]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w473_,
		_w483_,
		_w2867_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2653 (
		_w2750_,
		_w2781_,
		_w2866_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h0700)
	) name2654 (
		_w2750_,
		_w2781_,
		_w2866_,
		_w2867_,
		_w2869_
	);
	LUT3 #(
		.INIT('h02)
	) name2655 (
		_w2709_,
		_w2869_,
		_w2868_,
		_w2870_
	);
	LUT2 #(
		.INIT('h6)
	) name2656 (
		\reg1_reg[14]/NET0131 ,
		_w461_,
		_w2871_
	);
	LUT4 #(
		.INIT('h173f)
	) name2657 (
		\reg1_reg[12]/NET0131 ,
		\reg1_reg[13]/NET0131 ,
		_w473_,
		_w483_,
		_w2872_
	);
	LUT3 #(
		.INIT('h70)
	) name2658 (
		_w2758_,
		_w2766_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('h01)
	) name2659 (
		\addr[14]_pad ,
		_w275_,
		_w919_,
		_w2874_
	);
	LUT4 #(
		.INIT('h3031)
	) name2660 (
		_w275_,
		_w277_,
		_w461_,
		_w919_,
		_w2875_
	);
	LUT2 #(
		.INIT('h4)
	) name2661 (
		_w2874_,
		_w2875_,
		_w2876_
	);
	LUT4 #(
		.INIT('h007d)
	) name2662 (
		_w2737_,
		_w2871_,
		_w2873_,
		_w2876_,
		_w2877_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2663 (
		\reg3_reg[14]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2870_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h9996)
	) name2664 (
		\IR_reg[10]/NET0131 ,
		\reg2_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2879_
	);
	LUT3 #(
		.INIT('h28)
	) name2665 (
		_w2709_,
		_w2748_,
		_w2879_,
		_w2880_
	);
	LUT3 #(
		.INIT('h01)
	) name2666 (
		\addr[10]_pad ,
		_w275_,
		_w919_,
		_w2881_
	);
	LUT4 #(
		.INIT('h3031)
	) name2667 (
		_w275_,
		_w277_,
		_w507_,
		_w919_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name2668 (
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h9996)
	) name2669 (
		\IR_reg[10]/NET0131 ,
		\reg1_reg[10]/NET0131 ,
		_w505_,
		_w506_,
		_w2884_
	);
	LUT4 #(
		.INIT('h0d07)
	) name2670 (
		_w2737_,
		_w2756_,
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2671 (
		\reg3_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2880_,
		_w2885_,
		_w2886_
	);
	LUT4 #(
		.INIT('h008c)
	) name2672 (
		_w2736_,
		_w2766_,
		_w2767_,
		_w2768_,
		_w2887_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2673 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[13]/NET0131 ,
		_w237_,
		_w2888_
	);
	LUT4 #(
		.INIT('h00dc)
	) name2674 (
		_w2736_,
		_w2752_,
		_w2767_,
		_w2888_,
		_w2889_
	);
	LUT3 #(
		.INIT('h02)
	) name2675 (
		_w2737_,
		_w2889_,
		_w2887_,
		_w2890_
	);
	LUT4 #(
		.INIT('h008a)
	) name2676 (
		_w2781_,
		_w2783_,
		_w2784_,
		_w2785_,
		_w2891_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2677 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[13]/NET0131 ,
		_w237_,
		_w2892_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2678 (
		_w2744_,
		_w2783_,
		_w2784_,
		_w2892_,
		_w2893_
	);
	LUT3 #(
		.INIT('h01)
	) name2679 (
		\addr[13]_pad ,
		_w275_,
		_w919_,
		_w2894_
	);
	LUT4 #(
		.INIT('h3031)
	) name2680 (
		_w275_,
		_w277_,
		_w473_,
		_w919_,
		_w2895_
	);
	LUT2 #(
		.INIT('h4)
	) name2681 (
		_w2894_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2682 (
		_w2709_,
		_w2893_,
		_w2891_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2683 (
		\reg3_reg[13]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2890_,
		_w2897_,
		_w2898_
	);
	LUT4 #(
		.INIT('h4448)
	) name2684 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2899_
	);
	LUT4 #(
		.INIT('h2221)
	) name2685 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2900_
	);
	LUT4 #(
		.INIT('h9996)
	) name2686 (
		\IR_reg[18]/NET0131 ,
		\reg2_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2901_
	);
	LUT4 #(
		.INIT('h2033)
	) name2687 (
		_w2750_,
		_w2779_,
		_w2781_,
		_w2867_,
		_w2902_
	);
	LUT4 #(
		.INIT('h135f)
	) name2688 (
		\reg2_reg[14]/NET0131 ,
		\reg2_reg[15]/NET0131 ,
		_w461_,
		_w469_,
		_w2903_
	);
	LUT4 #(
		.INIT('h1011)
	) name2689 (
		_w2776_,
		_w2798_,
		_w2902_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w2795_,
		_w2797_,
		_w2905_
	);
	LUT4 #(
		.INIT('h4044)
	) name2691 (
		_w2794_,
		_w2901_,
		_w2904_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('h2322)
	) name2692 (
		_w2794_,
		_w2901_,
		_w2904_,
		_w2905_,
		_w2907_
	);
	LUT3 #(
		.INIT('h02)
	) name2693 (
		_w2709_,
		_w2907_,
		_w2906_,
		_w2908_
	);
	LUT4 #(
		.INIT('h4448)
	) name2694 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2909_
	);
	LUT4 #(
		.INIT('h2221)
	) name2695 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2910_
	);
	LUT4 #(
		.INIT('h9996)
	) name2696 (
		\IR_reg[18]/NET0131 ,
		\reg1_reg[18]/NET0131 ,
		_w414_,
		_w415_,
		_w2911_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2697 (
		_w2758_,
		_w2766_,
		_w2772_,
		_w2872_,
		_w2912_
	);
	LUT4 #(
		.INIT('h137f)
	) name2698 (
		\reg1_reg[14]/NET0131 ,
		\reg1_reg[15]/NET0131 ,
		_w461_,
		_w469_,
		_w2913_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w2803_,
		_w2806_,
		_w2914_
	);
	LUT4 #(
		.INIT('hba00)
	) name2700 (
		_w2805_,
		_w2912_,
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('ha082)
	) name2701 (
		_w2737_,
		_w2802_,
		_w2911_,
		_w2915_,
		_w2916_
	);
	LUT3 #(
		.INIT('h01)
	) name2702 (
		\addr[18]_pad ,
		_w275_,
		_w919_,
		_w2917_
	);
	LUT4 #(
		.INIT('h3031)
	) name2703 (
		_w275_,
		_w277_,
		_w416_,
		_w919_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name2704 (
		_w2917_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name2705 (
		_w2916_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2706 (
		\reg3_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2908_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w2802_,
		_w2910_,
		_w2922_
	);
	LUT4 #(
		.INIT('h010f)
	) name2708 (
		_w2803_,
		_w2808_,
		_w2909_,
		_w2922_,
		_w2923_
	);
	LUT4 #(
		.INIT('h6090)
	) name2709 (
		\reg1_reg[19]/NET0131 ,
		_w405_,
		_w2737_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w2794_,
		_w2900_,
		_w2925_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2711 (
		_w2795_,
		_w2797_,
		_w2800_,
		_w2925_,
		_w2926_
	);
	LUT3 #(
		.INIT('h96)
	) name2712 (
		\IR_reg[19]/NET0131 ,
		\reg2_reg[19]/NET0131 ,
		_w264_,
		_w2927_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2713 (
		_w2709_,
		_w2899_,
		_w2926_,
		_w2927_,
		_w2928_
	);
	LUT3 #(
		.INIT('h01)
	) name2714 (
		\addr[19]_pad ,
		_w275_,
		_w919_,
		_w2929_
	);
	LUT4 #(
		.INIT('h3031)
	) name2715 (
		_w275_,
		_w277_,
		_w405_,
		_w919_,
		_w2930_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		_w2929_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2717 (
		\state_reg[0]/NET0131 ,
		_w2928_,
		_w2931_,
		_w2924_,
		_w2932_
	);
	LUT2 #(
		.INIT('he)
	) name2718 (
		_w1451_,
		_w2932_,
		_w2933_
	);
	LUT3 #(
		.INIT('h96)
	) name2719 (
		\IR_reg[16]/NET0131 ,
		\reg2_reg[16]/NET0131 ,
		_w414_,
		_w2934_
	);
	LUT4 #(
		.INIT('h4500)
	) name2720 (
		_w2776_,
		_w2902_,
		_w2903_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('h00ba)
	) name2721 (
		_w2776_,
		_w2902_,
		_w2903_,
		_w2934_,
		_w2936_
	);
	LUT3 #(
		.INIT('h02)
	) name2722 (
		_w2709_,
		_w2936_,
		_w2935_,
		_w2937_
	);
	LUT3 #(
		.INIT('h01)
	) name2723 (
		\addr[16]_pad ,
		_w275_,
		_w919_,
		_w2938_
	);
	LUT4 #(
		.INIT('h3031)
	) name2724 (
		_w275_,
		_w277_,
		_w435_,
		_w919_,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name2725 (
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h96)
	) name2726 (
		\IR_reg[16]/NET0131 ,
		\reg1_reg[16]/NET0131 ,
		_w414_,
		_w2941_
	);
	LUT4 #(
		.INIT('h208a)
	) name2727 (
		_w2737_,
		_w2912_,
		_w2913_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h1)
	) name2728 (
		_w2940_,
		_w2942_,
		_w2943_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2729 (
		\reg3_reg[16]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2937_,
		_w2943_,
		_w2944_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2730 (
		\addr[1]_pad ,
		_w278_,
		_w589_,
		_w919_,
		_w2945_
	);
	LUT4 #(
		.INIT('h936c)
	) name2731 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg2_reg[1]/NET0131 ,
		_w2946_
	);
	LUT2 #(
		.INIT('h6)
	) name2732 (
		_w2692_,
		_w2946_,
		_w2947_
	);
	LUT3 #(
		.INIT('h80)
	) name2733 (
		_w275_,
		_w277_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('h936c)
	) name2734 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\reg1_reg[1]/NET0131 ,
		_w2949_
	);
	LUT2 #(
		.INIT('h6)
	) name2735 (
		_w2716_,
		_w2949_,
		_w2950_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name2736 (
		_w275_,
		_w277_,
		_w589_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w2948_,
		_w2951_,
		_w2952_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2738 (
		\reg3_reg[1]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2945_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2739 (
		\addr[2]_pad ,
		_w278_,
		_w573_,
		_w919_,
		_w2954_
	);
	LUT2 #(
		.INIT('h9)
	) name2740 (
		\reg1_reg[2]/NET0131 ,
		_w573_,
		_w2955_
	);
	LUT2 #(
		.INIT('h9)
	) name2741 (
		_w2717_,
		_w2955_,
		_w2956_
	);
	LUT3 #(
		.INIT('h40)
	) name2742 (
		_w275_,
		_w277_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('h9)
	) name2743 (
		\reg2_reg[2]/NET0131 ,
		_w573_,
		_w2958_
	);
	LUT2 #(
		.INIT('h9)
	) name2744 (
		_w2693_,
		_w2958_,
		_w2959_
	);
	LUT4 #(
		.INIT('h75fd)
	) name2745 (
		_w275_,
		_w277_,
		_w573_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h4)
	) name2746 (
		_w2957_,
		_w2960_,
		_w2961_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2747 (
		\reg3_reg[2]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2954_,
		_w2961_,
		_w2962_
	);
	LUT4 #(
		.INIT('hc088)
	) name2748 (
		\addr[3]_pad ,
		_w278_,
		_w581_,
		_w919_,
		_w2963_
	);
	LUT3 #(
		.INIT('h96)
	) name2749 (
		\IR_reg[3]/NET0131 ,
		\reg2_reg[3]/NET0131 ,
		_w580_,
		_w2964_
	);
	LUT4 #(
		.INIT('hd42b)
	) name2750 (
		\reg2_reg[2]/NET0131 ,
		_w573_,
		_w2693_,
		_w2964_,
		_w2965_
	);
	LUT3 #(
		.INIT('h80)
	) name2751 (
		_w275_,
		_w277_,
		_w2965_,
		_w2966_
	);
	LUT3 #(
		.INIT('h96)
	) name2752 (
		\IR_reg[3]/NET0131 ,
		\reg1_reg[3]/NET0131 ,
		_w580_,
		_w2967_
	);
	LUT4 #(
		.INIT('hd42b)
	) name2753 (
		\reg1_reg[2]/NET0131 ,
		_w573_,
		_w2717_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name2754 (
		_w275_,
		_w277_,
		_w581_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w2966_,
		_w2969_,
		_w2970_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2756 (
		\reg3_reg[3]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2963_,
		_w2970_,
		_w2971_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2757 (
		\addr[4]_pad ,
		_w278_,
		_w557_,
		_w919_,
		_w2972_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2758 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\reg2_reg[4]/NET0131 ,
		_w217_,
		_w2973_
	);
	LUT3 #(
		.INIT('he0)
	) name2759 (
		_w2690_,
		_w2694_,
		_w2973_,
		_w2974_
	);
	LUT3 #(
		.INIT('h01)
	) name2760 (
		_w2690_,
		_w2694_,
		_w2973_,
		_w2975_
	);
	LUT4 #(
		.INIT('h0008)
	) name2761 (
		_w275_,
		_w277_,
		_w2975_,
		_w2974_,
		_w2976_
	);
	LUT3 #(
		.INIT('h02)
	) name2762 (
		_w275_,
		_w277_,
		_w557_,
		_w2977_
	);
	LUT4 #(
		.INIT('h3c96)
	) name2763 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\reg1_reg[4]/NET0131 ,
		_w217_,
		_w2978_
	);
	LUT3 #(
		.INIT('he0)
	) name2764 (
		_w2714_,
		_w2718_,
		_w2978_,
		_w2979_
	);
	LUT3 #(
		.INIT('h01)
	) name2765 (
		_w2714_,
		_w2718_,
		_w2978_,
		_w2980_
	);
	LUT4 #(
		.INIT('h0004)
	) name2766 (
		_w275_,
		_w277_,
		_w2980_,
		_w2979_,
		_w2981_
	);
	LUT3 #(
		.INIT('h01)
	) name2767 (
		_w2977_,
		_w2981_,
		_w2976_,
		_w2982_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2768 (
		\reg3_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2972_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name2769 (
		\IR_reg[0]/NET0131 ,
		\addr[0]_pad ,
		_w278_,
		_w919_,
		_w2984_
	);
	LUT2 #(
		.INIT('h6)
	) name2770 (
		\IR_reg[0]/NET0131 ,
		\reg2_reg[0]/NET0131 ,
		_w2985_
	);
	LUT3 #(
		.INIT('h80)
	) name2771 (
		_w275_,
		_w277_,
		_w2985_,
		_w2986_
	);
	LUT4 #(
		.INIT('hf95f)
	) name2772 (
		\IR_reg[0]/NET0131 ,
		\reg1_reg[0]/NET0131 ,
		_w275_,
		_w277_,
		_w2987_
	);
	LUT2 #(
		.INIT('h4)
	) name2773 (
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('he2ee)
	) name2774 (
		\reg3_reg[0]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2984_,
		_w2988_,
		_w2989_
	);
	LUT3 #(
		.INIT('h57)
	) name2775 (
		\state_reg[0]/NET0131 ,
		_w278_,
		_w919_,
		_w2990_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		\state_reg[0]/NET0131 ,
		_w919_,
		_w2991_
	);
	LUT4 #(
		.INIT('ha060)
	) name2777 (
		\IR_reg[27]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w274_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name2778 (
		\datai[27]_pad ,
		\state_reg[0]/NET0131 ,
		_w2993_
	);
	LUT2 #(
		.INIT('he)
	) name2779 (
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h4448)
	) name2780 (
		\IR_reg[30]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w223_,
		_w233_,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name2781 (
		\datai[30]_pad ,
		\state_reg[0]/NET0131 ,
		_w2996_
	);
	LUT2 #(
		.INIT('he)
	) name2782 (
		_w2995_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h2)
	) name2783 (
		\datai[31]_pad ,
		\state_reg[0]/NET0131 ,
		_w2998_
	);
	LUT3 #(
		.INIT('h40)
	) name2784 (
		\IR_reg[30]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name2785 (
		_w231_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('hec)
	) name2786 (
		_w274_,
		_w2998_,
		_w3000_,
		_w3001_
	);
	LUT3 #(
		.INIT('he2)
	) name2787 (
		\datai[29]_pad ,
		\state_reg[0]/NET0131 ,
		_w243_,
		_w3002_
	);
	LUT4 #(
		.INIT('h4448)
	) name2788 (
		\IR_reg[28]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w271_,
		_w276_,
		_w3003_
	);
	LUT2 #(
		.INIT('h2)
	) name2789 (
		\datai[28]_pad ,
		\state_reg[0]/NET0131 ,
		_w3004_
	);
	LUT2 #(
		.INIT('he)
	) name2790 (
		_w3003_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2791 (
		\IR_reg[19]/NET0131 ,
		\datai[19]_pad ,
		\state_reg[0]/NET0131 ,
		_w264_,
		_w3006_
	);
	LUT4 #(
		.INIT('h4448)
	) name2792 (
		\IR_reg[22]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w271_,
		_w631_,
		_w3007_
	);
	LUT2 #(
		.INIT('h2)
	) name2793 (
		\datai[22]_pad ,
		\state_reg[0]/NET0131 ,
		_w3008_
	);
	LUT2 #(
		.INIT('he)
	) name2794 (
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT3 #(
		.INIT('he2)
	) name2795 (
		\datai[21]_pad ,
		\state_reg[0]/NET0131 ,
		_w630_,
		_w3010_
	);
	LUT3 #(
		.INIT('he2)
	) name2796 (
		\datai[17]_pad ,
		\state_reg[0]/NET0131 ,
		_w432_,
		_w3011_
	);
	LUT2 #(
		.INIT('h2)
	) name2797 (
		\datai[23]_pad ,
		\state_reg[0]/NET0131 ,
		_w3012_
	);
	LUT2 #(
		.INIT('he)
	) name2798 (
		_w269_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('h4448)
	) name2799 (
		\IR_reg[24]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w271_,
		_w768_,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name2800 (
		\datai[24]_pad ,
		\state_reg[0]/NET0131 ,
		_w3015_
	);
	LUT2 #(
		.INIT('he)
	) name2801 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT3 #(
		.INIT('he2)
	) name2802 (
		\datai[15]_pad ,
		\state_reg[0]/NET0131 ,
		_w469_,
		_w3017_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2803 (
		\IR_reg[20]/NET0131 ,
		\datai[20]_pad ,
		\state_reg[0]/NET0131 ,
		_w271_,
		_w3018_
	);
	LUT4 #(
		.INIT('ha060)
	) name2804 (
		\IR_reg[11]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w482_,
		_w3019_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		\datai[11]_pad ,
		\state_reg[0]/NET0131 ,
		_w3020_
	);
	LUT2 #(
		.INIT('he)
	) name2806 (
		_w3019_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2807 (
		\IR_reg[25]/NET0131 ,
		\datai[25]_pad ,
		\state_reg[0]/NET0131 ,
		_w774_,
		_w3022_
	);
	LUT4 #(
		.INIT('h4448)
	) name2808 (
		\IR_reg[18]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w414_,
		_w415_,
		_w3023_
	);
	LUT2 #(
		.INIT('h2)
	) name2809 (
		\datai[18]_pad ,
		\state_reg[0]/NET0131 ,
		_w3024_
	);
	LUT2 #(
		.INIT('he)
	) name2810 (
		_w3023_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2811 (
		\IR_reg[26]/NET0131 ,
		\datai[26]_pad ,
		\state_reg[0]/NET0131 ,
		_w770_,
		_w3026_
	);
	LUT3 #(
		.INIT('he2)
	) name2812 (
		\datai[14]_pad ,
		\state_reg[0]/NET0131 ,
		_w461_,
		_w3027_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2813 (
		\IR_reg[16]/NET0131 ,
		\datai[16]_pad ,
		\state_reg[0]/NET0131 ,
		_w414_,
		_w3028_
	);
	LUT4 #(
		.INIT('ha060)
	) name2814 (
		\IR_reg[13]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w237_,
		_w3029_
	);
	LUT2 #(
		.INIT('h2)
	) name2815 (
		\datai[13]_pad ,
		\state_reg[0]/NET0131 ,
		_w3030_
	);
	LUT2 #(
		.INIT('he)
	) name2816 (
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('hac5c)
	) name2817 (
		\IR_reg[7]/NET0131 ,
		\datai[7]_pad ,
		\state_reg[0]/NET0131 ,
		_w552_,
		_w3032_
	);
	LUT3 #(
		.INIT('he2)
	) name2818 (
		\datai[12]_pad ,
		\state_reg[0]/NET0131 ,
		_w483_,
		_w3033_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2819 (
		\IR_reg[9]/NET0131 ,
		\datai[9]_pad ,
		\state_reg[0]/NET0131 ,
		_w505_,
		_w3034_
	);
	LUT4 #(
		.INIT('h4448)
	) name2820 (
		\IR_reg[10]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w505_,
		_w506_,
		_w3035_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		\datai[10]_pad ,
		\state_reg[0]/NET0131 ,
		_w3036_
	);
	LUT2 #(
		.INIT('he)
	) name2822 (
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2823 (
		\IR_reg[8]/NET0131 ,
		\datai[8]_pad ,
		\state_reg[0]/NET0131 ,
		_w525_,
		_w3038_
	);
	LUT3 #(
		.INIT('he2)
	) name2824 (
		\datai[5]_pad ,
		\state_reg[0]/NET0131 ,
		_w565_,
		_w3039_
	);
	LUT3 #(
		.INIT('h2e)
	) name2825 (
		\datai[6]_pad ,
		\state_reg[0]/NET0131 ,
		_w539_,
		_w3040_
	);
	LUT4 #(
		.INIT('h5cac)
	) name2826 (
		\IR_reg[3]/NET0131 ,
		\datai[3]_pad ,
		\state_reg[0]/NET0131 ,
		_w580_,
		_w3041_
	);
	LUT4 #(
		.INIT('hc060)
	) name2827 (
		\IR_reg[31]/NET0131 ,
		\IR_reg[4]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w217_,
		_w3042_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		\datai[4]_pad ,
		\state_reg[0]/NET0131 ,
		_w3043_
	);
	LUT2 #(
		.INIT('he)
	) name2829 (
		_w3042_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2830 (
		\IR_reg[0]/NET0131 ,
		\IR_reg[1]/NET0131 ,
		\IR_reg[31]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w3045_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		\datai[1]_pad ,
		\state_reg[0]/NET0131 ,
		_w3046_
	);
	LUT2 #(
		.INIT('he)
	) name2832 (
		_w3045_,
		_w3046_,
		_w3047_
	);
	LUT3 #(
		.INIT('h2e)
	) name2833 (
		\datai[2]_pad ,
		\state_reg[0]/NET0131 ,
		_w573_,
		_w3048_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2834 (
		_w321_,
		_w772_,
		_w778_,
		_w780_,
		_w3049_
	);
	LUT4 #(
		.INIT('h007b)
	) name2835 (
		_w720_,
		_w781_,
		_w1125_,
		_w3049_,
		_w3050_
	);
	LUT4 #(
		.INIT('h8488)
	) name2836 (
		_w720_,
		_w781_,
		_w1134_,
		_w1137_,
		_w3051_
	);
	LUT3 #(
		.INIT('ha8)
	) name2837 (
		_w791_,
		_w3049_,
		_w3051_,
		_w3052_
	);
	LUT4 #(
		.INIT('h7020)
	) name2838 (
		_w277_,
		_w333_,
		_w781_,
		_w1141_,
		_w3053_
	);
	LUT4 #(
		.INIT('h8400)
	) name2839 (
		_w320_,
		_w781_,
		_w876_,
		_w878_,
		_w3054_
	);
	LUT3 #(
		.INIT('ha8)
	) name2840 (
		_w321_,
		_w909_,
		_w1441_,
		_w3055_
	);
	LUT3 #(
		.INIT('ha8)
	) name2841 (
		_w320_,
		_w906_,
		_w907_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w3055_,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('h4)
	) name2843 (
		_w3054_,
		_w3057_,
		_w3058_
	);
	LUT4 #(
		.INIT('h5700)
	) name2844 (
		_w904_,
		_w3049_,
		_w3053_,
		_w3058_,
		_w3059_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2845 (
		_w858_,
		_w3050_,
		_w3052_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('hdd95)
	) name2846 (
		\reg3_reg[27]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w311_,
		_w918_,
		_w3061_
	);
	LUT3 #(
		.INIT('h2f)
	) name2847 (
		_w1110_,
		_w3060_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		\reg3_reg[0]/NET0131 ,
		_w942_,
		_w3063_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		\reg3_reg[0]/NET0131 ,
		_w919_,
		_w3064_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2850 (
		\reg3_reg[0]/NET0131 ,
		_w772_,
		_w778_,
		_w780_,
		_w3065_
	);
	LUT4 #(
		.INIT('h4010)
	) name2851 (
		_w277_,
		_w587_,
		_w781_,
		_w880_,
		_w3066_
	);
	LUT3 #(
		.INIT('ha8)
	) name2852 (
		_w904_,
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('h003a)
	) name2853 (
		\reg3_reg[0]/NET0131 ,
		_w735_,
		_w781_,
		_w1642_,
		_w3068_
	);
	LUT4 #(
		.INIT('h0100)
	) name2854 (
		_w597_,
		_w772_,
		_w778_,
		_w780_,
		_w3069_
	);
	LUT4 #(
		.INIT('h0080)
	) name2855 (
		\reg3_reg[0]/NET0131 ,
		_w268_,
		_w632_,
		_w762_,
		_w3070_
	);
	LUT3 #(
		.INIT('h0b)
	) name2856 (
		_w597_,
		_w907_,
		_w3070_,
		_w3071_
	);
	LUT4 #(
		.INIT('hab00)
	) name2857 (
		_w1064_,
		_w3065_,
		_w3069_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h4)
	) name2858 (
		_w3068_,
		_w3072_,
		_w3073_
	);
	LUT4 #(
		.INIT('h1311)
	) name2859 (
		_w918_,
		_w3064_,
		_w3067_,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('hce)
	) name2860 (
		\state_reg[0]/NET0131 ,
		_w3063_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h0100)
	) name2861 (
		\reg3_reg[3]/NET0131 ,
		_w268_,
		_w272_,
		_w645_,
		_w3076_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2862 (
		_w925_,
		_w1801_,
		_w1803_,
		_w2312_,
		_w3077_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2863 (
		\reg2_reg[3]/NET0131 ,
		_w1358_,
		_w1549_,
		_w2029_,
		_w3078_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2864 (
		_w1110_,
		_w3076_,
		_w3077_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2865 (
		_w337_,
		_w772_,
		_w778_,
		_w780_,
		_w3080_
	);
	LUT4 #(
		.INIT('h8848)
	) name2866 (
		_w682_,
		_w781_,
		_w1046_,
		_w1650_,
		_w3081_
	);
	LUT3 #(
		.INIT('ha8)
	) name2867 (
		_w791_,
		_w3080_,
		_w3081_,
		_w3082_
	);
	LUT4 #(
		.INIT('h4484)
	) name2868 (
		_w682_,
		_w781_,
		_w1000_,
		_w1654_,
		_w3083_
	);
	LUT3 #(
		.INIT('ha8)
	) name2869 (
		_w858_,
		_w3080_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('he020)
	) name2870 (
		_w337_,
		_w781_,
		_w904_,
		_w1657_,
		_w3085_
	);
	LUT3 #(
		.INIT('ha8)
	) name2871 (
		_w337_,
		_w909_,
		_w1441_,
		_w3086_
	);
	LUT3 #(
		.INIT('ha8)
	) name2872 (
		_w336_,
		_w906_,
		_w907_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		_w3086_,
		_w3087_,
		_w3088_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2874 (
		_w781_,
		_w878_,
		_w1659_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h4)
	) name2875 (
		_w3085_,
		_w3089_,
		_w3090_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2876 (
		_w1110_,
		_w3082_,
		_w3084_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('hdd95)
	) name2877 (
		\reg3_reg[25]/NET0131 ,
		\state_reg[0]/NET0131 ,
		_w289_,
		_w918_,
		_w3092_
	);
	LUT2 #(
		.INIT('hb)
	) name2878 (
		_w3091_,
		_w3092_,
		_w3093_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g29_dup/_0_  = _w252_ ;
	assign \g33_dup47063/_0_  = _w261_ ;
	assign \g36117/_0_  = _w767_ ;
	assign \g36132/_0_  = _w924_ ;
	assign \g36133/_0_  = _w944_ ;
	assign \g36134/_0_  = _w1055_ ;
	assign \g36135/_0_  = _w1072_ ;
	assign \g36136/_0_  = _w1084_ ;
	assign \g36153/_0_  = _w1113_ ;
	assign \g36154/_0_  = _w1155_ ;
	assign \g36155/_0_  = _w1168_ ;
	assign \g36156/_0_  = _w1178_ ;
	assign \g36157/_0_  = _w1189_ ;
	assign \g36158/_0_  = _w1199_ ;
	assign \g36186/_0_  = _w1219_ ;
	assign \g36187/_0_  = _w1238_ ;
	assign \g36193/_0_  = _w1267_ ;
	assign \g36197/_0_  = _w1291_ ;
	assign \g36198/_0_  = _w1302_ ;
	assign \g36199/_0_  = _w1316_ ;
	assign \g36200/_0_  = _w1333_ ;
	assign \g36201/_0_  = _w1341_ ;
	assign \g36202/_0_  = _w1352_ ;
	assign \g36203/_0_  = _w1364_ ;
	assign \g36204/_0_  = _w1377_ ;
	assign \g36239/_0_  = _w1409_ ;
	assign \g36240/_0_  = _w1430_ ;
	assign \g36242/_0_  = _w1450_ ;
	assign \g36246/_0_  = _w1468_ ;
	assign \g36255/_0_  = _w1487_ ;
	assign \g36259/_0_  = _w1529_ ;
	assign \g36260/_0_  = _w1539_ ;
	assign \g36261/_0_  = _w1555_ ;
	assign \g36262/_0_  = _w1571_ ;
	assign \g36263/_0_  = _w1579_ ;
	assign \g36264/_0_  = _w1592_ ;
	assign \g36265/_0_  = _w1609_ ;
	assign \g36266/_0_  = _w1624_ ;
	assign \g36267/_0_  = _w1639_ ;
	assign \g36268/_0_  = _w1664_ ;
	assign \g36269/_0_  = _w1680_ ;
	assign \g36270/_0_  = _w1695_ ;
	assign \g36271/_0_  = _w1707_ ;
	assign \g36272/_0_  = _w1723_ ;
	assign \g36273/_0_  = _w1738_ ;
	assign \g36274/_0_  = _w1754_ ;
	assign \g36321/_0_  = _w1774_ ;
	assign \g36322/_0_  = _w1794_ ;
	assign \g36323/_0_  = _w1810_ ;
	assign \g36324/_0_  = _w1831_ ;
	assign \g36325/_0_  = _w1848_ ;
	assign \g36341/_0_  = _w1872_ ;
	assign \g36343/_0_  = _w1877_ ;
	assign \g36344/_0_  = _w1892_ ;
	assign \g36345/_0_  = _w1899_ ;
	assign \g36346/_0_  = _w1914_ ;
	assign \g36347/_0_  = _w1929_ ;
	assign \g36348/_0_  = _w1937_ ;
	assign \g36349/_0_  = _w1939_ ;
	assign \g36350/_0_  = _w1941_ ;
	assign \g36351/_0_  = _w1954_ ;
	assign \g36352/_0_  = _w1970_ ;
	assign \g36353/_0_  = _w1975_ ;
	assign \g36354/_0_  = _w1989_ ;
	assign \g36355/_0_  = _w2000_ ;
	assign \g36356/_0_  = _w2006_ ;
	assign \g36357/_0_  = _w2012_ ;
	assign \g36358/_0_  = _w2014_ ;
	assign \g36359/_0_  = _w2027_ ;
	assign \g36360/_0_  = _w2037_ ;
	assign \g36361/_0_  = _w2052_ ;
	assign \g36362/_0_  = _w2065_ ;
	assign \g36363/_0_  = _w2082_ ;
	assign \g36410/_0_  = _w2101_ ;
	assign \g36413/_0_  = _w2124_ ;
	assign \g36414/_0_  = _w2143_ ;
	assign \g36415/_0_  = _w2164_ ;
	assign \g36416/_0_  = _w2179_ ;
	assign \g36424/_0_  = _w2197_ ;
	assign \g36425/_0_  = _w2214_ ;
	assign \g36452/_0_  = _w2234_ ;
	assign \g36455/_0_  = _w2252_ ;
	assign \g36456/_0_  = _w2265_ ;
	assign \g36457/_0_  = _w2281_ ;
	assign \g36458/_0_  = _w2292_ ;
	assign \g36459/_0_  = _w2304_ ;
	assign \g36460/_0_  = _w2311_ ;
	assign \g36461/_0_  = _w2314_ ;
	assign \g36462/_0_  = _w2330_ ;
	assign \g36463/_0_  = _w2336_ ;
	assign \g36464/_0_  = _w2347_ ;
	assign \g36465/_0_  = _w2363_ ;
	assign \g36466/_0_  = _w2372_ ;
	assign \g36467/_0_  = _w2374_ ;
	assign \g36468/_0_  = _w2387_ ;
	assign \g36469/_0_  = _w2389_ ;
	assign \g36470/_0_  = _w2405_ ;
	assign \g36471/_0_  = _w2411_ ;
	assign \g36472/_0_  = _w2423_ ;
	assign \g36473/_0_  = _w2434_ ;
	assign \g36557/_0_  = _w2438_ ;
	assign \g36558/_0_  = _w2442_ ;
	assign \g36559/_0_  = _w2457_ ;
	assign \g36560/_0_  = _w2475_ ;
	assign \g36561/_0_  = _w2487_ ;
	assign \g36562/_0_  = _w2492_ ;
	assign \g36563/_0_  = _w2500_ ;
	assign \g36564/_0_  = _w2513_ ;
	assign \g36565/_0_  = _w2529_ ;
	assign \g36566/_0_  = _w2532_ ;
	assign \g36567/_0_  = _w2542_ ;
	assign \g36568/_0_  = _w2548_ ;
	assign \g36569/_0_  = _w2550_ ;
	assign \g36570/_0_  = _w2563_ ;
	assign \g36571/_0_  = _w2579_ ;
	assign \g36572/_0_  = _w2590_ ;
	assign \g36573/_0_  = _w2593_ ;
	assign \g36574/_0_  = _w2605_ ;
	assign \g36575/_0_  = _w2615_ ;
	assign \g36576/_0_  = _w2632_ ;
	assign \g36577/_0_  = _w2645_ ;
	assign \g36672/_0_  = _w2657_ ;
	assign \g36673/_0_  = _w2671_ ;
	assign \g36674/_0_  = _w2683_ ;
	assign \g38/_0_  = _w563_ ;
	assign \g38_dup47616/_1_  = _w352_ ;
	assign \g39789/u3_syn_4  = _w1110_ ;
	assign \g40089/_0_  = _w2743_ ;
	assign \g40090/_0_  = _w2763_ ;
	assign \g40092/_0_  = _w2793_ ;
	assign \g40093/_0_  = _w2813_ ;
	assign \g40095/_0_  = _w2822_ ;
	assign \g40096/_0_  = _w2834_ ;
	assign \g40097/_0_  = _w2842_ ;
	assign \g40098/_0_  = _w2851_ ;
	assign \g40099/_0_  = _w2865_ ;
	assign \g40100/_0_  = _w2878_ ;
	assign \g40105/_0_  = _w2886_ ;
	assign \g40106/_0_  = _w2898_ ;
	assign \g40108/_0_  = _w2921_ ;
	assign \g40109/_0_  = _w2933_ ;
	assign \g40219/_0_  = _w2944_ ;
	assign \g40220/_0_  = _w2953_ ;
	assign \g40221/_0_  = _w2962_ ;
	assign \g40222/_0_  = _w2971_ ;
	assign \g40223/_0_  = _w2983_ ;
	assign \g40228/_0_  = _w2989_ ;
	assign \g40434/_0_  = _w779_ ;
	assign \g40495/_0_  = _w2990_ ;
	assign \g40760/_0_  = _w780_ ;
	assign \g41149/u3_syn_4  = _w2991_ ;
	assign \g42397/_0_  = _w295_ ;
	assign \g42487/_0_  = _w307_ ;
	assign \g42553/_0_  = _w300_ ;
	assign \g43089/_0_  = _w430_ ;
	assign \g43163/_0_  = _w334_ ;
	assign \g43169/_0_  = _w378_ ;
	assign \g43180/_0_  = _w326_ ;
	assign \g43189_dup/_0_  = _w468_ ;
	assign \g43196/_0_  = _w498_ ;
	assign \g43217/_0_  = _w442_ ;
	assign \g43236/_0_  = _w579_ ;
	assign \g43251/_0_  = _w316_ ;
	assign \g43256/_0_  = _w481_ ;
	assign \g43272/_0_  = _w423_ ;
	assign \g43277/_0_  = _w588_ ;
	assign \g43324/_0_  = _w596_ ;
	assign \g43341/_0_  = _w460_ ;
	assign \g43350/_0_  = _w545_ ;
	assign \g43360/_0_  = _w551_ ;
	assign \g44419/_3_  = _w2994_ ;
	assign \g44452/_3_  = _w2997_ ;
	assign \g44514/_3_  = _w3001_ ;
	assign \g44515/_3_  = _w3002_ ;
	assign \g44516/_3_  = _w3005_ ;
	assign \g44583/_3_  = _w3006_ ;
	assign \g44586/_3_  = _w3009_ ;
	assign \g44587/_3_  = _w3010_ ;
	assign \g44588/_3_  = _w3011_ ;
	assign \g44589/_3_  = _w3013_ ;
	assign \g44590/_3_  = _w3016_ ;
	assign \g44591/_3_  = _w3017_ ;
	assign \g44679/_0_  = _w3018_ ;
	assign \g44680/_3_  = _w3021_ ;
	assign \g44681/_3_  = _w3022_ ;
	assign \g44682/_3_  = _w3025_ ;
	assign \g44686/_3_  = _w3026_ ;
	assign \g44687/_3_  = _w3027_ ;
	assign \g44688/_3_  = _w3028_ ;
	assign \g44689/_3_  = _w3031_ ;
	assign \g44771/_3_  = _w3032_ ;
	assign \g44785/_3_  = _w3033_ ;
	assign \g44795/_3_  = _w3034_ ;
	assign \g44796/_3_  = _w3037_ ;
	assign \g44906/_3_  = _w3038_ ;
	assign \g44968/_3_  = _w3039_ ;
	assign \g44984/_3_  = _w3040_ ;
	assign \g45042/_3_  = _w3041_ ;
	assign \g45044/_3_  = _w3044_ ;
	assign \g45115/_3_  = _w3047_ ;
	assign \g45116/_3_  = _w3048_ ;
	assign \g46478/_1_  = _w572_ ;
	assign \g46505/_0_  = _w3062_ ;
	assign \g46519/_0_  = _w342_ ;
	assign \g46696/_0_  = _w3075_ ;
	assign \g47017/_2_  = _w504_ ;
	assign \g47072_dup/_0_  = _w524_ ;
	assign \g47395/_0_  = _w387_ ;
	assign \g47397/_0_  = _w370_ ;
	assign \g47401/_0_  = _w395_ ;
	assign \g47404/_0_  = _w412_ ;
	assign \g47458/_0_  = _w3079_ ;
	assign \g47540/_0_  = _w3093_ ;
	assign \g47791/_0_  = _w517_ ;
	assign \state_reg[0]/NET0131_syn_2  = _w215_ ;
endmodule;