module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] , \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] , \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] , \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	output \sin[0]  ;
	output \sin[1]  ;
	output \sin[2]  ;
	output \sin[3]  ;
	output \sin[4]  ;
	output \sin[5]  ;
	output \sin[6]  ;
	output \sin[7]  ;
	output \sin[8]  ;
	output \sin[9]  ;
	output \sin[10]  ;
	output \sin[11]  ;
	output \sin[12]  ;
	output \sin[13]  ;
	output \sin[14]  ;
	output \sin[15]  ;
	output \sin[16]  ;
	output \sin[17]  ;
	output \sin[18]  ;
	output \sin[19]  ;
	output \sin[20]  ;
	output \sin[21]  ;
	output \sin[22]  ;
	output \sin[23]  ;
	output \sin[24]  ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\a[0] ,
		\a[1] ,
		_w26_
	);
	LUT3 #(
		.INIT('h01)
	) name1 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w27_
	);
	LUT4 #(
		.INIT('h0001)
	) name2 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[3] ,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\a[4] ,
		_w28_,
		_w29_
	);
	LUT4 #(
		.INIT('h393c)
	) name4 (
		\a[4] ,
		\a[5] ,
		\a[22] ,
		_w28_,
		_w30_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[22] ,
		_w31_
	);
	LUT2 #(
		.INIT('h9)
	) name6 (
		\a[3] ,
		_w31_,
		_w32_
	);
	LUT4 #(
		.INIT('h0fe1)
	) name7 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[22] ,
		_w33_
	);
	LUT3 #(
		.INIT('h69)
	) name8 (
		\a[3] ,
		_w31_,
		_w33_,
		_w34_
	);
	LUT3 #(
		.INIT('h56)
	) name9 (
		\a[4] ,
		\a[22] ,
		_w28_,
		_w35_
	);
	LUT4 #(
		.INIT('h6c66)
	) name10 (
		\a[4] ,
		\a[5] ,
		\a[22] ,
		_w28_,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w34_,
		_w36_,
		_w37_
	);
	LUT3 #(
		.INIT('h10)
	) name12 (
		\a[4] ,
		\a[5] ,
		_w28_,
		_w38_
	);
	LUT4 #(
		.INIT('h0100)
	) name13 (
		\a[4] ,
		\a[5] ,
		\a[6] ,
		_w28_,
		_w39_
	);
	LUT3 #(
		.INIT('h10)
	) name14 (
		\a[7] ,
		\a[8] ,
		_w39_,
		_w40_
	);
	LUT4 #(
		.INIT('h0100)
	) name15 (
		\a[7] ,
		\a[8] ,
		\a[9] ,
		_w39_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\a[10] ,
		_w41_,
		_w42_
	);
	LUT3 #(
		.INIT('h10)
	) name17 (
		\a[10] ,
		\a[11] ,
		_w41_,
		_w43_
	);
	LUT4 #(
		.INIT('h0100)
	) name18 (
		\a[10] ,
		\a[11] ,
		\a[12] ,
		_w41_,
		_w44_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name19 (
		\a[13] ,
		\a[14] ,
		\a[22] ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h6)
	) name20 (
		\a[15] ,
		_w45_,
		_w46_
	);
	LUT4 #(
		.INIT('h0100)
	) name21 (
		\a[13] ,
		\a[14] ,
		\a[15] ,
		_w44_,
		_w47_
	);
	LUT3 #(
		.INIT('h10)
	) name22 (
		\a[16] ,
		\a[17] ,
		_w47_,
		_w48_
	);
	LUT4 #(
		.INIT('h0100)
	) name23 (
		\a[16] ,
		\a[17] ,
		\a[18] ,
		_w47_,
		_w49_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name24 (
		\a[19] ,
		\a[20] ,
		\a[22] ,
		_w49_,
		_w50_
	);
	LUT4 #(
		.INIT('h393c)
	) name25 (
		\a[19] ,
		\a[20] ,
		\a[22] ,
		_w49_,
		_w51_
	);
	LUT2 #(
		.INIT('h6)
	) name26 (
		\a[21] ,
		_w50_,
		_w52_
	);
	LUT3 #(
		.INIT('h60)
	) name27 (
		\a[21] ,
		_w50_,
		_w51_,
		_w53_
	);
	LUT4 #(
		.INIT('h0060)
	) name28 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w54_
	);
	LUT4 #(
		.INIT('h2824)
	) name29 (
		\a[16] ,
		\a[17] ,
		\a[22] ,
		_w47_,
		_w55_
	);
	LUT3 #(
		.INIT('h56)
	) name30 (
		\a[18] ,
		\a[22] ,
		_w48_,
		_w56_
	);
	LUT3 #(
		.INIT('h56)
	) name31 (
		\a[19] ,
		\a[22] ,
		_w49_,
		_w57_
	);
	LUT4 #(
		.INIT('h2824)
	) name32 (
		\a[18] ,
		\a[19] ,
		\a[22] ,
		_w48_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w55_,
		_w58_,
		_w59_
	);
	LUT4 #(
		.INIT('h1118)
	) name34 (
		\a[18] ,
		\a[19] ,
		\a[22] ,
		_w48_,
		_w60_
	);
	LUT4 #(
		.INIT('h8281)
	) name35 (
		\a[16] ,
		\a[17] ,
		\a[22] ,
		_w47_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w53_,
		_w62_,
		_w63_
	);
	LUT3 #(
		.INIT('h40)
	) name38 (
		_w46_,
		_w53_,
		_w62_,
		_w64_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name39 (
		_w46_,
		_w53_,
		_w59_,
		_w62_,
		_w65_
	);
	LUT4 #(
		.INIT('h1118)
	) name40 (
		\a[16] ,
		\a[17] ,
		\a[22] ,
		_w47_,
		_w66_
	);
	LUT4 #(
		.INIT('h8281)
	) name41 (
		\a[18] ,
		\a[19] ,
		\a[22] ,
		_w48_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w54_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('h09)
	) name44 (
		\a[21] ,
		_w50_,
		_w51_,
		_w70_
	);
	LUT4 #(
		.INIT('h0900)
	) name45 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w55_,
		_w67_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT4 #(
		.INIT('h0777)
	) name48 (
		_w54_,
		_w68_,
		_w71_,
		_w72_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w65_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w60_,
		_w66_,
		_w76_
	);
	LUT4 #(
		.INIT('h0009)
	) name51 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w67_,
		_w61_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w79_,
		_w77_,
		_w80_
	);
	LUT4 #(
		.INIT('h4442)
	) name55 (
		\a[18] ,
		\a[19] ,
		\a[22] ,
		_w48_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w66_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w82_,
		_w71_,
		_w83_
	);
	LUT4 #(
		.INIT('h27ff)
	) name58 (
		_w46_,
		_w82_,
		_w79_,
		_w70_,
		_w84_
	);
	LUT4 #(
		.INIT('h6000)
	) name59 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w85_,
		_w68_,
		_w86_
	);
	LUT3 #(
		.INIT('h90)
	) name61 (
		\a[21] ,
		_w50_,
		_w51_,
		_w87_
	);
	LUT4 #(
		.INIT('h0090)
	) name62 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w88_,
		_w62_,
		_w89_
	);
	LUT4 #(
		.INIT('h135f)
	) name64 (
		_w88_,
		_w85_,
		_w62_,
		_w68_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w58_,
		_w61_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w88_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h0400)
	) name67 (
		_w78_,
		_w90_,
		_w92_,
		_w84_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w75_,
		_w93_,
		_w94_
	);
	LUT3 #(
		.INIT('h06)
	) name69 (
		\a[21] ,
		_w50_,
		_w51_,
		_w95_
	);
	LUT4 #(
		.INIT('h0600)
	) name70 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w96_
	);
	LUT4 #(
		.INIT('h4442)
	) name71 (
		\a[16] ,
		\a[17] ,
		\a[22] ,
		_w47_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w97_,
		_w58_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w96_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w66_,
		_w58_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w85_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w81_,
		_w61_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w85_,
		_w102_,
		_w103_
	);
	LUT3 #(
		.INIT('h57)
	) name78 (
		_w85_,
		_w102_,
		_w100_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w99_,
		_w104_,
		_w105_
	);
	LUT4 #(
		.INIT('h0006)
	) name80 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w82_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w79_,
		_w71_,
		_w108_
	);
	LUT4 #(
		.INIT('h0777)
	) name83 (
		_w82_,
		_w106_,
		_w79_,
		_w71_,
		_w109_
	);
	LUT3 #(
		.INIT('h80)
	) name84 (
		_w46_,
		_w53_,
		_w62_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w88_,
		_w68_,
		_w111_
	);
	LUT3 #(
		.INIT('h10)
	) name86 (
		_w110_,
		_w111_,
		_w109_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w81_,
		_w97_,
		_w113_
	);
	LUT4 #(
		.INIT('h153f)
	) name88 (
		_w113_,
		_w59_,
		_w85_,
		_w77_,
		_w114_
	);
	LUT3 #(
		.INIT('h80)
	) name89 (
		_w46_,
		_w53_,
		_w113_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w97_,
		_w67_,
		_w116_
	);
	LUT3 #(
		.INIT('h40)
	) name91 (
		_w46_,
		_w53_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w88_,
		_w82_,
		_w118_
	);
	LUT3 #(
		.INIT('h01)
	) name93 (
		_w117_,
		_w118_,
		_w115_,
		_w119_
	);
	LUT4 #(
		.INIT('h0002)
	) name94 (
		_w114_,
		_w117_,
		_w118_,
		_w115_,
		_w120_
	);
	LUT4 #(
		.INIT('h9000)
	) name95 (
		\a[21] ,
		_w50_,
		_w51_,
		_w46_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w121_,
		_w113_,
		_w122_
	);
	LUT4 #(
		.INIT('h0777)
	) name97 (
		_w121_,
		_w113_,
		_w106_,
		_w79_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w82_,
		_w77_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w55_,
		_w81_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w77_,
		_w125_,
		_w126_
	);
	LUT3 #(
		.INIT('h37)
	) name101 (
		_w82_,
		_w77_,
		_w125_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w71_,
		_w100_,
		_w128_
	);
	LUT3 #(
		.INIT('h20)
	) name103 (
		_w127_,
		_w128_,
		_w123_,
		_w129_
	);
	LUT4 #(
		.INIT('h8000)
	) name104 (
		_w120_,
		_w129_,
		_w105_,
		_w112_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w94_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h80)
	) name106 (
		_w87_,
		_w46_,
		_w102_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w53_,
		_w72_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w60_,
		_w97_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w88_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w54_,
		_w98_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w106_,
		_w116_,
		_w137_
	);
	LUT4 #(
		.INIT('h153f)
	) name112 (
		_w106_,
		_w54_,
		_w98_,
		_w116_,
		_w138_
	);
	LUT4 #(
		.INIT('h0100)
	) name113 (
		_w132_,
		_w133_,
		_w135_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w62_,
		_w71_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w121_,
		_w79_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w121_,
		_w62_,
		_w142_
	);
	LUT4 #(
		.INIT('h0757)
	) name117 (
		_w121_,
		_w79_,
		_w62_,
		_w71_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w79_,
		_w96_,
		_w144_
	);
	LUT3 #(
		.INIT('h80)
	) name119 (
		_w46_,
		_w95_,
		_w113_,
		_w145_
	);
	LUT3 #(
		.INIT('h80)
	) name120 (
		_w46_,
		_w95_,
		_w102_,
		_w146_
	);
	LUT4 #(
		.INIT('h777f)
	) name121 (
		_w46_,
		_w95_,
		_w113_,
		_w102_,
		_w147_
	);
	LUT3 #(
		.INIT('h20)
	) name122 (
		_w143_,
		_w144_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w139_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w106_,
		_w68_,
		_w150_
	);
	LUT4 #(
		.INIT('h135f)
	) name125 (
		_w106_,
		_w54_,
		_w68_,
		_w100_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w96_,
		_w68_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w54_,
		_w102_,
		_w153_
	);
	LUT4 #(
		.INIT('h0777)
	) name128 (
		_w54_,
		_w102_,
		_w96_,
		_w68_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		_w151_,
		_w154_,
		_w155_
	);
	LUT3 #(
		.INIT('h20)
	) name130 (
		_w87_,
		_w46_,
		_w102_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w125_,
		_w71_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w76_,
		_w71_,
		_w158_
	);
	LUT4 #(
		.INIT('h135f)
	) name133 (
		_w76_,
		_w96_,
		_w71_,
		_w72_,
		_w159_
	);
	LUT3 #(
		.INIT('h10)
	) name134 (
		_w156_,
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w95_,
		_w59_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w88_,
		_w79_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w121_,
		_w134_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w88_,
		_w98_,
		_w164_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name139 (
		_w87_,
		_w46_,
		_w134_,
		_w98_,
		_w165_
	);
	LUT3 #(
		.INIT('h10)
	) name140 (
		_w161_,
		_w162_,
		_w165_,
		_w166_
	);
	LUT3 #(
		.INIT('h80)
	) name141 (
		_w155_,
		_w160_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('h40)
	) name142 (
		_w46_,
		_w95_,
		_w113_,
		_w168_
	);
	LUT3 #(
		.INIT('h40)
	) name143 (
		_w46_,
		_w95_,
		_w102_,
		_w169_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name144 (
		_w46_,
		_w95_,
		_w113_,
		_w102_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w121_,
		_w91_,
		_w171_
	);
	LUT4 #(
		.INIT('h0777)
	) name146 (
		_w121_,
		_w91_,
		_w96_,
		_w116_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w59_,
		_w77_,
		_w173_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name148 (
		_w46_,
		_w59_,
		_w70_,
		_w116_,
		_w174_
	);
	LUT3 #(
		.INIT('h80)
	) name149 (
		_w172_,
		_w174_,
		_w170_,
		_w175_
	);
	LUT3 #(
		.INIT('h80)
	) name150 (
		_w46_,
		_w95_,
		_w125_,
		_w176_
	);
	LUT4 #(
		.INIT('h373f)
	) name151 (
		_w46_,
		_w95_,
		_w91_,
		_w125_,
		_w177_
	);
	LUT3 #(
		.INIT('h80)
	) name152 (
		_w46_,
		_w53_,
		_w116_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w121_,
		_w98_,
		_w179_
	);
	LUT3 #(
		.INIT('h10)
	) name154 (
		_w178_,
		_w179_,
		_w177_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w106_,
		_w72_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w77_,
		_w116_,
		_w182_
	);
	LUT4 #(
		.INIT('h153f)
	) name157 (
		_w106_,
		_w77_,
		_w116_,
		_w72_,
		_w183_
	);
	LUT3 #(
		.INIT('h40)
	) name158 (
		_w46_,
		_w95_,
		_w125_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w106_,
		_w98_,
		_w185_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name160 (
		_w46_,
		_w95_,
		_w125_,
		_w98_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w183_,
		_w186_,
		_w187_
	);
	LUT3 #(
		.INIT('h80)
	) name162 (
		_w175_,
		_w180_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w82_,
		_w96_,
		_w189_
	);
	LUT4 #(
		.INIT('h135f)
	) name164 (
		_w82_,
		_w77_,
		_w96_,
		_w100_,
		_w190_
	);
	LUT4 #(
		.INIT('h8000)
	) name165 (
		_w175_,
		_w180_,
		_w187_,
		_w190_,
		_w191_
	);
	LUT3 #(
		.INIT('h80)
	) name166 (
		_w149_,
		_w167_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w131_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w121_,
		_w116_,
		_w194_
	);
	LUT4 #(
		.INIT('h153f)
	) name169 (
		_w121_,
		_w76_,
		_w77_,
		_w116_,
		_w195_
	);
	LUT3 #(
		.INIT('h10)
	) name170 (
		_w171_,
		_w146_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w134_,
		_w96_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w96_,
		_w100_,
		_w198_
	);
	LUT3 #(
		.INIT('h37)
	) name173 (
		_w134_,
		_w96_,
		_w100_,
		_w199_
	);
	LUT3 #(
		.INIT('h57)
	) name174 (
		_w54_,
		_w59_,
		_w98_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w199_,
		_w200_,
		_w201_
	);
	LUT3 #(
		.INIT('h37)
	) name176 (
		_w88_,
		_w59_,
		_w85_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w106_,
		_w100_,
		_w203_
	);
	LUT4 #(
		.INIT('h153f)
	) name178 (
		_w106_,
		_w91_,
		_w77_,
		_w100_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w202_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w60_,
		_w55_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w206_,
		_w96_,
		_w207_
	);
	LUT3 #(
		.INIT('h37)
	) name182 (
		_w206_,
		_w96_,
		_w116_,
		_w208_
	);
	LUT3 #(
		.INIT('h40)
	) name183 (
		_w46_,
		_w95_,
		_w62_,
		_w209_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name184 (
		_w46_,
		_w95_,
		_w62_,
		_w116_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w91_,
		_w71_,
		_w211_
	);
	LUT4 #(
		.INIT('h1bff)
	) name186 (
		_w46_,
		_w113_,
		_w91_,
		_w70_,
		_w212_
	);
	LUT4 #(
		.INIT('h8000)
	) name187 (
		_w208_,
		_w170_,
		_w210_,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('h8000)
	) name188 (
		_w196_,
		_w201_,
		_w205_,
		_w213_,
		_w214_
	);
	LUT4 #(
		.INIT('h0777)
	) name189 (
		_w88_,
		_w82_,
		_w79_,
		_w96_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT4 #(
		.INIT('h1dff)
	) name191 (
		_w87_,
		_w46_,
		_w53_,
		_w116_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w77_,
		_w62_,
		_w218_
	);
	LUT3 #(
		.INIT('h40)
	) name193 (
		_w46_,
		_w53_,
		_w113_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w54_,
		_w72_,
		_w220_
	);
	LUT3 #(
		.INIT('h80)
	) name195 (
		_w46_,
		_w95_,
		_w62_,
		_w221_
	);
	LUT4 #(
		.INIT('h0001)
	) name196 (
		_w218_,
		_w219_,
		_w220_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w217_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w134_,
		_w106_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w134_,
		_w54_,
		_w225_
	);
	LUT3 #(
		.INIT('h01)
	) name200 (
		_w224_,
		_w225_,
		_w145_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w121_,
		_w125_,
		_w227_
	);
	LUT4 #(
		.INIT('h153f)
	) name202 (
		_w121_,
		_w79_,
		_w77_,
		_w125_,
		_w228_
	);
	LUT4 #(
		.INIT('h0777)
	) name203 (
		_w85_,
		_w68_,
		_w125_,
		_w71_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT3 #(
		.INIT('h01)
	) name205 (
		_w176_,
		_w108_,
		_w150_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w77_,
		_w68_,
		_w232_
	);
	LUT4 #(
		.INIT('h135f)
	) name207 (
		_w77_,
		_w96_,
		_w68_,
		_w72_,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w111_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('h8000)
	) name209 (
		_w226_,
		_w230_,
		_w231_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w134_,
		_w71_,
		_w236_
	);
	LUT3 #(
		.INIT('h1f)
	) name211 (
		_w134_,
		_w68_,
		_w71_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w206_,
		_w88_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w206_,
		_w85_,
		_w239_
	);
	LUT4 #(
		.INIT('h135f)
	) name214 (
		_w206_,
		_w88_,
		_w85_,
		_w62_,
		_w240_
	);
	LUT4 #(
		.INIT('h1357)
	) name215 (
		_w206_,
		_w88_,
		_w85_,
		_w62_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w134_,
		_w85_,
		_w242_
	);
	LUT4 #(
		.INIT('h135f)
	) name217 (
		_w121_,
		_w134_,
		_w59_,
		_w85_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w88_,
		_w113_,
		_w244_
	);
	LUT4 #(
		.INIT('h4000)
	) name219 (
		_w244_,
		_w174_,
		_w241_,
		_w243_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w237_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w134_,
		_w77_,
		_w247_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name222 (
		_w46_,
		_w134_,
		_w70_,
		_w100_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w85_,
		_w125_,
		_w249_
	);
	LUT4 #(
		.INIT('h153f)
	) name224 (
		_w85_,
		_w96_,
		_w68_,
		_w125_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w248_,
		_w250_,
		_w251_
	);
	LUT3 #(
		.INIT('h80)
	) name226 (
		_w46_,
		_w53_,
		_w82_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w85_,
		_w72_,
		_w253_
	);
	LUT4 #(
		.INIT('h37bf)
	) name228 (
		_w46_,
		_w53_,
		_w125_,
		_w72_,
		_w254_
	);
	LUT3 #(
		.INIT('h10)
	) name229 (
		_w252_,
		_w181_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w77_,
		_w72_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w121_,
		_w72_,
		_w257_
	);
	LUT3 #(
		.INIT('h57)
	) name232 (
		_w121_,
		_w62_,
		_w72_,
		_w258_
	);
	LUT3 #(
		.INIT('h10)
	) name233 (
		_w117_,
		_w256_,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('h0777)
	) name234 (
		_w206_,
		_w121_,
		_w106_,
		_w79_,
		_w260_
	);
	LUT3 #(
		.INIT('h10)
	) name235 (
		_w132_,
		_w158_,
		_w260_,
		_w261_
	);
	LUT4 #(
		.INIT('h8000)
	) name236 (
		_w259_,
		_w261_,
		_w251_,
		_w255_,
		_w262_
	);
	LUT4 #(
		.INIT('h8000)
	) name237 (
		_w246_,
		_w223_,
		_w235_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w216_,
		_w263_,
		_w264_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name239 (
		_w46_,
		_w53_,
		_w113_,
		_w68_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w106_,
		_w91_,
		_w266_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name241 (
		_w46_,
		_w82_,
		_w95_,
		_w91_,
		_w267_
	);
	LUT4 #(
		.INIT('h153f)
	) name242 (
		_w54_,
		_w59_,
		_w77_,
		_w98_,
		_w268_
	);
	LUT3 #(
		.INIT('h80)
	) name243 (
		_w267_,
		_w268_,
		_w265_,
		_w269_
	);
	LUT4 #(
		.INIT('h0777)
	) name244 (
		_w88_,
		_w91_,
		_w77_,
		_w116_,
		_w270_
	);
	LUT3 #(
		.INIT('h40)
	) name245 (
		_w46_,
		_w53_,
		_w82_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w88_,
		_w125_,
		_w272_
	);
	LUT4 #(
		.INIT('h135f)
	) name247 (
		_w88_,
		_w79_,
		_w125_,
		_w71_,
		_w273_
	);
	LUT4 #(
		.INIT('h1000)
	) name248 (
		_w271_,
		_w209_,
		_w270_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w88_,
		_w72_,
		_w275_
	);
	LUT4 #(
		.INIT('h153f)
	) name250 (
		_w82_,
		_w121_,
		_w98_,
		_w71_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w121_,
		_w100_,
		_w278_
	);
	LUT3 #(
		.INIT('h1f)
	) name253 (
		_w121_,
		_w54_,
		_w100_,
		_w279_
	);
	LUT4 #(
		.INIT('h115f)
	) name254 (
		_w121_,
		_w54_,
		_w59_,
		_w100_,
		_w280_
	);
	LUT3 #(
		.INIT('h40)
	) name255 (
		_w275_,
		_w276_,
		_w280_,
		_w281_
	);
	LUT3 #(
		.INIT('h80)
	) name256 (
		_w269_,
		_w274_,
		_w281_,
		_w282_
	);
	LUT3 #(
		.INIT('h37)
	) name257 (
		_w88_,
		_w82_,
		_w106_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w77_,
		_w98_,
		_w284_
	);
	LUT3 #(
		.INIT('h57)
	) name259 (
		_w77_,
		_w125_,
		_w98_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w206_,
		_w71_,
		_w286_
	);
	LUT4 #(
		.INIT('h153f)
	) name261 (
		_w206_,
		_w121_,
		_w116_,
		_w71_,
		_w287_
	);
	LUT3 #(
		.INIT('h80)
	) name262 (
		_w283_,
		_w285_,
		_w287_,
		_w288_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name263 (
		_w87_,
		_w46_,
		_w134_,
		_w116_,
		_w289_
	);
	LUT4 #(
		.INIT('h1000)
	) name264 (
		_w184_,
		_w211_,
		_w237_,
		_w289_,
		_w290_
	);
	LUT3 #(
		.INIT('h37)
	) name265 (
		_w59_,
		_w85_,
		_w100_,
		_w291_
	);
	LUT4 #(
		.INIT('h0777)
	) name266 (
		_w206_,
		_w121_,
		_w85_,
		_w102_,
		_w292_
	);
	LUT4 #(
		.INIT('h135f)
	) name267 (
		_w113_,
		_w85_,
		_w77_,
		_w125_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT4 #(
		.INIT('h4000)
	) name269 (
		_w158_,
		_w291_,
		_w292_,
		_w293_,
		_w295_
	);
	LUT3 #(
		.INIT('h80)
	) name270 (
		_w288_,
		_w290_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w206_,
		_w54_,
		_w297_
	);
	LUT3 #(
		.INIT('h37)
	) name272 (
		_w134_,
		_w85_,
		_w72_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w76_,
		_w96_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w98_,
		_w71_,
		_w301_
	);
	LUT4 #(
		.INIT('h153f)
	) name276 (
		_w96_,
		_w98_,
		_w71_,
		_w100_,
		_w302_
	);
	LUT4 #(
		.INIT('h135f)
	) name277 (
		_w53_,
		_w106_,
		_w116_,
		_w100_,
		_w303_
	);
	LUT4 #(
		.INIT('h1000)
	) name278 (
		_w300_,
		_w142_,
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w299_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w91_,
		_w96_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w156_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w85_,
		_w91_,
		_w308_
	);
	LUT4 #(
		.INIT('h0777)
	) name283 (
		_w85_,
		_w91_,
		_w77_,
		_w62_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w102_,
		_w70_,
		_w310_
	);
	LUT3 #(
		.INIT('h80)
	) name285 (
		_w46_,
		_w102_,
		_w70_,
		_w311_
	);
	LUT3 #(
		.INIT('h10)
	) name286 (
		_w141_,
		_w311_,
		_w309_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w307_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h0777)
	) name288 (
		_w88_,
		_w113_,
		_w77_,
		_w100_,
		_w314_
	);
	LUT4 #(
		.INIT('h135f)
	) name289 (
		_w88_,
		_w77_,
		_w68_,
		_w72_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w121_,
		_w76_,
		_w316_
	);
	LUT4 #(
		.INIT('h153f)
	) name291 (
		_w206_,
		_w121_,
		_w76_,
		_w106_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w76_,
		_w106_,
		_w318_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name293 (
		_w46_,
		_w76_,
		_w95_,
		_w62_,
		_w319_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		_w317_,
		_w319_,
		_w314_,
		_w315_,
		_w320_
	);
	LUT3 #(
		.INIT('h80)
	) name295 (
		_w307_,
		_w312_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		_w296_,
		_w282_,
		_w305_,
		_w321_,
		_w322_
	);
	LUT3 #(
		.INIT('h07)
	) name297 (
		_w216_,
		_w263_,
		_w322_,
		_w323_
	);
	LUT4 #(
		.INIT('h37bf)
	) name298 (
		_w46_,
		_w95_,
		_w102_,
		_w62_,
		_w324_
	);
	LUT4 #(
		.INIT('h0777)
	) name299 (
		_w95_,
		_w113_,
		_w85_,
		_w72_,
		_w325_
	);
	LUT4 #(
		.INIT('h1000)
	) name300 (
		_w209_,
		_w86_,
		_w324_,
		_w325_,
		_w326_
	);
	LUT3 #(
		.INIT('h57)
	) name301 (
		_w54_,
		_w68_,
		_w72_,
		_w327_
	);
	LUT4 #(
		.INIT('h135f)
	) name302 (
		_w106_,
		_w54_,
		_w91_,
		_w125_,
		_w328_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name303 (
		_w46_,
		_w95_,
		_w98_,
		_w100_,
		_w329_
	);
	LUT4 #(
		.INIT('h0777)
	) name304 (
		_w53_,
		_w82_,
		_w91_,
		_w96_,
		_w330_
	);
	LUT4 #(
		.INIT('h135f)
	) name305 (
		_w85_,
		_w96_,
		_w125_,
		_w100_,
		_w331_
	);
	LUT4 #(
		.INIT('h8000)
	) name306 (
		_w330_,
		_w328_,
		_w329_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name307 (
		_w46_,
		_w95_,
		_w125_,
		_w116_,
		_w333_
	);
	LUT3 #(
		.INIT('h37)
	) name308 (
		_w206_,
		_w106_,
		_w72_,
		_w334_
	);
	LUT4 #(
		.INIT('h0777)
	) name309 (
		_w76_,
		_w106_,
		_w85_,
		_w79_,
		_w335_
	);
	LUT3 #(
		.INIT('h37)
	) name310 (
		_w76_,
		_w96_,
		_w72_,
		_w336_
	);
	LUT4 #(
		.INIT('h8000)
	) name311 (
		_w335_,
		_w336_,
		_w333_,
		_w334_,
		_w337_
	);
	LUT4 #(
		.INIT('h8000)
	) name312 (
		_w332_,
		_w326_,
		_w327_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w54_,
		_w91_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w85_,
		_w98_,
		_w340_
	);
	LUT4 #(
		.INIT('h37bf)
	) name315 (
		_w46_,
		_w53_,
		_w91_,
		_w98_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w189_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('h373f)
	) name317 (
		_w46_,
		_w53_,
		_w113_,
		_w102_,
		_w343_
	);
	LUT3 #(
		.INIT('h40)
	) name318 (
		_w189_,
		_w341_,
		_w343_,
		_w344_
	);
	LUT4 #(
		.INIT('h0777)
	) name319 (
		_w82_,
		_w106_,
		_w54_,
		_w102_,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w184_,
		_w345_,
		_w346_
	);
	LUT3 #(
		.INIT('h80)
	) name321 (
		_w46_,
		_w95_,
		_w59_,
		_w347_
	);
	LUT3 #(
		.INIT('h40)
	) name322 (
		_w46_,
		_w95_,
		_w59_,
		_w348_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name323 (
		_w46_,
		_w95_,
		_w59_,
		_w98_,
		_w349_
	);
	LUT3 #(
		.INIT('h10)
	) name324 (
		_w308_,
		_w347_,
		_w349_,
		_w350_
	);
	LUT3 #(
		.INIT('h80)
	) name325 (
		_w346_,
		_w350_,
		_w344_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w54_,
		_w79_,
		_w352_
	);
	LUT4 #(
		.INIT('h153f)
	) name327 (
		_w53_,
		_w96_,
		_w68_,
		_w116_,
		_w353_
	);
	LUT4 #(
		.INIT('h0100)
	) name328 (
		_w352_,
		_w150_,
		_w146_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name329 (
		_w56_,
		_w57_,
		_w97_,
		_w61_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		_w95_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		_w208_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w354_,
		_w357_,
		_w358_
	);
	LUT3 #(
		.INIT('h80)
	) name333 (
		_w351_,
		_w338_,
		_w358_,
		_w359_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name334 (
		\a[7] ,
		\a[8] ,
		\a[22] ,
		_w39_,
		_w360_
	);
	LUT2 #(
		.INIT('h9)
	) name335 (
		\a[9] ,
		_w360_,
		_w361_
	);
	LUT4 #(
		.INIT('h007f)
	) name336 (
		_w351_,
		_w338_,
		_w358_,
		_w361_,
		_w362_
	);
	LUT3 #(
		.INIT('h56)
	) name337 (
		\a[10] ,
		\a[22] ,
		_w41_,
		_w363_
	);
	LUT4 #(
		.INIT('h007f)
	) name338 (
		_w351_,
		_w338_,
		_w358_,
		_w363_,
		_w364_
	);
	LUT4 #(
		.INIT('h011f)
	) name339 (
		_w193_,
		_w323_,
		_w362_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('h393c)
	) name340 (
		\a[10] ,
		\a[11] ,
		\a[22] ,
		_w41_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w76_,
		_w54_,
		_w367_
	);
	LUT3 #(
		.INIT('h1f)
	) name342 (
		_w206_,
		_w134_,
		_w85_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT4 #(
		.INIT('h37bf)
	) name344 (
		_w46_,
		_w53_,
		_w134_,
		_w62_,
		_w370_
	);
	LUT4 #(
		.INIT('h153f)
	) name345 (
		_w54_,
		_w79_,
		_w77_,
		_w98_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w76_,
		_w85_,
		_w372_
	);
	LUT4 #(
		.INIT('h0777)
	) name347 (
		_w76_,
		_w85_,
		_w77_,
		_w68_,
		_w373_
	);
	LUT3 #(
		.INIT('h80)
	) name348 (
		_w371_,
		_w373_,
		_w370_,
		_w374_
	);
	LUT3 #(
		.INIT('h37)
	) name349 (
		_w68_,
		_w71_,
		_w72_,
		_w375_
	);
	LUT4 #(
		.INIT('h337f)
	) name350 (
		_w46_,
		_w70_,
		_w68_,
		_w72_,
		_w376_
	);
	LUT4 #(
		.INIT('h1f3f)
	) name351 (
		_w46_,
		_w102_,
		_w70_,
		_w116_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w376_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w113_,
		_w71_,
		_w379_
	);
	LUT4 #(
		.INIT('h0777)
	) name354 (
		_w206_,
		_w54_,
		_w79_,
		_w71_,
		_w380_
	);
	LUT4 #(
		.INIT('h0100)
	) name355 (
		_w64_,
		_w182_,
		_w379_,
		_w380_,
		_w381_
	);
	LUT4 #(
		.INIT('h8000)
	) name356 (
		_w369_,
		_w378_,
		_w381_,
		_w374_,
		_w382_
	);
	LUT3 #(
		.INIT('h57)
	) name357 (
		_w54_,
		_w59_,
		_w100_,
		_w383_
	);
	LUT4 #(
		.INIT('h5d5f)
	) name358 (
		_w87_,
		_w46_,
		_w79_,
		_w116_,
		_w384_
	);
	LUT3 #(
		.INIT('h80)
	) name359 (
		_w195_,
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		_w121_,
		_w68_,
		_w386_
	);
	LUT3 #(
		.INIT('h57)
	) name361 (
		_w121_,
		_w68_,
		_w72_,
		_w387_
	);
	LUT4 #(
		.INIT('h557f)
	) name362 (
		_w87_,
		_w46_,
		_w68_,
		_w72_,
		_w388_
	);
	LUT3 #(
		.INIT('h40)
	) name363 (
		_w158_,
		_w291_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w385_,
		_w389_,
		_w390_
	);
	LUT4 #(
		.INIT('h557f)
	) name365 (
		_w87_,
		_w46_,
		_w113_,
		_w102_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w111_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		_w82_,
		_w121_,
		_w393_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name368 (
		_w87_,
		_w46_,
		_w82_,
		_w125_,
		_w394_
	);
	LUT4 #(
		.INIT('h57df)
	) name369 (
		_w87_,
		_w46_,
		_w113_,
		_w125_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT4 #(
		.INIT('h8000)
	) name371 (
		_w385_,
		_w389_,
		_w392_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w382_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w59_,
		_w71_,
		_w399_
	);
	LUT4 #(
		.INIT('h27ff)
	) name374 (
		_w46_,
		_w59_,
		_w91_,
		_w70_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w284_,
		_w400_,
		_w401_
	);
	LUT4 #(
		.INIT('h01ff)
	) name376 (
		_w82_,
		_w125_,
		_w98_,
		_w71_,
		_w402_
	);
	LUT3 #(
		.INIT('h80)
	) name377 (
		_w127_,
		_w212_,
		_w402_,
		_w403_
	);
	LUT4 #(
		.INIT('h333f)
	) name378 (
		_w46_,
		_w53_,
		_w59_,
		_w100_,
		_w404_
	);
	LUT3 #(
		.INIT('h80)
	) name379 (
		_w401_,
		_w403_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w382_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		_w206_,
		_w77_,
		_w407_
	);
	LUT4 #(
		.INIT('h4f5f)
	) name382 (
		_w206_,
		_w46_,
		_w70_,
		_w62_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w248_,
		_w408_,
		_w409_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name384 (
		_w46_,
		_w70_,
		_w62_,
		_w100_,
		_w410_
	);
	LUT4 #(
		.INIT('h0800)
	) name385 (
		_w248_,
		_w408_,
		_w236_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w173_,
		_w411_,
		_w412_
	);
	LUT3 #(
		.INIT('h80)
	) name387 (
		_w382_,
		_w405_,
		_w412_,
		_w413_
	);
	LUT4 #(
		.INIT('h5777)
	) name388 (
		_w382_,
		_w397_,
		_w405_,
		_w412_,
		_w414_
	);
	LUT4 #(
		.INIT('h8000)
	) name389 (
		_w382_,
		_w397_,
		_w405_,
		_w412_,
		_w415_
	);
	LUT4 #(
		.INIT('h2888)
	) name390 (
		_w382_,
		_w397_,
		_w405_,
		_w412_,
		_w416_
	);
	LUT4 #(
		.INIT('h5001)
	) name391 (
		_w366_,
		_w359_,
		_w398_,
		_w413_,
		_w417_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name392 (
		_w366_,
		_w359_,
		_w414_,
		_w415_,
		_w418_
	);
	LUT3 #(
		.INIT('h56)
	) name393 (
		\a[12] ,
		\a[22] ,
		_w43_,
		_w419_
	);
	LUT4 #(
		.INIT('h007f)
	) name394 (
		_w351_,
		_w338_,
		_w358_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('h7f80)
	) name395 (
		_w351_,
		_w338_,
		_w358_,
		_w419_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w416_,
		_w421_,
		_w422_
	);
	LUT3 #(
		.INIT('h01)
	) name397 (
		_w418_,
		_w417_,
		_w422_,
		_w423_
	);
	LUT4 #(
		.INIT('h393c)
	) name398 (
		\a[13] ,
		\a[14] ,
		\a[22] ,
		_w44_,
		_w424_
	);
	LUT4 #(
		.INIT('h777f)
	) name399 (
		_w46_,
		_w95_,
		_w125_,
		_w98_,
		_w425_
	);
	LUT4 #(
		.INIT('h135f)
	) name400 (
		_w88_,
		_w76_,
		_w98_,
		_w71_,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name402 (
		_w46_,
		_w82_,
		_w70_,
		_w98_,
		_w428_
	);
	LUT4 #(
		.INIT('h57df)
	) name403 (
		_w87_,
		_w46_,
		_w116_,
		_w100_,
		_w429_
	);
	LUT3 #(
		.INIT('h80)
	) name404 (
		_w429_,
		_w186_,
		_w428_,
		_w430_
	);
	LUT4 #(
		.INIT('h0777)
	) name405 (
		_w121_,
		_w59_,
		_w85_,
		_w100_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w88_,
		_w100_,
		_w432_
	);
	LUT4 #(
		.INIT('h153f)
	) name407 (
		_w88_,
		_w76_,
		_w85_,
		_w100_,
		_w433_
	);
	LUT4 #(
		.INIT('h1000)
	) name408 (
		_w386_,
		_w64_,
		_w431_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('h131f)
	) name409 (
		_w206_,
		_w82_,
		_w106_,
		_w77_,
		_w435_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name410 (
		_w46_,
		_w76_,
		_w95_,
		_w59_,
		_w436_
	);
	LUT4 #(
		.INIT('h0777)
	) name411 (
		_w91_,
		_w96_,
		_w125_,
		_w71_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT3 #(
		.INIT('h80)
	) name413 (
		_w435_,
		_w436_,
		_w437_,
		_w439_
	);
	LUT4 #(
		.INIT('h8000)
	) name414 (
		_w427_,
		_w430_,
		_w434_,
		_w439_,
		_w440_
	);
	LUT3 #(
		.INIT('h80)
	) name415 (
		_w214_,
		_w215_,
		_w440_,
		_w441_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name416 (
		_w206_,
		_w46_,
		_w53_,
		_w79_,
		_w442_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name417 (
		_w46_,
		_w95_,
		_w59_,
		_w72_,
		_w443_
	);
	LUT3 #(
		.INIT('h57)
	) name418 (
		_w121_,
		_w79_,
		_w98_,
		_w444_
	);
	LUT3 #(
		.INIT('h80)
	) name419 (
		_w442_,
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w221_,
		_w239_,
		_w446_
	);
	LUT3 #(
		.INIT('h80)
	) name421 (
		_w226_,
		_w445_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('h0777)
	) name422 (
		_w54_,
		_w79_,
		_w96_,
		_w68_,
		_w448_
	);
	LUT4 #(
		.INIT('h135f)
	) name423 (
		_w134_,
		_w106_,
		_w85_,
		_w79_,
		_w449_
	);
	LUT4 #(
		.INIT('h0777)
	) name424 (
		_w76_,
		_w106_,
		_w98_,
		_w71_,
		_w450_
	);
	LUT4 #(
		.INIT('h135f)
	) name425 (
		_w77_,
		_w96_,
		_w125_,
		_w72_,
		_w451_
	);
	LUT4 #(
		.INIT('h8000)
	) name426 (
		_w450_,
		_w451_,
		_w448_,
		_w449_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w257_,
		_w267_,
		_w453_
	);
	LUT3 #(
		.INIT('h57)
	) name428 (
		_w88_,
		_w79_,
		_w91_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w151_,
		_w454_,
		_w455_
	);
	LUT4 #(
		.INIT('h153f)
	) name430 (
		_w88_,
		_w76_,
		_w54_,
		_w72_,
		_w456_
	);
	LUT3 #(
		.INIT('h10)
	) name431 (
		_w399_,
		_w110_,
		_w456_,
		_w457_
	);
	LUT4 #(
		.INIT('h8000)
	) name432 (
		_w452_,
		_w453_,
		_w455_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w447_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w441_,
		_w459_,
		_w460_
	);
	LUT4 #(
		.INIT('h0777)
	) name435 (
		_w131_,
		_w192_,
		_w441_,
		_w459_,
		_w461_
	);
	LUT4 #(
		.INIT('h7888)
	) name436 (
		_w131_,
		_w192_,
		_w441_,
		_w459_,
		_w462_
	);
	LUT3 #(
		.INIT('h7b)
	) name437 (
		_w398_,
		_w462_,
		_w424_,
		_w463_
	);
	LUT3 #(
		.INIT('h56)
	) name438 (
		\a[13] ,
		\a[22] ,
		_w44_,
		_w464_
	);
	LUT4 #(
		.INIT('h6e76)
	) name439 (
		_w193_,
		_w460_,
		_w398_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w463_,
		_w465_,
		_w466_
	);
	LUT3 #(
		.INIT('h80)
	) name441 (
		_w423_,
		_w463_,
		_w465_,
		_w467_
	);
	LUT3 #(
		.INIT('h78)
	) name442 (
		_w216_,
		_w263_,
		_w322_,
		_w468_
	);
	LUT4 #(
		.INIT('h4552)
	) name443 (
		_w193_,
		_w424_,
		_w264_,
		_w322_,
		_w469_
	);
	LUT3 #(
		.INIT('h7b)
	) name444 (
		_w398_,
		_w462_,
		_w464_,
		_w470_
	);
	LUT4 #(
		.INIT('h6e76)
	) name445 (
		_w193_,
		_w460_,
		_w398_,
		_w419_,
		_w471_
	);
	LUT4 #(
		.INIT('h2bbb)
	) name446 (
		_w362_,
		_w469_,
		_w470_,
		_w471_,
		_w472_
	);
	LUT3 #(
		.INIT('h15)
	) name447 (
		_w423_,
		_w463_,
		_w465_,
		_w473_
	);
	LUT3 #(
		.INIT('h6a)
	) name448 (
		_w423_,
		_w463_,
		_w465_,
		_w474_
	);
	LUT3 #(
		.INIT('h54)
	) name449 (
		_w467_,
		_w472_,
		_w473_,
		_w475_
	);
	LUT4 #(
		.INIT('h4054)
	) name450 (
		_w365_,
		_w423_,
		_w466_,
		_w472_,
		_w476_
	);
	LUT4 #(
		.INIT('h1555)
	) name451 (
		_w366_,
		_w351_,
		_w338_,
		_w358_,
		_w477_
	);
	LUT4 #(
		.INIT('h0e16)
	) name452 (
		_w193_,
		_w460_,
		_w398_,
		_w424_,
		_w478_
	);
	LUT4 #(
		.INIT('h00c1)
	) name453 (
		_w359_,
		_w398_,
		_w413_,
		_w419_,
		_w479_
	);
	LUT4 #(
		.INIT('hec00)
	) name454 (
		_w359_,
		_w414_,
		_w415_,
		_w419_,
		_w480_
	);
	LUT4 #(
		.INIT('h007f)
	) name455 (
		_w351_,
		_w338_,
		_w358_,
		_w464_,
		_w481_
	);
	LUT4 #(
		.INIT('h7f80)
	) name456 (
		_w351_,
		_w338_,
		_w358_,
		_w464_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		_w416_,
		_w482_,
		_w483_
	);
	LUT3 #(
		.INIT('h01)
	) name458 (
		_w480_,
		_w479_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h69)
	) name459 (
		_w477_,
		_w478_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h2a02)
	) name460 (
		_w365_,
		_w423_,
		_w466_,
		_w472_,
		_w486_
	);
	LUT4 #(
		.INIT('h999a)
	) name461 (
		_w365_,
		_w467_,
		_w472_,
		_w473_,
		_w487_
	);
	LUT3 #(
		.INIT('h51)
	) name462 (
		_w476_,
		_w485_,
		_w486_,
		_w488_
	);
	LUT3 #(
		.INIT('h2b)
	) name463 (
		_w477_,
		_w478_,
		_w484_,
		_w489_
	);
	LUT4 #(
		.INIT('h00c1)
	) name464 (
		_w359_,
		_w398_,
		_w413_,
		_w464_,
		_w490_
	);
	LUT4 #(
		.INIT('hec00)
	) name465 (
		_w359_,
		_w414_,
		_w415_,
		_w464_,
		_w491_
	);
	LUT4 #(
		.INIT('h807f)
	) name466 (
		_w351_,
		_w338_,
		_w358_,
		_w424_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w416_,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h01)
	) name468 (
		_w491_,
		_w490_,
		_w493_,
		_w494_
	);
	LUT4 #(
		.INIT('hd400)
	) name469 (
		_w477_,
		_w478_,
		_w484_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h002b)
	) name470 (
		_w477_,
		_w478_,
		_w484_,
		_w494_,
		_w496_
	);
	LUT4 #(
		.INIT('h2bd4)
	) name471 (
		_w477_,
		_w478_,
		_w484_,
		_w494_,
		_w497_
	);
	LUT4 #(
		.INIT('ha956)
	) name472 (
		_w477_,
		_w461_,
		_w398_,
		_w420_,
		_w498_
	);
	LUT2 #(
		.INIT('h6)
	) name473 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('h7100)
	) name474 (
		_w365_,
		_w475_,
		_w485_,
		_w499_,
		_w500_
	);
	LUT3 #(
		.INIT('h56)
	) name475 (
		\a[7] ,
		\a[22] ,
		_w39_,
		_w501_
	);
	LUT4 #(
		.INIT('h007f)
	) name476 (
		_w351_,
		_w338_,
		_w358_,
		_w501_,
		_w502_
	);
	LUT3 #(
		.INIT('h57)
	) name477 (
		_w106_,
		_w68_,
		_w116_,
		_w503_
	);
	LUT4 #(
		.INIT('h0777)
	) name478 (
		_w106_,
		_w79_,
		_w71_,
		_w72_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT4 #(
		.INIT('h0777)
	) name480 (
		_w134_,
		_w54_,
		_w79_,
		_w77_,
		_w506_
	);
	LUT4 #(
		.INIT('h153f)
	) name481 (
		_w121_,
		_w134_,
		_w106_,
		_w125_,
		_w507_
	);
	LUT4 #(
		.INIT('h4000)
	) name482 (
		_w99_,
		_w394_,
		_w506_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('h37)
	) name483 (
		_w206_,
		_w106_,
		_w100_,
		_w509_
	);
	LUT4 #(
		.INIT('h135f)
	) name484 (
		_w82_,
		_w54_,
		_w96_,
		_w72_,
		_w510_
	);
	LUT3 #(
		.INIT('h40)
	) name485 (
		_w144_,
		_w509_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h0040)
	) name486 (
		_w117_,
		_w159_,
		_w442_,
		_w256_,
		_w512_
	);
	LUT4 #(
		.INIT('h8000)
	) name487 (
		_w511_,
		_w505_,
		_w512_,
		_w508_,
		_w513_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name488 (
		_w46_,
		_w82_,
		_w95_,
		_w68_,
		_w514_
	);
	LUT3 #(
		.INIT('h57)
	) name489 (
		_w88_,
		_w82_,
		_w91_,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT3 #(
		.INIT('h40)
	) name491 (
		_w46_,
		_w102_,
		_w70_,
		_w517_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name492 (
		_w46_,
		_w102_,
		_w70_,
		_w98_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		_w153_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h0100)
	) name494 (
		_w156_,
		_w101_,
		_w153_,
		_w518_,
		_w520_
	);
	LUT4 #(
		.INIT('h135f)
	) name495 (
		_w88_,
		_w54_,
		_w79_,
		_w125_,
		_w521_
	);
	LUT3 #(
		.INIT('h20)
	) name496 (
		_w186_,
		_w126_,
		_w521_,
		_w522_
	);
	LUT4 #(
		.INIT('h8000)
	) name497 (
		_w196_,
		_w201_,
		_w520_,
		_w522_,
		_w523_
	);
	LUT3 #(
		.INIT('h01)
	) name498 (
		_w110_,
		_w157_,
		_w311_,
		_w524_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name499 (
		_w46_,
		_w91_,
		_w70_,
		_w62_,
		_w525_
	);
	LUT4 #(
		.INIT('h153f)
	) name500 (
		_w77_,
		_w96_,
		_w116_,
		_w100_,
		_w526_
	);
	LUT3 #(
		.INIT('h80)
	) name501 (
		_w265_,
		_w525_,
		_w526_,
		_w527_
	);
	LUT4 #(
		.INIT('h37bf)
	) name502 (
		_w46_,
		_w53_,
		_w82_,
		_w116_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w244_,
		_w528_,
		_w529_
	);
	LUT3 #(
		.INIT('h57)
	) name504 (
		_w121_,
		_w113_,
		_w79_,
		_w530_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name505 (
		_w46_,
		_w53_,
		_w76_,
		_w91_,
		_w531_
	);
	LUT4 #(
		.INIT('h153f)
	) name506 (
		_w106_,
		_w77_,
		_w62_,
		_w72_,
		_w532_
	);
	LUT3 #(
		.INIT('h80)
	) name507 (
		_w531_,
		_w530_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w529_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('h8000)
	) name509 (
		_w524_,
		_w527_,
		_w529_,
		_w533_,
		_w535_
	);
	LUT4 #(
		.INIT('h8000)
	) name510 (
		_w513_,
		_w516_,
		_w523_,
		_w535_,
		_w536_
	);
	LUT4 #(
		.INIT('h135f)
	) name511 (
		_w134_,
		_w85_,
		_w96_,
		_w98_,
		_w537_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		_w137_,
		_w537_,
		_w538_
	);
	LUT3 #(
		.INIT('h37)
	) name513 (
		_w82_,
		_w77_,
		_w62_,
		_w539_
	);
	LUT4 #(
		.INIT('h37bf)
	) name514 (
		_w46_,
		_w53_,
		_w79_,
		_w91_,
		_w540_
	);
	LUT4 #(
		.INIT('h0008)
	) name515 (
		_w539_,
		_w540_,
		_w108_,
		_w347_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		_w538_,
		_w541_,
		_w542_
	);
	LUT3 #(
		.INIT('h01)
	) name517 (
		_w132_,
		_w181_,
		_w163_,
		_w543_
	);
	LUT4 #(
		.INIT('h0777)
	) name518 (
		_w76_,
		_w85_,
		_w77_,
		_w72_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		_w270_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w543_,
		_w545_,
		_w546_
	);
	LUT4 #(
		.INIT('h153f)
	) name521 (
		_w88_,
		_w54_,
		_w102_,
		_w68_,
		_w547_
	);
	LUT3 #(
		.INIT('h40)
	) name522 (
		_w219_,
		_w317_,
		_w547_,
		_w548_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name523 (
		_w46_,
		_w95_,
		_w79_,
		_w102_,
		_w549_
	);
	LUT3 #(
		.INIT('h1f)
	) name524 (
		_w206_,
		_w91_,
		_w71_,
		_w550_
	);
	LUT4 #(
		.INIT('h37bf)
	) name525 (
		_w46_,
		_w70_,
		_w68_,
		_w98_,
		_w551_
	);
	LUT4 #(
		.INIT('h135f)
	) name526 (
		_w121_,
		_w85_,
		_w91_,
		_w68_,
		_w552_
	);
	LUT4 #(
		.INIT('h8000)
	) name527 (
		_w551_,
		_w552_,
		_w549_,
		_w550_,
		_w553_
	);
	LUT4 #(
		.INIT('h8000)
	) name528 (
		_w548_,
		_w543_,
		_w545_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		_w542_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('h135f)
	) name530 (
		_w88_,
		_w113_,
		_w79_,
		_w77_,
		_w556_
	);
	LUT4 #(
		.INIT('h0400)
	) name531 (
		_w145_,
		_w330_,
		_w89_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		_w221_,
		_w451_,
		_w558_
	);
	LUT4 #(
		.INIT('h153f)
	) name533 (
		_w54_,
		_w59_,
		_w77_,
		_w125_,
		_w559_
	);
	LUT3 #(
		.INIT('h10)
	) name534 (
		_w339_,
		_w184_,
		_w559_,
		_w560_
	);
	LUT3 #(
		.INIT('h80)
	) name535 (
		_w143_,
		_w394_,
		_w506_,
		_w561_
	);
	LUT4 #(
		.INIT('h8000)
	) name536 (
		_w557_,
		_w558_,
		_w560_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('h0777)
	) name537 (
		_w88_,
		_w82_,
		_w96_,
		_w116_,
		_w563_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w198_,
		_w563_,
		_w564_
	);
	LUT3 #(
		.INIT('h01)
	) name539 (
		_w144_,
		_w194_,
		_w517_,
		_w565_
	);
	LUT3 #(
		.INIT('h80)
	) name540 (
		_w105_,
		_w565_,
		_w564_,
		_w566_
	);
	LUT3 #(
		.INIT('h01)
	) name541 (
		_w386_,
		_w115_,
		_w178_,
		_w567_
	);
	LUT3 #(
		.INIT('h57)
	) name542 (
		_w54_,
		_w68_,
		_w100_,
		_w568_
	);
	LUT4 #(
		.INIT('h0777)
	) name543 (
		_w206_,
		_w121_,
		_w76_,
		_w96_,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		_w567_,
		_w570_,
		_w571_
	);
	LUT4 #(
		.INIT('h0777)
	) name546 (
		_w88_,
		_w76_,
		_w85_,
		_w125_,
		_w572_
	);
	LUT3 #(
		.INIT('h57)
	) name547 (
		_w206_,
		_w88_,
		_w77_,
		_w573_
	);
	LUT3 #(
		.INIT('h37)
	) name548 (
		_w88_,
		_w134_,
		_w85_,
		_w574_
	);
	LUT4 #(
		.INIT('h0777)
	) name549 (
		_w85_,
		_w79_,
		_w71_,
		_w100_,
		_w575_
	);
	LUT4 #(
		.INIT('h8000)
	) name550 (
		_w572_,
		_w574_,
		_w575_,
		_w573_,
		_w576_
	);
	LUT3 #(
		.INIT('h80)
	) name551 (
		_w567_,
		_w570_,
		_w576_,
		_w577_
	);
	LUT3 #(
		.INIT('h80)
	) name552 (
		_w562_,
		_w566_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		_w555_,
		_w578_,
		_w579_
	);
	LUT4 #(
		.INIT('h5444)
	) name554 (
		_w322_,
		_w536_,
		_w555_,
		_w578_,
		_w580_
	);
	LUT4 #(
		.INIT('h393c)
	) name555 (
		\a[7] ,
		\a[8] ,
		\a[22] ,
		_w39_,
		_w581_
	);
	LUT4 #(
		.INIT('h007f)
	) name556 (
		_w351_,
		_w338_,
		_w358_,
		_w581_,
		_w582_
	);
	LUT3 #(
		.INIT('h4d)
	) name557 (
		_w502_,
		_w580_,
		_w582_,
		_w583_
	);
	LUT4 #(
		.INIT('h00c1)
	) name558 (
		_w359_,
		_w398_,
		_w413_,
		_w363_,
		_w584_
	);
	LUT4 #(
		.INIT('hec00)
	) name559 (
		_w359_,
		_w414_,
		_w415_,
		_w363_,
		_w585_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name560 (
		_w366_,
		_w351_,
		_w338_,
		_w358_,
		_w586_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w416_,
		_w586_,
		_w587_
	);
	LUT3 #(
		.INIT('h01)
	) name562 (
		_w585_,
		_w584_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w583_,
		_w588_,
		_w589_
	);
	LUT3 #(
		.INIT('h6f)
	) name564 (
		_w193_,
		_w424_,
		_w468_,
		_w590_
	);
	LUT4 #(
		.INIT('h4ff2)
	) name565 (
		_w193_,
		_w464_,
		_w264_,
		_w322_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name566 (
		_w590_,
		_w591_,
		_w592_
	);
	LUT3 #(
		.INIT('h7b)
	) name567 (
		_w398_,
		_w462_,
		_w419_,
		_w593_
	);
	LUT4 #(
		.INIT('h3dbc)
	) name568 (
		_w366_,
		_w193_,
		_w460_,
		_w398_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('h8000)
	) name570 (
		_w590_,
		_w591_,
		_w593_,
		_w594_,
		_w596_
	);
	LUT4 #(
		.INIT('h0777)
	) name571 (
		_w590_,
		_w591_,
		_w593_,
		_w594_,
		_w597_
	);
	LUT4 #(
		.INIT('h7888)
	) name572 (
		_w590_,
		_w591_,
		_w593_,
		_w594_,
		_w598_
	);
	LUT4 #(
		.INIT('h00c1)
	) name573 (
		_w359_,
		_w398_,
		_w413_,
		_w361_,
		_w599_
	);
	LUT4 #(
		.INIT('hec00)
	) name574 (
		_w359_,
		_w414_,
		_w415_,
		_w361_,
		_w600_
	);
	LUT4 #(
		.INIT('h7f80)
	) name575 (
		_w351_,
		_w338_,
		_w358_,
		_w363_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		_w416_,
		_w601_,
		_w602_
	);
	LUT3 #(
		.INIT('h01)
	) name577 (
		_w600_,
		_w599_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h9)
	) name578 (
		_w583_,
		_w588_,
		_w604_
	);
	LUT4 #(
		.INIT('he800)
	) name579 (
		_w592_,
		_w595_,
		_w603_,
		_w604_,
		_w605_
	);
	LUT4 #(
		.INIT('he11e)
	) name580 (
		_w193_,
		_w323_,
		_w362_,
		_w364_,
		_w606_
	);
	LUT2 #(
		.INIT('h9)
	) name581 (
		_w472_,
		_w474_,
		_w607_
	);
	LUT4 #(
		.INIT('h011f)
	) name582 (
		_w589_,
		_w605_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h6)
	) name583 (
		_w485_,
		_w487_,
		_w609_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w608_,
		_w609_,
		_w610_
	);
	LUT4 #(
		.INIT('h00c1)
	) name585 (
		_w359_,
		_w398_,
		_w413_,
		_w581_,
		_w611_
	);
	LUT4 #(
		.INIT('hec00)
	) name586 (
		_w359_,
		_w414_,
		_w415_,
		_w581_,
		_w612_
	);
	LUT4 #(
		.INIT('h7f80)
	) name587 (
		_w351_,
		_w338_,
		_w358_,
		_w361_,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		_w416_,
		_w613_,
		_w614_
	);
	LUT3 #(
		.INIT('h01)
	) name589 (
		_w612_,
		_w611_,
		_w614_,
		_w615_
	);
	LUT3 #(
		.INIT('h6f)
	) name590 (
		_w366_,
		_w398_,
		_w462_,
		_w616_
	);
	LUT4 #(
		.INIT('h6e76)
	) name591 (
		_w193_,
		_w460_,
		_w398_,
		_w363_,
		_w617_
	);
	LUT3 #(
		.INIT('h01)
	) name592 (
		_w117_,
		_w135_,
		_w372_,
		_w618_
	);
	LUT4 #(
		.INIT('h153f)
	) name593 (
		_w88_,
		_w77_,
		_w125_,
		_w72_,
		_w619_
	);
	LUT3 #(
		.INIT('h10)
	) name594 (
		_w152_,
		_w64_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('h153f)
	) name595 (
		_w206_,
		_w54_,
		_w98_,
		_w71_,
		_w621_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		_w407_,
		_w621_,
		_w622_
	);
	LUT3 #(
		.INIT('h80)
	) name597 (
		_w620_,
		_w622_,
		_w618_,
		_w623_
	);
	LUT4 #(
		.INIT('h135f)
	) name598 (
		_w54_,
		_w79_,
		_w91_,
		_w71_,
		_w624_
	);
	LUT3 #(
		.INIT('h80)
	) name599 (
		_w174_,
		_w123_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		_w511_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w623_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name602 (
		_w87_,
		_w46_,
		_w125_,
		_w100_,
		_w628_
	);
	LUT4 #(
		.INIT('h1000)
	) name603 (
		_w252_,
		_w185_,
		_w199_,
		_w628_,
		_w629_
	);
	LUT4 #(
		.INIT('h0777)
	) name604 (
		_w88_,
		_w91_,
		_w77_,
		_w72_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w236_,
		_w630_,
		_w631_
	);
	LUT3 #(
		.INIT('h04)
	) name606 (
		_w209_,
		_w572_,
		_w178_,
		_w632_
	);
	LUT3 #(
		.INIT('h80)
	) name607 (
		_w631_,
		_w632_,
		_w629_,
		_w633_
	);
	LUT3 #(
		.INIT('h37)
	) name608 (
		_w113_,
		_w71_,
		_w100_,
		_w634_
	);
	LUT4 #(
		.INIT('h135f)
	) name609 (
		_w53_,
		_w121_,
		_w113_,
		_w116_,
		_w635_
	);
	LUT3 #(
		.INIT('h40)
	) name610 (
		_w310_,
		_w635_,
		_w634_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w166_,
		_w636_,
		_w637_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name612 (
		_w46_,
		_w53_,
		_w134_,
		_w125_,
		_w638_
	);
	LUT3 #(
		.INIT('h10)
	) name613 (
		_w132_,
		_w83_,
		_w638_,
		_w639_
	);
	LUT4 #(
		.INIT('h0777)
	) name614 (
		_w91_,
		_w96_,
		_w68_,
		_w71_,
		_w640_
	);
	LUT4 #(
		.INIT('h8000)
	) name615 (
		_w551_,
		_w151_,
		_w431_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		_w639_,
		_w641_,
		_w642_
	);
	LUT4 #(
		.INIT('h135f)
	) name617 (
		_w54_,
		_w91_,
		_w68_,
		_w71_,
		_w643_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w393_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h0777)
	) name619 (
		_w121_,
		_w76_,
		_w134_,
		_w77_,
		_w645_
	);
	LUT3 #(
		.INIT('h80)
	) name620 (
		_w336_,
		_w370_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		_w644_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('h8000)
	) name622 (
		_w639_,
		_w641_,
		_w644_,
		_w646_,
		_w648_
	);
	LUT3 #(
		.INIT('h80)
	) name623 (
		_w633_,
		_w637_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		_w627_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h8000)
	) name625 (
		_w555_,
		_w578_,
		_w627_,
		_w649_,
		_w651_
	);
	LUT3 #(
		.INIT('h56)
	) name626 (
		\a[6] ,
		\a[22] ,
		_w38_,
		_w652_
	);
	LUT4 #(
		.INIT('h007f)
	) name627 (
		_w351_,
		_w338_,
		_w358_,
		_w652_,
		_w653_
	);
	LUT3 #(
		.INIT('h01)
	) name628 (
		_w168_,
		_w218_,
		_w137_,
		_w654_
	);
	LUT3 #(
		.INIT('h80)
	) name629 (
		_w453_,
		_w564_,
		_w654_,
		_w655_
	);
	LUT3 #(
		.INIT('h37)
	) name630 (
		_w79_,
		_w96_,
		_w98_,
		_w656_
	);
	LUT4 #(
		.INIT('h8000)
	) name631 (
		_w368_,
		_w250_,
		_w628_,
		_w656_,
		_w657_
	);
	LUT4 #(
		.INIT('h0777)
	) name632 (
		_w106_,
		_w79_,
		_w125_,
		_w71_,
		_w658_
	);
	LUT4 #(
		.INIT('h153f)
	) name633 (
		_w88_,
		_w76_,
		_w54_,
		_w59_,
		_w659_
	);
	LUT4 #(
		.INIT('h1000)
	) name634 (
		_w308_,
		_w347_,
		_w659_,
		_w658_,
		_w660_
	);
	LUT3 #(
		.INIT('h80)
	) name635 (
		_w636_,
		_w657_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		_w655_,
		_w661_,
		_w662_
	);
	LUT4 #(
		.INIT('h135f)
	) name637 (
		_w206_,
		_w54_,
		_w96_,
		_w98_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		_w547_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h135f)
	) name639 (
		_w88_,
		_w54_,
		_w91_,
		_w125_,
		_w665_
	);
	LUT4 #(
		.INIT('h0777)
	) name640 (
		_w76_,
		_w106_,
		_w54_,
		_w79_,
		_w666_
	);
	LUT3 #(
		.INIT('h80)
	) name641 (
		_w569_,
		_w666_,
		_w665_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		_w664_,
		_w667_,
		_w668_
	);
	LUT3 #(
		.INIT('h10)
	) name643 (
		_w132_,
		_w133_,
		_w291_,
		_w669_
	);
	LUT4 #(
		.INIT('h57df)
	) name644 (
		_w87_,
		_w46_,
		_w76_,
		_w91_,
		_w670_
	);
	LUT3 #(
		.INIT('h10)
	) name645 (
		_w238_,
		_w252_,
		_w670_,
		_w671_
	);
	LUT3 #(
		.INIT('h57)
	) name646 (
		_w121_,
		_w76_,
		_w100_,
		_w672_
	);
	LUT4 #(
		.INIT('h1000)
	) name647 (
		_w244_,
		_w103_,
		_w528_,
		_w672_,
		_w673_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		_w669_,
		_w671_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h153f)
	) name649 (
		_w106_,
		_w77_,
		_w116_,
		_w100_,
		_w675_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		_w232_,
		_w675_,
		_w676_
	);
	LUT4 #(
		.INIT('h1000)
	) name651 (
		_w407_,
		_w348_,
		_w324_,
		_w376_,
		_w677_
	);
	LUT3 #(
		.INIT('h1f)
	) name652 (
		_w76_,
		_w134_,
		_w77_,
		_w678_
	);
	LUT3 #(
		.INIT('h37)
	) name653 (
		_w91_,
		_w77_,
		_w100_,
		_w679_
	);
	LUT4 #(
		.INIT('h1000)
	) name654 (
		_w399_,
		_w110_,
		_w678_,
		_w679_,
		_w680_
	);
	LUT4 #(
		.INIT('h153f)
	) name655 (
		_w88_,
		_w79_,
		_w71_,
		_w72_,
		_w681_
	);
	LUT3 #(
		.INIT('h80)
	) name656 (
		_w186_,
		_w212_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h8000)
	) name657 (
		_w680_,
		_w676_,
		_w682_,
		_w677_,
		_w683_
	);
	LUT3 #(
		.INIT('h80)
	) name658 (
		_w668_,
		_w674_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		_w662_,
		_w684_,
		_w685_
	);
	LUT4 #(
		.INIT('h7000)
	) name660 (
		_w555_,
		_w578_,
		_w662_,
		_w684_,
		_w686_
	);
	LUT4 #(
		.INIT('h1303)
	) name661 (
		_w650_,
		_w651_,
		_w653_,
		_w686_,
		_w687_
	);
	LUT4 #(
		.INIT('h7f15)
	) name662 (
		_w615_,
		_w616_,
		_w617_,
		_w687_,
		_w688_
	);
	LUT3 #(
		.INIT('h6a)
	) name663 (
		_w536_,
		_w555_,
		_w578_,
		_w689_
	);
	LUT4 #(
		.INIT('h4111)
	) name664 (
		_w424_,
		_w536_,
		_w555_,
		_w578_,
		_w690_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name665 (
		_w322_,
		_w536_,
		_w555_,
		_w578_,
		_w691_
	);
	LUT4 #(
		.INIT('h5404)
	) name666 (
		_w502_,
		_w580_,
		_w690_,
		_w691_,
		_w692_
	);
	LUT4 #(
		.INIT('h02a2)
	) name667 (
		_w502_,
		_w580_,
		_w690_,
		_w691_,
		_w693_
	);
	LUT4 #(
		.INIT('ha959)
	) name668 (
		_w502_,
		_w580_,
		_w690_,
		_w691_,
		_w694_
	);
	LUT3 #(
		.INIT('h6f)
	) name669 (
		_w193_,
		_w464_,
		_w468_,
		_w695_
	);
	LUT4 #(
		.INIT('h4ff2)
	) name670 (
		_w193_,
		_w419_,
		_w264_,
		_w322_,
		_w696_
	);
	LUT4 #(
		.INIT('h4555)
	) name671 (
		_w692_,
		_w693_,
		_w695_,
		_w696_,
		_w697_
	);
	LUT3 #(
		.INIT('h69)
	) name672 (
		_w502_,
		_w580_,
		_w582_,
		_w698_
	);
	LUT4 #(
		.INIT('h6999)
	) name673 (
		_w362_,
		_w469_,
		_w470_,
		_w471_,
		_w699_
	);
	LUT4 #(
		.INIT('h7100)
	) name674 (
		_w688_,
		_w697_,
		_w698_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h008e)
	) name675 (
		_w688_,
		_w697_,
		_w698_,
		_w699_,
		_w701_
	);
	LUT4 #(
		.INIT('h8e71)
	) name676 (
		_w688_,
		_w697_,
		_w698_,
		_w699_,
		_w702_
	);
	LUT4 #(
		.INIT('h45ba)
	) name677 (
		_w596_,
		_w597_,
		_w603_,
		_w604_,
		_w703_
	);
	LUT3 #(
		.INIT('h45)
	) name678 (
		_w700_,
		_w701_,
		_w703_,
		_w704_
	);
	LUT4 #(
		.INIT('he11e)
	) name679 (
		_w589_,
		_w605_,
		_w606_,
		_w607_,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h6)
	) name681 (
		_w702_,
		_w703_,
		_w707_
	);
	LUT4 #(
		.INIT('h00c1)
	) name682 (
		_w359_,
		_w398_,
		_w413_,
		_w501_,
		_w708_
	);
	LUT4 #(
		.INIT('hec00)
	) name683 (
		_w359_,
		_w414_,
		_w415_,
		_w501_,
		_w709_
	);
	LUT4 #(
		.INIT('h7f80)
	) name684 (
		_w351_,
		_w338_,
		_w358_,
		_w581_,
		_w710_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		_w416_,
		_w710_,
		_w711_
	);
	LUT3 #(
		.INIT('h01)
	) name686 (
		_w709_,
		_w708_,
		_w711_,
		_w712_
	);
	LUT3 #(
		.INIT('h7b)
	) name687 (
		_w398_,
		_w462_,
		_w363_,
		_w713_
	);
	LUT4 #(
		.INIT('h6e76)
	) name688 (
		_w193_,
		_w460_,
		_w398_,
		_w361_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		_w713_,
		_w714_,
		_w715_
	);
	LUT3 #(
		.INIT('h80)
	) name690 (
		_w712_,
		_w713_,
		_w714_,
		_w716_
	);
	LUT3 #(
		.INIT('h15)
	) name691 (
		_w712_,
		_w713_,
		_w714_,
		_w717_
	);
	LUT3 #(
		.INIT('h6a)
	) name692 (
		_w712_,
		_w713_,
		_w714_,
		_w718_
	);
	LUT3 #(
		.INIT('h6f)
	) name693 (
		_w424_,
		_w322_,
		_w689_,
		_w719_
	);
	LUT4 #(
		.INIT('hc111)
	) name694 (
		_w322_,
		_w536_,
		_w555_,
		_w578_,
		_w720_
	);
	LUT4 #(
		.INIT('h8333)
	) name695 (
		_w322_,
		_w536_,
		_w555_,
		_w578_,
		_w721_
	);
	LUT3 #(
		.INIT('h1b)
	) name696 (
		_w464_,
		_w720_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		_w719_,
		_w722_,
		_w723_
	);
	LUT3 #(
		.INIT('h45)
	) name698 (
		_w716_,
		_w717_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h6a)
	) name699 (
		_w694_,
		_w695_,
		_w696_,
		_w725_
	);
	LUT4 #(
		.INIT('he800)
	) name700 (
		_w712_,
		_w715_,
		_w723_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('h6a95)
	) name701 (
		_w615_,
		_w616_,
		_w617_,
		_w687_,
		_w727_
	);
	LUT4 #(
		.INIT('h0017)
	) name702 (
		_w712_,
		_w715_,
		_w723_,
		_w725_,
		_w728_
	);
	LUT4 #(
		.INIT('h45ba)
	) name703 (
		_w716_,
		_w717_,
		_w723_,
		_w725_,
		_w729_
	);
	LUT3 #(
		.INIT('h51)
	) name704 (
		_w726_,
		_w727_,
		_w728_,
		_w730_
	);
	LUT2 #(
		.INIT('h6)
	) name705 (
		_w598_,
		_w603_,
		_w731_
	);
	LUT4 #(
		.INIT('h002b)
	) name706 (
		_w724_,
		_w725_,
		_w727_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('hd400)
	) name707 (
		_w724_,
		_w725_,
		_w727_,
		_w731_,
		_w733_
	);
	LUT3 #(
		.INIT('h96)
	) name708 (
		_w688_,
		_w697_,
		_w698_,
		_w734_
	);
	LUT3 #(
		.INIT('h54)
	) name709 (
		_w732_,
		_w733_,
		_w734_,
		_w735_
	);
	LUT4 #(
		.INIT('ha220)
	) name710 (
		_w707_,
		_w730_,
		_w731_,
		_w734_,
		_w736_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name711 (
		_w650_,
		_w651_,
		_w653_,
		_w686_,
		_w737_
	);
	LUT3 #(
		.INIT('h6f)
	) name712 (
		_w193_,
		_w419_,
		_w468_,
		_w738_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name713 (
		_w366_,
		_w193_,
		_w264_,
		_w322_,
		_w739_
	);
	LUT3 #(
		.INIT('h40)
	) name714 (
		_w737_,
		_w738_,
		_w739_,
		_w740_
	);
	LUT4 #(
		.INIT('h1555)
	) name715 (
		_w30_,
		_w351_,
		_w338_,
		_w358_,
		_w741_
	);
	LUT3 #(
		.INIT('h70)
	) name716 (
		_w627_,
		_w649_,
		_w741_,
		_w742_
	);
	LUT3 #(
		.INIT('h08)
	) name717 (
		_w627_,
		_w649_,
		_w741_,
		_w743_
	);
	LUT3 #(
		.INIT('h87)
	) name718 (
		_w627_,
		_w649_,
		_w741_,
		_w744_
	);
	LUT4 #(
		.INIT('h0777)
	) name719 (
		_w627_,
		_w649_,
		_w662_,
		_w684_,
		_w745_
	);
	LUT4 #(
		.INIT('h8000)
	) name720 (
		_w627_,
		_w649_,
		_w662_,
		_w684_,
		_w746_
	);
	LUT4 #(
		.INIT('h7888)
	) name721 (
		_w627_,
		_w649_,
		_w662_,
		_w684_,
		_w747_
	);
	LUT4 #(
		.INIT('h0243)
	) name722 (
		_w424_,
		_w579_,
		_w745_,
		_w746_,
		_w748_
	);
	LUT3 #(
		.INIT('h45)
	) name723 (
		_w742_,
		_w743_,
		_w748_,
		_w749_
	);
	LUT3 #(
		.INIT('h2a)
	) name724 (
		_w737_,
		_w738_,
		_w739_,
		_w750_
	);
	LUT3 #(
		.INIT('h95)
	) name725 (
		_w737_,
		_w738_,
		_w739_,
		_w751_
	);
	LUT3 #(
		.INIT('h54)
	) name726 (
		_w740_,
		_w749_,
		_w750_,
		_w752_
	);
	LUT3 #(
		.INIT('h6f)
	) name727 (
		_w464_,
		_w322_,
		_w689_,
		_w753_
	);
	LUT3 #(
		.INIT('h1b)
	) name728 (
		_w419_,
		_w720_,
		_w721_,
		_w754_
	);
	LUT3 #(
		.INIT('h6f)
	) name729 (
		_w366_,
		_w193_,
		_w468_,
		_w755_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name730 (
		_w193_,
		_w264_,
		_w322_,
		_w363_,
		_w756_
	);
	LUT4 #(
		.INIT('h8000)
	) name731 (
		_w753_,
		_w754_,
		_w755_,
		_w756_,
		_w757_
	);
	LUT4 #(
		.INIT('h0777)
	) name732 (
		_w753_,
		_w754_,
		_w755_,
		_w756_,
		_w758_
	);
	LUT4 #(
		.INIT('h7888)
	) name733 (
		_w753_,
		_w754_,
		_w755_,
		_w756_,
		_w759_
	);
	LUT3 #(
		.INIT('h7b)
	) name734 (
		_w398_,
		_w462_,
		_w361_,
		_w760_
	);
	LUT4 #(
		.INIT('h6e76)
	) name735 (
		_w193_,
		_w460_,
		_w398_,
		_w581_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		_w760_,
		_w761_,
		_w762_
	);
	LUT3 #(
		.INIT('h45)
	) name737 (
		_w757_,
		_w758_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h6)
	) name738 (
		_w718_,
		_w723_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w763_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('h007f)
	) name740 (
		_w351_,
		_w338_,
		_w358_,
		_w35_,
		_w766_
	);
	LUT3 #(
		.INIT('h70)
	) name741 (
		_w627_,
		_w649_,
		_w766_,
		_w767_
	);
	LUT3 #(
		.INIT('h08)
	) name742 (
		_w627_,
		_w649_,
		_w766_,
		_w768_
	);
	LUT3 #(
		.INIT('h87)
	) name743 (
		_w627_,
		_w649_,
		_w766_,
		_w769_
	);
	LUT3 #(
		.INIT('h6f)
	) name744 (
		_w424_,
		_w579_,
		_w747_,
		_w770_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name745 (
		_w464_,
		_w579_,
		_w650_,
		_w685_,
		_w771_
	);
	LUT4 #(
		.INIT('h4555)
	) name746 (
		_w767_,
		_w768_,
		_w770_,
		_w771_,
		_w772_
	);
	LUT4 #(
		.INIT('h00c1)
	) name747 (
		_w359_,
		_w398_,
		_w413_,
		_w652_,
		_w773_
	);
	LUT4 #(
		.INIT('hec00)
	) name748 (
		_w359_,
		_w414_,
		_w415_,
		_w652_,
		_w774_
	);
	LUT4 #(
		.INIT('h7f80)
	) name749 (
		_w351_,
		_w338_,
		_w358_,
		_w501_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w416_,
		_w775_,
		_w776_
	);
	LUT3 #(
		.INIT('h01)
	) name751 (
		_w774_,
		_w773_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w772_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h9)
	) name753 (
		_w772_,
		_w777_,
		_w779_
	);
	LUT3 #(
		.INIT('h6f)
	) name754 (
		_w193_,
		_w363_,
		_w468_,
		_w780_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name755 (
		_w193_,
		_w264_,
		_w322_,
		_w361_,
		_w781_
	);
	LUT3 #(
		.INIT('h6f)
	) name756 (
		_w419_,
		_w322_,
		_w689_,
		_w782_
	);
	LUT3 #(
		.INIT('h1b)
	) name757 (
		_w366_,
		_w720_,
		_w721_,
		_w783_
	);
	LUT4 #(
		.INIT('h8000)
	) name758 (
		_w780_,
		_w781_,
		_w782_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h0777)
	) name759 (
		_w780_,
		_w781_,
		_w782_,
		_w783_,
		_w785_
	);
	LUT4 #(
		.INIT('h7888)
	) name760 (
		_w780_,
		_w781_,
		_w782_,
		_w783_,
		_w786_
	);
	LUT3 #(
		.INIT('h7b)
	) name761 (
		_w398_,
		_w462_,
		_w581_,
		_w787_
	);
	LUT4 #(
		.INIT('h6e76)
	) name762 (
		_w193_,
		_w460_,
		_w398_,
		_w501_,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w787_,
		_w788_,
		_w789_
	);
	LUT3 #(
		.INIT('h45)
	) name764 (
		_w784_,
		_w785_,
		_w789_,
		_w790_
	);
	LUT3 #(
		.INIT('h51)
	) name765 (
		_w778_,
		_w779_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w763_,
		_w764_,
		_w792_
	);
	LUT2 #(
		.INIT('h9)
	) name767 (
		_w763_,
		_w764_,
		_w793_
	);
	LUT3 #(
		.INIT('h54)
	) name768 (
		_w765_,
		_w791_,
		_w792_,
		_w794_
	);
	LUT4 #(
		.INIT('h1051)
	) name769 (
		_w752_,
		_w763_,
		_w764_,
		_w791_,
		_w795_
	);
	LUT2 #(
		.INIT('h6)
	) name770 (
		_w727_,
		_w729_,
		_w796_
	);
	LUT4 #(
		.INIT('h8a08)
	) name771 (
		_w752_,
		_w763_,
		_w764_,
		_w791_,
		_w797_
	);
	LUT4 #(
		.INIT('h999a)
	) name772 (
		_w752_,
		_w765_,
		_w791_,
		_w792_,
		_w798_
	);
	LUT4 #(
		.INIT('h51ae)
	) name773 (
		_w726_,
		_w727_,
		_w728_,
		_w731_,
		_w799_
	);
	LUT2 #(
		.INIT('h9)
	) name774 (
		_w734_,
		_w799_,
		_w800_
	);
	LUT4 #(
		.INIT('h0071)
	) name775 (
		_w752_,
		_w794_,
		_w796_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h6)
	) name776 (
		_w744_,
		_w748_,
		_w802_
	);
	LUT3 #(
		.INIT('h60)
	) name777 (
		_w759_,
		_w762_,
		_w802_,
		_w803_
	);
	LUT4 #(
		.INIT('h007f)
	) name778 (
		_w351_,
		_w338_,
		_w358_,
		_w32_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		_w208_,
		_w456_,
		_w805_
	);
	LUT4 #(
		.INIT('h0001)
	) name780 (
		_w271_,
		_w107_,
		_w178_,
		_w300_,
		_w806_
	);
	LUT3 #(
		.INIT('h01)
	) name781 (
		_w218_,
		_w219_,
		_w99_,
		_w807_
	);
	LUT4 #(
		.INIT('h135f)
	) name782 (
		_w88_,
		_w54_,
		_w79_,
		_w72_,
		_w808_
	);
	LUT4 #(
		.INIT('h4000)
	) name783 (
		_w140_,
		_w65_,
		_w74_,
		_w808_,
		_w809_
	);
	LUT4 #(
		.INIT('h8000)
	) name784 (
		_w807_,
		_w805_,
		_w806_,
		_w809_,
		_w810_
	);
	LUT4 #(
		.INIT('h47ff)
	) name785 (
		_w87_,
		_w46_,
		_w95_,
		_w59_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w432_,
		_w811_,
		_w812_
	);
	LUT4 #(
		.INIT('h0777)
	) name787 (
		_w106_,
		_w68_,
		_w71_,
		_w100_,
		_w813_
	);
	LUT4 #(
		.INIT('h0777)
	) name788 (
		_w206_,
		_w88_,
		_w59_,
		_w71_,
		_w814_
	);
	LUT3 #(
		.INIT('h80)
	) name789 (
		_w429_,
		_w814_,
		_w813_,
		_w815_
	);
	LUT3 #(
		.INIT('h80)
	) name790 (
		_w326_,
		_w812_,
		_w815_,
		_w816_
	);
	LUT3 #(
		.INIT('h01)
	) name791 (
		_w386_,
		_w110_,
		_w372_,
		_w817_
	);
	LUT4 #(
		.INIT('h27ff)
	) name792 (
		_w46_,
		_w76_,
		_w113_,
		_w70_,
		_w818_
	);
	LUT3 #(
		.INIT('h37)
	) name793 (
		_w76_,
		_w77_,
		_w125_,
		_w819_
	);
	LUT3 #(
		.INIT('h80)
	) name794 (
		_w670_,
		_w819_,
		_w818_,
		_w820_
	);
	LUT4 #(
		.INIT('h37bf)
	) name795 (
		_w46_,
		_w53_,
		_w102_,
		_w125_,
		_w821_
	);
	LUT3 #(
		.INIT('h57)
	) name796 (
		_w88_,
		_w91_,
		_w62_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		_w821_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('h0777)
	) name798 (
		_w206_,
		_w85_,
		_w79_,
		_w77_,
		_w824_
	);
	LUT4 #(
		.INIT('h1000)
	) name799 (
		_w108_,
		_w347_,
		_w574_,
		_w824_,
		_w825_
	);
	LUT4 #(
		.INIT('h8000)
	) name800 (
		_w817_,
		_w820_,
		_w823_,
		_w825_,
		_w826_
	);
	LUT3 #(
		.INIT('h80)
	) name801 (
		_w810_,
		_w816_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('hd5c0)
	) name802 (
		_w424_,
		_w627_,
		_w649_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		_w804_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		_w804_,
		_w828_,
		_w830_
	);
	LUT2 #(
		.INIT('h9)
	) name805 (
		_w804_,
		_w828_,
		_w831_
	);
	LUT3 #(
		.INIT('h6f)
	) name806 (
		_w464_,
		_w579_,
		_w747_,
		_w832_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name807 (
		_w419_,
		_w579_,
		_w650_,
		_w685_,
		_w833_
	);
	LUT4 #(
		.INIT('h4555)
	) name808 (
		_w829_,
		_w830_,
		_w832_,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('h5001)
	) name809 (
		_w30_,
		_w359_,
		_w398_,
		_w413_,
		_w835_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name810 (
		_w30_,
		_w359_,
		_w414_,
		_w415_,
		_w836_
	);
	LUT4 #(
		.INIT('h7f80)
	) name811 (
		_w351_,
		_w338_,
		_w358_,
		_w652_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name812 (
		_w416_,
		_w837_,
		_w838_
	);
	LUT3 #(
		.INIT('h01)
	) name813 (
		_w836_,
		_w835_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w834_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h9)
	) name815 (
		_w834_,
		_w839_,
		_w841_
	);
	LUT3 #(
		.INIT('h6f)
	) name816 (
		_w193_,
		_w361_,
		_w468_,
		_w842_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name817 (
		_w193_,
		_w264_,
		_w322_,
		_w581_,
		_w843_
	);
	LUT3 #(
		.INIT('h6f)
	) name818 (
		_w366_,
		_w322_,
		_w689_,
		_w844_
	);
	LUT3 #(
		.INIT('h1b)
	) name819 (
		_w363_,
		_w720_,
		_w721_,
		_w845_
	);
	LUT4 #(
		.INIT('h8000)
	) name820 (
		_w842_,
		_w843_,
		_w844_,
		_w845_,
		_w846_
	);
	LUT4 #(
		.INIT('h0777)
	) name821 (
		_w842_,
		_w843_,
		_w844_,
		_w845_,
		_w847_
	);
	LUT4 #(
		.INIT('h7888)
	) name822 (
		_w842_,
		_w843_,
		_w844_,
		_w845_,
		_w848_
	);
	LUT3 #(
		.INIT('h7b)
	) name823 (
		_w398_,
		_w462_,
		_w501_,
		_w849_
	);
	LUT4 #(
		.INIT('h6e76)
	) name824 (
		_w193_,
		_w460_,
		_w398_,
		_w652_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w849_,
		_w850_,
		_w851_
	);
	LUT3 #(
		.INIT('h45)
	) name826 (
		_w846_,
		_w847_,
		_w851_,
		_w852_
	);
	LUT3 #(
		.INIT('h96)
	) name827 (
		_w759_,
		_w762_,
		_w802_,
		_w853_
	);
	LUT4 #(
		.INIT('h4d00)
	) name828 (
		_w834_,
		_w839_,
		_w852_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h9)
	) name829 (
		_w749_,
		_w751_,
		_w855_
	);
	LUT3 #(
		.INIT('he0)
	) name830 (
		_w803_,
		_w854_,
		_w855_,
		_w856_
	);
	LUT3 #(
		.INIT('h01)
	) name831 (
		_w803_,
		_w854_,
		_w855_,
		_w857_
	);
	LUT3 #(
		.INIT('h1e)
	) name832 (
		_w803_,
		_w854_,
		_w855_,
		_w858_
	);
	LUT2 #(
		.INIT('h9)
	) name833 (
		_w791_,
		_w793_,
		_w859_
	);
	LUT3 #(
		.INIT('h45)
	) name834 (
		_w856_,
		_w857_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h6)
	) name835 (
		_w796_,
		_w798_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		_w416_,
		_w32_,
		_w863_
	);
	LUT4 #(
		.INIT('h5440)
	) name838 (
		_w359_,
		_w398_,
		_w413_,
		_w32_,
		_w864_
	);
	LUT4 #(
		.INIT('h1555)
	) name839 (
		_w424_,
		_w810_,
		_w816_,
		_w826_,
		_w865_
	);
	LUT3 #(
		.INIT('h70)
	) name840 (
		_w627_,
		_w649_,
		_w865_,
		_w866_
	);
	LUT3 #(
		.INIT('h2a)
	) name841 (
		_w464_,
		_w627_,
		_w649_,
		_w867_
	);
	LUT4 #(
		.INIT('h00f8)
	) name842 (
		_w627_,
		_w649_,
		_w827_,
		_w865_,
		_w868_
	);
	LUT4 #(
		.INIT('h2022)
	) name843 (
		_w864_,
		_w866_,
		_w867_,
		_w868_,
		_w869_
	);
	LUT4 #(
		.INIT('h00c1)
	) name844 (
		_w359_,
		_w398_,
		_w413_,
		_w35_,
		_w870_
	);
	LUT4 #(
		.INIT('hec00)
	) name845 (
		_w359_,
		_w414_,
		_w415_,
		_w35_,
		_w871_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name846 (
		_w30_,
		_w351_,
		_w338_,
		_w358_,
		_w872_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w416_,
		_w872_,
		_w873_
	);
	LUT3 #(
		.INIT('h01)
	) name848 (
		_w871_,
		_w870_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		_w869_,
		_w874_,
		_w875_
	);
	LUT3 #(
		.INIT('h7b)
	) name850 (
		_w193_,
		_w468_,
		_w581_,
		_w876_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name851 (
		_w193_,
		_w264_,
		_w322_,
		_w501_,
		_w877_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		_w876_,
		_w877_,
		_w878_
	);
	LUT3 #(
		.INIT('h7b)
	) name853 (
		_w398_,
		_w462_,
		_w652_,
		_w879_
	);
	LUT4 #(
		.INIT('h3dbc)
	) name854 (
		_w30_,
		_w193_,
		_w460_,
		_w398_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT4 #(
		.INIT('h8000)
	) name856 (
		_w876_,
		_w877_,
		_w879_,
		_w880_,
		_w882_
	);
	LUT4 #(
		.INIT('h0777)
	) name857 (
		_w876_,
		_w877_,
		_w879_,
		_w880_,
		_w883_
	);
	LUT4 #(
		.INIT('h7888)
	) name858 (
		_w876_,
		_w877_,
		_w879_,
		_w880_,
		_w884_
	);
	LUT3 #(
		.INIT('h6f)
	) name859 (
		_w322_,
		_w363_,
		_w689_,
		_w885_
	);
	LUT3 #(
		.INIT('h1b)
	) name860 (
		_w361_,
		_w720_,
		_w721_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w885_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h6)
	) name862 (
		_w869_,
		_w874_,
		_w888_
	);
	LUT4 #(
		.INIT('he800)
	) name863 (
		_w878_,
		_w881_,
		_w887_,
		_w888_,
		_w889_
	);
	LUT3 #(
		.INIT('h6a)
	) name864 (
		_w769_,
		_w770_,
		_w771_,
		_w890_
	);
	LUT2 #(
		.INIT('h6)
	) name865 (
		_w786_,
		_w789_,
		_w891_
	);
	LUT4 #(
		.INIT('h011f)
	) name866 (
		_w875_,
		_w889_,
		_w890_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h9)
	) name867 (
		_w779_,
		_w790_,
		_w893_
	);
	LUT4 #(
		.INIT('h51ae)
	) name868 (
		_w840_,
		_w841_,
		_w852_,
		_w853_,
		_w894_
	);
	LUT3 #(
		.INIT('h2b)
	) name869 (
		_w892_,
		_w893_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h6)
	) name870 (
		_w858_,
		_w859_,
		_w896_
	);
	LUT3 #(
		.INIT('h06)
	) name871 (
		_w858_,
		_w859_,
		_w895_,
		_w897_
	);
	LUT3 #(
		.INIT('h6a)
	) name872 (
		_w831_,
		_w832_,
		_w833_,
		_w898_
	);
	LUT4 #(
		.INIT('h00c1)
	) name873 (
		_w359_,
		_w398_,
		_w413_,
		_w32_,
		_w899_
	);
	LUT4 #(
		.INIT('hec00)
	) name874 (
		_w359_,
		_w414_,
		_w415_,
		_w32_,
		_w900_
	);
	LUT4 #(
		.INIT('h7f80)
	) name875 (
		_w351_,
		_w338_,
		_w358_,
		_w35_,
		_w901_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		_w416_,
		_w901_,
		_w902_
	);
	LUT3 #(
		.INIT('h01)
	) name877 (
		_w900_,
		_w899_,
		_w902_,
		_w903_
	);
	LUT3 #(
		.INIT('h6f)
	) name878 (
		_w419_,
		_w579_,
		_w747_,
		_w904_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name879 (
		_w366_,
		_w579_,
		_w650_,
		_w685_,
		_w905_
	);
	LUT4 #(
		.INIT('h9a99)
	) name880 (
		_w864_,
		_w866_,
		_w867_,
		_w868_,
		_w906_
	);
	LUT4 #(
		.INIT('h157f)
	) name881 (
		_w903_,
		_w904_,
		_w905_,
		_w906_,
		_w907_
	);
	LUT4 #(
		.INIT('h60f6)
	) name882 (
		_w848_,
		_w851_,
		_w898_,
		_w907_,
		_w908_
	);
	LUT3 #(
		.INIT('h90)
	) name883 (
		_w841_,
		_w852_,
		_w908_,
		_w909_
	);
	LUT3 #(
		.INIT('h06)
	) name884 (
		_w841_,
		_w852_,
		_w908_,
		_w910_
	);
	LUT3 #(
		.INIT('h69)
	) name885 (
		_w841_,
		_w852_,
		_w908_,
		_w911_
	);
	LUT4 #(
		.INIT('he11e)
	) name886 (
		_w875_,
		_w889_,
		_w890_,
		_w891_,
		_w912_
	);
	LUT3 #(
		.INIT('h45)
	) name887 (
		_w909_,
		_w910_,
		_w912_,
		_w913_
	);
	LUT3 #(
		.INIT('h69)
	) name888 (
		_w892_,
		_w893_,
		_w894_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w913_,
		_w914_,
		_w915_
	);
	LUT3 #(
		.INIT('h6f)
	) name890 (
		_w322_,
		_w361_,
		_w689_,
		_w916_
	);
	LUT3 #(
		.INIT('h1b)
	) name891 (
		_w581_,
		_w720_,
		_w721_,
		_w917_
	);
	LUT3 #(
		.INIT('h7b)
	) name892 (
		_w193_,
		_w468_,
		_w501_,
		_w918_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name893 (
		_w193_,
		_w264_,
		_w322_,
		_w652_,
		_w919_
	);
	LUT4 #(
		.INIT('h8000)
	) name894 (
		_w916_,
		_w917_,
		_w918_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		_w462_,
		_w32_,
		_w921_
	);
	LUT4 #(
		.INIT('h0e08)
	) name896 (
		_w193_,
		_w460_,
		_w398_,
		_w32_,
		_w922_
	);
	LUT4 #(
		.INIT('h1555)
	) name897 (
		_w419_,
		_w810_,
		_w816_,
		_w826_,
		_w923_
	);
	LUT3 #(
		.INIT('h70)
	) name898 (
		_w627_,
		_w649_,
		_w923_,
		_w924_
	);
	LUT3 #(
		.INIT('h2a)
	) name899 (
		_w366_,
		_w627_,
		_w649_,
		_w925_
	);
	LUT4 #(
		.INIT('h00f8)
	) name900 (
		_w627_,
		_w649_,
		_w827_,
		_w923_,
		_w926_
	);
	LUT3 #(
		.INIT('h45)
	) name901 (
		_w924_,
		_w925_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		_w922_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h0777)
	) name903 (
		_w916_,
		_w917_,
		_w918_,
		_w919_,
		_w929_
	);
	LUT4 #(
		.INIT('h7888)
	) name904 (
		_w916_,
		_w917_,
		_w918_,
		_w919_,
		_w930_
	);
	LUT3 #(
		.INIT('h51)
	) name905 (
		_w920_,
		_w928_,
		_w929_,
		_w931_
	);
	LUT4 #(
		.INIT('h1555)
	) name906 (
		_w464_,
		_w810_,
		_w816_,
		_w826_,
		_w932_
	);
	LUT3 #(
		.INIT('h70)
	) name907 (
		_w627_,
		_w649_,
		_w932_,
		_w933_
	);
	LUT3 #(
		.INIT('h2a)
	) name908 (
		_w419_,
		_w627_,
		_w649_,
		_w934_
	);
	LUT4 #(
		.INIT('h00f8)
	) name909 (
		_w627_,
		_w649_,
		_w827_,
		_w932_,
		_w935_
	);
	LUT3 #(
		.INIT('h45)
	) name910 (
		_w933_,
		_w934_,
		_w935_,
		_w936_
	);
	LUT3 #(
		.INIT('h6f)
	) name911 (
		_w366_,
		_w579_,
		_w747_,
		_w937_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name912 (
		_w363_,
		_w579_,
		_w650_,
		_w685_,
		_w938_
	);
	LUT3 #(
		.INIT('h80)
	) name913 (
		_w936_,
		_w937_,
		_w938_,
		_w939_
	);
	LUT3 #(
		.INIT('h15)
	) name914 (
		_w936_,
		_w937_,
		_w938_,
		_w940_
	);
	LUT3 #(
		.INIT('h6a)
	) name915 (
		_w936_,
		_w937_,
		_w938_,
		_w941_
	);
	LUT3 #(
		.INIT('h6f)
	) name916 (
		_w30_,
		_w398_,
		_w462_,
		_w942_
	);
	LUT4 #(
		.INIT('h6e76)
	) name917 (
		_w193_,
		_w460_,
		_w398_,
		_w35_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		_w942_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('h45)
	) name919 (
		_w939_,
		_w940_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h6)
	) name920 (
		_w884_,
		_w887_,
		_w946_
	);
	LUT4 #(
		.INIT('h45ba)
	) name921 (
		_w882_,
		_w883_,
		_w887_,
		_w888_,
		_w947_
	);
	LUT4 #(
		.INIT('h7100)
	) name922 (
		_w931_,
		_w945_,
		_w946_,
		_w947_,
		_w948_
	);
	LUT4 #(
		.INIT('h008e)
	) name923 (
		_w931_,
		_w945_,
		_w946_,
		_w947_,
		_w949_
	);
	LUT4 #(
		.INIT('h8e71)
	) name924 (
		_w931_,
		_w945_,
		_w946_,
		_w947_,
		_w950_
	);
	LUT4 #(
		.INIT('h9669)
	) name925 (
		_w848_,
		_w851_,
		_w898_,
		_w907_,
		_w951_
	);
	LUT3 #(
		.INIT('h45)
	) name926 (
		_w948_,
		_w949_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h6)
	) name927 (
		_w911_,
		_w912_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name928 (
		_w952_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h9)
	) name929 (
		_w952_,
		_w953_,
		_w955_
	);
	LUT3 #(
		.INIT('h6f)
	) name930 (
		_w363_,
		_w579_,
		_w747_,
		_w956_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name931 (
		_w361_,
		_w579_,
		_w650_,
		_w685_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		_w956_,
		_w957_,
		_w958_
	);
	LUT3 #(
		.INIT('h7b)
	) name933 (
		_w193_,
		_w468_,
		_w652_,
		_w959_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name934 (
		_w30_,
		_w193_,
		_w264_,
		_w322_,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('h8000)
	) name936 (
		_w956_,
		_w957_,
		_w959_,
		_w960_,
		_w962_
	);
	LUT4 #(
		.INIT('h0777)
	) name937 (
		_w956_,
		_w957_,
		_w959_,
		_w960_,
		_w963_
	);
	LUT4 #(
		.INIT('h7888)
	) name938 (
		_w956_,
		_w957_,
		_w959_,
		_w960_,
		_w964_
	);
	LUT3 #(
		.INIT('h6f)
	) name939 (
		_w322_,
		_w581_,
		_w689_,
		_w965_
	);
	LUT3 #(
		.INIT('h1b)
	) name940 (
		_w501_,
		_w720_,
		_w721_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		_w965_,
		_w966_,
		_w967_
	);
	LUT3 #(
		.INIT('h45)
	) name942 (
		_w962_,
		_w963_,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('ha880)
	) name943 (
		_w863_,
		_w958_,
		_w961_,
		_w967_,
		_w969_
	);
	LUT2 #(
		.INIT('h6)
	) name944 (
		_w928_,
		_w930_,
		_w970_
	);
	LUT4 #(
		.INIT('h0115)
	) name945 (
		_w863_,
		_w958_,
		_w961_,
		_w967_,
		_w971_
	);
	LUT4 #(
		.INIT('h6566)
	) name946 (
		_w863_,
		_w962_,
		_w963_,
		_w967_,
		_w972_
	);
	LUT4 #(
		.INIT('h6a95)
	) name947 (
		_w903_,
		_w904_,
		_w905_,
		_w906_,
		_w973_
	);
	LUT4 #(
		.INIT('h00b2)
	) name948 (
		_w863_,
		_w968_,
		_w970_,
		_w973_,
		_w974_
	);
	LUT4 #(
		.INIT('h4d00)
	) name949 (
		_w863_,
		_w968_,
		_w970_,
		_w973_,
		_w975_
	);
	LUT4 #(
		.INIT('hae51)
	) name950 (
		_w969_,
		_w970_,
		_w971_,
		_w973_,
		_w976_
	);
	LUT3 #(
		.INIT('h96)
	) name951 (
		_w931_,
		_w945_,
		_w946_,
		_w977_
	);
	LUT3 #(
		.INIT('h45)
	) name952 (
		_w974_,
		_w975_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h6)
	) name953 (
		_w950_,
		_w951_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w978_,
		_w979_,
		_w981_
	);
	LUT2 #(
		.INIT('h6)
	) name956 (
		_w976_,
		_w977_,
		_w982_
	);
	LUT3 #(
		.INIT('h7b)
	) name957 (
		_w398_,
		_w462_,
		_w35_,
		_w983_
	);
	LUT4 #(
		.INIT('h6e76)
	) name958 (
		_w193_,
		_w460_,
		_w398_,
		_w32_,
		_w984_
	);
	LUT4 #(
		.INIT('h6000)
	) name959 (
		_w922_,
		_w927_,
		_w983_,
		_w984_,
		_w985_
	);
	LUT4 #(
		.INIT('h1555)
	) name960 (
		_w366_,
		_w810_,
		_w816_,
		_w826_,
		_w986_
	);
	LUT3 #(
		.INIT('h70)
	) name961 (
		_w627_,
		_w649_,
		_w986_,
		_w987_
	);
	LUT3 #(
		.INIT('h2a)
	) name962 (
		_w363_,
		_w627_,
		_w649_,
		_w988_
	);
	LUT4 #(
		.INIT('h00f8)
	) name963 (
		_w627_,
		_w649_,
		_w827_,
		_w986_,
		_w989_
	);
	LUT3 #(
		.INIT('h45)
	) name964 (
		_w987_,
		_w988_,
		_w989_,
		_w990_
	);
	LUT3 #(
		.INIT('h6f)
	) name965 (
		_w361_,
		_w579_,
		_w747_,
		_w991_
	);
	LUT4 #(
		.INIT('h4ff2)
	) name966 (
		_w579_,
		_w581_,
		_w650_,
		_w685_,
		_w992_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		_w991_,
		_w992_,
		_w993_
	);
	LUT3 #(
		.INIT('h80)
	) name968 (
		_w990_,
		_w991_,
		_w992_,
		_w994_
	);
	LUT3 #(
		.INIT('h15)
	) name969 (
		_w990_,
		_w991_,
		_w992_,
		_w995_
	);
	LUT3 #(
		.INIT('h6a)
	) name970 (
		_w990_,
		_w991_,
		_w992_,
		_w996_
	);
	LUT3 #(
		.INIT('h6f)
	) name971 (
		_w322_,
		_w501_,
		_w689_,
		_w997_
	);
	LUT3 #(
		.INIT('h1b)
	) name972 (
		_w652_,
		_w720_,
		_w721_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		_w997_,
		_w998_,
		_w999_
	);
	LUT4 #(
		.INIT('h9666)
	) name974 (
		_w922_,
		_w927_,
		_w983_,
		_w984_,
		_w1000_
	);
	LUT4 #(
		.INIT('he800)
	) name975 (
		_w990_,
		_w993_,
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h6)
	) name976 (
		_w941_,
		_w944_,
		_w1002_
	);
	LUT3 #(
		.INIT('he0)
	) name977 (
		_w985_,
		_w1001_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h6)
	) name978 (
		_w970_,
		_w972_,
		_w1004_
	);
	LUT3 #(
		.INIT('h01)
	) name979 (
		_w985_,
		_w1001_,
		_w1002_,
		_w1005_
	);
	LUT3 #(
		.INIT('h1e)
	) name980 (
		_w985_,
		_w1001_,
		_w1002_,
		_w1006_
	);
	LUT3 #(
		.INIT('h51)
	) name981 (
		_w1003_,
		_w1004_,
		_w1005_,
		_w1007_
	);
	LUT2 #(
		.INIT('h2)
	) name982 (
		_w982_,
		_w1007_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0078)
	) name983 (
		_w216_,
		_w263_,
		_w322_,
		_w32_,
		_w1009_
	);
	LUT3 #(
		.INIT('h01)
	) name984 (
		_w193_,
		_w323_,
		_w1009_,
		_w1010_
	);
	LUT4 #(
		.INIT('hd500)
	) name985 (
		_w361_,
		_w627_,
		_w649_,
		_w827_,
		_w1011_
	);
	LUT4 #(
		.INIT('h8095)
	) name986 (
		_w363_,
		_w627_,
		_w649_,
		_w827_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w1011_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h6)
	) name988 (
		_w1010_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('hd500)
	) name989 (
		_w581_,
		_w627_,
		_w649_,
		_w827_,
		_w1015_
	);
	LUT4 #(
		.INIT('h8095)
	) name990 (
		_w361_,
		_w627_,
		_w649_,
		_w827_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT3 #(
		.INIT('h6f)
	) name992 (
		_w501_,
		_w579_,
		_w747_,
		_w1018_
	);
	LUT4 #(
		.INIT('h73ce)
	) name993 (
		_w579_,
		_w650_,
		_w652_,
		_w685_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w1018_,
		_w1019_,
		_w1020_
	);
	LUT3 #(
		.INIT('h80)
	) name995 (
		_w1017_,
		_w1018_,
		_w1019_,
		_w1021_
	);
	LUT3 #(
		.INIT('h15)
	) name996 (
		_w1017_,
		_w1018_,
		_w1019_,
		_w1022_
	);
	LUT3 #(
		.INIT('h6a)
	) name997 (
		_w1017_,
		_w1018_,
		_w1019_,
		_w1023_
	);
	LUT3 #(
		.INIT('h6f)
	) name998 (
		_w30_,
		_w322_,
		_w689_,
		_w1024_
	);
	LUT3 #(
		.INIT('h35)
	) name999 (
		_w720_,
		_w721_,
		_w35_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT4 #(
		.INIT('ha880)
	) name1001 (
		_w1014_,
		_w1017_,
		_w1020_,
		_w1026_,
		_w1027_
	);
	LUT4 #(
		.INIT('h0115)
	) name1002 (
		_w1014_,
		_w1017_,
		_w1020_,
		_w1026_,
		_w1028_
	);
	LUT4 #(
		.INIT('h6566)
	) name1003 (
		_w1014_,
		_w1021_,
		_w1022_,
		_w1026_,
		_w1029_
	);
	LUT3 #(
		.INIT('h6f)
	) name1004 (
		_w579_,
		_w581_,
		_w747_,
		_w1030_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name1005 (
		_w501_,
		_w579_,
		_w650_,
		_w685_,
		_w1031_
	);
	LUT3 #(
		.INIT('h6f)
	) name1006 (
		_w322_,
		_w652_,
		_w689_,
		_w1032_
	);
	LUT3 #(
		.INIT('h1b)
	) name1007 (
		_w30_,
		_w720_,
		_w721_,
		_w1033_
	);
	LUT4 #(
		.INIT('h8000)
	) name1008 (
		_w1030_,
		_w1031_,
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('h0777)
	) name1009 (
		_w1030_,
		_w1031_,
		_w1032_,
		_w1033_,
		_w1035_
	);
	LUT4 #(
		.INIT('h7888)
	) name1010 (
		_w1030_,
		_w1031_,
		_w1032_,
		_w1033_,
		_w1036_
	);
	LUT3 #(
		.INIT('h7b)
	) name1011 (
		_w193_,
		_w468_,
		_w35_,
		_w1037_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name1012 (
		_w193_,
		_w264_,
		_w322_,
		_w32_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h6)
	) name1014 (
		_w1036_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h006a)
	) name1015 (
		_w536_,
		_w555_,
		_w578_,
		_w32_,
		_w1041_
	);
	LUT4 #(
		.INIT('hd500)
	) name1016 (
		_w501_,
		_w627_,
		_w649_,
		_w827_,
		_w1042_
	);
	LUT4 #(
		.INIT('h8095)
	) name1017 (
		_w581_,
		_w627_,
		_w649_,
		_w827_,
		_w1043_
	);
	LUT4 #(
		.INIT('h0002)
	) name1018 (
		_w580_,
		_w1041_,
		_w1042_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w1009_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h6)
	) name1020 (
		_w1009_,
		_w1044_,
		_w1046_
	);
	LUT3 #(
		.INIT('h6f)
	) name1021 (
		_w579_,
		_w652_,
		_w747_,
		_w1047_
	);
	LUT4 #(
		.INIT('h2ff4)
	) name1022 (
		_w30_,
		_w579_,
		_w650_,
		_w685_,
		_w1048_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT3 #(
		.INIT('h7b)
	) name1024 (
		_w322_,
		_w689_,
		_w35_,
		_w1050_
	);
	LUT3 #(
		.INIT('h35)
	) name1025 (
		_w720_,
		_w721_,
		_w32_,
		_w1051_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		_w1050_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h0777)
	) name1027 (
		_w1047_,
		_w1048_,
		_w1050_,
		_w1051_,
		_w1053_
	);
	LUT4 #(
		.INIT('h8000)
	) name1028 (
		_w1047_,
		_w1048_,
		_w1050_,
		_w1051_,
		_w1054_
	);
	LUT4 #(
		.INIT('h222d)
	) name1029 (
		_w580_,
		_w1041_,
		_w1042_,
		_w1043_,
		_w1055_
	);
	LUT4 #(
		.INIT('ha880)
	) name1030 (
		_w1046_,
		_w1049_,
		_w1052_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('h0009)
	) name1031 (
		_w1029_,
		_w1040_,
		_w1045_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h999a)
	) name1032 (
		_w1046_,
		_w1053_,
		_w1054_,
		_w1055_,
		_w1058_
	);
	LUT2 #(
		.INIT('h6)
	) name1033 (
		_w1023_,
		_w1026_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT4 #(
		.INIT('h5440)
	) name1035 (
		_w579_,
		_w650_,
		_w685_,
		_w32_,
		_w1061_
	);
	LUT4 #(
		.INIT('hd500)
	) name1036 (
		_w30_,
		_w627_,
		_w649_,
		_w827_,
		_w1062_
	);
	LUT4 #(
		.INIT('h8087)
	) name1037 (
		_w627_,
		_w649_,
		_w652_,
		_w827_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w1062_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		_w1061_,
		_w1064_,
		_w1065_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1040 (
		_w627_,
		_w649_,
		_w652_,
		_w827_,
		_w1066_
	);
	LUT4 #(
		.INIT('h8095)
	) name1041 (
		_w501_,
		_w627_,
		_w649_,
		_w827_,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1066_,
		_w1067_,
		_w1068_
	);
	LUT3 #(
		.INIT('h6f)
	) name1043 (
		_w30_,
		_w579_,
		_w747_,
		_w1069_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name1044 (
		_w579_,
		_w650_,
		_w685_,
		_w35_,
		_w1070_
	);
	LUT3 #(
		.INIT('h80)
	) name1045 (
		_w1068_,
		_w1069_,
		_w1070_,
		_w1071_
	);
	LUT3 #(
		.INIT('h15)
	) name1046 (
		_w1068_,
		_w1069_,
		_w1070_,
		_w1072_
	);
	LUT3 #(
		.INIT('h6a)
	) name1047 (
		_w1068_,
		_w1069_,
		_w1070_,
		_w1073_
	);
	LUT2 #(
		.INIT('h6)
	) name1048 (
		_w1065_,
		_w1073_,
		_w1074_
	);
	LUT4 #(
		.INIT('h1555)
	) name1049 (
		_w35_,
		_w810_,
		_w816_,
		_w826_,
		_w1075_
	);
	LUT4 #(
		.INIT('h0070)
	) name1050 (
		_w627_,
		_w649_,
		_w32_,
		_w1075_,
		_w1076_
	);
	LUT3 #(
		.INIT('h0d)
	) name1051 (
		_w747_,
		_w32_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h006a)
	) name1052 (
		_w30_,
		_w627_,
		_w649_,
		_w827_,
		_w1078_
	);
	LUT4 #(
		.INIT('h7000)
	) name1053 (
		_w627_,
		_w649_,
		_w35_,
		_w827_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		_w1077_,
		_w1080_,
		_w1081_
	);
	LUT3 #(
		.INIT('h7b)
	) name1056 (
		_w579_,
		_w747_,
		_w35_,
		_w1082_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name1057 (
		_w579_,
		_w650_,
		_w685_,
		_w32_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h6)
	) name1059 (
		_w1061_,
		_w1064_,
		_w1085_
	);
	LUT4 #(
		.INIT('ha880)
	) name1060 (
		_w1041_,
		_w1081_,
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1074_,
		_w1086_,
		_w1087_
	);
	LUT4 #(
		.INIT('h0115)
	) name1062 (
		_w1041_,
		_w1081_,
		_w1084_,
		_w1085_,
		_w1088_
	);
	LUT3 #(
		.INIT('h51)
	) name1063 (
		_w1071_,
		_w1065_,
		_w1072_,
		_w1089_
	);
	LUT3 #(
		.INIT('h1e)
	) name1064 (
		_w1053_,
		_w1054_,
		_w1055_,
		_w1090_
	);
	LUT3 #(
		.INIT('h07)
	) name1065 (
		_w1089_,
		_w1090_,
		_w1088_,
		_w1091_
	);
	LUT4 #(
		.INIT('h7770)
	) name1066 (
		_w1058_,
		_w1059_,
		_w1089_,
		_w1090_,
		_w1092_
	);
	LUT4 #(
		.INIT('h1055)
	) name1067 (
		_w1060_,
		_w1087_,
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT4 #(
		.INIT('h6660)
	) name1068 (
		_w1029_,
		_w1040_,
		_w1045_,
		_w1056_,
		_w1094_
	);
	LUT3 #(
		.INIT('h45)
	) name1069 (
		_w1027_,
		_w1028_,
		_w1040_,
		_w1095_
	);
	LUT3 #(
		.INIT('h6f)
	) name1070 (
		_w30_,
		_w193_,
		_w468_,
		_w1096_
	);
	LUT4 #(
		.INIT('h7c3e)
	) name1071 (
		_w193_,
		_w264_,
		_w322_,
		_w35_,
		_w1097_
	);
	LUT4 #(
		.INIT('h8000)
	) name1072 (
		_w1010_,
		_w1013_,
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h0777)
	) name1073 (
		_w1010_,
		_w1013_,
		_w1096_,
		_w1097_,
		_w1099_
	);
	LUT4 #(
		.INIT('h7888)
	) name1074 (
		_w1010_,
		_w1013_,
		_w1096_,
		_w1097_,
		_w1100_
	);
	LUT2 #(
		.INIT('h6)
	) name1075 (
		_w921_,
		_w1100_,
		_w1101_
	);
	LUT3 #(
		.INIT('h45)
	) name1076 (
		_w1034_,
		_w1035_,
		_w1039_,
		_w1102_
	);
	LUT2 #(
		.INIT('h6)
	) name1077 (
		_w996_,
		_w999_,
		_w1103_
	);
	LUT3 #(
		.INIT('h69)
	) name1078 (
		_w1102_,
		_w1103_,
		_w1101_,
		_w1104_
	);
	LUT3 #(
		.INIT('h45)
	) name1079 (
		_w1094_,
		_w1095_,
		_w1104_,
		_w1105_
	);
	LUT3 #(
		.INIT('h31)
	) name1080 (
		_w921_,
		_w1098_,
		_w1099_,
		_w1106_
	);
	LUT2 #(
		.INIT('h6)
	) name1081 (
		_w964_,
		_w967_,
		_w1107_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1082 (
		_w994_,
		_w995_,
		_w999_,
		_w1000_,
		_w1108_
	);
	LUT3 #(
		.INIT('h69)
	) name1083 (
		_w1106_,
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT3 #(
		.INIT('h2b)
	) name1084 (
		_w1102_,
		_w1103_,
		_w1101_,
		_w1110_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1085 (
		_w1109_,
		_w1110_,
		_w1095_,
		_w1104_,
		_w1111_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1086 (
		_w1057_,
		_w1093_,
		_w1105_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		_w1109_,
		_w1110_,
		_w1113_
	);
	LUT3 #(
		.INIT('h2b)
	) name1088 (
		_w1106_,
		_w1107_,
		_w1108_,
		_w1114_
	);
	LUT3 #(
		.INIT('h06)
	) name1089 (
		_w1004_,
		_w1006_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1113_,
		_w1115_,
		_w1116_
	);
	LUT3 #(
		.INIT('h90)
	) name1091 (
		_w1004_,
		_w1006_,
		_w1114_,
		_w1117_
	);
	LUT3 #(
		.INIT('h0b)
	) name1092 (
		_w982_,
		_w1007_,
		_w1117_,
		_w1118_
	);
	LUT4 #(
		.INIT('h1055)
	) name1093 (
		_w1008_,
		_w1112_,
		_w1116_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('h20a2)
	) name1094 (
		_w955_,
		_w978_,
		_w979_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		_w913_,
		_w914_,
		_w1121_
	);
	LUT2 #(
		.INIT('h9)
	) name1096 (
		_w913_,
		_w914_,
		_w1122_
	);
	LUT4 #(
		.INIT('h5501)
	) name1097 (
		_w915_,
		_w954_,
		_w1120_,
		_w1121_,
		_w1123_
	);
	LUT3 #(
		.INIT('h90)
	) name1098 (
		_w858_,
		_w859_,
		_w895_,
		_w1124_
	);
	LUT3 #(
		.INIT('h69)
	) name1099 (
		_w858_,
		_w859_,
		_w895_,
		_w1125_
	);
	LUT2 #(
		.INIT('h9)
	) name1100 (
		_w860_,
		_w861_,
		_w1126_
	);
	LUT4 #(
		.INIT('h4d00)
	) name1101 (
		_w895_,
		_w896_,
		_w1123_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('hae51)
	) name1102 (
		_w795_,
		_w796_,
		_w797_,
		_w800_,
		_w1128_
	);
	LUT4 #(
		.INIT('h0155)
	) name1103 (
		_w801_,
		_w862_,
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h0445)
	) name1104 (
		_w707_,
		_w730_,
		_w731_,
		_w734_,
		_w1130_
	);
	LUT4 #(
		.INIT('h999a)
	) name1105 (
		_w707_,
		_w732_,
		_w733_,
		_w734_,
		_w1131_
	);
	LUT2 #(
		.INIT('h9)
	) name1106 (
		_w704_,
		_w705_,
		_w1132_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1107 (
		_w707_,
		_w735_,
		_w1129_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name1108 (
		_w608_,
		_w609_,
		_w1134_
	);
	LUT2 #(
		.INIT('h9)
	) name1109 (
		_w608_,
		_w609_,
		_w1135_
	);
	LUT4 #(
		.INIT('h5501)
	) name1110 (
		_w610_,
		_w706_,
		_w1133_,
		_w1134_,
		_w1136_
	);
	LUT4 #(
		.INIT('h008e)
	) name1111 (
		_w365_,
		_w475_,
		_w485_,
		_w499_,
		_w1137_
	);
	LUT4 #(
		.INIT('h51ae)
	) name1112 (
		_w476_,
		_w485_,
		_w486_,
		_w499_,
		_w1138_
	);
	LUT4 #(
		.INIT('h0157)
	) name1113 (
		_w477_,
		_w461_,
		_w398_,
		_w420_,
		_w1139_
	);
	LUT4 #(
		.INIT('h5146)
	) name1114 (
		_w359_,
		_w398_,
		_w424_,
		_w413_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		_w481_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name1116 (
		_w481_,
		_w1140_,
		_w1142_
	);
	LUT2 #(
		.INIT('h9)
	) name1117 (
		_w481_,
		_w1140_,
		_w1143_
	);
	LUT2 #(
		.INIT('h9)
	) name1118 (
		_w1139_,
		_w1143_,
		_w1144_
	);
	LUT4 #(
		.INIT('hd400)
	) name1119 (
		_w489_,
		_w494_,
		_w498_,
		_w1144_,
		_w1145_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1120 (
		_w495_,
		_w496_,
		_w498_,
		_w1144_,
		_w1146_
	);
	LUT4 #(
		.INIT('h4d00)
	) name1121 (
		_w488_,
		_w499_,
		_w1136_,
		_w1146_,
		_w1147_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1122 (
		_w500_,
		_w1136_,
		_w1137_,
		_w1146_,
		_w1148_
	);
	LUT4 #(
		.INIT('h153f)
	) name1123 (
		_w106_,
		_w91_,
		_w77_,
		_w98_,
		_w1149_
	);
	LUT4 #(
		.INIT('h153f)
	) name1124 (
		_w206_,
		_w88_,
		_w134_,
		_w85_,
		_w1150_
	);
	LUT3 #(
		.INIT('h80)
	) name1125 (
		_w559_,
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		_w230_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h0777)
	) name1127 (
		_w88_,
		_w79_,
		_w91_,
		_w71_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		_w170_,
		_w1153_,
		_w1154_
	);
	LUT3 #(
		.INIT('h10)
	) name1129 (
		_w252_,
		_w181_,
		_w279_,
		_w1155_
	);
	LUT4 #(
		.INIT('h37bf)
	) name1130 (
		_w46_,
		_w95_,
		_w134_,
		_w62_,
		_w1156_
	);
	LUT3 #(
		.INIT('h10)
	) name1131 (
		_w176_,
		_w393_,
		_w1156_,
		_w1157_
	);
	LUT4 #(
		.INIT('h8000)
	) name1132 (
		_w342_,
		_w1157_,
		_w1154_,
		_w1155_,
		_w1158_
	);
	LUT3 #(
		.INIT('h80)
	) name1133 (
		_w313_,
		_w1152_,
		_w1158_,
		_w1159_
	);
	LUT3 #(
		.INIT('h1f)
	) name1134 (
		_w88_,
		_w54_,
		_w59_,
		_w1160_
	);
	LUT4 #(
		.INIT('h153f)
	) name1135 (
		_w121_,
		_w134_,
		_w77_,
		_w68_,
		_w1161_
	);
	LUT3 #(
		.INIT('h40)
	) name1136 (
		_w297_,
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT4 #(
		.INIT('h135f)
	) name1137 (
		_w88_,
		_w134_,
		_w62_,
		_w71_,
		_w1163_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w517_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name1139 (
		_w46_,
		_w53_,
		_w68_,
		_w116_,
		_w1165_
	);
	LUT3 #(
		.INIT('h80)
	) name1140 (
		_w292_,
		_w681_,
		_w1165_,
		_w1166_
	);
	LUT3 #(
		.INIT('h80)
	) name1141 (
		_w1162_,
		_w1164_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('h4000)
	) name1142 (
		_w158_,
		_w291_,
		_w503_,
		_w504_,
		_w1168_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name1143 (
		_w46_,
		_w59_,
		_w70_,
		_w116_,
		_w1169_
	);
	LUT4 #(
		.INIT('h4000)
	) name1144 (
		_w407_,
		_w528_,
		_w621_,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name1145 (
		_w46_,
		_w76_,
		_w70_,
		_w68_,
		_w1171_
	);
	LUT3 #(
		.INIT('h40)
	) name1146 (
		_w318_,
		_w436_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('h40)
	) name1147 (
		_w171_,
		_w165_,
		_w276_,
		_w1173_
	);
	LUT4 #(
		.INIT('h8000)
	) name1148 (
		_w1172_,
		_w1173_,
		_w1168_,
		_w1170_,
		_w1174_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		_w1167_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w1159_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w1148_,
		_w1176_,
		_w1177_
	);
	LUT4 #(
		.INIT('h0777)
	) name1152 (
		_w121_,
		_w62_,
		_w68_,
		_w71_,
		_w1178_
	);
	LUT4 #(
		.INIT('h8000)
	) name1153 (
		_w183_,
		_w195_,
		_w666_,
		_w1178_,
		_w1179_
	);
	LUT3 #(
		.INIT('h01)
	) name1154 (
		_w156_,
		_w247_,
		_w239_,
		_w1180_
	);
	LUT4 #(
		.INIT('h4000)
	) name1155 (
		_w111_,
		_w233_,
		_w292_,
		_w293_,
		_w1181_
	);
	LUT4 #(
		.INIT('h8000)
	) name1156 (
		_w538_,
		_w1180_,
		_w1179_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h8000)
	) name1157 (
		_w427_,
		_w430_,
		_w524_,
		_w527_,
		_w1183_
	);
	LUT4 #(
		.INIT('h8000)
	) name1158 (
		_w623_,
		_w626_,
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT3 #(
		.INIT('h06)
	) name1159 (
		_w1136_,
		_w1138_,
		_w1184_,
		_w1185_
	);
	LUT3 #(
		.INIT('h1e)
	) name1160 (
		_w706_,
		_w1133_,
		_w1135_,
		_w1186_
	);
	LUT4 #(
		.INIT('h37bf)
	) name1161 (
		_w46_,
		_w53_,
		_w59_,
		_w79_,
		_w1187_
	);
	LUT4 #(
		.INIT('h153f)
	) name1162 (
		_w134_,
		_w79_,
		_w96_,
		_w71_,
		_w1188_
	);
	LUT4 #(
		.INIT('h8000)
	) name1163 (
		_w1187_,
		_w528_,
		_w1169_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		_w1157_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		_w243_,
		_w666_,
		_w1191_
	);
	LUT4 #(
		.INIT('h135f)
	) name1166 (
		_w121_,
		_w62_,
		_w116_,
		_w71_,
		_w1192_
	);
	LUT3 #(
		.INIT('h10)
	) name1167 (
		_w347_,
		_w253_,
		_w1192_,
		_w1193_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		_w120_,
		_w1191_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		_w1190_,
		_w1194_,
		_w1195_
	);
	LUT4 #(
		.INIT('h0777)
	) name1170 (
		_w206_,
		_w54_,
		_w59_,
		_w77_,
		_w1196_
	);
	LUT4 #(
		.INIT('h0777)
	) name1171 (
		_w121_,
		_w134_,
		_w77_,
		_w68_,
		_w1197_
	);
	LUT4 #(
		.INIT('h4000)
	) name1172 (
		_w311_,
		_w544_,
		_w1197_,
		_w1196_,
		_w1198_
	);
	LUT4 #(
		.INIT('h0777)
	) name1173 (
		_w206_,
		_w121_,
		_w54_,
		_w72_,
		_w1199_
	);
	LUT3 #(
		.INIT('h10)
	) name1174 (
		_w249_,
		_w146_,
		_w1199_,
		_w1200_
	);
	LUT4 #(
		.INIT('h8000)
	) name1175 (
		_w129_,
		_w438_,
		_w1198_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h135f)
	) name1176 (
		_w121_,
		_w106_,
		_w79_,
		_w68_,
		_w1202_
	);
	LUT2 #(
		.INIT('h4)
	) name1177 (
		_w284_,
		_w1202_,
		_w1203_
	);
	LUT4 #(
		.INIT('h153f)
	) name1178 (
		_w88_,
		_w85_,
		_w91_,
		_w125_,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name1179 (
		_w301_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('h1000)
	) name1180 (
		_w252_,
		_w301_,
		_w172_,
		_w1204_,
		_w1206_
	);
	LUT2 #(
		.INIT('h8)
	) name1181 (
		_w1203_,
		_w1206_,
		_w1207_
	);
	LUT4 #(
		.INIT('h153f)
	) name1182 (
		_w88_,
		_w134_,
		_w96_,
		_w98_,
		_w1208_
	);
	LUT3 #(
		.INIT('h40)
	) name1183 (
		_w367_,
		_w388_,
		_w1208_,
		_w1209_
	);
	LUT3 #(
		.INIT('h80)
	) name1184 (
		_w105_,
		_w112_,
		_w1209_,
		_w1210_
	);
	LUT3 #(
		.INIT('h80)
	) name1185 (
		_w1201_,
		_w1207_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		_w1195_,
		_w1211_,
		_w1212_
	);
	LUT4 #(
		.INIT('h00e1)
	) name1187 (
		_w706_,
		_w1133_,
		_w1135_,
		_w1212_,
		_w1213_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1188 (
		_w736_,
		_w1129_,
		_w1130_,
		_w1132_,
		_w1214_
	);
	LUT4 #(
		.INIT('h777f)
	) name1189 (
		_w87_,
		_w46_,
		_w102_,
		_w100_,
		_w1215_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w169_,
		_w1215_,
		_w1216_
	);
	LUT3 #(
		.INIT('h80)
	) name1191 (
		_w1190_,
		_w1194_,
		_w1216_,
		_w1217_
	);
	LUT4 #(
		.INIT('h153f)
	) name1192 (
		_w206_,
		_w88_,
		_w79_,
		_w77_,
		_w1218_
	);
	LUT3 #(
		.INIT('h1f)
	) name1193 (
		_w88_,
		_w77_,
		_w100_,
		_w1219_
	);
	LUT3 #(
		.INIT('h80)
	) name1194 (
		_w210_,
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT3 #(
		.INIT('h40)
	) name1195 (
		_w184_,
		_w345_,
		_w376_,
		_w1221_
	);
	LUT3 #(
		.INIT('h80)
	) name1196 (
		_w1203_,
		_w1220_,
		_w1221_,
		_w1222_
	);
	LUT4 #(
		.INIT('h337f)
	) name1197 (
		_w46_,
		_w53_,
		_w91_,
		_w62_,
		_w1223_
	);
	LUT4 #(
		.INIT('h0777)
	) name1198 (
		_w85_,
		_w102_,
		_w96_,
		_w72_,
		_w1224_
	);
	LUT4 #(
		.INIT('h8000)
	) name1199 (
		_w572_,
		_w509_,
		_w1223_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('h57df)
	) name1200 (
		_w87_,
		_w46_,
		_w91_,
		_w62_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name1201 (
		_w311_,
		_w1226_,
		_w1227_
	);
	LUT3 #(
		.INIT('h80)
	) name1202 (
		_w807_,
		_w1227_,
		_w1225_,
		_w1228_
	);
	LUT3 #(
		.INIT('h80)
	) name1203 (
		_w1152_,
		_w1222_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		_w1217_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		_w1214_,
		_w1230_,
		_w1231_
	);
	LUT3 #(
		.INIT('h57)
	) name1206 (
		_w88_,
		_w59_,
		_w116_,
		_w1232_
	);
	LUT3 #(
		.INIT('h80)
	) name1207 (
		_w542_,
		_w554_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h1dff)
	) name1208 (
		_w87_,
		_w46_,
		_w95_,
		_w113_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name1209 (
		_w1234_,
		_w186_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		_w456_,
		_w628_,
		_w1236_
	);
	LUT3 #(
		.INIT('h10)
	) name1211 (
		_w107_,
		_w311_,
		_w824_,
		_w1237_
	);
	LUT3 #(
		.INIT('h80)
	) name1212 (
		_w1235_,
		_w1236_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		_w571_,
		_w1238_,
		_w1239_
	);
	LUT3 #(
		.INIT('h37)
	) name1214 (
		_w121_,
		_w59_,
		_w85_,
		_w1240_
	);
	LUT4 #(
		.INIT('h0777)
	) name1215 (
		_w82_,
		_w96_,
		_w116_,
		_w71_,
		_w1241_
	);
	LUT3 #(
		.INIT('h40)
	) name1216 (
		_w122_,
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT3 #(
		.INIT('h10)
	) name1217 (
		_w156_,
		_w266_,
		_w525_,
		_w1243_
	);
	LUT3 #(
		.INIT('h10)
	) name1218 (
		_w249_,
		_w146_,
		_w818_,
		_w1244_
	);
	LUT4 #(
		.INIT('h135f)
	) name1219 (
		_w82_,
		_w106_,
		_w71_,
		_w100_,
		_w1245_
	);
	LUT4 #(
		.INIT('h135f)
	) name1220 (
		_w206_,
		_w88_,
		_w96_,
		_w125_,
		_w1246_
	);
	LUT4 #(
		.INIT('h8000)
	) name1221 (
		_w375_,
		_w1156_,
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT4 #(
		.INIT('h8000)
	) name1222 (
		_w1243_,
		_w1244_,
		_w1242_,
		_w1247_,
		_w1248_
	);
	LUT3 #(
		.INIT('h80)
	) name1223 (
		_w571_,
		_w1238_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h8)
	) name1224 (
		_w1233_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('h06)
	) name1225 (
		_w1129_,
		_w1131_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h1e)
	) name1226 (
		_w862_,
		_w1127_,
		_w1128_,
		_w1252_
	);
	LUT4 #(
		.INIT('h0737)
	) name1227 (
		_w206_,
		_w121_,
		_w76_,
		_w54_,
		_w1253_
	);
	LUT3 #(
		.INIT('h40)
	) name1228 (
		_w284_,
		_w400_,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('h0777)
	) name1229 (
		_w106_,
		_w91_,
		_w116_,
		_w71_,
		_w1255_
	);
	LUT4 #(
		.INIT('h153f)
	) name1230 (
		_w206_,
		_w59_,
		_w85_,
		_w71_,
		_w1256_
	);
	LUT3 #(
		.INIT('h80)
	) name1231 (
		_w635_,
		_w1256_,
		_w1255_,
		_w1257_
	);
	LUT3 #(
		.INIT('h80)
	) name1232 (
		_w557_,
		_w1254_,
		_w1257_,
		_w1258_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name1233 (
		_w46_,
		_w82_,
		_w70_,
		_w125_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w551_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1235 (
		_w87_,
		_w46_,
		_w113_,
		_w59_,
		_w1261_
	);
	LUT3 #(
		.INIT('h10)
	) name1236 (
		_w339_,
		_w184_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('h80)
	) name1237 (
		_w280_,
		_w1260_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w136_,
		_w289_,
		_w1264_
	);
	LUT4 #(
		.INIT('h0001)
	) name1239 (
		_w386_,
		_w64_,
		_w169_,
		_w128_,
		_w1265_
	);
	LUT3 #(
		.INIT('h10)
	) name1240 (
		_w308_,
		_w347_,
		_w208_,
		_w1266_
	);
	LUT3 #(
		.INIT('h80)
	) name1241 (
		_w1264_,
		_w1265_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('h8000)
	) name1242 (
		_w513_,
		_w1263_,
		_w1267_,
		_w1258_,
		_w1268_
	);
	LUT4 #(
		.INIT('h00e1)
	) name1243 (
		_w862_,
		_w1127_,
		_w1128_,
		_w1268_,
		_w1269_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1244 (
		_w897_,
		_w1123_,
		_w1124_,
		_w1126_,
		_w1270_
	);
	LUT4 #(
		.INIT('h153f)
	) name1245 (
		_w88_,
		_w134_,
		_w54_,
		_w79_,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		_w1234_,
		_w1271_,
		_w1272_
	);
	LUT4 #(
		.INIT('h153f)
	) name1247 (
		_w121_,
		_w54_,
		_w102_,
		_w125_,
		_w1273_
	);
	LUT4 #(
		.INIT('h6fff)
	) name1248 (
		_w51_,
		_w52_,
		_w46_,
		_w116_,
		_w1274_
	);
	LUT3 #(
		.INIT('h80)
	) name1249 (
		_w429_,
		_w1273_,
		_w1274_,
		_w1275_
	);
	LUT4 #(
		.INIT('h8000)
	) name1250 (
		_w120_,
		_w1272_,
		_w680_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name1251 (
		_w219_,
		_w172_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name1252 (
		_w1276_,
		_w1277_,
		_w1278_
	);
	LUT4 #(
		.INIT('h153f)
	) name1253 (
		_w88_,
		_w85_,
		_w79_,
		_w98_,
		_w1279_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w73_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h153f)
	) name1255 (
		_w85_,
		_w77_,
		_w125_,
		_w100_,
		_w1281_
	);
	LUT3 #(
		.INIT('h10)
	) name1256 (
		_w339_,
		_w209_,
		_w1281_,
		_w1282_
	);
	LUT4 #(
		.INIT('h153f)
	) name1257 (
		_w206_,
		_w121_,
		_w62_,
		_w96_,
		_w1283_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		_w200_,
		_w1283_,
		_w1284_
	);
	LUT3 #(
		.INIT('h80)
	) name1259 (
		_w1280_,
		_w1282_,
		_w1284_,
		_w1285_
	);
	LUT4 #(
		.INIT('h0777)
	) name1260 (
		_w88_,
		_w134_,
		_w54_,
		_w72_,
		_w1286_
	);
	LUT4 #(
		.INIT('h135f)
	) name1261 (
		_w121_,
		_w113_,
		_w116_,
		_w71_,
		_w1287_
	);
	LUT4 #(
		.INIT('h8000)
	) name1262 (
		_w540_,
		_w186_,
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('haebf)
	) name1263 (
		_w51_,
		_w52_,
		_w79_,
		_w102_,
		_w1289_
	);
	LUT4 #(
		.INIT('h0100)
	) name1264 (
		_w80_,
		_w347_,
		_w103_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h80)
	) name1265 (
		_w277_,
		_w1288_,
		_w1290_,
		_w1291_
	);
	LUT3 #(
		.INIT('h80)
	) name1266 (
		_w546_,
		_w1285_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		_w1278_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name1268 (
		_w1270_,
		_w1293_,
		_w1294_
	);
	LUT4 #(
		.INIT('h135f)
	) name1269 (
		_w88_,
		_w82_,
		_w59_,
		_w77_,
		_w1295_
	);
	LUT4 #(
		.INIT('h1000)
	) name1270 (
		_w227_,
		_w110_,
		_w544_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h0800)
	) name1271 (
		_w328_,
		_w329_,
		_w144_,
		_w147_,
		_w1297_
	);
	LUT3 #(
		.INIT('h80)
	) name1272 (
		_w1205_,
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('hafff)
	) name1273 (
		_w51_,
		_w52_,
		_w46_,
		_w62_,
		_w1299_
	);
	LUT4 #(
		.INIT('h777f)
	) name1274 (
		_w87_,
		_w46_,
		_w102_,
		_w68_,
		_w1300_
	);
	LUT4 #(
		.INIT('h4000)
	) name1275 (
		_w164_,
		_w174_,
		_w1300_,
		_w1299_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		_w505_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h135f)
	) name1277 (
		_w88_,
		_w82_,
		_w79_,
		_w71_,
		_w1303_
	);
	LUT4 #(
		.INIT('h8000)
	) name1278 (
		_w335_,
		_w383_,
		_w634_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w117_,
		_w189_,
		_w1305_
	);
	LUT3 #(
		.INIT('h10)
	) name1280 (
		_w238_,
		_w252_,
		_w90_,
		_w1306_
	);
	LUT3 #(
		.INIT('h80)
	) name1281 (
		_w1304_,
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h8000)
	) name1282 (
		_w296_,
		_w1298_,
		_w1302_,
		_w1307_,
		_w1308_
	);
	LUT3 #(
		.INIT('h06)
	) name1283 (
		_w1123_,
		_w1125_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name1284 (
		_w247_,
		_w429_,
		_w1310_
	);
	LUT4 #(
		.INIT('h2000)
	) name1285 (
		_w394_,
		_w311_,
		_w506_,
		_w1226_,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT3 #(
		.INIT('h57)
	) name1287 (
		_w88_,
		_w134_,
		_w100_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w407_,
		_w1313_,
		_w1314_
	);
	LUT4 #(
		.INIT('h153f)
	) name1289 (
		_w121_,
		_w77_,
		_w68_,
		_w72_,
		_w1315_
	);
	LUT3 #(
		.INIT('h40)
	) name1290 (
		_w407_,
		_w1313_,
		_w1315_,
		_w1316_
	);
	LUT4 #(
		.INIT('h5557)
	) name1291 (
		_w121_,
		_w113_,
		_w79_,
		_w125_,
		_w1317_
	);
	LUT4 #(
		.INIT('h153f)
	) name1292 (
		_w88_,
		_w77_,
		_w100_,
		_w72_,
		_w1318_
	);
	LUT4 #(
		.INIT('h1000)
	) name1293 (
		_w132_,
		_w73_,
		_w1318_,
		_w1317_,
		_w1319_
	);
	LUT3 #(
		.INIT('h80)
	) name1294 (
		_w1254_,
		_w1316_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h8)
	) name1295 (
		_w1312_,
		_w1320_,
		_w1321_
	);
	LUT3 #(
		.INIT('h1f)
	) name1296 (
		_w82_,
		_w134_,
		_w106_,
		_w1322_
	);
	LUT4 #(
		.INIT('h0777)
	) name1297 (
		_w88_,
		_w82_,
		_w91_,
		_w71_,
		_w1323_
	);
	LUT4 #(
		.INIT('h1000)
	) name1298 (
		_w271_,
		_w300_,
		_w1323_,
		_w1322_,
		_w1324_
	);
	LUT4 #(
		.INIT('h37bf)
	) name1299 (
		_w46_,
		_w53_,
		_w102_,
		_w62_,
		_w1325_
	);
	LUT4 #(
		.INIT('h2000)
	) name1300 (
		_w572_,
		_w163_,
		_w254_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('h8000)
	) name1301 (
		_w511_,
		_w1304_,
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h80)
	) name1302 (
		_w542_,
		_w188_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name1303 (
		_w1321_,
		_w1328_,
		_w1329_
	);
	LUT4 #(
		.INIT('h00e1)
	) name1304 (
		_w954_,
		_w1120_,
		_w1122_,
		_w1329_,
		_w1330_
	);
	LUT4 #(
		.INIT('h9a99)
	) name1305 (
		_w955_,
		_w980_,
		_w981_,
		_w1119_,
		_w1331_
	);
	LUT4 #(
		.INIT('h37bf)
	) name1306 (
		_w46_,
		_w95_,
		_w59_,
		_w125_,
		_w1332_
	);
	LUT3 #(
		.INIT('h04)
	) name1307 (
		_w107_,
		_w1332_,
		_w115_,
		_w1333_
	);
	LUT3 #(
		.INIT('h10)
	) name1308 (
		_w132_,
		_w73_,
		_w195_,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name1309 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		_w249_,
		_w442_,
		_w1336_
	);
	LUT4 #(
		.INIT('h153f)
	) name1311 (
		_w88_,
		_w91_,
		_w77_,
		_w125_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name1312 (
		_w379_,
		_w1337_,
		_w1338_
	);
	LUT3 #(
		.INIT('h80)
	) name1313 (
		_w259_,
		_w1336_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h135f)
	) name1314 (
		_w95_,
		_w79_,
		_w102_,
		_w77_,
		_w1340_
	);
	LUT4 #(
		.INIT('h0100)
	) name1315 (
		_w252_,
		_w185_,
		_w164_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h135f)
	) name1316 (
		_w59_,
		_w96_,
		_w71_,
		_w72_,
		_w1342_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1317 (
		_w121_,
		_w54_,
		_w98_,
		_w355_,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name1319 (
		_w87_,
		_w91_,
		_w1345_
	);
	LUT4 #(
		.INIT('h0777)
	) name1320 (
		_w206_,
		_w85_,
		_w77_,
		_w100_,
		_w1346_
	);
	LUT3 #(
		.INIT('h10)
	) name1321 (
		_w64_,
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT3 #(
		.INIT('h80)
	) name1322 (
		_w1341_,
		_w1344_,
		_w1347_,
		_w1348_
	);
	LUT4 #(
		.INIT('h8000)
	) name1323 (
		_w1263_,
		_w1348_,
		_w1335_,
		_w1339_,
		_w1349_
	);
	LUT2 #(
		.INIT('h9)
	) name1324 (
		_w978_,
		_w979_,
		_w1350_
	);
	LUT3 #(
		.INIT('h80)
	) name1325 (
		_w299_,
		_w620_,
		_w1310_,
		_w1351_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1326 (
		_w46_,
		_w53_,
		_w113_,
		_w72_,
		_w1352_
	);
	LUT3 #(
		.INIT('h10)
	) name1327 (
		_w432_,
		_w517_,
		_w1352_,
		_w1353_
	);
	LUT3 #(
		.INIT('h80)
	) name1328 (
		_w294_,
		_w548_,
		_w1353_,
		_w1354_
	);
	LUT4 #(
		.INIT('h8000)
	) name1329 (
		_w1174_,
		_w1298_,
		_w1351_,
		_w1354_,
		_w1355_
	);
	LUT3 #(
		.INIT('h90)
	) name1330 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1356_
	);
	LUT3 #(
		.INIT('he8)
	) name1331 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1357_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1332 (
		_w954_,
		_w1120_,
		_w1122_,
		_w1329_,
		_w1358_
	);
	LUT4 #(
		.INIT('he11e)
	) name1333 (
		_w954_,
		_w1120_,
		_w1122_,
		_w1329_,
		_w1359_
	);
	LUT3 #(
		.INIT('h54)
	) name1334 (
		_w1330_,
		_w1357_,
		_w1358_,
		_w1360_
	);
	LUT3 #(
		.INIT('h90)
	) name1335 (
		_w1123_,
		_w1125_,
		_w1308_,
		_w1361_
	);
	LUT3 #(
		.INIT('h69)
	) name1336 (
		_w1123_,
		_w1125_,
		_w1308_,
		_w1362_
	);
	LUT3 #(
		.INIT('h54)
	) name1337 (
		_w1309_,
		_w1360_,
		_w1361_,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		_w1270_,
		_w1293_,
		_w1364_
	);
	LUT2 #(
		.INIT('h6)
	) name1339 (
		_w1270_,
		_w1293_,
		_w1365_
	);
	LUT3 #(
		.INIT('h54)
	) name1340 (
		_w1294_,
		_w1363_,
		_w1364_,
		_w1366_
	);
	LUT4 #(
		.INIT('he11e)
	) name1341 (
		_w862_,
		_w1127_,
		_w1128_,
		_w1268_,
		_w1367_
	);
	LUT4 #(
		.INIT('h1700)
	) name1342 (
		_w1270_,
		_w1293_,
		_w1363_,
		_w1367_,
		_w1368_
	);
	LUT3 #(
		.INIT('h69)
	) name1343 (
		_w1129_,
		_w1131_,
		_w1250_,
		_w1369_
	);
	LUT4 #(
		.INIT('h0155)
	) name1344 (
		_w1251_,
		_w1269_,
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1345 (
		_w1214_,
		_w1230_,
		_w1371_
	);
	LUT2 #(
		.INIT('h6)
	) name1346 (
		_w1214_,
		_w1230_,
		_w1372_
	);
	LUT3 #(
		.INIT('h54)
	) name1347 (
		_w1231_,
		_w1370_,
		_w1371_,
		_w1373_
	);
	LUT4 #(
		.INIT('he11e)
	) name1348 (
		_w706_,
		_w1133_,
		_w1135_,
		_w1212_,
		_w1374_
	);
	LUT4 #(
		.INIT('h1700)
	) name1349 (
		_w1214_,
		_w1230_,
		_w1370_,
		_w1374_,
		_w1375_
	);
	LUT3 #(
		.INIT('h69)
	) name1350 (
		_w1136_,
		_w1138_,
		_w1184_,
		_w1376_
	);
	LUT4 #(
		.INIT('h0155)
	) name1351 (
		_w1185_,
		_w1213_,
		_w1375_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		_w1148_,
		_w1176_,
		_w1378_
	);
	LUT2 #(
		.INIT('h6)
	) name1353 (
		_w1148_,
		_w1176_,
		_w1379_
	);
	LUT3 #(
		.INIT('h54)
	) name1354 (
		_w1177_,
		_w1377_,
		_w1378_,
		_w1380_
	);
	LUT4 #(
		.INIT('h0001)
	) name1355 (
		_w238_,
		_w271_,
		_w316_,
		_w168_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w1332_,
		_w572_,
		_w1382_
	);
	LUT3 #(
		.INIT('h02)
	) name1357 (
		_w371_,
		_w386_,
		_w64_,
		_w1383_
	);
	LUT3 #(
		.INIT('h80)
	) name1358 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT4 #(
		.INIT('h135f)
	) name1359 (
		_w88_,
		_w54_,
		_w59_,
		_w91_,
		_w1385_
	);
	LUT4 #(
		.INIT('h0040)
	) name1360 (
		_w224_,
		_w1187_,
		_w1385_,
		_w156_,
		_w1386_
	);
	LUT4 #(
		.INIT('h0010)
	) name1361 (
		_w407_,
		_w209_,
		_w514_,
		_w252_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h8000)
	) name1363 (
		_w538_,
		_w541_,
		_w639_,
		_w641_,
		_w1389_
	);
	LUT3 #(
		.INIT('h80)
	) name1364 (
		_w1384_,
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		_w1278_,
		_w1390_,
		_w1391_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1366 (
		\a[13] ,
		\a[14] ,
		\a[22] ,
		_w44_,
		_w1392_
	);
	LUT3 #(
		.INIT('h41)
	) name1367 (
		_w359_,
		_w414_,
		_w1392_,
		_w1393_
	);
	LUT4 #(
		.INIT('h32cd)
	) name1368 (
		_w1139_,
		_w1141_,
		_w1142_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h1e)
	) name1369 (
		_w1145_,
		_w1147_,
		_w1394_,
		_w1395_
	);
	LUT4 #(
		.INIT('h0154)
	) name1370 (
		_w1391_,
		_w1145_,
		_w1147_,
		_w1394_,
		_w1396_
	);
	LUT4 #(
		.INIT('h56a9)
	) name1371 (
		_w1391_,
		_w1145_,
		_w1147_,
		_w1394_,
		_w1397_
	);
	LUT4 #(
		.INIT('h1700)
	) name1372 (
		_w1148_,
		_w1176_,
		_w1377_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1373 (
		_w1148_,
		_w1176_,
		_w1377_,
		_w1397_,
		_w1399_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1374 (
		_w1177_,
		_w1377_,
		_w1378_,
		_w1397_,
		_w1400_
	);
	LUT4 #(
		.INIT('h6801)
	) name1375 (
		_w1148_,
		_w1176_,
		_w1377_,
		_w1397_,
		_w1401_
	);
	LUT3 #(
		.INIT('h1e)
	) name1376 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1402_
	);
	LUT3 #(
		.INIT('h90)
	) name1377 (
		_w1377_,
		_w1379_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1378 (
		_w1214_,
		_w1230_,
		_w1370_,
		_w1374_,
		_w1404_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1379 (
		_w1231_,
		_w1370_,
		_w1371_,
		_w1374_,
		_w1405_
	);
	LUT4 #(
		.INIT('h6801)
	) name1380 (
		_w1186_,
		_w1212_,
		_w1373_,
		_w1376_,
		_w1406_
	);
	LUT4 #(
		.INIT('h6801)
	) name1381 (
		_w1214_,
		_w1230_,
		_w1370_,
		_w1374_,
		_w1407_
	);
	LUT3 #(
		.INIT('h1e)
	) name1382 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1408_
	);
	LUT3 #(
		.INIT('h90)
	) name1383 (
		_w1370_,
		_w1372_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1384 (
		_w1270_,
		_w1293_,
		_w1363_,
		_w1367_,
		_w1410_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1385 (
		_w1294_,
		_w1363_,
		_w1364_,
		_w1367_,
		_w1411_
	);
	LUT4 #(
		.INIT('h6801)
	) name1386 (
		_w1252_,
		_w1268_,
		_w1366_,
		_w1369_,
		_w1412_
	);
	LUT4 #(
		.INIT('h6801)
	) name1387 (
		_w1270_,
		_w1293_,
		_w1363_,
		_w1367_,
		_w1413_
	);
	LUT2 #(
		.INIT('h9)
	) name1388 (
		_w1360_,
		_w1362_,
		_w1414_
	);
	LUT2 #(
		.INIT('h9)
	) name1389 (
		_w1357_,
		_w1359_,
		_w1415_
	);
	LUT3 #(
		.INIT('h06)
	) name1390 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1416_
	);
	LUT3 #(
		.INIT('h69)
	) name1391 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1417_
	);
	LUT3 #(
		.INIT('h69)
	) name1392 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1418_
	);
	LUT4 #(
		.INIT('h9f00)
	) name1393 (
		_w1357_,
		_w1359_,
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT4 #(
		.INIT('h066f)
	) name1394 (
		_w1360_,
		_w1362_,
		_w1415_,
		_w1419_,
		_w1420_
	);
	LUT4 #(
		.INIT('h6f06)
	) name1395 (
		_w1363_,
		_w1365_,
		_w1414_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('h1680)
	) name1396 (
		_w1270_,
		_w1293_,
		_w1363_,
		_w1367_,
		_w1422_
	);
	LUT4 #(
		.INIT('h629d)
	) name1397 (
		_w1294_,
		_w1363_,
		_w1364_,
		_w1367_,
		_w1423_
	);
	LUT3 #(
		.INIT('h54)
	) name1398 (
		_w1413_,
		_w1421_,
		_w1422_,
		_w1424_
	);
	LUT4 #(
		.INIT('h1680)
	) name1399 (
		_w1252_,
		_w1268_,
		_w1366_,
		_w1369_,
		_w1425_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name1400 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1410_,
		_w1426_
	);
	LUT3 #(
		.INIT('h54)
	) name1401 (
		_w1412_,
		_w1424_,
		_w1425_,
		_w1427_
	);
	LUT3 #(
		.INIT('h06)
	) name1402 (
		_w1370_,
		_w1372_,
		_w1408_,
		_w1428_
	);
	LUT3 #(
		.INIT('h69)
	) name1403 (
		_w1370_,
		_w1372_,
		_w1408_,
		_w1429_
	);
	LUT4 #(
		.INIT('h629d)
	) name1404 (
		_w1231_,
		_w1370_,
		_w1371_,
		_w1374_,
		_w1430_
	);
	LUT4 #(
		.INIT('hba00)
	) name1405 (
		_w1409_,
		_w1427_,
		_w1429_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name1406 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1404_,
		_w1432_
	);
	LUT4 #(
		.INIT('h0155)
	) name1407 (
		_w1406_,
		_w1407_,
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT3 #(
		.INIT('h06)
	) name1408 (
		_w1377_,
		_w1379_,
		_w1402_,
		_w1434_
	);
	LUT3 #(
		.INIT('h69)
	) name1409 (
		_w1377_,
		_w1379_,
		_w1402_,
		_w1435_
	);
	LUT4 #(
		.INIT('h629d)
	) name1410 (
		_w1177_,
		_w1377_,
		_w1378_,
		_w1397_,
		_w1436_
	);
	LUT4 #(
		.INIT('hba00)
	) name1411 (
		_w1403_,
		_w1433_,
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h0400)
	) name1412 (
		_w144_,
		_w387_,
		_w517_,
		_w665_,
		_w1438_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1413 (
		_w87_,
		_w46_,
		_w125_,
		_w98_,
		_w1439_
	);
	LUT4 #(
		.INIT('h4000)
	) name1414 (
		_w407_,
		_w174_,
		_w621_,
		_w1439_,
		_w1440_
	);
	LUT4 #(
		.INIT('h8000)
	) name1415 (
		_w226_,
		_w445_,
		_w1438_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h1bff)
	) name1416 (
		_w46_,
		_w53_,
		_w95_,
		_w102_,
		_w1442_
	);
	LUT4 #(
		.INIT('h0100)
	) name1417 (
		_w209_,
		_w244_,
		_w203_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		_w231_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h8000)
	) name1419 (
		_w810_,
		_w1263_,
		_w1444_,
		_w1441_,
		_w1445_
	);
	LUT3 #(
		.INIT('h10)
	) name1420 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1446_
	);
	LUT4 #(
		.INIT('h9204)
	) name1421 (
		_w1391_,
		_w1395_,
		_w1380_,
		_w1445_,
		_w1447_
	);
	LUT4 #(
		.INIT('h1e2d)
	) name1422 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1399_,
		_w1448_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1423 (
		_w37_,
		_w1401_,
		_w1437_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h2)
	) name1424 (
		_w34_,
		_w36_,
		_w1450_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1425 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1450_,
		_w1451_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1426 (
		\a[3] ,
		\a[4] ,
		\a[22] ,
		_w27_,
		_w1452_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		_w34_,
		_w1452_,
		_w1453_
	);
	LUT3 #(
		.INIT('h04)
	) name1428 (
		_w34_,
		_w36_,
		_w1452_,
		_w1454_
	);
	LUT3 #(
		.INIT('h90)
	) name1429 (
		_w1377_,
		_w1379_,
		_w1454_,
		_w1455_
	);
	LUT3 #(
		.INIT('h07)
	) name1430 (
		_w1400_,
		_w1453_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		_w1451_,
		_w1456_,
		_w1457_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1432 (
		\a[10] ,
		\a[11] ,
		\a[22] ,
		_w41_,
		_w1458_
	);
	LUT3 #(
		.INIT('h69)
	) name1433 (
		\a[9] ,
		_w360_,
		_w581_,
		_w1459_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		_w1458_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h6996)
	) name1435 (
		_w1363_,
		_w1365_,
		_w1414_,
		_w1420_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w1458_,
		_w1459_,
		_w1462_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1437 (
		\a[9] ,
		\a[10] ,
		\a[22] ,
		_w40_,
		_w1463_
	);
	LUT3 #(
		.INIT('h02)
	) name1438 (
		_w1458_,
		_w1459_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h90)
	) name1439 (
		_w1357_,
		_w1359_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name1440 (
		_w1459_,
		_w1463_,
		_w1466_
	);
	LUT4 #(
		.INIT('h060f)
	) name1441 (
		_w1360_,
		_w1362_,
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1442 (
		_w1363_,
		_w1365_,
		_w1462_,
		_w1467_,
		_w1468_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1443 (
		_w366_,
		_w1460_,
		_w1461_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1444 (
		\a[11] ,
		\a[12] ,
		\a[22] ,
		_w42_,
		_w1470_
	);
	LUT4 #(
		.INIT('h4114)
	) name1445 (
		_w424_,
		_w1119_,
		_w1350_,
		_w1355_,
		_w1471_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('h90)
	) name1447 (
		_w1331_,
		_w1349_,
		_w1417_,
		_w1473_
	);
	LUT4 #(
		.INIT('h6966)
	) name1448 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1416_,
		_w1474_
	);
	LUT2 #(
		.INIT('h8)
	) name1449 (
		_w1392_,
		_w1470_,
		_w1475_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1450 (
		\a[12] ,
		\a[13] ,
		\a[22] ,
		_w43_,
		_w1476_
	);
	LUT2 #(
		.INIT('h4)
	) name1451 (
		_w1470_,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('h9600)
	) name1452 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w1392_,
		_w1470_,
		_w1479_
	);
	LUT4 #(
		.INIT('h6900)
	) name1454 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1479_,
		_w1480_
	);
	LUT4 #(
		.INIT('h000b)
	) name1455 (
		_w1474_,
		_w1475_,
		_w1478_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h9)
	) name1456 (
		_w1472_,
		_w1481_,
		_w1482_
	);
	LUT4 #(
		.INIT('h9600)
	) name1457 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1470_,
		_w1483_
	);
	LUT4 #(
		.INIT('h9600)
	) name1458 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1466_,
		_w1484_
	);
	LUT4 #(
		.INIT('h6900)
	) name1459 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1462_,
		_w1485_
	);
	LUT4 #(
		.INIT('h000d)
	) name1460 (
		_w1460_,
		_w1474_,
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h9600)
	) name1461 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1459_,
		_w1487_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w366_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		_w1486_,
		_w1488_,
		_w1489_
	);
	LUT4 #(
		.INIT('h6090)
	) name1464 (
		_w1357_,
		_w1359_,
		_w1460_,
		_w1473_,
		_w1490_
	);
	LUT3 #(
		.INIT('h90)
	) name1465 (
		_w1357_,
		_w1359_,
		_w1462_,
		_w1491_
	);
	LUT4 #(
		.INIT('h9600)
	) name1466 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1464_,
		_w1492_
	);
	LUT4 #(
		.INIT('h6900)
	) name1467 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1466_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('h10)
	) name1469 (
		_w1491_,
		_w1490_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h80)
	) name1470 (
		_w1483_,
		_w1489_,
		_w1495_,
		_w1496_
	);
	LUT4 #(
		.INIT('h9669)
	) name1471 (
		_w1360_,
		_w1362_,
		_w1415_,
		_w1419_,
		_w1497_
	);
	LUT4 #(
		.INIT('h6900)
	) name1472 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1464_,
		_w1498_
	);
	LUT4 #(
		.INIT('h006f)
	) name1473 (
		_w1357_,
		_w1359_,
		_w1466_,
		_w1498_,
		_w1499_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1474 (
		_w1360_,
		_w1362_,
		_w1462_,
		_w1499_,
		_w1500_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1475 (
		_w366_,
		_w1460_,
		_w1497_,
		_w1500_,
		_w1501_
	);
	LUT3 #(
		.INIT('h15)
	) name1476 (
		_w1483_,
		_w1489_,
		_w1495_,
		_w1502_
	);
	LUT3 #(
		.INIT('h6a)
	) name1477 (
		_w1483_,
		_w1489_,
		_w1495_,
		_w1503_
	);
	LUT3 #(
		.INIT('h51)
	) name1478 (
		_w1496_,
		_w1501_,
		_w1502_,
		_w1504_
	);
	LUT3 #(
		.INIT('h71)
	) name1479 (
		_w1469_,
		_w1482_,
		_w1504_,
		_w1505_
	);
	LUT3 #(
		.INIT('h90)
	) name1480 (
		_w1421_,
		_w1423_,
		_w1460_,
		_w1506_
	);
	LUT3 #(
		.INIT('h90)
	) name1481 (
		_w1360_,
		_w1362_,
		_w1464_,
		_w1507_
	);
	LUT4 #(
		.INIT('h006f)
	) name1482 (
		_w1363_,
		_w1365_,
		_w1466_,
		_w1507_,
		_w1508_
	);
	LUT3 #(
		.INIT('h70)
	) name1483 (
		_w1411_,
		_w1462_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name1484 (
		_w1481_,
		_w1483_,
		_w1510_
	);
	LUT3 #(
		.INIT('h51)
	) name1485 (
		_w424_,
		_w1481_,
		_w1483_,
		_w1511_
	);
	LUT4 #(
		.INIT('h6900)
	) name1486 (
		_w1357_,
		_w1359_,
		_w1473_,
		_w1475_,
		_w1512_
	);
	LUT3 #(
		.INIT('h90)
	) name1487 (
		_w1357_,
		_w1359_,
		_w1479_,
		_w1513_
	);
	LUT3 #(
		.INIT('h02)
	) name1488 (
		_w1392_,
		_w1470_,
		_w1476_,
		_w1514_
	);
	LUT4 #(
		.INIT('h9600)
	) name1489 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1514_,
		_w1515_
	);
	LUT4 #(
		.INIT('h6900)
	) name1490 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1477_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name1491 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT3 #(
		.INIT('h10)
	) name1492 (
		_w1513_,
		_w1512_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h9)
	) name1493 (
		_w1511_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1494 (
		_w366_,
		_w1506_,
		_w1509_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0065)
	) name1495 (
		_w366_,
		_w1506_,
		_w1509_,
		_w1519_,
		_w1521_
	);
	LUT4 #(
		.INIT('h659a)
	) name1496 (
		_w366_,
		_w1506_,
		_w1509_,
		_w1519_,
		_w1522_
	);
	LUT2 #(
		.INIT('h9)
	) name1497 (
		_w1505_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1498 (
		\a[5] ,
		\a[6] ,
		\a[22] ,
		_w29_,
		_w1524_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1499 (
		\a[7] ,
		\a[8] ,
		\a[22] ,
		_w39_,
		_w1525_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1501 (
		_w1409_,
		_w1427_,
		_w1428_,
		_w1430_,
		_w1527_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		_w1524_,
		_w1525_,
		_w1528_
	);
	LUT4 #(
		.INIT('h6c66)
	) name1503 (
		\a[6] ,
		\a[7] ,
		\a[22] ,
		_w38_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w1524_,
		_w1529_,
		_w1530_
	);
	LUT3 #(
		.INIT('h04)
	) name1505 (
		_w1524_,
		_w1525_,
		_w1529_,
		_w1531_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1506 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1531_,
		_w1532_
	);
	LUT4 #(
		.INIT('h006f)
	) name1507 (
		_w1370_,
		_w1372_,
		_w1530_,
		_w1532_,
		_w1533_
	);
	LUT3 #(
		.INIT('h70)
	) name1508 (
		_w1405_,
		_w1528_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1509 (
		_w581_,
		_w1526_,
		_w1527_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		_w1523_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w1523_,
		_w1535_,
		_w1537_
	);
	LUT2 #(
		.INIT('h6)
	) name1512 (
		_w1523_,
		_w1535_,
		_w1538_
	);
	LUT3 #(
		.INIT('h90)
	) name1513 (
		_w1427_,
		_w1429_,
		_w1526_,
		_w1539_
	);
	LUT3 #(
		.INIT('h90)
	) name1514 (
		_w1370_,
		_w1372_,
		_w1528_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name1515 (
		_w1411_,
		_w1531_,
		_w1541_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1516 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1530_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		_w1540_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h69)
	) name1519 (
		_w1469_,
		_w1482_,
		_w1504_,
		_w1545_
	);
	LUT4 #(
		.INIT('h0065)
	) name1520 (
		_w581_,
		_w1539_,
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1521 (
		_w581_,
		_w1539_,
		_w1544_,
		_w1545_,
		_w1547_
	);
	LUT3 #(
		.INIT('h90)
	) name1522 (
		_w1424_,
		_w1426_,
		_w1526_,
		_w1548_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1523 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1528_,
		_w1549_
	);
	LUT3 #(
		.INIT('h90)
	) name1524 (
		_w1363_,
		_w1365_,
		_w1531_,
		_w1550_
	);
	LUT3 #(
		.INIT('h07)
	) name1525 (
		_w1411_,
		_w1530_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		_w1549_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h6)
	) name1527 (
		_w1501_,
		_w1503_,
		_w1553_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1528 (
		_w581_,
		_w1548_,
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h0065)
	) name1529 (
		_w581_,
		_w1548_,
		_w1552_,
		_w1553_,
		_w1555_
	);
	LUT4 #(
		.INIT('h659a)
	) name1530 (
		_w581_,
		_w1548_,
		_w1552_,
		_w1553_,
		_w1556_
	);
	LUT3 #(
		.INIT('h90)
	) name1531 (
		_w1421_,
		_w1423_,
		_w1526_,
		_w1557_
	);
	LUT3 #(
		.INIT('h90)
	) name1532 (
		_w1360_,
		_w1362_,
		_w1531_,
		_w1558_
	);
	LUT4 #(
		.INIT('h006f)
	) name1533 (
		_w1363_,
		_w1365_,
		_w1530_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h70)
	) name1534 (
		_w1411_,
		_w1528_,
		_w1559_,
		_w1560_
	);
	LUT3 #(
		.INIT('h45)
	) name1535 (
		_w366_,
		_w1487_,
		_w1486_,
		_w1561_
	);
	LUT2 #(
		.INIT('h9)
	) name1536 (
		_w1495_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('h0065)
	) name1537 (
		_w581_,
		_w1557_,
		_w1560_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1538 (
		_w581_,
		_w1557_,
		_w1560_,
		_w1562_,
		_w1564_
	);
	LUT3 #(
		.INIT('h90)
	) name1539 (
		_w1357_,
		_w1359_,
		_w1531_,
		_w1565_
	);
	LUT4 #(
		.INIT('h006f)
	) name1540 (
		_w1360_,
		_w1362_,
		_w1530_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1541 (
		_w1363_,
		_w1365_,
		_w1528_,
		_w1566_,
		_w1567_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1542 (
		_w581_,
		_w1461_,
		_w1526_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name1543 (
		_w366_,
		_w1487_,
		_w1569_
	);
	LUT2 #(
		.INIT('h9)
	) name1544 (
		_w1486_,
		_w1569_,
		_w1570_
	);
	LUT4 #(
		.INIT('h9600)
	) name1545 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1530_,
		_w1571_
	);
	LUT4 #(
		.INIT('h6900)
	) name1546 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1528_,
		_w1572_
	);
	LUT4 #(
		.INIT('h000b)
	) name1547 (
		_w1474_,
		_w1526_,
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('h9600)
	) name1548 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1524_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		_w581_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h8)
	) name1550 (
		_w1573_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h6900)
	) name1551 (
		_w1357_,
		_w1359_,
		_w1473_,
		_w1526_,
		_w1577_
	);
	LUT3 #(
		.INIT('h90)
	) name1552 (
		_w1357_,
		_w1359_,
		_w1528_,
		_w1578_
	);
	LUT4 #(
		.INIT('h9600)
	) name1553 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1531_,
		_w1579_
	);
	LUT4 #(
		.INIT('h6900)
	) name1554 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1530_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h10)
	) name1556 (
		_w1578_,
		_w1577_,
		_w1581_,
		_w1582_
	);
	LUT3 #(
		.INIT('h80)
	) name1557 (
		_w1487_,
		_w1576_,
		_w1582_,
		_w1583_
	);
	LUT4 #(
		.INIT('h6900)
	) name1558 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1531_,
		_w1584_
	);
	LUT4 #(
		.INIT('h006f)
	) name1559 (
		_w1357_,
		_w1359_,
		_w1530_,
		_w1584_,
		_w1585_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1560 (
		_w1360_,
		_w1362_,
		_w1528_,
		_w1585_,
		_w1586_
	);
	LUT4 #(
		.INIT('h6a55)
	) name1561 (
		_w581_,
		_w1497_,
		_w1526_,
		_w1586_,
		_w1587_
	);
	LUT3 #(
		.INIT('h15)
	) name1562 (
		_w1487_,
		_w1576_,
		_w1582_,
		_w1588_
	);
	LUT3 #(
		.INIT('h6a)
	) name1563 (
		_w1487_,
		_w1576_,
		_w1582_,
		_w1589_
	);
	LUT3 #(
		.INIT('h54)
	) name1564 (
		_w1583_,
		_w1587_,
		_w1588_,
		_w1590_
	);
	LUT3 #(
		.INIT('h71)
	) name1565 (
		_w1568_,
		_w1570_,
		_w1590_,
		_w1591_
	);
	LUT3 #(
		.INIT('h45)
	) name1566 (
		_w1563_,
		_w1564_,
		_w1591_,
		_w1592_
	);
	LUT3 #(
		.INIT('h45)
	) name1567 (
		_w1554_,
		_w1555_,
		_w1592_,
		_w1593_
	);
	LUT3 #(
		.INIT('h45)
	) name1568 (
		_w1546_,
		_w1547_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h32)
	) name1569 (
		_w1505_,
		_w1520_,
		_w1521_,
		_w1595_
	);
	LUT3 #(
		.INIT('h90)
	) name1570 (
		_w1424_,
		_w1426_,
		_w1460_,
		_w1596_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1571 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1462_,
		_w1597_
	);
	LUT3 #(
		.INIT('h90)
	) name1572 (
		_w1363_,
		_w1365_,
		_w1464_,
		_w1598_
	);
	LUT3 #(
		.INIT('h07)
	) name1573 (
		_w1411_,
		_w1466_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h4)
	) name1574 (
		_w1597_,
		_w1599_,
		_w1600_
	);
	LUT3 #(
		.INIT('h80)
	) name1575 (
		_w1471_,
		_w1510_,
		_w1518_,
		_w1601_
	);
	LUT4 #(
		.INIT('h1444)
	) name1576 (
		_w424_,
		_w1417_,
		_w1510_,
		_w1518_,
		_w1602_
	);
	LUT4 #(
		.INIT('h6900)
	) name1577 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1514_,
		_w1603_
	);
	LUT4 #(
		.INIT('h006f)
	) name1578 (
		_w1357_,
		_w1359_,
		_w1477_,
		_w1603_,
		_w1604_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1579 (
		_w1360_,
		_w1362_,
		_w1479_,
		_w1604_,
		_w1605_
	);
	LUT3 #(
		.INIT('h70)
	) name1580 (
		_w1475_,
		_w1497_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h9)
	) name1581 (
		_w1602_,
		_w1606_,
		_w1607_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1582 (
		_w366_,
		_w1596_,
		_w1600_,
		_w1607_,
		_w1608_
	);
	LUT4 #(
		.INIT('h0065)
	) name1583 (
		_w366_,
		_w1596_,
		_w1600_,
		_w1607_,
		_w1609_
	);
	LUT4 #(
		.INIT('h659a)
	) name1584 (
		_w366_,
		_w1596_,
		_w1600_,
		_w1607_,
		_w1610_
	);
	LUT2 #(
		.INIT('h9)
	) name1585 (
		_w1595_,
		_w1610_,
		_w1611_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1586 (
		_w1407_,
		_w1431_,
		_w1432_,
		_w1526_,
		_w1612_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1587 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1528_,
		_w1613_
	);
	LUT3 #(
		.INIT('h90)
	) name1588 (
		_w1370_,
		_w1372_,
		_w1531_,
		_w1614_
	);
	LUT3 #(
		.INIT('h07)
	) name1589 (
		_w1405_,
		_w1530_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name1590 (
		_w1613_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('h8488)
	) name1591 (
		_w581_,
		_w1611_,
		_w1612_,
		_w1616_,
		_w1617_
	);
	LUT4 #(
		.INIT('h6966)
	) name1592 (
		_w581_,
		_w1611_,
		_w1612_,
		_w1616_,
		_w1618_
	);
	LUT4 #(
		.INIT('he800)
	) name1593 (
		_w1523_,
		_w1535_,
		_w1594_,
		_w1618_,
		_w1619_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1594 (
		_w1536_,
		_w1537_,
		_w1594_,
		_w1618_,
		_w1620_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1595 (
		_w30_,
		_w1449_,
		_w1457_,
		_w1620_,
		_w1621_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1596 (
		_w1403_,
		_w1433_,
		_w1434_,
		_w1436_,
		_w1622_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1597 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1454_,
		_w1623_
	);
	LUT4 #(
		.INIT('h006f)
	) name1598 (
		_w1377_,
		_w1379_,
		_w1453_,
		_w1623_,
		_w1624_
	);
	LUT3 #(
		.INIT('h70)
	) name1599 (
		_w1450_,
		_w1400_,
		_w1624_,
		_w1625_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1600 (
		_w30_,
		_w37_,
		_w1622_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h6)
	) name1601 (
		_w1538_,
		_w1594_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h82)
	) name1603 (
		_w37_,
		_w1433_,
		_w1435_,
		_w1629_
	);
	LUT3 #(
		.INIT('h90)
	) name1604 (
		_w1377_,
		_w1379_,
		_w1450_,
		_w1630_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1605 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1453_,
		_w1631_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		_w1454_,
		_w1405_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h4)
	) name1608 (
		_w1630_,
		_w1633_,
		_w1634_
	);
	LUT4 #(
		.INIT('h659a)
	) name1609 (
		_w581_,
		_w1539_,
		_w1544_,
		_w1545_,
		_w1635_
	);
	LUT2 #(
		.INIT('h6)
	) name1610 (
		_w1593_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h009a)
	) name1611 (
		_w30_,
		_w1629_,
		_w1634_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1612 (
		_w37_,
		_w1407_,
		_w1431_,
		_w1432_,
		_w1638_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1613 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1450_,
		_w1639_
	);
	LUT3 #(
		.INIT('h90)
	) name1614 (
		_w1370_,
		_w1372_,
		_w1454_,
		_w1640_
	);
	LUT3 #(
		.INIT('h07)
	) name1615 (
		_w1453_,
		_w1405_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w1639_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h6)
	) name1617 (
		_w1556_,
		_w1592_,
		_w1643_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1618 (
		_w30_,
		_w1638_,
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1619 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1454_,
		_w1645_
	);
	LUT4 #(
		.INIT('h006f)
	) name1620 (
		_w1370_,
		_w1372_,
		_w1453_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h70)
	) name1621 (
		_w1450_,
		_w1405_,
		_w1646_,
		_w1647_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1622 (
		_w30_,
		_w37_,
		_w1527_,
		_w1647_,
		_w1648_
	);
	LUT4 #(
		.INIT('h659a)
	) name1623 (
		_w581_,
		_w1557_,
		_w1560_,
		_w1562_,
		_w1649_
	);
	LUT2 #(
		.INIT('h6)
	) name1624 (
		_w1591_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		_w1648_,
		_w1650_,
		_w1651_
	);
	LUT3 #(
		.INIT('h82)
	) name1626 (
		_w37_,
		_w1427_,
		_w1429_,
		_w1652_
	);
	LUT3 #(
		.INIT('h90)
	) name1627 (
		_w1370_,
		_w1372_,
		_w1450_,
		_w1653_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w1454_,
		_w1411_,
		_w1654_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1629 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1453_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h4)
	) name1631 (
		_w1653_,
		_w1656_,
		_w1657_
	);
	LUT3 #(
		.INIT('h69)
	) name1632 (
		_w1568_,
		_w1570_,
		_w1590_,
		_w1658_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1633 (
		_w30_,
		_w1652_,
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT3 #(
		.INIT('h82)
	) name1634 (
		_w37_,
		_w1424_,
		_w1426_,
		_w1660_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1635 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1450_,
		_w1661_
	);
	LUT3 #(
		.INIT('h90)
	) name1636 (
		_w1363_,
		_w1365_,
		_w1454_,
		_w1662_
	);
	LUT3 #(
		.INIT('h07)
	) name1637 (
		_w1453_,
		_w1411_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h4)
	) name1638 (
		_w1661_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h9)
	) name1639 (
		_w1587_,
		_w1589_,
		_w1665_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1640 (
		_w30_,
		_w1660_,
		_w1664_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('h82)
	) name1641 (
		_w37_,
		_w1421_,
		_w1423_,
		_w1667_
	);
	LUT3 #(
		.INIT('h90)
	) name1642 (
		_w1360_,
		_w1362_,
		_w1454_,
		_w1668_
	);
	LUT4 #(
		.INIT('h006f)
	) name1643 (
		_w1363_,
		_w1365_,
		_w1453_,
		_w1668_,
		_w1669_
	);
	LUT3 #(
		.INIT('h70)
	) name1644 (
		_w1450_,
		_w1411_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('h45)
	) name1645 (
		_w581_,
		_w1574_,
		_w1573_,
		_w1671_
	);
	LUT2 #(
		.INIT('h9)
	) name1646 (
		_w1582_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1647 (
		_w30_,
		_w1667_,
		_w1670_,
		_w1672_,
		_w1673_
	);
	LUT3 #(
		.INIT('h90)
	) name1648 (
		_w1357_,
		_w1359_,
		_w1454_,
		_w1674_
	);
	LUT4 #(
		.INIT('h006f)
	) name1649 (
		_w1360_,
		_w1362_,
		_w1453_,
		_w1674_,
		_w1675_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1650 (
		_w1363_,
		_w1365_,
		_w1450_,
		_w1675_,
		_w1676_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1651 (
		_w30_,
		_w37_,
		_w1461_,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h4)
	) name1652 (
		_w581_,
		_w1574_,
		_w1678_
	);
	LUT2 #(
		.INIT('h9)
	) name1653 (
		_w1573_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h9600)
	) name1654 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1453_,
		_w1680_
	);
	LUT4 #(
		.INIT('h6900)
	) name1655 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1450_,
		_w1681_
	);
	LUT4 #(
		.INIT('h000d)
	) name1656 (
		_w37_,
		_w1474_,
		_w1680_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h9600)
	) name1657 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w34_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w30_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		_w1682_,
		_w1684_,
		_w1685_
	);
	LUT4 #(
		.INIT('h6090)
	) name1660 (
		_w1357_,
		_w1359_,
		_w37_,
		_w1473_,
		_w1686_
	);
	LUT3 #(
		.INIT('h90)
	) name1661 (
		_w1357_,
		_w1359_,
		_w1450_,
		_w1687_
	);
	LUT4 #(
		.INIT('h9600)
	) name1662 (
		_w1119_,
		_w1350_,
		_w1355_,
		_w1454_,
		_w1688_
	);
	LUT4 #(
		.INIT('h6900)
	) name1663 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1453_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w1688_,
		_w1689_,
		_w1690_
	);
	LUT3 #(
		.INIT('h10)
	) name1665 (
		_w1687_,
		_w1686_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h80)
	) name1666 (
		_w1574_,
		_w1685_,
		_w1691_,
		_w1692_
	);
	LUT4 #(
		.INIT('h6900)
	) name1667 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1454_,
		_w1693_
	);
	LUT4 #(
		.INIT('h006f)
	) name1668 (
		_w1357_,
		_w1359_,
		_w1453_,
		_w1693_,
		_w1694_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1669 (
		_w1360_,
		_w1362_,
		_w1450_,
		_w1694_,
		_w1695_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1670 (
		_w30_,
		_w37_,
		_w1497_,
		_w1695_,
		_w1696_
	);
	LUT3 #(
		.INIT('h15)
	) name1671 (
		_w1574_,
		_w1685_,
		_w1691_,
		_w1697_
	);
	LUT3 #(
		.INIT('h6a)
	) name1672 (
		_w1574_,
		_w1685_,
		_w1691_,
		_w1698_
	);
	LUT3 #(
		.INIT('h51)
	) name1673 (
		_w1692_,
		_w1696_,
		_w1697_,
		_w1699_
	);
	LUT3 #(
		.INIT('h71)
	) name1674 (
		_w1677_,
		_w1679_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h0065)
	) name1675 (
		_w30_,
		_w1667_,
		_w1670_,
		_w1672_,
		_w1701_
	);
	LUT4 #(
		.INIT('h659a)
	) name1676 (
		_w30_,
		_w1667_,
		_w1670_,
		_w1672_,
		_w1702_
	);
	LUT3 #(
		.INIT('h54)
	) name1677 (
		_w1673_,
		_w1700_,
		_w1701_,
		_w1703_
	);
	LUT4 #(
		.INIT('h0065)
	) name1678 (
		_w30_,
		_w1660_,
		_w1664_,
		_w1665_,
		_w1704_
	);
	LUT4 #(
		.INIT('h659a)
	) name1679 (
		_w30_,
		_w1660_,
		_w1664_,
		_w1665_,
		_w1705_
	);
	LUT3 #(
		.INIT('h54)
	) name1680 (
		_w1666_,
		_w1703_,
		_w1704_,
		_w1706_
	);
	LUT4 #(
		.INIT('h0065)
	) name1681 (
		_w30_,
		_w1652_,
		_w1657_,
		_w1658_,
		_w1707_
	);
	LUT4 #(
		.INIT('h659a)
	) name1682 (
		_w30_,
		_w1652_,
		_w1657_,
		_w1658_,
		_w1708_
	);
	LUT3 #(
		.INIT('h54)
	) name1683 (
		_w1659_,
		_w1706_,
		_w1707_,
		_w1709_
	);
	LUT2 #(
		.INIT('h4)
	) name1684 (
		_w1648_,
		_w1650_,
		_w1710_
	);
	LUT2 #(
		.INIT('h9)
	) name1685 (
		_w1648_,
		_w1650_,
		_w1711_
	);
	LUT4 #(
		.INIT('h659a)
	) name1686 (
		_w30_,
		_w1638_,
		_w1642_,
		_w1643_,
		_w1712_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1687 (
		_w1648_,
		_w1650_,
		_w1709_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h9a65)
	) name1688 (
		_w30_,
		_w1629_,
		_w1634_,
		_w1636_,
		_w1714_
	);
	LUT4 #(
		.INIT('h0155)
	) name1689 (
		_w1637_,
		_w1644_,
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		_w1626_,
		_w1627_,
		_w1716_
	);
	LUT2 #(
		.INIT('h6)
	) name1691 (
		_w1626_,
		_w1627_,
		_w1717_
	);
	LUT4 #(
		.INIT('h659a)
	) name1692 (
		_w30_,
		_w1449_,
		_w1457_,
		_w1620_,
		_w1718_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1693 (
		_w1626_,
		_w1627_,
		_w1715_,
		_w1718_,
		_w1719_
	);
	LUT4 #(
		.INIT('h010f)
	) name1694 (
		_w1401_,
		_w1437_,
		_w1447_,
		_w1448_,
		_w1720_
	);
	LUT3 #(
		.INIT('h01)
	) name1695 (
		_w252_,
		_w242_,
		_w181_,
		_w1721_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name1696 (
		_w46_,
		_w53_,
		_w134_,
		_w116_,
		_w1722_
	);
	LUT4 #(
		.INIT('h1bff)
	) name1697 (
		_w46_,
		_w134_,
		_w102_,
		_w70_,
		_w1723_
	);
	LUT4 #(
		.INIT('h8000)
	) name1698 (
		_w319_,
		_w659_,
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT4 #(
		.INIT('h777f)
	) name1699 (
		_w46_,
		_w53_,
		_w113_,
		_w100_,
		_w1725_
	);
	LUT4 #(
		.INIT('h4f7f)
	) name1700 (
		_w206_,
		_w46_,
		_w95_,
		_w79_,
		_w1726_
	);
	LUT3 #(
		.INIT('h40)
	) name1701 (
		_w517_,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h153f)
	) name1702 (
		_w88_,
		_w82_,
		_w77_,
		_w116_,
		_w1728_
	);
	LUT4 #(
		.INIT('h135f)
	) name1703 (
		_w206_,
		_w121_,
		_w77_,
		_w68_,
		_w1729_
	);
	LUT4 #(
		.INIT('h1000)
	) name1704 (
		_w176_,
		_w393_,
		_w1729_,
		_w1728_,
		_w1730_
	);
	LUT4 #(
		.INIT('h8000)
	) name1705 (
		_w1727_,
		_w1721_,
		_w1730_,
		_w1724_,
		_w1731_
	);
	LUT3 #(
		.INIT('h01)
	) name1706 (
		_w348_,
		_w340_,
		_w236_,
		_w1732_
	);
	LUT4 #(
		.INIT('h777f)
	) name1707 (
		_w46_,
		_w95_,
		_w102_,
		_w98_,
		_w1733_
	);
	LUT4 #(
		.INIT('h153f)
	) name1708 (
		_w121_,
		_w76_,
		_w85_,
		_w72_,
		_w1734_
	);
	LUT4 #(
		.INIT('h4000)
	) name1709 (
		_w73_,
		_w1279_,
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('h0400)
	) name1710 (
		_w168_,
		_w172_,
		_w86_,
		_w1342_,
		_w1736_
	);
	LUT4 #(
		.INIT('h8000)
	) name1711 (
		_w288_,
		_w1732_,
		_w1736_,
		_w1735_,
		_w1737_
	);
	LUT3 #(
		.INIT('h80)
	) name1712 (
		_w282_,
		_w1731_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h1000)
	) name1713 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1739_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1714 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1740_
	);
	LUT4 #(
		.INIT('hef10)
	) name1715 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1741_
	);
	LUT4 #(
		.INIT('h100e)
	) name1716 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1742_
	);
	LUT4 #(
		.INIT('he100)
	) name1717 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1743_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name1718 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1738_,
		_w1744_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w1400_,
		_w1454_,
		_w1745_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1720 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1453_,
		_w1746_
	);
	LUT4 #(
		.INIT('h000d)
	) name1721 (
		_w1450_,
		_w1741_,
		_w1745_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1722 (
		_w37_,
		_w1720_,
		_w1744_,
		_w1747_,
		_w1748_
	);
	LUT3 #(
		.INIT('h90)
	) name1723 (
		_w1433_,
		_w1435_,
		_w1526_,
		_w1749_
	);
	LUT3 #(
		.INIT('h90)
	) name1724 (
		_w1377_,
		_w1379_,
		_w1528_,
		_w1750_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1725 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1530_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		_w1405_,
		_w1531_,
		_w1752_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w1751_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h4)
	) name1728 (
		_w1750_,
		_w1753_,
		_w1754_
	);
	LUT3 #(
		.INIT('h32)
	) name1729 (
		_w1595_,
		_w1608_,
		_w1609_,
		_w1755_
	);
	LUT3 #(
		.INIT('h90)
	) name1730 (
		_w1427_,
		_w1429_,
		_w1460_,
		_w1756_
	);
	LUT3 #(
		.INIT('h90)
	) name1731 (
		_w1370_,
		_w1372_,
		_w1462_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		_w1411_,
		_w1464_,
		_w1758_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1733 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1466_,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h4)
	) name1735 (
		_w1757_,
		_w1760_,
		_w1761_
	);
	LUT4 #(
		.INIT('h4114)
	) name1736 (
		_w424_,
		_w1331_,
		_w1349_,
		_w1356_,
		_w1762_
	);
	LUT3 #(
		.INIT('h90)
	) name1737 (
		_w1357_,
		_w1359_,
		_w1514_,
		_w1763_
	);
	LUT4 #(
		.INIT('h006f)
	) name1738 (
		_w1360_,
		_w1362_,
		_w1477_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1739 (
		_w1363_,
		_w1365_,
		_w1479_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('h780f)
	) name1740 (
		_w1461_,
		_w1475_,
		_w1762_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('h5111)
	) name1741 (
		_w424_,
		_w1417_,
		_w1510_,
		_w1518_,
		_w1767_
	);
	LUT3 #(
		.INIT('h15)
	) name1742 (
		_w1601_,
		_w1606_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h9)
	) name1743 (
		_w1766_,
		_w1768_,
		_w1769_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1744 (
		_w366_,
		_w1756_,
		_w1761_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h0065)
	) name1745 (
		_w366_,
		_w1756_,
		_w1761_,
		_w1769_,
		_w1771_
	);
	LUT4 #(
		.INIT('h659a)
	) name1746 (
		_w366_,
		_w1756_,
		_w1761_,
		_w1769_,
		_w1772_
	);
	LUT2 #(
		.INIT('h9)
	) name1747 (
		_w1755_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1748 (
		_w581_,
		_w1749_,
		_w1754_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h659a)
	) name1749 (
		_w581_,
		_w1749_,
		_w1754_,
		_w1773_,
		_w1775_
	);
	LUT3 #(
		.INIT('h1e)
	) name1750 (
		_w1617_,
		_w1619_,
		_w1775_,
		_w1776_
	);
	LUT3 #(
		.INIT('h60)
	) name1751 (
		_w30_,
		_w1748_,
		_w1776_,
		_w1777_
	);
	LUT3 #(
		.INIT('h96)
	) name1752 (
		_w30_,
		_w1748_,
		_w1776_,
		_w1778_
	);
	LUT3 #(
		.INIT('h1e)
	) name1753 (
		_w1621_,
		_w1719_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('h2828)
	) name1754 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[22] ,
		_w1780_
	);
	LUT3 #(
		.INIT('h80)
	) name1755 (
		_w518_,
		_w1178_,
		_w1313_,
		_w1781_
	);
	LUT4 #(
		.INIT('h0777)
	) name1756 (
		_w88_,
		_w76_,
		_w79_,
		_w71_,
		_w1782_
	);
	LUT3 #(
		.INIT('h40)
	) name1757 (
		_w211_,
		_w241_,
		_w1782_,
		_w1783_
	);
	LUT4 #(
		.INIT('h8000)
	) name1758 (
		_w1198_,
		_w1254_,
		_w1781_,
		_w1783_,
		_w1784_
	);
	LUT3 #(
		.INIT('h80)
	) name1759 (
		_w338_,
		_w390_,
		_w1784_,
		_w1785_
	);
	LUT4 #(
		.INIT('h777f)
	) name1760 (
		_w46_,
		_w95_,
		_w125_,
		_w100_,
		_w1786_
	);
	LUT3 #(
		.INIT('h80)
	) name1761 (
		_w371_,
		_w341_,
		_w1786_,
		_w1787_
	);
	LUT3 #(
		.INIT('h80)
	) name1762 (
		_w350_,
		_w676_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w354_,
		_w378_,
		_w1789_
	);
	LUT4 #(
		.INIT('h8000)
	) name1764 (
		_w326_,
		_w327_,
		_w385_,
		_w389_,
		_w1790_
	);
	LUT4 #(
		.INIT('h8000)
	) name1765 (
		_w411_,
		_w1788_,
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT3 #(
		.INIT('h81)
	) name1766 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1792_
	);
	LUT3 #(
		.INIT('h21)
	) name1767 (
		_w1739_,
		_w1741_,
		_w1785_,
		_w1793_
	);
	LUT3 #(
		.INIT('h4b)
	) name1768 (
		_w1739_,
		_w1740_,
		_w1785_,
		_w1794_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1769 (
		_w1720_,
		_w1742_,
		_w1744_,
		_w1794_,
		_w1795_
	);
	LUT3 #(
		.INIT('h60)
	) name1770 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1796_
	);
	LUT3 #(
		.INIT('h1e)
	) name1771 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1797_
	);
	LUT4 #(
		.INIT('h5501)
	) name1772 (
		_w1792_,
		_w1793_,
		_w1795_,
		_w1796_,
		_w1798_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w411_,
		_w268_,
		_w1799_
	);
	LUT4 #(
		.INIT('h135f)
	) name1774 (
		_w95_,
		_w113_,
		_w62_,
		_w71_,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		_w332_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h8000)
	) name1776 (
		_w385_,
		_w389_,
		_w401_,
		_w403_,
		_w1802_
	);
	LUT4 #(
		.INIT('h8000)
	) name1777 (
		_w351_,
		_w1799_,
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT4 #(
		.INIT('h007f)
	) name1778 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('h8000)
	) name1779 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1805_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1780 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1806_
	);
	LUT4 #(
		.INIT('h8007)
	) name1781 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1807_
	);
	LUT4 #(
		.INIT('h7800)
	) name1782 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1808_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1783 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1803_,
		_w1809_
	);
	LUT4 #(
		.INIT('h8282)
	) name1784 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		\a[22] ,
		_w1810_
	);
	LUT3 #(
		.INIT('h10)
	) name1785 (
		\a[0] ,
		\a[1] ,
		\a[2] ,
		_w1811_
	);
	LUT3 #(
		.INIT('h90)
	) name1786 (
		_w1739_,
		_w1785_,
		_w1811_,
		_w1812_
	);
	LUT3 #(
		.INIT('h44)
	) name1787 (
		\a[0] ,
		\a[1] ,
		\a[22] ,
		_w1813_
	);
	LUT4 #(
		.INIT('h8700)
	) name1788 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1813_,
		_w1814_
	);
	LUT4 #(
		.INIT('h000b)
	) name1789 (
		_w1806_,
		_w1810_,
		_w1812_,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1790 (
		_w1780_,
		_w1798_,
		_w1809_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h6)
	) name1791 (
		_w33_,
		_w1816_,
		_w1817_
	);
	LUT3 #(
		.INIT('h48)
	) name1792 (
		_w33_,
		_w1779_,
		_w1816_,
		_w1818_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1793 (
		_w1628_,
		_w1715_,
		_w1716_,
		_w1718_,
		_w1819_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1794 (
		_w1780_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w1820_
	);
	LUT4 #(
		.INIT('h8700)
	) name1795 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1810_,
		_w1821_
	);
	LUT2 #(
		.INIT('h4)
	) name1796 (
		_w1741_,
		_w1811_,
		_w1822_
	);
	LUT3 #(
		.INIT('h90)
	) name1797 (
		_w1739_,
		_w1785_,
		_w1813_,
		_w1823_
	);
	LUT3 #(
		.INIT('h01)
	) name1798 (
		_w1821_,
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT4 #(
		.INIT('h8488)
	) name1799 (
		_w33_,
		_w1819_,
		_w1820_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h9)
	) name1800 (
		_w1715_,
		_w1717_,
		_w1826_
	);
	LUT4 #(
		.INIT('h32cd)
	) name1801 (
		_w1720_,
		_w1742_,
		_w1743_,
		_w1794_,
		_w1827_
	);
	LUT3 #(
		.INIT('h90)
	) name1802 (
		_w1739_,
		_w1785_,
		_w1810_,
		_w1828_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1803 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1811_,
		_w1829_
	);
	LUT3 #(
		.INIT('h0b)
	) name1804 (
		_w1741_,
		_w1813_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h4)
	) name1805 (
		_w1828_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1806 (
		_w33_,
		_w1780_,
		_w1827_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name1807 (
		_w1826_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h6)
	) name1808 (
		_w1826_,
		_w1832_,
		_w1834_
	);
	LUT3 #(
		.INIT('h1e)
	) name1809 (
		_w1644_,
		_w1713_,
		_w1714_,
		_w1835_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1810 (
		_w1651_,
		_w1709_,
		_w1710_,
		_w1712_,
		_w1836_
	);
	LUT3 #(
		.INIT('h90)
	) name1811 (
		_w1377_,
		_w1379_,
		_w1811_,
		_w1837_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1812 (
		_w1401_,
		_w1437_,
		_w1448_,
		_w1780_,
		_w1838_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1813 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1810_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		_w1400_,
		_w1813_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT4 #(
		.INIT('ha1aa)
	) name1816 (
		_w33_,
		_w1837_,
		_w1838_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w1836_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w1836_,
		_w1842_,
		_w1844_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1819 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1811_,
		_w1845_
	);
	LUT4 #(
		.INIT('h006f)
	) name1820 (
		_w1377_,
		_w1379_,
		_w1813_,
		_w1845_,
		_w1846_
	);
	LUT3 #(
		.INIT('h70)
	) name1821 (
		_w1400_,
		_w1810_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h6a55)
	) name1822 (
		_w33_,
		_w1622_,
		_w1780_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h9)
	) name1823 (
		_w1709_,
		_w1711_,
		_w1849_
	);
	LUT2 #(
		.INIT('h2)
	) name1824 (
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h9)
	) name1825 (
		_w1706_,
		_w1708_,
		_w1851_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1826 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1813_,
		_w1852_
	);
	LUT4 #(
		.INIT('h006f)
	) name1827 (
		_w1377_,
		_w1379_,
		_w1810_,
		_w1852_,
		_w1853_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1828 (
		_w1433_,
		_w1435_,
		_w1780_,
		_w1853_,
		_w1854_
	);
	LUT3 #(
		.INIT('h15)
	) name1829 (
		_w33_,
		_w1405_,
		_w1811_,
		_w1855_
	);
	LUT4 #(
		.INIT('h0131)
	) name1830 (
		_w33_,
		_w1851_,
		_w1854_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h9)
	) name1831 (
		_w1703_,
		_w1705_,
		_w1857_
	);
	LUT2 #(
		.INIT('h9)
	) name1832 (
		_w1700_,
		_w1702_,
		_w1858_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1833 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1811_,
		_w1859_
	);
	LUT2 #(
		.INIT('h1)
	) name1834 (
		_w33_,
		_w1859_,
		_w1860_
	);
	LUT3 #(
		.INIT('h90)
	) name1835 (
		_w1370_,
		_w1372_,
		_w1813_,
		_w1861_
	);
	LUT3 #(
		.INIT('h07)
	) name1836 (
		_w1405_,
		_w1810_,
		_w1861_,
		_w1862_
	);
	LUT4 #(
		.INIT('h0700)
	) name1837 (
		_w1527_,
		_w1780_,
		_w1860_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('h4055)
	) name1838 (
		_w33_,
		_w1527_,
		_w1780_,
		_w1862_,
		_w1864_
	);
	LUT3 #(
		.INIT('h54)
	) name1839 (
		_w1858_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h6)
	) name1840 (
		_w1696_,
		_w1698_,
		_w1866_
	);
	LUT3 #(
		.INIT('h45)
	) name1841 (
		_w30_,
		_w1683_,
		_w1682_,
		_w1867_
	);
	LUT2 #(
		.INIT('h9)
	) name1842 (
		_w1691_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w30_,
		_w1683_,
		_w1869_
	);
	LUT2 #(
		.INIT('h9)
	) name1844 (
		_w1682_,
		_w1869_,
		_w1870_
	);
	LUT4 #(
		.INIT('h9f00)
	) name1845 (
		_w1357_,
		_w1359_,
		_w1474_,
		_w1780_,
		_w1871_
	);
	LUT4 #(
		.INIT('hf900)
	) name1846 (
		_w1357_,
		_w1359_,
		_w1418_,
		_w1810_,
		_w1872_
	);
	LUT4 #(
		.INIT('h6900)
	) name1847 (
		_w1331_,
		_w1349_,
		_w1356_,
		_w1813_,
		_w1873_
	);
	LUT4 #(
		.INIT('h4114)
	) name1848 (
		_w27_,
		_w1119_,
		_w1350_,
		_w1355_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w33_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name1850 (
		_w1873_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('h0200)
	) name1851 (
		_w1683_,
		_w1872_,
		_w1871_,
		_w1876_,
		_w1877_
	);
	LUT4 #(
		.INIT('h5455)
	) name1852 (
		_w1683_,
		_w1872_,
		_w1871_,
		_w1876_,
		_w1878_
	);
	LUT3 #(
		.INIT('h90)
	) name1853 (
		_w1357_,
		_w1359_,
		_w1813_,
		_w1879_
	);
	LUT4 #(
		.INIT('h006f)
	) name1854 (
		_w1360_,
		_w1362_,
		_w1810_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1855 (
		_w33_,
		_w1497_,
		_w1780_,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('h2882)
	) name1856 (
		_w26_,
		_w1331_,
		_w1349_,
		_w1356_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w33_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('h7000)
	) name1858 (
		_w1497_,
		_w1780_,
		_w1880_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('h4445)
	) name1859 (
		_w1877_,
		_w1878_,
		_w1881_,
		_w1884_,
		_w1885_
	);
	LUT3 #(
		.INIT('h90)
	) name1860 (
		_w1357_,
		_w1359_,
		_w1811_,
		_w1886_
	);
	LUT4 #(
		.INIT('h006f)
	) name1861 (
		_w1360_,
		_w1362_,
		_w1813_,
		_w1886_,
		_w1887_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1862 (
		_w1363_,
		_w1365_,
		_w1810_,
		_w1887_,
		_w1888_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1863 (
		_w33_,
		_w1461_,
		_w1780_,
		_w1888_,
		_w1889_
	);
	LUT3 #(
		.INIT('h4d)
	) name1864 (
		_w1870_,
		_w1885_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h90)
	) name1865 (
		_w1421_,
		_w1423_,
		_w1780_,
		_w1891_
	);
	LUT3 #(
		.INIT('h90)
	) name1866 (
		_w1360_,
		_w1362_,
		_w1811_,
		_w1892_
	);
	LUT4 #(
		.INIT('h006f)
	) name1867 (
		_w1363_,
		_w1365_,
		_w1813_,
		_w1892_,
		_w1893_
	);
	LUT3 #(
		.INIT('h70)
	) name1868 (
		_w1411_,
		_w1810_,
		_w1893_,
		_w1894_
	);
	LUT3 #(
		.INIT('h65)
	) name1869 (
		_w33_,
		_w1891_,
		_w1894_,
		_w1895_
	);
	LUT4 #(
		.INIT('h088a)
	) name1870 (
		_w1866_,
		_w1868_,
		_w1890_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h90)
	) name1871 (
		_w1424_,
		_w1426_,
		_w1780_,
		_w1897_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1872 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1810_,
		_w1898_
	);
	LUT3 #(
		.INIT('h90)
	) name1873 (
		_w1363_,
		_w1365_,
		_w1811_,
		_w1899_
	);
	LUT3 #(
		.INIT('h07)
	) name1874 (
		_w1411_,
		_w1813_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h4)
	) name1875 (
		_w1898_,
		_w1900_,
		_w1901_
	);
	LUT3 #(
		.INIT('h65)
	) name1876 (
		_w33_,
		_w1897_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1877 (
		_w1896_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('h5110)
	) name1878 (
		_w1866_,
		_w1868_,
		_w1890_,
		_w1895_,
		_w1904_
	);
	LUT3 #(
		.INIT('h69)
	) name1879 (
		_w1677_,
		_w1679_,
		_w1699_,
		_w1905_
	);
	LUT3 #(
		.INIT('h90)
	) name1880 (
		_w1427_,
		_w1429_,
		_w1780_,
		_w1906_
	);
	LUT3 #(
		.INIT('h90)
	) name1881 (
		_w1370_,
		_w1372_,
		_w1810_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		_w1411_,
		_w1811_,
		_w1908_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1883 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1813_,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h4)
	) name1885 (
		_w1907_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('h1211)
	) name1886 (
		_w33_,
		_w1905_,
		_w1906_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('h01)
	) name1887 (
		_w1904_,
		_w1912_,
		_w1903_,
		_w1913_
	);
	LUT4 #(
		.INIT('h8488)
	) name1888 (
		_w33_,
		_w1905_,
		_w1906_,
		_w1911_,
		_w1914_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1889 (
		_w1858_,
		_w1863_,
		_w1864_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('h45)
	) name1890 (
		_w1865_,
		_w1913_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1891 (
		_w1407_,
		_w1431_,
		_w1432_,
		_w1780_,
		_w1917_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1892 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1810_,
		_w1918_
	);
	LUT3 #(
		.INIT('h90)
	) name1893 (
		_w1370_,
		_w1372_,
		_w1811_,
		_w1919_
	);
	LUT3 #(
		.INIT('h07)
	) name1894 (
		_w1405_,
		_w1813_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		_w1918_,
		_w1920_,
		_w1921_
	);
	LUT3 #(
		.INIT('h9a)
	) name1896 (
		_w33_,
		_w1917_,
		_w1921_,
		_w1922_
	);
	LUT4 #(
		.INIT('hc808)
	) name1897 (
		_w33_,
		_w1851_,
		_w1854_,
		_w1855_,
		_w1923_
	);
	LUT4 #(
		.INIT('h0107)
	) name1898 (
		_w1857_,
		_w1916_,
		_w1923_,
		_w1922_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w1848_,
		_w1849_,
		_w1925_
	);
	LUT4 #(
		.INIT('h5501)
	) name1900 (
		_w1850_,
		_w1856_,
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT3 #(
		.INIT('h54)
	) name1901 (
		_w1843_,
		_w1844_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		_w1400_,
		_w1811_,
		_w1928_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1903 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1813_,
		_w1929_
	);
	LUT4 #(
		.INIT('h000b)
	) name1904 (
		_w1741_,
		_w1810_,
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1905 (
		_w1720_,
		_w1744_,
		_w1780_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('h9)
	) name1906 (
		_w33_,
		_w1931_,
		_w1932_
	);
	LUT4 #(
		.INIT('h80a8)
	) name1907 (
		_w1834_,
		_w1835_,
		_w1927_,
		_w1932_,
		_w1933_
	);
	LUT4 #(
		.INIT('h6966)
	) name1908 (
		_w33_,
		_w1819_,
		_w1820_,
		_w1824_,
		_w1934_
	);
	LUT4 #(
		.INIT('h0155)
	) name1909 (
		_w1825_,
		_w1833_,
		_w1933_,
		_w1934_,
		_w1935_
	);
	LUT3 #(
		.INIT('h21)
	) name1910 (
		_w33_,
		_w1779_,
		_w1816_,
		_w1936_
	);
	LUT3 #(
		.INIT('h96)
	) name1911 (
		_w33_,
		_w1779_,
		_w1816_,
		_w1937_
	);
	LUT3 #(
		.INIT('h57)
	) name1912 (
		_w85_,
		_w125_,
		_w98_,
		_w1938_
	);
	LUT4 #(
		.INIT('h47ff)
	) name1913 (
		_w87_,
		_w46_,
		_w53_,
		_w113_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT3 #(
		.INIT('h57)
	) name1915 (
		_w121_,
		_w134_,
		_w62_,
		_w1941_
	);
	LUT3 #(
		.INIT('h80)
	) name1916 (
		_w90_,
		_w1204_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		_w1940_,
		_w1942_,
		_w1943_
	);
	LUT3 #(
		.INIT('h57)
	) name1918 (
		_w121_,
		_w59_,
		_w125_,
		_w1944_
	);
	LUT4 #(
		.INIT('h8000)
	) name1919 (
		_w568_,
		_w1208_,
		_w1313_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('h135f)
	) name1920 (
		_w206_,
		_w121_,
		_w106_,
		_w98_,
		_w1946_
	);
	LUT2 #(
		.INIT('h4)
	) name1921 (
		_w393_,
		_w1946_,
		_w1947_
	);
	LUT4 #(
		.INIT('h8000)
	) name1922 (
		_w1386_,
		_w119_,
		_w1947_,
		_w1945_,
		_w1948_
	);
	LUT4 #(
		.INIT('h8000)
	) name1923 (
		_w668_,
		_w674_,
		_w1943_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h6)
	) name1924 (
		_w1805_,
		_w1949_,
		_w1950_
	);
	LUT3 #(
		.INIT('h21)
	) name1925 (
		_w1805_,
		_w1806_,
		_w1949_,
		_w1951_
	);
	LUT3 #(
		.INIT('h2d)
	) name1926 (
		_w1804_,
		_w1805_,
		_w1949_,
		_w1952_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1927 (
		_w1798_,
		_w1807_,
		_w1809_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('h32cd)
	) name1928 (
		_w1798_,
		_w1807_,
		_w1808_,
		_w1952_,
		_w1954_
	);
	LUT3 #(
		.INIT('h84)
	) name1929 (
		_w1805_,
		_w1810_,
		_w1949_,
		_w1955_
	);
	LUT4 #(
		.INIT('h8700)
	) name1930 (
		_w1739_,
		_w1785_,
		_w1791_,
		_w1811_,
		_w1956_
	);
	LUT3 #(
		.INIT('h0b)
	) name1931 (
		_w1806_,
		_w1813_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w1955_,
		_w1957_,
		_w1958_
	);
	LUT4 #(
		.INIT('h6a55)
	) name1933 (
		_w33_,
		_w1780_,
		_w1954_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h010f)
	) name1934 (
		_w1621_,
		_w1719_,
		_w1777_,
		_w1778_,
		_w1960_
	);
	LUT4 #(
		.INIT('h010f)
	) name1935 (
		_w1617_,
		_w1619_,
		_w1774_,
		_w1775_,
		_w1961_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1936 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1531_,
		_w1962_
	);
	LUT4 #(
		.INIT('h006f)
	) name1937 (
		_w1377_,
		_w1379_,
		_w1530_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('h70)
	) name1938 (
		_w1400_,
		_w1528_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h6a55)
	) name1939 (
		_w581_,
		_w1526_,
		_w1622_,
		_w1964_,
		_w1965_
	);
	LUT3 #(
		.INIT('h32)
	) name1940 (
		_w1755_,
		_w1770_,
		_w1771_,
		_w1966_
	);
	LUT3 #(
		.INIT('h14)
	) name1941 (
		_w424_,
		_w1357_,
		_w1359_,
		_w1967_
	);
	LUT3 #(
		.INIT('h90)
	) name1942 (
		_w1421_,
		_w1423_,
		_w1475_,
		_w1968_
	);
	LUT3 #(
		.INIT('h90)
	) name1943 (
		_w1360_,
		_w1362_,
		_w1514_,
		_w1969_
	);
	LUT4 #(
		.INIT('h006f)
	) name1944 (
		_w1363_,
		_w1365_,
		_w1477_,
		_w1969_,
		_w1970_
	);
	LUT3 #(
		.INIT('h70)
	) name1945 (
		_w1411_,
		_w1479_,
		_w1970_,
		_w1971_
	);
	LUT3 #(
		.INIT('h65)
	) name1946 (
		_w1967_,
		_w1968_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h1441)
	) name1947 (
		_w424_,
		_w1331_,
		_w1349_,
		_w1356_,
		_w1973_
	);
	LUT4 #(
		.INIT('h7000)
	) name1948 (
		_w1461_,
		_w1475_,
		_w1765_,
		_w1973_,
		_w1974_
	);
	LUT3 #(
		.INIT('h0d)
	) name1949 (
		_w1766_,
		_w1768_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h9)
	) name1950 (
		_w1972_,
		_w1975_,
		_w1976_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1951 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1464_,
		_w1977_
	);
	LUT4 #(
		.INIT('h006f)
	) name1952 (
		_w1370_,
		_w1372_,
		_w1466_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('h70)
	) name1953 (
		_w1405_,
		_w1462_,
		_w1978_,
		_w1979_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1954 (
		_w366_,
		_w1460_,
		_w1527_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		_w1976_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w1976_,
		_w1980_,
		_w1982_
	);
	LUT2 #(
		.INIT('h6)
	) name1957 (
		_w1976_,
		_w1980_,
		_w1983_
	);
	LUT2 #(
		.INIT('h9)
	) name1958 (
		_w1966_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h4)
	) name1959 (
		_w1965_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		_w1965_,
		_w1984_,
		_w1986_
	);
	LUT2 #(
		.INIT('h9)
	) name1961 (
		_w1965_,
		_w1984_,
		_w1987_
	);
	LUT2 #(
		.INIT('h9)
	) name1962 (
		_w1961_,
		_w1987_,
		_w1988_
	);
	LUT3 #(
		.INIT('h82)
	) name1963 (
		_w1450_,
		_w1739_,
		_w1785_,
		_w1989_
	);
	LUT4 #(
		.INIT('h1e00)
	) name1964 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1454_,
		_w1990_
	);
	LUT3 #(
		.INIT('h0d)
	) name1965 (
		_w1453_,
		_w1741_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w1989_,
		_w1991_,
		_w1992_
	);
	LUT4 #(
		.INIT('h95aa)
	) name1967 (
		_w30_,
		_w37_,
		_w1827_,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		_w1988_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		_w1988_,
		_w1993_,
		_w1995_
	);
	LUT2 #(
		.INIT('h6)
	) name1970 (
		_w1988_,
		_w1993_,
		_w1996_
	);
	LUT2 #(
		.INIT('h9)
	) name1971 (
		_w1960_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h4)
	) name1972 (
		_w1959_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h9)
	) name1973 (
		_w1959_,
		_w1997_,
		_w1999_
	);
	LUT4 #(
		.INIT('h8e00)
	) name1974 (
		_w1779_,
		_w1817_,
		_w1935_,
		_w1999_,
		_w2000_
	);
	LUT4 #(
		.INIT('h54ab)
	) name1975 (
		_w1818_,
		_w1935_,
		_w1936_,
		_w1999_,
		_w2001_
	);
	LUT3 #(
		.INIT('h80)
	) name1976 (
		_w618_,
		_w807_,
		_w1732_,
		_w2002_
	);
	LUT4 #(
		.INIT('h0777)
	) name1977 (
		_w121_,
		_w76_,
		_w85_,
		_w79_,
		_w2003_
	);
	LUT4 #(
		.INIT('h4000)
	) name1978 (
		_w173_,
		_w254_,
		_w1941_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		_w452_,
		_w2004_,
		_w2005_
	);
	LUT3 #(
		.INIT('h80)
	) name1980 (
		_w214_,
		_w2002_,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w1239_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name1982 (
		_w2001_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w2001_,
		_w2007_,
		_w2009_
	);
	LUT2 #(
		.INIT('h9)
	) name1984 (
		_w2001_,
		_w2007_,
		_w2010_
	);
	LUT4 #(
		.INIT('h135f)
	) name1985 (
		_w113_,
		_w85_,
		_w71_,
		_w72_,
		_w2011_
	);
	LUT3 #(
		.INIT('h10)
	) name1986 (
		_w227_,
		_w146_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1987 (
		_w1305_,
		_w2012_,
		_w2013_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1988 (
		_w206_,
		_w46_,
		_w95_,
		_w98_,
		_w2014_
	);
	LUT3 #(
		.INIT('h10)
	) name1989 (
		_w347_,
		_w278_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1990 (
		_w114_,
		_w1192_,
		_w2016_
	);
	LUT3 #(
		.INIT('h10)
	) name1991 (
		_w69_,
		_w221_,
		_w1941_,
		_w2017_
	);
	LUT3 #(
		.INIT('h80)
	) name1992 (
		_w2015_,
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT4 #(
		.INIT('h0777)
	) name1993 (
		_w121_,
		_w59_,
		_w79_,
		_w71_,
		_w2019_
	);
	LUT3 #(
		.INIT('h57)
	) name1994 (
		_w76_,
		_w54_,
		_w96_,
		_w2020_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT3 #(
		.INIT('h80)
	) name1996 (
		_w2013_,
		_w2018_,
		_w2021_,
		_w2022_
	);
	LUT4 #(
		.INIT('h0777)
	) name1997 (
		_w85_,
		_w102_,
		_w77_,
		_w72_,
		_w2023_
	);
	LUT3 #(
		.INIT('h10)
	) name1998 (
		_w209_,
		_w86_,
		_w2023_,
		_w2024_
	);
	LUT4 #(
		.INIT('h8000)
	) name1999 (
		_w155_,
		_w160_,
		_w1727_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('h0001)
	) name2000 (
		_w348_,
		_w340_,
		_w128_,
		_w236_,
		_w2026_
	);
	LUT4 #(
		.INIT('h153f)
	) name2001 (
		_w106_,
		_w77_,
		_w68_,
		_w116_,
		_w2027_
	);
	LUT2 #(
		.INIT('h4)
	) name2002 (
		_w145_,
		_w2027_,
		_w2028_
	);
	LUT3 #(
		.INIT('h10)
	) name2003 (
		_w238_,
		_w271_,
		_w1728_,
		_w2029_
	);
	LUT4 #(
		.INIT('h8000)
	) name2004 (
		_w1336_,
		_w2026_,
		_w2028_,
		_w2029_,
		_w2030_
	);
	LUT3 #(
		.INIT('h80)
	) name2005 (
		_w188_,
		_w2025_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		_w2022_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('h60)
	) name2007 (
		_w1935_,
		_w1937_,
		_w2032_,
		_w2033_
	);
	LUT3 #(
		.INIT('h09)
	) name2008 (
		_w1935_,
		_w1937_,
		_w2032_,
		_w2034_
	);
	LUT3 #(
		.INIT('h1e)
	) name2009 (
		_w1833_,
		_w1933_,
		_w1934_,
		_w2035_
	);
	LUT4 #(
		.INIT('h1501)
	) name2010 (
		_w1834_,
		_w1835_,
		_w1927_,
		_w1932_,
		_w2036_
	);
	LUT3 #(
		.INIT('h1f)
	) name2011 (
		_w121_,
		_w106_,
		_w72_,
		_w2037_
	);
	LUT3 #(
		.INIT('h80)
	) name2012 (
		_w341_,
		_w819_,
		_w2037_,
		_w2038_
	);
	LUT4 #(
		.INIT('h8000)
	) name2013 (
		_w1227_,
		_w1243_,
		_w1244_,
		_w2038_,
		_w2039_
	);
	LUT3 #(
		.INIT('h37)
	) name2014 (
		_w91_,
		_w96_,
		_w116_,
		_w2040_
	);
	LUT3 #(
		.INIT('h80)
	) name2015 (
		_w1387_,
		_w245_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('h10)
	) name2016 (
		_w132_,
		_w73_,
		_w370_,
		_w2042_
	);
	LUT3 #(
		.INIT('h10)
	) name2017 (
		_w69_,
		_w221_,
		_w1323_,
		_w2043_
	);
	LUT4 #(
		.INIT('h37bf)
	) name2018 (
		_w46_,
		_w95_,
		_w113_,
		_w134_,
		_w2044_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w153_,
		_w2044_,
		_w2045_
	);
	LUT3 #(
		.INIT('h10)
	) name2020 (
		_w386_,
		_w64_,
		_w450_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8000)
	) name2021 (
		_w2045_,
		_w2046_,
		_w2042_,
		_w2043_,
		_w2047_
	);
	LUT4 #(
		.INIT('h8000)
	) name2022 (
		_w1288_,
		_w2041_,
		_w2039_,
		_w2047_,
		_w2048_
	);
	LUT3 #(
		.INIT('h01)
	) name2023 (
		_w1933_,
		_w2048_,
		_w2036_,
		_w2049_
	);
	LUT4 #(
		.INIT('h153f)
	) name2024 (
		_w121_,
		_w85_,
		_w79_,
		_w100_,
		_w2050_
	);
	LUT3 #(
		.INIT('h80)
	) name2025 (
		_w212_,
		_w1256_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('h57df)
	) name2026 (
		_w87_,
		_w46_,
		_w134_,
		_w79_,
		_w2052_
	);
	LUT4 #(
		.INIT('h0800)
	) name2027 (
		_w1234_,
		_w1271_,
		_w272_,
		_w2052_,
		_w2053_
	);
	LUT3 #(
		.INIT('h80)
	) name2028 (
		_w657_,
		_w2051_,
		_w2053_,
		_w2054_
	);
	LUT4 #(
		.INIT('h135f)
	) name2029 (
		_w82_,
		_w54_,
		_w71_,
		_w72_,
		_w2055_
	);
	LUT4 #(
		.INIT('h1000)
	) name2030 (
		_w117_,
		_w256_,
		_w258_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h8000)
	) name2031 (
		_w657_,
		_w2051_,
		_w2053_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('h0777)
	) name2032 (
		_w206_,
		_w121_,
		_w77_,
		_w98_,
		_w2058_
	);
	LUT4 #(
		.INIT('h0100)
	) name2033 (
		_w124_,
		_w132_,
		_w171_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h0777)
	) name2034 (
		_w85_,
		_w91_,
		_w77_,
		_w100_,
		_w2060_
	);
	LUT3 #(
		.INIT('h10)
	) name2035 (
		_w184_,
		_w182_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h1000)
	) name2036 (
		_w168_,
		_w86_,
		_w254_,
		_w217_,
		_w2062_
	);
	LUT3 #(
		.INIT('h80)
	) name2037 (
		_w2059_,
		_w2061_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h0777)
	) name2038 (
		_w88_,
		_w68_,
		_w116_,
		_w71_,
		_w2064_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		_w297_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h8000)
	) name2040 (
		_w640_,
		_w509_,
		_w531_,
		_w1729_,
		_w2066_
	);
	LUT3 #(
		.INIT('h80)
	) name2041 (
		_w1341_,
		_w2065_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h80)
	) name2042 (
		_w2063_,
		_w2057_,
		_w2067_,
		_w2068_
	);
	LUT3 #(
		.INIT('h8e)
	) name2043 (
		_w2035_,
		_w2049_,
		_w2068_,
		_w2069_
	);
	LUT3 #(
		.INIT('h54)
	) name2044 (
		_w2033_,
		_w2034_,
		_w2069_,
		_w2070_
	);
	LUT3 #(
		.INIT('h96)
	) name2045 (
		_w1935_,
		_w1937_,
		_w2032_,
		_w2071_
	);
	LUT2 #(
		.INIT('h9)
	) name2046 (
		_w2069_,
		_w2071_,
		_w2072_
	);
	LUT3 #(
		.INIT('h06)
	) name2047 (
		_w2010_,
		_w2070_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('h90)
	) name2048 (
		_w2010_,
		_w2070_,
		_w2072_,
		_w2074_
	);
	LUT3 #(
		.INIT('h69)
	) name2049 (
		_w2010_,
		_w2070_,
		_w2072_,
		_w2075_
	);
	LUT2 #(
		.INIT('h9)
	) name2050 (
		\a[22] ,
		\a[23] ,
		_w2076_
	);
	LUT4 #(
		.INIT('h0069)
	) name2051 (
		_w2010_,
		_w2070_,
		_w2072_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name2052 (
		_w46_,
		_w70_,
		_w100_,
		_w72_,
		_w2078_
	);
	LUT3 #(
		.INIT('h10)
	) name2053 (
		_w156_,
		_w157_,
		_w2078_,
		_w2079_
	);
	LUT3 #(
		.INIT('h80)
	) name2054 (
		_w276_,
		_w1192_,
		_w1323_,
		_w2080_
	);
	LUT3 #(
		.INIT('h80)
	) name2055 (
		_w381_,
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		_w539_,
		_w518_,
		_w2082_
	);
	LUT3 #(
		.INIT('h57)
	) name2057 (
		_w88_,
		_w59_,
		_w68_,
		_w2083_
	);
	LUT4 #(
		.INIT('h0400)
	) name2058 (
		_w162_,
		_w165_,
		_w286_,
		_w2083_,
		_w2084_
	);
	LUT4 #(
		.INIT('h8000)
	) name2059 (
		_w817_,
		_w820_,
		_w2082_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('h80)
	) name2060 (
		_w246_,
		_w2081_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		_w1321_,
		_w2086_,
		_w2087_
	);
	LUT3 #(
		.INIT('h1e)
	) name2062 (
		_w1805_,
		_w1949_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2063 (
		_w1780_,
		_w1951_,
		_w1953_,
		_w2088_,
		_w2089_
	);
	LUT3 #(
		.INIT('h87)
	) name2064 (
		_w1805_,
		_w1949_,
		_w2087_,
		_w2090_
	);
	LUT4 #(
		.INIT('h804c)
	) name2065 (
		_w1805_,
		_w1810_,
		_w1949_,
		_w2087_,
		_w2091_
	);
	LUT2 #(
		.INIT('h4)
	) name2066 (
		_w1806_,
		_w1811_,
		_w2092_
	);
	LUT3 #(
		.INIT('h84)
	) name2067 (
		_w1805_,
		_w1813_,
		_w1949_,
		_w2093_
	);
	LUT3 #(
		.INIT('h01)
	) name2068 (
		_w2091_,
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2069 (
		_w1401_,
		_w1437_,
		_w1448_,
		_w1526_,
		_w2095_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2070 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1528_,
		_w2096_
	);
	LUT3 #(
		.INIT('h90)
	) name2071 (
		_w1377_,
		_w1379_,
		_w1531_,
		_w2097_
	);
	LUT3 #(
		.INIT('h07)
	) name2072 (
		_w1400_,
		_w1530_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w2096_,
		_w2098_,
		_w2099_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2074 (
		_w1407_,
		_w1431_,
		_w1432_,
		_w1460_,
		_w2100_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2075 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1462_,
		_w2101_
	);
	LUT3 #(
		.INIT('h90)
	) name2076 (
		_w1370_,
		_w1372_,
		_w1464_,
		_w2102_
	);
	LUT3 #(
		.INIT('h07)
	) name2077 (
		_w1405_,
		_w1466_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h4)
	) name2078 (
		_w2101_,
		_w2103_,
		_w2104_
	);
	LUT3 #(
		.INIT('h14)
	) name2079 (
		_w424_,
		_w1360_,
		_w1362_,
		_w2105_
	);
	LUT3 #(
		.INIT('h90)
	) name2080 (
		_w1424_,
		_w1426_,
		_w1475_,
		_w2106_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2081 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1479_,
		_w2107_
	);
	LUT3 #(
		.INIT('h90)
	) name2082 (
		_w1363_,
		_w1365_,
		_w1514_,
		_w2108_
	);
	LUT3 #(
		.INIT('h07)
	) name2083 (
		_w1411_,
		_w1477_,
		_w2108_,
		_w2109_
	);
	LUT2 #(
		.INIT('h4)
	) name2084 (
		_w2107_,
		_w2109_,
		_w2110_
	);
	LUT3 #(
		.INIT('h65)
	) name2085 (
		_w2105_,
		_w2106_,
		_w2110_,
		_w2111_
	);
	LUT3 #(
		.INIT('h41)
	) name2086 (
		_w424_,
		_w1357_,
		_w1359_,
		_w2112_
	);
	LUT3 #(
		.INIT('h40)
	) name2087 (
		_w1968_,
		_w1971_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h0d)
	) name2088 (
		_w1972_,
		_w1975_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h9)
	) name2089 (
		_w2111_,
		_w2114_,
		_w2115_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2090 (
		_w366_,
		_w2100_,
		_w2104_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('h659a)
	) name2091 (
		_w366_,
		_w2100_,
		_w2104_,
		_w2115_,
		_w2117_
	);
	LUT4 #(
		.INIT('hd400)
	) name2092 (
		_w1966_,
		_w1976_,
		_w1980_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2093 (
		_w1966_,
		_w1981_,
		_w1982_,
		_w2117_,
		_w2119_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2094 (
		_w581_,
		_w2095_,
		_w2099_,
		_w2119_,
		_w2120_
	);
	LUT4 #(
		.INIT('h659a)
	) name2095 (
		_w581_,
		_w2095_,
		_w2099_,
		_w2119_,
		_w2121_
	);
	LUT4 #(
		.INIT('h7100)
	) name2096 (
		_w1961_,
		_w1965_,
		_w1984_,
		_w2121_,
		_w2122_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2097 (
		_w1961_,
		_w1985_,
		_w1986_,
		_w2121_,
		_w2123_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2098 (
		_w37_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w2124_
	);
	LUT4 #(
		.INIT('h802a)
	) name2099 (
		_w1450_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w1454_,
		_w1741_,
		_w2126_
	);
	LUT3 #(
		.INIT('h82)
	) name2101 (
		_w1453_,
		_w1739_,
		_w1785_,
		_w2127_
	);
	LUT3 #(
		.INIT('h01)
	) name2102 (
		_w2125_,
		_w2126_,
		_w2127_,
		_w2128_
	);
	LUT4 #(
		.INIT('h8488)
	) name2103 (
		_w30_,
		_w2123_,
		_w2124_,
		_w2128_,
		_w2129_
	);
	LUT4 #(
		.INIT('h6966)
	) name2104 (
		_w30_,
		_w2123_,
		_w2124_,
		_w2128_,
		_w2130_
	);
	LUT4 #(
		.INIT('hd400)
	) name2105 (
		_w1960_,
		_w1988_,
		_w1993_,
		_w2130_,
		_w2131_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2106 (
		_w1960_,
		_w1994_,
		_w1995_,
		_w2130_,
		_w2132_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2107 (
		_w33_,
		_w2089_,
		_w2094_,
		_w2132_,
		_w2133_
	);
	LUT4 #(
		.INIT('h659a)
	) name2108 (
		_w33_,
		_w2089_,
		_w2094_,
		_w2132_,
		_w2134_
	);
	LUT4 #(
		.INIT('h153f)
	) name2109 (
		_w85_,
		_w96_,
		_w116_,
		_w100_,
		_w2135_
	);
	LUT4 #(
		.INIT('h4000)
	) name2110 (
		_w272_,
		_w276_,
		_w666_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h4)
	) name2111 (
		_w152_,
		_w1255_,
		_w2137_
	);
	LUT4 #(
		.INIT('h37bf)
	) name2112 (
		_w46_,
		_w95_,
		_w98_,
		_w100_,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		_w814_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h4000)
	) name2114 (
		_w152_,
		_w814_,
		_w1255_,
		_w2138_,
		_w2140_
	);
	LUT4 #(
		.INIT('h0002)
	) name2115 (
		_w1385_,
		_w252_,
		_w242_,
		_w181_,
		_w2141_
	);
	LUT4 #(
		.INIT('h8000)
	) name2116 (
		_w2026_,
		_w2141_,
		_w2136_,
		_w2140_,
		_w2142_
	);
	LUT4 #(
		.INIT('h8000)
	) name2117 (
		_w1222_,
		_w2013_,
		_w2018_,
		_w2142_,
		_w2143_
	);
	LUT4 #(
		.INIT('h001e)
	) name2118 (
		_w1998_,
		_w2000_,
		_w2134_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2119 (
		_w1998_,
		_w2000_,
		_w2134_,
		_w2143_,
		_w2145_
	);
	LUT4 #(
		.INIT('hb200)
	) name2120 (
		_w2001_,
		_w2007_,
		_w2070_,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h23dc)
	) name2121 (
		_w2008_,
		_w2009_,
		_w2070_,
		_w2145_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		_w2073_,
		_w2147_,
		_w2148_
	);
	LUT3 #(
		.INIT('h1e)
	) name2123 (
		_w2073_,
		_w2077_,
		_w2147_,
		_w2149_
	);
	LUT4 #(
		.INIT('h010f)
	) name2124 (
		_w1998_,
		_w2000_,
		_w2133_,
		_w2134_,
		_w2150_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2125 (
		_w1951_,
		_w1953_,
		_w2090_,
		_w2088_,
		_w2151_
	);
	LUT3 #(
		.INIT('h02)
	) name2126 (
		_w1950_,
		_w1953_,
		_w2087_,
		_w2152_
	);
	LUT3 #(
		.INIT('h84)
	) name2127 (
		_w1805_,
		_w1811_,
		_w1949_,
		_w2153_
	);
	LUT4 #(
		.INIT('h804c)
	) name2128 (
		_w1805_,
		_w1813_,
		_w1949_,
		_w2087_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name2129 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h5700)
	) name2130 (
		_w1780_,
		_w2151_,
		_w2152_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h9)
	) name2131 (
		_w33_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		_w1400_,
		_w1531_,
		_w2158_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2133 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1530_,
		_w2159_
	);
	LUT4 #(
		.INIT('h000d)
	) name2134 (
		_w1528_,
		_w1741_,
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2135 (
		_w1526_,
		_w1720_,
		_w1744_,
		_w2160_,
		_w2161_
	);
	LUT3 #(
		.INIT('h90)
	) name2136 (
		_w1433_,
		_w1435_,
		_w1460_,
		_w2162_
	);
	LUT3 #(
		.INIT('h90)
	) name2137 (
		_w1377_,
		_w1379_,
		_w1462_,
		_w2163_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2138 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1466_,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		_w1405_,
		_w1464_,
		_w2165_
	);
	LUT2 #(
		.INIT('h1)
	) name2140 (
		_w2164_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w2163_,
		_w2166_,
		_w2167_
	);
	LUT3 #(
		.INIT('h14)
	) name2142 (
		_w424_,
		_w1363_,
		_w1365_,
		_w2168_
	);
	LUT3 #(
		.INIT('h90)
	) name2143 (
		_w1427_,
		_w1429_,
		_w1475_,
		_w2169_
	);
	LUT3 #(
		.INIT('h90)
	) name2144 (
		_w1370_,
		_w1372_,
		_w1479_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		_w1411_,
		_w1514_,
		_w2171_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2146 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1477_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name2148 (
		_w2170_,
		_w2173_,
		_w2174_
	);
	LUT3 #(
		.INIT('h65)
	) name2149 (
		_w2168_,
		_w2169_,
		_w2174_,
		_w2175_
	);
	LUT3 #(
		.INIT('h41)
	) name2150 (
		_w424_,
		_w1360_,
		_w1362_,
		_w2176_
	);
	LUT3 #(
		.INIT('h40)
	) name2151 (
		_w2106_,
		_w2110_,
		_w2176_,
		_w2177_
	);
	LUT3 #(
		.INIT('h0d)
	) name2152 (
		_w2111_,
		_w2114_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h9)
	) name2153 (
		_w2175_,
		_w2178_,
		_w2179_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2154 (
		_w366_,
		_w2162_,
		_w2167_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h659a)
	) name2155 (
		_w366_,
		_w2162_,
		_w2167_,
		_w2179_,
		_w2181_
	);
	LUT3 #(
		.INIT('h1e)
	) name2156 (
		_w2116_,
		_w2118_,
		_w2181_,
		_w2182_
	);
	LUT3 #(
		.INIT('h60)
	) name2157 (
		_w581_,
		_w2161_,
		_w2182_,
		_w2183_
	);
	LUT3 #(
		.INIT('h96)
	) name2158 (
		_w581_,
		_w2161_,
		_w2182_,
		_w2184_
	);
	LUT3 #(
		.INIT('h1e)
	) name2159 (
		_w2120_,
		_w2122_,
		_w2184_,
		_w2185_
	);
	LUT3 #(
		.INIT('h82)
	) name2160 (
		_w1454_,
		_w1739_,
		_w1785_,
		_w2186_
	);
	LUT4 #(
		.INIT('h802a)
	) name2161 (
		_w1453_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2187_
	);
	LUT4 #(
		.INIT('h000d)
	) name2162 (
		_w1450_,
		_w1806_,
		_w2186_,
		_w2187_,
		_w2188_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2163 (
		_w37_,
		_w1798_,
		_w1809_,
		_w2188_,
		_w2189_
	);
	LUT3 #(
		.INIT('h48)
	) name2164 (
		_w30_,
		_w2185_,
		_w2189_,
		_w2190_
	);
	LUT3 #(
		.INIT('h96)
	) name2165 (
		_w30_,
		_w2185_,
		_w2189_,
		_w2191_
	);
	LUT3 #(
		.INIT('h1e)
	) name2166 (
		_w2129_,
		_w2131_,
		_w2191_,
		_w2192_
	);
	LUT3 #(
		.INIT('h60)
	) name2167 (
		_w33_,
		_w2156_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('h09)
	) name2168 (
		_w33_,
		_w2156_,
		_w2192_,
		_w2194_
	);
	LUT3 #(
		.INIT('h96)
	) name2169 (
		_w33_,
		_w2156_,
		_w2192_,
		_w2195_
	);
	LUT4 #(
		.INIT('h2f7f)
	) name2170 (
		_w46_,
		_w82_,
		_w95_,
		_w116_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name2171 (
		_w179_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h10)
	) name2172 (
		_w316_,
		_w168_,
		_w675_,
		_w2198_
	);
	LUT4 #(
		.INIT('h0777)
	) name2173 (
		_w88_,
		_w59_,
		_w85_,
		_w91_,
		_w2199_
	);
	LUT3 #(
		.INIT('h80)
	) name2174 (
		_w335_,
		_w428_,
		_w2199_,
		_w2200_
	);
	LUT4 #(
		.INIT('h0777)
	) name2175 (
		_w206_,
		_w85_,
		_w116_,
		_w71_,
		_w2201_
	);
	LUT3 #(
		.INIT('h20)
	) name2176 (
		_w435_,
		_w211_,
		_w2201_,
		_w2202_
	);
	LUT4 #(
		.INIT('h8000)
	) name2177 (
		_w2197_,
		_w2198_,
		_w2200_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h8000)
	) name2178 (
		_w223_,
		_w235_,
		_w2039_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h09)
	) name2179 (
		_w2150_,
		_w2195_,
		_w2204_,
		_w2205_
	);
	LUT3 #(
		.INIT('h96)
	) name2180 (
		_w2150_,
		_w2195_,
		_w2204_,
		_w2206_
	);
	LUT3 #(
		.INIT('h1e)
	) name2181 (
		_w2144_,
		_w2146_,
		_w2206_,
		_w2207_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		_w2148_,
		_w2207_,
		_w2208_
	);
	LUT3 #(
		.INIT('h21)
	) name2183 (
		_w2073_,
		_w2075_,
		_w2147_,
		_w2209_
	);
	LUT4 #(
		.INIT('h050b)
	) name2184 (
		_w2073_,
		_w2074_,
		_w2076_,
		_w2147_,
		_w2210_
	);
	LUT3 #(
		.INIT('h96)
	) name2185 (
		_w2148_,
		_w2207_,
		_w2210_,
		_w2211_
	);
	LUT3 #(
		.INIT('h90)
	) name2186 (
		_w2148_,
		_w2207_,
		_w2209_,
		_w2212_
	);
	LUT4 #(
		.INIT('h1455)
	) name2187 (
		_w2076_,
		_w2148_,
		_w2207_,
		_w2209_,
		_w2213_
	);
	LUT4 #(
		.INIT('h010f)
	) name2188 (
		_w2144_,
		_w2146_,
		_w2205_,
		_w2206_,
		_w2214_
	);
	LUT4 #(
		.INIT('h010f)
	) name2189 (
		_w2129_,
		_w2131_,
		_w2190_,
		_w2191_,
		_w2215_
	);
	LUT4 #(
		.INIT('h1151)
	) name2190 (
		_w1811_,
		_w1780_,
		_w1950_,
		_w1953_,
		_w2216_
	);
	LUT3 #(
		.INIT('ha6)
	) name2191 (
		_w33_,
		_w2090_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h010f)
	) name2192 (
		_w2120_,
		_w2122_,
		_w2183_,
		_w2184_,
		_w2218_
	);
	LUT3 #(
		.INIT('h82)
	) name2193 (
		_w1528_,
		_w1739_,
		_w1785_,
		_w2219_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2194 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1531_,
		_w2220_
	);
	LUT3 #(
		.INIT('h0d)
	) name2195 (
		_w1530_,
		_w1741_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h4)
	) name2196 (
		_w2219_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h6a55)
	) name2197 (
		_w581_,
		_w1526_,
		_w1827_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h010f)
	) name2198 (
		_w2116_,
		_w2118_,
		_w2180_,
		_w2181_,
		_w2224_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2199 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1464_,
		_w2225_
	);
	LUT4 #(
		.INIT('h006f)
	) name2200 (
		_w1377_,
		_w1379_,
		_w1466_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h70)
	) name2201 (
		_w1400_,
		_w1462_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2202 (
		_w366_,
		_w1460_,
		_w1622_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w424_,
		_w1411_,
		_w2229_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2204 (
		_w1269_,
		_w1368_,
		_w1369_,
		_w1514_,
		_w2230_
	);
	LUT4 #(
		.INIT('h006f)
	) name2205 (
		_w1370_,
		_w1372_,
		_w1477_,
		_w2230_,
		_w2231_
	);
	LUT3 #(
		.INIT('h70)
	) name2206 (
		_w1405_,
		_w1479_,
		_w2231_,
		_w2232_
	);
	LUT4 #(
		.INIT('h780f)
	) name2207 (
		_w1475_,
		_w1527_,
		_w2229_,
		_w2232_,
		_w2233_
	);
	LUT3 #(
		.INIT('h41)
	) name2208 (
		_w424_,
		_w1363_,
		_w1365_,
		_w2234_
	);
	LUT3 #(
		.INIT('h40)
	) name2209 (
		_w2169_,
		_w2174_,
		_w2234_,
		_w2235_
	);
	LUT4 #(
		.INIT('hf020)
	) name2210 (
		_w2175_,
		_w2178_,
		_w2233_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h0fd2)
	) name2211 (
		_w2175_,
		_w2178_,
		_w2233_,
		_w2235_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		_w2228_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w2228_,
		_w2237_,
		_w2239_
	);
	LUT2 #(
		.INIT('h6)
	) name2214 (
		_w2228_,
		_w2237_,
		_w2240_
	);
	LUT2 #(
		.INIT('h9)
	) name2215 (
		_w2224_,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w2223_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name2217 (
		_w2223_,
		_w2241_,
		_w2243_
	);
	LUT2 #(
		.INIT('h9)
	) name2218 (
		_w2223_,
		_w2241_,
		_w2244_
	);
	LUT2 #(
		.INIT('h9)
	) name2219 (
		_w2218_,
		_w2244_,
		_w2245_
	);
	LUT3 #(
		.INIT('h82)
	) name2220 (
		_w1450_,
		_w1805_,
		_w1949_,
		_w2246_
	);
	LUT4 #(
		.INIT('h802a)
	) name2221 (
		_w1454_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2247_
	);
	LUT3 #(
		.INIT('h0d)
	) name2222 (
		_w1453_,
		_w1806_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name2223 (
		_w2246_,
		_w2248_,
		_w2249_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2224 (
		_w30_,
		_w37_,
		_w1954_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w2245_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name2226 (
		_w2245_,
		_w2250_,
		_w2252_
	);
	LUT2 #(
		.INIT('h6)
	) name2227 (
		_w2245_,
		_w2250_,
		_w2253_
	);
	LUT3 #(
		.INIT('h41)
	) name2228 (
		_w2215_,
		_w2217_,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('h96)
	) name2229 (
		_w2215_,
		_w2217_,
		_w2253_,
		_w2255_
	);
	LUT4 #(
		.INIT('h7100)
	) name2230 (
		_w2150_,
		_w2157_,
		_w2192_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2231 (
		_w2150_,
		_w2193_,
		_w2194_,
		_w2255_,
		_w2257_
	);
	LUT3 #(
		.INIT('h80)
	) name2232 (
		_w120_,
		_w320_,
		_w2059_,
		_w2258_
	);
	LUT4 #(
		.INIT('h0777)
	) name2233 (
		_w206_,
		_w88_,
		_w54_,
		_w91_,
		_w2259_
	);
	LUT4 #(
		.INIT('h2000)
	) name2234 (
		_w537_,
		_w225_,
		_w1197_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('h80)
	) name2235 (
		_w565_,
		_w2137_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h8000)
	) name2236 (
		_w810_,
		_w1152_,
		_w2261_,
		_w2258_,
		_w2262_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w2257_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w2257_,
		_w2262_,
		_w2264_
	);
	LUT2 #(
		.INIT('h9)
	) name2239 (
		_w2257_,
		_w2262_,
		_w2265_
	);
	LUT2 #(
		.INIT('h9)
	) name2240 (
		_w2214_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h8008)
	) name2241 (
		_w2148_,
		_w2207_,
		_w2214_,
		_w2265_,
		_w2267_
	);
	LUT4 #(
		.INIT('h7887)
	) name2242 (
		_w2148_,
		_w2207_,
		_w2214_,
		_w2265_,
		_w2268_
	);
	LUT2 #(
		.INIT('h6)
	) name2243 (
		_w2213_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2244 (
		_w1526_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w2270_
	);
	LUT4 #(
		.INIT('h802a)
	) name2245 (
		_w1528_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		_w1531_,
		_w1741_,
		_w2272_
	);
	LUT3 #(
		.INIT('h82)
	) name2247 (
		_w1530_,
		_w1739_,
		_w1785_,
		_w2273_
	);
	LUT3 #(
		.INIT('h01)
	) name2248 (
		_w2271_,
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2249 (
		_w1401_,
		_w1437_,
		_w1448_,
		_w1460_,
		_w2275_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2250 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1462_,
		_w2276_
	);
	LUT3 #(
		.INIT('h90)
	) name2251 (
		_w1377_,
		_w1379_,
		_w1464_,
		_w2277_
	);
	LUT3 #(
		.INIT('h07)
	) name2252 (
		_w1400_,
		_w1466_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name2253 (
		_w2276_,
		_w2278_,
		_w2279_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2254 (
		_w1407_,
		_w1431_,
		_w1432_,
		_w1475_,
		_w2280_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2255 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1479_,
		_w2281_
	);
	LUT3 #(
		.INIT('h90)
	) name2256 (
		_w1370_,
		_w1372_,
		_w1514_,
		_w2282_
	);
	LUT3 #(
		.INIT('h07)
	) name2257 (
		_w1405_,
		_w1477_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h4)
	) name2258 (
		_w2281_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h0154)
	) name2259 (
		_w424_,
		_w1269_,
		_w1368_,
		_w1369_,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name2260 (
		_w33_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h9)
	) name2261 (
		_w33_,
		_w2285_,
		_w2287_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2262 (
		_w424_,
		_w2280_,
		_w2284_,
		_w2287_,
		_w2288_
	);
	LUT4 #(
		.INIT('h659a)
	) name2263 (
		_w424_,
		_w2280_,
		_w2284_,
		_w2287_,
		_w2289_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		_w424_,
		_w1411_,
		_w2290_
	);
	LUT4 #(
		.INIT('h7000)
	) name2265 (
		_w1475_,
		_w1527_,
		_w2232_,
		_w2290_,
		_w2291_
	);
	LUT3 #(
		.INIT('hc8)
	) name2266 (
		_w2236_,
		_w2289_,
		_w2291_,
		_w2292_
	);
	LUT3 #(
		.INIT('h36)
	) name2267 (
		_w2236_,
		_w2289_,
		_w2291_,
		_w2293_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2268 (
		_w366_,
		_w2275_,
		_w2279_,
		_w2293_,
		_w2294_
	);
	LUT4 #(
		.INIT('h659a)
	) name2269 (
		_w366_,
		_w2275_,
		_w2279_,
		_w2293_,
		_w2295_
	);
	LUT4 #(
		.INIT('hd400)
	) name2270 (
		_w2224_,
		_w2228_,
		_w2237_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2271 (
		_w2224_,
		_w2238_,
		_w2239_,
		_w2295_,
		_w2297_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2272 (
		_w581_,
		_w2270_,
		_w2274_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('h659a)
	) name2273 (
		_w581_,
		_w2270_,
		_w2274_,
		_w2297_,
		_w2299_
	);
	LUT4 #(
		.INIT('h7100)
	) name2274 (
		_w2218_,
		_w2223_,
		_w2241_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2275 (
		_w2218_,
		_w2242_,
		_w2243_,
		_w2299_,
		_w2301_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2276 (
		_w37_,
		_w1951_,
		_w1953_,
		_w2088_,
		_w2302_
	);
	LUT4 #(
		.INIT('h802a)
	) name2277 (
		_w1450_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name2278 (
		_w1454_,
		_w1806_,
		_w2304_
	);
	LUT3 #(
		.INIT('h82)
	) name2279 (
		_w1453_,
		_w1805_,
		_w1949_,
		_w2305_
	);
	LUT3 #(
		.INIT('h01)
	) name2280 (
		_w2303_,
		_w2304_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('h8488)
	) name2281 (
		_w30_,
		_w2301_,
		_w2302_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('h6966)
	) name2282 (
		_w30_,
		_w2301_,
		_w2302_,
		_w2306_,
		_w2308_
	);
	LUT4 #(
		.INIT('hd400)
	) name2283 (
		_w2217_,
		_w2245_,
		_w2250_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('h002b)
	) name2284 (
		_w2217_,
		_w2245_,
		_w2250_,
		_w2308_,
		_w2310_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2285 (
		_w2217_,
		_w2251_,
		_w2252_,
		_w2308_,
		_w2311_
	);
	LUT3 #(
		.INIT('h80)
	) name2286 (
		_w456_,
		_w243_,
		_w813_,
		_w2312_
	);
	LUT4 #(
		.INIT('h153f)
	) name2287 (
		_w206_,
		_w88_,
		_w62_,
		_w96_,
		_w2313_
	);
	LUT3 #(
		.INIT('h10)
	) name2288 (
		_w316_,
		_w168_,
		_w2313_,
		_w2314_
	);
	LUT3 #(
		.INIT('h80)
	) name2289 (
		_w1314_,
		_w2314_,
		_w2312_,
		_w2315_
	);
	LUT4 #(
		.INIT('h8000)
	) name2290 (
		_w296_,
		_w534_,
		_w1348_,
		_w2315_,
		_w2316_
	);
	LUT4 #(
		.INIT('h001e)
	) name2291 (
		_w2254_,
		_w2256_,
		_w2311_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2292 (
		_w2254_,
		_w2256_,
		_w2311_,
		_w2316_,
		_w2318_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2293 (
		_w2214_,
		_w2257_,
		_w2262_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2294 (
		_w2214_,
		_w2263_,
		_w2264_,
		_w2318_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		_w2267_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h6)
	) name2296 (
		_w2267_,
		_w2320_,
		_w2322_
	);
	LUT3 #(
		.INIT('h51)
	) name2297 (
		_w2076_,
		_w2212_,
		_w2268_,
		_w2323_
	);
	LUT2 #(
		.INIT('h6)
	) name2298 (
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2299 (
		_w2254_,
		_w2256_,
		_w2309_,
		_w2310_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w2300_,
		_w2307_,
		_w2326_
	);
	LUT3 #(
		.INIT('h82)
	) name2301 (
		_w1454_,
		_w1805_,
		_w1949_,
		_w2327_
	);
	LUT4 #(
		.INIT('h802a)
	) name2302 (
		_w1453_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w2327_,
		_w2328_,
		_w2329_
	);
	LUT4 #(
		.INIT('h5700)
	) name2304 (
		_w37_,
		_w2151_,
		_w2152_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		_w2296_,
		_w2298_,
		_w2331_
	);
	LUT3 #(
		.INIT('h82)
	) name2306 (
		_w1531_,
		_w1739_,
		_w1785_,
		_w2332_
	);
	LUT4 #(
		.INIT('h802a)
	) name2307 (
		_w1530_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2333_
	);
	LUT4 #(
		.INIT('h000d)
	) name2308 (
		_w1528_,
		_w1806_,
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2309 (
		_w1526_,
		_w1798_,
		_w1809_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name2310 (
		_w2292_,
		_w2294_,
		_w2336_
	);
	LUT2 #(
		.INIT('h8)
	) name2311 (
		_w1400_,
		_w1464_,
		_w2337_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2312 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1466_,
		_w2338_
	);
	LUT4 #(
		.INIT('h000d)
	) name2313 (
		_w1462_,
		_w1741_,
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2314 (
		_w1460_,
		_w1720_,
		_w1744_,
		_w2339_,
		_w2340_
	);
	LUT3 #(
		.INIT('h90)
	) name2315 (
		_w1433_,
		_w1435_,
		_w1475_,
		_w2341_
	);
	LUT3 #(
		.INIT('h90)
	) name2316 (
		_w1377_,
		_w1379_,
		_w1479_,
		_w2342_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2317 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1477_,
		_w2343_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		_w1405_,
		_w1514_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w2343_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name2320 (
		_w2342_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h9a)
	) name2321 (
		_w424_,
		_w2341_,
		_w2346_,
		_w2347_
	);
	LUT4 #(
		.INIT('h0041)
	) name2322 (
		_w424_,
		_w1370_,
		_w1372_,
		_w33_,
		_w2348_
	);
	LUT4 #(
		.INIT('h41be)
	) name2323 (
		_w424_,
		_w1370_,
		_w1372_,
		_w33_,
		_w2349_
	);
	LUT3 #(
		.INIT('h1e)
	) name2324 (
		_w2286_,
		_w2288_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		_w2347_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w2347_,
		_w2350_,
		_w2352_
	);
	LUT2 #(
		.INIT('h6)
	) name2327 (
		_w2347_,
		_w2350_,
		_w2353_
	);
	LUT3 #(
		.INIT('h96)
	) name2328 (
		_w366_,
		_w2340_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name2329 (
		_w2336_,
		_w2354_,
		_w2355_
	);
	LUT2 #(
		.INIT('h2)
	) name2330 (
		_w2336_,
		_w2354_,
		_w2356_
	);
	LUT2 #(
		.INIT('h9)
	) name2331 (
		_w2336_,
		_w2354_,
		_w2357_
	);
	LUT3 #(
		.INIT('h96)
	) name2332 (
		_w581_,
		_w2335_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name2333 (
		_w2331_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w2331_,
		_w2358_,
		_w2360_
	);
	LUT2 #(
		.INIT('h9)
	) name2335 (
		_w2331_,
		_w2358_,
		_w2361_
	);
	LUT3 #(
		.INIT('h96)
	) name2336 (
		_w30_,
		_w2330_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h4)
	) name2337 (
		_w2326_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w2326_,
		_w2362_,
		_w2364_
	);
	LUT2 #(
		.INIT('h9)
	) name2339 (
		_w2326_,
		_w2362_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		_w197_,
		_w1318_,
		_w2366_
	);
	LUT3 #(
		.INIT('h04)
	) name2341 (
		_w209_,
		_w1234_,
		_w86_,
		_w2367_
	);
	LUT3 #(
		.INIT('h80)
	) name2342 (
		_w2139_,
		_w2367_,
		_w2366_,
		_w2368_
	);
	LUT4 #(
		.INIT('h135f)
	) name2343 (
		_w106_,
		_w54_,
		_w68_,
		_w125_,
		_w2369_
	);
	LUT4 #(
		.INIT('h135f)
	) name2344 (
		_w121_,
		_w54_,
		_w62_,
		_w72_,
		_w2370_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT3 #(
		.INIT('h10)
	) name2346 (
		_w308_,
		_w347_,
		_w250_,
		_w2372_
	);
	LUT3 #(
		.INIT('h80)
	) name2347 (
		_w1242_,
		_w2371_,
		_w2372_,
		_w2373_
	);
	LUT4 #(
		.INIT('h8000)
	) name2348 (
		_w1731_,
		_w2081_,
		_w2368_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('h09)
	) name2349 (
		_w2325_,
		_w2365_,
		_w2374_,
		_w2375_
	);
	LUT3 #(
		.INIT('h96)
	) name2350 (
		_w2325_,
		_w2365_,
		_w2374_,
		_w2376_
	);
	LUT3 #(
		.INIT('h1e)
	) name2351 (
		_w2317_,
		_w2319_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w2321_,
		_w2377_,
		_w2378_
	);
	LUT4 #(
		.INIT('h8004)
	) name2353 (
		_w2208_,
		_w2212_,
		_w2266_,
		_w2320_,
		_w2379_
	);
	LUT4 #(
		.INIT('h3c69)
	) name2354 (
		_w2076_,
		_w2321_,
		_w2377_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h010f)
	) name2355 (
		_w2317_,
		_w2319_,
		_w2375_,
		_w2376_,
		_w2381_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2356 (
		_w30_,
		_w2330_,
		_w2359_,
		_w2360_,
		_w2382_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2357 (
		_w581_,
		_w2335_,
		_w2355_,
		_w2356_,
		_w2383_
	);
	LUT4 #(
		.INIT('h1151)
	) name2358 (
		_w1454_,
		_w37_,
		_w1950_,
		_w1953_,
		_w2384_
	);
	LUT4 #(
		.INIT('h0509)
	) name2359 (
		_w30_,
		_w2090_,
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT4 #(
		.INIT('ha060)
	) name2360 (
		_w30_,
		_w2090_,
		_w2383_,
		_w2384_,
		_w2386_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2361 (
		_w30_,
		_w2090_,
		_w2383_,
		_w2384_,
		_w2387_
	);
	LUT3 #(
		.INIT('h82)
	) name2362 (
		_w1528_,
		_w1805_,
		_w1949_,
		_w2388_
	);
	LUT4 #(
		.INIT('h802a)
	) name2363 (
		_w1531_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2389_
	);
	LUT3 #(
		.INIT('h0d)
	) name2364 (
		_w1530_,
		_w1806_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h4)
	) name2365 (
		_w2388_,
		_w2390_,
		_w2391_
	);
	LUT4 #(
		.INIT('h6a55)
	) name2366 (
		_w581_,
		_w1526_,
		_w1954_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2367 (
		_w366_,
		_w2340_,
		_w2351_,
		_w2352_,
		_w2393_
	);
	LUT3 #(
		.INIT('h82)
	) name2368 (
		_w1462_,
		_w1739_,
		_w1785_,
		_w2394_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2369 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1464_,
		_w2395_
	);
	LUT3 #(
		.INIT('h0d)
	) name2370 (
		_w1466_,
		_w1741_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name2371 (
		_w2394_,
		_w2396_,
		_w2397_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2372 (
		_w366_,
		_w1460_,
		_w1827_,
		_w2397_,
		_w2398_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2373 (
		_w1213_,
		_w1375_,
		_w1376_,
		_w1514_,
		_w2399_
	);
	LUT4 #(
		.INIT('h006f)
	) name2374 (
		_w1377_,
		_w1379_,
		_w1477_,
		_w2399_,
		_w2400_
	);
	LUT3 #(
		.INIT('h70)
	) name2375 (
		_w1400_,
		_w1479_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2376 (
		_w424_,
		_w1475_,
		_w1622_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('h010f)
	) name2377 (
		_w2286_,
		_w2288_,
		_w2348_,
		_w2349_,
		_w2403_
	);
	LUT3 #(
		.INIT('h10)
	) name2378 (
		_w424_,
		_w33_,
		_w1405_,
		_w2404_
	);
	LUT3 #(
		.INIT('h8c)
	) name2379 (
		_w424_,
		_w33_,
		_w1405_,
		_w2405_
	);
	LUT3 #(
		.INIT('h63)
	) name2380 (
		_w424_,
		_w33_,
		_w1405_,
		_w2406_
	);
	LUT3 #(
		.INIT('h82)
	) name2381 (
		_w2402_,
		_w2403_,
		_w2406_,
		_w2407_
	);
	LUT3 #(
		.INIT('h14)
	) name2382 (
		_w2402_,
		_w2403_,
		_w2406_,
		_w2408_
	);
	LUT3 #(
		.INIT('h69)
	) name2383 (
		_w2402_,
		_w2403_,
		_w2406_,
		_w2409_
	);
	LUT3 #(
		.INIT('h14)
	) name2384 (
		_w2393_,
		_w2398_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('h82)
	) name2385 (
		_w2393_,
		_w2398_,
		_w2409_,
		_w2411_
	);
	LUT3 #(
		.INIT('h69)
	) name2386 (
		_w2393_,
		_w2398_,
		_w2409_,
		_w2412_
	);
	LUT2 #(
		.INIT('h9)
	) name2387 (
		_w2392_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h6)
	) name2388 (
		_w2387_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h4)
	) name2389 (
		_w2382_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h9)
	) name2390 (
		_w2382_,
		_w2414_,
		_w2416_
	);
	LUT4 #(
		.INIT('h7100)
	) name2391 (
		_w2325_,
		_w2326_,
		_w2362_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2392 (
		_w2325_,
		_w2363_,
		_w2364_,
		_w2416_,
		_w2418_
	);
	LUT4 #(
		.INIT('h0400)
	) name2393 (
		_w252_,
		_w172_,
		_w78_,
		_w84_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name2394 (
		_w1234_,
		_w1149_,
		_w1255_,
		_w2420_
	);
	LUT4 #(
		.INIT('h8000)
	) name2395 (
		_w1316_,
		_w2082_,
		_w2420_,
		_w2419_,
		_w2421_
	);
	LUT4 #(
		.INIT('h1000)
	) name2396 (
		_w107_,
		_w311_,
		_w530_,
		_w1786_,
		_w2422_
	);
	LUT4 #(
		.INIT('h27ff)
	) name2397 (
		_w46_,
		_w76_,
		_w59_,
		_w70_,
		_w2423_
	);
	LUT3 #(
		.INIT('h10)
	) name2398 (
		_w168_,
		_w157_,
		_w2423_,
		_w2424_
	);
	LUT3 #(
		.INIT('h80)
	) name2399 (
		_w1344_,
		_w2424_,
		_w2422_,
		_w2425_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		_w2421_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		_w2022_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h4)
	) name2402 (
		_w2418_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h2)
	) name2403 (
		_w2418_,
		_w2427_,
		_w2429_
	);
	LUT2 #(
		.INIT('h9)
	) name2404 (
		_w2418_,
		_w2427_,
		_w2430_
	);
	LUT2 #(
		.INIT('h9)
	) name2405 (
		_w2381_,
		_w2430_,
		_w2431_
	);
	LUT4 #(
		.INIT('h8008)
	) name2406 (
		_w2321_,
		_w2377_,
		_w2381_,
		_w2430_,
		_w2432_
	);
	LUT4 #(
		.INIT('h7887)
	) name2407 (
		_w2321_,
		_w2377_,
		_w2381_,
		_w2430_,
		_w2433_
	);
	LUT3 #(
		.INIT('h90)
	) name2408 (
		_w2321_,
		_w2377_,
		_w2379_,
		_w2434_
	);
	LUT4 #(
		.INIT('h1455)
	) name2409 (
		_w2076_,
		_w2321_,
		_w2377_,
		_w2379_,
		_w2435_
	);
	LUT2 #(
		.INIT('h6)
	) name2410 (
		_w2433_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h45)
	) name2411 (
		_w2385_,
		_w2386_,
		_w2413_,
		_w2437_
	);
	LUT3 #(
		.INIT('h32)
	) name2412 (
		_w2392_,
		_w2410_,
		_w2411_,
		_w2438_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2413 (
		_w1526_,
		_w1951_,
		_w1953_,
		_w2088_,
		_w2439_
	);
	LUT4 #(
		.INIT('h802a)
	) name2414 (
		_w1528_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		_w1531_,
		_w1806_,
		_w2441_
	);
	LUT3 #(
		.INIT('h82)
	) name2416 (
		_w1530_,
		_w1805_,
		_w1949_,
		_w2442_
	);
	LUT3 #(
		.INIT('h01)
	) name2417 (
		_w2440_,
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT3 #(
		.INIT('h9a)
	) name2418 (
		_w581_,
		_w2439_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('h31)
	) name2419 (
		_w2398_,
		_w2407_,
		_w2408_,
		_w2445_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2420 (
		_w1460_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w2446_
	);
	LUT4 #(
		.INIT('h802a)
	) name2421 (
		_w1462_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2447_
	);
	LUT2 #(
		.INIT('h2)
	) name2422 (
		_w1464_,
		_w1741_,
		_w2448_
	);
	LUT3 #(
		.INIT('h82)
	) name2423 (
		_w1466_,
		_w1739_,
		_w1785_,
		_w2449_
	);
	LUT3 #(
		.INIT('h01)
	) name2424 (
		_w2447_,
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('h32)
	) name2425 (
		_w2403_,
		_w2404_,
		_w2405_,
		_w2451_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2426 (
		_w1401_,
		_w1437_,
		_w1448_,
		_w1475_,
		_w2452_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2427 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1479_,
		_w2453_
	);
	LUT3 #(
		.INIT('h90)
	) name2428 (
		_w1377_,
		_w1379_,
		_w1514_,
		_w2454_
	);
	LUT3 #(
		.INIT('h07)
	) name2429 (
		_w1400_,
		_w1477_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h0154)
	) name2431 (
		_w424_,
		_w1213_,
		_w1375_,
		_w1376_,
		_w2457_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		_w30_,
		_w33_,
		_w2458_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		_w30_,
		_w33_,
		_w2459_
	);
	LUT2 #(
		.INIT('h6)
	) name2434 (
		_w30_,
		_w33_,
		_w2460_
	);
	LUT2 #(
		.INIT('h6)
	) name2435 (
		_w2457_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2436 (
		_w424_,
		_w2452_,
		_w2456_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('h0065)
	) name2437 (
		_w424_,
		_w2452_,
		_w2456_,
		_w2461_,
		_w2463_
	);
	LUT4 #(
		.INIT('h659a)
	) name2438 (
		_w424_,
		_w2452_,
		_w2456_,
		_w2461_,
		_w2464_
	);
	LUT2 #(
		.INIT('h9)
	) name2439 (
		_w2451_,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2440 (
		_w366_,
		_w2446_,
		_w2450_,
		_w2465_,
		_w2466_
	);
	LUT4 #(
		.INIT('h0065)
	) name2441 (
		_w366_,
		_w2446_,
		_w2450_,
		_w2465_,
		_w2467_
	);
	LUT4 #(
		.INIT('h659a)
	) name2442 (
		_w366_,
		_w2446_,
		_w2450_,
		_w2465_,
		_w2468_
	);
	LUT2 #(
		.INIT('h9)
	) name2443 (
		_w2445_,
		_w2468_,
		_w2469_
	);
	LUT3 #(
		.INIT('h69)
	) name2444 (
		_w2438_,
		_w2444_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w2437_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h2)
	) name2446 (
		_w2437_,
		_w2470_,
		_w2472_
	);
	LUT2 #(
		.INIT('h9)
	) name2447 (
		_w2437_,
		_w2470_,
		_w2473_
	);
	LUT4 #(
		.INIT('h0001)
	) name2448 (
		_w339_,
		_w156_,
		_w306_,
		_w184_,
		_w2474_
	);
	LUT4 #(
		.INIT('h135f)
	) name2449 (
		_w206_,
		_w54_,
		_w96_,
		_w68_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		_w621_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h135f)
	) name2451 (
		_w88_,
		_w106_,
		_w125_,
		_w116_,
		_w2477_
	);
	LUT4 #(
		.INIT('h4000)
	) name2452 (
		_w197_,
		_w240_,
		_w1318_,
		_w2477_,
		_w2478_
	);
	LUT3 #(
		.INIT('h80)
	) name2453 (
		_w2474_,
		_w2476_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w2421_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		_w1217_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h001e)
	) name2456 (
		_w2415_,
		_w2417_,
		_w2473_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2457 (
		_w2415_,
		_w2417_,
		_w2473_,
		_w2481_,
		_w2483_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2458 (
		_w2381_,
		_w2418_,
		_w2427_,
		_w2483_,
		_w2484_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name2459 (
		_w2381_,
		_w2428_,
		_w2429_,
		_w2483_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		_w2432_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h6)
	) name2461 (
		_w2432_,
		_w2485_,
		_w2487_
	);
	LUT3 #(
		.INIT('h45)
	) name2462 (
		_w2076_,
		_w2433_,
		_w2434_,
		_w2488_
	);
	LUT2 #(
		.INIT('h6)
	) name2463 (
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2464 (
		_w2415_,
		_w2417_,
		_w2471_,
		_w2472_,
		_w2490_
	);
	LUT3 #(
		.INIT('h2b)
	) name2465 (
		_w2438_,
		_w2444_,
		_w2469_,
		_w2491_
	);
	LUT3 #(
		.INIT('h82)
	) name2466 (
		_w1531_,
		_w1805_,
		_w1949_,
		_w2492_
	);
	LUT4 #(
		.INIT('h802a)
	) name2467 (
		_w1530_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('h5700)
	) name2469 (
		_w1526_,
		_w2151_,
		_w2152_,
		_w2494_,
		_w2495_
	);
	LUT3 #(
		.INIT('h32)
	) name2470 (
		_w2445_,
		_w2466_,
		_w2467_,
		_w2496_
	);
	LUT3 #(
		.INIT('h82)
	) name2471 (
		_w1464_,
		_w1739_,
		_w1785_,
		_w2497_
	);
	LUT4 #(
		.INIT('h802a)
	) name2472 (
		_w1466_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2498_
	);
	LUT4 #(
		.INIT('h000d)
	) name2473 (
		_w1462_,
		_w1806_,
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2474 (
		_w1460_,
		_w1798_,
		_w1809_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h32)
	) name2475 (
		_w2451_,
		_w2462_,
		_w2463_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		_w1400_,
		_w1514_,
		_w2502_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2477 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1477_,
		_w2503_
	);
	LUT4 #(
		.INIT('h000d)
	) name2478 (
		_w1479_,
		_w1741_,
		_w2502_,
		_w2503_,
		_w2504_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2479 (
		_w1475_,
		_w1720_,
		_w1744_,
		_w2504_,
		_w2505_
	);
	LUT3 #(
		.INIT('h41)
	) name2480 (
		_w424_,
		_w1377_,
		_w1379_,
		_w2506_
	);
	LUT3 #(
		.INIT('h31)
	) name2481 (
		_w2457_,
		_w2458_,
		_w2459_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w2506_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		_w2506_,
		_w2507_,
		_w2509_
	);
	LUT2 #(
		.INIT('h6)
	) name2484 (
		_w2506_,
		_w2507_,
		_w2510_
	);
	LUT3 #(
		.INIT('h96)
	) name2485 (
		_w424_,
		_w2505_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h4)
	) name2486 (
		_w2501_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h2)
	) name2487 (
		_w2501_,
		_w2511_,
		_w2513_
	);
	LUT2 #(
		.INIT('h9)
	) name2488 (
		_w2501_,
		_w2511_,
		_w2514_
	);
	LUT3 #(
		.INIT('h96)
	) name2489 (
		_w366_,
		_w2500_,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name2490 (
		_w2496_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		_w2496_,
		_w2515_,
		_w2517_
	);
	LUT2 #(
		.INIT('h9)
	) name2492 (
		_w2496_,
		_w2515_,
		_w2518_
	);
	LUT3 #(
		.INIT('h96)
	) name2493 (
		_w581_,
		_w2495_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w2491_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name2495 (
		_w2491_,
		_w2519_,
		_w2521_
	);
	LUT2 #(
		.INIT('h9)
	) name2496 (
		_w2491_,
		_w2519_,
		_w2522_
	);
	LUT4 #(
		.INIT('h0777)
	) name2497 (
		_w121_,
		_w59_,
		_w85_,
		_w102_,
		_w2523_
	);
	LUT2 #(
		.INIT('h4)
	) name2498 (
		_w221_,
		_w2523_,
		_w2524_
	);
	LUT4 #(
		.INIT('h1000)
	) name2499 (
		_w347_,
		_w253_,
		_w199_,
		_w373_,
		_w2525_
	);
	LUT3 #(
		.INIT('h80)
	) name2500 (
		_w1172_,
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		_w188_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h153f)
	) name2502 (
		_w106_,
		_w59_,
		_w71_,
		_w100_,
		_w2528_
	);
	LUT4 #(
		.INIT('h37bf)
	) name2503 (
		_w46_,
		_w53_,
		_w82_,
		_w98_,
		_w2529_
	);
	LUT4 #(
		.INIT('h4000)
	) name2504 (
		_w379_,
		_w1261_,
		_w2529_,
		_w2528_,
		_w2530_
	);
	LUT4 #(
		.INIT('h8000)
	) name2505 (
		_w520_,
		_w524_,
		_w1264_,
		_w2530_,
		_w2531_
	);
	LUT4 #(
		.INIT('h8000)
	) name2506 (
		_w188_,
		_w2057_,
		_w2526_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('h09)
	) name2507 (
		_w2490_,
		_w2522_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h96)
	) name2508 (
		_w2490_,
		_w2522_,
		_w2532_,
		_w2534_
	);
	LUT3 #(
		.INIT('h1e)
	) name2509 (
		_w2482_,
		_w2484_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		_w2486_,
		_w2535_,
		_w2536_
	);
	LUT4 #(
		.INIT('h8010)
	) name2511 (
		_w2378_,
		_w2431_,
		_w2434_,
		_w2485_,
		_w2537_
	);
	LUT4 #(
		.INIT('h3c69)
	) name2512 (
		_w2076_,
		_w2486_,
		_w2535_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('h010f)
	) name2513 (
		_w2482_,
		_w2484_,
		_w2533_,
		_w2534_,
		_w2539_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2514 (
		_w581_,
		_w2495_,
		_w2516_,
		_w2517_,
		_w2540_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2515 (
		_w366_,
		_w2500_,
		_w2512_,
		_w2513_,
		_w2541_
	);
	LUT4 #(
		.INIT('h1151)
	) name2516 (
		_w1531_,
		_w1526_,
		_w1950_,
		_w1953_,
		_w2542_
	);
	LUT4 #(
		.INIT('h0509)
	) name2517 (
		_w581_,
		_w2090_,
		_w2541_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('ha060)
	) name2518 (
		_w581_,
		_w2090_,
		_w2541_,
		_w2542_,
		_w2544_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2519 (
		_w581_,
		_w2090_,
		_w2541_,
		_w2542_,
		_w2545_
	);
	LUT3 #(
		.INIT('h82)
	) name2520 (
		_w1462_,
		_w1805_,
		_w1949_,
		_w2546_
	);
	LUT4 #(
		.INIT('h802a)
	) name2521 (
		_w1464_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2547_
	);
	LUT3 #(
		.INIT('h0d)
	) name2522 (
		_w1466_,
		_w1806_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h4)
	) name2523 (
		_w2546_,
		_w2548_,
		_w2549_
	);
	LUT4 #(
		.INIT('h95aa)
	) name2524 (
		_w366_,
		_w1460_,
		_w1954_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2525 (
		_w424_,
		_w2505_,
		_w2508_,
		_w2509_,
		_w2551_
	);
	LUT3 #(
		.INIT('h82)
	) name2526 (
		_w1479_,
		_w1739_,
		_w1785_,
		_w2552_
	);
	LUT4 #(
		.INIT('h1e00)
	) name2527 (
		_w1396_,
		_w1398_,
		_w1445_,
		_w1514_,
		_w2553_
	);
	LUT3 #(
		.INIT('h0d)
	) name2528 (
		_w1477_,
		_w1741_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h4)
	) name2529 (
		_w2552_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h6a55)
	) name2530 (
		_w424_,
		_w1475_,
		_w1827_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		_w424_,
		_w1436_,
		_w2557_
	);
	LUT3 #(
		.INIT('h14)
	) name2532 (
		_w2551_,
		_w2556_,
		_w2557_,
		_w2558_
	);
	LUT3 #(
		.INIT('h82)
	) name2533 (
		_w2551_,
		_w2556_,
		_w2557_,
		_w2559_
	);
	LUT3 #(
		.INIT('h69)
	) name2534 (
		_w2551_,
		_w2556_,
		_w2557_,
		_w2560_
	);
	LUT2 #(
		.INIT('h6)
	) name2535 (
		_w2550_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h6)
	) name2536 (
		_w2545_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name2537 (
		_w2540_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h9)
	) name2538 (
		_w2540_,
		_w2562_,
		_w2564_
	);
	LUT4 #(
		.INIT('h7100)
	) name2539 (
		_w2490_,
		_w2491_,
		_w2519_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2540 (
		_w2490_,
		_w2520_,
		_w2521_,
		_w2564_,
		_w2566_
	);
	LUT3 #(
		.INIT('h1f)
	) name2541 (
		_w76_,
		_w113_,
		_w77_,
		_w2567_
	);
	LUT4 #(
		.INIT('h153f)
	) name2542 (
		_w85_,
		_w62_,
		_w71_,
		_w72_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('h1000)
	) name2544 (
		_w107_,
		_w178_,
		_w240_,
		_w1786_,
		_w2570_
	);
	LUT4 #(
		.INIT('h8000)
	) name2545 (
		_w269_,
		_w2141_,
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('h8000)
	) name2546 (
		_w1312_,
		_w1320_,
		_w2025_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h4)
	) name2547 (
		_w2566_,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h2)
	) name2548 (
		_w2566_,
		_w2572_,
		_w2574_
	);
	LUT2 #(
		.INIT('h9)
	) name2549 (
		_w2566_,
		_w2572_,
		_w2575_
	);
	LUT2 #(
		.INIT('h9)
	) name2550 (
		_w2539_,
		_w2575_,
		_w2576_
	);
	LUT4 #(
		.INIT('h8008)
	) name2551 (
		_w2486_,
		_w2535_,
		_w2539_,
		_w2575_,
		_w2577_
	);
	LUT4 #(
		.INIT('h7887)
	) name2552 (
		_w2486_,
		_w2535_,
		_w2539_,
		_w2575_,
		_w2578_
	);
	LUT3 #(
		.INIT('h90)
	) name2553 (
		_w2486_,
		_w2535_,
		_w2537_,
		_w2579_
	);
	LUT4 #(
		.INIT('h1455)
	) name2554 (
		_w2076_,
		_w2486_,
		_w2535_,
		_w2537_,
		_w2580_
	);
	LUT2 #(
		.INIT('h6)
	) name2555 (
		_w2578_,
		_w2580_,
		_w2581_
	);
	LUT3 #(
		.INIT('h45)
	) name2556 (
		_w2543_,
		_w2544_,
		_w2561_,
		_w2582_
	);
	LUT3 #(
		.INIT('h31)
	) name2557 (
		_w2550_,
		_w2558_,
		_w2559_,
		_w2583_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2558 (
		_w1460_,
		_w1951_,
		_w1953_,
		_w2088_,
		_w2584_
	);
	LUT4 #(
		.INIT('h802a)
	) name2559 (
		_w1462_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2585_
	);
	LUT2 #(
		.INIT('h2)
	) name2560 (
		_w1464_,
		_w1806_,
		_w2586_
	);
	LUT3 #(
		.INIT('h82)
	) name2561 (
		_w1466_,
		_w1805_,
		_w1949_,
		_w2587_
	);
	LUT3 #(
		.INIT('h01)
	) name2562 (
		_w2585_,
		_w2586_,
		_w2587_,
		_w2588_
	);
	LUT3 #(
		.INIT('h9a)
	) name2563 (
		_w366_,
		_w2584_,
		_w2588_,
		_w2589_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2564 (
		_w1475_,
		_w1793_,
		_w1795_,
		_w1797_,
		_w2590_
	);
	LUT4 #(
		.INIT('h802a)
	) name2565 (
		_w1479_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2591_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		_w1514_,
		_w1741_,
		_w2592_
	);
	LUT3 #(
		.INIT('h82)
	) name2567 (
		_w1477_,
		_w1739_,
		_w1785_,
		_w2593_
	);
	LUT3 #(
		.INIT('h01)
	) name2568 (
		_w2591_,
		_w2592_,
		_w2593_,
		_w2594_
	);
	LUT3 #(
		.INIT('h65)
	) name2569 (
		_w424_,
		_w2590_,
		_w2594_,
		_w2595_
	);
	LUT4 #(
		.INIT('h0154)
	) name2570 (
		_w424_,
		_w1396_,
		_w1398_,
		_w1445_,
		_w2596_
	);
	LUT3 #(
		.INIT('h69)
	) name2571 (
		_w581_,
		_w2506_,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('h14)
	) name2572 (
		_w424_,
		_w1377_,
		_w1379_,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		_w1400_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2574 (
		_w2556_,
		_w2557_,
		_w2597_,
		_w2599_,
		_w2600_
	);
	LUT4 #(
		.INIT('h00e0)
	) name2575 (
		_w2556_,
		_w2557_,
		_w2597_,
		_w2599_,
		_w2601_
	);
	LUT4 #(
		.INIT('hf01e)
	) name2576 (
		_w2556_,
		_w2557_,
		_w2597_,
		_w2599_,
		_w2602_
	);
	LUT2 #(
		.INIT('h9)
	) name2577 (
		_w2595_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('h69)
	) name2578 (
		_w2583_,
		_w2589_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h4)
	) name2579 (
		_w2582_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w2582_,
		_w2604_,
		_w2606_
	);
	LUT2 #(
		.INIT('h9)
	) name2581 (
		_w2582_,
		_w2604_,
		_w2607_
	);
	LUT4 #(
		.INIT('h1000)
	) name2582 (
		_w238_,
		_w271_,
		_w212_,
		_w1786_,
		_w2608_
	);
	LUT4 #(
		.INIT('h0777)
	) name2583 (
		_w54_,
		_w79_,
		_w77_,
		_w62_,
		_w2609_
	);
	LUT4 #(
		.INIT('h1000)
	) name2584 (
		_w115_,
		_w158_,
		_w291_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h8000)
	) name2585 (
		_w519_,
		_w1732_,
		_w2608_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name2586 (
		_w447_,
		_w2611_,
		_w2612_
	);
	LUT3 #(
		.INIT('h80)
	) name2587 (
		_w623_,
		_w626_,
		_w2063_,
		_w2613_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT4 #(
		.INIT('h001e)
	) name2589 (
		_w2563_,
		_w2565_,
		_w2607_,
		_w2614_,
		_w2615_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2590 (
		_w2563_,
		_w2565_,
		_w2607_,
		_w2614_,
		_w2616_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2591 (
		_w2539_,
		_w2566_,
		_w2572_,
		_w2616_,
		_w2617_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name2592 (
		_w2539_,
		_w2573_,
		_w2574_,
		_w2616_,
		_w2618_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		_w2577_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h6)
	) name2594 (
		_w2577_,
		_w2618_,
		_w2620_
	);
	LUT3 #(
		.INIT('h45)
	) name2595 (
		_w2076_,
		_w2578_,
		_w2579_,
		_w2621_
	);
	LUT2 #(
		.INIT('h6)
	) name2596 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2597 (
		_w2563_,
		_w2565_,
		_w2605_,
		_w2606_,
		_w2623_
	);
	LUT3 #(
		.INIT('h2b)
	) name2598 (
		_w2583_,
		_w2589_,
		_w2603_,
		_w2624_
	);
	LUT3 #(
		.INIT('h82)
	) name2599 (
		_w1464_,
		_w1805_,
		_w1949_,
		_w2625_
	);
	LUT4 #(
		.INIT('h802a)
	) name2600 (
		_w1466_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name2601 (
		_w2625_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('h5700)
	) name2602 (
		_w1460_,
		_w2151_,
		_w2152_,
		_w2627_,
		_w2628_
	);
	LUT3 #(
		.INIT('h82)
	) name2603 (
		_w1514_,
		_w1739_,
		_w1785_,
		_w2629_
	);
	LUT4 #(
		.INIT('h802a)
	) name2604 (
		_w1477_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2630_
	);
	LUT4 #(
		.INIT('h000d)
	) name2605 (
		_w1479_,
		_w1806_,
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2606 (
		_w1475_,
		_w1798_,
		_w1809_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w424_,
		_w1741_,
		_w2633_
	);
	LUT3 #(
		.INIT('he8)
	) name2608 (
		_w581_,
		_w2506_,
		_w2596_,
		_w2634_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		_w2633_,
		_w2634_,
		_w2636_
	);
	LUT2 #(
		.INIT('h9)
	) name2611 (
		_w2633_,
		_w2634_,
		_w2637_
	);
	LUT3 #(
		.INIT('h96)
	) name2612 (
		_w424_,
		_w2632_,
		_w2637_,
		_w2638_
	);
	LUT3 #(
		.INIT('h32)
	) name2613 (
		_w2595_,
		_w2600_,
		_w2601_,
		_w2639_
	);
	LUT2 #(
		.INIT('h2)
	) name2614 (
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w2638_,
		_w2639_,
		_w2641_
	);
	LUT2 #(
		.INIT('h9)
	) name2616 (
		_w2638_,
		_w2639_,
		_w2642_
	);
	LUT3 #(
		.INIT('h96)
	) name2617 (
		_w366_,
		_w2628_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h4)
	) name2618 (
		_w2624_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		_w2624_,
		_w2643_,
		_w2645_
	);
	LUT2 #(
		.INIT('h9)
	) name2620 (
		_w2624_,
		_w2643_,
		_w2646_
	);
	LUT4 #(
		.INIT('h1000)
	) name2621 (
		_w252_,
		_w244_,
		_w528_,
		_w547_,
		_w2647_
	);
	LUT3 #(
		.INIT('h80)
	) name2622 (
		_w378_,
		_w409_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		_w1943_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name2624 (
		_w441_,
		_w2649_,
		_w2650_
	);
	LUT3 #(
		.INIT('h09)
	) name2625 (
		_w2623_,
		_w2646_,
		_w2650_,
		_w2651_
	);
	LUT3 #(
		.INIT('h96)
	) name2626 (
		_w2623_,
		_w2646_,
		_w2650_,
		_w2652_
	);
	LUT3 #(
		.INIT('h1e)
	) name2627 (
		_w2615_,
		_w2617_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		_w2619_,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h8010)
	) name2629 (
		_w2536_,
		_w2576_,
		_w2579_,
		_w2618_,
		_w2655_
	);
	LUT4 #(
		.INIT('h3c69)
	) name2630 (
		_w2076_,
		_w2619_,
		_w2653_,
		_w2655_,
		_w2656_
	);
	LUT4 #(
		.INIT('h010f)
	) name2631 (
		_w2615_,
		_w2617_,
		_w2651_,
		_w2652_,
		_w2657_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2632 (
		_w366_,
		_w2628_,
		_w2640_,
		_w2641_,
		_w2658_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2633 (
		_w424_,
		_w2632_,
		_w2635_,
		_w2636_,
		_w2659_
	);
	LUT4 #(
		.INIT('h4010)
	) name2634 (
		_w424_,
		_w1739_,
		_w1741_,
		_w1785_,
		_w2660_
	);
	LUT4 #(
		.INIT('h0140)
	) name2635 (
		_w424_,
		_w1446_,
		_w1738_,
		_w1785_,
		_w2661_
	);
	LUT4 #(
		.INIT('hefba)
	) name2636 (
		_w424_,
		_w1739_,
		_w1740_,
		_w1785_,
		_w2662_
	);
	LUT2 #(
		.INIT('h9)
	) name2637 (
		_w2659_,
		_w2662_,
		_w2663_
	);
	LUT3 #(
		.INIT('h82)
	) name2638 (
		_w1479_,
		_w1805_,
		_w1949_,
		_w2664_
	);
	LUT4 #(
		.INIT('h802a)
	) name2639 (
		_w1514_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2665_
	);
	LUT3 #(
		.INIT('h0d)
	) name2640 (
		_w1477_,
		_w1806_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h4)
	) name2641 (
		_w2664_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h6a55)
	) name2642 (
		_w424_,
		_w1475_,
		_w1954_,
		_w2667_,
		_w2668_
	);
	LUT4 #(
		.INIT('h1151)
	) name2643 (
		_w1464_,
		_w1460_,
		_w1950_,
		_w1953_,
		_w2669_
	);
	LUT4 #(
		.INIT('h0509)
	) name2644 (
		_w366_,
		_w2090_,
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('ha060)
	) name2645 (
		_w366_,
		_w2090_,
		_w2668_,
		_w2669_,
		_w2671_
	);
	LUT4 #(
		.INIT('h5a96)
	) name2646 (
		_w366_,
		_w2090_,
		_w2668_,
		_w2669_,
		_w2672_
	);
	LUT2 #(
		.INIT('h6)
	) name2647 (
		_w2663_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w2658_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h9)
	) name2649 (
		_w2658_,
		_w2673_,
		_w2675_
	);
	LUT4 #(
		.INIT('h7100)
	) name2650 (
		_w2623_,
		_w2624_,
		_w2643_,
		_w2675_,
		_w2676_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2651 (
		_w2623_,
		_w2644_,
		_w2645_,
		_w2675_,
		_w2677_
	);
	LUT4 #(
		.INIT('h135f)
	) name2652 (
		_w206_,
		_w85_,
		_w77_,
		_w98_,
		_w2678_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name2653 (
		_w46_,
		_w53_,
		_w68_,
		_w100_,
		_w2679_
	);
	LUT3 #(
		.INIT('h40)
	) name2654 (
		_w140_,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h135f)
	) name2655 (
		_w121_,
		_w95_,
		_w59_,
		_w125_,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		_w1283_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('h8000)
	) name2657 (
		_w565_,
		_w2197_,
		_w2198_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('h8000)
	) name2658 (
		_w1276_,
		_w1201_,
		_w2680_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h4)
	) name2659 (
		_w2677_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h2)
	) name2660 (
		_w2677_,
		_w2684_,
		_w2686_
	);
	LUT2 #(
		.INIT('h9)
	) name2661 (
		_w2677_,
		_w2684_,
		_w2687_
	);
	LUT2 #(
		.INIT('h9)
	) name2662 (
		_w2657_,
		_w2687_,
		_w2688_
	);
	LUT4 #(
		.INIT('h8008)
	) name2663 (
		_w2619_,
		_w2653_,
		_w2657_,
		_w2687_,
		_w2689_
	);
	LUT4 #(
		.INIT('h7887)
	) name2664 (
		_w2619_,
		_w2653_,
		_w2657_,
		_w2687_,
		_w2690_
	);
	LUT3 #(
		.INIT('h90)
	) name2665 (
		_w2619_,
		_w2653_,
		_w2655_,
		_w2691_
	);
	LUT4 #(
		.INIT('h1455)
	) name2666 (
		_w2076_,
		_w2619_,
		_w2653_,
		_w2655_,
		_w2692_
	);
	LUT2 #(
		.INIT('h6)
	) name2667 (
		_w2690_,
		_w2692_,
		_w2693_
	);
	LUT3 #(
		.INIT('h31)
	) name2668 (
		_w2663_,
		_w2670_,
		_w2671_,
		_w2694_
	);
	LUT3 #(
		.INIT('h0e)
	) name2669 (
		_w2659_,
		_w2660_,
		_w2661_,
		_w2695_
	);
	LUT4 #(
		.INIT('h02a8)
	) name2670 (
		_w1475_,
		_w1951_,
		_w1953_,
		_w2088_,
		_w2696_
	);
	LUT4 #(
		.INIT('h802a)
	) name2671 (
		_w1479_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2697_
	);
	LUT2 #(
		.INIT('h2)
	) name2672 (
		_w1514_,
		_w1806_,
		_w2698_
	);
	LUT3 #(
		.INIT('h82)
	) name2673 (
		_w1477_,
		_w1805_,
		_w1949_,
		_w2699_
	);
	LUT3 #(
		.INIT('h01)
	) name2674 (
		_w2697_,
		_w2698_,
		_w2699_,
		_w2700_
	);
	LUT4 #(
		.INIT('h2002)
	) name2675 (
		_w366_,
		_w424_,
		_w1739_,
		_w1785_,
		_w2701_
	);
	LUT4 #(
		.INIT('h4554)
	) name2676 (
		_w366_,
		_w424_,
		_w1739_,
		_w1785_,
		_w2702_
	);
	LUT4 #(
		.INIT('h9aa9)
	) name2677 (
		_w366_,
		_w424_,
		_w1739_,
		_w1785_,
		_w2703_
	);
	LUT4 #(
		.INIT('h4015)
	) name2678 (
		_w424_,
		_w1739_,
		_w1785_,
		_w1791_,
		_w2704_
	);
	LUT2 #(
		.INIT('h6)
	) name2679 (
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2680 (
		_w424_,
		_w2696_,
		_w2700_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h0065)
	) name2681 (
		_w424_,
		_w2696_,
		_w2700_,
		_w2705_,
		_w2707_
	);
	LUT4 #(
		.INIT('h659a)
	) name2682 (
		_w424_,
		_w2696_,
		_w2700_,
		_w2705_,
		_w2708_
	);
	LUT2 #(
		.INIT('h9)
	) name2683 (
		_w2695_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h4)
	) name2684 (
		_w2694_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name2685 (
		_w2694_,
		_w2709_,
		_w2711_
	);
	LUT2 #(
		.INIT('h9)
	) name2686 (
		_w2694_,
		_w2709_,
		_w2712_
	);
	LUT4 #(
		.INIT('h0100)
	) name2687 (
		_w110_,
		_w207_,
		_w144_,
		_w575_,
		_w2713_
	);
	LUT3 #(
		.INIT('h04)
	) name2688 (
		_w64_,
		_w172_,
		_w182_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		_w509_,
		_w658_,
		_w2715_
	);
	LUT4 #(
		.INIT('hcdff)
	) name2690 (
		_w87_,
		_w46_,
		_w53_,
		_w82_,
		_w2716_
	);
	LUT4 #(
		.INIT('h4000)
	) name2691 (
		_w111_,
		_w814_,
		_w2138_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('h8000)
	) name2692 (
		_w2713_,
		_w2714_,
		_w2715_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h8000)
	) name2693 (
		_w642_,
		_w1167_,
		_w2039_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h001e)
	) name2694 (
		_w2674_,
		_w2676_,
		_w2712_,
		_w2719_,
		_w2720_
	);
	LUT4 #(
		.INIT('h1ee1)
	) name2695 (
		_w2674_,
		_w2676_,
		_w2712_,
		_w2719_,
		_w2721_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2696 (
		_w2657_,
		_w2677_,
		_w2684_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h0ef1)
	) name2697 (
		_w2657_,
		_w2685_,
		_w2686_,
		_w2721_,
		_w2723_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		_w2689_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h6)
	) name2699 (
		_w2689_,
		_w2723_,
		_w2725_
	);
	LUT3 #(
		.INIT('h45)
	) name2700 (
		_w2076_,
		_w2690_,
		_w2691_,
		_w2726_
	);
	LUT2 #(
		.INIT('h6)
	) name2701 (
		_w2725_,
		_w2726_,
		_w2727_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2702 (
		_w2674_,
		_w2676_,
		_w2710_,
		_w2711_,
		_w2728_
	);
	LUT3 #(
		.INIT('h32)
	) name2703 (
		_w2695_,
		_w2706_,
		_w2707_,
		_w2729_
	);
	LUT3 #(
		.INIT('h82)
	) name2704 (
		_w1514_,
		_w1805_,
		_w1949_,
		_w2730_
	);
	LUT4 #(
		.INIT('h802a)
	) name2705 (
		_w1477_,
		_w1805_,
		_w1949_,
		_w2087_,
		_w2731_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w2730_,
		_w2731_,
		_w2732_
	);
	LUT4 #(
		.INIT('h5700)
	) name2707 (
		_w1475_,
		_w2151_,
		_w2152_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w424_,
		_w1806_,
		_w2734_
	);
	LUT3 #(
		.INIT('h45)
	) name2709 (
		_w2701_,
		_w2702_,
		_w2704_,
		_w2735_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		_w2734_,
		_w2735_,
		_w2737_
	);
	LUT2 #(
		.INIT('h6)
	) name2712 (
		_w2734_,
		_w2735_,
		_w2738_
	);
	LUT3 #(
		.INIT('h96)
	) name2713 (
		_w424_,
		_w2733_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w2729_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h2)
	) name2715 (
		_w2729_,
		_w2739_,
		_w2741_
	);
	LUT2 #(
		.INIT('h9)
	) name2716 (
		_w2729_,
		_w2739_,
		_w2742_
	);
	LUT4 #(
		.INIT('h8000)
	) name2717 (
		_w383_,
		_w1283_,
		_w1323_,
		_w1786_,
		_w2743_
	);
	LUT4 #(
		.INIT('h37bf)
	) name2718 (
		_w46_,
		_w95_,
		_w91_,
		_w72_,
		_w2744_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w284_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name2720 (
		_w46_,
		_w53_,
		_w82_,
		_w62_,
		_w2746_
	);
	LUT3 #(
		.INIT('h10)
	) name2721 (
		_w225_,
		_w145_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h8000)
	) name2722 (
		_w511_,
		_w2745_,
		_w2747_,
		_w2743_,
		_w2748_
	);
	LUT4 #(
		.INIT('h8000)
	) name2723 (
		_w524_,
		_w527_,
		_w823_,
		_w825_,
		_w2749_
	);
	LUT3 #(
		.INIT('h80)
	) name2724 (
		_w1174_,
		_w2748_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('h09)
	) name2725 (
		_w2728_,
		_w2742_,
		_w2750_,
		_w2751_
	);
	LUT3 #(
		.INIT('h96)
	) name2726 (
		_w2728_,
		_w2742_,
		_w2750_,
		_w2752_
	);
	LUT3 #(
		.INIT('h1e)
	) name2727 (
		_w2720_,
		_w2722_,
		_w2752_,
		_w2753_
	);
	LUT4 #(
		.INIT('h8010)
	) name2728 (
		_w2654_,
		_w2688_,
		_w2691_,
		_w2723_,
		_w2754_
	);
	LUT4 #(
		.INIT('h3c69)
	) name2729 (
		_w2076_,
		_w2724_,
		_w2753_,
		_w2754_,
		_w2755_
	);
	LUT4 #(
		.INIT('h010f)
	) name2730 (
		_w2720_,
		_w2722_,
		_w2751_,
		_w2752_,
		_w2756_
	);
	LUT4 #(
		.INIT('h0f09)
	) name2731 (
		_w424_,
		_w2733_,
		_w2736_,
		_w2737_,
		_w2757_
	);
	LUT4 #(
		.INIT('h1131)
	) name2732 (
		_w1475_,
		_w1514_,
		_w1950_,
		_w1953_,
		_w2758_
	);
	LUT4 #(
		.INIT('h11a1)
	) name2733 (
		_w424_,
		_w1952_,
		_w2090_,
		_w2758_,
		_w2759_
	);
	LUT4 #(
		.INIT('hee1e)
	) name2734 (
		_w424_,
		_w1952_,
		_w2090_,
		_w2758_,
		_w2760_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w2757_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h9)
	) name2736 (
		_w2757_,
		_w2760_,
		_w2762_
	);
	LUT4 #(
		.INIT('h7100)
	) name2737 (
		_w2728_,
		_w2729_,
		_w2739_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('h32cd)
	) name2738 (
		_w2728_,
		_w2740_,
		_w2741_,
		_w2762_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name2739 (
		_w297_,
		_w1322_,
		_w2765_
	);
	LUT3 #(
		.INIT('h80)
	) name2740 (
		_w655_,
		_w661_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name2741 (
		_w46_,
		_w53_,
		_w59_,
		_w116_,
		_w2767_
	);
	LUT3 #(
		.INIT('h10)
	) name2742 (
		_w145_,
		_w78_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('h1000)
	) name2743 (
		_w386_,
		_w64_,
		_w530_,
		_w2058_,
		_w2769_
	);
	LUT3 #(
		.INIT('h80)
	) name2744 (
		_w2680_,
		_w2768_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('h8000)
	) name2745 (
		_w546_,
		_w647_,
		_w1285_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		_w2766_,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		_w2764_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h4)
	) name2748 (
		_w2764_,
		_w2772_,
		_w2774_
	);
	LUT2 #(
		.INIT('h9)
	) name2749 (
		_w2764_,
		_w2772_,
		_w2775_
	);
	LUT4 #(
		.INIT('h8008)
	) name2750 (
		_w2724_,
		_w2753_,
		_w2756_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('h7887)
	) name2751 (
		_w2724_,
		_w2753_,
		_w2756_,
		_w2775_,
		_w2777_
	);
	LUT3 #(
		.INIT('h90)
	) name2752 (
		_w2724_,
		_w2753_,
		_w2754_,
		_w2778_
	);
	LUT4 #(
		.INIT('h1455)
	) name2753 (
		_w2076_,
		_w2724_,
		_w2753_,
		_w2754_,
		_w2779_
	);
	LUT2 #(
		.INIT('h6)
	) name2754 (
		_w2777_,
		_w2779_,
		_w2780_
	);
	LUT3 #(
		.INIT('h32)
	) name2755 (
		_w2756_,
		_w2773_,
		_w2774_,
		_w2781_
	);
	LUT3 #(
		.INIT('h01)
	) name2756 (
		_w348_,
		_w257_,
		_w311_,
		_w2782_
	);
	LUT2 #(
		.INIT('h8)
	) name2757 (
		_w451_,
		_w291_,
		_w2783_
	);
	LUT3 #(
		.INIT('h80)
	) name2758 (
		_w1203_,
		_w2782_,
		_w2783_,
		_w2784_
	);
	LUT3 #(
		.INIT('h80)
	) name2759 (
		_w1305_,
		_w2012_,
		_w2713_,
		_w2785_
	);
	LUT3 #(
		.INIT('h80)
	) name2760 (
		_w2041_,
		_w2784_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		_w1233_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		_w424_,
		_w1949_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name2763 (
		_w1806_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w2759_,
		_w2789_,
		_w2790_
	);
	LUT4 #(
		.INIT('h1320)
	) name2765 (
		_w1805_,
		_w1806_,
		_w1949_,
		_w2087_,
		_w2791_
	);
	LUT3 #(
		.INIT('h51)
	) name2766 (
		_w424_,
		_w1806_,
		_w2087_,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name2767 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT4 #(
		.INIT('he11e)
	) name2768 (
		_w2761_,
		_w2763_,
		_w2790_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name2769 (
		_w2787_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h4)
	) name2770 (
		_w2787_,
		_w2794_,
		_w2796_
	);
	LUT2 #(
		.INIT('h9)
	) name2771 (
		_w2787_,
		_w2794_,
		_w2797_
	);
	LUT3 #(
		.INIT('h14)
	) name2772 (
		_w2776_,
		_w2781_,
		_w2797_,
		_w2798_
	);
	LUT3 #(
		.INIT('h82)
	) name2773 (
		_w2776_,
		_w2781_,
		_w2797_,
		_w2799_
	);
	LUT3 #(
		.INIT('h69)
	) name2774 (
		_w2776_,
		_w2781_,
		_w2797_,
		_w2800_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		_w2777_,
		_w2778_,
		_w2801_
	);
	LUT3 #(
		.INIT('h45)
	) name2776 (
		_w2076_,
		_w2777_,
		_w2778_,
		_w2802_
	);
	LUT2 #(
		.INIT('h6)
	) name2777 (
		_w2800_,
		_w2802_,
		_w2803_
	);
	LUT3 #(
		.INIT('h45)
	) name2778 (
		_w2076_,
		_w2800_,
		_w2801_,
		_w2804_
	);
	LUT4 #(
		.INIT('h135f)
	) name2779 (
		_w85_,
		_w68_,
		_w98_,
		_w71_,
		_w2805_
	);
	LUT3 #(
		.INIT('h10)
	) name2780 (
		_w238_,
		_w271_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h8)
	) name2781 (
		_w509_,
		_w544_,
		_w2807_
	);
	LUT4 #(
		.INIT('h57df)
	) name2782 (
		_w87_,
		_w46_,
		_w113_,
		_w100_,
		_w2808_
	);
	LUT4 #(
		.INIT('h1000)
	) name2783 (
		_w184_,
		_w300_,
		_w302_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('h8000)
	) name2784 (
		_w175_,
		_w2806_,
		_w2807_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('h8000)
	) name2785 (
		_w149_,
		_w167_,
		_w1731_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h0071)
	) name2786 (
		_w2781_,
		_w2787_,
		_w2794_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('h8e00)
	) name2787 (
		_w2781_,
		_w2787_,
		_w2794_,
		_w2811_,
		_w2813_
	);
	LUT4 #(
		.INIT('h31ce)
	) name2788 (
		_w2781_,
		_w2795_,
		_w2796_,
		_w2811_,
		_w2814_
	);
	LUT2 #(
		.INIT('h6)
	) name2789 (
		_w2799_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h6)
	) name2790 (
		_w2804_,
		_w2815_,
		_w2816_
	);
	LUT4 #(
		.INIT('hc020)
	) name2791 (
		_w2798_,
		_w2799_,
		_w2801_,
		_w2814_,
		_w2817_
	);
	LUT4 #(
		.INIT('h153f)
	) name2792 (
		_w85_,
		_w91_,
		_w77_,
		_w98_,
		_w2818_
	);
	LUT4 #(
		.INIT('h777f)
	) name2793 (
		_w46_,
		_w95_,
		_w102_,
		_w72_,
		_w2819_
	);
	LUT3 #(
		.INIT('h40)
	) name2794 (
		_w163_,
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT3 #(
		.INIT('h80)
	) name2795 (
		_w435_,
		_w503_,
		_w504_,
		_w2821_
	);
	LUT4 #(
		.INIT('h8000)
	) name2796 (
		_w636_,
		_w1162_,
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('h8000)
	) name2797 (
		_w191_,
		_w668_,
		_w2054_,
		_w2822_,
		_w2823_
	);
	LUT4 #(
		.INIT('h31ce)
	) name2798 (
		_w2799_,
		_w2812_,
		_w2813_,
		_w2823_,
		_w2824_
	);
	LUT3 #(
		.INIT('h1e)
	) name2799 (
		_w2076_,
		_w2817_,
		_w2824_,
		_w2825_
	);
	LUT4 #(
		.INIT('h153f)
	) name2800 (
		_w82_,
		_w106_,
		_w98_,
		_w71_,
		_w2826_
	);
	LUT4 #(
		.INIT('h0400)
	) name2801 (
		_w348_,
		_w429_,
		_w236_,
		_w2826_,
		_w2827_
	);
	LUT4 #(
		.INIT('hbbbf)
	) name2802 (
		_w46_,
		_w95_,
		_w102_,
		_w72_,
		_w2828_
	);
	LUT4 #(
		.INIT('h1000)
	) name2803 (
		_w197_,
		_w372_,
		_w1318_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h8000)
	) name2804 (
		_w231_,
		_w1443_,
		_w2827_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h8)
	) name2805 (
		_w562_,
		_w2830_,
		_w2831_
	);
	LUT2 #(
		.INIT('h8)
	) name2806 (
		_w2766_,
		_w2831_,
		_w2832_
	);
	LUT3 #(
		.INIT('hd0)
	) name2807 (
		_w2812_,
		_w2823_,
		_w2832_,
		_w2833_
	);
	LUT3 #(
		.INIT('h02)
	) name2808 (
		_w2812_,
		_w2823_,
		_w2832_,
		_w2834_
	);
	LUT3 #(
		.INIT('h2d)
	) name2809 (
		_w2812_,
		_w2823_,
		_w2832_,
		_w2835_
	);
	LUT3 #(
		.INIT('h08)
	) name2810 (
		_w2799_,
		_w2814_,
		_w2823_,
		_w2836_
	);
	LUT2 #(
		.INIT('h6)
	) name2811 (
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('h15)
	) name2812 (
		_w2076_,
		_w2817_,
		_w2824_,
		_w2838_
	);
	LUT2 #(
		.INIT('h6)
	) name2813 (
		_w2837_,
		_w2838_,
		_w2839_
	);
	LUT4 #(
		.INIT('h8008)
	) name2814 (
		_w2817_,
		_w2824_,
		_w2835_,
		_w2836_,
		_w2840_
	);
	LUT4 #(
		.INIT('h135f)
	) name2815 (
		_w88_,
		_w79_,
		_w98_,
		_w71_,
		_w2841_
	);
	LUT4 #(
		.INIT('h1000)
	) name2816 (
		_w352_,
		_w146_,
		_w2475_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('h8000)
	) name2817 (
		_w369_,
		_w411_,
		_w2367_,
		_w2842_,
		_w2843_
	);
	LUT3 #(
		.INIT('h80)
	) name2818 (
		_w513_,
		_w516_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		_w2527_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('h23dc)
	) name2820 (
		_w2833_,
		_w2834_,
		_w2836_,
		_w2845_,
		_w2846_
	);
	LUT3 #(
		.INIT('h1e)
	) name2821 (
		_w2076_,
		_w2840_,
		_w2846_,
		_w2847_
	);
	LUT4 #(
		.INIT('h0002)
	) name2822 (
		_w2812_,
		_w2823_,
		_w2832_,
		_w2845_,
		_w2848_
	);
	LUT4 #(
		.INIT('h4000)
	) name2823 (
		_w63_,
		_w385_,
		_w389_,
		_w392_,
		_w2849_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w1799_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		_w359_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h4)
	) name2826 (
		_w2848_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h2)
	) name2827 (
		_w2848_,
		_w2851_,
		_w2853_
	);
	LUT2 #(
		.INIT('h9)
	) name2828 (
		_w2848_,
		_w2851_,
		_w2854_
	);
	LUT3 #(
		.INIT('h08)
	) name2829 (
		_w2835_,
		_w2836_,
		_w2845_,
		_w2855_
	);
	LUT2 #(
		.INIT('h6)
	) name2830 (
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT3 #(
		.INIT('h15)
	) name2831 (
		_w2076_,
		_w2840_,
		_w2846_,
		_w2857_
	);
	LUT2 #(
		.INIT('h6)
	) name2832 (
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT4 #(
		.INIT('h8008)
	) name2833 (
		_w2840_,
		_w2846_,
		_w2854_,
		_w2855_,
		_w2859_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		_w359_,
		_w406_,
		_w2860_
	);
	LUT4 #(
		.INIT('h00b2)
	) name2835 (
		_w2848_,
		_w2851_,
		_w2855_,
		_w2860_,
		_w2861_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2836 (
		_w2848_,
		_w2851_,
		_w2855_,
		_w2860_,
		_w2862_
	);
	LUT4 #(
		.INIT('hdc23)
	) name2837 (
		_w2852_,
		_w2853_,
		_w2855_,
		_w2860_,
		_w2863_
	);
	LUT3 #(
		.INIT('he1)
	) name2838 (
		_w2076_,
		_w2859_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('he0)
	) name2839 (
		_w2076_,
		_w2859_,
		_w2861_,
		_w2865_
	);
	LUT4 #(
		.INIT('h0105)
	) name2840 (
		_w2076_,
		_w2859_,
		_w2861_,
		_w2862_,
		_w2866_
	);
	LUT2 #(
		.INIT('h1)
	) name2841 (
		\a[21] ,
		\a[22] ,
		_w2867_
	);
	LUT4 #(
		.INIT('h1000)
	) name2842 (
		\a[19] ,
		\a[20] ,
		_w49_,
		_w2867_,
		_w2868_
	);
	LUT3 #(
		.INIT('hfe)
	) name2843 (
		_w2866_,
		_w2865_,
		_w2868_,
		_w2869_
	);
	LUT3 #(
		.INIT('h02)
	) name2844 (
		_w2848_,
		_w2851_,
		_w2860_,
		_w2870_
	);
	LUT3 #(
		.INIT('h80)
	) name2845 (
		_w2854_,
		_w2855_,
		_w2870_,
		_w2871_
	);
	LUT3 #(
		.INIT('h0d)
	) name2846 (
		_w2859_,
		_w2863_,
		_w2871_,
		_w2872_
	);
	LUT3 #(
		.INIT('h07)
	) name2847 (
		_w2859_,
		_w2861_,
		_w2868_,
		_w2873_
	);
	LUT3 #(
		.INIT('h45)
	) name2848 (
		_w2076_,
		_w2872_,
		_w2873_,
		_w2874_
	);
	assign \sin[0]  = _w2075_ ;
	assign \sin[1]  = _w2149_ ;
	assign \sin[2]  = _w2211_ ;
	assign \sin[3]  = _w2269_ ;
	assign \sin[4]  = _w2324_ ;
	assign \sin[5]  = _w2380_ ;
	assign \sin[6]  = _w2436_ ;
	assign \sin[7]  = _w2489_ ;
	assign \sin[8]  = _w2538_ ;
	assign \sin[9]  = _w2581_ ;
	assign \sin[10]  = _w2622_ ;
	assign \sin[11]  = _w2656_ ;
	assign \sin[12]  = _w2693_ ;
	assign \sin[13]  = _w2727_ ;
	assign \sin[14]  = _w2755_ ;
	assign \sin[15]  = _w2780_ ;
	assign \sin[16]  = _w2803_ ;
	assign \sin[17]  = _w2816_ ;
	assign \sin[18]  = _w2825_ ;
	assign \sin[19]  = _w2839_ ;
	assign \sin[20]  = _w2847_ ;
	assign \sin[21]  = _w2858_ ;
	assign \sin[22]  = _w2864_ ;
	assign \sin[23]  = _w2869_ ;
	assign \sin[24]  = _w2874_ ;
endmodule;