module top( a_pad , b_pad , d_pad , \e0_pad  , f_pad , \g0_pad  , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , \a0_pad  , \b0_pad  , \c0_pad  , \d0_pad  , \f0_pad  , \h0_pad  , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad );
  input a_pad ;
  input b_pad ;
  input d_pad ;
  input \e0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  output \a0_pad  ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \d0_pad  ;
  output \f0_pad  ;
  output \h0_pad  ;
  output t_pad ;
  output u_pad ;
  output v_pad ;
  output w_pad ;
  output x_pad ;
  output y_pad ;
  output z_pad ;
  wire n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 ;
  assign n20 = g_pad & h_pad ;
  assign n21 = i_pad & n20 ;
  assign n22 = ~j_pad & n21 ;
  assign n25 = ~k_pad & n22 ;
  assign n26 = l_pad & ~n25 ;
  assign n23 = ~k_pad & ~l_pad ;
  assign n24 = n22 & n23 ;
  assign n27 = ~d_pad & \e0_pad  ;
  assign n28 = q_pad & ~n27 ;
  assign n29 = \g0_pad  & ~n28 ;
  assign n30 = ~n24 & n29 ;
  assign n31 = ~n26 & n30 ;
  assign n33 = m_pad & ~n24 ;
  assign n32 = ~m_pad & n24 ;
  assign n34 = n29 & ~n32 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = n_pad & ~n32 ;
  assign n37 = ~m_pad & ~n_pad ;
  assign n38 = n23 & n37 ;
  assign n39 = n22 & n38 ;
  assign n40 = n29 & ~n39 ;
  assign n41 = ~n36 & n40 ;
  assign n42 = o_pad & n28 ;
  assign n43 = ~a_pad & ~n38 ;
  assign n44 = n22 & ~n28 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = ~n42 & ~n45 ;
  assign n47 = \g0_pad  & ~n46 ;
  assign n48 = ~\e0_pad  & q_pad ;
  assign n49 = ~d_pad & ~n48 ;
  assign n50 = \g0_pad  & ~n49 ;
  assign n51 = \g0_pad  & r_pad ;
  assign n52 = b_pad & \e0_pad  ;
  assign n53 = ~b_pad & o_pad ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = ~p_pad & s_pad ;
  assign n56 = ~f_pad & ~n55 ;
  assign n57 = f_pad & ~\g0_pad  ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = ~g_pad & n29 ;
  assign n60 = ~g_pad & ~h_pad ;
  assign n61 = ~n20 & ~n60 ;
  assign n62 = n29 & n61 ;
  assign n63 = ~i_pad & ~n20 ;
  assign n64 = ~n21 & ~n63 ;
  assign n65 = n29 & n64 ;
  assign n66 = j_pad & ~n21 ;
  assign n67 = ~n22 & n29 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = k_pad & n67 ;
  assign n70 = ~n25 & n29 ;
  assign n71 = ~n69 & n70 ;
  assign \a0_pad  = ~n31 ;
  assign \b0_pad  = ~n35 ;
  assign \c0_pad  = ~n41 ;
  assign \d0_pad  = n47 ;
  assign \f0_pad  = n50 ;
  assign \h0_pad  = n51 ;
  assign t_pad = n54 ;
  assign u_pad = ~n58 ;
  assign v_pad = n59 ;
  assign w_pad = n62 ;
  assign x_pad = n65 ;
  assign y_pad = ~n68 ;
  assign z_pad = ~n71 ;
endmodule
