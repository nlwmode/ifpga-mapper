module top( \adr_i[0]_pad  , \adr_i[10]_pad  , \adr_i[1]_pad  , \adr_i[2]_pad  , \adr_i[3]_pad  , \adr_i[4]_pad  , \adr_i[5]_pad  , \adr_i[6]_pad  , \adr_i[7]_pad  , \adr_i[8]_pad  , \adr_i[9]_pad  , \adr_set_reg/NET0131  , \bits_transfered_reg[0]/NET0131  , \bits_transfered_reg[1]/NET0131  , \bits_transfered_reg[2]/NET0131  , \bits_transfered_reg[3]/NET0131  , \clk_gen_cnt_reg[0]/NET0131  , \clk_gen_cnt_reg[1]/NET0131  , \clk_gen_cnt_reg[2]/NET0131  , \clk_gen_cnt_reg[3]/NET0131  , \clk_gen_cnt_reg[4]/NET0131  , \clk_gen_cnt_reg[5]/NET0131  , \clk_gen_cnt_reg[6]/NET0131  , \clk_gen_cnt_reg[7]/NET0131  , \clk_gen_cnt_reg[8]/NET0131  , \dat_i[0]_pad  , \dat_i[1]_pad  , \dat_i[2]_pad  , \dat_i[3]_pad  , \dat_i[4]_pad  , \dat_i[5]_pad  , \dat_i[6]_pad  , \dat_i[7]_pad  , dat_rdy_o_pad , do_rnd_read_i_pad , do_seq_read_i_pad , do_write_i_pad , \doing_read_reg/NET0131  , \doing_seq_read_reg/NET0131  , \doing_write_reg/NET0131  , no_ack_o_pad , pci_spoci_sda_oe_o_pad , \rec_ack_reg/NET0131  , \rec_bit_reg/NET0131  , \rw_seq_state_reg[0]/NET0131  , \rw_seq_state_reg[1]/NET0131  , \rw_seq_state_reg[2]/NET0131  , \rw_seq_state_reg[3]/NET0131  , \rw_seq_state_reg[4]/NET0131  , \sda_i_reg_reg/NET0131  , \send_ack_reg/NET0131  , \send_bit_reg/NET0131  , \send_nack_reg/NET0131  , \send_start_reg/NET0131  , \send_stop_reg/NET0131  , \tx_rx_state_reg[0]/NET0131  , \tx_rx_state_reg[1]/NET0131  , \tx_rx_state_reg[2]/NET0131  , \tx_rx_state_reg[3]/NET0131  , \tx_rx_state_reg[4]/NET0131  , \tx_rx_state_reg[5]/NET0131  , \tx_rx_state_reg[6]/NET0131  , \tx_rx_state_reg[7]/NET0131  , \tx_rx_state_reg[8]/NET0131  , \tx_shift_reg_reg[0]/NET0131  , \tx_shift_reg_reg[1]/NET0131  , \tx_shift_reg_reg[2]/NET0131  , \tx_shift_reg_reg[3]/NET0131  , \tx_shift_reg_reg[4]/NET0131  , \tx_shift_reg_reg[5]/NET0131  , \tx_shift_reg_reg[6]/NET0131  , \tx_shift_reg_reg[7]/NET0131  , write_done_o_pad , \_al_n0  , \_al_n1  , \g4613/_2_  , \g4620/_0_  , \g4621/_0_  , \g4627/_0_  , \g4628/_0_  , \g4630/_0_  , \g4631/_0_  , \g4632/_0_  , \g4657/_0_  , \g4672/_0_  , \g4673/_0_  , \g4674/_0_  , \g4675/_0_  , \g4676/_0_  , \g4677/_0_  , \g4679/_0_  , \g4680/_0_  , \g4684/_0_  , \g4685/_0_  , \g4696/_0_  , \g4697/_0_  , \g4699/_0_  , \g4700/_0_  , \g4743/_0_  , \g4768/_0_  , \g4769/_0_  , \g4770/_0_  , \g4771/_0_  , \g4785/_0_  , \g4790/_0_  , \g4792/_0_  , \g4810/_0_  , \g4830/_0_  , \g4831/_0_  , \g4870/_0_  , \g4891/_0_  , \g4898/_0_  , \g4903/_0_  , \g4951/_2__syn_2  , \g4991/_3_  , \g5054/_0_  , \g5064/_0_  , \g5068/u3_syn_4  , \g5085/_1_  , \g5290/_0_  , \g5524/_0_  , \g5574/_2_  , \g57/_0_  , \g6488/_0_  , \g6585/_0_  , \g6602/_0_  , \g6658/_0_  , \g6720/_0_  , \g6767/_0_  , \g6827/_0_  );
  input \adr_i[0]_pad  ;
  input \adr_i[10]_pad  ;
  input \adr_i[1]_pad  ;
  input \adr_i[2]_pad  ;
  input \adr_i[3]_pad  ;
  input \adr_i[4]_pad  ;
  input \adr_i[5]_pad  ;
  input \adr_i[6]_pad  ;
  input \adr_i[7]_pad  ;
  input \adr_i[8]_pad  ;
  input \adr_i[9]_pad  ;
  input \adr_set_reg/NET0131  ;
  input \bits_transfered_reg[0]/NET0131  ;
  input \bits_transfered_reg[1]/NET0131  ;
  input \bits_transfered_reg[2]/NET0131  ;
  input \bits_transfered_reg[3]/NET0131  ;
  input \clk_gen_cnt_reg[0]/NET0131  ;
  input \clk_gen_cnt_reg[1]/NET0131  ;
  input \clk_gen_cnt_reg[2]/NET0131  ;
  input \clk_gen_cnt_reg[3]/NET0131  ;
  input \clk_gen_cnt_reg[4]/NET0131  ;
  input \clk_gen_cnt_reg[5]/NET0131  ;
  input \clk_gen_cnt_reg[6]/NET0131  ;
  input \clk_gen_cnt_reg[7]/NET0131  ;
  input \clk_gen_cnt_reg[8]/NET0131  ;
  input \dat_i[0]_pad  ;
  input \dat_i[1]_pad  ;
  input \dat_i[2]_pad  ;
  input \dat_i[3]_pad  ;
  input \dat_i[4]_pad  ;
  input \dat_i[5]_pad  ;
  input \dat_i[6]_pad  ;
  input \dat_i[7]_pad  ;
  input dat_rdy_o_pad ;
  input do_rnd_read_i_pad ;
  input do_seq_read_i_pad ;
  input do_write_i_pad ;
  input \doing_read_reg/NET0131  ;
  input \doing_seq_read_reg/NET0131  ;
  input \doing_write_reg/NET0131  ;
  input no_ack_o_pad ;
  input pci_spoci_sda_oe_o_pad ;
  input \rec_ack_reg/NET0131  ;
  input \rec_bit_reg/NET0131  ;
  input \rw_seq_state_reg[0]/NET0131  ;
  input \rw_seq_state_reg[1]/NET0131  ;
  input \rw_seq_state_reg[2]/NET0131  ;
  input \rw_seq_state_reg[3]/NET0131  ;
  input \rw_seq_state_reg[4]/NET0131  ;
  input \sda_i_reg_reg/NET0131  ;
  input \send_ack_reg/NET0131  ;
  input \send_bit_reg/NET0131  ;
  input \send_nack_reg/NET0131  ;
  input \send_start_reg/NET0131  ;
  input \send_stop_reg/NET0131  ;
  input \tx_rx_state_reg[0]/NET0131  ;
  input \tx_rx_state_reg[1]/NET0131  ;
  input \tx_rx_state_reg[2]/NET0131  ;
  input \tx_rx_state_reg[3]/NET0131  ;
  input \tx_rx_state_reg[4]/NET0131  ;
  input \tx_rx_state_reg[5]/NET0131  ;
  input \tx_rx_state_reg[6]/NET0131  ;
  input \tx_rx_state_reg[7]/NET0131  ;
  input \tx_rx_state_reg[8]/NET0131  ;
  input \tx_shift_reg_reg[0]/NET0131  ;
  input \tx_shift_reg_reg[1]/NET0131  ;
  input \tx_shift_reg_reg[2]/NET0131  ;
  input \tx_shift_reg_reg[3]/NET0131  ;
  input \tx_shift_reg_reg[4]/NET0131  ;
  input \tx_shift_reg_reg[5]/NET0131  ;
  input \tx_shift_reg_reg[6]/NET0131  ;
  input \tx_shift_reg_reg[7]/NET0131  ;
  input write_done_o_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g4613/_2_  ;
  output \g4620/_0_  ;
  output \g4621/_0_  ;
  output \g4627/_0_  ;
  output \g4628/_0_  ;
  output \g4630/_0_  ;
  output \g4631/_0_  ;
  output \g4632/_0_  ;
  output \g4657/_0_  ;
  output \g4672/_0_  ;
  output \g4673/_0_  ;
  output \g4674/_0_  ;
  output \g4675/_0_  ;
  output \g4676/_0_  ;
  output \g4677/_0_  ;
  output \g4679/_0_  ;
  output \g4680/_0_  ;
  output \g4684/_0_  ;
  output \g4685/_0_  ;
  output \g4696/_0_  ;
  output \g4697/_0_  ;
  output \g4699/_0_  ;
  output \g4700/_0_  ;
  output \g4743/_0_  ;
  output \g4768/_0_  ;
  output \g4769/_0_  ;
  output \g4770/_0_  ;
  output \g4771/_0_  ;
  output \g4785/_0_  ;
  output \g4790/_0_  ;
  output \g4792/_0_  ;
  output \g4810/_0_  ;
  output \g4830/_0_  ;
  output \g4831/_0_  ;
  output \g4870/_0_  ;
  output \g4891/_0_  ;
  output \g4898/_0_  ;
  output \g4903/_0_  ;
  output \g4951/_2__syn_2  ;
  output \g4991/_3_  ;
  output \g5054/_0_  ;
  output \g5064/_0_  ;
  output \g5068/u3_syn_4  ;
  output \g5085/_1_  ;
  output \g5290/_0_  ;
  output \g5524/_0_  ;
  output \g5574/_2_  ;
  output \g57/_0_  ;
  output \g6488/_0_  ;
  output \g6585/_0_  ;
  output \g6602/_0_  ;
  output \g6658/_0_  ;
  output \g6720/_0_  ;
  output \g6767/_0_  ;
  output \g6827/_0_  ;
  wire n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 ;
  assign n74 = \clk_gen_cnt_reg[3]/NET0131  & \clk_gen_cnt_reg[4]/NET0131  ;
  assign n75 = \clk_gen_cnt_reg[5]/NET0131  & \clk_gen_cnt_reg[6]/NET0131  ;
  assign n76 = n74 & n75 ;
  assign n77 = \clk_gen_cnt_reg[7]/NET0131  & n76 ;
  assign n78 = ~\clk_gen_cnt_reg[0]/NET0131  & \clk_gen_cnt_reg[1]/NET0131  ;
  assign n79 = ~\clk_gen_cnt_reg[2]/NET0131  & ~\clk_gen_cnt_reg[8]/NET0131  ;
  assign n80 = n78 & n79 ;
  assign n81 = n77 & n80 ;
  assign n82 = ~\tx_rx_state_reg[1]/NET0131  & ~\tx_rx_state_reg[4]/NET0131  ;
  assign n83 = ~\tx_rx_state_reg[2]/NET0131  & ~\tx_rx_state_reg[3]/NET0131  ;
  assign n84 = n82 & n83 ;
  assign n85 = ~\tx_rx_state_reg[7]/NET0131  & ~\tx_rx_state_reg[8]/NET0131  ;
  assign n86 = n84 & n85 ;
  assign n87 = ~\tx_rx_state_reg[0]/NET0131  & ~\tx_rx_state_reg[5]/NET0131  ;
  assign n88 = \tx_rx_state_reg[6]/NET0131  & n87 ;
  assign n89 = n86 & n88 ;
  assign n90 = n81 & n89 ;
  assign n91 = ~\send_stop_reg/NET0131  & ~n90 ;
  assign n92 = \rec_ack_reg/NET0131  & ~\send_bit_reg/NET0131  ;
  assign n93 = ~\sda_i_reg_reg/NET0131  & n80 ;
  assign n94 = n77 & n93 ;
  assign n95 = n89 & n94 ;
  assign n96 = n92 & ~n95 ;
  assign n97 = ~n91 & n96 ;
  assign n98 = ~\rw_seq_state_reg[2]/NET0131  & ~\rw_seq_state_reg[4]/NET0131  ;
  assign n99 = \rw_seq_state_reg[1]/NET0131  & n98 ;
  assign n100 = \send_start_reg/NET0131  & ~\send_stop_reg/NET0131  ;
  assign n101 = ~\rw_seq_state_reg[0]/NET0131  & ~\rw_seq_state_reg[3]/NET0131  ;
  assign n102 = ~n100 & n101 ;
  assign n103 = n99 & n102 ;
  assign n104 = ~\rw_seq_state_reg[1]/NET0131  & n101 ;
  assign n105 = \rw_seq_state_reg[2]/NET0131  & ~\rw_seq_state_reg[4]/NET0131  ;
  assign n106 = n104 & n105 ;
  assign n107 = ~n103 & ~n106 ;
  assign n108 = n97 & ~n107 ;
  assign n109 = ~\clk_gen_cnt_reg[4]/NET0131  & ~\clk_gen_cnt_reg[7]/NET0131  ;
  assign n110 = \clk_gen_cnt_reg[8]/NET0131  & n109 ;
  assign n111 = ~\clk_gen_cnt_reg[5]/NET0131  & \clk_gen_cnt_reg[6]/NET0131  ;
  assign n112 = \clk_gen_cnt_reg[2]/NET0131  & \clk_gen_cnt_reg[3]/NET0131  ;
  assign n113 = n78 & n112 ;
  assign n114 = n111 & n113 ;
  assign n115 = n110 & n114 ;
  assign n116 = ~\tx_rx_state_reg[7]/NET0131  & n84 ;
  assign n117 = ~\tx_rx_state_reg[0]/NET0131  & ~\tx_rx_state_reg[6]/NET0131  ;
  assign n118 = ~\tx_rx_state_reg[5]/NET0131  & \tx_rx_state_reg[8]/NET0131  ;
  assign n119 = n117 & n118 ;
  assign n120 = n116 & n119 ;
  assign n121 = n115 & n120 ;
  assign n122 = ~\rec_ack_reg/NET0131  & ~\send_bit_reg/NET0131  ;
  assign n123 = n121 & n122 ;
  assign n124 = ~n96 & ~n123 ;
  assign n125 = \send_stop_reg/NET0131  & ~n107 ;
  assign n126 = n124 & n125 ;
  assign n127 = ~n108 & ~n126 ;
  assign n128 = ~n91 & n92 ;
  assign n129 = \send_bit_reg/NET0131  & \send_stop_reg/NET0131  ;
  assign n130 = ~\rec_ack_reg/NET0131  & \send_stop_reg/NET0131  ;
  assign n131 = ~n121 & n130 ;
  assign n132 = ~n129 & ~n131 ;
  assign n133 = ~n128 & n132 ;
  assign n134 = ~\rw_seq_state_reg[1]/NET0131  & n98 ;
  assign n135 = ~\rw_seq_state_reg[0]/NET0131  & \rw_seq_state_reg[3]/NET0131  ;
  assign n136 = n134 & n135 ;
  assign n137 = ~n133 & n136 ;
  assign n138 = ~\clk_gen_cnt_reg[7]/NET0131  & n79 ;
  assign n139 = \clk_gen_cnt_reg[0]/NET0131  & \clk_gen_cnt_reg[1]/NET0131  ;
  assign n140 = ~\clk_gen_cnt_reg[3]/NET0131  & \clk_gen_cnt_reg[4]/NET0131  ;
  assign n141 = n111 & n140 ;
  assign n142 = n139 & n141 ;
  assign n143 = n138 & n142 ;
  assign n144 = \tx_rx_state_reg[7]/NET0131  & ~\tx_rx_state_reg[8]/NET0131  ;
  assign n145 = n84 & n144 ;
  assign n146 = ~\tx_rx_state_reg[5]/NET0131  & n117 ;
  assign n147 = ~\rec_bit_reg/NET0131  & \send_nack_reg/NET0131  ;
  assign n148 = n146 & n147 ;
  assign n149 = n145 & n148 ;
  assign n150 = n143 & n149 ;
  assign n151 = ~\rw_seq_state_reg[2]/NET0131  & \rw_seq_state_reg[4]/NET0131  ;
  assign n152 = n104 & n151 ;
  assign n153 = n150 & n152 ;
  assign n154 = ~\rec_bit_reg/NET0131  & ~\send_ack_reg/NET0131  ;
  assign n155 = ~\send_nack_reg/NET0131  & n154 ;
  assign n156 = n110 & n155 ;
  assign n157 = n114 & n156 ;
  assign n158 = n120 & n157 ;
  assign n159 = \send_stop_reg/NET0131  & n152 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = ~n153 & ~n160 ;
  assign n162 = ~n106 & ~n136 ;
  assign n163 = n99 & n101 ;
  assign n164 = ~n152 & ~n163 ;
  assign n165 = n162 & n164 ;
  assign n166 = \send_start_reg/NET0131  & n101 ;
  assign n167 = n99 & n166 ;
  assign n168 = ~n165 & ~n167 ;
  assign n169 = \send_stop_reg/NET0131  & ~n168 ;
  assign n170 = n161 & ~n169 ;
  assign n171 = ~n137 & n170 ;
  assign n172 = n127 & n171 ;
  assign n173 = \send_start_reg/NET0131  & \tx_shift_reg_reg[2]/NET0131  ;
  assign n174 = \adr_set_reg/NET0131  & ~\doing_write_reg/NET0131  ;
  assign n175 = \rec_ack_reg/NET0131  & ~n174 ;
  assign n176 = n95 & n175 ;
  assign n177 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[2]/NET0131  ;
  assign n178 = ~n176 & n177 ;
  assign n179 = ~n173 & ~n178 ;
  assign n180 = n163 & ~n179 ;
  assign n181 = \adr_i[2]_pad  & n92 ;
  assign n182 = ~n174 & n181 ;
  assign n183 = n95 & n182 ;
  assign n184 = ~\tx_rx_state_reg[5]/NET0131  & ~\tx_rx_state_reg[7]/NET0131  ;
  assign n185 = ~\tx_rx_state_reg[6]/NET0131  & ~\tx_rx_state_reg[8]/NET0131  ;
  assign n186 = n184 & n185 ;
  assign n187 = n82 & n186 ;
  assign n188 = ~\tx_rx_state_reg[0]/NET0131  & ~\tx_rx_state_reg[2]/NET0131  ;
  assign n189 = \tx_rx_state_reg[3]/NET0131  & n188 ;
  assign n190 = n187 & n189 ;
  assign n191 = n143 & n190 ;
  assign n192 = ~\tx_shift_reg_reg[2]/NET0131  & ~n191 ;
  assign n193 = ~\tx_shift_reg_reg[1]/NET0131  & n138 ;
  assign n194 = n142 & n193 ;
  assign n195 = n190 & n194 ;
  assign n196 = \send_bit_reg/NET0131  & ~n195 ;
  assign n197 = ~n192 & n196 ;
  assign n198 = ~n183 & ~n197 ;
  assign n199 = ~\send_start_reg/NET0131  & n163 ;
  assign n200 = ~n198 & n199 ;
  assign n201 = ~n180 & ~n200 ;
  assign n202 = \dat_i[2]_pad  & \doing_write_reg/NET0131  ;
  assign n203 = n95 & n202 ;
  assign n204 = n92 & n203 ;
  assign n205 = ~\doing_read_reg/NET0131  & ~\doing_seq_read_reg/NET0131  ;
  assign n206 = ~\doing_write_reg/NET0131  & n205 ;
  assign n207 = n95 & ~n206 ;
  assign n208 = \tx_shift_reg_reg[2]/NET0131  & n92 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = ~n204 & ~n209 ;
  assign n211 = ~\rec_ack_reg/NET0131  & n177 ;
  assign n212 = ~n197 & ~n211 ;
  assign n213 = n210 & n212 ;
  assign n214 = n106 & ~n213 ;
  assign n215 = ~n177 & ~n197 ;
  assign n216 = n136 & ~n215 ;
  assign n217 = \rw_seq_state_reg[0]/NET0131  & ~\rw_seq_state_reg[3]/NET0131  ;
  assign n218 = n134 & n217 ;
  assign n219 = ~n163 & ~n218 ;
  assign n220 = n162 & n219 ;
  assign n221 = \tx_shift_reg_reg[2]/NET0131  & n220 ;
  assign n222 = \adr_i[9]_pad  & n217 ;
  assign n223 = n134 & n222 ;
  assign n224 = ~n221 & ~n223 ;
  assign n225 = ~n216 & n224 ;
  assign n226 = ~n214 & n225 ;
  assign n227 = n201 & n226 ;
  assign n228 = \dat_i[4]_pad  & \rec_ack_reg/NET0131  ;
  assign n229 = \doing_write_reg/NET0131  & n228 ;
  assign n230 = n95 & n229 ;
  assign n231 = ~\send_bit_reg/NET0131  & n230 ;
  assign n232 = \rec_ack_reg/NET0131  & ~n206 ;
  assign n233 = n95 & n232 ;
  assign n234 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[4]/NET0131  ;
  assign n235 = ~n233 & n234 ;
  assign n236 = ~n231 & ~n235 ;
  assign n237 = ~\tx_shift_reg_reg[4]/NET0131  & ~n191 ;
  assign n238 = ~\tx_shift_reg_reg[3]/NET0131  & n138 ;
  assign n239 = n142 & n238 ;
  assign n240 = n190 & n239 ;
  assign n241 = \send_bit_reg/NET0131  & ~n240 ;
  assign n242 = ~n237 & n241 ;
  assign n243 = n236 & ~n242 ;
  assign n244 = n106 & ~n243 ;
  assign n245 = ~\adr_i[4]_pad  & ~n174 ;
  assign n246 = n95 & n245 ;
  assign n247 = ~\send_bit_reg/NET0131  & ~\send_start_reg/NET0131  ;
  assign n248 = \rec_ack_reg/NET0131  & n247 ;
  assign n249 = \tx_shift_reg_reg[4]/NET0131  & n248 ;
  assign n250 = ~n174 & n248 ;
  assign n251 = n95 & n250 ;
  assign n252 = ~n249 & ~n251 ;
  assign n253 = ~n246 & ~n252 ;
  assign n254 = \send_bit_reg/NET0131  & ~\send_start_reg/NET0131  ;
  assign n255 = ~n240 & n254 ;
  assign n256 = ~n237 & n255 ;
  assign n257 = ~\send_start_reg/NET0131  & ~n122 ;
  assign n258 = \tx_shift_reg_reg[4]/NET0131  & ~n257 ;
  assign n259 = ~n256 & ~n258 ;
  assign n260 = ~n253 & n259 ;
  assign n261 = n163 & ~n260 ;
  assign n262 = \tx_shift_reg_reg[4]/NET0131  & n220 ;
  assign n263 = ~n136 & ~n262 ;
  assign n264 = ~n234 & ~n262 ;
  assign n265 = ~n242 & n264 ;
  assign n266 = ~n263 & ~n265 ;
  assign n267 = ~n261 & ~n266 ;
  assign n268 = ~n244 & n267 ;
  assign n269 = \send_start_reg/NET0131  & \tx_shift_reg_reg[1]/NET0131  ;
  assign n270 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[1]/NET0131  ;
  assign n271 = ~n176 & n270 ;
  assign n272 = ~n269 & ~n271 ;
  assign n273 = n163 & ~n272 ;
  assign n274 = \adr_i[1]_pad  & n92 ;
  assign n275 = ~n174 & n274 ;
  assign n276 = n95 & n275 ;
  assign n277 = ~\tx_shift_reg_reg[1]/NET0131  & ~n191 ;
  assign n278 = ~\tx_shift_reg_reg[0]/NET0131  & n138 ;
  assign n279 = n142 & n278 ;
  assign n280 = n190 & n279 ;
  assign n281 = \send_bit_reg/NET0131  & ~n280 ;
  assign n282 = ~n277 & n281 ;
  assign n283 = ~n276 & ~n282 ;
  assign n284 = n199 & ~n283 ;
  assign n285 = ~n273 & ~n284 ;
  assign n286 = \dat_i[1]_pad  & \doing_write_reg/NET0131  ;
  assign n287 = n95 & n286 ;
  assign n288 = n92 & n287 ;
  assign n289 = \tx_shift_reg_reg[1]/NET0131  & n92 ;
  assign n290 = ~n207 & n289 ;
  assign n291 = ~n288 & ~n290 ;
  assign n292 = ~\rec_ack_reg/NET0131  & n270 ;
  assign n293 = ~n282 & ~n292 ;
  assign n294 = n291 & n293 ;
  assign n295 = n106 & ~n294 ;
  assign n296 = ~n270 & ~n282 ;
  assign n297 = n136 & ~n296 ;
  assign n298 = \tx_shift_reg_reg[1]/NET0131  & n220 ;
  assign n299 = \adr_i[8]_pad  & n217 ;
  assign n300 = n134 & n299 ;
  assign n301 = ~n298 & ~n300 ;
  assign n302 = ~n297 & n301 ;
  assign n303 = ~n295 & n302 ;
  assign n304 = n285 & n303 ;
  assign n305 = \send_start_reg/NET0131  & \tx_shift_reg_reg[3]/NET0131  ;
  assign n306 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[3]/NET0131  ;
  assign n307 = ~n176 & n306 ;
  assign n308 = ~n305 & ~n307 ;
  assign n309 = n163 & ~n308 ;
  assign n310 = \adr_i[3]_pad  & n92 ;
  assign n311 = ~n174 & n310 ;
  assign n312 = n95 & n311 ;
  assign n313 = ~\tx_shift_reg_reg[3]/NET0131  & ~n191 ;
  assign n314 = ~\tx_shift_reg_reg[2]/NET0131  & n138 ;
  assign n315 = n142 & n314 ;
  assign n316 = n190 & n315 ;
  assign n317 = \send_bit_reg/NET0131  & ~n316 ;
  assign n318 = ~n313 & n317 ;
  assign n319 = ~n312 & ~n318 ;
  assign n320 = n199 & ~n319 ;
  assign n321 = ~n309 & ~n320 ;
  assign n322 = \dat_i[3]_pad  & \doing_write_reg/NET0131  ;
  assign n323 = n95 & n322 ;
  assign n324 = n92 & n323 ;
  assign n325 = \tx_shift_reg_reg[3]/NET0131  & n92 ;
  assign n326 = ~n207 & n325 ;
  assign n327 = ~n324 & ~n326 ;
  assign n328 = ~\rec_ack_reg/NET0131  & n306 ;
  assign n329 = ~n318 & ~n328 ;
  assign n330 = n327 & n329 ;
  assign n331 = n106 & ~n330 ;
  assign n332 = ~n306 & ~n318 ;
  assign n333 = n136 & ~n332 ;
  assign n334 = \tx_shift_reg_reg[3]/NET0131  & n220 ;
  assign n335 = \adr_i[10]_pad  & n217 ;
  assign n336 = n134 & n335 ;
  assign n337 = ~n334 & ~n336 ;
  assign n338 = ~n333 & n337 ;
  assign n339 = ~n331 & n338 ;
  assign n340 = n321 & n339 ;
  assign n341 = n162 & ~n163 ;
  assign n342 = \send_stop_reg/NET0131  & n122 ;
  assign n343 = ~n167 & n342 ;
  assign n344 = ~n341 & n343 ;
  assign n345 = no_ack_o_pad & ~n344 ;
  assign n346 = ~\send_start_reg/NET0131  & n101 ;
  assign n347 = n99 & n346 ;
  assign n348 = n162 & ~n347 ;
  assign n349 = \sda_i_reg_reg/NET0131  & n92 ;
  assign n350 = ~n348 & n349 ;
  assign n351 = n90 & n350 ;
  assign n352 = ~n345 & ~n351 ;
  assign n353 = ~\tx_shift_reg_reg[5]/NET0131  & ~n191 ;
  assign n354 = ~\tx_shift_reg_reg[4]/NET0131  & n138 ;
  assign n355 = n142 & n354 ;
  assign n356 = n190 & n355 ;
  assign n357 = n254 & ~n356 ;
  assign n358 = ~n353 & n357 ;
  assign n359 = ~\tx_shift_reg_reg[5]/NET0131  & ~n176 ;
  assign n360 = ~\adr_i[5]_pad  & \rec_ack_reg/NET0131  ;
  assign n361 = ~n174 & n360 ;
  assign n362 = n95 & n361 ;
  assign n363 = n247 & ~n362 ;
  assign n364 = ~n359 & n363 ;
  assign n365 = ~n358 & ~n364 ;
  assign n366 = n163 & ~n365 ;
  assign n367 = ~\tx_shift_reg_reg[5]/NET0131  & ~n207 ;
  assign n368 = ~\dat_i[5]_pad  & \doing_write_reg/NET0131  ;
  assign n369 = n95 & n368 ;
  assign n370 = n92 & ~n369 ;
  assign n371 = ~n367 & n370 ;
  assign n372 = \send_bit_reg/NET0131  & ~n356 ;
  assign n373 = ~n353 & n372 ;
  assign n374 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[5]/NET0131  ;
  assign n375 = ~\rec_ack_reg/NET0131  & n374 ;
  assign n376 = ~n373 & ~n375 ;
  assign n377 = ~n371 & n376 ;
  assign n378 = n106 & ~n377 ;
  assign n379 = ~n373 & ~n374 ;
  assign n380 = n136 & ~n379 ;
  assign n381 = \tx_shift_reg_reg[5]/NET0131  & n167 ;
  assign n382 = \tx_shift_reg_reg[5]/NET0131  & ~n163 ;
  assign n383 = n162 & n382 ;
  assign n384 = ~n381 & ~n383 ;
  assign n385 = ~n218 & n384 ;
  assign n386 = ~n380 & n385 ;
  assign n387 = ~n378 & n386 ;
  assign n388 = ~n366 & n387 ;
  assign n389 = \send_start_reg/NET0131  & \tx_shift_reg_reg[7]/NET0131  ;
  assign n390 = ~\send_bit_reg/NET0131  & \tx_shift_reg_reg[7]/NET0131  ;
  assign n391 = ~n176 & n390 ;
  assign n392 = ~n389 & ~n391 ;
  assign n393 = n163 & ~n392 ;
  assign n394 = \adr_i[7]_pad  & n92 ;
  assign n395 = ~n174 & n394 ;
  assign n396 = n95 & n395 ;
  assign n397 = ~\tx_shift_reg_reg[7]/NET0131  & ~n191 ;
  assign n398 = ~\tx_shift_reg_reg[6]/NET0131  & n138 ;
  assign n399 = n142 & n398 ;
  assign n400 = n190 & n399 ;
  assign n401 = \send_bit_reg/NET0131  & ~n400 ;
  assign n402 = ~n397 & n401 ;
  assign n403 = ~n396 & ~n402 ;
  assign n404 = n199 & ~n403 ;
  assign n405 = ~n393 & ~n404 ;
  assign n406 = ~\tx_shift_reg_reg[7]/NET0131  & ~n207 ;
  assign n407 = ~\dat_i[7]_pad  & \doing_write_reg/NET0131  ;
  assign n408 = n95 & n407 ;
  assign n409 = n92 & ~n408 ;
  assign n410 = ~n406 & n409 ;
  assign n411 = ~\rec_ack_reg/NET0131  & n390 ;
  assign n412 = ~n402 & ~n411 ;
  assign n413 = ~n410 & n412 ;
  assign n414 = n106 & ~n413 ;
  assign n415 = \tx_shift_reg_reg[7]/NET0131  & ~n163 ;
  assign n416 = n162 & n415 ;
  assign n417 = ~n218 & ~n416 ;
  assign n418 = ~n136 & n417 ;
  assign n419 = ~n390 & n417 ;
  assign n420 = ~n402 & n419 ;
  assign n421 = ~n418 & ~n420 ;
  assign n422 = ~n414 & ~n421 ;
  assign n423 = n405 & n422 ;
  assign n424 = n110 & n122 ;
  assign n425 = n114 & n424 ;
  assign n426 = n190 & n425 ;
  assign n427 = ~n143 & ~n426 ;
  assign n428 = n145 & n146 ;
  assign n429 = ~n89 & ~n428 ;
  assign n430 = \tx_rx_state_reg[4]/NET0131  & n186 ;
  assign n431 = ~\tx_rx_state_reg[1]/NET0131  & ~\tx_rx_state_reg[3]/NET0131  ;
  assign n432 = n188 & n431 ;
  assign n433 = n430 & n432 ;
  assign n434 = ~n190 & ~n433 ;
  assign n435 = n429 & n434 ;
  assign n436 = \tx_rx_state_reg[5]/NET0131  & \tx_rx_state_reg[8]/NET0131  ;
  assign n437 = ~\tx_rx_state_reg[5]/NET0131  & ~\tx_rx_state_reg[8]/NET0131  ;
  assign n438 = n117 & ~n437 ;
  assign n439 = ~n436 & n438 ;
  assign n440 = n116 & n439 ;
  assign n441 = ~\tx_rx_state_reg[0]/NET0131  & \tx_rx_state_reg[2]/NET0131  ;
  assign n442 = ~\tx_rx_state_reg[3]/NET0131  & n441 ;
  assign n443 = n187 & n442 ;
  assign n444 = ~n440 & ~n443 ;
  assign n445 = n435 & n444 ;
  assign n446 = ~n427 & ~n445 ;
  assign n447 = ~\tx_rx_state_reg[3]/NET0131  & n188 ;
  assign n448 = \tx_rx_state_reg[1]/NET0131  & ~\tx_rx_state_reg[4]/NET0131  ;
  assign n449 = n447 & n448 ;
  assign n450 = n186 & n449 ;
  assign n451 = \clk_gen_cnt_reg[2]/NET0131  & n139 ;
  assign n452 = ~\clk_gen_cnt_reg[3]/NET0131  & ~\clk_gen_cnt_reg[4]/NET0131  ;
  assign n453 = \clk_gen_cnt_reg[5]/NET0131  & ~\clk_gen_cnt_reg[6]/NET0131  ;
  assign n454 = \clk_gen_cnt_reg[7]/NET0131  & ~\clk_gen_cnt_reg[8]/NET0131  ;
  assign n455 = n453 & n454 ;
  assign n456 = n452 & n455 ;
  assign n457 = n451 & n456 ;
  assign n458 = n450 & n457 ;
  assign n459 = ~n115 & n458 ;
  assign n460 = \tx_rx_state_reg[5]/NET0131  & n117 ;
  assign n461 = n86 & n460 ;
  assign n462 = ~\rec_bit_reg/NET0131  & n110 ;
  assign n463 = n114 & n462 ;
  assign n464 = n461 & n463 ;
  assign n465 = ~n459 & ~n464 ;
  assign n466 = ~\send_bit_reg/NET0131  & n110 ;
  assign n467 = n114 & n466 ;
  assign n468 = n450 & n467 ;
  assign n469 = ~n121 & ~n468 ;
  assign n470 = pci_spoci_sda_oe_o_pad & n469 ;
  assign n471 = n465 & n470 ;
  assign n472 = ~n446 & n471 ;
  assign n473 = n465 & n469 ;
  assign n474 = ~n446 & n473 ;
  assign n475 = n450 & ~n467 ;
  assign n476 = ~\tx_shift_reg_reg[7]/NET0131  & n189 ;
  assign n477 = n187 & n476 ;
  assign n478 = ~n440 & ~n477 ;
  assign n479 = n143 & ~n478 ;
  assign n480 = ~n475 & ~n479 ;
  assign n481 = ~n474 & n480 ;
  assign n482 = ~n472 & ~n481 ;
  assign n483 = \doing_write_reg/NET0131  & n92 ;
  assign n484 = n95 & n483 ;
  assign n485 = n106 & n484 ;
  assign n486 = n92 & n95 ;
  assign n487 = \send_stop_reg/NET0131  & n110 ;
  assign n488 = n114 & n487 ;
  assign n489 = n120 & n488 ;
  assign n490 = n122 & n489 ;
  assign n491 = ~n486 & ~n490 ;
  assign n492 = ~\rec_ack_reg/NET0131  & n489 ;
  assign n493 = n205 & ~n492 ;
  assign n494 = ~n491 & ~n493 ;
  assign n495 = \rw_seq_state_reg[3]/NET0131  & n106 ;
  assign n496 = ~n494 & n495 ;
  assign n497 = ~n485 & ~n496 ;
  assign n498 = \rw_seq_state_reg[3]/NET0131  & n165 ;
  assign n499 = n110 & n342 ;
  assign n500 = n114 & n499 ;
  assign n501 = n120 & n500 ;
  assign n502 = n136 & ~n501 ;
  assign n503 = ~n498 & ~n502 ;
  assign n504 = n497 & n503 ;
  assign n505 = \tx_rx_state_reg[0]/NET0131  & n84 ;
  assign n506 = n186 & n505 ;
  assign n507 = ~n450 & ~n506 ;
  assign n508 = n444 & n507 ;
  assign n509 = n435 & n508 ;
  assign n510 = \clk_gen_cnt_reg[0]/NET0131  & ~n506 ;
  assign n511 = ~n509 & n510 ;
  assign n512 = ~\clk_gen_cnt_reg[1]/NET0131  & ~n511 ;
  assign n513 = n139 & ~n506 ;
  assign n514 = ~n509 & n513 ;
  assign n515 = ~n450 & ~n461 ;
  assign n516 = n435 & n515 ;
  assign n517 = n115 & ~n516 ;
  assign n518 = n443 & n457 ;
  assign n519 = \send_start_reg/NET0131  & n186 ;
  assign n520 = n505 & n519 ;
  assign n521 = ~n518 & ~n520 ;
  assign n522 = ~n517 & n521 ;
  assign n523 = ~n514 & n522 ;
  assign n524 = ~n512 & n523 ;
  assign n525 = ~\clk_gen_cnt_reg[2]/NET0131  & ~n514 ;
  assign n526 = n451 & ~n506 ;
  assign n527 = ~n509 & n526 ;
  assign n528 = n522 & ~n527 ;
  assign n529 = ~n525 & n528 ;
  assign n530 = \clk_gen_cnt_reg[3]/NET0131  & n451 ;
  assign n531 = ~n506 & n530 ;
  assign n532 = ~n509 & n531 ;
  assign n533 = ~\clk_gen_cnt_reg[3]/NET0131  & ~n527 ;
  assign n534 = n522 & ~n533 ;
  assign n535 = ~n532 & n534 ;
  assign n536 = ~\clk_gen_cnt_reg[4]/NET0131  & ~n532 ;
  assign n537 = n74 & n451 ;
  assign n538 = ~n506 & n537 ;
  assign n539 = ~n509 & n538 ;
  assign n540 = n522 & ~n539 ;
  assign n541 = ~n536 & n540 ;
  assign n542 = \clk_gen_cnt_reg[5]/NET0131  & n539 ;
  assign n543 = ~\clk_gen_cnt_reg[5]/NET0131  & ~n539 ;
  assign n544 = n522 & ~n543 ;
  assign n545 = ~n542 & n544 ;
  assign n546 = n76 & n451 ;
  assign n547 = ~n506 & n546 ;
  assign n548 = ~n509 & n547 ;
  assign n549 = ~\clk_gen_cnt_reg[7]/NET0131  & ~n548 ;
  assign n550 = n77 & n451 ;
  assign n551 = ~n506 & n550 ;
  assign n552 = ~n509 & n551 ;
  assign n553 = n522 & ~n552 ;
  assign n554 = ~n549 & n553 ;
  assign n555 = \clk_gen_cnt_reg[8]/NET0131  & n552 ;
  assign n556 = ~\clk_gen_cnt_reg[8]/NET0131  & ~n552 ;
  assign n557 = n522 & ~n556 ;
  assign n558 = ~n555 & n557 ;
  assign n559 = n165 & ~n218 ;
  assign n560 = \rw_seq_state_reg[1]/NET0131  & n559 ;
  assign n561 = ~n106 & ~n347 ;
  assign n562 = \rw_seq_state_reg[1]/NET0131  & ~n561 ;
  assign n563 = n491 & n562 ;
  assign n564 = ~n560 & ~n563 ;
  assign n565 = \rec_ack_reg/NET0131  & n105 ;
  assign n566 = n104 & n565 ;
  assign n567 = ~\rw_seq_state_reg[1]/NET0131  & n205 ;
  assign n568 = ~\send_bit_reg/NET0131  & ~n567 ;
  assign n569 = n566 & n568 ;
  assign n570 = ~\doing_write_reg/NET0131  & n569 ;
  assign n571 = n95 & n570 ;
  assign n572 = n206 & n218 ;
  assign n573 = ~do_rnd_read_i_pad & ~do_seq_read_i_pad ;
  assign n574 = ~do_write_i_pad & n573 ;
  assign n575 = n186 & ~n574 ;
  assign n576 = n505 & n575 ;
  assign n577 = n572 & n576 ;
  assign n578 = ~n167 & ~n577 ;
  assign n579 = ~n571 & n578 ;
  assign n580 = n564 & n579 ;
  assign n581 = ~\bits_transfered_reg[0]/NET0131  & ~\bits_transfered_reg[1]/NET0131  ;
  assign n582 = ~\bits_transfered_reg[2]/NET0131  & \bits_transfered_reg[3]/NET0131  ;
  assign n583 = n581 & n582 ;
  assign n584 = \send_bit_reg/NET0131  & ~n583 ;
  assign n585 = ~n484 & ~n584 ;
  assign n586 = n106 & ~n585 ;
  assign n587 = ~\send_bit_reg/NET0131  & ~n176 ;
  assign n588 = \send_bit_reg/NET0131  & n583 ;
  assign n589 = n347 & ~n588 ;
  assign n590 = ~n587 & n589 ;
  assign n591 = n167 & n458 ;
  assign n592 = n136 & ~n583 ;
  assign n593 = ~n167 & ~n592 ;
  assign n594 = ~n341 & n593 ;
  assign n595 = \send_bit_reg/NET0131  & ~n594 ;
  assign n596 = ~n591 & ~n595 ;
  assign n597 = ~n590 & n596 ;
  assign n598 = ~n586 & n597 ;
  assign n599 = \bits_transfered_reg[0]/NET0131  & \bits_transfered_reg[1]/NET0131  ;
  assign n600 = \bits_transfered_reg[2]/NET0131  & n599 ;
  assign n601 = \bits_transfered_reg[3]/NET0131  & ~n600 ;
  assign n602 = \bits_transfered_reg[2]/NET0131  & ~\bits_transfered_reg[3]/NET0131  ;
  assign n603 = n599 & n602 ;
  assign n604 = ~n601 & ~n603 ;
  assign n605 = \send_bit_reg/NET0131  & ~n604 ;
  assign n606 = n191 & n605 ;
  assign n607 = ~n348 & n606 ;
  assign n608 = ~\send_bit_reg/NET0131  & ~n122 ;
  assign n609 = ~n122 & n604 ;
  assign n610 = n191 & n609 ;
  assign n611 = ~n608 & ~n610 ;
  assign n612 = \bits_transfered_reg[3]/NET0131  & ~n348 ;
  assign n613 = n611 & n612 ;
  assign n614 = ~n607 & ~n613 ;
  assign n615 = \bits_transfered_reg[3]/NET0131  & n165 ;
  assign n616 = ~n152 & ~n615 ;
  assign n617 = n81 & n433 ;
  assign n618 = \bits_transfered_reg[3]/NET0131  & \rec_bit_reg/NET0131  ;
  assign n619 = ~n617 & n618 ;
  assign n620 = \rec_bit_reg/NET0131  & ~n604 ;
  assign n621 = n617 & n620 ;
  assign n622 = ~n619 & ~n621 ;
  assign n623 = \bits_transfered_reg[3]/NET0131  & ~\send_nack_reg/NET0131  ;
  assign n624 = n154 & n623 ;
  assign n625 = ~n615 & ~n624 ;
  assign n626 = n622 & n625 ;
  assign n627 = ~n616 & ~n626 ;
  assign n628 = n614 & ~n627 ;
  assign n629 = n443 & ~n457 ;
  assign n630 = ~n506 & ~n629 ;
  assign n631 = ~n509 & n630 ;
  assign n632 = \tx_rx_state_reg[1]/NET0131  & ~n631 ;
  assign n633 = ~n115 & n450 ;
  assign n634 = ~n506 & ~n518 ;
  assign n635 = \send_start_reg/NET0131  & ~n634 ;
  assign n636 = ~n633 & ~n635 ;
  assign n637 = ~n632 & n636 ;
  assign n638 = n175 & n247 ;
  assign n639 = n95 & n638 ;
  assign n640 = n163 & n639 ;
  assign n641 = n206 & n566 ;
  assign n642 = ~n220 & ~n641 ;
  assign n643 = \rw_seq_state_reg[2]/NET0131  & ~n642 ;
  assign n644 = \rw_seq_state_reg[2]/NET0131  & ~n561 ;
  assign n645 = n491 & n644 ;
  assign n646 = ~n643 & ~n645 ;
  assign n647 = ~n640 & n646 ;
  assign n648 = n92 & n174 ;
  assign n649 = n95 & n648 ;
  assign n650 = n347 & n649 ;
  assign n651 = \rw_seq_state_reg[4]/NET0131  & n347 ;
  assign n652 = n491 & n651 ;
  assign n653 = ~n650 & ~n652 ;
  assign n654 = \rw_seq_state_reg[4]/NET0131  & ~n218 ;
  assign n655 = n165 & n654 ;
  assign n656 = n155 & n489 ;
  assign n657 = n152 & ~n656 ;
  assign n658 = ~n655 & ~n657 ;
  assign n659 = n653 & n658 ;
  assign n660 = ~n348 & n588 ;
  assign n661 = ~n167 & ~n341 ;
  assign n662 = ~\send_bit_reg/NET0131  & n80 ;
  assign n663 = n77 & n662 ;
  assign n664 = n89 & n663 ;
  assign n665 = n661 & n664 ;
  assign n666 = \rec_ack_reg/NET0131  & ~n665 ;
  assign n667 = ~n660 & ~n666 ;
  assign n668 = \adr_set_reg/NET0131  & ~n218 ;
  assign n669 = \adr_set_reg/NET0131  & n106 ;
  assign n670 = n92 & n106 ;
  assign n671 = n95 & n670 ;
  assign n672 = ~n669 & ~n671 ;
  assign n673 = ~n668 & n672 ;
  assign n674 = \bits_transfered_reg[1]/NET0131  & n122 ;
  assign n675 = ~n581 & ~n599 ;
  assign n676 = n138 & ~n675 ;
  assign n677 = n142 & n676 ;
  assign n678 = n190 & n677 ;
  assign n679 = \bits_transfered_reg[1]/NET0131  & \send_bit_reg/NET0131  ;
  assign n680 = ~n678 & n679 ;
  assign n681 = ~n674 & ~n680 ;
  assign n682 = \send_bit_reg/NET0131  & n675 ;
  assign n683 = n191 & n682 ;
  assign n684 = n681 & ~n683 ;
  assign n685 = ~n348 & ~n684 ;
  assign n686 = \bits_transfered_reg[1]/NET0131  & n165 ;
  assign n687 = ~n152 & ~n686 ;
  assign n688 = ~\bits_transfered_reg[1]/NET0131  & ~n617 ;
  assign n689 = n80 & ~n675 ;
  assign n690 = n77 & n689 ;
  assign n691 = n433 & n690 ;
  assign n692 = \rec_bit_reg/NET0131  & ~n691 ;
  assign n693 = ~n688 & n692 ;
  assign n694 = \bits_transfered_reg[1]/NET0131  & ~\send_nack_reg/NET0131  ;
  assign n695 = n154 & n694 ;
  assign n696 = ~n686 & ~n695 ;
  assign n697 = ~n693 & n696 ;
  assign n698 = ~n687 & ~n697 ;
  assign n699 = ~n685 & ~n698 ;
  assign n700 = ~\bits_transfered_reg[2]/NET0131  & ~n599 ;
  assign n701 = ~n600 & ~n700 ;
  assign n702 = \send_bit_reg/NET0131  & n701 ;
  assign n703 = n191 & n702 ;
  assign n704 = ~n348 & n703 ;
  assign n705 = ~n122 & ~n701 ;
  assign n706 = n191 & n705 ;
  assign n707 = ~n608 & ~n706 ;
  assign n708 = \bits_transfered_reg[2]/NET0131  & ~n348 ;
  assign n709 = n707 & n708 ;
  assign n710 = ~n704 & ~n709 ;
  assign n711 = \bits_transfered_reg[2]/NET0131  & n165 ;
  assign n712 = ~n152 & ~n711 ;
  assign n713 = \bits_transfered_reg[2]/NET0131  & \rec_bit_reg/NET0131  ;
  assign n714 = ~n617 & n713 ;
  assign n715 = \rec_bit_reg/NET0131  & n701 ;
  assign n716 = n617 & n715 ;
  assign n717 = ~n714 & ~n716 ;
  assign n718 = \bits_transfered_reg[2]/NET0131  & ~\send_nack_reg/NET0131  ;
  assign n719 = n154 & n718 ;
  assign n720 = ~n711 & ~n719 ;
  assign n721 = n717 & n720 ;
  assign n722 = ~n712 & ~n721 ;
  assign n723 = n710 & ~n722 ;
  assign n724 = \send_bit_reg/NET0131  & n138 ;
  assign n725 = n142 & n724 ;
  assign n726 = n190 & n725 ;
  assign n727 = ~n348 & n726 ;
  assign n728 = \rec_bit_reg/NET0131  & n151 ;
  assign n729 = n104 & n728 ;
  assign n730 = n617 & n729 ;
  assign n731 = ~n727 & ~n730 ;
  assign n732 = ~\bits_transfered_reg[0]/NET0131  & n731 ;
  assign n733 = ~n92 & ~n348 ;
  assign n734 = ~n726 & n733 ;
  assign n735 = ~n165 & ~n734 ;
  assign n736 = n152 & n155 ;
  assign n737 = \rec_bit_reg/NET0131  & n152 ;
  assign n738 = ~n617 & n737 ;
  assign n739 = ~n736 & ~n738 ;
  assign n740 = \bits_transfered_reg[0]/NET0131  & n739 ;
  assign n741 = n735 & n740 ;
  assign n742 = ~n732 & ~n741 ;
  assign n743 = ~n428 & ~n440 ;
  assign n744 = ~n115 & ~n743 ;
  assign n745 = ~n509 & ~n744 ;
  assign n746 = \tx_rx_state_reg[8]/NET0131  & ~n745 ;
  assign n747 = ~\send_bit_reg/NET0131  & n88 ;
  assign n748 = n86 & n747 ;
  assign n749 = n463 & n748 ;
  assign n750 = n115 & n428 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = \send_stop_reg/NET0131  & ~n751 ;
  assign n753 = ~n746 & ~n752 ;
  assign n754 = \tx_rx_state_reg[4]/NET0131  & n509 ;
  assign n755 = \send_bit_reg/NET0131  & n110 ;
  assign n756 = n114 & n755 ;
  assign n757 = n89 & ~n756 ;
  assign n758 = ~n461 & ~n757 ;
  assign n759 = ~\tx_rx_state_reg[4]/NET0131  & ~n115 ;
  assign n760 = ~n463 & ~n759 ;
  assign n761 = ~n758 & n760 ;
  assign n762 = n433 & ~n463 ;
  assign n763 = ~n761 & ~n762 ;
  assign n764 = ~n754 & n763 ;
  assign n765 = \tx_rx_state_reg[2]/NET0131  & n509 ;
  assign n766 = n100 & n749 ;
  assign n767 = ~n629 & ~n766 ;
  assign n768 = ~n765 & n767 ;
  assign n769 = ~n115 & ~n429 ;
  assign n770 = ~n762 & ~n769 ;
  assign n771 = ~n509 & n770 ;
  assign n772 = \tx_rx_state_reg[7]/NET0131  & ~n771 ;
  assign n773 = ~\send_ack_reg/NET0131  & n147 ;
  assign n774 = n110 & n773 ;
  assign n775 = n114 & n774 ;
  assign n776 = n433 & n775 ;
  assign n777 = ~n772 & ~n776 ;
  assign n778 = \tx_rx_state_reg[3]/NET0131  & n509 ;
  assign n779 = ~n89 & ~n450 ;
  assign n780 = ~\tx_rx_state_reg[3]/NET0131  & ~n115 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = ~n190 & ~n781 ;
  assign n783 = ~n467 & ~n782 ;
  assign n784 = ~n778 & ~n783 ;
  assign n785 = \tx_rx_state_reg[5]/NET0131  & n509 ;
  assign n786 = ~n115 & n461 ;
  assign n787 = \rec_bit_reg/NET0131  & ~\tx_rx_state_reg[5]/NET0131  ;
  assign n788 = ~n154 & ~n787 ;
  assign n789 = n110 & n788 ;
  assign n790 = n114 & n789 ;
  assign n791 = n433 & n790 ;
  assign n792 = ~n786 & ~n791 ;
  assign n793 = ~n785 & n792 ;
  assign n794 = ~\rec_bit_reg/NET0131  & ~\send_nack_reg/NET0131  ;
  assign n795 = n151 & n794 ;
  assign n796 = n104 & n795 ;
  assign n797 = \send_ack_reg/NET0131  & ~n796 ;
  assign n798 = n143 & n461 ;
  assign n799 = do_seq_read_i_pad & \send_ack_reg/NET0131  ;
  assign n800 = ~n798 & n799 ;
  assign n801 = ~n797 & ~n800 ;
  assign n802 = \rec_bit_reg/NET0131  & n583 ;
  assign n803 = ~\doing_read_reg/NET0131  & n151 ;
  assign n804 = n104 & n803 ;
  assign n805 = n802 & n804 ;
  assign n806 = n801 & ~n805 ;
  assign n807 = \send_bit_reg/NET0131  & ~\tx_rx_state_reg[6]/NET0131  ;
  assign n808 = ~n122 & ~n807 ;
  assign n809 = n110 & n808 ;
  assign n810 = n114 & n809 ;
  assign n811 = n190 & n810 ;
  assign n812 = ~\tx_rx_state_reg[6]/NET0131  & ~n811 ;
  assign n813 = ~n769 & ~n811 ;
  assign n814 = ~n509 & n813 ;
  assign n815 = ~n812 & ~n814 ;
  assign n816 = \doing_read_reg/NET0131  & ~n218 ;
  assign n817 = ~do_rnd_read_i_pad & ~\doing_read_reg/NET0131  ;
  assign n818 = ~do_write_i_pad & ~n817 ;
  assign n819 = n186 & n818 ;
  assign n820 = n505 & n819 ;
  assign n821 = n572 & n820 ;
  assign n822 = ~n816 & ~n821 ;
  assign n823 = n136 & n342 ;
  assign n824 = write_done_o_pad & ~n823 ;
  assign n825 = n92 & n136 ;
  assign n826 = n95 & n825 ;
  assign n827 = ~n824 & ~n826 ;
  assign n828 = ~\clk_gen_cnt_reg[0]/NET0131  & ~\clk_gen_cnt_reg[1]/NET0131  ;
  assign n829 = ~\clk_gen_cnt_reg[5]/NET0131  & ~\clk_gen_cnt_reg[6]/NET0131  ;
  assign n830 = n828 & n829 ;
  assign n831 = n452 & n830 ;
  assign n832 = n138 & n831 ;
  assign n833 = ~n457 & ~n832 ;
  assign n834 = ~n445 & ~n833 ;
  assign n835 = \doing_seq_read_reg/NET0131  & ~n218 ;
  assign n836 = n506 & n572 ;
  assign n837 = ~do_rnd_read_i_pad & do_seq_read_i_pad ;
  assign n838 = ~\doing_seq_read_reg/NET0131  & ~n837 ;
  assign n839 = ~do_write_i_pad & ~n838 ;
  assign n840 = n836 & n839 ;
  assign n841 = ~n835 & ~n840 ;
  assign n842 = n143 & n428 ;
  assign n843 = \send_nack_reg/NET0131  & ~n842 ;
  assign n844 = \rec_bit_reg/NET0131  & \send_nack_reg/NET0131  ;
  assign n845 = \doing_read_reg/NET0131  & \rec_bit_reg/NET0131  ;
  assign n846 = n583 & n845 ;
  assign n847 = ~n844 & ~n846 ;
  assign n848 = ~do_seq_read_i_pad & \send_ack_reg/NET0131  ;
  assign n849 = n794 & n848 ;
  assign n850 = n847 & ~n849 ;
  assign n851 = ~n843 & n850 ;
  assign n852 = \doing_write_reg/NET0131  & ~n218 ;
  assign n853 = do_write_i_pad & n186 ;
  assign n854 = n505 & n853 ;
  assign n855 = n572 & n854 ;
  assign n856 = ~n852 & ~n855 ;
  assign n857 = ~n445 & n832 ;
  assign n858 = ~\tx_rx_state_reg[8]/NET0131  & n184 ;
  assign n859 = ~\tx_rx_state_reg[4]/NET0131  & ~\tx_rx_state_reg[6]/NET0131  ;
  assign n860 = \tx_rx_state_reg[4]/NET0131  & \tx_rx_state_reg[6]/NET0131  ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = n858 & n861 ;
  assign n863 = n432 & n862 ;
  assign n864 = ~\send_ack_reg/NET0131  & ~\send_nack_reg/NET0131  ;
  assign n865 = ~\rec_bit_reg/NET0131  & ~n864 ;
  assign n866 = dat_rdy_o_pad & ~n865 ;
  assign n867 = ~n802 & ~n866 ;
  assign n868 = \rw_seq_state_reg[0]/NET0131  & n165 ;
  assign n869 = ~n218 & ~n868 ;
  assign n870 = ~n577 & ~n869 ;
  assign n871 = ~\rw_seq_state_reg[0]/NET0131  & ~n489 ;
  assign n872 = n122 & ~n162 ;
  assign n873 = ~\rw_seq_state_reg[0]/NET0131  & ~n155 ;
  assign n874 = n152 & ~n873 ;
  assign n875 = ~n872 & ~n874 ;
  assign n876 = ~n871 & ~n875 ;
  assign n877 = ~n870 & ~n876 ;
  assign n878 = \send_bit_reg/NET0131  & ~n561 ;
  assign n879 = \rw_seq_state_reg[0]/NET0131  & n878 ;
  assign n880 = \rw_seq_state_reg[0]/NET0131  & n566 ;
  assign n881 = ~n207 & n880 ;
  assign n882 = ~n879 & ~n881 ;
  assign n883 = ~\rw_seq_state_reg[0]/NET0131  & ~n492 ;
  assign n884 = \rec_ack_reg/NET0131  & n95 ;
  assign n885 = n101 & n247 ;
  assign n886 = n99 & n885 ;
  assign n887 = ~n884 & n886 ;
  assign n888 = ~n883 & n887 ;
  assign n889 = n882 & ~n888 ;
  assign n890 = n877 & n889 ;
  assign n891 = \tx_shift_reg_reg[0]/NET0131  & n163 ;
  assign n892 = ~n639 & n891 ;
  assign n893 = \adr_i[0]_pad  & n163 ;
  assign n894 = n639 & n893 ;
  assign n895 = ~n892 & ~n894 ;
  assign n896 = ~n136 & ~n220 ;
  assign n897 = \tx_shift_reg_reg[0]/NET0131  & ~n896 ;
  assign n898 = n92 & ~n206 ;
  assign n899 = n95 & n898 ;
  assign n900 = ~\tx_shift_reg_reg[0]/NET0131  & ~n899 ;
  assign n901 = ~\dat_i[0]_pad  & \doing_write_reg/NET0131  ;
  assign n902 = n92 & n901 ;
  assign n903 = n95 & n902 ;
  assign n904 = n106 & ~n903 ;
  assign n905 = ~n900 & n904 ;
  assign n906 = ~n897 & ~n905 ;
  assign n907 = n895 & n906 ;
  assign n908 = ~\clk_gen_cnt_reg[6]/NET0131  & ~n542 ;
  assign n909 = n522 & ~n548 ;
  assign n910 = ~n908 & n909 ;
  assign n911 = ~n506 & ~n509 ;
  assign n912 = ~\clk_gen_cnt_reg[0]/NET0131  & ~n911 ;
  assign n913 = ~n511 & n522 ;
  assign n914 = ~n912 & n913 ;
  assign n915 = \dat_i[6]_pad  & \doing_write_reg/NET0131  ;
  assign n916 = n95 & n915 ;
  assign n917 = n106 & n916 ;
  assign n918 = \tx_shift_reg_reg[6]/NET0131  & n106 ;
  assign n919 = ~n207 & n918 ;
  assign n920 = ~n917 & ~n919 ;
  assign n921 = ~\adr_i[6]_pad  & ~n174 ;
  assign n922 = n95 & n921 ;
  assign n923 = \tx_shift_reg_reg[6]/NET0131  & n347 ;
  assign n924 = ~n174 & n347 ;
  assign n925 = n95 & n924 ;
  assign n926 = ~n923 & ~n925 ;
  assign n927 = ~n922 & ~n926 ;
  assign n928 = n920 & ~n927 ;
  assign n929 = n92 & ~n928 ;
  assign n930 = ~n167 & ~n220 ;
  assign n931 = \tx_shift_reg_reg[6]/NET0131  & ~n930 ;
  assign n932 = \tx_shift_reg_reg[6]/NET0131  & n92 ;
  assign n933 = ~n136 & n932 ;
  assign n934 = ~\tx_shift_reg_reg[5]/NET0131  & ~n933 ;
  assign n935 = n726 & n934 ;
  assign n936 = \tx_shift_reg_reg[6]/NET0131  & ~n92 ;
  assign n937 = \tx_shift_reg_reg[6]/NET0131  & n135 ;
  assign n938 = n134 & n937 ;
  assign n939 = ~n936 & ~n938 ;
  assign n940 = ~n726 & n939 ;
  assign n941 = ~n348 & ~n940 ;
  assign n942 = ~n935 & n941 ;
  assign n943 = ~n931 & ~n942 ;
  assign n944 = ~n929 & n943 ;
  assign n945 = n92 & ~n205 ;
  assign n946 = ~\doing_write_reg/NET0131  & n945 ;
  assign n947 = n95 & n946 ;
  assign n948 = ~\send_start_reg/NET0131  & ~n947 ;
  assign n949 = n106 & ~n948 ;
  assign n950 = n163 & n458 ;
  assign n951 = \send_start_reg/NET0131  & ~n950 ;
  assign n952 = ~n577 & ~n951 ;
  assign n953 = ~n949 & n952 ;
  assign n954 = \rec_bit_reg/NET0131  & n163 ;
  assign n955 = n174 & n248 ;
  assign n956 = n163 & n955 ;
  assign n957 = n95 & n956 ;
  assign n958 = ~n954 & ~n957 ;
  assign n959 = n152 & n583 ;
  assign n960 = \rec_bit_reg/NET0131  & ~n959 ;
  assign n961 = n796 & n799 ;
  assign n962 = n798 & n961 ;
  assign n963 = ~n960 & ~n962 ;
  assign n964 = n958 & n963 ;
  assign n965 = \tx_rx_state_reg[0]/NET0131  & n509 ;
  assign n966 = ~\send_start_reg/NET0131  & \tx_rx_state_reg[0]/NET0131  ;
  assign n967 = n506 & n966 ;
  assign n968 = ~n965 & ~n967 ;
  assign n969 = n115 & n433 ;
  assign n970 = \rec_bit_reg/NET0131  & ~\tx_rx_state_reg[0]/NET0131  ;
  assign n971 = ~n865 & ~n970 ;
  assign n972 = n969 & n971 ;
  assign n973 = \send_bit_reg/NET0131  & ~\tx_rx_state_reg[0]/NET0131  ;
  assign n974 = ~n92 & ~n973 ;
  assign n975 = n110 & n974 ;
  assign n976 = n114 & n975 ;
  assign n977 = n190 & n976 ;
  assign n978 = ~\send_stop_reg/NET0131  & n247 ;
  assign n979 = n88 & n978 ;
  assign n980 = n86 & n979 ;
  assign n981 = n463 & n980 ;
  assign n982 = ~n977 & ~n981 ;
  assign n983 = ~n972 & n982 ;
  assign n984 = ~\tx_rx_state_reg[0]/NET0131  & ~n115 ;
  assign n985 = n428 & ~n488 ;
  assign n986 = \rec_bit_reg/NET0131  & n110 ;
  assign n987 = n114 & n986 ;
  assign n988 = n461 & ~n987 ;
  assign n989 = ~n985 & ~n988 ;
  assign n990 = ~n984 & ~n989 ;
  assign n991 = ~\tx_rx_state_reg[0]/NET0131  & ~n457 ;
  assign n992 = \send_start_reg/NET0131  & n451 ;
  assign n993 = n456 & n992 ;
  assign n994 = n443 & ~n993 ;
  assign n995 = ~n991 & n994 ;
  assign n996 = n469 & ~n995 ;
  assign n997 = ~n990 & n996 ;
  assign n998 = n983 & n997 ;
  assign n999 = n968 & n998 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g4613/_2_  = ~n172 ;
  assign \g4620/_0_  = ~n227 ;
  assign \g4621/_0_  = ~n268 ;
  assign \g4627/_0_  = ~n304 ;
  assign \g4628/_0_  = ~n340 ;
  assign \g4630/_0_  = ~n352 ;
  assign \g4631/_0_  = ~n388 ;
  assign \g4632/_0_  = ~n423 ;
  assign \g4657/_0_  = ~n482 ;
  assign \g4672/_0_  = ~n504 ;
  assign \g4673/_0_  = n524 ;
  assign \g4674/_0_  = n529 ;
  assign \g4675/_0_  = n535 ;
  assign \g4676/_0_  = n541 ;
  assign \g4677/_0_  = n545 ;
  assign \g4679/_0_  = n554 ;
  assign \g4680/_0_  = n558 ;
  assign \g4684/_0_  = ~n580 ;
  assign \g4685/_0_  = ~n598 ;
  assign \g4696/_0_  = ~n628 ;
  assign \g4697/_0_  = ~n637 ;
  assign \g4699/_0_  = ~n647 ;
  assign \g4700/_0_  = ~n659 ;
  assign \g4743/_0_  = ~n667 ;
  assign \g4768/_0_  = ~n673 ;
  assign \g4769/_0_  = ~n699 ;
  assign \g4770/_0_  = ~n723 ;
  assign \g4771/_0_  = n742 ;
  assign \g4785/_0_  = ~n753 ;
  assign \g4790/_0_  = ~n764 ;
  assign \g4792/_0_  = ~n768 ;
  assign \g4810/_0_  = ~n777 ;
  assign \g4830/_0_  = ~n784 ;
  assign \g4831/_0_  = ~n793 ;
  assign \g4870/_0_  = ~n806 ;
  assign \g4891/_0_  = n815 ;
  assign \g4898/_0_  = ~n822 ;
  assign \g4903/_0_  = ~n827 ;
  assign \g4951/_2__syn_2  = n834 ;
  assign \g4991/_3_  = ~n841 ;
  assign \g5054/_0_  = ~n851 ;
  assign \g5064/_0_  = ~n856 ;
  assign \g5068/u3_syn_4  = n730 ;
  assign \g5085/_1_  = ~n857 ;
  assign \g5290/_0_  = n863 ;
  assign \g5524/_0_  = ~n867 ;
  assign \g5574/_2_  = n152 ;
  assign \g57/_0_  = ~n890 ;
  assign \g6488/_0_  = ~n907 ;
  assign \g6585/_0_  = n910 ;
  assign \g6602/_0_  = n914 ;
  assign \g6658/_0_  = ~n944 ;
  assign \g6720/_0_  = ~n953 ;
  assign \g6767/_0_  = ~n964 ;
  assign \g6827/_0_  = ~n999 ;
endmodule
