module top( \a0_pad  , a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , \h0_pad  , h_pad , \i0_pad  , i_pad , \j0_pad  , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , \u0_pad  , \v0_pad  , \w0_pad  , \x0_pad  , \y0_pad  , \z0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output \u0_pad  ;
  output \v0_pad  ;
  output \w0_pad  ;
  output \x0_pad  ;
  output \y0_pad  ;
  output \z0_pad  ;
  wire n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 ;
  assign n36 = ~r_pad & ~u_pad ;
  assign n37 = r_pad & u_pad ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = q_pad & ~n38 ;
  assign n40 = ~p_pad & ~q_pad ;
  assign n41 = ~s_pad & ~n40 ;
  assign n42 = ~n39 & n41 ;
  assign n43 = q_pad & v_pad ;
  assign n44 = ~n36 & n43 ;
  assign n45 = q_pad & ~v_pad ;
  assign n46 = n36 & n45 ;
  assign n47 = ~n44 & ~n46 ;
  assign n48 = ~o_pad & ~q_pad ;
  assign n49 = ~s_pad & ~n48 ;
  assign n50 = n47 & n49 ;
  assign n51 = ~v_pad & n36 ;
  assign n52 = q_pad & w_pad ;
  assign n53 = ~n51 & n52 ;
  assign n54 = q_pad & ~w_pad ;
  assign n55 = n51 & n54 ;
  assign n56 = ~n53 & ~n55 ;
  assign n57 = ~n_pad & ~q_pad ;
  assign n58 = ~s_pad & ~n57 ;
  assign n59 = n56 & n58 ;
  assign n60 = ~v_pad & ~w_pad ;
  assign n61 = n36 & n60 ;
  assign n62 = q_pad & x_pad ;
  assign n63 = ~n61 & n62 ;
  assign n64 = q_pad & ~x_pad ;
  assign n65 = n61 & n64 ;
  assign n66 = ~n63 & ~n65 ;
  assign n67 = ~m_pad & ~q_pad ;
  assign n68 = ~s_pad & ~n67 ;
  assign n69 = n66 & n68 ;
  assign n70 = ~x_pad & n61 ;
  assign n71 = q_pad & y_pad ;
  assign n72 = ~n70 & n71 ;
  assign n73 = q_pad & ~y_pad ;
  assign n74 = ~x_pad & n73 ;
  assign n75 = n61 & n74 ;
  assign n76 = ~l_pad & ~q_pad ;
  assign n77 = ~s_pad & ~n76 ;
  assign n78 = ~n75 & n77 ;
  assign n79 = ~n72 & n78 ;
  assign n80 = ~x_pad & ~y_pad ;
  assign n81 = n61 & n80 ;
  assign n82 = q_pad & z_pad ;
  assign n83 = ~n81 & n82 ;
  assign n84 = q_pad & ~z_pad ;
  assign n85 = n80 & n84 ;
  assign n86 = n61 & n85 ;
  assign n87 = ~k_pad & ~q_pad ;
  assign n88 = ~s_pad & ~n87 ;
  assign n89 = ~n86 & n88 ;
  assign n90 = ~n83 & n89 ;
  assign n91 = ~x_pad & ~z_pad ;
  assign n92 = ~y_pad & n91 ;
  assign n93 = n61 & n92 ;
  assign n94 = ~\a0_pad  & q_pad ;
  assign n95 = ~j_pad & ~q_pad ;
  assign n96 = ~s_pad & ~n95 ;
  assign n97 = ~n94 & n96 ;
  assign n98 = n93 & n97 ;
  assign n99 = \a0_pad  & q_pad ;
  assign n100 = n96 & ~n99 ;
  assign n101 = ~n93 & n100 ;
  assign n102 = ~n98 & ~n101 ;
  assign n103 = ~\a0_pad  & ~y_pad ;
  assign n104 = n91 & n103 ;
  assign n105 = n61 & n104 ;
  assign n106 = ~\b0_pad  & q_pad ;
  assign n107 = ~i_pad & ~q_pad ;
  assign n108 = ~s_pad & ~n107 ;
  assign n109 = ~n106 & n108 ;
  assign n110 = n105 & n109 ;
  assign n111 = \b0_pad  & q_pad ;
  assign n112 = n108 & ~n111 ;
  assign n113 = ~n105 & n112 ;
  assign n114 = ~n110 & ~n113 ;
  assign n115 = ~\a0_pad  & ~\b0_pad  ;
  assign n116 = n93 & n115 ;
  assign n117 = \c0_pad  & q_pad ;
  assign n118 = ~n116 & n117 ;
  assign n119 = ~\c0_pad  & q_pad ;
  assign n120 = n115 & n119 ;
  assign n121 = n93 & n120 ;
  assign n122 = ~h_pad & ~q_pad ;
  assign n123 = ~s_pad & ~n122 ;
  assign n124 = ~n121 & n123 ;
  assign n125 = ~n118 & n124 ;
  assign n126 = ~\a0_pad  & ~\c0_pad  ;
  assign n127 = ~\b0_pad  & n126 ;
  assign n128 = n93 & n127 ;
  assign n129 = \d0_pad  & q_pad ;
  assign n130 = ~n128 & n129 ;
  assign n131 = ~\d0_pad  & q_pad ;
  assign n132 = n127 & n131 ;
  assign n133 = n93 & n132 ;
  assign n134 = ~g_pad & ~q_pad ;
  assign n135 = ~s_pad & ~n134 ;
  assign n136 = ~n133 & n135 ;
  assign n137 = ~n130 & n136 ;
  assign n138 = ~\d0_pad  & n127 ;
  assign n139 = n93 & n138 ;
  assign n140 = \e0_pad  & q_pad ;
  assign n141 = ~n139 & n140 ;
  assign n142 = ~\e0_pad  & q_pad ;
  assign n143 = ~\d0_pad  & n142 ;
  assign n144 = n127 & n143 ;
  assign n145 = n93 & n144 ;
  assign n146 = ~f_pad & ~q_pad ;
  assign n147 = ~s_pad & ~n146 ;
  assign n148 = ~n145 & n147 ;
  assign n149 = ~n141 & n148 ;
  assign n150 = ~\d0_pad  & ~\e0_pad  ;
  assign n151 = n127 & n150 ;
  assign n152 = n93 & n151 ;
  assign n153 = \f0_pad  & q_pad ;
  assign n154 = ~n152 & n153 ;
  assign n155 = ~\f0_pad  & q_pad ;
  assign n156 = n150 & n155 ;
  assign n157 = n127 & n156 ;
  assign n158 = n93 & n157 ;
  assign n159 = ~e_pad & ~q_pad ;
  assign n160 = ~s_pad & ~n159 ;
  assign n161 = ~n158 & n160 ;
  assign n162 = ~n154 & n161 ;
  assign n163 = ~\d0_pad  & ~\f0_pad  ;
  assign n164 = ~\e0_pad  & n163 ;
  assign n165 = n127 & n164 ;
  assign n166 = n93 & n165 ;
  assign n167 = ~\g0_pad  & q_pad ;
  assign n168 = ~d_pad & ~q_pad ;
  assign n169 = ~s_pad & ~n168 ;
  assign n170 = ~n167 & n169 ;
  assign n171 = n166 & n170 ;
  assign n172 = \g0_pad  & q_pad ;
  assign n173 = n169 & ~n172 ;
  assign n174 = ~n166 & n173 ;
  assign n175 = ~n171 & ~n174 ;
  assign n176 = ~\g0_pad  & n166 ;
  assign n177 = \h0_pad  & q_pad ;
  assign n178 = ~n176 & n177 ;
  assign n179 = ~\h0_pad  & q_pad ;
  assign n180 = ~\g0_pad  & n179 ;
  assign n181 = n166 & n180 ;
  assign n182 = ~c_pad & ~q_pad ;
  assign n183 = ~s_pad & ~n182 ;
  assign n184 = ~n181 & n183 ;
  assign n185 = ~n178 & n184 ;
  assign n186 = ~\g0_pad  & ~\h0_pad  ;
  assign n187 = n166 & n186 ;
  assign n188 = \i0_pad  & q_pad ;
  assign n189 = ~n187 & n188 ;
  assign n190 = ~\i0_pad  & q_pad ;
  assign n191 = n186 & n190 ;
  assign n192 = n166 & n191 ;
  assign n193 = ~b_pad & ~q_pad ;
  assign n194 = ~s_pad & ~n193 ;
  assign n195 = ~n192 & n194 ;
  assign n196 = ~n189 & n195 ;
  assign n197 = ~\g0_pad  & ~\i0_pad  ;
  assign n198 = ~\h0_pad  & n197 ;
  assign n199 = n166 & n198 ;
  assign n200 = \j0_pad  & q_pad ;
  assign n201 = ~n199 & n200 ;
  assign n202 = ~\j0_pad  & q_pad ;
  assign n203 = n198 & n202 ;
  assign n204 = n166 & n203 ;
  assign n205 = ~a_pad & ~q_pad ;
  assign n206 = ~s_pad & ~n205 ;
  assign n207 = ~n204 & n206 ;
  assign n208 = ~n201 & n207 ;
  assign \k0_pad  = ~n42 ;
  assign \l0_pad  = ~n50 ;
  assign \m0_pad  = ~n59 ;
  assign \n0_pad  = ~n69 ;
  assign \o0_pad  = ~n79 ;
  assign \p0_pad  = ~n90 ;
  assign \q0_pad  = n102 ;
  assign \r0_pad  = n114 ;
  assign \s0_pad  = ~n125 ;
  assign \t0_pad  = ~n137 ;
  assign \u0_pad  = ~n149 ;
  assign \v0_pad  = ~n162 ;
  assign \w0_pad  = n175 ;
  assign \x0_pad  = ~n185 ;
  assign \y0_pad  = ~n196 ;
  assign \z0_pad  = ~n208 ;
endmodule
