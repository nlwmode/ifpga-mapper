module top (\d_in_reg[0]/NET0131 , \d_in_reg[1]/NET0131 , \d_in_reg[2]/NET0131 , \d_in_reg[3]/NET0131 , \d_in_reg[4]/NET0131 , \d_in_reg[5]/NET0131 , \d_in_reg[6]/NET0131 , \d_in_reg[7]/NET0131 , \d_in_reg[8]/NET0131 , \d_out_reg[0]/NET0131 , \d_out_reg[1]/NET0131 , \d_out_reg[2]/NET0131 , \d_out_reg[3]/NET0131 , \d_out_reg[4]/NET0131 , \d_out_reg[5]/NET0131 , \d_out_reg[6]/NET0131 , \d_out_reg[7]/NET0131 , \old_reg[0]/NET0131 , \old_reg[1]/NET0131 , \old_reg[2]/NET0131 , \old_reg[3]/NET0131 , \old_reg[4]/NET0131 , \old_reg[5]/NET0131 , \old_reg[6]/NET0131 , \old_reg[7]/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , x_pad, y_pad, \_al_n0 , \_al_n1 , \g1026/_0_ , \g1035/_0_ , \g41/_0_ , \g708/_0_ , \g709/_0_ , \g711/_0_ , \g712/_0_ , \g714/_0_ , \g716/_0_ , \g718/_0_ , \g728/_0_ , \g770/_0_ , \g771/_0_ , \g772/_0_ , \g773/_0_ , \g774/_0_ , \g775/_0_ , \g776/_0_ , \g777/_0_ , \g782/_0_ , \g783/_0_ , \g784/_0_ , \g785/_0_ , \g786/_0_ , \g787/_0_ , \g788/_0_ , \g789/_0_ , \g806/_0_ );
	input \d_in_reg[0]/NET0131  ;
	input \d_in_reg[1]/NET0131  ;
	input \d_in_reg[2]/NET0131  ;
	input \d_in_reg[3]/NET0131  ;
	input \d_in_reg[4]/NET0131  ;
	input \d_in_reg[5]/NET0131  ;
	input \d_in_reg[6]/NET0131  ;
	input \d_in_reg[7]/NET0131  ;
	input \d_in_reg[8]/NET0131  ;
	input \d_out_reg[0]/NET0131  ;
	input \d_out_reg[1]/NET0131  ;
	input \d_out_reg[2]/NET0131  ;
	input \d_out_reg[3]/NET0131  ;
	input \d_out_reg[4]/NET0131  ;
	input \d_out_reg[5]/NET0131  ;
	input \d_out_reg[6]/NET0131  ;
	input \d_out_reg[7]/NET0131  ;
	input \old_reg[0]/NET0131  ;
	input \old_reg[1]/NET0131  ;
	input \old_reg[2]/NET0131  ;
	input \old_reg[3]/NET0131  ;
	input \old_reg[4]/NET0131  ;
	input \old_reg[5]/NET0131  ;
	input \old_reg[6]/NET0131  ;
	input \old_reg[7]/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input x_pad ;
	input y_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1026/_0_  ;
	output \g1035/_0_  ;
	output \g41/_0_  ;
	output \g708/_0_  ;
	output \g709/_0_  ;
	output \g711/_0_  ;
	output \g712/_0_  ;
	output \g714/_0_  ;
	output \g716/_0_  ;
	output \g718/_0_  ;
	output \g728/_0_  ;
	output \g770/_0_  ;
	output \g771/_0_  ;
	output \g772/_0_  ;
	output \g773/_0_  ;
	output \g774/_0_  ;
	output \g775/_0_  ;
	output \g776/_0_  ;
	output \g777/_0_  ;
	output \g782/_0_  ;
	output \g783/_0_  ;
	output \g784/_0_  ;
	output \g785/_0_  ;
	output \g786/_0_  ;
	output \g787/_0_  ;
	output \g788/_0_  ;
	output \g789/_0_  ;
	output \g806/_0_  ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\d_in_reg[0]/NET0131 ,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\d_in_reg[3]/NET0131 ,
		\old_reg[2]/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\d_in_reg[3]/NET0131 ,
		\old_reg[2]/NET0131 ,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\d_in_reg[2]/NET0131 ,
		\old_reg[1]/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\d_in_reg[2]/NET0131 ,
		\old_reg[1]/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w34_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\d_in_reg[1]/NET0131 ,
		\old_reg[0]/NET0131 ,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\d_in_reg[1]/NET0131 ,
		\old_reg[0]/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\d_in_reg[4]/NET0131 ,
		\old_reg[3]/NET0131 ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\d_in_reg[4]/NET0131 ,
		\old_reg[3]/NET0131 ,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\d_in_reg[6]/NET0131 ,
		\old_reg[5]/NET0131 ,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\d_in_reg[6]/NET0131 ,
		\old_reg[5]/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\d_in_reg[5]/NET0131 ,
		\old_reg[4]/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\d_in_reg[5]/NET0131 ,
		\old_reg[4]/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\d_in_reg[8]/NET0131 ,
		\old_reg[7]/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\d_in_reg[8]/NET0131 ,
		\old_reg[7]/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\d_in_reg[7]/NET0131 ,
		\old_reg[6]/NET0131 ,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\d_in_reg[7]/NET0131 ,
		\old_reg[6]/NET0131 ,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w32_,
		_w33_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w43_,
		_w44_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w36_,
		_w39_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w42_,
		_w47_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w50_,
		_w53_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w56_,
		_w57_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\d_in_reg[1]/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\d_out_reg[0]/NET0131 ,
		_w62_,
		_w64_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w31_,
		_w63_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w64_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[1]/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\d_in_reg[0]/NET0131 ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\d_out_reg[1]/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\d_in_reg[0]/NET0131 ,
		_w67_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\d_in_reg[0]/NET0131 ,
		_w30_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\d_in_reg[0]/NET0131 ,
		_w70_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w73_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\d_out_reg[0]/NET0131 ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w69_,
		_w72_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w66_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\d_in_reg[2]/NET0131 ,
		_w62_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		\d_out_reg[1]/NET0131 ,
		_w62_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		_w31_,
		_w82_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w67_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\d_out_reg[2]/NET0131 ,
		_w71_,
		_w88_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\d_out_reg[1]/NET0131 ,
		_w77_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w87_,
		_w88_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w85_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\d_out_reg[7]/NET0131 ,
		_w77_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w67_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\d_in_reg[8]/NET0131 ,
		_w62_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\d_out_reg[7]/NET0131 ,
		_w62_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w31_,
		_w96_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w93_,
		_w95_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w70_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		x_pad,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\stato_reg[1]/NET0131 ,
		_w62_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w104_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\d_in_reg[4]/NET0131 ,
		_w62_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		\d_out_reg[3]/NET0131 ,
		_w62_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w31_,
		_w109_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\d_out_reg[3]/NET0131 ,
		_w76_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[3]/NET0131 ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[4]/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w67_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\d_out_reg[4]/NET0131 ,
		_w71_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w113_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w112_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\d_in_reg[5]/NET0131 ,
		_w62_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\d_out_reg[4]/NET0131 ,
		_w62_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w31_,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w67_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\d_out_reg[5]/NET0131 ,
		_w71_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\d_out_reg[4]/NET0131 ,
		_w77_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w127_,
		_w128_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w125_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\d_in_reg[6]/NET0131 ,
		_w62_,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\d_out_reg[5]/NET0131 ,
		_w62_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		_w31_,
		_w133_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w67_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\d_out_reg[6]/NET0131 ,
		_w71_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		\d_out_reg[5]/NET0131 ,
		_w77_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w138_,
		_w139_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w136_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\d_in_reg[7]/NET0131 ,
		_w62_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\d_out_reg[6]/NET0131 ,
		_w62_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		_w31_,
		_w144_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[7]/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w67_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\d_out_reg[7]/NET0131 ,
		_w71_,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\d_out_reg[6]/NET0131 ,
		_w77_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w149_,
		_w150_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w147_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w70_,
		_w114_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\d_out_reg[2]/NET0131 ,
		_w77_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\d_in_reg[0]/NET0131 ,
		_w67_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\d_in_reg[3]/NET0131 ,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\d_in_reg[3]/NET0131 ,
		_w62_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		\d_out_reg[2]/NET0131 ,
		_w62_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w31_,
		_w159_,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w155_,
		_w158_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w156_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w162_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w71_,
		_w107_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		_w31_,
		_w62_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\d_in_reg[0]/NET0131 ,
		y_pad,
		_w168_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		_w67_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\d_out_reg[0]/NET0131 ,
		_w71_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w167_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\d_in_reg[2]/NET0131 ,
		_w103_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\d_in_reg[7]/NET0131 ,
		_w103_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\d_in_reg[8]/NET0131 ,
		_w103_,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\d_in_reg[1]/NET0131 ,
		_w103_,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\d_in_reg[6]/NET0131 ,
		_w103_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\d_in_reg[3]/NET0131 ,
		_w103_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		\d_in_reg[4]/NET0131 ,
		_w103_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\d_in_reg[5]/NET0131 ,
		_w103_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[5]/NET0131 ,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w137_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\stato_reg[0]/NET0131 ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\old_reg[5]/NET0131 ,
		_w70_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[6]/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w148_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\stato_reg[0]/NET0131 ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\old_reg[6]/NET0131 ,
		_w70_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[7]/NET0131 ,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w94_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\stato_reg[0]/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\old_reg[7]/NET0131 ,
		_w70_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w193_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[0]/NET0131 ,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w68_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\stato_reg[0]/NET0131 ,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\old_reg[0]/NET0131 ,
		_w70_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w198_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[1]/NET0131 ,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w86_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\stato_reg[0]/NET0131 ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\old_reg[1]/NET0131 ,
		_w70_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\d_in_reg[3]/NET0131 ,
		_w105_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\old_reg[2]/NET0131 ,
		_w103_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[3]/NET0131 ,
		_w209_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w115_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\stato_reg[0]/NET0131 ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\old_reg[3]/NET0131 ,
		_w70_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[4]/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w126_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\stato_reg[0]/NET0131 ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		\old_reg[4]/NET0131 ,
		_w70_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w30_,
		_w70_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w157_,
		_w219_,
		_w220_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1026/_0_  = _w81_ ;
	assign \g1035/_0_  = _w92_ ;
	assign \g41/_0_  = _w101_ ;
	assign \g708/_0_  = _w108_ ;
	assign \g709/_0_  = _w121_ ;
	assign \g711/_0_  = _w132_ ;
	assign \g712/_0_  = _w143_ ;
	assign \g714/_0_  = _w154_ ;
	assign \g716/_0_  = _w165_ ;
	assign \g718/_0_  = _w166_ ;
	assign \g728/_0_  = _w172_ ;
	assign \g770/_0_  = _w173_ ;
	assign \g771/_0_  = _w174_ ;
	assign \g772/_0_  = _w175_ ;
	assign \g773/_0_  = _w176_ ;
	assign \g774/_0_  = _w177_ ;
	assign \g775/_0_  = _w178_ ;
	assign \g776/_0_  = _w179_ ;
	assign \g777/_0_  = _w180_ ;
	assign \g782/_0_  = _w185_ ;
	assign \g783/_0_  = _w190_ ;
	assign \g784/_0_  = _w195_ ;
	assign \g785/_0_  = _w200_ ;
	assign \g786/_0_  = _w205_ ;
	assign \g787/_0_  = _w208_ ;
	assign \g788/_0_  = _w213_ ;
	assign \g789/_0_  = _w218_ ;
	assign \g806/_0_  = _w220_ ;
endmodule;