module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  output m_pad ;
  output n_pad ;
  wire n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 ;
  assign n24 = a_pad & ~i_pad ;
  assign n23 = b_pad & i_pad ;
  assign n25 = ~j_pad & ~n23 ;
  assign n26 = ~n24 & n25 ;
  assign n28 = c_pad & ~i_pad ;
  assign n27 = d_pad & i_pad ;
  assign n29 = j_pad & ~n27 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = ~n26 & ~n30 ;
  assign n32 = ~k_pad & ~n31 ;
  assign n14 = e_pad & ~i_pad ;
  assign n13 = f_pad & i_pad ;
  assign n15 = ~j_pad & ~n13 ;
  assign n16 = ~n14 & n15 ;
  assign n18 = g_pad & ~i_pad ;
  assign n17 = h_pad & i_pad ;
  assign n19 = j_pad & ~n17 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = ~n16 & ~n20 ;
  assign n22 = k_pad & ~n21 ;
  assign n33 = ~l_pad & ~n22 ;
  assign n34 = ~n32 & n33 ;
  assign m_pad = n34 ;
  assign n_pad = ~n34 ;
endmodule
