module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \a0_pad , \b0_pad , \c0_pad , \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad );
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a0_pad  ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		a_pad,
		i_pad,
		_w18_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		i_pad,
		s_pad,
		_w19_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w18_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		b_pad,
		i_pad,
		_w21_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		i_pad,
		t_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w21_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		c_pad,
		i_pad,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		i_pad,
		u_pad,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w24_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		d_pad,
		i_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		i_pad,
		v_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		e_pad,
		i_pad,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		i_pad,
		w_pad,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w30_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		f_pad,
		i_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		i_pad,
		x_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		g_pad,
		i_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		i_pad,
		y_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w36_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		h_pad,
		i_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		i_pad,
		z_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w39_,
		_w40_,
		_w41_
	);
	assign \a0_pad  = _w20_ ;
	assign \b0_pad  = _w23_ ;
	assign \c0_pad  = _w26_ ;
	assign \d0_pad  = _w29_ ;
	assign \e0_pad  = _w32_ ;
	assign \f0_pad  = _w35_ ;
	assign \g0_pad  = _w38_ ;
	assign \h0_pad  = _w41_ ;
endmodule;