module top (\dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4] , \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9] , \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] , \dest_x[14] , \dest_x[15] , \dest_x[16] , \dest_x[17] , \dest_x[18] , \dest_x[19] , \dest_x[20] , \dest_x[21] , \dest_x[22] , \dest_x[23] , \dest_x[24] , \dest_x[25] , \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] , \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] , \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] , \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] , \dest_y[14] , \dest_y[15] , \dest_y[16] , \dest_y[17] , \dest_y[18] , \dest_y[19] , \dest_y[20] , \dest_y[21] , \dest_y[22] , \dest_y[23] , \dest_y[24] , \dest_y[25] , \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] , \outport[0] , \outport[1] , \outport[2] , \outport[3] , \outport[4] , \outport[5] , \outport[6] , \outport[7] , \outport[8] , \outport[9] , \outport[10] , \outport[11] , \outport[12] , \outport[13] , \outport[14] , \outport[15] , \outport[16] , \outport[17] , \outport[18] , \outport[19] , \outport[20] , \outport[21] , \outport[22] , \outport[23] , \outport[24] , \outport[25] , \outport[26] , \outport[27] , \outport[28] , \outport[29] );
	input \dest_x[0]  ;
	input \dest_x[1]  ;
	input \dest_x[2]  ;
	input \dest_x[3]  ;
	input \dest_x[4]  ;
	input \dest_x[5]  ;
	input \dest_x[6]  ;
	input \dest_x[7]  ;
	input \dest_x[8]  ;
	input \dest_x[9]  ;
	input \dest_x[10]  ;
	input \dest_x[11]  ;
	input \dest_x[12]  ;
	input \dest_x[13]  ;
	input \dest_x[14]  ;
	input \dest_x[15]  ;
	input \dest_x[16]  ;
	input \dest_x[17]  ;
	input \dest_x[18]  ;
	input \dest_x[19]  ;
	input \dest_x[20]  ;
	input \dest_x[21]  ;
	input \dest_x[22]  ;
	input \dest_x[23]  ;
	input \dest_x[24]  ;
	input \dest_x[25]  ;
	input \dest_x[26]  ;
	input \dest_x[27]  ;
	input \dest_x[28]  ;
	input \dest_x[29]  ;
	input \dest_y[0]  ;
	input \dest_y[1]  ;
	input \dest_y[2]  ;
	input \dest_y[3]  ;
	input \dest_y[4]  ;
	input \dest_y[5]  ;
	input \dest_y[6]  ;
	input \dest_y[7]  ;
	input \dest_y[8]  ;
	input \dest_y[9]  ;
	input \dest_y[10]  ;
	input \dest_y[11]  ;
	input \dest_y[12]  ;
	input \dest_y[13]  ;
	input \dest_y[14]  ;
	input \dest_y[15]  ;
	input \dest_y[16]  ;
	input \dest_y[17]  ;
	input \dest_y[18]  ;
	input \dest_y[19]  ;
	input \dest_y[20]  ;
	input \dest_y[21]  ;
	input \dest_y[22]  ;
	input \dest_y[23]  ;
	input \dest_y[24]  ;
	input \dest_y[25]  ;
	input \dest_y[26]  ;
	input \dest_y[27]  ;
	input \dest_y[28]  ;
	input \dest_y[29]  ;
	output \outport[0]  ;
	output \outport[1]  ;
	output \outport[2]  ;
	output \outport[3]  ;
	output \outport[4]  ;
	output \outport[5]  ;
	output \outport[6]  ;
	output \outport[7]  ;
	output \outport[8]  ;
	output \outport[9]  ;
	output \outport[10]  ;
	output \outport[11]  ;
	output \outport[12]  ;
	output \outport[13]  ;
	output \outport[14]  ;
	output \outport[15]  ;
	output \outport[16]  ;
	output \outport[17]  ;
	output \outport[18]  ;
	output \outport[19]  ;
	output \outport[20]  ;
	output \outport[21]  ;
	output \outport[22]  ;
	output \outport[23]  ;
	output \outport[24]  ;
	output \outport[25]  ;
	output \outport[26]  ;
	output \outport[27]  ;
	output \outport[28]  ;
	output \outport[29]  ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\dest_x[9] ,
		\dest_x[10] ,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\dest_x[11] ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\dest_x[12] ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\dest_x[13] ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\dest_x[14] ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\dest_x[15] ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\dest_x[16] ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\dest_x[17] ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\dest_x[18] ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\dest_x[19] ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\dest_x[20] ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\dest_x[21] ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\dest_x[22] ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\dest_x[23] ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\dest_x[24] ,
		\dest_x[25] ,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\dest_x[26] ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\dest_x[27] ,
		\dest_x[28] ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\dest_x[29] ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w77_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\dest_x[13] ,
		_w63_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\dest_x[14] ,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\dest_x[20] ,
		\dest_x[21] ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w75_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\dest_x[17] ,
		\dest_x[18] ,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\dest_x[22] ,
		_w72_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\dest_x[23] ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\dest_x[0] ,
		\dest_x[1] ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\dest_x[2] ,
		\dest_x[3] ,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\dest_x[4] ,
		\dest_x[5] ,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\dest_x[6] ,
		\dest_x[7] ,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\dest_x[8] ,
		\dest_x[11] ,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\dest_x[12] ,
		\dest_x[15] ,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\dest_x[19] ,
		\dest_x[26] ,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w93_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w91_,
		_w92_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w89_,
		_w90_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w61_,
		_w88_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w85_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w96_,
		_w97_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w79_,
		_w95_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w84_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w99_,
		_w100_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w65_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w82_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w67_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w74_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w87_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w80_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\dest_x[14] ,
		\dest_x[15] ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w63_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\dest_x[16] ,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\dest_x[26] ,
		_w76_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\dest_x[1] ,
		\dest_x[2] ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		\dest_x[3] ,
		\dest_x[4] ,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\dest_x[5] ,
		\dest_x[6] ,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\dest_x[7] ,
		\dest_x[8] ,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\dest_x[9] ,
		\dest_x[10] ,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\dest_x[11] ,
		\dest_x[12] ,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		\dest_x[13] ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w118_,
		_w119_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w116_,
		_w117_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w85_,
		_w115_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w121_,
		_w122_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w84_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w125_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w113_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w67_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w70_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w86_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w74_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w114_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		_w80_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w110_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\dest_y[9] ,
		\dest_y[10] ,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\dest_y[11] ,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\dest_y[12] ,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\dest_y[13] ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\dest_y[14] ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\dest_y[15] ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\dest_y[16] ,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\dest_y[17] ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\dest_y[18] ,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\dest_y[19] ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\dest_y[20] ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\dest_y[21] ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\dest_y[22] ,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\dest_y[23] ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\dest_y[24] ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\dest_y[25] ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\dest_y[26] ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\dest_y[27] ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\dest_y[28] ,
		\dest_y[29] ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\dest_y[24] ,
		_w150_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w151_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\dest_y[11] ,
		\dest_y[12] ,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\dest_y[15] ,
		\dest_y[16] ,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\dest_y[18] ,
		\dest_y[19] ,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		\dest_y[22] ,
		\dest_y[23] ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w161_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w159_,
		_w160_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\dest_y[13] ,
		_w139_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\dest_y[20] ,
		_w146_,
		_w167_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\dest_y[21] ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\dest_y[25] ,
		_w151_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w152_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\dest_y[26] ,
		_w152_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\dest_y[1] ,
		\dest_y[2] ,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\dest_y[3] ,
		\dest_y[4] ,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\dest_y[5] ,
		\dest_y[6] ,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\dest_y[7] ,
		\dest_y[8] ,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\dest_y[9] ,
		\dest_y[10] ,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\dest_y[17] ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w174_,
		_w175_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w172_,
		_w173_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w177_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w165_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w166_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w141_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w148_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w168_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w158_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w170_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w171_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\dest_x[0] ,
		\dest_y[0] ,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w156_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\dest_y[17] ,
		_w141_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\dest_y[27] ,
		_w171_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\dest_y[17] ,
		_w141_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\dest_y[0] ,
		\dest_y[1] ,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\dest_y[2] ,
		\dest_y[3] ,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		\dest_y[4] ,
		\dest_y[5] ,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\dest_y[6] ,
		\dest_y[7] ,
		_w199_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\dest_y[8] ,
		\dest_y[13] ,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\dest_y[14] ,
		\dest_y[21] ,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w198_,
		_w199_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w196_,
		_w197_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w137_,
		_w155_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w202_,
		_w203_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w165_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w193_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w195_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w147_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w167_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w158_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w170_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w154_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w194_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w192_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\dest_x[0] ,
		_w156_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w110_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w218_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w135_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\dest_x[0] ,
		\dest_y[0] ,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		_w154_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w189_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w136_,
		_w156_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w225_,
		_w226_,
		_w227_
	);
	assign \outport[0]  = _w136_ ;
	assign \outport[1]  = _w222_ ;
	assign \outport[2]  = _w227_ ;
	assign \outport[3]  = 1'b0;
	assign \outport[4]  = 1'b0;
	assign \outport[5]  = 1'b0;
	assign \outport[6]  = 1'b0;
	assign \outport[7]  = 1'b0;
	assign \outport[8]  = 1'b0;
	assign \outport[9]  = 1'b0;
	assign \outport[10]  = 1'b0;
	assign \outport[11]  = 1'b0;
	assign \outport[12]  = 1'b0;
	assign \outport[13]  = 1'b0;
	assign \outport[14]  = 1'b0;
	assign \outport[15]  = 1'b0;
	assign \outport[16]  = 1'b0;
	assign \outport[17]  = 1'b0;
	assign \outport[18]  = 1'b0;
	assign \outport[19]  = 1'b0;
	assign \outport[20]  = 1'b0;
	assign \outport[21]  = 1'b0;
	assign \outport[22]  = 1'b0;
	assign \outport[23]  = 1'b0;
	assign \outport[24]  = 1'b0;
	assign \outport[25]  = 1'b0;
	assign \outport[26]  = 1'b0;
	assign \outport[27]  = 1'b0;
	assign \outport[28]  = 1'b0;
	assign \outport[29]  = 1'b0;
endmodule;