module top (\P1_BE_n_reg[0]/NET0131 , \P1_BE_n_reg[1]/NET0131 , \P1_BE_n_reg[2]/NET0131 , \P1_BE_n_reg[3]/NET0131 , \P1_ByteEnable_reg[0]/NET0131 , \P1_ByteEnable_reg[1]/NET0131 , \P1_ByteEnable_reg[2]/NET0131 , \P1_ByteEnable_reg[3]/NET0131 , \P1_CodeFetch_reg/NET0131 , \P1_D_C_n_reg/NET0131 , \P1_DataWidth_reg[0]/NET0131 , \P1_DataWidth_reg[1]/NET0131 , \P1_Datao_reg[0]/NET0131 , \P1_Datao_reg[10]/NET0131 , \P1_Datao_reg[11]/NET0131 , \P1_Datao_reg[12]/NET0131 , \P1_Datao_reg[13]/NET0131 , \P1_Datao_reg[14]/NET0131 , \P1_Datao_reg[15]/NET0131 , \P1_Datao_reg[16]/NET0131 , \P1_Datao_reg[17]/NET0131 , \P1_Datao_reg[18]/NET0131 , \P1_Datao_reg[19]/NET0131 , \P1_Datao_reg[1]/NET0131 , \P1_Datao_reg[20]/NET0131 , \P1_Datao_reg[21]/NET0131 , \P1_Datao_reg[22]/NET0131 , \P1_Datao_reg[23]/NET0131 , \P1_Datao_reg[24]/NET0131 , \P1_Datao_reg[25]/NET0131 , \P1_Datao_reg[26]/NET0131 , \P1_Datao_reg[27]/NET0131 , \P1_Datao_reg[28]/NET0131 , \P1_Datao_reg[29]/NET0131 , \P1_Datao_reg[2]/NET0131 , \P1_Datao_reg[30]/NET0131 , \P1_Datao_reg[3]/NET0131 , \P1_Datao_reg[4]/NET0131 , \P1_Datao_reg[5]/NET0131 , \P1_Datao_reg[6]/NET0131 , \P1_Datao_reg[7]/NET0131 , \P1_Datao_reg[8]/NET0131 , \P1_Datao_reg[9]/NET0131 , \P1_EAX_reg[0]/NET0131 , \P1_EAX_reg[10]/NET0131 , \P1_EAX_reg[11]/NET0131 , \P1_EAX_reg[12]/NET0131 , \P1_EAX_reg[13]/NET0131 , \P1_EAX_reg[14]/NET0131 , \P1_EAX_reg[15]/NET0131 , \P1_EAX_reg[16]/NET0131 , \P1_EAX_reg[17]/NET0131 , \P1_EAX_reg[18]/NET0131 , \P1_EAX_reg[19]/NET0131 , \P1_EAX_reg[1]/NET0131 , \P1_EAX_reg[20]/NET0131 , \P1_EAX_reg[21]/NET0131 , \P1_EAX_reg[22]/NET0131 , \P1_EAX_reg[23]/NET0131 , \P1_EAX_reg[24]/NET0131 , \P1_EAX_reg[25]/NET0131 , \P1_EAX_reg[26]/NET0131 , \P1_EAX_reg[27]/NET0131 , \P1_EAX_reg[28]/NET0131 , \P1_EAX_reg[29]/NET0131 , \P1_EAX_reg[2]/NET0131 , \P1_EAX_reg[30]/NET0131 , \P1_EAX_reg[31]/NET0131 , \P1_EAX_reg[3]/NET0131 , \P1_EAX_reg[4]/NET0131 , \P1_EAX_reg[5]/NET0131 , \P1_EAX_reg[6]/NET0131 , \P1_EAX_reg[7]/NET0131 , \P1_EAX_reg[8]/NET0131 , \P1_EAX_reg[9]/NET0131 , \P1_EBX_reg[0]/NET0131 , \P1_EBX_reg[10]/NET0131 , \P1_EBX_reg[11]/NET0131 , \P1_EBX_reg[12]/NET0131 , \P1_EBX_reg[13]/NET0131 , \P1_EBX_reg[14]/NET0131 , \P1_EBX_reg[15]/NET0131 , \P1_EBX_reg[16]/NET0131 , \P1_EBX_reg[17]/NET0131 , \P1_EBX_reg[18]/NET0131 , \P1_EBX_reg[19]/NET0131 , \P1_EBX_reg[1]/NET0131 , \P1_EBX_reg[20]/NET0131 , \P1_EBX_reg[21]/NET0131 , \P1_EBX_reg[22]/NET0131 , \P1_EBX_reg[23]/NET0131 , \P1_EBX_reg[24]/NET0131 , \P1_EBX_reg[25]/NET0131 , \P1_EBX_reg[26]/NET0131 , \P1_EBX_reg[27]/NET0131 , \P1_EBX_reg[28]/NET0131 , \P1_EBX_reg[29]/NET0131 , \P1_EBX_reg[2]/NET0131 , \P1_EBX_reg[30]/NET0131 , \P1_EBX_reg[31]/NET0131 , \P1_EBX_reg[3]/NET0131 , \P1_EBX_reg[4]/NET0131 , \P1_EBX_reg[5]/NET0131 , \P1_EBX_reg[6]/NET0131 , \P1_EBX_reg[7]/NET0131 , \P1_EBX_reg[8]/NET0131 , \P1_EBX_reg[9]/NET0131 , \P1_Flush_reg/NET0131 , \P1_InstAddrPointer_reg[0]/NET0131 , \P1_InstAddrPointer_reg[10]/NET0131 , \P1_InstAddrPointer_reg[11]/NET0131 , \P1_InstAddrPointer_reg[12]/NET0131 , \P1_InstAddrPointer_reg[13]/NET0131 , \P1_InstAddrPointer_reg[14]/NET0131 , \P1_InstAddrPointer_reg[15]/NET0131 , \P1_InstAddrPointer_reg[16]/NET0131 , \P1_InstAddrPointer_reg[17]/NET0131 , \P1_InstAddrPointer_reg[18]/NET0131 , \P1_InstAddrPointer_reg[19]/NET0131 , \P1_InstAddrPointer_reg[1]/NET0131 , \P1_InstAddrPointer_reg[20]/NET0131 , \P1_InstAddrPointer_reg[21]/NET0131 , \P1_InstAddrPointer_reg[22]/NET0131 , \P1_InstAddrPointer_reg[23]/NET0131 , \P1_InstAddrPointer_reg[24]/NET0131 , \P1_InstAddrPointer_reg[25]/NET0131 , \P1_InstAddrPointer_reg[26]/NET0131 , \P1_InstAddrPointer_reg[27]/NET0131 , \P1_InstAddrPointer_reg[28]/NET0131 , \P1_InstAddrPointer_reg[29]/NET0131 , \P1_InstAddrPointer_reg[2]/NET0131 , \P1_InstAddrPointer_reg[30]/NET0131 , \P1_InstAddrPointer_reg[31]/NET0131 , \P1_InstAddrPointer_reg[3]/NET0131 , \P1_InstAddrPointer_reg[4]/NET0131 , \P1_InstAddrPointer_reg[5]/NET0131 , \P1_InstAddrPointer_reg[6]/NET0131 , \P1_InstAddrPointer_reg[7]/NET0131 , \P1_InstAddrPointer_reg[8]/NET0131 , \P1_InstAddrPointer_reg[9]/NET0131 , \P1_InstQueueRd_Addr_reg[0]/NET0131 , \P1_InstQueueRd_Addr_reg[1]/NET0131 , \P1_InstQueueRd_Addr_reg[2]/NET0131 , \P1_InstQueueRd_Addr_reg[3]/NET0131 , \P1_InstQueueWr_Addr_reg[0]/NET0131 , \P1_InstQueueWr_Addr_reg[1]/NET0131 , \P1_InstQueueWr_Addr_reg[2]/NET0131 , \P1_InstQueueWr_Addr_reg[3]/NET0131 , \P1_InstQueue_reg[0][0]/NET0131 , \P1_InstQueue_reg[0][1]/NET0131 , \P1_InstQueue_reg[0][2]/NET0131 , \P1_InstQueue_reg[0][3]/NET0131 , \P1_InstQueue_reg[0][4]/NET0131 , \P1_InstQueue_reg[0][5]/NET0131 , \P1_InstQueue_reg[0][6]/NET0131 , \P1_InstQueue_reg[0][7]/NET0131 , \P1_InstQueue_reg[10][0]/NET0131 , \P1_InstQueue_reg[10][1]/NET0131 , \P1_InstQueue_reg[10][2]/NET0131 , \P1_InstQueue_reg[10][3]/NET0131 , \P1_InstQueue_reg[10][4]/NET0131 , \P1_InstQueue_reg[10][5]/NET0131 , \P1_InstQueue_reg[10][6]/NET0131 , \P1_InstQueue_reg[10][7]/NET0131 , \P1_InstQueue_reg[11][0]/NET0131 , \P1_InstQueue_reg[11][1]/NET0131 , \P1_InstQueue_reg[11][2]/NET0131 , \P1_InstQueue_reg[11][3]/NET0131 , \P1_InstQueue_reg[11][4]/NET0131 , \P1_InstQueue_reg[11][5]/NET0131 , \P1_InstQueue_reg[11][6]/NET0131 , \P1_InstQueue_reg[11][7]/NET0131 , \P1_InstQueue_reg[12][0]/NET0131 , \P1_InstQueue_reg[12][1]/NET0131 , \P1_InstQueue_reg[12][2]/NET0131 , \P1_InstQueue_reg[12][3]/NET0131 , \P1_InstQueue_reg[12][4]/NET0131 , \P1_InstQueue_reg[12][5]/NET0131 , \P1_InstQueue_reg[12][6]/NET0131 , \P1_InstQueue_reg[12][7]/NET0131 , \P1_InstQueue_reg[13][0]/NET0131 , \P1_InstQueue_reg[13][1]/NET0131 , \P1_InstQueue_reg[13][2]/NET0131 , \P1_InstQueue_reg[13][3]/NET0131 , \P1_InstQueue_reg[13][4]/NET0131 , \P1_InstQueue_reg[13][5]/NET0131 , \P1_InstQueue_reg[13][6]/NET0131 , \P1_InstQueue_reg[13][7]/NET0131 , \P1_InstQueue_reg[14][0]/NET0131 , \P1_InstQueue_reg[14][1]/NET0131 , \P1_InstQueue_reg[14][2]/NET0131 , \P1_InstQueue_reg[14][3]/NET0131 , \P1_InstQueue_reg[14][4]/NET0131 , \P1_InstQueue_reg[14][5]/NET0131 , \P1_InstQueue_reg[14][6]/NET0131 , \P1_InstQueue_reg[14][7]/NET0131 , \P1_InstQueue_reg[15][0]/NET0131 , \P1_InstQueue_reg[15][1]/NET0131 , \P1_InstQueue_reg[15][2]/NET0131 , \P1_InstQueue_reg[15][3]/NET0131 , \P1_InstQueue_reg[15][4]/NET0131 , \P1_InstQueue_reg[15][5]/NET0131 , \P1_InstQueue_reg[15][6]/NET0131 , \P1_InstQueue_reg[15][7]/NET0131 , \P1_InstQueue_reg[1][0]/NET0131 , \P1_InstQueue_reg[1][1]/NET0131 , \P1_InstQueue_reg[1][2]/NET0131 , \P1_InstQueue_reg[1][3]/NET0131 , \P1_InstQueue_reg[1][4]/NET0131 , \P1_InstQueue_reg[1][5]/NET0131 , \P1_InstQueue_reg[1][6]/NET0131 , \P1_InstQueue_reg[1][7]/NET0131 , \P1_InstQueue_reg[2][0]/NET0131 , \P1_InstQueue_reg[2][1]/NET0131 , \P1_InstQueue_reg[2][2]/NET0131 , \P1_InstQueue_reg[2][3]/NET0131 , \P1_InstQueue_reg[2][4]/NET0131 , \P1_InstQueue_reg[2][5]/NET0131 , \P1_InstQueue_reg[2][6]/NET0131 , \P1_InstQueue_reg[2][7]/NET0131 , \P1_InstQueue_reg[3][0]/NET0131 , \P1_InstQueue_reg[3][1]/NET0131 , \P1_InstQueue_reg[3][2]/NET0131 , \P1_InstQueue_reg[3][3]/NET0131 , \P1_InstQueue_reg[3][4]/NET0131 , \P1_InstQueue_reg[3][5]/NET0131 , \P1_InstQueue_reg[3][6]/NET0131 , \P1_InstQueue_reg[3][7]/NET0131 , \P1_InstQueue_reg[4][0]/NET0131 , \P1_InstQueue_reg[4][1]/NET0131 , \P1_InstQueue_reg[4][2]/NET0131 , \P1_InstQueue_reg[4][3]/NET0131 , \P1_InstQueue_reg[4][4]/NET0131 , \P1_InstQueue_reg[4][5]/NET0131 , \P1_InstQueue_reg[4][6]/NET0131 , \P1_InstQueue_reg[4][7]/NET0131 , \P1_InstQueue_reg[5][0]/NET0131 , \P1_InstQueue_reg[5][1]/NET0131 , \P1_InstQueue_reg[5][2]/NET0131 , \P1_InstQueue_reg[5][3]/NET0131 , \P1_InstQueue_reg[5][4]/NET0131 , \P1_InstQueue_reg[5][5]/NET0131 , \P1_InstQueue_reg[5][6]/NET0131 , \P1_InstQueue_reg[5][7]/NET0131 , \P1_InstQueue_reg[6][0]/NET0131 , \P1_InstQueue_reg[6][1]/NET0131 , \P1_InstQueue_reg[6][2]/NET0131 , \P1_InstQueue_reg[6][3]/NET0131 , \P1_InstQueue_reg[6][4]/NET0131 , \P1_InstQueue_reg[6][5]/NET0131 , \P1_InstQueue_reg[6][6]/NET0131 , \P1_InstQueue_reg[6][7]/NET0131 , \P1_InstQueue_reg[7][0]/NET0131 , \P1_InstQueue_reg[7][1]/NET0131 , \P1_InstQueue_reg[7][2]/NET0131 , \P1_InstQueue_reg[7][3]/NET0131 , \P1_InstQueue_reg[7][4]/NET0131 , \P1_InstQueue_reg[7][5]/NET0131 , \P1_InstQueue_reg[7][6]/NET0131 , \P1_InstQueue_reg[7][7]/NET0131 , \P1_InstQueue_reg[8][0]/NET0131 , \P1_InstQueue_reg[8][1]/NET0131 , \P1_InstQueue_reg[8][2]/NET0131 , \P1_InstQueue_reg[8][3]/NET0131 , \P1_InstQueue_reg[8][4]/NET0131 , \P1_InstQueue_reg[8][5]/NET0131 , \P1_InstQueue_reg[8][6]/NET0131 , \P1_InstQueue_reg[8][7]/NET0131 , \P1_InstQueue_reg[9][0]/NET0131 , \P1_InstQueue_reg[9][1]/NET0131 , \P1_InstQueue_reg[9][2]/NET0131 , \P1_InstQueue_reg[9][3]/NET0131 , \P1_InstQueue_reg[9][4]/NET0131 , \P1_InstQueue_reg[9][5]/NET0131 , \P1_InstQueue_reg[9][6]/NET0131 , \P1_InstQueue_reg[9][7]/NET0131 , \P1_M_IO_n_reg/NET0131 , \P1_MemoryFetch_reg/NET0131 , \P1_More_reg/NET0131 , \P1_PhyAddrPointer_reg[0]/NET0131 , \P1_PhyAddrPointer_reg[10]/NET0131 , \P1_PhyAddrPointer_reg[11]/NET0131 , \P1_PhyAddrPointer_reg[12]/NET0131 , \P1_PhyAddrPointer_reg[13]/NET0131 , \P1_PhyAddrPointer_reg[14]/NET0131 , \P1_PhyAddrPointer_reg[15]/NET0131 , \P1_PhyAddrPointer_reg[16]/NET0131 , \P1_PhyAddrPointer_reg[17]/NET0131 , \P1_PhyAddrPointer_reg[18]/NET0131 , \P1_PhyAddrPointer_reg[19]/NET0131 , \P1_PhyAddrPointer_reg[1]/NET0131 , \P1_PhyAddrPointer_reg[20]/NET0131 , \P1_PhyAddrPointer_reg[21]/NET0131 , \P1_PhyAddrPointer_reg[22]/NET0131 , \P1_PhyAddrPointer_reg[23]/NET0131 , \P1_PhyAddrPointer_reg[24]/NET0131 , \P1_PhyAddrPointer_reg[25]/NET0131 , \P1_PhyAddrPointer_reg[26]/NET0131 , \P1_PhyAddrPointer_reg[27]/NET0131 , \P1_PhyAddrPointer_reg[28]/NET0131 , \P1_PhyAddrPointer_reg[29]/NET0131 , \P1_PhyAddrPointer_reg[2]/NET0131 , \P1_PhyAddrPointer_reg[30]/NET0131 , \P1_PhyAddrPointer_reg[31]/NET0131 , \P1_PhyAddrPointer_reg[3]/NET0131 , \P1_PhyAddrPointer_reg[4]/NET0131 , \P1_PhyAddrPointer_reg[5]/NET0131 , \P1_PhyAddrPointer_reg[6]/NET0131 , \P1_PhyAddrPointer_reg[7]/NET0131 , \P1_PhyAddrPointer_reg[8]/NET0131 , \P1_PhyAddrPointer_reg[9]/NET0131 , \P1_ReadRequest_reg/NET0131 , \P1_RequestPending_reg/NET0131 , \P1_State2_reg[0]/NET0131 , \P1_State2_reg[1]/NET0131 , \P1_State2_reg[2]/NET0131 , \P1_State2_reg[3]/NET0131 , \P1_State_reg[0]/NET0131 , \P1_State_reg[1]/NET0131 , \P1_State_reg[2]/NET0131 , \P1_W_R_n_reg/NET0131 , \P1_lWord_reg[0]/NET0131 , \P1_lWord_reg[10]/NET0131 , \P1_lWord_reg[11]/NET0131 , \P1_lWord_reg[12]/NET0131 , \P1_lWord_reg[13]/NET0131 , \P1_lWord_reg[14]/NET0131 , \P1_lWord_reg[15]/NET0131 , \P1_lWord_reg[1]/NET0131 , \P1_lWord_reg[2]/NET0131 , \P1_lWord_reg[3]/NET0131 , \P1_lWord_reg[4]/NET0131 , \P1_lWord_reg[5]/NET0131 , \P1_lWord_reg[6]/NET0131 , \P1_lWord_reg[7]/NET0131 , \P1_lWord_reg[8]/NET0131 , \P1_lWord_reg[9]/NET0131 , \P1_rEIP_reg[0]/NET0131 , \P1_rEIP_reg[10]/NET0131 , \P1_rEIP_reg[11]/NET0131 , \P1_rEIP_reg[12]/NET0131 , \P1_rEIP_reg[13]/NET0131 , \P1_rEIP_reg[14]/NET0131 , \P1_rEIP_reg[15]/NET0131 , \P1_rEIP_reg[16]/NET0131 , \P1_rEIP_reg[17]/NET0131 , \P1_rEIP_reg[18]/NET0131 , \P1_rEIP_reg[19]/NET0131 , \P1_rEIP_reg[1]/NET0131 , \P1_rEIP_reg[20]/NET0131 , \P1_rEIP_reg[21]/NET0131 , \P1_rEIP_reg[22]/NET0131 , \P1_rEIP_reg[23]/NET0131 , \P1_rEIP_reg[24]/NET0131 , \P1_rEIP_reg[25]/NET0131 , \P1_rEIP_reg[26]/NET0131 , \P1_rEIP_reg[27]/NET0131 , \P1_rEIP_reg[28]/NET0131 , \P1_rEIP_reg[29]/NET0131 , \P1_rEIP_reg[2]/NET0131 , \P1_rEIP_reg[30]/NET0131 , \P1_rEIP_reg[31]/NET0131 , \P1_rEIP_reg[3]/NET0131 , \P1_rEIP_reg[4]/NET0131 , \P1_rEIP_reg[5]/NET0131 , \P1_rEIP_reg[6]/NET0131 , \P1_rEIP_reg[7]/NET0131 , \P1_rEIP_reg[8]/NET0131 , \P1_rEIP_reg[9]/NET0131 , \P1_uWord_reg[0]/NET0131 , \P1_uWord_reg[10]/NET0131 , \P1_uWord_reg[11]/NET0131 , \P1_uWord_reg[12]/NET0131 , \P1_uWord_reg[13]/NET0131 , \P1_uWord_reg[14]/NET0131 , \P1_uWord_reg[1]/NET0131 , \P1_uWord_reg[2]/NET0131 , \P1_uWord_reg[3]/NET0131 , \P1_uWord_reg[4]/NET0131 , \P1_uWord_reg[5]/NET0131 , \P1_uWord_reg[6]/NET0131 , \P1_uWord_reg[7]/NET0131 , \P1_uWord_reg[8]/NET0131 , \P1_uWord_reg[9]/NET0131 , \P2_ADS_n_reg/NET0131 , \P2_Address_reg[0]/NET0131 , \P2_Address_reg[10]/NET0131 , \P2_Address_reg[11]/NET0131 , \P2_Address_reg[12]/NET0131 , \P2_Address_reg[13]/NET0131 , \P2_Address_reg[14]/NET0131 , \P2_Address_reg[15]/NET0131 , \P2_Address_reg[16]/NET0131 , \P2_Address_reg[17]/NET0131 , \P2_Address_reg[18]/NET0131 , \P2_Address_reg[19]/NET0131 , \P2_Address_reg[1]/NET0131 , \P2_Address_reg[20]/NET0131 , \P2_Address_reg[21]/NET0131 , \P2_Address_reg[22]/NET0131 , \P2_Address_reg[23]/NET0131 , \P2_Address_reg[24]/NET0131 , \P2_Address_reg[25]/NET0131 , \P2_Address_reg[26]/NET0131 , \P2_Address_reg[27]/NET0131 , \P2_Address_reg[28]/NET0131 , \P2_Address_reg[29]/NET0131 , \P2_Address_reg[2]/NET0131 , \P2_Address_reg[3]/NET0131 , \P2_Address_reg[4]/NET0131 , \P2_Address_reg[5]/NET0131 , \P2_Address_reg[6]/NET0131 , \P2_Address_reg[7]/NET0131 , \P2_Address_reg[8]/NET0131 , \P2_Address_reg[9]/NET0131 , \P2_BE_n_reg[0]/NET0131 , \P2_BE_n_reg[1]/NET0131 , \P2_BE_n_reg[2]/NET0131 , \P2_BE_n_reg[3]/NET0131 , \P2_ByteEnable_reg[0]/NET0131 , \P2_ByteEnable_reg[1]/NET0131 , \P2_ByteEnable_reg[2]/NET0131 , \P2_ByteEnable_reg[3]/NET0131 , \P2_CodeFetch_reg/NET0131 , \P2_D_C_n_reg/NET0131 , \P2_DataWidth_reg[0]/NET0131 , \P2_DataWidth_reg[1]/NET0131 , \P2_Datao_reg[0]/NET0131 , \P2_Datao_reg[10]/NET0131 , \P2_Datao_reg[11]/NET0131 , \P2_Datao_reg[12]/NET0131 , \P2_Datao_reg[13]/NET0131 , \P2_Datao_reg[14]/NET0131 , \P2_Datao_reg[15]/NET0131 , \P2_Datao_reg[16]/NET0131 , \P2_Datao_reg[17]/NET0131 , \P2_Datao_reg[18]/NET0131 , \P2_Datao_reg[19]/NET0131 , \P2_Datao_reg[1]/NET0131 , \P2_Datao_reg[20]/NET0131 , \P2_Datao_reg[21]/NET0131 , \P2_Datao_reg[22]/NET0131 , \P2_Datao_reg[23]/NET0131 , \P2_Datao_reg[24]/NET0131 , \P2_Datao_reg[25]/NET0131 , \P2_Datao_reg[26]/NET0131 , \P2_Datao_reg[27]/NET0131 , \P2_Datao_reg[28]/NET0131 , \P2_Datao_reg[29]/NET0131 , \P2_Datao_reg[2]/NET0131 , \P2_Datao_reg[30]/NET0131 , \P2_Datao_reg[3]/NET0131 , \P2_Datao_reg[4]/NET0131 , \P2_Datao_reg[5]/NET0131 , \P2_Datao_reg[6]/NET0131 , \P2_Datao_reg[7]/NET0131 , \P2_Datao_reg[8]/NET0131 , \P2_Datao_reg[9]/NET0131 , \P2_EAX_reg[0]/NET0131 , \P2_EAX_reg[10]/NET0131 , \P2_EAX_reg[11]/NET0131 , \P2_EAX_reg[12]/NET0131 , \P2_EAX_reg[13]/NET0131 , \P2_EAX_reg[14]/NET0131 , \P2_EAX_reg[15]/NET0131 , \P2_EAX_reg[16]/NET0131 , \P2_EAX_reg[17]/NET0131 , \P2_EAX_reg[18]/NET0131 , \P2_EAX_reg[19]/NET0131 , \P2_EAX_reg[1]/NET0131 , \P2_EAX_reg[20]/NET0131 , \P2_EAX_reg[21]/NET0131 , \P2_EAX_reg[22]/NET0131 , \P2_EAX_reg[23]/NET0131 , \P2_EAX_reg[24]/NET0131 , \P2_EAX_reg[25]/NET0131 , \P2_EAX_reg[26]/NET0131 , \P2_EAX_reg[27]/NET0131 , \P2_EAX_reg[28]/NET0131 , \P2_EAX_reg[29]/NET0131 , \P2_EAX_reg[2]/NET0131 , \P2_EAX_reg[30]/NET0131 , \P2_EAX_reg[31]/NET0131 , \P2_EAX_reg[3]/NET0131 , \P2_EAX_reg[4]/NET0131 , \P2_EAX_reg[5]/NET0131 , \P2_EAX_reg[6]/NET0131 , \P2_EAX_reg[7]/NET0131 , \P2_EAX_reg[8]/NET0131 , \P2_EAX_reg[9]/NET0131 , \P2_EBX_reg[0]/NET0131 , \P2_EBX_reg[10]/NET0131 , \P2_EBX_reg[11]/NET0131 , \P2_EBX_reg[12]/NET0131 , \P2_EBX_reg[13]/NET0131 , \P2_EBX_reg[14]/NET0131 , \P2_EBX_reg[15]/NET0131 , \P2_EBX_reg[16]/NET0131 , \P2_EBX_reg[17]/NET0131 , \P2_EBX_reg[18]/NET0131 , \P2_EBX_reg[19]/NET0131 , \P2_EBX_reg[1]/NET0131 , \P2_EBX_reg[20]/NET0131 , \P2_EBX_reg[21]/NET0131 , \P2_EBX_reg[22]/NET0131 , \P2_EBX_reg[23]/NET0131 , \P2_EBX_reg[24]/NET0131 , \P2_EBX_reg[25]/NET0131 , \P2_EBX_reg[26]/NET0131 , \P2_EBX_reg[27]/NET0131 , \P2_EBX_reg[28]/NET0131 , \P2_EBX_reg[29]/NET0131 , \P2_EBX_reg[2]/NET0131 , \P2_EBX_reg[30]/NET0131 , \P2_EBX_reg[31]/NET0131 , \P2_EBX_reg[3]/NET0131 , \P2_EBX_reg[4]/NET0131 , \P2_EBX_reg[5]/NET0131 , \P2_EBX_reg[6]/NET0131 , \P2_EBX_reg[7]/NET0131 , \P2_EBX_reg[8]/NET0131 , \P2_EBX_reg[9]/NET0131 , \P2_Flush_reg/NET0131 , \P2_InstAddrPointer_reg[0]/NET0131 , \P2_InstAddrPointer_reg[10]/NET0131 , \P2_InstAddrPointer_reg[11]/NET0131 , \P2_InstAddrPointer_reg[12]/NET0131 , \P2_InstAddrPointer_reg[13]/NET0131 , \P2_InstAddrPointer_reg[14]/NET0131 , \P2_InstAddrPointer_reg[15]/NET0131 , \P2_InstAddrPointer_reg[16]/NET0131 , \P2_InstAddrPointer_reg[17]/NET0131 , \P2_InstAddrPointer_reg[18]/NET0131 , \P2_InstAddrPointer_reg[19]/NET0131 , \P2_InstAddrPointer_reg[1]/NET0131 , \P2_InstAddrPointer_reg[20]/NET0131 , \P2_InstAddrPointer_reg[21]/NET0131 , \P2_InstAddrPointer_reg[22]/NET0131 , \P2_InstAddrPointer_reg[23]/NET0131 , \P2_InstAddrPointer_reg[24]/NET0131 , \P2_InstAddrPointer_reg[25]/NET0131 , \P2_InstAddrPointer_reg[26]/NET0131 , \P2_InstAddrPointer_reg[27]/NET0131 , \P2_InstAddrPointer_reg[28]/NET0131 , \P2_InstAddrPointer_reg[29]/NET0131 , \P2_InstAddrPointer_reg[2]/NET0131 , \P2_InstAddrPointer_reg[30]/NET0131 , \P2_InstAddrPointer_reg[31]/NET0131 , \P2_InstAddrPointer_reg[3]/NET0131 , \P2_InstAddrPointer_reg[4]/NET0131 , \P2_InstAddrPointer_reg[5]/NET0131 , \P2_InstAddrPointer_reg[6]/NET0131 , \P2_InstAddrPointer_reg[7]/NET0131 , \P2_InstAddrPointer_reg[8]/NET0131 , \P2_InstAddrPointer_reg[9]/NET0131 , \P2_InstQueueRd_Addr_reg[0]/NET0131 , \P2_InstQueueRd_Addr_reg[1]/NET0131 , \P2_InstQueueRd_Addr_reg[2]/NET0131 , \P2_InstQueueRd_Addr_reg[3]/NET0131 , \P2_InstQueueWr_Addr_reg[0]/NET0131 , \P2_InstQueueWr_Addr_reg[1]/NET0131 , \P2_InstQueueWr_Addr_reg[2]/NET0131 , \P2_InstQueueWr_Addr_reg[3]/NET0131 , \P2_InstQueue_reg[0][0]/NET0131 , \P2_InstQueue_reg[0][1]/NET0131 , \P2_InstQueue_reg[0][2]/NET0131 , \P2_InstQueue_reg[0][3]/NET0131 , \P2_InstQueue_reg[0][4]/NET0131 , \P2_InstQueue_reg[0][5]/NET0131 , \P2_InstQueue_reg[0][6]/NET0131 , \P2_InstQueue_reg[0][7]/NET0131 , \P2_InstQueue_reg[10][0]/NET0131 , \P2_InstQueue_reg[10][1]/NET0131 , \P2_InstQueue_reg[10][2]/NET0131 , \P2_InstQueue_reg[10][3]/NET0131 , \P2_InstQueue_reg[10][4]/NET0131 , \P2_InstQueue_reg[10][5]/NET0131 , \P2_InstQueue_reg[10][6]/NET0131 , \P2_InstQueue_reg[10][7]/NET0131 , \P2_InstQueue_reg[11][0]/NET0131 , \P2_InstQueue_reg[11][1]/NET0131 , \P2_InstQueue_reg[11][2]/NET0131 , \P2_InstQueue_reg[11][3]/NET0131 , \P2_InstQueue_reg[11][4]/NET0131 , \P2_InstQueue_reg[11][5]/NET0131 , \P2_InstQueue_reg[11][6]/NET0131 , \P2_InstQueue_reg[11][7]/NET0131 , \P2_InstQueue_reg[12][0]/NET0131 , \P2_InstQueue_reg[12][1]/NET0131 , \P2_InstQueue_reg[12][2]/NET0131 , \P2_InstQueue_reg[12][3]/NET0131 , \P2_InstQueue_reg[12][4]/NET0131 , \P2_InstQueue_reg[12][5]/NET0131 , \P2_InstQueue_reg[12][6]/NET0131 , \P2_InstQueue_reg[12][7]/NET0131 , \P2_InstQueue_reg[13][0]/NET0131 , \P2_InstQueue_reg[13][1]/NET0131 , \P2_InstQueue_reg[13][2]/NET0131 , \P2_InstQueue_reg[13][3]/NET0131 , \P2_InstQueue_reg[13][4]/NET0131 , \P2_InstQueue_reg[13][5]/NET0131 , \P2_InstQueue_reg[13][6]/NET0131 , \P2_InstQueue_reg[13][7]/NET0131 , \P2_InstQueue_reg[14][0]/NET0131 , \P2_InstQueue_reg[14][1]/NET0131 , \P2_InstQueue_reg[14][2]/NET0131 , \P2_InstQueue_reg[14][3]/NET0131 , \P2_InstQueue_reg[14][4]/NET0131 , \P2_InstQueue_reg[14][5]/NET0131 , \P2_InstQueue_reg[14][6]/NET0131 , \P2_InstQueue_reg[14][7]/NET0131 , \P2_InstQueue_reg[15][0]/NET0131 , \P2_InstQueue_reg[15][1]/NET0131 , \P2_InstQueue_reg[15][2]/NET0131 , \P2_InstQueue_reg[15][3]/NET0131 , \P2_InstQueue_reg[15][4]/NET0131 , \P2_InstQueue_reg[15][5]/NET0131 , \P2_InstQueue_reg[15][6]/NET0131 , \P2_InstQueue_reg[15][7]/NET0131 , \P2_InstQueue_reg[1][0]/NET0131 , \P2_InstQueue_reg[1][1]/NET0131 , \P2_InstQueue_reg[1][2]/NET0131 , \P2_InstQueue_reg[1][3]/NET0131 , \P2_InstQueue_reg[1][4]/NET0131 , \P2_InstQueue_reg[1][5]/NET0131 , \P2_InstQueue_reg[1][6]/NET0131 , \P2_InstQueue_reg[1][7]/NET0131 , \P2_InstQueue_reg[2][0]/NET0131 , \P2_InstQueue_reg[2][1]/NET0131 , \P2_InstQueue_reg[2][2]/NET0131 , \P2_InstQueue_reg[2][3]/NET0131 , \P2_InstQueue_reg[2][4]/NET0131 , \P2_InstQueue_reg[2][5]/NET0131 , \P2_InstQueue_reg[2][6]/NET0131 , \P2_InstQueue_reg[2][7]/NET0131 , \P2_InstQueue_reg[3][0]/NET0131 , \P2_InstQueue_reg[3][1]/NET0131 , \P2_InstQueue_reg[3][2]/NET0131 , \P2_InstQueue_reg[3][3]/NET0131 , \P2_InstQueue_reg[3][4]/NET0131 , \P2_InstQueue_reg[3][5]/NET0131 , \P2_InstQueue_reg[3][6]/NET0131 , \P2_InstQueue_reg[3][7]/NET0131 , \P2_InstQueue_reg[4][0]/NET0131 , \P2_InstQueue_reg[4][1]/NET0131 , \P2_InstQueue_reg[4][2]/NET0131 , \P2_InstQueue_reg[4][3]/NET0131 , \P2_InstQueue_reg[4][4]/NET0131 , \P2_InstQueue_reg[4][5]/NET0131 , \P2_InstQueue_reg[4][6]/NET0131 , \P2_InstQueue_reg[4][7]/NET0131 , \P2_InstQueue_reg[5][0]/NET0131 , \P2_InstQueue_reg[5][1]/NET0131 , \P2_InstQueue_reg[5][2]/NET0131 , \P2_InstQueue_reg[5][3]/NET0131 , \P2_InstQueue_reg[5][4]/NET0131 , \P2_InstQueue_reg[5][5]/NET0131 , \P2_InstQueue_reg[5][6]/NET0131 , \P2_InstQueue_reg[5][7]/NET0131 , \P2_InstQueue_reg[6][0]/NET0131 , \P2_InstQueue_reg[6][1]/NET0131 , \P2_InstQueue_reg[6][2]/NET0131 , \P2_InstQueue_reg[6][3]/NET0131 , \P2_InstQueue_reg[6][4]/NET0131 , \P2_InstQueue_reg[6][5]/NET0131 , \P2_InstQueue_reg[6][6]/NET0131 , \P2_InstQueue_reg[6][7]/NET0131 , \P2_InstQueue_reg[7][0]/NET0131 , \P2_InstQueue_reg[7][1]/NET0131 , \P2_InstQueue_reg[7][2]/NET0131 , \P2_InstQueue_reg[7][3]/NET0131 , \P2_InstQueue_reg[7][4]/NET0131 , \P2_InstQueue_reg[7][5]/NET0131 , \P2_InstQueue_reg[7][6]/NET0131 , \P2_InstQueue_reg[7][7]/NET0131 , \P2_InstQueue_reg[8][0]/NET0131 , \P2_InstQueue_reg[8][1]/NET0131 , \P2_InstQueue_reg[8][2]/NET0131 , \P2_InstQueue_reg[8][3]/NET0131 , \P2_InstQueue_reg[8][4]/NET0131 , \P2_InstQueue_reg[8][5]/NET0131 , \P2_InstQueue_reg[8][6]/NET0131 , \P2_InstQueue_reg[8][7]/NET0131 , \P2_InstQueue_reg[9][0]/NET0131 , \P2_InstQueue_reg[9][1]/NET0131 , \P2_InstQueue_reg[9][2]/NET0131 , \P2_InstQueue_reg[9][3]/NET0131 , \P2_InstQueue_reg[9][4]/NET0131 , \P2_InstQueue_reg[9][5]/NET0131 , \P2_InstQueue_reg[9][6]/NET0131 , \P2_InstQueue_reg[9][7]/NET0131 , \P2_M_IO_n_reg/NET0131 , \P2_MemoryFetch_reg/NET0131 , \P2_More_reg/NET0131 , \P2_PhyAddrPointer_reg[0]/NET0131 , \P2_PhyAddrPointer_reg[10]/NET0131 , \P2_PhyAddrPointer_reg[11]/NET0131 , \P2_PhyAddrPointer_reg[12]/NET0131 , \P2_PhyAddrPointer_reg[13]/NET0131 , \P2_PhyAddrPointer_reg[14]/NET0131 , \P2_PhyAddrPointer_reg[15]/NET0131 , \P2_PhyAddrPointer_reg[16]/NET0131 , \P2_PhyAddrPointer_reg[17]/NET0131 , \P2_PhyAddrPointer_reg[18]/NET0131 , \P2_PhyAddrPointer_reg[19]/NET0131 , \P2_PhyAddrPointer_reg[1]/NET0131 , \P2_PhyAddrPointer_reg[20]/NET0131 , \P2_PhyAddrPointer_reg[21]/NET0131 , \P2_PhyAddrPointer_reg[22]/NET0131 , \P2_PhyAddrPointer_reg[23]/NET0131 , \P2_PhyAddrPointer_reg[24]/NET0131 , \P2_PhyAddrPointer_reg[25]/NET0131 , \P2_PhyAddrPointer_reg[26]/NET0131 , \P2_PhyAddrPointer_reg[27]/NET0131 , \P2_PhyAddrPointer_reg[28]/NET0131 , \P2_PhyAddrPointer_reg[29]/NET0131 , \P2_PhyAddrPointer_reg[2]/NET0131 , \P2_PhyAddrPointer_reg[30]/NET0131 , \P2_PhyAddrPointer_reg[31]/NET0131 , \P2_PhyAddrPointer_reg[3]/NET0131 , \P2_PhyAddrPointer_reg[4]/NET0131 , \P2_PhyAddrPointer_reg[5]/NET0131 , \P2_PhyAddrPointer_reg[6]/NET0131 , \P2_PhyAddrPointer_reg[7]/NET0131 , \P2_PhyAddrPointer_reg[8]/NET0131 , \P2_PhyAddrPointer_reg[9]/NET0131 , \P2_ReadRequest_reg/NET0131 , \P2_RequestPending_reg/NET0131 , \P2_State2_reg[0]/NET0131 , \P2_State2_reg[1]/NET0131 , \P2_State2_reg[2]/NET0131 , \P2_State2_reg[3]/NET0131 , \P2_State_reg[0]/NET0131 , \P2_State_reg[1]/NET0131 , \P2_State_reg[2]/NET0131 , \P2_W_R_n_reg/NET0131 , \P2_lWord_reg[0]/NET0131 , \P2_lWord_reg[10]/NET0131 , \P2_lWord_reg[11]/NET0131 , \P2_lWord_reg[12]/NET0131 , \P2_lWord_reg[13]/NET0131 , \P2_lWord_reg[14]/NET0131 , \P2_lWord_reg[15]/NET0131 , \P2_lWord_reg[1]/NET0131 , \P2_lWord_reg[2]/NET0131 , \P2_lWord_reg[3]/NET0131 , \P2_lWord_reg[4]/NET0131 , \P2_lWord_reg[5]/NET0131 , \P2_lWord_reg[6]/NET0131 , \P2_lWord_reg[7]/NET0131 , \P2_lWord_reg[8]/NET0131 , \P2_lWord_reg[9]/NET0131 , \P2_rEIP_reg[0]/NET0131 , \P2_rEIP_reg[10]/NET0131 , \P2_rEIP_reg[11]/NET0131 , \P2_rEIP_reg[12]/NET0131 , \P2_rEIP_reg[13]/NET0131 , \P2_rEIP_reg[14]/NET0131 , \P2_rEIP_reg[15]/NET0131 , \P2_rEIP_reg[16]/NET0131 , \P2_rEIP_reg[17]/NET0131 , \P2_rEIP_reg[18]/NET0131 , \P2_rEIP_reg[19]/NET0131 , \P2_rEIP_reg[1]/NET0131 , \P2_rEIP_reg[20]/NET0131 , \P2_rEIP_reg[21]/NET0131 , \P2_rEIP_reg[22]/NET0131 , \P2_rEIP_reg[23]/NET0131 , \P2_rEIP_reg[24]/NET0131 , \P2_rEIP_reg[25]/NET0131 , \P2_rEIP_reg[26]/NET0131 , \P2_rEIP_reg[27]/NET0131 , \P2_rEIP_reg[28]/NET0131 , \P2_rEIP_reg[29]/NET0131 , \P2_rEIP_reg[2]/NET0131 , \P2_rEIP_reg[30]/NET0131 , \P2_rEIP_reg[31]/NET0131 , \P2_rEIP_reg[3]/NET0131 , \P2_rEIP_reg[4]/NET0131 , \P2_rEIP_reg[5]/NET0131 , \P2_rEIP_reg[6]/NET0131 , \P2_rEIP_reg[7]/NET0131 , \P2_rEIP_reg[8]/NET0131 , \P2_rEIP_reg[9]/NET0131 , \P2_uWord_reg[0]/NET0131 , \P2_uWord_reg[10]/NET0131 , \P2_uWord_reg[11]/NET0131 , \P2_uWord_reg[12]/NET0131 , \P2_uWord_reg[13]/NET0131 , \P2_uWord_reg[14]/NET0131 , \P2_uWord_reg[1]/NET0131 , \P2_uWord_reg[2]/NET0131 , \P2_uWord_reg[3]/NET0131 , \P2_uWord_reg[4]/NET0131 , \P2_uWord_reg[5]/NET0131 , \P2_uWord_reg[6]/NET0131 , \P2_uWord_reg[7]/NET0131 , \P2_uWord_reg[8]/NET0131 , \P2_uWord_reg[9]/NET0131 , \P3_Address_reg[0]/NET0131 , \P3_Address_reg[10]/NET0131 , \P3_Address_reg[11]/NET0131 , \P3_Address_reg[12]/NET0131 , \P3_Address_reg[13]/NET0131 , \P3_Address_reg[14]/NET0131 , \P3_Address_reg[15]/NET0131 , \P3_Address_reg[16]/NET0131 , \P3_Address_reg[17]/NET0131 , \P3_Address_reg[18]/NET0131 , \P3_Address_reg[19]/NET0131 , \P3_Address_reg[1]/NET0131 , \P3_Address_reg[20]/NET0131 , \P3_Address_reg[21]/NET0131 , \P3_Address_reg[22]/NET0131 , \P3_Address_reg[23]/NET0131 , \P3_Address_reg[24]/NET0131 , \P3_Address_reg[25]/NET0131 , \P3_Address_reg[26]/NET0131 , \P3_Address_reg[27]/NET0131 , \P3_Address_reg[28]/NET0131 , \P3_Address_reg[29]/NET0131 , \P3_Address_reg[2]/NET0131 , \P3_Address_reg[3]/NET0131 , \P3_Address_reg[4]/NET0131 , \P3_Address_reg[5]/NET0131 , \P3_Address_reg[6]/NET0131 , \P3_Address_reg[7]/NET0131 , \P3_Address_reg[8]/NET0131 , \P3_Address_reg[9]/NET0131 , \P3_BE_n_reg[0]/NET0131 , \P3_BE_n_reg[1]/NET0131 , \P3_BE_n_reg[2]/NET0131 , \P3_BE_n_reg[3]/NET0131 , \P3_ByteEnable_reg[0]/NET0131 , \P3_ByteEnable_reg[1]/NET0131 , \P3_ByteEnable_reg[2]/NET0131 , \P3_ByteEnable_reg[3]/NET0131 , \P3_CodeFetch_reg/NET0131 , \P3_DataWidth_reg[0]/NET0131 , \P3_DataWidth_reg[1]/NET0131 , \P3_EAX_reg[0]/NET0131 , \P3_EAX_reg[10]/NET0131 , \P3_EAX_reg[11]/NET0131 , \P3_EAX_reg[12]/NET0131 , \P3_EAX_reg[13]/NET0131 , \P3_EAX_reg[14]/NET0131 , \P3_EAX_reg[15]/NET0131 , \P3_EAX_reg[16]/NET0131 , \P3_EAX_reg[17]/NET0131 , \P3_EAX_reg[18]/NET0131 , \P3_EAX_reg[19]/NET0131 , \P3_EAX_reg[1]/NET0131 , \P3_EAX_reg[20]/NET0131 , \P3_EAX_reg[21]/NET0131 , \P3_EAX_reg[22]/NET0131 , \P3_EAX_reg[23]/NET0131 , \P3_EAX_reg[24]/NET0131 , \P3_EAX_reg[25]/NET0131 , \P3_EAX_reg[26]/NET0131 , \P3_EAX_reg[27]/NET0131 , \P3_EAX_reg[28]/NET0131 , \P3_EAX_reg[29]/NET0131 , \P3_EAX_reg[2]/NET0131 , \P3_EAX_reg[30]/NET0131 , \P3_EAX_reg[31]/NET0131 , \P3_EAX_reg[3]/NET0131 , \P3_EAX_reg[4]/NET0131 , \P3_EAX_reg[5]/NET0131 , \P3_EAX_reg[6]/NET0131 , \P3_EAX_reg[7]/NET0131 , \P3_EAX_reg[8]/NET0131 , \P3_EAX_reg[9]/NET0131 , \P3_EBX_reg[0]/NET0131 , \P3_EBX_reg[10]/NET0131 , \P3_EBX_reg[11]/NET0131 , \P3_EBX_reg[12]/NET0131 , \P3_EBX_reg[13]/NET0131 , \P3_EBX_reg[14]/NET0131 , \P3_EBX_reg[15]/NET0131 , \P3_EBX_reg[16]/NET0131 , \P3_EBX_reg[17]/NET0131 , \P3_EBX_reg[18]/NET0131 , \P3_EBX_reg[19]/NET0131 , \P3_EBX_reg[1]/NET0131 , \P3_EBX_reg[20]/NET0131 , \P3_EBX_reg[21]/NET0131 , \P3_EBX_reg[22]/NET0131 , \P3_EBX_reg[23]/NET0131 , \P3_EBX_reg[24]/NET0131 , \P3_EBX_reg[25]/NET0131 , \P3_EBX_reg[26]/NET0131 , \P3_EBX_reg[27]/NET0131 , \P3_EBX_reg[28]/NET0131 , \P3_EBX_reg[29]/NET0131 , \P3_EBX_reg[2]/NET0131 , \P3_EBX_reg[30]/NET0131 , \P3_EBX_reg[31]/NET0131 , \P3_EBX_reg[3]/NET0131 , \P3_EBX_reg[4]/NET0131 , \P3_EBX_reg[5]/NET0131 , \P3_EBX_reg[6]/NET0131 , \P3_EBX_reg[7]/NET0131 , \P3_EBX_reg[8]/NET0131 , \P3_EBX_reg[9]/NET0131 , \P3_Flush_reg/NET0131 , \P3_InstAddrPointer_reg[0]/NET0131 , \P3_InstAddrPointer_reg[10]/NET0131 , \P3_InstAddrPointer_reg[11]/NET0131 , \P3_InstAddrPointer_reg[12]/NET0131 , \P3_InstAddrPointer_reg[13]/NET0131 , \P3_InstAddrPointer_reg[14]/NET0131 , \P3_InstAddrPointer_reg[15]/NET0131 , \P3_InstAddrPointer_reg[16]/NET0131 , \P3_InstAddrPointer_reg[17]/NET0131 , \P3_InstAddrPointer_reg[18]/NET0131 , \P3_InstAddrPointer_reg[19]/NET0131 , \P3_InstAddrPointer_reg[1]/NET0131 , \P3_InstAddrPointer_reg[20]/NET0131 , \P3_InstAddrPointer_reg[21]/NET0131 , \P3_InstAddrPointer_reg[22]/NET0131 , \P3_InstAddrPointer_reg[23]/NET0131 , \P3_InstAddrPointer_reg[24]/NET0131 , \P3_InstAddrPointer_reg[25]/NET0131 , \P3_InstAddrPointer_reg[26]/NET0131 , \P3_InstAddrPointer_reg[27]/NET0131 , \P3_InstAddrPointer_reg[28]/NET0131 , \P3_InstAddrPointer_reg[29]/NET0131 , \P3_InstAddrPointer_reg[2]/NET0131 , \P3_InstAddrPointer_reg[30]/NET0131 , \P3_InstAddrPointer_reg[31]/NET0131 , \P3_InstAddrPointer_reg[3]/NET0131 , \P3_InstAddrPointer_reg[4]/NET0131 , \P3_InstAddrPointer_reg[5]/NET0131 , \P3_InstAddrPointer_reg[6]/NET0131 , \P3_InstAddrPointer_reg[7]/NET0131 , \P3_InstAddrPointer_reg[8]/NET0131 , \P3_InstAddrPointer_reg[9]/NET0131 , \P3_InstQueueRd_Addr_reg[0]/NET0131 , \P3_InstQueueRd_Addr_reg[1]/NET0131 , \P3_InstQueueRd_Addr_reg[2]/NET0131 , \P3_InstQueueRd_Addr_reg[3]/NET0131 , \P3_InstQueueWr_Addr_reg[0]/NET0131 , \P3_InstQueueWr_Addr_reg[1]/NET0131 , \P3_InstQueueWr_Addr_reg[2]/NET0131 , \P3_InstQueueWr_Addr_reg[3]/NET0131 , \P3_InstQueue_reg[0][0]/NET0131 , \P3_InstQueue_reg[0][1]/NET0131 , \P3_InstQueue_reg[0][2]/NET0131 , \P3_InstQueue_reg[0][3]/NET0131 , \P3_InstQueue_reg[0][4]/NET0131 , \P3_InstQueue_reg[0][5]/NET0131 , \P3_InstQueue_reg[0][6]/NET0131 , \P3_InstQueue_reg[0][7]/NET0131 , \P3_InstQueue_reg[10][0]/NET0131 , \P3_InstQueue_reg[10][1]/NET0131 , \P3_InstQueue_reg[10][2]/NET0131 , \P3_InstQueue_reg[10][3]/NET0131 , \P3_InstQueue_reg[10][4]/NET0131 , \P3_InstQueue_reg[10][5]/NET0131 , \P3_InstQueue_reg[10][6]/NET0131 , \P3_InstQueue_reg[10][7]/NET0131 , \P3_InstQueue_reg[11][0]/NET0131 , \P3_InstQueue_reg[11][1]/NET0131 , \P3_InstQueue_reg[11][2]/NET0131 , \P3_InstQueue_reg[11][3]/NET0131 , \P3_InstQueue_reg[11][4]/NET0131 , \P3_InstQueue_reg[11][5]/NET0131 , \P3_InstQueue_reg[11][6]/NET0131 , \P3_InstQueue_reg[11][7]/NET0131 , \P3_InstQueue_reg[12][0]/NET0131 , \P3_InstQueue_reg[12][1]/NET0131 , \P3_InstQueue_reg[12][2]/NET0131 , \P3_InstQueue_reg[12][3]/NET0131 , \P3_InstQueue_reg[12][4]/NET0131 , \P3_InstQueue_reg[12][5]/NET0131 , \P3_InstQueue_reg[12][6]/NET0131 , \P3_InstQueue_reg[12][7]/NET0131 , \P3_InstQueue_reg[13][0]/NET0131 , \P3_InstQueue_reg[13][1]/NET0131 , \P3_InstQueue_reg[13][2]/NET0131 , \P3_InstQueue_reg[13][3]/NET0131 , \P3_InstQueue_reg[13][4]/NET0131 , \P3_InstQueue_reg[13][5]/NET0131 , \P3_InstQueue_reg[13][6]/NET0131 , \P3_InstQueue_reg[13][7]/NET0131 , \P3_InstQueue_reg[14][0]/NET0131 , \P3_InstQueue_reg[14][1]/NET0131 , \P3_InstQueue_reg[14][2]/NET0131 , \P3_InstQueue_reg[14][3]/NET0131 , \P3_InstQueue_reg[14][4]/NET0131 , \P3_InstQueue_reg[14][5]/NET0131 , \P3_InstQueue_reg[14][6]/NET0131 , \P3_InstQueue_reg[14][7]/NET0131 , \P3_InstQueue_reg[15][0]/NET0131 , \P3_InstQueue_reg[15][1]/NET0131 , \P3_InstQueue_reg[15][2]/NET0131 , \P3_InstQueue_reg[15][3]/NET0131 , \P3_InstQueue_reg[15][4]/NET0131 , \P3_InstQueue_reg[15][5]/NET0131 , \P3_InstQueue_reg[15][6]/NET0131 , \P3_InstQueue_reg[15][7]/NET0131 , \P3_InstQueue_reg[1][0]/NET0131 , \P3_InstQueue_reg[1][1]/NET0131 , \P3_InstQueue_reg[1][2]/NET0131 , \P3_InstQueue_reg[1][3]/NET0131 , \P3_InstQueue_reg[1][4]/NET0131 , \P3_InstQueue_reg[1][5]/NET0131 , \P3_InstQueue_reg[1][6]/NET0131 , \P3_InstQueue_reg[1][7]/NET0131 , \P3_InstQueue_reg[2][0]/NET0131 , \P3_InstQueue_reg[2][1]/NET0131 , \P3_InstQueue_reg[2][2]/NET0131 , \P3_InstQueue_reg[2][3]/NET0131 , \P3_InstQueue_reg[2][4]/NET0131 , \P3_InstQueue_reg[2][5]/NET0131 , \P3_InstQueue_reg[2][6]/NET0131 , \P3_InstQueue_reg[2][7]/NET0131 , \P3_InstQueue_reg[3][0]/NET0131 , \P3_InstQueue_reg[3][1]/NET0131 , \P3_InstQueue_reg[3][2]/NET0131 , \P3_InstQueue_reg[3][3]/NET0131 , \P3_InstQueue_reg[3][4]/NET0131 , \P3_InstQueue_reg[3][5]/NET0131 , \P3_InstQueue_reg[3][6]/NET0131 , \P3_InstQueue_reg[3][7]/NET0131 , \P3_InstQueue_reg[4][0]/NET0131 , \P3_InstQueue_reg[4][1]/NET0131 , \P3_InstQueue_reg[4][2]/NET0131 , \P3_InstQueue_reg[4][3]/NET0131 , \P3_InstQueue_reg[4][4]/NET0131 , \P3_InstQueue_reg[4][5]/NET0131 , \P3_InstQueue_reg[4][6]/NET0131 , \P3_InstQueue_reg[4][7]/NET0131 , \P3_InstQueue_reg[5][0]/NET0131 , \P3_InstQueue_reg[5][1]/NET0131 , \P3_InstQueue_reg[5][2]/NET0131 , \P3_InstQueue_reg[5][3]/NET0131 , \P3_InstQueue_reg[5][4]/NET0131 , \P3_InstQueue_reg[5][5]/NET0131 , \P3_InstQueue_reg[5][6]/NET0131 , \P3_InstQueue_reg[5][7]/NET0131 , \P3_InstQueue_reg[6][0]/NET0131 , \P3_InstQueue_reg[6][1]/NET0131 , \P3_InstQueue_reg[6][2]/NET0131 , \P3_InstQueue_reg[6][3]/NET0131 , \P3_InstQueue_reg[6][4]/NET0131 , \P3_InstQueue_reg[6][5]/NET0131 , \P3_InstQueue_reg[6][6]/NET0131 , \P3_InstQueue_reg[6][7]/NET0131 , \P3_InstQueue_reg[7][0]/NET0131 , \P3_InstQueue_reg[7][1]/NET0131 , \P3_InstQueue_reg[7][2]/NET0131 , \P3_InstQueue_reg[7][3]/NET0131 , \P3_InstQueue_reg[7][4]/NET0131 , \P3_InstQueue_reg[7][5]/NET0131 , \P3_InstQueue_reg[7][6]/NET0131 , \P3_InstQueue_reg[7][7]/NET0131 , \P3_InstQueue_reg[8][0]/NET0131 , \P3_InstQueue_reg[8][1]/NET0131 , \P3_InstQueue_reg[8][2]/NET0131 , \P3_InstQueue_reg[8][3]/NET0131 , \P3_InstQueue_reg[8][4]/NET0131 , \P3_InstQueue_reg[8][5]/NET0131 , \P3_InstQueue_reg[8][6]/NET0131 , \P3_InstQueue_reg[8][7]/NET0131 , \P3_InstQueue_reg[9][0]/NET0131 , \P3_InstQueue_reg[9][1]/NET0131 , \P3_InstQueue_reg[9][2]/NET0131 , \P3_InstQueue_reg[9][3]/NET0131 , \P3_InstQueue_reg[9][4]/NET0131 , \P3_InstQueue_reg[9][5]/NET0131 , \P3_InstQueue_reg[9][6]/NET0131 , \P3_InstQueue_reg[9][7]/NET0131 , \P3_MemoryFetch_reg/NET0131 , \P3_More_reg/NET0131 , \P3_PhyAddrPointer_reg[0]/NET0131 , \P3_PhyAddrPointer_reg[10]/NET0131 , \P3_PhyAddrPointer_reg[11]/NET0131 , \P3_PhyAddrPointer_reg[12]/NET0131 , \P3_PhyAddrPointer_reg[13]/NET0131 , \P3_PhyAddrPointer_reg[14]/NET0131 , \P3_PhyAddrPointer_reg[15]/NET0131 , \P3_PhyAddrPointer_reg[16]/NET0131 , \P3_PhyAddrPointer_reg[17]/NET0131 , \P3_PhyAddrPointer_reg[18]/NET0131 , \P3_PhyAddrPointer_reg[19]/NET0131 , \P3_PhyAddrPointer_reg[1]/NET0131 , \P3_PhyAddrPointer_reg[20]/NET0131 , \P3_PhyAddrPointer_reg[21]/NET0131 , \P3_PhyAddrPointer_reg[22]/NET0131 , \P3_PhyAddrPointer_reg[23]/NET0131 , \P3_PhyAddrPointer_reg[24]/NET0131 , \P3_PhyAddrPointer_reg[25]/NET0131 , \P3_PhyAddrPointer_reg[26]/NET0131 , \P3_PhyAddrPointer_reg[27]/NET0131 , \P3_PhyAddrPointer_reg[28]/NET0131 , \P3_PhyAddrPointer_reg[29]/NET0131 , \P3_PhyAddrPointer_reg[2]/NET0131 , \P3_PhyAddrPointer_reg[30]/NET0131 , \P3_PhyAddrPointer_reg[31]/NET0131 , \P3_PhyAddrPointer_reg[3]/NET0131 , \P3_PhyAddrPointer_reg[4]/NET0131 , \P3_PhyAddrPointer_reg[5]/NET0131 , \P3_PhyAddrPointer_reg[6]/NET0131 , \P3_PhyAddrPointer_reg[7]/NET0131 , \P3_PhyAddrPointer_reg[8]/NET0131 , \P3_PhyAddrPointer_reg[9]/NET0131 , \P3_ReadRequest_reg/NET0131 , \P3_RequestPending_reg/NET0131 , \P3_State2_reg[0]/NET0131 , \P3_State2_reg[1]/NET0131 , \P3_State2_reg[2]/NET0131 , \P3_State2_reg[3]/NET0131 , \P3_State_reg[0]/NET0131 , \P3_State_reg[1]/NET0131 , \P3_State_reg[2]/NET0131 , \P3_lWord_reg[0]/NET0131 , \P3_lWord_reg[10]/NET0131 , \P3_lWord_reg[11]/NET0131 , \P3_lWord_reg[12]/NET0131 , \P3_lWord_reg[13]/NET0131 , \P3_lWord_reg[14]/NET0131 , \P3_lWord_reg[15]/NET0131 , \P3_lWord_reg[1]/NET0131 , \P3_lWord_reg[2]/NET0131 , \P3_lWord_reg[3]/NET0131 , \P3_lWord_reg[4]/NET0131 , \P3_lWord_reg[5]/NET0131 , \P3_lWord_reg[6]/NET0131 , \P3_lWord_reg[7]/NET0131 , \P3_lWord_reg[8]/NET0131 , \P3_lWord_reg[9]/NET0131 , \P3_rEIP_reg[0]/NET0131 , \P3_rEIP_reg[10]/NET0131 , \P3_rEIP_reg[11]/NET0131 , \P3_rEIP_reg[12]/NET0131 , \P3_rEIP_reg[13]/NET0131 , \P3_rEIP_reg[14]/NET0131 , \P3_rEIP_reg[15]/NET0131 , \P3_rEIP_reg[16]/NET0131 , \P3_rEIP_reg[17]/NET0131 , \P3_rEIP_reg[18]/NET0131 , \P3_rEIP_reg[19]/NET0131 , \P3_rEIP_reg[1]/NET0131 , \P3_rEIP_reg[20]/NET0131 , \P3_rEIP_reg[21]/NET0131 , \P3_rEIP_reg[22]/NET0131 , \P3_rEIP_reg[23]/NET0131 , \P3_rEIP_reg[24]/NET0131 , \P3_rEIP_reg[25]/NET0131 , \P3_rEIP_reg[26]/NET0131 , \P3_rEIP_reg[27]/NET0131 , \P3_rEIP_reg[28]/NET0131 , \P3_rEIP_reg[29]/NET0131 , \P3_rEIP_reg[2]/NET0131 , \P3_rEIP_reg[30]/NET0131 , \P3_rEIP_reg[31]/NET0131 , \P3_rEIP_reg[3]/NET0131 , \P3_rEIP_reg[4]/NET0131 , \P3_rEIP_reg[5]/NET0131 , \P3_rEIP_reg[6]/NET0131 , \P3_rEIP_reg[7]/NET0131 , \P3_rEIP_reg[8]/NET0131 , \P3_rEIP_reg[9]/NET0131 , \P3_uWord_reg[0]/NET0131 , \P3_uWord_reg[10]/NET0131 , \P3_uWord_reg[11]/NET0131 , \P3_uWord_reg[12]/NET0131 , \P3_uWord_reg[13]/NET0131 , \P3_uWord_reg[14]/NET0131 , \P3_uWord_reg[1]/NET0131 , \P3_uWord_reg[2]/NET0131 , \P3_uWord_reg[3]/NET0131 , \P3_uWord_reg[4]/NET0131 , \P3_uWord_reg[5]/NET0131 , \P3_uWord_reg[6]/NET0131 , \P3_uWord_reg[7]/NET0131 , \P3_uWord_reg[8]/NET0131 , \P3_uWord_reg[9]/NET0131 , \address1[0]_pad , \address1[10]_pad , \address1[11]_pad , \address1[12]_pad , \address1[13]_pad , \address1[14]_pad , \address1[15]_pad , \address1[16]_pad , \address1[17]_pad , \address1[18]_pad , \address1[19]_pad , \address1[1]_pad , \address1[20]_pad , \address1[21]_pad , \address1[22]_pad , \address1[23]_pad , \address1[24]_pad , \address1[25]_pad , \address1[26]_pad , \address1[27]_pad , \address1[28]_pad , \address1[29]_pad , \address1[2]_pad , \address1[3]_pad , \address1[4]_pad , \address1[5]_pad , \address1[6]_pad , \address1[7]_pad , \address1[8]_pad , \address1[9]_pad , \ast1_pad , \ast2_pad , \bs16_pad , \buf1_reg[0]/NET0131 , \buf1_reg[10]/NET0131 , \buf1_reg[11]/NET0131 , \buf1_reg[12]/NET0131 , \buf1_reg[13]/NET0131 , \buf1_reg[14]/NET0131 , \buf1_reg[15]/NET0131 , \buf1_reg[16]/NET0131 , \buf1_reg[17]/NET0131 , \buf1_reg[18]/NET0131 , \buf1_reg[19]/NET0131 , \buf1_reg[1]/NET0131 , \buf1_reg[20]/NET0131 , \buf1_reg[21]/NET0131 , \buf1_reg[22]/NET0131 , \buf1_reg[23]/NET0131 , \buf1_reg[24]/NET0131 , \buf1_reg[25]/NET0131 , \buf1_reg[26]/NET0131 , \buf1_reg[27]/NET0131 , \buf1_reg[28]/NET0131 , \buf1_reg[29]/NET0131 , \buf1_reg[2]/NET0131 , \buf1_reg[30]/NET0131 , \buf1_reg[3]/NET0131 , \buf1_reg[4]/NET0131 , \buf1_reg[5]/NET0131 , \buf1_reg[6]/NET0131 , \buf1_reg[7]/NET0131 , \buf1_reg[8]/NET0131 , \buf1_reg[9]/NET0131 , \buf2_reg[0]/NET0131 , \buf2_reg[10]/NET0131 , \buf2_reg[11]/NET0131 , \buf2_reg[12]/NET0131 , \buf2_reg[13]/NET0131 , \buf2_reg[14]/NET0131 , \buf2_reg[15]/NET0131 , \buf2_reg[16]/NET0131 , \buf2_reg[17]/NET0131 , \buf2_reg[18]/NET0131 , \buf2_reg[19]/NET0131 , \buf2_reg[1]/NET0131 , \buf2_reg[20]/NET0131 , \buf2_reg[21]/NET0131 , \buf2_reg[22]/NET0131 , \buf2_reg[23]/NET0131 , \buf2_reg[24]/NET0131 , \buf2_reg[25]/NET0131 , \buf2_reg[26]/NET0131 , \buf2_reg[27]/NET0131 , \buf2_reg[28]/NET0131 , \buf2_reg[29]/NET0131 , \buf2_reg[2]/NET0131 , \buf2_reg[30]/NET0131 , \buf2_reg[3]/NET0131 , \buf2_reg[4]/NET0131 , \buf2_reg[5]/NET0131 , \buf2_reg[6]/NET0131 , \buf2_reg[7]/NET0131 , \buf2_reg[8]/NET0131 , \buf2_reg[9]/NET0131 , \datai[0]_pad , \datai[10]_pad , \datai[11]_pad , \datai[12]_pad , \datai[13]_pad , \datai[14]_pad , \datai[15]_pad , \datai[16]_pad , \datai[17]_pad , \datai[18]_pad , \datai[19]_pad , \datai[1]_pad , \datai[20]_pad , \datai[21]_pad , \datai[22]_pad , \datai[23]_pad , \datai[24]_pad , \datai[25]_pad , \datai[26]_pad , \datai[27]_pad , \datai[28]_pad , \datai[29]_pad , \datai[2]_pad , \datai[30]_pad , \datai[31]_pad , \datai[3]_pad , \datai[4]_pad , \datai[5]_pad , \datai[6]_pad , \datai[7]_pad , \datai[8]_pad , \datai[9]_pad , \datao[0]_pad , \datao[10]_pad , \datao[11]_pad , \datao[12]_pad , \datao[13]_pad , \datao[14]_pad , \datao[15]_pad , \datao[16]_pad , \datao[17]_pad , \datao[18]_pad , \datao[19]_pad , \datao[1]_pad , \datao[20]_pad , \datao[21]_pad , \datao[22]_pad , \datao[23]_pad , \datao[24]_pad , \datao[25]_pad , \datao[26]_pad , \datao[27]_pad , \datao[28]_pad , \datao[29]_pad , \datao[2]_pad , \datao[30]_pad , \datao[3]_pad , \datao[4]_pad , \datao[5]_pad , \datao[6]_pad , \datao[7]_pad , \datao[8]_pad , \datao[9]_pad , dc_pad, hold_pad, mio_pad, na_pad, \ready11_reg/NET0131 , \ready12_reg/NET0131 , \ready1_pad , \ready21_reg/NET0131 , \ready22_reg/NET0131 , \ready2_pad , wr_pad, \_al_n0 , \_al_n1 , \address2[0]_pad , \address2[10]_pad , \address2[11]_pad , \address2[12]_pad , \address2[13]_pad , \address2[14]_pad , \address2[15]_pad , \address2[16]_pad , \address2[17]_pad , \address2[18]_pad , \address2[19]_pad , \address2[1]_pad , \address2[20]_pad , \address2[21]_pad , \address2[22]_pad , \address2[23]_pad , \address2[24]_pad , \address2[25]_pad , \address2[26]_pad , \address2[27]_pad , \address2[28]_pad , \address2[29]_pad , \address2[2]_pad , \address2[3]_pad , \address2[4]_pad , \address2[5]_pad , \address2[6]_pad , \address2[7]_pad , \address2[8]_pad , \address2[9]_pad , \g133468/_2_ , \g133469/_2_ , \g133470/_2_ , \g133475/_0_ , \g133476/_2_ , \g133515/_0_ , \g133516/_0_ , \g133517/_0_ , \g133518/_0_ , \g133523/_0_ , \g133524/_0_ , \g133528/_0_ , \g133529/_0_ , \g133531/_0_ , \g133532/_0_ , \g133533/_0_ , \g133534/_0_ , \g133535/_0_ , \g133536/_0_ , \g133537/_0_ , \g133538/_0_ , \g133539/_0_ , \g133540/_0_ , \g133541/_0_ , \g133542/_0_ , \g133543/_0_ , \g133544/_0_ , \g133545/_0_ , \g133546/_0_ , \g133547/_0_ , \g133548/_0_ , \g133549/_0_ , \g133550/_0_ , \g133551/_0_ , \g133552/_0_ , \g133553/_0_ , \g133554/_0_ , \g133555/_0_ , \g133556/_0_ , \g133557/_0_ , \g133558/_0_ , \g133559/_0_ , \g133560/_0_ , \g133561/_0_ , \g133566/_0_ , \g133619/_0_ , \g133659/_0_ , \g133660/_0_ , \g133662/_0_ , \g133663/_0_ , \g133664/_0_ , \g133665/_0_ , \g133666/_0_ , \g133667/_0_ , \g133668/_0_ , \g133669/_0_ , \g133670/_0_ , \g133671/_0_ , \g133672/_0_ , \g133673/_0_ , \g133674/_0_ , \g133675/_0_ , \g133676/_0_ , \g133677/_0_ , \g133678/_0_ , \g133679/_0_ , \g133680/_0_ , \g133681/_0_ , \g133682/_0_ , \g133683/_0_ , \g133684/_0_ , \g133685/_0_ , \g133686/_0_ , \g133687/_0_ , \g133688/_0_ , \g133689/_0_ , \g133690/_0_ , \g133691/_0_ , \g133694/_0_ , \g133697/_0_ , \g133702/_0_ , \g133703/_0_ , \g133756/_0_ , \g133792/_0_ , \g133793/_0_ , \g133794/_0_ , \g133796/_0_ , \g133797/_0_ , \g133798/_0_ , \g133799/_0_ , \g133800/_0_ , \g133801/_0_ , \g133802/_0_ , \g133803/_0_ , \g133804/_0_ , \g133806/_0_ , \g133807/_0_ , \g133808/_0_ , \g133812/_0_ , \g133813/_0_ , \g133814/_0_ , \g133817/_0_ , \g133821/_0_ , \g133824/_0_ , \g133826/_0_ , \g133828/_0_ , \g133864/_0_ , \g133865/_0_ , \g133867/_0_ , \g133868/_0_ , \g133869/_0_ , \g133871/_0_ , \g133872/_0_ , \g133873/_0_ , \g133874/_0_ , \g133875/_0_ , \g133876/_0_ , \g133877/_0_ , \g133878/_0_ , \g133879/_0_ , \g133881/_0_ , \g133882/_0_ , \g133883/_0_ , \g133884/_0_ , \g133885/_0_ , \g133886/_0_ , \g133887/_0_ , \g133888/_0_ , \g133889/_0_ , \g133890/_0_ , \g133891/_0_ , \g133892/_0_ , \g133893/_0_ , \g133894/_0_ , \g133895/_0_ , \g133896/_0_ , \g133897/_0_ , \g133898/_0_ , \g133910/_0_ , \g133911/_0_ , \g133912/_0_ , \g133915/_0_ , \g133917/_0_ , \g133929/_0_ , \g134014/_0_ , \g134040/_0_ , \g134041/_0_ , \g134042/_0_ , \g134043/_0_ , \g134044/_0_ , \g134045/_0_ , \g134046/_0_ , \g134047/_0_ , \g134048/_0_ , \g134049/_0_ , \g134050/_0_ , \g134051/_0_ , \g134052/_0_ , \g134053/_0_ , \g134054/_0_ , \g134056/_0_ , \g134059/_0_ , \g134064/_0_ , \g134067/_0_ , \g134068/_0_ , \g134069/_0_ , \g134070/_0_ , \g134071/_0_ , \g134073/_0_ , \g134076/_0_ , \g134131/_0_ , \g134132/_0_ , \g134156/_0_ , \g134157/_0_ , \g134158/_0_ , \g134159/_0_ , \g134163/_0_ , \g134164/_0_ , \g134165/_0_ , \g134166/_0_ , \g134167/_0_ , \g134168/_0_ , \g134169/_0_ , \g134170/_0_ , \g134171/_0_ , \g134172/_0_ , \g134173/_0_ , \g134174/_0_ , \g134176/_0_ , \g134177/_0_ , \g134178/_0_ , \g134179/_0_ , \g134181/_0_ , \g134183/_0_ , \g134184/_0_ , \g134185/_0_ , \g134186/_0_ , \g134187/_0_ , \g134188/_0_ , \g134189/_0_ , \g134190/_0_ , \g134191/_0_ , \g134194/_0_ , \g134202/_0_ , \g134207/_0_ , \g134214/_0_ , \g134216/_0_ , \g134226/_0_ , \g134228/_0_ , \g134360/_0_ , \g134383/_0_ , \g134412/_0_ , \g134413/_0_ , \g134419/_0_ , \g134420/_0_ , \g134421/_0_ , \g134422/_0_ , \g134423/_0_ , \g134424/_0_ , \g134426/_0_ , \g134429/_0_ , \g134431/_0_ , \g134433/_0_ , \g134434/_0_ , \g134435/_0_ , \g134436/_0_ , \g134438/_0_ , \g134439/_0_ , \g134441/_0_ , \g134442/_0_ , \g134443/_0_ , \g134445/_0_ , \g134446/_0_ , \g134447/_0_ , \g134448/_0_ , \g134449/_0_ , \g134450/_0_ , \g134451/_0_ , \g134453/_0_ , \g134454/_0_ , \g134455/_0_ , \g134457/_0_ , \g134458/_0_ , \g134459/_0_ , \g134460/_0_ , \g134469/_0_ , \g134470/_0_ , \g134471/_0_ , \g134472/_0_ , \g134479/_0_ , \g134480/_0_ , \g134481/_0_ , \g134482/_0_ , \g134490/_0_ , \g134491/_0_ , \g134496/_0_ , \g134506/_0_ , \g134508/_0_ , \g134579/_0_ , \g134603/_0_ , \g134604/_0_ , \g134605/_0_ , \g134606/_0_ , \g134607/_0_ , \g134608/_0_ , \g134609/_0_ , \g134610/_0_ , \g134611/_0_ , \g134612/_0_ , \g134613/_0_ , \g134614/_0_ , \g134615/_0_ , \g134616/_0_ , \g134617/_0_ , \g134618/_0_ , \g134619/_0_ , \g134620/_0_ , \g134621/_0_ , \g134632/_0_ , \g134633/_0_ , \g134636/_0_ , \g134637/_0_ , \g134638/_0_ , \g134639/_0_ , \g134645/_0_ , \g134646/_0_ , \g134648/_0_ , \g134649/_0_ , \g134650/_0_ , \g134651/_0_ , \g134652/_0_ , \g134656/_0_ , \g134657/_0_ , \g134658/_0_ , \g134664/_0_ , \g134665/_0_ , \g134671/_0_ , \g134672/_0_ , \g134686/_0_ , \g134687/_0_ , \g134735/_0_ , \g134908/_0_ , \g134909/_0_ , \g134910/_0_ , \g134920/_0_ , \g134921/_0_ , \g134922/_0_ , \g134923/_0_ , \g134925/_0_ , \g134926/_0_ , \g134928/_0_ , \g134929/_0_ , \g134933/_0_ , \g134934/_0_ , \g134935/_0_ , \g134936/_0_ , \g134937/_0_ , \g134938/_0_ , \g134940/_0_ , \g134941/_0_ , \g134943/_0_ , \g134945/_0_ , \g134946/_0_ , \g134947/_0_ , \g134948/_0_ , \g134949/_0_ , \g134950/_0_ , \g134959/_0_ , \g134960/_0_ , \g134961/_0_ , \g134979/_0_ , \g134980/_0_ , \g135054/_0_ , \g135061/_0_ , \g135072/_0_ , \g135100/_0_ , \g135127/_0_ , \g135128/_0_ , \g135129/_0_ , \g135130/_0_ , \g135132/_0_ , \g135133/_0_ , \g135134/_0_ , \g135135/_0_ , \g135136/_0_ , \g135137/_0_ , \g135138/_0_ , \g135139/_0_ , \g135140/_0_ , \g135141/_0_ , \g135142/_0_ , \g135145/_0_ , \g135146/_0_ , \g135151/_0_ , \g135154/_0_ , \g135155/_0_ , \g135158/_0_ , \g135163/_0_ , \g135164/_0_ , \g135165/_0_ , \g135192/_0_ , \g135197/_0_ , \g135217/_0_ , \g135225/_0_ , \g135231/_0_ , \g135272/_0_ , \g135290/_0_ , \g135291/_0_ , \g135293/_0_ , \g135294/_0_ , \g135295/_0_ , \g135296/_0_ , \g135297/_0_ , \g135412/_0_ , \g135437/_0_ , \g135438/_0_ , \g135443/_0_ , \g135444/_0_ , \g135445/_0_ , \g135446/_0_ , \g135447/_0_ , \g135448/_0_ , \g135449/_0_ , \g135450/_0_ , \g135451/_0_ , \g135452/_0_ , \g135454/_0_ , \g135455/_0_ , \g135456/_0_ , \g135457/_0_ , \g135458/_0_ , \g135463/_0_ , \g135466/_0_ , \g135473/_0_ , \g135481/_0_ , \g135497/_0_ , \g135503/_0_ , \g135505/_0_ , \g135506/_0_ , \g135557/_0_ , \g135558/_0_ , \g135569/_0_ , \g135570/_0_ , \g135571/_0_ , \g135572/_0_ , \g135573/_0_ , \g135575/_0_ , \g135578/_0_ , \g135754/_0_ , \g135755/_0_ , \g135756/_0_ , \g135767/_0_ , \g135768/_0_ , \g135769/_0_ , \g135777/_0_ , \g135778/_0_ , \g135779/_0_ , \g135872/_0_ , \g135873/_0_ , \g135875/_0_ , \g135877/_0_ , \g135878/_0_ , \g135879/_0_ , \g135880/_0_ , \g136087/_0_ , \g136118/_0_ , \g136119/_0_ , \g136120/_0_ , \g136121/_0_ , \g136122/_0_ , \g136123/_0_ , \g136124/_0_ , \g136125/_0_ , \g136126/_0_ , \g136127/_0_ , \g136128/_0_ , \g136129/_0_ , \g136130/_0_ , \g136131/_0_ , \g136132/_0_ , \g136133/_0_ , \g136172/_0_ , \g136173/_0_ , \g136174/_0_ , \g136175/_0_ , \g136177/_0_ , \g136178/_0_ , \g136242/_0_ , \g136243/_0_ , \g136244/_0_ , \g136246/_0_ , \g136248/_0_ , \g136249/_0_ , \g136250/_0_ , \g136251/_0_ , \g136252/_0_ , \g136253/_0_ , \g136254/_0_ , \g136255/_0_ , \g136256/_0_ , \g136257/_0_ , \g136258/_0_ , \g136259/_0_ , \g136260/_0_ , \g136261/_0_ , \g136262/_0_ , \g136263/_0_ , \g136264/_0_ , \g136265/_0_ , \g136266/_0_ , \g136267/_0_ , \g136268/_0_ , \g136269/_0_ , \g136270/_0_ , \g136271/_0_ , \g136272/_0_ , \g136273/_0_ , \g136274/_0_ , \g136275/_0_ , \g136276/_0_ , \g136277/_0_ , \g136279/_0_ , \g136280/_0_ , \g136281/_0_ , \g136282/_0_ , \g136283/_0_ , \g136285/_0_ , \g136286/_0_ , \g136287/_0_ , \g136288/_0_ , \g136289/_0_ , \g136290/_0_ , \g136291/_0_ , \g136292/_0_ , \g136293/_0_ , \g136295/_0_ , \g136467/_0_ , \g136468/_0_ , \g136469/_0_ , \g136470/_0_ , \g136472/_0_ , \g136473/_0_ , \g136474/_0_ , \g136476/_0_ , \g136479/_0_ , \g136480/_0_ , \g136481/_0_ , \g136482/_0_ , \g136483/_0_ , \g136484/_0_ , \g136485/_0_ , \g136486/_0_ , \g136528/_0_ , \g136529/_0_ , \g136530/_0_ , \g136531/_0_ , \g136532/_0_ , \g136533/_0_ , \g136534/_0_ , \g136535/_0_ , \g136536/_0_ , \g136537/_0_ , \g136538/_0_ , \g136539/_0_ , \g136540/_0_ , \g136541/_0_ , \g136542/_0_ , \g136543/_0_ , \g136544/_0_ , \g136545/_0_ , \g136546/_0_ , \g136547/_0_ , \g136548/_0_ , \g136549/_0_ , \g136550/_0_ , \g136551/_0_ , \g136552/_0_ , \g136553/_0_ , \g136554/_0_ , \g136555/_0_ , \g136556/_0_ , \g136557/_0_ , \g136558/_0_ , \g136559/_0_ , \g136560/_0_ , \g136561/_0_ , \g136562/_0_ , \g136563/_0_ , \g136564/_0_ , \g136565/_0_ , \g136566/_0_ , \g136567/_0_ , \g136568/_0_ , \g136570/_0_ , \g136571/_0_ , \g136572/_0_ , \g136573/_0_ , \g136574/_0_ , \g136575/_0_ , \g136576/_0_ , \g136577/_0_ , \g136578/_0_ , \g136579/_0_ , \g136580/_0_ , \g136582/_0_ , \g136583/_0_ , \g136584/_0_ , \g136585/_0_ , \g136586/_0_ , \g136587/_0_ , \g136588/_0_ , \g136589/_0_ , \g136590/_0_ , \g136591/_0_ , \g136592/_0_ , \g136593/_0_ , \g136594/_0_ , \g136595/_0_ , \g136596/_0_ , \g136597/_0_ , \g136598/_0_ , \g136599/_0_ , \g136600/_0_ , \g136601/_0_ , \g136602/_0_ , \g136603/_0_ , \g136604/_0_ , \g136605/_0_ , \g136606/_0_ , \g136607/_0_ , \g136609/_0_ , \g136610/_0_ , \g136611/_0_ , \g136616/_0_ , \g136617/_0_ , \g136618/_0_ , \g136619/_0_ , \g136626/_0_ , \g136628/_0_ , \g136646/_0_ , \g136649/_0_ , \g136662/_0_ , \g136666/_0_ , \g136695/_0_ , \g136696/_0_ , \g136699/_0_ , \g136762/_0_ , \g136763/_0_ , \g136764/_0_ , \g136765/_0_ , \g136768/_0_ , \g136769/_0_ , \g137051/_0_ , \g137052/_0_ , \g137053/_0_ , \g137054/_0_ , \g137055/_0_ , \g137056/_0_ , \g137057/_0_ , \g137060/_0_ , \g137061/_0_ , \g137063/_0_ , \g137064/_0_ , \g137065/_0_ , \g137067/_0_ , \g137069/_0_ , \g137072/_0_ , \g137073/_0_ , \g137075/_0_ , \g137111/_0_ , \g137122/_0_ , \g137133/_0_ , \g137134/_0_ , \g137135/_0_ , \g137136/_0_ , \g137137/_0_ , \g137138/_0_ , \g137144/_0_ , \g137145/_0_ , \g137146/_0_ , \g137149/_0_ , \g137234/_0_ , \g137237/_0_ , \g137238/_0_ , \g137294/_0_ , \g137295/_0_ , \g137296/_0_ , \g137297/_0_ , \g137298/_0_ , \g137299/_0_ , \g137300/_0_ , \g137301/_0_ , \g137302/_0_ , \g137303/_0_ , \g137304/_0_ , \g137305/_0_ , \g137306/_0_ , \g137307/_0_ , \g137308/_0_ , \g137309/_0_ , \g137310/_0_ , \g137311/_0_ , \g137312/_0_ , \g137313/_0_ , \g137314/_0_ , \g137315/_0_ , \g137316/_0_ , \g137317/_0_ , \g137318/_0_ , \g137319/_0_ , \g137320/_0_ , \g137321/_0_ , \g137322/_0_ , \g137323/_0_ , \g137324/_0_ , \g137325/_0_ , \g137327/_0_ , \g137328/_0_ , \g137329/_0_ , \g137330/_0_ , \g137331/_0_ , \g137332/_0_ , \g137333/_0_ , \g137334/_0_ , \g137335/_0_ , \g137336/_0_ , \g137337/_0_ , \g137338/_0_ , \g137339/_0_ , \g137340/_0_ , \g137341/_0_ , \g137342/_0_ , \g137343/_0_ , \g137344/_0_ , \g137345/_0_ , \g137346/_0_ , \g137347/_0_ , \g137349/_0_ , \g137350/_0_ , \g137351/_0_ , \g137352/_0_ , \g137353/_0_ , \g137354/_0_ , \g137448/_0_ , \g137483/_0_ , \g137484/_0_ , \g137485/_0_ , \g137486/_0_ , \g137487/_0_ , \g137488/_0_ , \g137491/_0_ , \g137492/_0_ , \g137493/_0_ , \g137494/_0_ , \g137495/_0_ , \g137496/_0_ , \g137497/_0_ , \g137499/_0_ , \g137501/_0_ , \g137502/_0_ , \g137503/_0_ , \g137504/_0_ , \g137505/_0_ , \g137506/_0_ , \g137507/_0_ , \g137508/_0_ , \g137509/_0_ , \g137511/_0_ , \g137512/_0_ , \g137513/_0_ , \g137514/_0_ , \g137515/_0_ , \g137516/_0_ , \g137517/_0_ , \g137519/_0_ , \g137520/_0_ , \g137521/_0_ , \g137524/_0_ , \g137541/_0_ , \g137547/_0_ , \g137554/_0_ , \g137559/_0_ , \g137566/_0_ , \g137571/_0_ , \g137778/_0_ , \g137782/_0_ , \g137783/_0_ , \g137784/_0_ , \g137785/_0_ , \g137786/_0_ , \g137820/_0_ , \g137821/_0_ , \g137822/_0_ , \g137823/_0_ , \g137824/_0_ , \g137825/_0_ , \g137826/_0_ , \g137827/_0_ , \g137828/_0_ , \g137829/_0_ , \g137830/_0_ , \g137831/_0_ , \g137832/_0_ , \g137833/_0_ , \g137834/_0_ , \g137835/_0_ , \g137836/_0_ , \g137837/_0_ , \g137838/_0_ , \g137839/_0_ , \g137840/_0_ , \g137841/_0_ , \g137842/_0_ , \g137843/_0_ , \g137844/_0_ , \g137845/_0_ , \g137846/_0_ , \g137847/_0_ , \g137848/_0_ , \g137849/_0_ , \g137850/_0_ , \g137851/_0_ , \g137852/_0_ , \g137853/_0_ , \g137854/_0_ , \g137855/_0_ , \g137856/_0_ , \g137857/_0_ , \g137858/_0_ , \g137859/_0_ , \g137860/_0_ , \g137861/_0_ , \g137862/_0_ , \g137863/_0_ , \g137864/_0_ , \g137865/_0_ , \g137866/_0_ , \g137867/_0_ , \g137868/_0_ , \g137869/_0_ , \g137870/_0_ , \g137871/_0_ , \g137872/_0_ , \g137873/_0_ , \g137874/_0_ , \g137875/_0_ , \g137876/_0_ , \g137877/_0_ , \g137878/_0_ , \g137879/_0_ , \g137880/_0_ , \g137881/_0_ , \g137882/_0_ , \g137883/_0_ , \g137884/_0_ , \g137885/_0_ , \g137886/_0_ , \g137887/_0_ , \g137888/_0_ , \g137889/_0_ , \g137890/_0_ , \g137891/_0_ , \g137892/_0_ , \g137893/_0_ , \g137894/_0_ , \g137895/_0_ , \g137896/_0_ , \g137897/_0_ , \g137898/_0_ , \g137899/_0_ , \g137900/_0_ , \g137901/_0_ , \g137902/_0_ , \g137903/_0_ , \g138338/_0_ , \g138340/_0_ , \g138341/_0_ , \g138346/_0_ , \g138347/_0_ , \g138375/_0_ , \g138395/_0_ , \g138396/_0_ , \g138397/_0_ , \g138398/_0_ , \g138400/_0_ , \g138401/_0_ , \g138402/_0_ , \g138403/_0_ , \g138404/_0_ , \g138405/_0_ , \g138406/_0_ , \g138407/_0_ , \g138408/_0_ , \g138409/_0_ , \g138410/_0_ , \g138411/_0_ , \g138412/_0_ , \g138419/_0_ , \g138420/_0_ , \g138421/_0_ , \g138422/_0_ , \g138423/_0_ , \g138424/_0_ , \g138425/_0_ , \g138426/_0_ , \g138427/_0_ , \g138428/_0_ , \g138429/_0_ , \g138430/_0_ , \g138431/_0_ , \g138432/_0_ , \g138433/_0_ , \g138434/_0_ , \g138435/_0_ , \g138436/_0_ , \g138437/_0_ , \g138438/_0_ , \g138439/_0_ , \g138440/_0_ , \g138441/_0_ , \g138442/_0_ , \g138443/_0_ , \g138908/_0_ , \g138909/_0_ , \g138910/_0_ , \g138914/_0_ , \g138915/_0_ , \g138917/_0_ , \g138918/_0_ , \g138919/_0_ , \g138920/_0_ , \g138921/_0_ , \g138925/_0_ , \g138926/_0_ , \g138927/_0_ , \g138930/_0_ , \g138931/_0_ , \g138932/_0_ , \g138960/_0_ , \g138962/_0_ , \g139037/_0_ , \g139038/_0_ , \g139040/_0_ , \g139043/_0_ , \g139044/_0_ , \g139045/_0_ , \g139046/_0_ , \g139047/_0_ , \g139048/_0_ , \g139049/_0_ , \g139050/_0_ , \g139051/_0_ , \g139053/_0_ , \g139054/_0_ , \g139055/_0_ , \g139056/_0_ , \g139057/_0_ , \g139058/_0_ , \g139059/_0_ , \g139060/_0_ , \g139062/_0_ , \g139063/_0_ , \g139064/_0_ , \g139099/_0_ , \g139126/_0_ , \g139127/_0_ , \g139128/_0_ , \g139129/_0_ , \g139130/_0_ , \g139131/_0_ , \g139132/_0_ , \g139133/_0_ , \g139134/_0_ , \g139135/_0_ , \g139136/_0_ , \g139137/_0_ , \g139138/_0_ , \g139139/_0_ , \g139140/_0_ , \g139141/_0_ , \g139260/_0_ , \g139263/_0_ , \g139267/_0_ , \g139270/_0_ , \g139273/_0_ , \g139276/_0_ , \g139279/_0_ , \g139283/_0_ , \g139286/_0_ , \g139289/_0_ , \g139292/_0_ , \g139295/_0_ , \g139298/_0_ , \g139302/_0_ , \g139305/_0_ , \g139309/_0_ , \g139871/_0_ , \g139872/_0_ , \g139873/_0_ , \g139874/_0_ , \g139875/_0_ , \g139876/_0_ , \g139877/_0_ , \g139878/_0_ , \g139879/_0_ , \g139880/_0_ , \g139881/_0_ , \g139882/_0_ , \g139883/_0_ , \g139884/_0_ , \g139885/_0_ , \g139886/_0_ , \g139887/_0_ , \g139888/_0_ , \g139889/_0_ , \g139890/_0_ , \g139891/_0_ , \g139892/_0_ , \g139893/_0_ , \g139895/_0_ , \g139896/_0_ , \g139899/_0_ , \g139901/_0_ , \g139902/_0_ , \g139903/_0_ , \g139904/_0_ , \g140285/_0_ , \g140288/_0_ , \g140329/_0_ , \g140774/_0_ , \g140832/_0_ , \g140834/_0_ , \g140836/_0_ , \g140838/_0_ , \g140840/_0_ , \g140842/_0_ , \g140844/_0_ , \g140846/_0_ , \g140847/_0_ , \g140848/_0_ , \g140850/_0_ , \g140851/_0_ , \g140852/_0_ , \g140853/_0_ , \g140855/_0_ , \g140857/_0_ , \g140861/_0_ , \g140923/_0_ , \g141178/_0_ , \g141179/_0_ , \g141180/_0_ , \g141480/_0_ , \g141495/_0_ , \g141497/_0_ , \g141562/_0_ , \g141563/_0_ , \g141564/_0_ , \g141589/_0_ , \g141617/_0_ , \g141618/_0_ , \g141621/_0_ , \g141625/_0_ , \g141626/_0_ , \g141630/_0_ , \g141634/_0_ , \g141638/_0_ , \g141642/_0_ , \g141646/_0_ , \g141649/_0_ , \g141651/_0_ , \g141652/_0_ , \g141655/_0_ , \g141658/_0_ , \g141661/_0_ , \g141663/_0_ , \g141664/_0_ , \g141667/_0_ , \g141671/_0_ , \g141706/_0_ , \g141976/_0_ , \g141977/_0_ , \g141994/_0_ , \g142246/_0_ , \g142247/_0_ , \g142253/_0_ , \g142689/_0_ , \g142693/_0_ , \g142701/_0_ , \g142704/_0_ , \g142707/_0_ , \g142710/_0_ , \g142713/_0_ , \g142714/_0_ , \g142717/_0_ , \g142720/_0_ , \g142723/_0_ , \g142727/_0_ , \g142734/_0_ , \g143080/_0_ , \g143081/_0_ , \g143083/_0_ , \g143149/_0_ , \g143150/_0_ , \g143153/_0_ , \g143752/_0_ , \g143753/_0_ , \g143759/_0_ , \g144242/_0_ , \g144243/_0_ , \g144244/_0_ , \g144245/_0_ , \g144246/_0_ , \g144249/_0_ , \g145699/_0_ , \g145700/_0_ , \g145702/_0_ , \g145756/_0_ , \g145757/_0_ , \g145758/_0_ , \g146850/_0_ , \g146851/_0_ , \g146864/_0_ , \g147277/_0_ , \g147278/_0_ , \g147279/_0_ , \g147304/_0_ , \g147305/_0_ , \g147306/_0_ , \g147338/_3_ , \g147339/_3_ , \g147340/_3_ , \g147341/_3_ , \g147342/_3_ , \g147343/_3_ , \g147344/_3_ , \g147345/_3_ , \g147346/_3_ , \g147347/_3_ , \g147348/_3_ , \g147349/_3_ , \g147350/_3_ , \g147351/_3_ , \g147352/_3_ , \g147353/_3_ , \g147354/_3_ , \g147355/_3_ , \g147356/_3_ , \g147357/_3_ , \g147358/_3_ , \g147359/_3_ , \g147360/_3_ , \g147362/_3_ , \g147363/_3_ , \g147364/_3_ , \g147365/_3_ , \g147366/_3_ , \g147367/_3_ , \g147368/_3_ , \g147369/_3_ , \g148630/_0_ , \g148631/_0_ , \g148676/_0_ , \g148785/_0_ , \g148788/_0_ , \g148789/_0_ , \g148834/_0_ , \g148836/_0_ , \g148838/_0_ , \g149836/_0_ , \g149837/_0_ , \g149838/_0_ , \g150142/_0_ , \g152366/_0_ , \g152367/_0_ , \g152368/_0_ , \g152426/_0_ , \g152427/_0_ , \g152428/_0_ , \g152586/_0_ , \g152587/_0_ , \g152588/_0_ , \g153217/_0_ , \g154117/_0_ , \g154118/_0_ , \g154130/_0_ , \g154269/_0_ , \g154270/_0_ , \g154284/_0_ , \g154682/_0_ , \g155004/_0_ , \g155020/_0_ , \g155121/_0_ , \g155124/_0_ , \g155126/_0_ , \g155228/_0_ , \g155229/_0_ , \g155230/_0_ , \g155326/_0_ , \g155327/_0_ , \g155330/_0_ , \g155353/_0_ , \g155354/_0_ , \g155356/_0_ , \g155602/_0_ , \g155633/_0_ , \g155634/_0_ , \g155699/_0_ , \g155708/_0_ , \g155715/_0_ , \g156008/_0_ , \g156013/_0_ , \g156019/_0_ , \g156352/_0_ , \g156353/_0_ , \g156356/_0_ , \g156359/_0_ , \g156360/_0_ , \g156361/_0_ , \g156464/_0_ , \g156465/_0_ , \g156469/_0_ , \g156777/_0_ , \g156778/_0_ , \g156789/_0_ , \g158956/_0_ , \g158957/_0_ , \g158966/_0_ , \g159429/_1_ , \g159477/_1_ , \g159500/_1_ , \g159681/_0_ , \g159890/_0_ , \g159950/_0_ , \g160246/_0_ , \g160846/_0_ , \g160860/_0_ , \g160961/_0_ , \g160987/_0_ , \g161000/_0_ , \g161005/_0_ , \g161042/_0_ , \g161119/_0_ , \g161143/_0_ , \g161150/_0_ , \g161172/_0_ , \g161207/_0_ , \g161315/_0_ , \g161332/_0_ , \g161421/_0_ , \g161492/_0_ , \g161541/_0_ , \g161623/_0_ , \g161655/_0_ , \g161678/_0_ , \g161709/_0_ , \g161737/_0_ , \g161751/_0_ , \g161756/_0_ , \g162016/_0_ , \g162020/_0_ , \g162024/_0_ , \g163326/_0_ , \g163326/_3_ , \g174072/_1_ , \g174360/_1_ , \g174391/_0_ , \g180307/_0_ , \g180335/_0_ , \g180369/_0_ , \g180385/_0_ , \g180395/_0_ , \g180442/_0_ , \g180453/_0_ , \g180524/_0_ , \g180586/_0_ , \g180596/_0_ , \g180606/_0_ , \g180654/_0_ , \g180715/_0_ , \g180805/_0_ , \g180836/_0_ , \g180929/_0_ , \g180944/_0_ , \g180975/_0_ , \g181036/_0_ , \g181072/_0_ , \g181083/_0_ , \g181093/_0_ , \g181127/_0_ , \g181137/_0_ , \g181150/_0_ , \g181160/_0_ , \g181180/_0_ , \g181191/_0_ , \g181238/_0_ , \g181262/_0_ , \g181270/_0_ , \g181280/_0_ , \g181315/_0_ , \g181366/_0_ , \g181385/_0_ , \g181458/_0_ , \g181464/_0_ , \g181478/_0_ , \g181522/_0_ , \g181537/_0_ , \g181584/_0_ , \g181669/_0_ , \g181681/_0_ , \g181719/_0_ , \g181778/_0_ , \g181840/_0_ , \g181936/_0_ , \g181986/_0_ , \g182000/_0_ , \g182083/_0_ , \g182179/_0_ , \g182201/_0_ , \g182227/_0_ , \g182316/_0_ , \g182358/_0_ , \g182473/_0_ , \g182678/_0_ , \g53/_0_ );
	input \P1_BE_n_reg[0]/NET0131  ;
	input \P1_BE_n_reg[1]/NET0131  ;
	input \P1_BE_n_reg[2]/NET0131  ;
	input \P1_BE_n_reg[3]/NET0131  ;
	input \P1_ByteEnable_reg[0]/NET0131  ;
	input \P1_ByteEnable_reg[1]/NET0131  ;
	input \P1_ByteEnable_reg[2]/NET0131  ;
	input \P1_ByteEnable_reg[3]/NET0131  ;
	input \P1_CodeFetch_reg/NET0131  ;
	input \P1_D_C_n_reg/NET0131  ;
	input \P1_DataWidth_reg[0]/NET0131  ;
	input \P1_DataWidth_reg[1]/NET0131  ;
	input \P1_Datao_reg[0]/NET0131  ;
	input \P1_Datao_reg[10]/NET0131  ;
	input \P1_Datao_reg[11]/NET0131  ;
	input \P1_Datao_reg[12]/NET0131  ;
	input \P1_Datao_reg[13]/NET0131  ;
	input \P1_Datao_reg[14]/NET0131  ;
	input \P1_Datao_reg[15]/NET0131  ;
	input \P1_Datao_reg[16]/NET0131  ;
	input \P1_Datao_reg[17]/NET0131  ;
	input \P1_Datao_reg[18]/NET0131  ;
	input \P1_Datao_reg[19]/NET0131  ;
	input \P1_Datao_reg[1]/NET0131  ;
	input \P1_Datao_reg[20]/NET0131  ;
	input \P1_Datao_reg[21]/NET0131  ;
	input \P1_Datao_reg[22]/NET0131  ;
	input \P1_Datao_reg[23]/NET0131  ;
	input \P1_Datao_reg[24]/NET0131  ;
	input \P1_Datao_reg[25]/NET0131  ;
	input \P1_Datao_reg[26]/NET0131  ;
	input \P1_Datao_reg[27]/NET0131  ;
	input \P1_Datao_reg[28]/NET0131  ;
	input \P1_Datao_reg[29]/NET0131  ;
	input \P1_Datao_reg[2]/NET0131  ;
	input \P1_Datao_reg[30]/NET0131  ;
	input \P1_Datao_reg[3]/NET0131  ;
	input \P1_Datao_reg[4]/NET0131  ;
	input \P1_Datao_reg[5]/NET0131  ;
	input \P1_Datao_reg[6]/NET0131  ;
	input \P1_Datao_reg[7]/NET0131  ;
	input \P1_Datao_reg[8]/NET0131  ;
	input \P1_Datao_reg[9]/NET0131  ;
	input \P1_EAX_reg[0]/NET0131  ;
	input \P1_EAX_reg[10]/NET0131  ;
	input \P1_EAX_reg[11]/NET0131  ;
	input \P1_EAX_reg[12]/NET0131  ;
	input \P1_EAX_reg[13]/NET0131  ;
	input \P1_EAX_reg[14]/NET0131  ;
	input \P1_EAX_reg[15]/NET0131  ;
	input \P1_EAX_reg[16]/NET0131  ;
	input \P1_EAX_reg[17]/NET0131  ;
	input \P1_EAX_reg[18]/NET0131  ;
	input \P1_EAX_reg[19]/NET0131  ;
	input \P1_EAX_reg[1]/NET0131  ;
	input \P1_EAX_reg[20]/NET0131  ;
	input \P1_EAX_reg[21]/NET0131  ;
	input \P1_EAX_reg[22]/NET0131  ;
	input \P1_EAX_reg[23]/NET0131  ;
	input \P1_EAX_reg[24]/NET0131  ;
	input \P1_EAX_reg[25]/NET0131  ;
	input \P1_EAX_reg[26]/NET0131  ;
	input \P1_EAX_reg[27]/NET0131  ;
	input \P1_EAX_reg[28]/NET0131  ;
	input \P1_EAX_reg[29]/NET0131  ;
	input \P1_EAX_reg[2]/NET0131  ;
	input \P1_EAX_reg[30]/NET0131  ;
	input \P1_EAX_reg[31]/NET0131  ;
	input \P1_EAX_reg[3]/NET0131  ;
	input \P1_EAX_reg[4]/NET0131  ;
	input \P1_EAX_reg[5]/NET0131  ;
	input \P1_EAX_reg[6]/NET0131  ;
	input \P1_EAX_reg[7]/NET0131  ;
	input \P1_EAX_reg[8]/NET0131  ;
	input \P1_EAX_reg[9]/NET0131  ;
	input \P1_EBX_reg[0]/NET0131  ;
	input \P1_EBX_reg[10]/NET0131  ;
	input \P1_EBX_reg[11]/NET0131  ;
	input \P1_EBX_reg[12]/NET0131  ;
	input \P1_EBX_reg[13]/NET0131  ;
	input \P1_EBX_reg[14]/NET0131  ;
	input \P1_EBX_reg[15]/NET0131  ;
	input \P1_EBX_reg[16]/NET0131  ;
	input \P1_EBX_reg[17]/NET0131  ;
	input \P1_EBX_reg[18]/NET0131  ;
	input \P1_EBX_reg[19]/NET0131  ;
	input \P1_EBX_reg[1]/NET0131  ;
	input \P1_EBX_reg[20]/NET0131  ;
	input \P1_EBX_reg[21]/NET0131  ;
	input \P1_EBX_reg[22]/NET0131  ;
	input \P1_EBX_reg[23]/NET0131  ;
	input \P1_EBX_reg[24]/NET0131  ;
	input \P1_EBX_reg[25]/NET0131  ;
	input \P1_EBX_reg[26]/NET0131  ;
	input \P1_EBX_reg[27]/NET0131  ;
	input \P1_EBX_reg[28]/NET0131  ;
	input \P1_EBX_reg[29]/NET0131  ;
	input \P1_EBX_reg[2]/NET0131  ;
	input \P1_EBX_reg[30]/NET0131  ;
	input \P1_EBX_reg[31]/NET0131  ;
	input \P1_EBX_reg[3]/NET0131  ;
	input \P1_EBX_reg[4]/NET0131  ;
	input \P1_EBX_reg[5]/NET0131  ;
	input \P1_EBX_reg[6]/NET0131  ;
	input \P1_EBX_reg[7]/NET0131  ;
	input \P1_EBX_reg[8]/NET0131  ;
	input \P1_EBX_reg[9]/NET0131  ;
	input \P1_Flush_reg/NET0131  ;
	input \P1_InstAddrPointer_reg[0]/NET0131  ;
	input \P1_InstAddrPointer_reg[10]/NET0131  ;
	input \P1_InstAddrPointer_reg[11]/NET0131  ;
	input \P1_InstAddrPointer_reg[12]/NET0131  ;
	input \P1_InstAddrPointer_reg[13]/NET0131  ;
	input \P1_InstAddrPointer_reg[14]/NET0131  ;
	input \P1_InstAddrPointer_reg[15]/NET0131  ;
	input \P1_InstAddrPointer_reg[16]/NET0131  ;
	input \P1_InstAddrPointer_reg[17]/NET0131  ;
	input \P1_InstAddrPointer_reg[18]/NET0131  ;
	input \P1_InstAddrPointer_reg[19]/NET0131  ;
	input \P1_InstAddrPointer_reg[1]/NET0131  ;
	input \P1_InstAddrPointer_reg[20]/NET0131  ;
	input \P1_InstAddrPointer_reg[21]/NET0131  ;
	input \P1_InstAddrPointer_reg[22]/NET0131  ;
	input \P1_InstAddrPointer_reg[23]/NET0131  ;
	input \P1_InstAddrPointer_reg[24]/NET0131  ;
	input \P1_InstAddrPointer_reg[25]/NET0131  ;
	input \P1_InstAddrPointer_reg[26]/NET0131  ;
	input \P1_InstAddrPointer_reg[27]/NET0131  ;
	input \P1_InstAddrPointer_reg[28]/NET0131  ;
	input \P1_InstAddrPointer_reg[29]/NET0131  ;
	input \P1_InstAddrPointer_reg[2]/NET0131  ;
	input \P1_InstAddrPointer_reg[30]/NET0131  ;
	input \P1_InstAddrPointer_reg[31]/NET0131  ;
	input \P1_InstAddrPointer_reg[3]/NET0131  ;
	input \P1_InstAddrPointer_reg[4]/NET0131  ;
	input \P1_InstAddrPointer_reg[5]/NET0131  ;
	input \P1_InstAddrPointer_reg[6]/NET0131  ;
	input \P1_InstAddrPointer_reg[7]/NET0131  ;
	input \P1_InstAddrPointer_reg[8]/NET0131  ;
	input \P1_InstAddrPointer_reg[9]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P1_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P1_InstQueue_reg[0][0]/NET0131  ;
	input \P1_InstQueue_reg[0][1]/NET0131  ;
	input \P1_InstQueue_reg[0][2]/NET0131  ;
	input \P1_InstQueue_reg[0][3]/NET0131  ;
	input \P1_InstQueue_reg[0][4]/NET0131  ;
	input \P1_InstQueue_reg[0][5]/NET0131  ;
	input \P1_InstQueue_reg[0][6]/NET0131  ;
	input \P1_InstQueue_reg[0][7]/NET0131  ;
	input \P1_InstQueue_reg[10][0]/NET0131  ;
	input \P1_InstQueue_reg[10][1]/NET0131  ;
	input \P1_InstQueue_reg[10][2]/NET0131  ;
	input \P1_InstQueue_reg[10][3]/NET0131  ;
	input \P1_InstQueue_reg[10][4]/NET0131  ;
	input \P1_InstQueue_reg[10][5]/NET0131  ;
	input \P1_InstQueue_reg[10][6]/NET0131  ;
	input \P1_InstQueue_reg[10][7]/NET0131  ;
	input \P1_InstQueue_reg[11][0]/NET0131  ;
	input \P1_InstQueue_reg[11][1]/NET0131  ;
	input \P1_InstQueue_reg[11][2]/NET0131  ;
	input \P1_InstQueue_reg[11][3]/NET0131  ;
	input \P1_InstQueue_reg[11][4]/NET0131  ;
	input \P1_InstQueue_reg[11][5]/NET0131  ;
	input \P1_InstQueue_reg[11][6]/NET0131  ;
	input \P1_InstQueue_reg[11][7]/NET0131  ;
	input \P1_InstQueue_reg[12][0]/NET0131  ;
	input \P1_InstQueue_reg[12][1]/NET0131  ;
	input \P1_InstQueue_reg[12][2]/NET0131  ;
	input \P1_InstQueue_reg[12][3]/NET0131  ;
	input \P1_InstQueue_reg[12][4]/NET0131  ;
	input \P1_InstQueue_reg[12][5]/NET0131  ;
	input \P1_InstQueue_reg[12][6]/NET0131  ;
	input \P1_InstQueue_reg[12][7]/NET0131  ;
	input \P1_InstQueue_reg[13][0]/NET0131  ;
	input \P1_InstQueue_reg[13][1]/NET0131  ;
	input \P1_InstQueue_reg[13][2]/NET0131  ;
	input \P1_InstQueue_reg[13][3]/NET0131  ;
	input \P1_InstQueue_reg[13][4]/NET0131  ;
	input \P1_InstQueue_reg[13][5]/NET0131  ;
	input \P1_InstQueue_reg[13][6]/NET0131  ;
	input \P1_InstQueue_reg[13][7]/NET0131  ;
	input \P1_InstQueue_reg[14][0]/NET0131  ;
	input \P1_InstQueue_reg[14][1]/NET0131  ;
	input \P1_InstQueue_reg[14][2]/NET0131  ;
	input \P1_InstQueue_reg[14][3]/NET0131  ;
	input \P1_InstQueue_reg[14][4]/NET0131  ;
	input \P1_InstQueue_reg[14][5]/NET0131  ;
	input \P1_InstQueue_reg[14][6]/NET0131  ;
	input \P1_InstQueue_reg[14][7]/NET0131  ;
	input \P1_InstQueue_reg[15][0]/NET0131  ;
	input \P1_InstQueue_reg[15][1]/NET0131  ;
	input \P1_InstQueue_reg[15][2]/NET0131  ;
	input \P1_InstQueue_reg[15][3]/NET0131  ;
	input \P1_InstQueue_reg[15][4]/NET0131  ;
	input \P1_InstQueue_reg[15][5]/NET0131  ;
	input \P1_InstQueue_reg[15][6]/NET0131  ;
	input \P1_InstQueue_reg[15][7]/NET0131  ;
	input \P1_InstQueue_reg[1][0]/NET0131  ;
	input \P1_InstQueue_reg[1][1]/NET0131  ;
	input \P1_InstQueue_reg[1][2]/NET0131  ;
	input \P1_InstQueue_reg[1][3]/NET0131  ;
	input \P1_InstQueue_reg[1][4]/NET0131  ;
	input \P1_InstQueue_reg[1][5]/NET0131  ;
	input \P1_InstQueue_reg[1][6]/NET0131  ;
	input \P1_InstQueue_reg[1][7]/NET0131  ;
	input \P1_InstQueue_reg[2][0]/NET0131  ;
	input \P1_InstQueue_reg[2][1]/NET0131  ;
	input \P1_InstQueue_reg[2][2]/NET0131  ;
	input \P1_InstQueue_reg[2][3]/NET0131  ;
	input \P1_InstQueue_reg[2][4]/NET0131  ;
	input \P1_InstQueue_reg[2][5]/NET0131  ;
	input \P1_InstQueue_reg[2][6]/NET0131  ;
	input \P1_InstQueue_reg[2][7]/NET0131  ;
	input \P1_InstQueue_reg[3][0]/NET0131  ;
	input \P1_InstQueue_reg[3][1]/NET0131  ;
	input \P1_InstQueue_reg[3][2]/NET0131  ;
	input \P1_InstQueue_reg[3][3]/NET0131  ;
	input \P1_InstQueue_reg[3][4]/NET0131  ;
	input \P1_InstQueue_reg[3][5]/NET0131  ;
	input \P1_InstQueue_reg[3][6]/NET0131  ;
	input \P1_InstQueue_reg[3][7]/NET0131  ;
	input \P1_InstQueue_reg[4][0]/NET0131  ;
	input \P1_InstQueue_reg[4][1]/NET0131  ;
	input \P1_InstQueue_reg[4][2]/NET0131  ;
	input \P1_InstQueue_reg[4][3]/NET0131  ;
	input \P1_InstQueue_reg[4][4]/NET0131  ;
	input \P1_InstQueue_reg[4][5]/NET0131  ;
	input \P1_InstQueue_reg[4][6]/NET0131  ;
	input \P1_InstQueue_reg[4][7]/NET0131  ;
	input \P1_InstQueue_reg[5][0]/NET0131  ;
	input \P1_InstQueue_reg[5][1]/NET0131  ;
	input \P1_InstQueue_reg[5][2]/NET0131  ;
	input \P1_InstQueue_reg[5][3]/NET0131  ;
	input \P1_InstQueue_reg[5][4]/NET0131  ;
	input \P1_InstQueue_reg[5][5]/NET0131  ;
	input \P1_InstQueue_reg[5][6]/NET0131  ;
	input \P1_InstQueue_reg[5][7]/NET0131  ;
	input \P1_InstQueue_reg[6][0]/NET0131  ;
	input \P1_InstQueue_reg[6][1]/NET0131  ;
	input \P1_InstQueue_reg[6][2]/NET0131  ;
	input \P1_InstQueue_reg[6][3]/NET0131  ;
	input \P1_InstQueue_reg[6][4]/NET0131  ;
	input \P1_InstQueue_reg[6][5]/NET0131  ;
	input \P1_InstQueue_reg[6][6]/NET0131  ;
	input \P1_InstQueue_reg[6][7]/NET0131  ;
	input \P1_InstQueue_reg[7][0]/NET0131  ;
	input \P1_InstQueue_reg[7][1]/NET0131  ;
	input \P1_InstQueue_reg[7][2]/NET0131  ;
	input \P1_InstQueue_reg[7][3]/NET0131  ;
	input \P1_InstQueue_reg[7][4]/NET0131  ;
	input \P1_InstQueue_reg[7][5]/NET0131  ;
	input \P1_InstQueue_reg[7][6]/NET0131  ;
	input \P1_InstQueue_reg[7][7]/NET0131  ;
	input \P1_InstQueue_reg[8][0]/NET0131  ;
	input \P1_InstQueue_reg[8][1]/NET0131  ;
	input \P1_InstQueue_reg[8][2]/NET0131  ;
	input \P1_InstQueue_reg[8][3]/NET0131  ;
	input \P1_InstQueue_reg[8][4]/NET0131  ;
	input \P1_InstQueue_reg[8][5]/NET0131  ;
	input \P1_InstQueue_reg[8][6]/NET0131  ;
	input \P1_InstQueue_reg[8][7]/NET0131  ;
	input \P1_InstQueue_reg[9][0]/NET0131  ;
	input \P1_InstQueue_reg[9][1]/NET0131  ;
	input \P1_InstQueue_reg[9][2]/NET0131  ;
	input \P1_InstQueue_reg[9][3]/NET0131  ;
	input \P1_InstQueue_reg[9][4]/NET0131  ;
	input \P1_InstQueue_reg[9][5]/NET0131  ;
	input \P1_InstQueue_reg[9][6]/NET0131  ;
	input \P1_InstQueue_reg[9][7]/NET0131  ;
	input \P1_M_IO_n_reg/NET0131  ;
	input \P1_MemoryFetch_reg/NET0131  ;
	input \P1_More_reg/NET0131  ;
	input \P1_PhyAddrPointer_reg[0]/NET0131  ;
	input \P1_PhyAddrPointer_reg[10]/NET0131  ;
	input \P1_PhyAddrPointer_reg[11]/NET0131  ;
	input \P1_PhyAddrPointer_reg[12]/NET0131  ;
	input \P1_PhyAddrPointer_reg[13]/NET0131  ;
	input \P1_PhyAddrPointer_reg[14]/NET0131  ;
	input \P1_PhyAddrPointer_reg[15]/NET0131  ;
	input \P1_PhyAddrPointer_reg[16]/NET0131  ;
	input \P1_PhyAddrPointer_reg[17]/NET0131  ;
	input \P1_PhyAddrPointer_reg[18]/NET0131  ;
	input \P1_PhyAddrPointer_reg[19]/NET0131  ;
	input \P1_PhyAddrPointer_reg[1]/NET0131  ;
	input \P1_PhyAddrPointer_reg[20]/NET0131  ;
	input \P1_PhyAddrPointer_reg[21]/NET0131  ;
	input \P1_PhyAddrPointer_reg[22]/NET0131  ;
	input \P1_PhyAddrPointer_reg[23]/NET0131  ;
	input \P1_PhyAddrPointer_reg[24]/NET0131  ;
	input \P1_PhyAddrPointer_reg[25]/NET0131  ;
	input \P1_PhyAddrPointer_reg[26]/NET0131  ;
	input \P1_PhyAddrPointer_reg[27]/NET0131  ;
	input \P1_PhyAddrPointer_reg[28]/NET0131  ;
	input \P1_PhyAddrPointer_reg[29]/NET0131  ;
	input \P1_PhyAddrPointer_reg[2]/NET0131  ;
	input \P1_PhyAddrPointer_reg[30]/NET0131  ;
	input \P1_PhyAddrPointer_reg[31]/NET0131  ;
	input \P1_PhyAddrPointer_reg[3]/NET0131  ;
	input \P1_PhyAddrPointer_reg[4]/NET0131  ;
	input \P1_PhyAddrPointer_reg[5]/NET0131  ;
	input \P1_PhyAddrPointer_reg[6]/NET0131  ;
	input \P1_PhyAddrPointer_reg[7]/NET0131  ;
	input \P1_PhyAddrPointer_reg[8]/NET0131  ;
	input \P1_PhyAddrPointer_reg[9]/NET0131  ;
	input \P1_ReadRequest_reg/NET0131  ;
	input \P1_RequestPending_reg/NET0131  ;
	input \P1_State2_reg[0]/NET0131  ;
	input \P1_State2_reg[1]/NET0131  ;
	input \P1_State2_reg[2]/NET0131  ;
	input \P1_State2_reg[3]/NET0131  ;
	input \P1_State_reg[0]/NET0131  ;
	input \P1_State_reg[1]/NET0131  ;
	input \P1_State_reg[2]/NET0131  ;
	input \P1_W_R_n_reg/NET0131  ;
	input \P1_lWord_reg[0]/NET0131  ;
	input \P1_lWord_reg[10]/NET0131  ;
	input \P1_lWord_reg[11]/NET0131  ;
	input \P1_lWord_reg[12]/NET0131  ;
	input \P1_lWord_reg[13]/NET0131  ;
	input \P1_lWord_reg[14]/NET0131  ;
	input \P1_lWord_reg[15]/NET0131  ;
	input \P1_lWord_reg[1]/NET0131  ;
	input \P1_lWord_reg[2]/NET0131  ;
	input \P1_lWord_reg[3]/NET0131  ;
	input \P1_lWord_reg[4]/NET0131  ;
	input \P1_lWord_reg[5]/NET0131  ;
	input \P1_lWord_reg[6]/NET0131  ;
	input \P1_lWord_reg[7]/NET0131  ;
	input \P1_lWord_reg[8]/NET0131  ;
	input \P1_lWord_reg[9]/NET0131  ;
	input \P1_rEIP_reg[0]/NET0131  ;
	input \P1_rEIP_reg[10]/NET0131  ;
	input \P1_rEIP_reg[11]/NET0131  ;
	input \P1_rEIP_reg[12]/NET0131  ;
	input \P1_rEIP_reg[13]/NET0131  ;
	input \P1_rEIP_reg[14]/NET0131  ;
	input \P1_rEIP_reg[15]/NET0131  ;
	input \P1_rEIP_reg[16]/NET0131  ;
	input \P1_rEIP_reg[17]/NET0131  ;
	input \P1_rEIP_reg[18]/NET0131  ;
	input \P1_rEIP_reg[19]/NET0131  ;
	input \P1_rEIP_reg[1]/NET0131  ;
	input \P1_rEIP_reg[20]/NET0131  ;
	input \P1_rEIP_reg[21]/NET0131  ;
	input \P1_rEIP_reg[22]/NET0131  ;
	input \P1_rEIP_reg[23]/NET0131  ;
	input \P1_rEIP_reg[24]/NET0131  ;
	input \P1_rEIP_reg[25]/NET0131  ;
	input \P1_rEIP_reg[26]/NET0131  ;
	input \P1_rEIP_reg[27]/NET0131  ;
	input \P1_rEIP_reg[28]/NET0131  ;
	input \P1_rEIP_reg[29]/NET0131  ;
	input \P1_rEIP_reg[2]/NET0131  ;
	input \P1_rEIP_reg[30]/NET0131  ;
	input \P1_rEIP_reg[31]/NET0131  ;
	input \P1_rEIP_reg[3]/NET0131  ;
	input \P1_rEIP_reg[4]/NET0131  ;
	input \P1_rEIP_reg[5]/NET0131  ;
	input \P1_rEIP_reg[6]/NET0131  ;
	input \P1_rEIP_reg[7]/NET0131  ;
	input \P1_rEIP_reg[8]/NET0131  ;
	input \P1_rEIP_reg[9]/NET0131  ;
	input \P1_uWord_reg[0]/NET0131  ;
	input \P1_uWord_reg[10]/NET0131  ;
	input \P1_uWord_reg[11]/NET0131  ;
	input \P1_uWord_reg[12]/NET0131  ;
	input \P1_uWord_reg[13]/NET0131  ;
	input \P1_uWord_reg[14]/NET0131  ;
	input \P1_uWord_reg[1]/NET0131  ;
	input \P1_uWord_reg[2]/NET0131  ;
	input \P1_uWord_reg[3]/NET0131  ;
	input \P1_uWord_reg[4]/NET0131  ;
	input \P1_uWord_reg[5]/NET0131  ;
	input \P1_uWord_reg[6]/NET0131  ;
	input \P1_uWord_reg[7]/NET0131  ;
	input \P1_uWord_reg[8]/NET0131  ;
	input \P1_uWord_reg[9]/NET0131  ;
	input \P2_ADS_n_reg/NET0131  ;
	input \P2_Address_reg[0]/NET0131  ;
	input \P2_Address_reg[10]/NET0131  ;
	input \P2_Address_reg[11]/NET0131  ;
	input \P2_Address_reg[12]/NET0131  ;
	input \P2_Address_reg[13]/NET0131  ;
	input \P2_Address_reg[14]/NET0131  ;
	input \P2_Address_reg[15]/NET0131  ;
	input \P2_Address_reg[16]/NET0131  ;
	input \P2_Address_reg[17]/NET0131  ;
	input \P2_Address_reg[18]/NET0131  ;
	input \P2_Address_reg[19]/NET0131  ;
	input \P2_Address_reg[1]/NET0131  ;
	input \P2_Address_reg[20]/NET0131  ;
	input \P2_Address_reg[21]/NET0131  ;
	input \P2_Address_reg[22]/NET0131  ;
	input \P2_Address_reg[23]/NET0131  ;
	input \P2_Address_reg[24]/NET0131  ;
	input \P2_Address_reg[25]/NET0131  ;
	input \P2_Address_reg[26]/NET0131  ;
	input \P2_Address_reg[27]/NET0131  ;
	input \P2_Address_reg[28]/NET0131  ;
	input \P2_Address_reg[29]/NET0131  ;
	input \P2_Address_reg[2]/NET0131  ;
	input \P2_Address_reg[3]/NET0131  ;
	input \P2_Address_reg[4]/NET0131  ;
	input \P2_Address_reg[5]/NET0131  ;
	input \P2_Address_reg[6]/NET0131  ;
	input \P2_Address_reg[7]/NET0131  ;
	input \P2_Address_reg[8]/NET0131  ;
	input \P2_Address_reg[9]/NET0131  ;
	input \P2_BE_n_reg[0]/NET0131  ;
	input \P2_BE_n_reg[1]/NET0131  ;
	input \P2_BE_n_reg[2]/NET0131  ;
	input \P2_BE_n_reg[3]/NET0131  ;
	input \P2_ByteEnable_reg[0]/NET0131  ;
	input \P2_ByteEnable_reg[1]/NET0131  ;
	input \P2_ByteEnable_reg[2]/NET0131  ;
	input \P2_ByteEnable_reg[3]/NET0131  ;
	input \P2_CodeFetch_reg/NET0131  ;
	input \P2_D_C_n_reg/NET0131  ;
	input \P2_DataWidth_reg[0]/NET0131  ;
	input \P2_DataWidth_reg[1]/NET0131  ;
	input \P2_Datao_reg[0]/NET0131  ;
	input \P2_Datao_reg[10]/NET0131  ;
	input \P2_Datao_reg[11]/NET0131  ;
	input \P2_Datao_reg[12]/NET0131  ;
	input \P2_Datao_reg[13]/NET0131  ;
	input \P2_Datao_reg[14]/NET0131  ;
	input \P2_Datao_reg[15]/NET0131  ;
	input \P2_Datao_reg[16]/NET0131  ;
	input \P2_Datao_reg[17]/NET0131  ;
	input \P2_Datao_reg[18]/NET0131  ;
	input \P2_Datao_reg[19]/NET0131  ;
	input \P2_Datao_reg[1]/NET0131  ;
	input \P2_Datao_reg[20]/NET0131  ;
	input \P2_Datao_reg[21]/NET0131  ;
	input \P2_Datao_reg[22]/NET0131  ;
	input \P2_Datao_reg[23]/NET0131  ;
	input \P2_Datao_reg[24]/NET0131  ;
	input \P2_Datao_reg[25]/NET0131  ;
	input \P2_Datao_reg[26]/NET0131  ;
	input \P2_Datao_reg[27]/NET0131  ;
	input \P2_Datao_reg[28]/NET0131  ;
	input \P2_Datao_reg[29]/NET0131  ;
	input \P2_Datao_reg[2]/NET0131  ;
	input \P2_Datao_reg[30]/NET0131  ;
	input \P2_Datao_reg[3]/NET0131  ;
	input \P2_Datao_reg[4]/NET0131  ;
	input \P2_Datao_reg[5]/NET0131  ;
	input \P2_Datao_reg[6]/NET0131  ;
	input \P2_Datao_reg[7]/NET0131  ;
	input \P2_Datao_reg[8]/NET0131  ;
	input \P2_Datao_reg[9]/NET0131  ;
	input \P2_EAX_reg[0]/NET0131  ;
	input \P2_EAX_reg[10]/NET0131  ;
	input \P2_EAX_reg[11]/NET0131  ;
	input \P2_EAX_reg[12]/NET0131  ;
	input \P2_EAX_reg[13]/NET0131  ;
	input \P2_EAX_reg[14]/NET0131  ;
	input \P2_EAX_reg[15]/NET0131  ;
	input \P2_EAX_reg[16]/NET0131  ;
	input \P2_EAX_reg[17]/NET0131  ;
	input \P2_EAX_reg[18]/NET0131  ;
	input \P2_EAX_reg[19]/NET0131  ;
	input \P2_EAX_reg[1]/NET0131  ;
	input \P2_EAX_reg[20]/NET0131  ;
	input \P2_EAX_reg[21]/NET0131  ;
	input \P2_EAX_reg[22]/NET0131  ;
	input \P2_EAX_reg[23]/NET0131  ;
	input \P2_EAX_reg[24]/NET0131  ;
	input \P2_EAX_reg[25]/NET0131  ;
	input \P2_EAX_reg[26]/NET0131  ;
	input \P2_EAX_reg[27]/NET0131  ;
	input \P2_EAX_reg[28]/NET0131  ;
	input \P2_EAX_reg[29]/NET0131  ;
	input \P2_EAX_reg[2]/NET0131  ;
	input \P2_EAX_reg[30]/NET0131  ;
	input \P2_EAX_reg[31]/NET0131  ;
	input \P2_EAX_reg[3]/NET0131  ;
	input \P2_EAX_reg[4]/NET0131  ;
	input \P2_EAX_reg[5]/NET0131  ;
	input \P2_EAX_reg[6]/NET0131  ;
	input \P2_EAX_reg[7]/NET0131  ;
	input \P2_EAX_reg[8]/NET0131  ;
	input \P2_EAX_reg[9]/NET0131  ;
	input \P2_EBX_reg[0]/NET0131  ;
	input \P2_EBX_reg[10]/NET0131  ;
	input \P2_EBX_reg[11]/NET0131  ;
	input \P2_EBX_reg[12]/NET0131  ;
	input \P2_EBX_reg[13]/NET0131  ;
	input \P2_EBX_reg[14]/NET0131  ;
	input \P2_EBX_reg[15]/NET0131  ;
	input \P2_EBX_reg[16]/NET0131  ;
	input \P2_EBX_reg[17]/NET0131  ;
	input \P2_EBX_reg[18]/NET0131  ;
	input \P2_EBX_reg[19]/NET0131  ;
	input \P2_EBX_reg[1]/NET0131  ;
	input \P2_EBX_reg[20]/NET0131  ;
	input \P2_EBX_reg[21]/NET0131  ;
	input \P2_EBX_reg[22]/NET0131  ;
	input \P2_EBX_reg[23]/NET0131  ;
	input \P2_EBX_reg[24]/NET0131  ;
	input \P2_EBX_reg[25]/NET0131  ;
	input \P2_EBX_reg[26]/NET0131  ;
	input \P2_EBX_reg[27]/NET0131  ;
	input \P2_EBX_reg[28]/NET0131  ;
	input \P2_EBX_reg[29]/NET0131  ;
	input \P2_EBX_reg[2]/NET0131  ;
	input \P2_EBX_reg[30]/NET0131  ;
	input \P2_EBX_reg[31]/NET0131  ;
	input \P2_EBX_reg[3]/NET0131  ;
	input \P2_EBX_reg[4]/NET0131  ;
	input \P2_EBX_reg[5]/NET0131  ;
	input \P2_EBX_reg[6]/NET0131  ;
	input \P2_EBX_reg[7]/NET0131  ;
	input \P2_EBX_reg[8]/NET0131  ;
	input \P2_EBX_reg[9]/NET0131  ;
	input \P2_Flush_reg/NET0131  ;
	input \P2_InstAddrPointer_reg[0]/NET0131  ;
	input \P2_InstAddrPointer_reg[10]/NET0131  ;
	input \P2_InstAddrPointer_reg[11]/NET0131  ;
	input \P2_InstAddrPointer_reg[12]/NET0131  ;
	input \P2_InstAddrPointer_reg[13]/NET0131  ;
	input \P2_InstAddrPointer_reg[14]/NET0131  ;
	input \P2_InstAddrPointer_reg[15]/NET0131  ;
	input \P2_InstAddrPointer_reg[16]/NET0131  ;
	input \P2_InstAddrPointer_reg[17]/NET0131  ;
	input \P2_InstAddrPointer_reg[18]/NET0131  ;
	input \P2_InstAddrPointer_reg[19]/NET0131  ;
	input \P2_InstAddrPointer_reg[1]/NET0131  ;
	input \P2_InstAddrPointer_reg[20]/NET0131  ;
	input \P2_InstAddrPointer_reg[21]/NET0131  ;
	input \P2_InstAddrPointer_reg[22]/NET0131  ;
	input \P2_InstAddrPointer_reg[23]/NET0131  ;
	input \P2_InstAddrPointer_reg[24]/NET0131  ;
	input \P2_InstAddrPointer_reg[25]/NET0131  ;
	input \P2_InstAddrPointer_reg[26]/NET0131  ;
	input \P2_InstAddrPointer_reg[27]/NET0131  ;
	input \P2_InstAddrPointer_reg[28]/NET0131  ;
	input \P2_InstAddrPointer_reg[29]/NET0131  ;
	input \P2_InstAddrPointer_reg[2]/NET0131  ;
	input \P2_InstAddrPointer_reg[30]/NET0131  ;
	input \P2_InstAddrPointer_reg[31]/NET0131  ;
	input \P2_InstAddrPointer_reg[3]/NET0131  ;
	input \P2_InstAddrPointer_reg[4]/NET0131  ;
	input \P2_InstAddrPointer_reg[5]/NET0131  ;
	input \P2_InstAddrPointer_reg[6]/NET0131  ;
	input \P2_InstAddrPointer_reg[7]/NET0131  ;
	input \P2_InstAddrPointer_reg[8]/NET0131  ;
	input \P2_InstAddrPointer_reg[9]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P2_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P2_InstQueue_reg[0][0]/NET0131  ;
	input \P2_InstQueue_reg[0][1]/NET0131  ;
	input \P2_InstQueue_reg[0][2]/NET0131  ;
	input \P2_InstQueue_reg[0][3]/NET0131  ;
	input \P2_InstQueue_reg[0][4]/NET0131  ;
	input \P2_InstQueue_reg[0][5]/NET0131  ;
	input \P2_InstQueue_reg[0][6]/NET0131  ;
	input \P2_InstQueue_reg[0][7]/NET0131  ;
	input \P2_InstQueue_reg[10][0]/NET0131  ;
	input \P2_InstQueue_reg[10][1]/NET0131  ;
	input \P2_InstQueue_reg[10][2]/NET0131  ;
	input \P2_InstQueue_reg[10][3]/NET0131  ;
	input \P2_InstQueue_reg[10][4]/NET0131  ;
	input \P2_InstQueue_reg[10][5]/NET0131  ;
	input \P2_InstQueue_reg[10][6]/NET0131  ;
	input \P2_InstQueue_reg[10][7]/NET0131  ;
	input \P2_InstQueue_reg[11][0]/NET0131  ;
	input \P2_InstQueue_reg[11][1]/NET0131  ;
	input \P2_InstQueue_reg[11][2]/NET0131  ;
	input \P2_InstQueue_reg[11][3]/NET0131  ;
	input \P2_InstQueue_reg[11][4]/NET0131  ;
	input \P2_InstQueue_reg[11][5]/NET0131  ;
	input \P2_InstQueue_reg[11][6]/NET0131  ;
	input \P2_InstQueue_reg[11][7]/NET0131  ;
	input \P2_InstQueue_reg[12][0]/NET0131  ;
	input \P2_InstQueue_reg[12][1]/NET0131  ;
	input \P2_InstQueue_reg[12][2]/NET0131  ;
	input \P2_InstQueue_reg[12][3]/NET0131  ;
	input \P2_InstQueue_reg[12][4]/NET0131  ;
	input \P2_InstQueue_reg[12][5]/NET0131  ;
	input \P2_InstQueue_reg[12][6]/NET0131  ;
	input \P2_InstQueue_reg[12][7]/NET0131  ;
	input \P2_InstQueue_reg[13][0]/NET0131  ;
	input \P2_InstQueue_reg[13][1]/NET0131  ;
	input \P2_InstQueue_reg[13][2]/NET0131  ;
	input \P2_InstQueue_reg[13][3]/NET0131  ;
	input \P2_InstQueue_reg[13][4]/NET0131  ;
	input \P2_InstQueue_reg[13][5]/NET0131  ;
	input \P2_InstQueue_reg[13][6]/NET0131  ;
	input \P2_InstQueue_reg[13][7]/NET0131  ;
	input \P2_InstQueue_reg[14][0]/NET0131  ;
	input \P2_InstQueue_reg[14][1]/NET0131  ;
	input \P2_InstQueue_reg[14][2]/NET0131  ;
	input \P2_InstQueue_reg[14][3]/NET0131  ;
	input \P2_InstQueue_reg[14][4]/NET0131  ;
	input \P2_InstQueue_reg[14][5]/NET0131  ;
	input \P2_InstQueue_reg[14][6]/NET0131  ;
	input \P2_InstQueue_reg[14][7]/NET0131  ;
	input \P2_InstQueue_reg[15][0]/NET0131  ;
	input \P2_InstQueue_reg[15][1]/NET0131  ;
	input \P2_InstQueue_reg[15][2]/NET0131  ;
	input \P2_InstQueue_reg[15][3]/NET0131  ;
	input \P2_InstQueue_reg[15][4]/NET0131  ;
	input \P2_InstQueue_reg[15][5]/NET0131  ;
	input \P2_InstQueue_reg[15][6]/NET0131  ;
	input \P2_InstQueue_reg[15][7]/NET0131  ;
	input \P2_InstQueue_reg[1][0]/NET0131  ;
	input \P2_InstQueue_reg[1][1]/NET0131  ;
	input \P2_InstQueue_reg[1][2]/NET0131  ;
	input \P2_InstQueue_reg[1][3]/NET0131  ;
	input \P2_InstQueue_reg[1][4]/NET0131  ;
	input \P2_InstQueue_reg[1][5]/NET0131  ;
	input \P2_InstQueue_reg[1][6]/NET0131  ;
	input \P2_InstQueue_reg[1][7]/NET0131  ;
	input \P2_InstQueue_reg[2][0]/NET0131  ;
	input \P2_InstQueue_reg[2][1]/NET0131  ;
	input \P2_InstQueue_reg[2][2]/NET0131  ;
	input \P2_InstQueue_reg[2][3]/NET0131  ;
	input \P2_InstQueue_reg[2][4]/NET0131  ;
	input \P2_InstQueue_reg[2][5]/NET0131  ;
	input \P2_InstQueue_reg[2][6]/NET0131  ;
	input \P2_InstQueue_reg[2][7]/NET0131  ;
	input \P2_InstQueue_reg[3][0]/NET0131  ;
	input \P2_InstQueue_reg[3][1]/NET0131  ;
	input \P2_InstQueue_reg[3][2]/NET0131  ;
	input \P2_InstQueue_reg[3][3]/NET0131  ;
	input \P2_InstQueue_reg[3][4]/NET0131  ;
	input \P2_InstQueue_reg[3][5]/NET0131  ;
	input \P2_InstQueue_reg[3][6]/NET0131  ;
	input \P2_InstQueue_reg[3][7]/NET0131  ;
	input \P2_InstQueue_reg[4][0]/NET0131  ;
	input \P2_InstQueue_reg[4][1]/NET0131  ;
	input \P2_InstQueue_reg[4][2]/NET0131  ;
	input \P2_InstQueue_reg[4][3]/NET0131  ;
	input \P2_InstQueue_reg[4][4]/NET0131  ;
	input \P2_InstQueue_reg[4][5]/NET0131  ;
	input \P2_InstQueue_reg[4][6]/NET0131  ;
	input \P2_InstQueue_reg[4][7]/NET0131  ;
	input \P2_InstQueue_reg[5][0]/NET0131  ;
	input \P2_InstQueue_reg[5][1]/NET0131  ;
	input \P2_InstQueue_reg[5][2]/NET0131  ;
	input \P2_InstQueue_reg[5][3]/NET0131  ;
	input \P2_InstQueue_reg[5][4]/NET0131  ;
	input \P2_InstQueue_reg[5][5]/NET0131  ;
	input \P2_InstQueue_reg[5][6]/NET0131  ;
	input \P2_InstQueue_reg[5][7]/NET0131  ;
	input \P2_InstQueue_reg[6][0]/NET0131  ;
	input \P2_InstQueue_reg[6][1]/NET0131  ;
	input \P2_InstQueue_reg[6][2]/NET0131  ;
	input \P2_InstQueue_reg[6][3]/NET0131  ;
	input \P2_InstQueue_reg[6][4]/NET0131  ;
	input \P2_InstQueue_reg[6][5]/NET0131  ;
	input \P2_InstQueue_reg[6][6]/NET0131  ;
	input \P2_InstQueue_reg[6][7]/NET0131  ;
	input \P2_InstQueue_reg[7][0]/NET0131  ;
	input \P2_InstQueue_reg[7][1]/NET0131  ;
	input \P2_InstQueue_reg[7][2]/NET0131  ;
	input \P2_InstQueue_reg[7][3]/NET0131  ;
	input \P2_InstQueue_reg[7][4]/NET0131  ;
	input \P2_InstQueue_reg[7][5]/NET0131  ;
	input \P2_InstQueue_reg[7][6]/NET0131  ;
	input \P2_InstQueue_reg[7][7]/NET0131  ;
	input \P2_InstQueue_reg[8][0]/NET0131  ;
	input \P2_InstQueue_reg[8][1]/NET0131  ;
	input \P2_InstQueue_reg[8][2]/NET0131  ;
	input \P2_InstQueue_reg[8][3]/NET0131  ;
	input \P2_InstQueue_reg[8][4]/NET0131  ;
	input \P2_InstQueue_reg[8][5]/NET0131  ;
	input \P2_InstQueue_reg[8][6]/NET0131  ;
	input \P2_InstQueue_reg[8][7]/NET0131  ;
	input \P2_InstQueue_reg[9][0]/NET0131  ;
	input \P2_InstQueue_reg[9][1]/NET0131  ;
	input \P2_InstQueue_reg[9][2]/NET0131  ;
	input \P2_InstQueue_reg[9][3]/NET0131  ;
	input \P2_InstQueue_reg[9][4]/NET0131  ;
	input \P2_InstQueue_reg[9][5]/NET0131  ;
	input \P2_InstQueue_reg[9][6]/NET0131  ;
	input \P2_InstQueue_reg[9][7]/NET0131  ;
	input \P2_M_IO_n_reg/NET0131  ;
	input \P2_MemoryFetch_reg/NET0131  ;
	input \P2_More_reg/NET0131  ;
	input \P2_PhyAddrPointer_reg[0]/NET0131  ;
	input \P2_PhyAddrPointer_reg[10]/NET0131  ;
	input \P2_PhyAddrPointer_reg[11]/NET0131  ;
	input \P2_PhyAddrPointer_reg[12]/NET0131  ;
	input \P2_PhyAddrPointer_reg[13]/NET0131  ;
	input \P2_PhyAddrPointer_reg[14]/NET0131  ;
	input \P2_PhyAddrPointer_reg[15]/NET0131  ;
	input \P2_PhyAddrPointer_reg[16]/NET0131  ;
	input \P2_PhyAddrPointer_reg[17]/NET0131  ;
	input \P2_PhyAddrPointer_reg[18]/NET0131  ;
	input \P2_PhyAddrPointer_reg[19]/NET0131  ;
	input \P2_PhyAddrPointer_reg[1]/NET0131  ;
	input \P2_PhyAddrPointer_reg[20]/NET0131  ;
	input \P2_PhyAddrPointer_reg[21]/NET0131  ;
	input \P2_PhyAddrPointer_reg[22]/NET0131  ;
	input \P2_PhyAddrPointer_reg[23]/NET0131  ;
	input \P2_PhyAddrPointer_reg[24]/NET0131  ;
	input \P2_PhyAddrPointer_reg[25]/NET0131  ;
	input \P2_PhyAddrPointer_reg[26]/NET0131  ;
	input \P2_PhyAddrPointer_reg[27]/NET0131  ;
	input \P2_PhyAddrPointer_reg[28]/NET0131  ;
	input \P2_PhyAddrPointer_reg[29]/NET0131  ;
	input \P2_PhyAddrPointer_reg[2]/NET0131  ;
	input \P2_PhyAddrPointer_reg[30]/NET0131  ;
	input \P2_PhyAddrPointer_reg[31]/NET0131  ;
	input \P2_PhyAddrPointer_reg[3]/NET0131  ;
	input \P2_PhyAddrPointer_reg[4]/NET0131  ;
	input \P2_PhyAddrPointer_reg[5]/NET0131  ;
	input \P2_PhyAddrPointer_reg[6]/NET0131  ;
	input \P2_PhyAddrPointer_reg[7]/NET0131  ;
	input \P2_PhyAddrPointer_reg[8]/NET0131  ;
	input \P2_PhyAddrPointer_reg[9]/NET0131  ;
	input \P2_ReadRequest_reg/NET0131  ;
	input \P2_RequestPending_reg/NET0131  ;
	input \P2_State2_reg[0]/NET0131  ;
	input \P2_State2_reg[1]/NET0131  ;
	input \P2_State2_reg[2]/NET0131  ;
	input \P2_State2_reg[3]/NET0131  ;
	input \P2_State_reg[0]/NET0131  ;
	input \P2_State_reg[1]/NET0131  ;
	input \P2_State_reg[2]/NET0131  ;
	input \P2_W_R_n_reg/NET0131  ;
	input \P2_lWord_reg[0]/NET0131  ;
	input \P2_lWord_reg[10]/NET0131  ;
	input \P2_lWord_reg[11]/NET0131  ;
	input \P2_lWord_reg[12]/NET0131  ;
	input \P2_lWord_reg[13]/NET0131  ;
	input \P2_lWord_reg[14]/NET0131  ;
	input \P2_lWord_reg[15]/NET0131  ;
	input \P2_lWord_reg[1]/NET0131  ;
	input \P2_lWord_reg[2]/NET0131  ;
	input \P2_lWord_reg[3]/NET0131  ;
	input \P2_lWord_reg[4]/NET0131  ;
	input \P2_lWord_reg[5]/NET0131  ;
	input \P2_lWord_reg[6]/NET0131  ;
	input \P2_lWord_reg[7]/NET0131  ;
	input \P2_lWord_reg[8]/NET0131  ;
	input \P2_lWord_reg[9]/NET0131  ;
	input \P2_rEIP_reg[0]/NET0131  ;
	input \P2_rEIP_reg[10]/NET0131  ;
	input \P2_rEIP_reg[11]/NET0131  ;
	input \P2_rEIP_reg[12]/NET0131  ;
	input \P2_rEIP_reg[13]/NET0131  ;
	input \P2_rEIP_reg[14]/NET0131  ;
	input \P2_rEIP_reg[15]/NET0131  ;
	input \P2_rEIP_reg[16]/NET0131  ;
	input \P2_rEIP_reg[17]/NET0131  ;
	input \P2_rEIP_reg[18]/NET0131  ;
	input \P2_rEIP_reg[19]/NET0131  ;
	input \P2_rEIP_reg[1]/NET0131  ;
	input \P2_rEIP_reg[20]/NET0131  ;
	input \P2_rEIP_reg[21]/NET0131  ;
	input \P2_rEIP_reg[22]/NET0131  ;
	input \P2_rEIP_reg[23]/NET0131  ;
	input \P2_rEIP_reg[24]/NET0131  ;
	input \P2_rEIP_reg[25]/NET0131  ;
	input \P2_rEIP_reg[26]/NET0131  ;
	input \P2_rEIP_reg[27]/NET0131  ;
	input \P2_rEIP_reg[28]/NET0131  ;
	input \P2_rEIP_reg[29]/NET0131  ;
	input \P2_rEIP_reg[2]/NET0131  ;
	input \P2_rEIP_reg[30]/NET0131  ;
	input \P2_rEIP_reg[31]/NET0131  ;
	input \P2_rEIP_reg[3]/NET0131  ;
	input \P2_rEIP_reg[4]/NET0131  ;
	input \P2_rEIP_reg[5]/NET0131  ;
	input \P2_rEIP_reg[6]/NET0131  ;
	input \P2_rEIP_reg[7]/NET0131  ;
	input \P2_rEIP_reg[8]/NET0131  ;
	input \P2_rEIP_reg[9]/NET0131  ;
	input \P2_uWord_reg[0]/NET0131  ;
	input \P2_uWord_reg[10]/NET0131  ;
	input \P2_uWord_reg[11]/NET0131  ;
	input \P2_uWord_reg[12]/NET0131  ;
	input \P2_uWord_reg[13]/NET0131  ;
	input \P2_uWord_reg[14]/NET0131  ;
	input \P2_uWord_reg[1]/NET0131  ;
	input \P2_uWord_reg[2]/NET0131  ;
	input \P2_uWord_reg[3]/NET0131  ;
	input \P2_uWord_reg[4]/NET0131  ;
	input \P2_uWord_reg[5]/NET0131  ;
	input \P2_uWord_reg[6]/NET0131  ;
	input \P2_uWord_reg[7]/NET0131  ;
	input \P2_uWord_reg[8]/NET0131  ;
	input \P2_uWord_reg[9]/NET0131  ;
	input \P3_Address_reg[0]/NET0131  ;
	input \P3_Address_reg[10]/NET0131  ;
	input \P3_Address_reg[11]/NET0131  ;
	input \P3_Address_reg[12]/NET0131  ;
	input \P3_Address_reg[13]/NET0131  ;
	input \P3_Address_reg[14]/NET0131  ;
	input \P3_Address_reg[15]/NET0131  ;
	input \P3_Address_reg[16]/NET0131  ;
	input \P3_Address_reg[17]/NET0131  ;
	input \P3_Address_reg[18]/NET0131  ;
	input \P3_Address_reg[19]/NET0131  ;
	input \P3_Address_reg[1]/NET0131  ;
	input \P3_Address_reg[20]/NET0131  ;
	input \P3_Address_reg[21]/NET0131  ;
	input \P3_Address_reg[22]/NET0131  ;
	input \P3_Address_reg[23]/NET0131  ;
	input \P3_Address_reg[24]/NET0131  ;
	input \P3_Address_reg[25]/NET0131  ;
	input \P3_Address_reg[26]/NET0131  ;
	input \P3_Address_reg[27]/NET0131  ;
	input \P3_Address_reg[28]/NET0131  ;
	input \P3_Address_reg[29]/NET0131  ;
	input \P3_Address_reg[2]/NET0131  ;
	input \P3_Address_reg[3]/NET0131  ;
	input \P3_Address_reg[4]/NET0131  ;
	input \P3_Address_reg[5]/NET0131  ;
	input \P3_Address_reg[6]/NET0131  ;
	input \P3_Address_reg[7]/NET0131  ;
	input \P3_Address_reg[8]/NET0131  ;
	input \P3_Address_reg[9]/NET0131  ;
	input \P3_BE_n_reg[0]/NET0131  ;
	input \P3_BE_n_reg[1]/NET0131  ;
	input \P3_BE_n_reg[2]/NET0131  ;
	input \P3_BE_n_reg[3]/NET0131  ;
	input \P3_ByteEnable_reg[0]/NET0131  ;
	input \P3_ByteEnable_reg[1]/NET0131  ;
	input \P3_ByteEnable_reg[2]/NET0131  ;
	input \P3_ByteEnable_reg[3]/NET0131  ;
	input \P3_CodeFetch_reg/NET0131  ;
	input \P3_DataWidth_reg[0]/NET0131  ;
	input \P3_DataWidth_reg[1]/NET0131  ;
	input \P3_EAX_reg[0]/NET0131  ;
	input \P3_EAX_reg[10]/NET0131  ;
	input \P3_EAX_reg[11]/NET0131  ;
	input \P3_EAX_reg[12]/NET0131  ;
	input \P3_EAX_reg[13]/NET0131  ;
	input \P3_EAX_reg[14]/NET0131  ;
	input \P3_EAX_reg[15]/NET0131  ;
	input \P3_EAX_reg[16]/NET0131  ;
	input \P3_EAX_reg[17]/NET0131  ;
	input \P3_EAX_reg[18]/NET0131  ;
	input \P3_EAX_reg[19]/NET0131  ;
	input \P3_EAX_reg[1]/NET0131  ;
	input \P3_EAX_reg[20]/NET0131  ;
	input \P3_EAX_reg[21]/NET0131  ;
	input \P3_EAX_reg[22]/NET0131  ;
	input \P3_EAX_reg[23]/NET0131  ;
	input \P3_EAX_reg[24]/NET0131  ;
	input \P3_EAX_reg[25]/NET0131  ;
	input \P3_EAX_reg[26]/NET0131  ;
	input \P3_EAX_reg[27]/NET0131  ;
	input \P3_EAX_reg[28]/NET0131  ;
	input \P3_EAX_reg[29]/NET0131  ;
	input \P3_EAX_reg[2]/NET0131  ;
	input \P3_EAX_reg[30]/NET0131  ;
	input \P3_EAX_reg[31]/NET0131  ;
	input \P3_EAX_reg[3]/NET0131  ;
	input \P3_EAX_reg[4]/NET0131  ;
	input \P3_EAX_reg[5]/NET0131  ;
	input \P3_EAX_reg[6]/NET0131  ;
	input \P3_EAX_reg[7]/NET0131  ;
	input \P3_EAX_reg[8]/NET0131  ;
	input \P3_EAX_reg[9]/NET0131  ;
	input \P3_EBX_reg[0]/NET0131  ;
	input \P3_EBX_reg[10]/NET0131  ;
	input \P3_EBX_reg[11]/NET0131  ;
	input \P3_EBX_reg[12]/NET0131  ;
	input \P3_EBX_reg[13]/NET0131  ;
	input \P3_EBX_reg[14]/NET0131  ;
	input \P3_EBX_reg[15]/NET0131  ;
	input \P3_EBX_reg[16]/NET0131  ;
	input \P3_EBX_reg[17]/NET0131  ;
	input \P3_EBX_reg[18]/NET0131  ;
	input \P3_EBX_reg[19]/NET0131  ;
	input \P3_EBX_reg[1]/NET0131  ;
	input \P3_EBX_reg[20]/NET0131  ;
	input \P3_EBX_reg[21]/NET0131  ;
	input \P3_EBX_reg[22]/NET0131  ;
	input \P3_EBX_reg[23]/NET0131  ;
	input \P3_EBX_reg[24]/NET0131  ;
	input \P3_EBX_reg[25]/NET0131  ;
	input \P3_EBX_reg[26]/NET0131  ;
	input \P3_EBX_reg[27]/NET0131  ;
	input \P3_EBX_reg[28]/NET0131  ;
	input \P3_EBX_reg[29]/NET0131  ;
	input \P3_EBX_reg[2]/NET0131  ;
	input \P3_EBX_reg[30]/NET0131  ;
	input \P3_EBX_reg[31]/NET0131  ;
	input \P3_EBX_reg[3]/NET0131  ;
	input \P3_EBX_reg[4]/NET0131  ;
	input \P3_EBX_reg[5]/NET0131  ;
	input \P3_EBX_reg[6]/NET0131  ;
	input \P3_EBX_reg[7]/NET0131  ;
	input \P3_EBX_reg[8]/NET0131  ;
	input \P3_EBX_reg[9]/NET0131  ;
	input \P3_Flush_reg/NET0131  ;
	input \P3_InstAddrPointer_reg[0]/NET0131  ;
	input \P3_InstAddrPointer_reg[10]/NET0131  ;
	input \P3_InstAddrPointer_reg[11]/NET0131  ;
	input \P3_InstAddrPointer_reg[12]/NET0131  ;
	input \P3_InstAddrPointer_reg[13]/NET0131  ;
	input \P3_InstAddrPointer_reg[14]/NET0131  ;
	input \P3_InstAddrPointer_reg[15]/NET0131  ;
	input \P3_InstAddrPointer_reg[16]/NET0131  ;
	input \P3_InstAddrPointer_reg[17]/NET0131  ;
	input \P3_InstAddrPointer_reg[18]/NET0131  ;
	input \P3_InstAddrPointer_reg[19]/NET0131  ;
	input \P3_InstAddrPointer_reg[1]/NET0131  ;
	input \P3_InstAddrPointer_reg[20]/NET0131  ;
	input \P3_InstAddrPointer_reg[21]/NET0131  ;
	input \P3_InstAddrPointer_reg[22]/NET0131  ;
	input \P3_InstAddrPointer_reg[23]/NET0131  ;
	input \P3_InstAddrPointer_reg[24]/NET0131  ;
	input \P3_InstAddrPointer_reg[25]/NET0131  ;
	input \P3_InstAddrPointer_reg[26]/NET0131  ;
	input \P3_InstAddrPointer_reg[27]/NET0131  ;
	input \P3_InstAddrPointer_reg[28]/NET0131  ;
	input \P3_InstAddrPointer_reg[29]/NET0131  ;
	input \P3_InstAddrPointer_reg[2]/NET0131  ;
	input \P3_InstAddrPointer_reg[30]/NET0131  ;
	input \P3_InstAddrPointer_reg[31]/NET0131  ;
	input \P3_InstAddrPointer_reg[3]/NET0131  ;
	input \P3_InstAddrPointer_reg[4]/NET0131  ;
	input \P3_InstAddrPointer_reg[5]/NET0131  ;
	input \P3_InstAddrPointer_reg[6]/NET0131  ;
	input \P3_InstAddrPointer_reg[7]/NET0131  ;
	input \P3_InstAddrPointer_reg[8]/NET0131  ;
	input \P3_InstAddrPointer_reg[9]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[0]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[2]/NET0131  ;
	input \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[0]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[2]/NET0131  ;
	input \P3_InstQueueWr_Addr_reg[3]/NET0131  ;
	input \P3_InstQueue_reg[0][0]/NET0131  ;
	input \P3_InstQueue_reg[0][1]/NET0131  ;
	input \P3_InstQueue_reg[0][2]/NET0131  ;
	input \P3_InstQueue_reg[0][3]/NET0131  ;
	input \P3_InstQueue_reg[0][4]/NET0131  ;
	input \P3_InstQueue_reg[0][5]/NET0131  ;
	input \P3_InstQueue_reg[0][6]/NET0131  ;
	input \P3_InstQueue_reg[0][7]/NET0131  ;
	input \P3_InstQueue_reg[10][0]/NET0131  ;
	input \P3_InstQueue_reg[10][1]/NET0131  ;
	input \P3_InstQueue_reg[10][2]/NET0131  ;
	input \P3_InstQueue_reg[10][3]/NET0131  ;
	input \P3_InstQueue_reg[10][4]/NET0131  ;
	input \P3_InstQueue_reg[10][5]/NET0131  ;
	input \P3_InstQueue_reg[10][6]/NET0131  ;
	input \P3_InstQueue_reg[10][7]/NET0131  ;
	input \P3_InstQueue_reg[11][0]/NET0131  ;
	input \P3_InstQueue_reg[11][1]/NET0131  ;
	input \P3_InstQueue_reg[11][2]/NET0131  ;
	input \P3_InstQueue_reg[11][3]/NET0131  ;
	input \P3_InstQueue_reg[11][4]/NET0131  ;
	input \P3_InstQueue_reg[11][5]/NET0131  ;
	input \P3_InstQueue_reg[11][6]/NET0131  ;
	input \P3_InstQueue_reg[11][7]/NET0131  ;
	input \P3_InstQueue_reg[12][0]/NET0131  ;
	input \P3_InstQueue_reg[12][1]/NET0131  ;
	input \P3_InstQueue_reg[12][2]/NET0131  ;
	input \P3_InstQueue_reg[12][3]/NET0131  ;
	input \P3_InstQueue_reg[12][4]/NET0131  ;
	input \P3_InstQueue_reg[12][5]/NET0131  ;
	input \P3_InstQueue_reg[12][6]/NET0131  ;
	input \P3_InstQueue_reg[12][7]/NET0131  ;
	input \P3_InstQueue_reg[13][0]/NET0131  ;
	input \P3_InstQueue_reg[13][1]/NET0131  ;
	input \P3_InstQueue_reg[13][2]/NET0131  ;
	input \P3_InstQueue_reg[13][3]/NET0131  ;
	input \P3_InstQueue_reg[13][4]/NET0131  ;
	input \P3_InstQueue_reg[13][5]/NET0131  ;
	input \P3_InstQueue_reg[13][6]/NET0131  ;
	input \P3_InstQueue_reg[13][7]/NET0131  ;
	input \P3_InstQueue_reg[14][0]/NET0131  ;
	input \P3_InstQueue_reg[14][1]/NET0131  ;
	input \P3_InstQueue_reg[14][2]/NET0131  ;
	input \P3_InstQueue_reg[14][3]/NET0131  ;
	input \P3_InstQueue_reg[14][4]/NET0131  ;
	input \P3_InstQueue_reg[14][5]/NET0131  ;
	input \P3_InstQueue_reg[14][6]/NET0131  ;
	input \P3_InstQueue_reg[14][7]/NET0131  ;
	input \P3_InstQueue_reg[15][0]/NET0131  ;
	input \P3_InstQueue_reg[15][1]/NET0131  ;
	input \P3_InstQueue_reg[15][2]/NET0131  ;
	input \P3_InstQueue_reg[15][3]/NET0131  ;
	input \P3_InstQueue_reg[15][4]/NET0131  ;
	input \P3_InstQueue_reg[15][5]/NET0131  ;
	input \P3_InstQueue_reg[15][6]/NET0131  ;
	input \P3_InstQueue_reg[15][7]/NET0131  ;
	input \P3_InstQueue_reg[1][0]/NET0131  ;
	input \P3_InstQueue_reg[1][1]/NET0131  ;
	input \P3_InstQueue_reg[1][2]/NET0131  ;
	input \P3_InstQueue_reg[1][3]/NET0131  ;
	input \P3_InstQueue_reg[1][4]/NET0131  ;
	input \P3_InstQueue_reg[1][5]/NET0131  ;
	input \P3_InstQueue_reg[1][6]/NET0131  ;
	input \P3_InstQueue_reg[1][7]/NET0131  ;
	input \P3_InstQueue_reg[2][0]/NET0131  ;
	input \P3_InstQueue_reg[2][1]/NET0131  ;
	input \P3_InstQueue_reg[2][2]/NET0131  ;
	input \P3_InstQueue_reg[2][3]/NET0131  ;
	input \P3_InstQueue_reg[2][4]/NET0131  ;
	input \P3_InstQueue_reg[2][5]/NET0131  ;
	input \P3_InstQueue_reg[2][6]/NET0131  ;
	input \P3_InstQueue_reg[2][7]/NET0131  ;
	input \P3_InstQueue_reg[3][0]/NET0131  ;
	input \P3_InstQueue_reg[3][1]/NET0131  ;
	input \P3_InstQueue_reg[3][2]/NET0131  ;
	input \P3_InstQueue_reg[3][3]/NET0131  ;
	input \P3_InstQueue_reg[3][4]/NET0131  ;
	input \P3_InstQueue_reg[3][5]/NET0131  ;
	input \P3_InstQueue_reg[3][6]/NET0131  ;
	input \P3_InstQueue_reg[3][7]/NET0131  ;
	input \P3_InstQueue_reg[4][0]/NET0131  ;
	input \P3_InstQueue_reg[4][1]/NET0131  ;
	input \P3_InstQueue_reg[4][2]/NET0131  ;
	input \P3_InstQueue_reg[4][3]/NET0131  ;
	input \P3_InstQueue_reg[4][4]/NET0131  ;
	input \P3_InstQueue_reg[4][5]/NET0131  ;
	input \P3_InstQueue_reg[4][6]/NET0131  ;
	input \P3_InstQueue_reg[4][7]/NET0131  ;
	input \P3_InstQueue_reg[5][0]/NET0131  ;
	input \P3_InstQueue_reg[5][1]/NET0131  ;
	input \P3_InstQueue_reg[5][2]/NET0131  ;
	input \P3_InstQueue_reg[5][3]/NET0131  ;
	input \P3_InstQueue_reg[5][4]/NET0131  ;
	input \P3_InstQueue_reg[5][5]/NET0131  ;
	input \P3_InstQueue_reg[5][6]/NET0131  ;
	input \P3_InstQueue_reg[5][7]/NET0131  ;
	input \P3_InstQueue_reg[6][0]/NET0131  ;
	input \P3_InstQueue_reg[6][1]/NET0131  ;
	input \P3_InstQueue_reg[6][2]/NET0131  ;
	input \P3_InstQueue_reg[6][3]/NET0131  ;
	input \P3_InstQueue_reg[6][4]/NET0131  ;
	input \P3_InstQueue_reg[6][5]/NET0131  ;
	input \P3_InstQueue_reg[6][6]/NET0131  ;
	input \P3_InstQueue_reg[6][7]/NET0131  ;
	input \P3_InstQueue_reg[7][0]/NET0131  ;
	input \P3_InstQueue_reg[7][1]/NET0131  ;
	input \P3_InstQueue_reg[7][2]/NET0131  ;
	input \P3_InstQueue_reg[7][3]/NET0131  ;
	input \P3_InstQueue_reg[7][4]/NET0131  ;
	input \P3_InstQueue_reg[7][5]/NET0131  ;
	input \P3_InstQueue_reg[7][6]/NET0131  ;
	input \P3_InstQueue_reg[7][7]/NET0131  ;
	input \P3_InstQueue_reg[8][0]/NET0131  ;
	input \P3_InstQueue_reg[8][1]/NET0131  ;
	input \P3_InstQueue_reg[8][2]/NET0131  ;
	input \P3_InstQueue_reg[8][3]/NET0131  ;
	input \P3_InstQueue_reg[8][4]/NET0131  ;
	input \P3_InstQueue_reg[8][5]/NET0131  ;
	input \P3_InstQueue_reg[8][6]/NET0131  ;
	input \P3_InstQueue_reg[8][7]/NET0131  ;
	input \P3_InstQueue_reg[9][0]/NET0131  ;
	input \P3_InstQueue_reg[9][1]/NET0131  ;
	input \P3_InstQueue_reg[9][2]/NET0131  ;
	input \P3_InstQueue_reg[9][3]/NET0131  ;
	input \P3_InstQueue_reg[9][4]/NET0131  ;
	input \P3_InstQueue_reg[9][5]/NET0131  ;
	input \P3_InstQueue_reg[9][6]/NET0131  ;
	input \P3_InstQueue_reg[9][7]/NET0131  ;
	input \P3_MemoryFetch_reg/NET0131  ;
	input \P3_More_reg/NET0131  ;
	input \P3_PhyAddrPointer_reg[0]/NET0131  ;
	input \P3_PhyAddrPointer_reg[10]/NET0131  ;
	input \P3_PhyAddrPointer_reg[11]/NET0131  ;
	input \P3_PhyAddrPointer_reg[12]/NET0131  ;
	input \P3_PhyAddrPointer_reg[13]/NET0131  ;
	input \P3_PhyAddrPointer_reg[14]/NET0131  ;
	input \P3_PhyAddrPointer_reg[15]/NET0131  ;
	input \P3_PhyAddrPointer_reg[16]/NET0131  ;
	input \P3_PhyAddrPointer_reg[17]/NET0131  ;
	input \P3_PhyAddrPointer_reg[18]/NET0131  ;
	input \P3_PhyAddrPointer_reg[19]/NET0131  ;
	input \P3_PhyAddrPointer_reg[1]/NET0131  ;
	input \P3_PhyAddrPointer_reg[20]/NET0131  ;
	input \P3_PhyAddrPointer_reg[21]/NET0131  ;
	input \P3_PhyAddrPointer_reg[22]/NET0131  ;
	input \P3_PhyAddrPointer_reg[23]/NET0131  ;
	input \P3_PhyAddrPointer_reg[24]/NET0131  ;
	input \P3_PhyAddrPointer_reg[25]/NET0131  ;
	input \P3_PhyAddrPointer_reg[26]/NET0131  ;
	input \P3_PhyAddrPointer_reg[27]/NET0131  ;
	input \P3_PhyAddrPointer_reg[28]/NET0131  ;
	input \P3_PhyAddrPointer_reg[29]/NET0131  ;
	input \P3_PhyAddrPointer_reg[2]/NET0131  ;
	input \P3_PhyAddrPointer_reg[30]/NET0131  ;
	input \P3_PhyAddrPointer_reg[31]/NET0131  ;
	input \P3_PhyAddrPointer_reg[3]/NET0131  ;
	input \P3_PhyAddrPointer_reg[4]/NET0131  ;
	input \P3_PhyAddrPointer_reg[5]/NET0131  ;
	input \P3_PhyAddrPointer_reg[6]/NET0131  ;
	input \P3_PhyAddrPointer_reg[7]/NET0131  ;
	input \P3_PhyAddrPointer_reg[8]/NET0131  ;
	input \P3_PhyAddrPointer_reg[9]/NET0131  ;
	input \P3_ReadRequest_reg/NET0131  ;
	input \P3_RequestPending_reg/NET0131  ;
	input \P3_State2_reg[0]/NET0131  ;
	input \P3_State2_reg[1]/NET0131  ;
	input \P3_State2_reg[2]/NET0131  ;
	input \P3_State2_reg[3]/NET0131  ;
	input \P3_State_reg[0]/NET0131  ;
	input \P3_State_reg[1]/NET0131  ;
	input \P3_State_reg[2]/NET0131  ;
	input \P3_lWord_reg[0]/NET0131  ;
	input \P3_lWord_reg[10]/NET0131  ;
	input \P3_lWord_reg[11]/NET0131  ;
	input \P3_lWord_reg[12]/NET0131  ;
	input \P3_lWord_reg[13]/NET0131  ;
	input \P3_lWord_reg[14]/NET0131  ;
	input \P3_lWord_reg[15]/NET0131  ;
	input \P3_lWord_reg[1]/NET0131  ;
	input \P3_lWord_reg[2]/NET0131  ;
	input \P3_lWord_reg[3]/NET0131  ;
	input \P3_lWord_reg[4]/NET0131  ;
	input \P3_lWord_reg[5]/NET0131  ;
	input \P3_lWord_reg[6]/NET0131  ;
	input \P3_lWord_reg[7]/NET0131  ;
	input \P3_lWord_reg[8]/NET0131  ;
	input \P3_lWord_reg[9]/NET0131  ;
	input \P3_rEIP_reg[0]/NET0131  ;
	input \P3_rEIP_reg[10]/NET0131  ;
	input \P3_rEIP_reg[11]/NET0131  ;
	input \P3_rEIP_reg[12]/NET0131  ;
	input \P3_rEIP_reg[13]/NET0131  ;
	input \P3_rEIP_reg[14]/NET0131  ;
	input \P3_rEIP_reg[15]/NET0131  ;
	input \P3_rEIP_reg[16]/NET0131  ;
	input \P3_rEIP_reg[17]/NET0131  ;
	input \P3_rEIP_reg[18]/NET0131  ;
	input \P3_rEIP_reg[19]/NET0131  ;
	input \P3_rEIP_reg[1]/NET0131  ;
	input \P3_rEIP_reg[20]/NET0131  ;
	input \P3_rEIP_reg[21]/NET0131  ;
	input \P3_rEIP_reg[22]/NET0131  ;
	input \P3_rEIP_reg[23]/NET0131  ;
	input \P3_rEIP_reg[24]/NET0131  ;
	input \P3_rEIP_reg[25]/NET0131  ;
	input \P3_rEIP_reg[26]/NET0131  ;
	input \P3_rEIP_reg[27]/NET0131  ;
	input \P3_rEIP_reg[28]/NET0131  ;
	input \P3_rEIP_reg[29]/NET0131  ;
	input \P3_rEIP_reg[2]/NET0131  ;
	input \P3_rEIP_reg[30]/NET0131  ;
	input \P3_rEIP_reg[31]/NET0131  ;
	input \P3_rEIP_reg[3]/NET0131  ;
	input \P3_rEIP_reg[4]/NET0131  ;
	input \P3_rEIP_reg[5]/NET0131  ;
	input \P3_rEIP_reg[6]/NET0131  ;
	input \P3_rEIP_reg[7]/NET0131  ;
	input \P3_rEIP_reg[8]/NET0131  ;
	input \P3_rEIP_reg[9]/NET0131  ;
	input \P3_uWord_reg[0]/NET0131  ;
	input \P3_uWord_reg[10]/NET0131  ;
	input \P3_uWord_reg[11]/NET0131  ;
	input \P3_uWord_reg[12]/NET0131  ;
	input \P3_uWord_reg[13]/NET0131  ;
	input \P3_uWord_reg[14]/NET0131  ;
	input \P3_uWord_reg[1]/NET0131  ;
	input \P3_uWord_reg[2]/NET0131  ;
	input \P3_uWord_reg[3]/NET0131  ;
	input \P3_uWord_reg[4]/NET0131  ;
	input \P3_uWord_reg[5]/NET0131  ;
	input \P3_uWord_reg[6]/NET0131  ;
	input \P3_uWord_reg[7]/NET0131  ;
	input \P3_uWord_reg[8]/NET0131  ;
	input \P3_uWord_reg[9]/NET0131  ;
	input \address1[0]_pad  ;
	input \address1[10]_pad  ;
	input \address1[11]_pad  ;
	input \address1[12]_pad  ;
	input \address1[13]_pad  ;
	input \address1[14]_pad  ;
	input \address1[15]_pad  ;
	input \address1[16]_pad  ;
	input \address1[17]_pad  ;
	input \address1[18]_pad  ;
	input \address1[19]_pad  ;
	input \address1[1]_pad  ;
	input \address1[20]_pad  ;
	input \address1[21]_pad  ;
	input \address1[22]_pad  ;
	input \address1[23]_pad  ;
	input \address1[24]_pad  ;
	input \address1[25]_pad  ;
	input \address1[26]_pad  ;
	input \address1[27]_pad  ;
	input \address1[28]_pad  ;
	input \address1[29]_pad  ;
	input \address1[2]_pad  ;
	input \address1[3]_pad  ;
	input \address1[4]_pad  ;
	input \address1[5]_pad  ;
	input \address1[6]_pad  ;
	input \address1[7]_pad  ;
	input \address1[8]_pad  ;
	input \address1[9]_pad  ;
	input \ast1_pad  ;
	input \ast2_pad  ;
	input \bs16_pad  ;
	input \buf1_reg[0]/NET0131  ;
	input \buf1_reg[10]/NET0131  ;
	input \buf1_reg[11]/NET0131  ;
	input \buf1_reg[12]/NET0131  ;
	input \buf1_reg[13]/NET0131  ;
	input \buf1_reg[14]/NET0131  ;
	input \buf1_reg[15]/NET0131  ;
	input \buf1_reg[16]/NET0131  ;
	input \buf1_reg[17]/NET0131  ;
	input \buf1_reg[18]/NET0131  ;
	input \buf1_reg[19]/NET0131  ;
	input \buf1_reg[1]/NET0131  ;
	input \buf1_reg[20]/NET0131  ;
	input \buf1_reg[21]/NET0131  ;
	input \buf1_reg[22]/NET0131  ;
	input \buf1_reg[23]/NET0131  ;
	input \buf1_reg[24]/NET0131  ;
	input \buf1_reg[25]/NET0131  ;
	input \buf1_reg[26]/NET0131  ;
	input \buf1_reg[27]/NET0131  ;
	input \buf1_reg[28]/NET0131  ;
	input \buf1_reg[29]/NET0131  ;
	input \buf1_reg[2]/NET0131  ;
	input \buf1_reg[30]/NET0131  ;
	input \buf1_reg[3]/NET0131  ;
	input \buf1_reg[4]/NET0131  ;
	input \buf1_reg[5]/NET0131  ;
	input \buf1_reg[6]/NET0131  ;
	input \buf1_reg[7]/NET0131  ;
	input \buf1_reg[8]/NET0131  ;
	input \buf1_reg[9]/NET0131  ;
	input \buf2_reg[0]/NET0131  ;
	input \buf2_reg[10]/NET0131  ;
	input \buf2_reg[11]/NET0131  ;
	input \buf2_reg[12]/NET0131  ;
	input \buf2_reg[13]/NET0131  ;
	input \buf2_reg[14]/NET0131  ;
	input \buf2_reg[15]/NET0131  ;
	input \buf2_reg[16]/NET0131  ;
	input \buf2_reg[17]/NET0131  ;
	input \buf2_reg[18]/NET0131  ;
	input \buf2_reg[19]/NET0131  ;
	input \buf2_reg[1]/NET0131  ;
	input \buf2_reg[20]/NET0131  ;
	input \buf2_reg[21]/NET0131  ;
	input \buf2_reg[22]/NET0131  ;
	input \buf2_reg[23]/NET0131  ;
	input \buf2_reg[24]/NET0131  ;
	input \buf2_reg[25]/NET0131  ;
	input \buf2_reg[26]/NET0131  ;
	input \buf2_reg[27]/NET0131  ;
	input \buf2_reg[28]/NET0131  ;
	input \buf2_reg[29]/NET0131  ;
	input \buf2_reg[2]/NET0131  ;
	input \buf2_reg[30]/NET0131  ;
	input \buf2_reg[3]/NET0131  ;
	input \buf2_reg[4]/NET0131  ;
	input \buf2_reg[5]/NET0131  ;
	input \buf2_reg[6]/NET0131  ;
	input \buf2_reg[7]/NET0131  ;
	input \buf2_reg[8]/NET0131  ;
	input \buf2_reg[9]/NET0131  ;
	input \datai[0]_pad  ;
	input \datai[10]_pad  ;
	input \datai[11]_pad  ;
	input \datai[12]_pad  ;
	input \datai[13]_pad  ;
	input \datai[14]_pad  ;
	input \datai[15]_pad  ;
	input \datai[16]_pad  ;
	input \datai[17]_pad  ;
	input \datai[18]_pad  ;
	input \datai[19]_pad  ;
	input \datai[1]_pad  ;
	input \datai[20]_pad  ;
	input \datai[21]_pad  ;
	input \datai[22]_pad  ;
	input \datai[23]_pad  ;
	input \datai[24]_pad  ;
	input \datai[25]_pad  ;
	input \datai[26]_pad  ;
	input \datai[27]_pad  ;
	input \datai[28]_pad  ;
	input \datai[29]_pad  ;
	input \datai[2]_pad  ;
	input \datai[30]_pad  ;
	input \datai[31]_pad  ;
	input \datai[3]_pad  ;
	input \datai[4]_pad  ;
	input \datai[5]_pad  ;
	input \datai[6]_pad  ;
	input \datai[7]_pad  ;
	input \datai[8]_pad  ;
	input \datai[9]_pad  ;
	input \datao[0]_pad  ;
	input \datao[10]_pad  ;
	input \datao[11]_pad  ;
	input \datao[12]_pad  ;
	input \datao[13]_pad  ;
	input \datao[14]_pad  ;
	input \datao[15]_pad  ;
	input \datao[16]_pad  ;
	input \datao[17]_pad  ;
	input \datao[18]_pad  ;
	input \datao[19]_pad  ;
	input \datao[1]_pad  ;
	input \datao[20]_pad  ;
	input \datao[21]_pad  ;
	input \datao[22]_pad  ;
	input \datao[23]_pad  ;
	input \datao[24]_pad  ;
	input \datao[25]_pad  ;
	input \datao[26]_pad  ;
	input \datao[27]_pad  ;
	input \datao[28]_pad  ;
	input \datao[29]_pad  ;
	input \datao[2]_pad  ;
	input \datao[30]_pad  ;
	input \datao[3]_pad  ;
	input \datao[4]_pad  ;
	input \datao[5]_pad  ;
	input \datao[6]_pad  ;
	input \datao[7]_pad  ;
	input \datao[8]_pad  ;
	input \datao[9]_pad  ;
	input dc_pad ;
	input hold_pad ;
	input mio_pad ;
	input na_pad ;
	input \ready11_reg/NET0131  ;
	input \ready12_reg/NET0131  ;
	input \ready1_pad  ;
	input \ready21_reg/NET0131  ;
	input \ready22_reg/NET0131  ;
	input \ready2_pad  ;
	input wr_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \address2[0]_pad  ;
	output \address2[10]_pad  ;
	output \address2[11]_pad  ;
	output \address2[12]_pad  ;
	output \address2[13]_pad  ;
	output \address2[14]_pad  ;
	output \address2[15]_pad  ;
	output \address2[16]_pad  ;
	output \address2[17]_pad  ;
	output \address2[18]_pad  ;
	output \address2[19]_pad  ;
	output \address2[1]_pad  ;
	output \address2[20]_pad  ;
	output \address2[21]_pad  ;
	output \address2[22]_pad  ;
	output \address2[23]_pad  ;
	output \address2[24]_pad  ;
	output \address2[25]_pad  ;
	output \address2[26]_pad  ;
	output \address2[27]_pad  ;
	output \address2[28]_pad  ;
	output \address2[29]_pad  ;
	output \address2[2]_pad  ;
	output \address2[3]_pad  ;
	output \address2[4]_pad  ;
	output \address2[5]_pad  ;
	output \address2[6]_pad  ;
	output \address2[7]_pad  ;
	output \address2[8]_pad  ;
	output \address2[9]_pad  ;
	output \g133468/_2_  ;
	output \g133469/_2_  ;
	output \g133470/_2_  ;
	output \g133475/_0_  ;
	output \g133476/_2_  ;
	output \g133515/_0_  ;
	output \g133516/_0_  ;
	output \g133517/_0_  ;
	output \g133518/_0_  ;
	output \g133523/_0_  ;
	output \g133524/_0_  ;
	output \g133528/_0_  ;
	output \g133529/_0_  ;
	output \g133531/_0_  ;
	output \g133532/_0_  ;
	output \g133533/_0_  ;
	output \g133534/_0_  ;
	output \g133535/_0_  ;
	output \g133536/_0_  ;
	output \g133537/_0_  ;
	output \g133538/_0_  ;
	output \g133539/_0_  ;
	output \g133540/_0_  ;
	output \g133541/_0_  ;
	output \g133542/_0_  ;
	output \g133543/_0_  ;
	output \g133544/_0_  ;
	output \g133545/_0_  ;
	output \g133546/_0_  ;
	output \g133547/_0_  ;
	output \g133548/_0_  ;
	output \g133549/_0_  ;
	output \g133550/_0_  ;
	output \g133551/_0_  ;
	output \g133552/_0_  ;
	output \g133553/_0_  ;
	output \g133554/_0_  ;
	output \g133555/_0_  ;
	output \g133556/_0_  ;
	output \g133557/_0_  ;
	output \g133558/_0_  ;
	output \g133559/_0_  ;
	output \g133560/_0_  ;
	output \g133561/_0_  ;
	output \g133566/_0_  ;
	output \g133619/_0_  ;
	output \g133659/_0_  ;
	output \g133660/_0_  ;
	output \g133662/_0_  ;
	output \g133663/_0_  ;
	output \g133664/_0_  ;
	output \g133665/_0_  ;
	output \g133666/_0_  ;
	output \g133667/_0_  ;
	output \g133668/_0_  ;
	output \g133669/_0_  ;
	output \g133670/_0_  ;
	output \g133671/_0_  ;
	output \g133672/_0_  ;
	output \g133673/_0_  ;
	output \g133674/_0_  ;
	output \g133675/_0_  ;
	output \g133676/_0_  ;
	output \g133677/_0_  ;
	output \g133678/_0_  ;
	output \g133679/_0_  ;
	output \g133680/_0_  ;
	output \g133681/_0_  ;
	output \g133682/_0_  ;
	output \g133683/_0_  ;
	output \g133684/_0_  ;
	output \g133685/_0_  ;
	output \g133686/_0_  ;
	output \g133687/_0_  ;
	output \g133688/_0_  ;
	output \g133689/_0_  ;
	output \g133690/_0_  ;
	output \g133691/_0_  ;
	output \g133694/_0_  ;
	output \g133697/_0_  ;
	output \g133702/_0_  ;
	output \g133703/_0_  ;
	output \g133756/_0_  ;
	output \g133792/_0_  ;
	output \g133793/_0_  ;
	output \g133794/_0_  ;
	output \g133796/_0_  ;
	output \g133797/_0_  ;
	output \g133798/_0_  ;
	output \g133799/_0_  ;
	output \g133800/_0_  ;
	output \g133801/_0_  ;
	output \g133802/_0_  ;
	output \g133803/_0_  ;
	output \g133804/_0_  ;
	output \g133806/_0_  ;
	output \g133807/_0_  ;
	output \g133808/_0_  ;
	output \g133812/_0_  ;
	output \g133813/_0_  ;
	output \g133814/_0_  ;
	output \g133817/_0_  ;
	output \g133821/_0_  ;
	output \g133824/_0_  ;
	output \g133826/_0_  ;
	output \g133828/_0_  ;
	output \g133864/_0_  ;
	output \g133865/_0_  ;
	output \g133867/_0_  ;
	output \g133868/_0_  ;
	output \g133869/_0_  ;
	output \g133871/_0_  ;
	output \g133872/_0_  ;
	output \g133873/_0_  ;
	output \g133874/_0_  ;
	output \g133875/_0_  ;
	output \g133876/_0_  ;
	output \g133877/_0_  ;
	output \g133878/_0_  ;
	output \g133879/_0_  ;
	output \g133881/_0_  ;
	output \g133882/_0_  ;
	output \g133883/_0_  ;
	output \g133884/_0_  ;
	output \g133885/_0_  ;
	output \g133886/_0_  ;
	output \g133887/_0_  ;
	output \g133888/_0_  ;
	output \g133889/_0_  ;
	output \g133890/_0_  ;
	output \g133891/_0_  ;
	output \g133892/_0_  ;
	output \g133893/_0_  ;
	output \g133894/_0_  ;
	output \g133895/_0_  ;
	output \g133896/_0_  ;
	output \g133897/_0_  ;
	output \g133898/_0_  ;
	output \g133910/_0_  ;
	output \g133911/_0_  ;
	output \g133912/_0_  ;
	output \g133915/_0_  ;
	output \g133917/_0_  ;
	output \g133929/_0_  ;
	output \g134014/_0_  ;
	output \g134040/_0_  ;
	output \g134041/_0_  ;
	output \g134042/_0_  ;
	output \g134043/_0_  ;
	output \g134044/_0_  ;
	output \g134045/_0_  ;
	output \g134046/_0_  ;
	output \g134047/_0_  ;
	output \g134048/_0_  ;
	output \g134049/_0_  ;
	output \g134050/_0_  ;
	output \g134051/_0_  ;
	output \g134052/_0_  ;
	output \g134053/_0_  ;
	output \g134054/_0_  ;
	output \g134056/_0_  ;
	output \g134059/_0_  ;
	output \g134064/_0_  ;
	output \g134067/_0_  ;
	output \g134068/_0_  ;
	output \g134069/_0_  ;
	output \g134070/_0_  ;
	output \g134071/_0_  ;
	output \g134073/_0_  ;
	output \g134076/_0_  ;
	output \g134131/_0_  ;
	output \g134132/_0_  ;
	output \g134156/_0_  ;
	output \g134157/_0_  ;
	output \g134158/_0_  ;
	output \g134159/_0_  ;
	output \g134163/_0_  ;
	output \g134164/_0_  ;
	output \g134165/_0_  ;
	output \g134166/_0_  ;
	output \g134167/_0_  ;
	output \g134168/_0_  ;
	output \g134169/_0_  ;
	output \g134170/_0_  ;
	output \g134171/_0_  ;
	output \g134172/_0_  ;
	output \g134173/_0_  ;
	output \g134174/_0_  ;
	output \g134176/_0_  ;
	output \g134177/_0_  ;
	output \g134178/_0_  ;
	output \g134179/_0_  ;
	output \g134181/_0_  ;
	output \g134183/_0_  ;
	output \g134184/_0_  ;
	output \g134185/_0_  ;
	output \g134186/_0_  ;
	output \g134187/_0_  ;
	output \g134188/_0_  ;
	output \g134189/_0_  ;
	output \g134190/_0_  ;
	output \g134191/_0_  ;
	output \g134194/_0_  ;
	output \g134202/_0_  ;
	output \g134207/_0_  ;
	output \g134214/_0_  ;
	output \g134216/_0_  ;
	output \g134226/_0_  ;
	output \g134228/_0_  ;
	output \g134360/_0_  ;
	output \g134383/_0_  ;
	output \g134412/_0_  ;
	output \g134413/_0_  ;
	output \g134419/_0_  ;
	output \g134420/_0_  ;
	output \g134421/_0_  ;
	output \g134422/_0_  ;
	output \g134423/_0_  ;
	output \g134424/_0_  ;
	output \g134426/_0_  ;
	output \g134429/_0_  ;
	output \g134431/_0_  ;
	output \g134433/_0_  ;
	output \g134434/_0_  ;
	output \g134435/_0_  ;
	output \g134436/_0_  ;
	output \g134438/_0_  ;
	output \g134439/_0_  ;
	output \g134441/_0_  ;
	output \g134442/_0_  ;
	output \g134443/_0_  ;
	output \g134445/_0_  ;
	output \g134446/_0_  ;
	output \g134447/_0_  ;
	output \g134448/_0_  ;
	output \g134449/_0_  ;
	output \g134450/_0_  ;
	output \g134451/_0_  ;
	output \g134453/_0_  ;
	output \g134454/_0_  ;
	output \g134455/_0_  ;
	output \g134457/_0_  ;
	output \g134458/_0_  ;
	output \g134459/_0_  ;
	output \g134460/_0_  ;
	output \g134469/_0_  ;
	output \g134470/_0_  ;
	output \g134471/_0_  ;
	output \g134472/_0_  ;
	output \g134479/_0_  ;
	output \g134480/_0_  ;
	output \g134481/_0_  ;
	output \g134482/_0_  ;
	output \g134490/_0_  ;
	output \g134491/_0_  ;
	output \g134496/_0_  ;
	output \g134506/_0_  ;
	output \g134508/_0_  ;
	output \g134579/_0_  ;
	output \g134603/_0_  ;
	output \g134604/_0_  ;
	output \g134605/_0_  ;
	output \g134606/_0_  ;
	output \g134607/_0_  ;
	output \g134608/_0_  ;
	output \g134609/_0_  ;
	output \g134610/_0_  ;
	output \g134611/_0_  ;
	output \g134612/_0_  ;
	output \g134613/_0_  ;
	output \g134614/_0_  ;
	output \g134615/_0_  ;
	output \g134616/_0_  ;
	output \g134617/_0_  ;
	output \g134618/_0_  ;
	output \g134619/_0_  ;
	output \g134620/_0_  ;
	output \g134621/_0_  ;
	output \g134632/_0_  ;
	output \g134633/_0_  ;
	output \g134636/_0_  ;
	output \g134637/_0_  ;
	output \g134638/_0_  ;
	output \g134639/_0_  ;
	output \g134645/_0_  ;
	output \g134646/_0_  ;
	output \g134648/_0_  ;
	output \g134649/_0_  ;
	output \g134650/_0_  ;
	output \g134651/_0_  ;
	output \g134652/_0_  ;
	output \g134656/_0_  ;
	output \g134657/_0_  ;
	output \g134658/_0_  ;
	output \g134664/_0_  ;
	output \g134665/_0_  ;
	output \g134671/_0_  ;
	output \g134672/_0_  ;
	output \g134686/_0_  ;
	output \g134687/_0_  ;
	output \g134735/_0_  ;
	output \g134908/_0_  ;
	output \g134909/_0_  ;
	output \g134910/_0_  ;
	output \g134920/_0_  ;
	output \g134921/_0_  ;
	output \g134922/_0_  ;
	output \g134923/_0_  ;
	output \g134925/_0_  ;
	output \g134926/_0_  ;
	output \g134928/_0_  ;
	output \g134929/_0_  ;
	output \g134933/_0_  ;
	output \g134934/_0_  ;
	output \g134935/_0_  ;
	output \g134936/_0_  ;
	output \g134937/_0_  ;
	output \g134938/_0_  ;
	output \g134940/_0_  ;
	output \g134941/_0_  ;
	output \g134943/_0_  ;
	output \g134945/_0_  ;
	output \g134946/_0_  ;
	output \g134947/_0_  ;
	output \g134948/_0_  ;
	output \g134949/_0_  ;
	output \g134950/_0_  ;
	output \g134959/_0_  ;
	output \g134960/_0_  ;
	output \g134961/_0_  ;
	output \g134979/_0_  ;
	output \g134980/_0_  ;
	output \g135054/_0_  ;
	output \g135061/_0_  ;
	output \g135072/_0_  ;
	output \g135100/_0_  ;
	output \g135127/_0_  ;
	output \g135128/_0_  ;
	output \g135129/_0_  ;
	output \g135130/_0_  ;
	output \g135132/_0_  ;
	output \g135133/_0_  ;
	output \g135134/_0_  ;
	output \g135135/_0_  ;
	output \g135136/_0_  ;
	output \g135137/_0_  ;
	output \g135138/_0_  ;
	output \g135139/_0_  ;
	output \g135140/_0_  ;
	output \g135141/_0_  ;
	output \g135142/_0_  ;
	output \g135145/_0_  ;
	output \g135146/_0_  ;
	output \g135151/_0_  ;
	output \g135154/_0_  ;
	output \g135155/_0_  ;
	output \g135158/_0_  ;
	output \g135163/_0_  ;
	output \g135164/_0_  ;
	output \g135165/_0_  ;
	output \g135192/_0_  ;
	output \g135197/_0_  ;
	output \g135217/_0_  ;
	output \g135225/_0_  ;
	output \g135231/_0_  ;
	output \g135272/_0_  ;
	output \g135290/_0_  ;
	output \g135291/_0_  ;
	output \g135293/_0_  ;
	output \g135294/_0_  ;
	output \g135295/_0_  ;
	output \g135296/_0_  ;
	output \g135297/_0_  ;
	output \g135412/_0_  ;
	output \g135437/_0_  ;
	output \g135438/_0_  ;
	output \g135443/_0_  ;
	output \g135444/_0_  ;
	output \g135445/_0_  ;
	output \g135446/_0_  ;
	output \g135447/_0_  ;
	output \g135448/_0_  ;
	output \g135449/_0_  ;
	output \g135450/_0_  ;
	output \g135451/_0_  ;
	output \g135452/_0_  ;
	output \g135454/_0_  ;
	output \g135455/_0_  ;
	output \g135456/_0_  ;
	output \g135457/_0_  ;
	output \g135458/_0_  ;
	output \g135463/_0_  ;
	output \g135466/_0_  ;
	output \g135473/_0_  ;
	output \g135481/_0_  ;
	output \g135497/_0_  ;
	output \g135503/_0_  ;
	output \g135505/_0_  ;
	output \g135506/_0_  ;
	output \g135557/_0_  ;
	output \g135558/_0_  ;
	output \g135569/_0_  ;
	output \g135570/_0_  ;
	output \g135571/_0_  ;
	output \g135572/_0_  ;
	output \g135573/_0_  ;
	output \g135575/_0_  ;
	output \g135578/_0_  ;
	output \g135754/_0_  ;
	output \g135755/_0_  ;
	output \g135756/_0_  ;
	output \g135767/_0_  ;
	output \g135768/_0_  ;
	output \g135769/_0_  ;
	output \g135777/_0_  ;
	output \g135778/_0_  ;
	output \g135779/_0_  ;
	output \g135872/_0_  ;
	output \g135873/_0_  ;
	output \g135875/_0_  ;
	output \g135877/_0_  ;
	output \g135878/_0_  ;
	output \g135879/_0_  ;
	output \g135880/_0_  ;
	output \g136087/_0_  ;
	output \g136118/_0_  ;
	output \g136119/_0_  ;
	output \g136120/_0_  ;
	output \g136121/_0_  ;
	output \g136122/_0_  ;
	output \g136123/_0_  ;
	output \g136124/_0_  ;
	output \g136125/_0_  ;
	output \g136126/_0_  ;
	output \g136127/_0_  ;
	output \g136128/_0_  ;
	output \g136129/_0_  ;
	output \g136130/_0_  ;
	output \g136131/_0_  ;
	output \g136132/_0_  ;
	output \g136133/_0_  ;
	output \g136172/_0_  ;
	output \g136173/_0_  ;
	output \g136174/_0_  ;
	output \g136175/_0_  ;
	output \g136177/_0_  ;
	output \g136178/_0_  ;
	output \g136242/_0_  ;
	output \g136243/_0_  ;
	output \g136244/_0_  ;
	output \g136246/_0_  ;
	output \g136248/_0_  ;
	output \g136249/_0_  ;
	output \g136250/_0_  ;
	output \g136251/_0_  ;
	output \g136252/_0_  ;
	output \g136253/_0_  ;
	output \g136254/_0_  ;
	output \g136255/_0_  ;
	output \g136256/_0_  ;
	output \g136257/_0_  ;
	output \g136258/_0_  ;
	output \g136259/_0_  ;
	output \g136260/_0_  ;
	output \g136261/_0_  ;
	output \g136262/_0_  ;
	output \g136263/_0_  ;
	output \g136264/_0_  ;
	output \g136265/_0_  ;
	output \g136266/_0_  ;
	output \g136267/_0_  ;
	output \g136268/_0_  ;
	output \g136269/_0_  ;
	output \g136270/_0_  ;
	output \g136271/_0_  ;
	output \g136272/_0_  ;
	output \g136273/_0_  ;
	output \g136274/_0_  ;
	output \g136275/_0_  ;
	output \g136276/_0_  ;
	output \g136277/_0_  ;
	output \g136279/_0_  ;
	output \g136280/_0_  ;
	output \g136281/_0_  ;
	output \g136282/_0_  ;
	output \g136283/_0_  ;
	output \g136285/_0_  ;
	output \g136286/_0_  ;
	output \g136287/_0_  ;
	output \g136288/_0_  ;
	output \g136289/_0_  ;
	output \g136290/_0_  ;
	output \g136291/_0_  ;
	output \g136292/_0_  ;
	output \g136293/_0_  ;
	output \g136295/_0_  ;
	output \g136467/_0_  ;
	output \g136468/_0_  ;
	output \g136469/_0_  ;
	output \g136470/_0_  ;
	output \g136472/_0_  ;
	output \g136473/_0_  ;
	output \g136474/_0_  ;
	output \g136476/_0_  ;
	output \g136479/_0_  ;
	output \g136480/_0_  ;
	output \g136481/_0_  ;
	output \g136482/_0_  ;
	output \g136483/_0_  ;
	output \g136484/_0_  ;
	output \g136485/_0_  ;
	output \g136486/_0_  ;
	output \g136528/_0_  ;
	output \g136529/_0_  ;
	output \g136530/_0_  ;
	output \g136531/_0_  ;
	output \g136532/_0_  ;
	output \g136533/_0_  ;
	output \g136534/_0_  ;
	output \g136535/_0_  ;
	output \g136536/_0_  ;
	output \g136537/_0_  ;
	output \g136538/_0_  ;
	output \g136539/_0_  ;
	output \g136540/_0_  ;
	output \g136541/_0_  ;
	output \g136542/_0_  ;
	output \g136543/_0_  ;
	output \g136544/_0_  ;
	output \g136545/_0_  ;
	output \g136546/_0_  ;
	output \g136547/_0_  ;
	output \g136548/_0_  ;
	output \g136549/_0_  ;
	output \g136550/_0_  ;
	output \g136551/_0_  ;
	output \g136552/_0_  ;
	output \g136553/_0_  ;
	output \g136554/_0_  ;
	output \g136555/_0_  ;
	output \g136556/_0_  ;
	output \g136557/_0_  ;
	output \g136558/_0_  ;
	output \g136559/_0_  ;
	output \g136560/_0_  ;
	output \g136561/_0_  ;
	output \g136562/_0_  ;
	output \g136563/_0_  ;
	output \g136564/_0_  ;
	output \g136565/_0_  ;
	output \g136566/_0_  ;
	output \g136567/_0_  ;
	output \g136568/_0_  ;
	output \g136570/_0_  ;
	output \g136571/_0_  ;
	output \g136572/_0_  ;
	output \g136573/_0_  ;
	output \g136574/_0_  ;
	output \g136575/_0_  ;
	output \g136576/_0_  ;
	output \g136577/_0_  ;
	output \g136578/_0_  ;
	output \g136579/_0_  ;
	output \g136580/_0_  ;
	output \g136582/_0_  ;
	output \g136583/_0_  ;
	output \g136584/_0_  ;
	output \g136585/_0_  ;
	output \g136586/_0_  ;
	output \g136587/_0_  ;
	output \g136588/_0_  ;
	output \g136589/_0_  ;
	output \g136590/_0_  ;
	output \g136591/_0_  ;
	output \g136592/_0_  ;
	output \g136593/_0_  ;
	output \g136594/_0_  ;
	output \g136595/_0_  ;
	output \g136596/_0_  ;
	output \g136597/_0_  ;
	output \g136598/_0_  ;
	output \g136599/_0_  ;
	output \g136600/_0_  ;
	output \g136601/_0_  ;
	output \g136602/_0_  ;
	output \g136603/_0_  ;
	output \g136604/_0_  ;
	output \g136605/_0_  ;
	output \g136606/_0_  ;
	output \g136607/_0_  ;
	output \g136609/_0_  ;
	output \g136610/_0_  ;
	output \g136611/_0_  ;
	output \g136616/_0_  ;
	output \g136617/_0_  ;
	output \g136618/_0_  ;
	output \g136619/_0_  ;
	output \g136626/_0_  ;
	output \g136628/_0_  ;
	output \g136646/_0_  ;
	output \g136649/_0_  ;
	output \g136662/_0_  ;
	output \g136666/_0_  ;
	output \g136695/_0_  ;
	output \g136696/_0_  ;
	output \g136699/_0_  ;
	output \g136762/_0_  ;
	output \g136763/_0_  ;
	output \g136764/_0_  ;
	output \g136765/_0_  ;
	output \g136768/_0_  ;
	output \g136769/_0_  ;
	output \g137051/_0_  ;
	output \g137052/_0_  ;
	output \g137053/_0_  ;
	output \g137054/_0_  ;
	output \g137055/_0_  ;
	output \g137056/_0_  ;
	output \g137057/_0_  ;
	output \g137060/_0_  ;
	output \g137061/_0_  ;
	output \g137063/_0_  ;
	output \g137064/_0_  ;
	output \g137065/_0_  ;
	output \g137067/_0_  ;
	output \g137069/_0_  ;
	output \g137072/_0_  ;
	output \g137073/_0_  ;
	output \g137075/_0_  ;
	output \g137111/_0_  ;
	output \g137122/_0_  ;
	output \g137133/_0_  ;
	output \g137134/_0_  ;
	output \g137135/_0_  ;
	output \g137136/_0_  ;
	output \g137137/_0_  ;
	output \g137138/_0_  ;
	output \g137144/_0_  ;
	output \g137145/_0_  ;
	output \g137146/_0_  ;
	output \g137149/_0_  ;
	output \g137234/_0_  ;
	output \g137237/_0_  ;
	output \g137238/_0_  ;
	output \g137294/_0_  ;
	output \g137295/_0_  ;
	output \g137296/_0_  ;
	output \g137297/_0_  ;
	output \g137298/_0_  ;
	output \g137299/_0_  ;
	output \g137300/_0_  ;
	output \g137301/_0_  ;
	output \g137302/_0_  ;
	output \g137303/_0_  ;
	output \g137304/_0_  ;
	output \g137305/_0_  ;
	output \g137306/_0_  ;
	output \g137307/_0_  ;
	output \g137308/_0_  ;
	output \g137309/_0_  ;
	output \g137310/_0_  ;
	output \g137311/_0_  ;
	output \g137312/_0_  ;
	output \g137313/_0_  ;
	output \g137314/_0_  ;
	output \g137315/_0_  ;
	output \g137316/_0_  ;
	output \g137317/_0_  ;
	output \g137318/_0_  ;
	output \g137319/_0_  ;
	output \g137320/_0_  ;
	output \g137321/_0_  ;
	output \g137322/_0_  ;
	output \g137323/_0_  ;
	output \g137324/_0_  ;
	output \g137325/_0_  ;
	output \g137327/_0_  ;
	output \g137328/_0_  ;
	output \g137329/_0_  ;
	output \g137330/_0_  ;
	output \g137331/_0_  ;
	output \g137332/_0_  ;
	output \g137333/_0_  ;
	output \g137334/_0_  ;
	output \g137335/_0_  ;
	output \g137336/_0_  ;
	output \g137337/_0_  ;
	output \g137338/_0_  ;
	output \g137339/_0_  ;
	output \g137340/_0_  ;
	output \g137341/_0_  ;
	output \g137342/_0_  ;
	output \g137343/_0_  ;
	output \g137344/_0_  ;
	output \g137345/_0_  ;
	output \g137346/_0_  ;
	output \g137347/_0_  ;
	output \g137349/_0_  ;
	output \g137350/_0_  ;
	output \g137351/_0_  ;
	output \g137352/_0_  ;
	output \g137353/_0_  ;
	output \g137354/_0_  ;
	output \g137448/_0_  ;
	output \g137483/_0_  ;
	output \g137484/_0_  ;
	output \g137485/_0_  ;
	output \g137486/_0_  ;
	output \g137487/_0_  ;
	output \g137488/_0_  ;
	output \g137491/_0_  ;
	output \g137492/_0_  ;
	output \g137493/_0_  ;
	output \g137494/_0_  ;
	output \g137495/_0_  ;
	output \g137496/_0_  ;
	output \g137497/_0_  ;
	output \g137499/_0_  ;
	output \g137501/_0_  ;
	output \g137502/_0_  ;
	output \g137503/_0_  ;
	output \g137504/_0_  ;
	output \g137505/_0_  ;
	output \g137506/_0_  ;
	output \g137507/_0_  ;
	output \g137508/_0_  ;
	output \g137509/_0_  ;
	output \g137511/_0_  ;
	output \g137512/_0_  ;
	output \g137513/_0_  ;
	output \g137514/_0_  ;
	output \g137515/_0_  ;
	output \g137516/_0_  ;
	output \g137517/_0_  ;
	output \g137519/_0_  ;
	output \g137520/_0_  ;
	output \g137521/_0_  ;
	output \g137524/_0_  ;
	output \g137541/_0_  ;
	output \g137547/_0_  ;
	output \g137554/_0_  ;
	output \g137559/_0_  ;
	output \g137566/_0_  ;
	output \g137571/_0_  ;
	output \g137778/_0_  ;
	output \g137782/_0_  ;
	output \g137783/_0_  ;
	output \g137784/_0_  ;
	output \g137785/_0_  ;
	output \g137786/_0_  ;
	output \g137820/_0_  ;
	output \g137821/_0_  ;
	output \g137822/_0_  ;
	output \g137823/_0_  ;
	output \g137824/_0_  ;
	output \g137825/_0_  ;
	output \g137826/_0_  ;
	output \g137827/_0_  ;
	output \g137828/_0_  ;
	output \g137829/_0_  ;
	output \g137830/_0_  ;
	output \g137831/_0_  ;
	output \g137832/_0_  ;
	output \g137833/_0_  ;
	output \g137834/_0_  ;
	output \g137835/_0_  ;
	output \g137836/_0_  ;
	output \g137837/_0_  ;
	output \g137838/_0_  ;
	output \g137839/_0_  ;
	output \g137840/_0_  ;
	output \g137841/_0_  ;
	output \g137842/_0_  ;
	output \g137843/_0_  ;
	output \g137844/_0_  ;
	output \g137845/_0_  ;
	output \g137846/_0_  ;
	output \g137847/_0_  ;
	output \g137848/_0_  ;
	output \g137849/_0_  ;
	output \g137850/_0_  ;
	output \g137851/_0_  ;
	output \g137852/_0_  ;
	output \g137853/_0_  ;
	output \g137854/_0_  ;
	output \g137855/_0_  ;
	output \g137856/_0_  ;
	output \g137857/_0_  ;
	output \g137858/_0_  ;
	output \g137859/_0_  ;
	output \g137860/_0_  ;
	output \g137861/_0_  ;
	output \g137862/_0_  ;
	output \g137863/_0_  ;
	output \g137864/_0_  ;
	output \g137865/_0_  ;
	output \g137866/_0_  ;
	output \g137867/_0_  ;
	output \g137868/_0_  ;
	output \g137869/_0_  ;
	output \g137870/_0_  ;
	output \g137871/_0_  ;
	output \g137872/_0_  ;
	output \g137873/_0_  ;
	output \g137874/_0_  ;
	output \g137875/_0_  ;
	output \g137876/_0_  ;
	output \g137877/_0_  ;
	output \g137878/_0_  ;
	output \g137879/_0_  ;
	output \g137880/_0_  ;
	output \g137881/_0_  ;
	output \g137882/_0_  ;
	output \g137883/_0_  ;
	output \g137884/_0_  ;
	output \g137885/_0_  ;
	output \g137886/_0_  ;
	output \g137887/_0_  ;
	output \g137888/_0_  ;
	output \g137889/_0_  ;
	output \g137890/_0_  ;
	output \g137891/_0_  ;
	output \g137892/_0_  ;
	output \g137893/_0_  ;
	output \g137894/_0_  ;
	output \g137895/_0_  ;
	output \g137896/_0_  ;
	output \g137897/_0_  ;
	output \g137898/_0_  ;
	output \g137899/_0_  ;
	output \g137900/_0_  ;
	output \g137901/_0_  ;
	output \g137902/_0_  ;
	output \g137903/_0_  ;
	output \g138338/_0_  ;
	output \g138340/_0_  ;
	output \g138341/_0_  ;
	output \g138346/_0_  ;
	output \g138347/_0_  ;
	output \g138375/_0_  ;
	output \g138395/_0_  ;
	output \g138396/_0_  ;
	output \g138397/_0_  ;
	output \g138398/_0_  ;
	output \g138400/_0_  ;
	output \g138401/_0_  ;
	output \g138402/_0_  ;
	output \g138403/_0_  ;
	output \g138404/_0_  ;
	output \g138405/_0_  ;
	output \g138406/_0_  ;
	output \g138407/_0_  ;
	output \g138408/_0_  ;
	output \g138409/_0_  ;
	output \g138410/_0_  ;
	output \g138411/_0_  ;
	output \g138412/_0_  ;
	output \g138419/_0_  ;
	output \g138420/_0_  ;
	output \g138421/_0_  ;
	output \g138422/_0_  ;
	output \g138423/_0_  ;
	output \g138424/_0_  ;
	output \g138425/_0_  ;
	output \g138426/_0_  ;
	output \g138427/_0_  ;
	output \g138428/_0_  ;
	output \g138429/_0_  ;
	output \g138430/_0_  ;
	output \g138431/_0_  ;
	output \g138432/_0_  ;
	output \g138433/_0_  ;
	output \g138434/_0_  ;
	output \g138435/_0_  ;
	output \g138436/_0_  ;
	output \g138437/_0_  ;
	output \g138438/_0_  ;
	output \g138439/_0_  ;
	output \g138440/_0_  ;
	output \g138441/_0_  ;
	output \g138442/_0_  ;
	output \g138443/_0_  ;
	output \g138908/_0_  ;
	output \g138909/_0_  ;
	output \g138910/_0_  ;
	output \g138914/_0_  ;
	output \g138915/_0_  ;
	output \g138917/_0_  ;
	output \g138918/_0_  ;
	output \g138919/_0_  ;
	output \g138920/_0_  ;
	output \g138921/_0_  ;
	output \g138925/_0_  ;
	output \g138926/_0_  ;
	output \g138927/_0_  ;
	output \g138930/_0_  ;
	output \g138931/_0_  ;
	output \g138932/_0_  ;
	output \g138960/_0_  ;
	output \g138962/_0_  ;
	output \g139037/_0_  ;
	output \g139038/_0_  ;
	output \g139040/_0_  ;
	output \g139043/_0_  ;
	output \g139044/_0_  ;
	output \g139045/_0_  ;
	output \g139046/_0_  ;
	output \g139047/_0_  ;
	output \g139048/_0_  ;
	output \g139049/_0_  ;
	output \g139050/_0_  ;
	output \g139051/_0_  ;
	output \g139053/_0_  ;
	output \g139054/_0_  ;
	output \g139055/_0_  ;
	output \g139056/_0_  ;
	output \g139057/_0_  ;
	output \g139058/_0_  ;
	output \g139059/_0_  ;
	output \g139060/_0_  ;
	output \g139062/_0_  ;
	output \g139063/_0_  ;
	output \g139064/_0_  ;
	output \g139099/_0_  ;
	output \g139126/_0_  ;
	output \g139127/_0_  ;
	output \g139128/_0_  ;
	output \g139129/_0_  ;
	output \g139130/_0_  ;
	output \g139131/_0_  ;
	output \g139132/_0_  ;
	output \g139133/_0_  ;
	output \g139134/_0_  ;
	output \g139135/_0_  ;
	output \g139136/_0_  ;
	output \g139137/_0_  ;
	output \g139138/_0_  ;
	output \g139139/_0_  ;
	output \g139140/_0_  ;
	output \g139141/_0_  ;
	output \g139260/_0_  ;
	output \g139263/_0_  ;
	output \g139267/_0_  ;
	output \g139270/_0_  ;
	output \g139273/_0_  ;
	output \g139276/_0_  ;
	output \g139279/_0_  ;
	output \g139283/_0_  ;
	output \g139286/_0_  ;
	output \g139289/_0_  ;
	output \g139292/_0_  ;
	output \g139295/_0_  ;
	output \g139298/_0_  ;
	output \g139302/_0_  ;
	output \g139305/_0_  ;
	output \g139309/_0_  ;
	output \g139871/_0_  ;
	output \g139872/_0_  ;
	output \g139873/_0_  ;
	output \g139874/_0_  ;
	output \g139875/_0_  ;
	output \g139876/_0_  ;
	output \g139877/_0_  ;
	output \g139878/_0_  ;
	output \g139879/_0_  ;
	output \g139880/_0_  ;
	output \g139881/_0_  ;
	output \g139882/_0_  ;
	output \g139883/_0_  ;
	output \g139884/_0_  ;
	output \g139885/_0_  ;
	output \g139886/_0_  ;
	output \g139887/_0_  ;
	output \g139888/_0_  ;
	output \g139889/_0_  ;
	output \g139890/_0_  ;
	output \g139891/_0_  ;
	output \g139892/_0_  ;
	output \g139893/_0_  ;
	output \g139895/_0_  ;
	output \g139896/_0_  ;
	output \g139899/_0_  ;
	output \g139901/_0_  ;
	output \g139902/_0_  ;
	output \g139903/_0_  ;
	output \g139904/_0_  ;
	output \g140285/_0_  ;
	output \g140288/_0_  ;
	output \g140329/_0_  ;
	output \g140774/_0_  ;
	output \g140832/_0_  ;
	output \g140834/_0_  ;
	output \g140836/_0_  ;
	output \g140838/_0_  ;
	output \g140840/_0_  ;
	output \g140842/_0_  ;
	output \g140844/_0_  ;
	output \g140846/_0_  ;
	output \g140847/_0_  ;
	output \g140848/_0_  ;
	output \g140850/_0_  ;
	output \g140851/_0_  ;
	output \g140852/_0_  ;
	output \g140853/_0_  ;
	output \g140855/_0_  ;
	output \g140857/_0_  ;
	output \g140861/_0_  ;
	output \g140923/_0_  ;
	output \g141178/_0_  ;
	output \g141179/_0_  ;
	output \g141180/_0_  ;
	output \g141480/_0_  ;
	output \g141495/_0_  ;
	output \g141497/_0_  ;
	output \g141562/_0_  ;
	output \g141563/_0_  ;
	output \g141564/_0_  ;
	output \g141589/_0_  ;
	output \g141617/_0_  ;
	output \g141618/_0_  ;
	output \g141621/_0_  ;
	output \g141625/_0_  ;
	output \g141626/_0_  ;
	output \g141630/_0_  ;
	output \g141634/_0_  ;
	output \g141638/_0_  ;
	output \g141642/_0_  ;
	output \g141646/_0_  ;
	output \g141649/_0_  ;
	output \g141651/_0_  ;
	output \g141652/_0_  ;
	output \g141655/_0_  ;
	output \g141658/_0_  ;
	output \g141661/_0_  ;
	output \g141663/_0_  ;
	output \g141664/_0_  ;
	output \g141667/_0_  ;
	output \g141671/_0_  ;
	output \g141706/_0_  ;
	output \g141976/_0_  ;
	output \g141977/_0_  ;
	output \g141994/_0_  ;
	output \g142246/_0_  ;
	output \g142247/_0_  ;
	output \g142253/_0_  ;
	output \g142689/_0_  ;
	output \g142693/_0_  ;
	output \g142701/_0_  ;
	output \g142704/_0_  ;
	output \g142707/_0_  ;
	output \g142710/_0_  ;
	output \g142713/_0_  ;
	output \g142714/_0_  ;
	output \g142717/_0_  ;
	output \g142720/_0_  ;
	output \g142723/_0_  ;
	output \g142727/_0_  ;
	output \g142734/_0_  ;
	output \g143080/_0_  ;
	output \g143081/_0_  ;
	output \g143083/_0_  ;
	output \g143149/_0_  ;
	output \g143150/_0_  ;
	output \g143153/_0_  ;
	output \g143752/_0_  ;
	output \g143753/_0_  ;
	output \g143759/_0_  ;
	output \g144242/_0_  ;
	output \g144243/_0_  ;
	output \g144244/_0_  ;
	output \g144245/_0_  ;
	output \g144246/_0_  ;
	output \g144249/_0_  ;
	output \g145699/_0_  ;
	output \g145700/_0_  ;
	output \g145702/_0_  ;
	output \g145756/_0_  ;
	output \g145757/_0_  ;
	output \g145758/_0_  ;
	output \g146850/_0_  ;
	output \g146851/_0_  ;
	output \g146864/_0_  ;
	output \g147277/_0_  ;
	output \g147278/_0_  ;
	output \g147279/_0_  ;
	output \g147304/_0_  ;
	output \g147305/_0_  ;
	output \g147306/_0_  ;
	output \g147338/_3_  ;
	output \g147339/_3_  ;
	output \g147340/_3_  ;
	output \g147341/_3_  ;
	output \g147342/_3_  ;
	output \g147343/_3_  ;
	output \g147344/_3_  ;
	output \g147345/_3_  ;
	output \g147346/_3_  ;
	output \g147347/_3_  ;
	output \g147348/_3_  ;
	output \g147349/_3_  ;
	output \g147350/_3_  ;
	output \g147351/_3_  ;
	output \g147352/_3_  ;
	output \g147353/_3_  ;
	output \g147354/_3_  ;
	output \g147355/_3_  ;
	output \g147356/_3_  ;
	output \g147357/_3_  ;
	output \g147358/_3_  ;
	output \g147359/_3_  ;
	output \g147360/_3_  ;
	output \g147362/_3_  ;
	output \g147363/_3_  ;
	output \g147364/_3_  ;
	output \g147365/_3_  ;
	output \g147366/_3_  ;
	output \g147367/_3_  ;
	output \g147368/_3_  ;
	output \g147369/_3_  ;
	output \g148630/_0_  ;
	output \g148631/_0_  ;
	output \g148676/_0_  ;
	output \g148785/_0_  ;
	output \g148788/_0_  ;
	output \g148789/_0_  ;
	output \g148834/_0_  ;
	output \g148836/_0_  ;
	output \g148838/_0_  ;
	output \g149836/_0_  ;
	output \g149837/_0_  ;
	output \g149838/_0_  ;
	output \g150142/_0_  ;
	output \g152366/_0_  ;
	output \g152367/_0_  ;
	output \g152368/_0_  ;
	output \g152426/_0_  ;
	output \g152427/_0_  ;
	output \g152428/_0_  ;
	output \g152586/_0_  ;
	output \g152587/_0_  ;
	output \g152588/_0_  ;
	output \g153217/_0_  ;
	output \g154117/_0_  ;
	output \g154118/_0_  ;
	output \g154130/_0_  ;
	output \g154269/_0_  ;
	output \g154270/_0_  ;
	output \g154284/_0_  ;
	output \g154682/_0_  ;
	output \g155004/_0_  ;
	output \g155020/_0_  ;
	output \g155121/_0_  ;
	output \g155124/_0_  ;
	output \g155126/_0_  ;
	output \g155228/_0_  ;
	output \g155229/_0_  ;
	output \g155230/_0_  ;
	output \g155326/_0_  ;
	output \g155327/_0_  ;
	output \g155330/_0_  ;
	output \g155353/_0_  ;
	output \g155354/_0_  ;
	output \g155356/_0_  ;
	output \g155602/_0_  ;
	output \g155633/_0_  ;
	output \g155634/_0_  ;
	output \g155699/_0_  ;
	output \g155708/_0_  ;
	output \g155715/_0_  ;
	output \g156008/_0_  ;
	output \g156013/_0_  ;
	output \g156019/_0_  ;
	output \g156352/_0_  ;
	output \g156353/_0_  ;
	output \g156356/_0_  ;
	output \g156359/_0_  ;
	output \g156360/_0_  ;
	output \g156361/_0_  ;
	output \g156464/_0_  ;
	output \g156465/_0_  ;
	output \g156469/_0_  ;
	output \g156777/_0_  ;
	output \g156778/_0_  ;
	output \g156789/_0_  ;
	output \g158956/_0_  ;
	output \g158957/_0_  ;
	output \g158966/_0_  ;
	output \g159429/_1_  ;
	output \g159477/_1_  ;
	output \g159500/_1_  ;
	output \g159681/_0_  ;
	output \g159890/_0_  ;
	output \g159950/_0_  ;
	output \g160246/_0_  ;
	output \g160846/_0_  ;
	output \g160860/_0_  ;
	output \g160961/_0_  ;
	output \g160987/_0_  ;
	output \g161000/_0_  ;
	output \g161005/_0_  ;
	output \g161042/_0_  ;
	output \g161119/_0_  ;
	output \g161143/_0_  ;
	output \g161150/_0_  ;
	output \g161172/_0_  ;
	output \g161207/_0_  ;
	output \g161315/_0_  ;
	output \g161332/_0_  ;
	output \g161421/_0_  ;
	output \g161492/_0_  ;
	output \g161541/_0_  ;
	output \g161623/_0_  ;
	output \g161655/_0_  ;
	output \g161678/_0_  ;
	output \g161709/_0_  ;
	output \g161737/_0_  ;
	output \g161751/_0_  ;
	output \g161756/_0_  ;
	output \g162016/_0_  ;
	output \g162020/_0_  ;
	output \g162024/_0_  ;
	output \g163326/_0_  ;
	output \g163326/_3_  ;
	output \g174072/_1_  ;
	output \g174360/_1_  ;
	output \g174391/_0_  ;
	output \g180307/_0_  ;
	output \g180335/_0_  ;
	output \g180369/_0_  ;
	output \g180385/_0_  ;
	output \g180395/_0_  ;
	output \g180442/_0_  ;
	output \g180453/_0_  ;
	output \g180524/_0_  ;
	output \g180586/_0_  ;
	output \g180596/_0_  ;
	output \g180606/_0_  ;
	output \g180654/_0_  ;
	output \g180715/_0_  ;
	output \g180805/_0_  ;
	output \g180836/_0_  ;
	output \g180929/_0_  ;
	output \g180944/_0_  ;
	output \g180975/_0_  ;
	output \g181036/_0_  ;
	output \g181072/_0_  ;
	output \g181083/_0_  ;
	output \g181093/_0_  ;
	output \g181127/_0_  ;
	output \g181137/_0_  ;
	output \g181150/_0_  ;
	output \g181160/_0_  ;
	output \g181180/_0_  ;
	output \g181191/_0_  ;
	output \g181238/_0_  ;
	output \g181262/_0_  ;
	output \g181270/_0_  ;
	output \g181280/_0_  ;
	output \g181315/_0_  ;
	output \g181366/_0_  ;
	output \g181385/_0_  ;
	output \g181458/_0_  ;
	output \g181464/_0_  ;
	output \g181478/_0_  ;
	output \g181522/_0_  ;
	output \g181537/_0_  ;
	output \g181584/_0_  ;
	output \g181669/_0_  ;
	output \g181681/_0_  ;
	output \g181719/_0_  ;
	output \g181778/_0_  ;
	output \g181840/_0_  ;
	output \g181936/_0_  ;
	output \g181986/_0_  ;
	output \g182000/_0_  ;
	output \g182083/_0_  ;
	output \g182179/_0_  ;
	output \g182201/_0_  ;
	output \g182227/_0_  ;
	output \g182316/_0_  ;
	output \g182358/_0_  ;
	output \g182473/_0_  ;
	output \g182678/_0_  ;
	output \g53/_0_  ;
	wire _w17089_ ;
	wire _w17088_ ;
	wire _w17087_ ;
	wire _w17086_ ;
	wire _w17085_ ;
	wire _w17084_ ;
	wire _w17083_ ;
	wire _w17082_ ;
	wire _w17081_ ;
	wire _w17080_ ;
	wire _w17079_ ;
	wire _w17078_ ;
	wire _w17077_ ;
	wire _w17076_ ;
	wire _w17075_ ;
	wire _w17074_ ;
	wire _w17073_ ;
	wire _w17072_ ;
	wire _w17071_ ;
	wire _w17070_ ;
	wire _w17069_ ;
	wire _w17068_ ;
	wire _w17067_ ;
	wire _w17066_ ;
	wire _w17065_ ;
	wire _w17064_ ;
	wire _w17063_ ;
	wire _w17062_ ;
	wire _w17061_ ;
	wire _w17060_ ;
	wire _w17059_ ;
	wire _w17058_ ;
	wire _w17057_ ;
	wire _w17056_ ;
	wire _w17055_ ;
	wire _w17054_ ;
	wire _w17053_ ;
	wire _w17052_ ;
	wire _w17051_ ;
	wire _w17050_ ;
	wire _w17049_ ;
	wire _w17048_ ;
	wire _w17047_ ;
	wire _w17046_ ;
	wire _w17045_ ;
	wire _w17044_ ;
	wire _w17043_ ;
	wire _w17042_ ;
	wire _w17041_ ;
	wire _w17040_ ;
	wire _w17039_ ;
	wire _w17038_ ;
	wire _w17037_ ;
	wire _w17036_ ;
	wire _w17035_ ;
	wire _w17034_ ;
	wire _w17033_ ;
	wire _w17032_ ;
	wire _w17031_ ;
	wire _w17030_ ;
	wire _w17029_ ;
	wire _w17028_ ;
	wire _w17027_ ;
	wire _w17026_ ;
	wire _w17025_ ;
	wire _w17024_ ;
	wire _w17023_ ;
	wire _w17022_ ;
	wire _w17021_ ;
	wire _w17020_ ;
	wire _w17019_ ;
	wire _w17018_ ;
	wire _w17017_ ;
	wire _w17016_ ;
	wire _w17015_ ;
	wire _w17014_ ;
	wire _w17013_ ;
	wire _w17012_ ;
	wire _w17011_ ;
	wire _w17010_ ;
	wire _w17009_ ;
	wire _w17008_ ;
	wire _w17007_ ;
	wire _w17006_ ;
	wire _w17005_ ;
	wire _w17004_ ;
	wire _w17003_ ;
	wire _w17002_ ;
	wire _w17001_ ;
	wire _w17000_ ;
	wire _w16999_ ;
	wire _w16998_ ;
	wire _w16997_ ;
	wire _w16996_ ;
	wire _w16995_ ;
	wire _w16994_ ;
	wire _w16993_ ;
	wire _w16992_ ;
	wire _w16991_ ;
	wire _w16990_ ;
	wire _w16989_ ;
	wire _w16988_ ;
	wire _w16987_ ;
	wire _w16986_ ;
	wire _w16985_ ;
	wire _w16984_ ;
	wire _w16983_ ;
	wire _w16982_ ;
	wire _w16981_ ;
	wire _w16980_ ;
	wire _w16979_ ;
	wire _w16978_ ;
	wire _w16977_ ;
	wire _w16976_ ;
	wire _w16975_ ;
	wire _w16974_ ;
	wire _w16973_ ;
	wire _w16972_ ;
	wire _w16971_ ;
	wire _w16970_ ;
	wire _w16969_ ;
	wire _w16968_ ;
	wire _w16967_ ;
	wire _w16966_ ;
	wire _w16965_ ;
	wire _w16964_ ;
	wire _w16963_ ;
	wire _w16962_ ;
	wire _w16961_ ;
	wire _w16960_ ;
	wire _w16959_ ;
	wire _w16958_ ;
	wire _w16957_ ;
	wire _w16956_ ;
	wire _w16955_ ;
	wire _w16954_ ;
	wire _w16953_ ;
	wire _w16952_ ;
	wire _w16951_ ;
	wire _w16950_ ;
	wire _w16949_ ;
	wire _w16948_ ;
	wire _w16947_ ;
	wire _w16946_ ;
	wire _w16945_ ;
	wire _w16944_ ;
	wire _w16943_ ;
	wire _w16942_ ;
	wire _w16941_ ;
	wire _w16940_ ;
	wire _w16939_ ;
	wire _w16938_ ;
	wire _w16937_ ;
	wire _w16936_ ;
	wire _w16935_ ;
	wire _w16934_ ;
	wire _w16933_ ;
	wire _w16932_ ;
	wire _w16931_ ;
	wire _w16930_ ;
	wire _w16929_ ;
	wire _w16928_ ;
	wire _w16927_ ;
	wire _w16926_ ;
	wire _w16925_ ;
	wire _w16924_ ;
	wire _w16923_ ;
	wire _w16922_ ;
	wire _w16921_ ;
	wire _w16920_ ;
	wire _w16919_ ;
	wire _w16918_ ;
	wire _w16917_ ;
	wire _w16916_ ;
	wire _w16915_ ;
	wire _w16914_ ;
	wire _w16913_ ;
	wire _w16912_ ;
	wire _w16911_ ;
	wire _w16910_ ;
	wire _w16909_ ;
	wire _w16908_ ;
	wire _w16907_ ;
	wire _w16906_ ;
	wire _w16905_ ;
	wire _w16904_ ;
	wire _w16903_ ;
	wire _w16902_ ;
	wire _w16901_ ;
	wire _w16900_ ;
	wire _w16899_ ;
	wire _w16898_ ;
	wire _w16897_ ;
	wire _w16896_ ;
	wire _w16895_ ;
	wire _w16894_ ;
	wire _w16893_ ;
	wire _w16892_ ;
	wire _w16891_ ;
	wire _w16890_ ;
	wire _w16889_ ;
	wire _w16888_ ;
	wire _w16887_ ;
	wire _w16886_ ;
	wire _w16885_ ;
	wire _w16884_ ;
	wire _w16883_ ;
	wire _w16882_ ;
	wire _w16881_ ;
	wire _w16880_ ;
	wire _w16879_ ;
	wire _w16878_ ;
	wire _w16877_ ;
	wire _w16876_ ;
	wire _w16875_ ;
	wire _w16874_ ;
	wire _w16873_ ;
	wire _w16872_ ;
	wire _w16871_ ;
	wire _w16870_ ;
	wire _w16869_ ;
	wire _w16868_ ;
	wire _w16867_ ;
	wire _w16866_ ;
	wire _w16865_ ;
	wire _w16864_ ;
	wire _w16863_ ;
	wire _w16862_ ;
	wire _w16861_ ;
	wire _w16860_ ;
	wire _w16859_ ;
	wire _w16858_ ;
	wire _w16857_ ;
	wire _w16856_ ;
	wire _w16855_ ;
	wire _w16854_ ;
	wire _w16853_ ;
	wire _w16852_ ;
	wire _w16851_ ;
	wire _w16850_ ;
	wire _w16849_ ;
	wire _w16848_ ;
	wire _w16847_ ;
	wire _w16846_ ;
	wire _w16845_ ;
	wire _w16844_ ;
	wire _w16843_ ;
	wire _w16842_ ;
	wire _w16841_ ;
	wire _w16840_ ;
	wire _w16839_ ;
	wire _w16838_ ;
	wire _w16837_ ;
	wire _w16836_ ;
	wire _w16835_ ;
	wire _w16834_ ;
	wire _w16833_ ;
	wire _w16832_ ;
	wire _w16831_ ;
	wire _w16830_ ;
	wire _w16829_ ;
	wire _w16828_ ;
	wire _w16827_ ;
	wire _w16826_ ;
	wire _w16825_ ;
	wire _w16824_ ;
	wire _w16823_ ;
	wire _w16822_ ;
	wire _w16821_ ;
	wire _w16820_ ;
	wire _w16819_ ;
	wire _w16818_ ;
	wire _w16817_ ;
	wire _w16816_ ;
	wire _w16815_ ;
	wire _w16814_ ;
	wire _w16813_ ;
	wire _w16812_ ;
	wire _w16811_ ;
	wire _w16810_ ;
	wire _w16809_ ;
	wire _w16808_ ;
	wire _w16807_ ;
	wire _w16806_ ;
	wire _w16805_ ;
	wire _w16804_ ;
	wire _w16803_ ;
	wire _w16802_ ;
	wire _w16801_ ;
	wire _w16800_ ;
	wire _w16799_ ;
	wire _w16798_ ;
	wire _w16797_ ;
	wire _w16796_ ;
	wire _w16795_ ;
	wire _w16794_ ;
	wire _w16793_ ;
	wire _w16792_ ;
	wire _w16791_ ;
	wire _w16790_ ;
	wire _w16789_ ;
	wire _w16788_ ;
	wire _w16787_ ;
	wire _w16786_ ;
	wire _w16785_ ;
	wire _w16784_ ;
	wire _w16783_ ;
	wire _w16782_ ;
	wire _w16781_ ;
	wire _w16780_ ;
	wire _w16779_ ;
	wire _w16778_ ;
	wire _w16777_ ;
	wire _w16776_ ;
	wire _w16775_ ;
	wire _w16774_ ;
	wire _w16773_ ;
	wire _w16772_ ;
	wire _w16771_ ;
	wire _w16770_ ;
	wire _w16769_ ;
	wire _w16768_ ;
	wire _w16767_ ;
	wire _w16766_ ;
	wire _w16765_ ;
	wire _w16764_ ;
	wire _w16763_ ;
	wire _w16762_ ;
	wire _w16761_ ;
	wire _w16760_ ;
	wire _w16759_ ;
	wire _w16758_ ;
	wire _w16757_ ;
	wire _w16756_ ;
	wire _w16755_ ;
	wire _w16754_ ;
	wire _w16753_ ;
	wire _w16752_ ;
	wire _w16751_ ;
	wire _w16750_ ;
	wire _w16749_ ;
	wire _w16748_ ;
	wire _w16747_ ;
	wire _w16746_ ;
	wire _w16745_ ;
	wire _w16744_ ;
	wire _w16743_ ;
	wire _w16742_ ;
	wire _w16741_ ;
	wire _w16740_ ;
	wire _w16739_ ;
	wire _w16738_ ;
	wire _w16737_ ;
	wire _w16736_ ;
	wire _w16735_ ;
	wire _w16734_ ;
	wire _w16733_ ;
	wire _w16732_ ;
	wire _w16731_ ;
	wire _w16730_ ;
	wire _w16729_ ;
	wire _w16728_ ;
	wire _w16727_ ;
	wire _w16726_ ;
	wire _w16725_ ;
	wire _w16724_ ;
	wire _w16723_ ;
	wire _w16722_ ;
	wire _w16721_ ;
	wire _w16720_ ;
	wire _w16719_ ;
	wire _w16718_ ;
	wire _w16717_ ;
	wire _w16716_ ;
	wire _w16715_ ;
	wire _w16714_ ;
	wire _w16713_ ;
	wire _w16712_ ;
	wire _w16711_ ;
	wire _w16710_ ;
	wire _w16709_ ;
	wire _w16708_ ;
	wire _w16707_ ;
	wire _w16706_ ;
	wire _w16705_ ;
	wire _w16704_ ;
	wire _w16703_ ;
	wire _w16702_ ;
	wire _w16701_ ;
	wire _w16700_ ;
	wire _w16699_ ;
	wire _w16698_ ;
	wire _w16697_ ;
	wire _w16696_ ;
	wire _w16695_ ;
	wire _w16694_ ;
	wire _w16693_ ;
	wire _w16692_ ;
	wire _w16691_ ;
	wire _w16690_ ;
	wire _w16689_ ;
	wire _w16688_ ;
	wire _w16687_ ;
	wire _w16686_ ;
	wire _w16685_ ;
	wire _w16684_ ;
	wire _w16683_ ;
	wire _w16682_ ;
	wire _w16681_ ;
	wire _w16680_ ;
	wire _w16679_ ;
	wire _w16678_ ;
	wire _w16677_ ;
	wire _w16676_ ;
	wire _w16675_ ;
	wire _w16674_ ;
	wire _w16673_ ;
	wire _w16672_ ;
	wire _w16671_ ;
	wire _w16670_ ;
	wire _w16669_ ;
	wire _w16668_ ;
	wire _w16667_ ;
	wire _w16666_ ;
	wire _w16665_ ;
	wire _w16664_ ;
	wire _w16663_ ;
	wire _w16662_ ;
	wire _w16661_ ;
	wire _w16660_ ;
	wire _w16659_ ;
	wire _w16658_ ;
	wire _w16657_ ;
	wire _w16656_ ;
	wire _w16655_ ;
	wire _w16654_ ;
	wire _w16653_ ;
	wire _w16652_ ;
	wire _w16651_ ;
	wire _w16650_ ;
	wire _w16649_ ;
	wire _w16648_ ;
	wire _w16647_ ;
	wire _w16646_ ;
	wire _w16645_ ;
	wire _w16644_ ;
	wire _w16643_ ;
	wire _w16642_ ;
	wire _w16641_ ;
	wire _w16640_ ;
	wire _w16639_ ;
	wire _w16638_ ;
	wire _w16637_ ;
	wire _w16636_ ;
	wire _w16635_ ;
	wire _w16634_ ;
	wire _w16633_ ;
	wire _w16632_ ;
	wire _w16631_ ;
	wire _w16630_ ;
	wire _w16629_ ;
	wire _w16628_ ;
	wire _w16627_ ;
	wire _w16626_ ;
	wire _w16625_ ;
	wire _w16624_ ;
	wire _w16623_ ;
	wire _w16622_ ;
	wire _w16621_ ;
	wire _w16620_ ;
	wire _w16619_ ;
	wire _w16618_ ;
	wire _w16617_ ;
	wire _w16616_ ;
	wire _w16615_ ;
	wire _w16614_ ;
	wire _w16613_ ;
	wire _w16612_ ;
	wire _w16611_ ;
	wire _w16610_ ;
	wire _w16609_ ;
	wire _w16608_ ;
	wire _w16607_ ;
	wire _w16606_ ;
	wire _w16605_ ;
	wire _w16604_ ;
	wire _w16603_ ;
	wire _w16602_ ;
	wire _w16601_ ;
	wire _w16600_ ;
	wire _w16599_ ;
	wire _w16598_ ;
	wire _w16597_ ;
	wire _w16596_ ;
	wire _w16595_ ;
	wire _w16594_ ;
	wire _w16593_ ;
	wire _w16592_ ;
	wire _w16591_ ;
	wire _w16590_ ;
	wire _w16589_ ;
	wire _w16588_ ;
	wire _w16587_ ;
	wire _w16586_ ;
	wire _w16585_ ;
	wire _w16584_ ;
	wire _w16583_ ;
	wire _w16582_ ;
	wire _w16581_ ;
	wire _w16580_ ;
	wire _w16579_ ;
	wire _w16578_ ;
	wire _w16577_ ;
	wire _w16576_ ;
	wire _w16575_ ;
	wire _w16574_ ;
	wire _w16573_ ;
	wire _w16572_ ;
	wire _w16571_ ;
	wire _w16570_ ;
	wire _w16569_ ;
	wire _w16568_ ;
	wire _w16567_ ;
	wire _w16566_ ;
	wire _w16565_ ;
	wire _w16564_ ;
	wire _w16563_ ;
	wire _w16562_ ;
	wire _w16561_ ;
	wire _w16560_ ;
	wire _w16559_ ;
	wire _w16558_ ;
	wire _w16557_ ;
	wire _w16556_ ;
	wire _w16555_ ;
	wire _w16554_ ;
	wire _w16553_ ;
	wire _w16552_ ;
	wire _w16551_ ;
	wire _w16550_ ;
	wire _w16549_ ;
	wire _w16548_ ;
	wire _w16547_ ;
	wire _w16546_ ;
	wire _w16545_ ;
	wire _w16544_ ;
	wire _w16543_ ;
	wire _w16542_ ;
	wire _w16541_ ;
	wire _w16540_ ;
	wire _w16539_ ;
	wire _w16538_ ;
	wire _w16537_ ;
	wire _w16536_ ;
	wire _w16535_ ;
	wire _w16534_ ;
	wire _w16533_ ;
	wire _w16532_ ;
	wire _w16531_ ;
	wire _w16530_ ;
	wire _w16529_ ;
	wire _w16528_ ;
	wire _w16527_ ;
	wire _w16526_ ;
	wire _w16525_ ;
	wire _w16524_ ;
	wire _w16523_ ;
	wire _w16522_ ;
	wire _w16521_ ;
	wire _w16520_ ;
	wire _w16519_ ;
	wire _w16518_ ;
	wire _w16517_ ;
	wire _w16516_ ;
	wire _w16515_ ;
	wire _w16514_ ;
	wire _w16513_ ;
	wire _w16512_ ;
	wire _w16511_ ;
	wire _w16510_ ;
	wire _w16509_ ;
	wire _w16508_ ;
	wire _w16507_ ;
	wire _w16506_ ;
	wire _w16505_ ;
	wire _w16504_ ;
	wire _w16503_ ;
	wire _w16502_ ;
	wire _w16501_ ;
	wire _w16500_ ;
	wire _w16499_ ;
	wire _w16498_ ;
	wire _w16497_ ;
	wire _w16496_ ;
	wire _w16495_ ;
	wire _w16494_ ;
	wire _w16493_ ;
	wire _w16492_ ;
	wire _w16491_ ;
	wire _w16490_ ;
	wire _w16489_ ;
	wire _w16488_ ;
	wire _w16487_ ;
	wire _w16486_ ;
	wire _w16485_ ;
	wire _w16484_ ;
	wire _w16483_ ;
	wire _w16482_ ;
	wire _w16481_ ;
	wire _w16480_ ;
	wire _w16479_ ;
	wire _w16478_ ;
	wire _w16477_ ;
	wire _w16476_ ;
	wire _w16475_ ;
	wire _w16474_ ;
	wire _w16473_ ;
	wire _w16472_ ;
	wire _w16471_ ;
	wire _w16470_ ;
	wire _w16469_ ;
	wire _w16468_ ;
	wire _w16467_ ;
	wire _w16466_ ;
	wire _w16465_ ;
	wire _w16464_ ;
	wire _w16463_ ;
	wire _w16462_ ;
	wire _w16461_ ;
	wire _w16460_ ;
	wire _w16459_ ;
	wire _w16458_ ;
	wire _w16457_ ;
	wire _w16456_ ;
	wire _w16455_ ;
	wire _w16454_ ;
	wire _w16453_ ;
	wire _w16452_ ;
	wire _w16451_ ;
	wire _w16450_ ;
	wire _w16449_ ;
	wire _w16448_ ;
	wire _w16447_ ;
	wire _w16446_ ;
	wire _w16445_ ;
	wire _w16444_ ;
	wire _w16443_ ;
	wire _w16442_ ;
	wire _w16441_ ;
	wire _w16440_ ;
	wire _w16439_ ;
	wire _w16438_ ;
	wire _w16437_ ;
	wire _w16436_ ;
	wire _w16435_ ;
	wire _w16434_ ;
	wire _w16433_ ;
	wire _w16432_ ;
	wire _w16431_ ;
	wire _w16430_ ;
	wire _w16429_ ;
	wire _w16428_ ;
	wire _w16427_ ;
	wire _w16426_ ;
	wire _w16425_ ;
	wire _w16424_ ;
	wire _w16423_ ;
	wire _w16422_ ;
	wire _w16421_ ;
	wire _w16420_ ;
	wire _w16419_ ;
	wire _w16418_ ;
	wire _w16417_ ;
	wire _w16416_ ;
	wire _w16415_ ;
	wire _w16414_ ;
	wire _w16413_ ;
	wire _w16412_ ;
	wire _w16411_ ;
	wire _w16410_ ;
	wire _w16409_ ;
	wire _w16408_ ;
	wire _w16407_ ;
	wire _w16406_ ;
	wire _w16405_ ;
	wire _w16404_ ;
	wire _w16403_ ;
	wire _w16402_ ;
	wire _w16401_ ;
	wire _w16400_ ;
	wire _w16399_ ;
	wire _w16398_ ;
	wire _w16397_ ;
	wire _w16396_ ;
	wire _w16395_ ;
	wire _w16394_ ;
	wire _w16393_ ;
	wire _w16392_ ;
	wire _w16391_ ;
	wire _w16390_ ;
	wire _w16389_ ;
	wire _w16388_ ;
	wire _w16387_ ;
	wire _w16386_ ;
	wire _w16385_ ;
	wire _w16384_ ;
	wire _w16383_ ;
	wire _w16382_ ;
	wire _w16381_ ;
	wire _w16380_ ;
	wire _w16379_ ;
	wire _w16378_ ;
	wire _w16377_ ;
	wire _w16376_ ;
	wire _w16375_ ;
	wire _w16374_ ;
	wire _w16373_ ;
	wire _w16372_ ;
	wire _w16371_ ;
	wire _w16370_ ;
	wire _w16369_ ;
	wire _w16368_ ;
	wire _w16367_ ;
	wire _w16366_ ;
	wire _w16365_ ;
	wire _w16364_ ;
	wire _w16363_ ;
	wire _w16362_ ;
	wire _w16361_ ;
	wire _w16360_ ;
	wire _w16359_ ;
	wire _w16358_ ;
	wire _w16357_ ;
	wire _w16356_ ;
	wire _w16355_ ;
	wire _w16354_ ;
	wire _w16353_ ;
	wire _w16352_ ;
	wire _w16351_ ;
	wire _w16350_ ;
	wire _w16349_ ;
	wire _w16348_ ;
	wire _w16347_ ;
	wire _w16346_ ;
	wire _w16345_ ;
	wire _w16344_ ;
	wire _w16343_ ;
	wire _w16342_ ;
	wire _w16341_ ;
	wire _w16340_ ;
	wire _w16339_ ;
	wire _w16338_ ;
	wire _w16337_ ;
	wire _w16336_ ;
	wire _w16335_ ;
	wire _w16334_ ;
	wire _w16333_ ;
	wire _w16332_ ;
	wire _w16331_ ;
	wire _w16330_ ;
	wire _w16329_ ;
	wire _w16328_ ;
	wire _w16327_ ;
	wire _w16326_ ;
	wire _w16325_ ;
	wire _w16324_ ;
	wire _w16323_ ;
	wire _w16322_ ;
	wire _w16321_ ;
	wire _w16320_ ;
	wire _w16319_ ;
	wire _w16318_ ;
	wire _w16317_ ;
	wire _w16316_ ;
	wire _w16315_ ;
	wire _w16314_ ;
	wire _w16313_ ;
	wire _w16312_ ;
	wire _w16311_ ;
	wire _w16310_ ;
	wire _w16309_ ;
	wire _w16308_ ;
	wire _w16307_ ;
	wire _w16306_ ;
	wire _w16305_ ;
	wire _w16304_ ;
	wire _w16303_ ;
	wire _w16302_ ;
	wire _w16301_ ;
	wire _w16300_ ;
	wire _w16299_ ;
	wire _w16298_ ;
	wire _w16297_ ;
	wire _w16296_ ;
	wire _w16295_ ;
	wire _w16294_ ;
	wire _w16293_ ;
	wire _w16292_ ;
	wire _w16291_ ;
	wire _w16290_ ;
	wire _w16289_ ;
	wire _w16288_ ;
	wire _w16287_ ;
	wire _w16286_ ;
	wire _w16285_ ;
	wire _w16284_ ;
	wire _w16283_ ;
	wire _w16282_ ;
	wire _w16281_ ;
	wire _w16280_ ;
	wire _w16279_ ;
	wire _w16278_ ;
	wire _w16277_ ;
	wire _w16276_ ;
	wire _w16275_ ;
	wire _w16274_ ;
	wire _w16273_ ;
	wire _w16272_ ;
	wire _w16271_ ;
	wire _w16270_ ;
	wire _w16269_ ;
	wire _w16268_ ;
	wire _w16267_ ;
	wire _w16266_ ;
	wire _w16265_ ;
	wire _w16264_ ;
	wire _w16263_ ;
	wire _w16262_ ;
	wire _w16261_ ;
	wire _w16260_ ;
	wire _w16259_ ;
	wire _w16258_ ;
	wire _w16257_ ;
	wire _w16256_ ;
	wire _w16255_ ;
	wire _w16254_ ;
	wire _w16253_ ;
	wire _w16252_ ;
	wire _w16251_ ;
	wire _w16250_ ;
	wire _w16249_ ;
	wire _w16248_ ;
	wire _w16247_ ;
	wire _w16246_ ;
	wire _w16245_ ;
	wire _w16244_ ;
	wire _w16243_ ;
	wire _w16242_ ;
	wire _w16241_ ;
	wire _w16240_ ;
	wire _w16239_ ;
	wire _w16238_ ;
	wire _w16237_ ;
	wire _w16236_ ;
	wire _w16235_ ;
	wire _w16234_ ;
	wire _w16233_ ;
	wire _w16232_ ;
	wire _w16231_ ;
	wire _w16230_ ;
	wire _w16229_ ;
	wire _w16228_ ;
	wire _w16227_ ;
	wire _w16226_ ;
	wire _w16225_ ;
	wire _w16224_ ;
	wire _w16223_ ;
	wire _w16222_ ;
	wire _w16221_ ;
	wire _w16220_ ;
	wire _w16219_ ;
	wire _w16218_ ;
	wire _w16217_ ;
	wire _w16216_ ;
	wire _w16215_ ;
	wire _w16214_ ;
	wire _w16213_ ;
	wire _w16212_ ;
	wire _w16211_ ;
	wire _w16210_ ;
	wire _w16209_ ;
	wire _w16208_ ;
	wire _w16207_ ;
	wire _w16206_ ;
	wire _w16205_ ;
	wire _w16204_ ;
	wire _w16203_ ;
	wire _w16202_ ;
	wire _w16201_ ;
	wire _w16200_ ;
	wire _w16199_ ;
	wire _w16198_ ;
	wire _w16197_ ;
	wire _w16196_ ;
	wire _w16195_ ;
	wire _w16194_ ;
	wire _w16193_ ;
	wire _w16192_ ;
	wire _w16191_ ;
	wire _w16190_ ;
	wire _w16189_ ;
	wire _w16188_ ;
	wire _w16187_ ;
	wire _w16186_ ;
	wire _w16185_ ;
	wire _w16184_ ;
	wire _w16183_ ;
	wire _w16182_ ;
	wire _w16181_ ;
	wire _w16180_ ;
	wire _w16179_ ;
	wire _w16178_ ;
	wire _w16177_ ;
	wire _w16176_ ;
	wire _w16175_ ;
	wire _w16174_ ;
	wire _w16173_ ;
	wire _w16172_ ;
	wire _w16171_ ;
	wire _w16170_ ;
	wire _w16169_ ;
	wire _w16168_ ;
	wire _w16167_ ;
	wire _w16166_ ;
	wire _w16165_ ;
	wire _w16164_ ;
	wire _w16163_ ;
	wire _w16162_ ;
	wire _w16161_ ;
	wire _w16160_ ;
	wire _w16159_ ;
	wire _w16158_ ;
	wire _w16157_ ;
	wire _w16156_ ;
	wire _w16155_ ;
	wire _w16154_ ;
	wire _w16153_ ;
	wire _w16152_ ;
	wire _w16151_ ;
	wire _w16150_ ;
	wire _w16149_ ;
	wire _w16148_ ;
	wire _w16147_ ;
	wire _w16146_ ;
	wire _w16145_ ;
	wire _w16144_ ;
	wire _w16143_ ;
	wire _w16142_ ;
	wire _w16141_ ;
	wire _w16140_ ;
	wire _w16139_ ;
	wire _w16138_ ;
	wire _w16137_ ;
	wire _w16136_ ;
	wire _w16135_ ;
	wire _w16134_ ;
	wire _w16133_ ;
	wire _w16132_ ;
	wire _w16131_ ;
	wire _w16130_ ;
	wire _w16129_ ;
	wire _w16128_ ;
	wire _w16127_ ;
	wire _w16126_ ;
	wire _w16125_ ;
	wire _w16124_ ;
	wire _w16123_ ;
	wire _w16122_ ;
	wire _w16121_ ;
	wire _w16120_ ;
	wire _w16119_ ;
	wire _w16118_ ;
	wire _w16117_ ;
	wire _w16116_ ;
	wire _w16115_ ;
	wire _w16114_ ;
	wire _w16113_ ;
	wire _w16112_ ;
	wire _w16111_ ;
	wire _w16110_ ;
	wire _w16109_ ;
	wire _w16108_ ;
	wire _w16107_ ;
	wire _w16106_ ;
	wire _w16105_ ;
	wire _w16104_ ;
	wire _w16103_ ;
	wire _w16102_ ;
	wire _w16101_ ;
	wire _w16100_ ;
	wire _w16099_ ;
	wire _w16098_ ;
	wire _w16097_ ;
	wire _w16096_ ;
	wire _w16095_ ;
	wire _w16094_ ;
	wire _w16093_ ;
	wire _w16092_ ;
	wire _w16091_ ;
	wire _w16090_ ;
	wire _w16089_ ;
	wire _w16088_ ;
	wire _w16087_ ;
	wire _w16086_ ;
	wire _w16085_ ;
	wire _w16084_ ;
	wire _w16083_ ;
	wire _w16082_ ;
	wire _w16081_ ;
	wire _w16080_ ;
	wire _w16079_ ;
	wire _w16078_ ;
	wire _w16077_ ;
	wire _w16076_ ;
	wire _w16075_ ;
	wire _w16074_ ;
	wire _w16073_ ;
	wire _w16072_ ;
	wire _w16071_ ;
	wire _w16070_ ;
	wire _w16069_ ;
	wire _w16068_ ;
	wire _w16067_ ;
	wire _w16066_ ;
	wire _w16065_ ;
	wire _w16064_ ;
	wire _w16063_ ;
	wire _w16062_ ;
	wire _w16061_ ;
	wire _w16060_ ;
	wire _w16059_ ;
	wire _w16058_ ;
	wire _w16057_ ;
	wire _w16056_ ;
	wire _w16055_ ;
	wire _w16054_ ;
	wire _w16053_ ;
	wire _w16052_ ;
	wire _w16051_ ;
	wire _w16050_ ;
	wire _w16049_ ;
	wire _w16048_ ;
	wire _w16047_ ;
	wire _w16046_ ;
	wire _w16045_ ;
	wire _w16044_ ;
	wire _w16043_ ;
	wire _w16042_ ;
	wire _w16041_ ;
	wire _w16040_ ;
	wire _w16039_ ;
	wire _w16038_ ;
	wire _w16037_ ;
	wire _w16036_ ;
	wire _w16035_ ;
	wire _w16034_ ;
	wire _w16033_ ;
	wire _w16032_ ;
	wire _w16031_ ;
	wire _w16030_ ;
	wire _w16029_ ;
	wire _w16028_ ;
	wire _w16027_ ;
	wire _w16026_ ;
	wire _w16025_ ;
	wire _w16024_ ;
	wire _w16023_ ;
	wire _w16022_ ;
	wire _w16021_ ;
	wire _w16020_ ;
	wire _w16019_ ;
	wire _w16018_ ;
	wire _w16017_ ;
	wire _w16016_ ;
	wire _w16015_ ;
	wire _w16014_ ;
	wire _w16013_ ;
	wire _w16012_ ;
	wire _w16011_ ;
	wire _w16010_ ;
	wire _w16009_ ;
	wire _w16008_ ;
	wire _w16007_ ;
	wire _w16006_ ;
	wire _w16005_ ;
	wire _w16004_ ;
	wire _w16003_ ;
	wire _w16002_ ;
	wire _w16001_ ;
	wire _w16000_ ;
	wire _w15999_ ;
	wire _w15998_ ;
	wire _w15997_ ;
	wire _w15996_ ;
	wire _w15995_ ;
	wire _w15994_ ;
	wire _w15993_ ;
	wire _w15992_ ;
	wire _w15991_ ;
	wire _w15990_ ;
	wire _w15989_ ;
	wire _w15988_ ;
	wire _w15987_ ;
	wire _w15986_ ;
	wire _w15985_ ;
	wire _w15984_ ;
	wire _w15983_ ;
	wire _w15982_ ;
	wire _w15981_ ;
	wire _w15980_ ;
	wire _w15979_ ;
	wire _w15978_ ;
	wire _w15977_ ;
	wire _w15976_ ;
	wire _w15975_ ;
	wire _w15974_ ;
	wire _w15973_ ;
	wire _w15972_ ;
	wire _w15971_ ;
	wire _w15970_ ;
	wire _w15969_ ;
	wire _w15968_ ;
	wire _w15967_ ;
	wire _w15966_ ;
	wire _w15965_ ;
	wire _w15964_ ;
	wire _w15963_ ;
	wire _w15962_ ;
	wire _w15961_ ;
	wire _w15960_ ;
	wire _w15959_ ;
	wire _w15958_ ;
	wire _w15957_ ;
	wire _w15956_ ;
	wire _w15955_ ;
	wire _w15954_ ;
	wire _w15953_ ;
	wire _w15952_ ;
	wire _w15951_ ;
	wire _w15950_ ;
	wire _w15949_ ;
	wire _w15948_ ;
	wire _w15947_ ;
	wire _w15946_ ;
	wire _w15945_ ;
	wire _w15944_ ;
	wire _w15943_ ;
	wire _w15942_ ;
	wire _w15941_ ;
	wire _w15940_ ;
	wire _w15939_ ;
	wire _w15938_ ;
	wire _w15937_ ;
	wire _w15936_ ;
	wire _w15935_ ;
	wire _w15934_ ;
	wire _w15933_ ;
	wire _w15932_ ;
	wire _w15931_ ;
	wire _w15930_ ;
	wire _w15929_ ;
	wire _w15928_ ;
	wire _w15927_ ;
	wire _w15926_ ;
	wire _w15925_ ;
	wire _w15924_ ;
	wire _w15923_ ;
	wire _w15922_ ;
	wire _w15921_ ;
	wire _w15920_ ;
	wire _w15919_ ;
	wire _w15918_ ;
	wire _w15917_ ;
	wire _w15916_ ;
	wire _w15915_ ;
	wire _w15914_ ;
	wire _w15913_ ;
	wire _w15912_ ;
	wire _w15911_ ;
	wire _w15910_ ;
	wire _w15909_ ;
	wire _w15908_ ;
	wire _w15907_ ;
	wire _w15906_ ;
	wire _w15905_ ;
	wire _w15904_ ;
	wire _w15903_ ;
	wire _w15902_ ;
	wire _w15901_ ;
	wire _w15900_ ;
	wire _w15899_ ;
	wire _w15898_ ;
	wire _w15897_ ;
	wire _w15896_ ;
	wire _w15895_ ;
	wire _w15894_ ;
	wire _w15893_ ;
	wire _w15892_ ;
	wire _w15891_ ;
	wire _w15890_ ;
	wire _w15889_ ;
	wire _w15888_ ;
	wire _w15887_ ;
	wire _w15886_ ;
	wire _w15885_ ;
	wire _w15884_ ;
	wire _w15883_ ;
	wire _w15882_ ;
	wire _w15881_ ;
	wire _w15880_ ;
	wire _w15879_ ;
	wire _w15878_ ;
	wire _w15877_ ;
	wire _w15876_ ;
	wire _w15875_ ;
	wire _w15874_ ;
	wire _w15873_ ;
	wire _w15872_ ;
	wire _w15871_ ;
	wire _w15870_ ;
	wire _w15869_ ;
	wire _w15868_ ;
	wire _w15867_ ;
	wire _w15866_ ;
	wire _w15865_ ;
	wire _w15864_ ;
	wire _w15863_ ;
	wire _w15862_ ;
	wire _w15861_ ;
	wire _w15860_ ;
	wire _w15859_ ;
	wire _w15858_ ;
	wire _w15857_ ;
	wire _w15856_ ;
	wire _w15855_ ;
	wire _w15854_ ;
	wire _w15853_ ;
	wire _w15852_ ;
	wire _w15851_ ;
	wire _w15850_ ;
	wire _w15849_ ;
	wire _w15848_ ;
	wire _w15847_ ;
	wire _w15846_ ;
	wire _w15845_ ;
	wire _w15844_ ;
	wire _w15843_ ;
	wire _w15842_ ;
	wire _w15841_ ;
	wire _w15840_ ;
	wire _w15839_ ;
	wire _w15838_ ;
	wire _w15837_ ;
	wire _w15836_ ;
	wire _w15835_ ;
	wire _w15834_ ;
	wire _w15833_ ;
	wire _w15832_ ;
	wire _w15831_ ;
	wire _w15830_ ;
	wire _w15829_ ;
	wire _w15828_ ;
	wire _w15827_ ;
	wire _w15826_ ;
	wire _w15825_ ;
	wire _w15824_ ;
	wire _w15823_ ;
	wire _w15822_ ;
	wire _w15821_ ;
	wire _w15820_ ;
	wire _w15819_ ;
	wire _w15818_ ;
	wire _w15817_ ;
	wire _w15816_ ;
	wire _w15815_ ;
	wire _w15814_ ;
	wire _w15813_ ;
	wire _w15812_ ;
	wire _w15811_ ;
	wire _w15810_ ;
	wire _w15809_ ;
	wire _w15808_ ;
	wire _w15807_ ;
	wire _w15806_ ;
	wire _w15805_ ;
	wire _w15804_ ;
	wire _w15803_ ;
	wire _w15802_ ;
	wire _w15801_ ;
	wire _w15800_ ;
	wire _w15799_ ;
	wire _w15798_ ;
	wire _w15797_ ;
	wire _w15796_ ;
	wire _w15795_ ;
	wire _w15794_ ;
	wire _w15793_ ;
	wire _w15792_ ;
	wire _w15791_ ;
	wire _w15790_ ;
	wire _w15789_ ;
	wire _w15788_ ;
	wire _w15787_ ;
	wire _w15786_ ;
	wire _w15785_ ;
	wire _w15784_ ;
	wire _w15783_ ;
	wire _w15782_ ;
	wire _w15781_ ;
	wire _w15780_ ;
	wire _w15779_ ;
	wire _w15778_ ;
	wire _w15777_ ;
	wire _w15776_ ;
	wire _w15775_ ;
	wire _w15774_ ;
	wire _w15773_ ;
	wire _w15772_ ;
	wire _w15771_ ;
	wire _w15770_ ;
	wire _w15769_ ;
	wire _w15768_ ;
	wire _w15767_ ;
	wire _w15766_ ;
	wire _w15765_ ;
	wire _w15764_ ;
	wire _w15763_ ;
	wire _w15762_ ;
	wire _w15761_ ;
	wire _w15760_ ;
	wire _w15759_ ;
	wire _w15758_ ;
	wire _w15757_ ;
	wire _w15756_ ;
	wire _w15755_ ;
	wire _w15754_ ;
	wire _w15753_ ;
	wire _w15752_ ;
	wire _w15751_ ;
	wire _w15750_ ;
	wire _w15749_ ;
	wire _w15748_ ;
	wire _w15747_ ;
	wire _w15746_ ;
	wire _w15745_ ;
	wire _w15744_ ;
	wire _w15743_ ;
	wire _w15742_ ;
	wire _w15741_ ;
	wire _w15740_ ;
	wire _w15739_ ;
	wire _w15738_ ;
	wire _w15737_ ;
	wire _w15736_ ;
	wire _w15735_ ;
	wire _w15734_ ;
	wire _w15733_ ;
	wire _w15732_ ;
	wire _w15731_ ;
	wire _w15730_ ;
	wire _w15729_ ;
	wire _w15728_ ;
	wire _w15727_ ;
	wire _w15726_ ;
	wire _w15725_ ;
	wire _w15724_ ;
	wire _w15723_ ;
	wire _w15722_ ;
	wire _w15721_ ;
	wire _w15720_ ;
	wire _w15719_ ;
	wire _w15718_ ;
	wire _w15717_ ;
	wire _w15716_ ;
	wire _w15715_ ;
	wire _w15714_ ;
	wire _w15713_ ;
	wire _w15712_ ;
	wire _w15711_ ;
	wire _w15710_ ;
	wire _w15709_ ;
	wire _w15708_ ;
	wire _w15707_ ;
	wire _w15706_ ;
	wire _w15705_ ;
	wire _w15704_ ;
	wire _w15703_ ;
	wire _w15702_ ;
	wire _w15701_ ;
	wire _w15700_ ;
	wire _w15699_ ;
	wire _w15698_ ;
	wire _w15697_ ;
	wire _w15696_ ;
	wire _w15695_ ;
	wire _w15694_ ;
	wire _w15693_ ;
	wire _w15692_ ;
	wire _w15691_ ;
	wire _w15690_ ;
	wire _w15689_ ;
	wire _w15688_ ;
	wire _w15687_ ;
	wire _w15686_ ;
	wire _w15685_ ;
	wire _w15684_ ;
	wire _w15683_ ;
	wire _w15682_ ;
	wire _w15681_ ;
	wire _w15680_ ;
	wire _w15679_ ;
	wire _w15678_ ;
	wire _w15677_ ;
	wire _w15676_ ;
	wire _w15675_ ;
	wire _w15674_ ;
	wire _w15673_ ;
	wire _w15672_ ;
	wire _w15671_ ;
	wire _w15670_ ;
	wire _w15669_ ;
	wire _w15668_ ;
	wire _w15667_ ;
	wire _w15666_ ;
	wire _w15665_ ;
	wire _w15664_ ;
	wire _w15663_ ;
	wire _w15662_ ;
	wire _w15661_ ;
	wire _w15660_ ;
	wire _w15659_ ;
	wire _w15658_ ;
	wire _w15657_ ;
	wire _w15656_ ;
	wire _w15655_ ;
	wire _w15654_ ;
	wire _w15653_ ;
	wire _w15652_ ;
	wire _w15651_ ;
	wire _w15650_ ;
	wire _w15649_ ;
	wire _w15648_ ;
	wire _w15647_ ;
	wire _w15646_ ;
	wire _w15645_ ;
	wire _w15644_ ;
	wire _w15643_ ;
	wire _w15642_ ;
	wire _w15641_ ;
	wire _w15640_ ;
	wire _w15639_ ;
	wire _w15638_ ;
	wire _w15637_ ;
	wire _w15636_ ;
	wire _w15635_ ;
	wire _w15634_ ;
	wire _w15633_ ;
	wire _w15632_ ;
	wire _w15631_ ;
	wire _w15630_ ;
	wire _w15629_ ;
	wire _w15628_ ;
	wire _w15627_ ;
	wire _w15626_ ;
	wire _w15625_ ;
	wire _w15624_ ;
	wire _w15623_ ;
	wire _w15622_ ;
	wire _w15621_ ;
	wire _w15620_ ;
	wire _w15619_ ;
	wire _w15618_ ;
	wire _w15617_ ;
	wire _w15616_ ;
	wire _w15615_ ;
	wire _w15614_ ;
	wire _w15613_ ;
	wire _w15612_ ;
	wire _w15611_ ;
	wire _w15610_ ;
	wire _w15609_ ;
	wire _w15608_ ;
	wire _w15607_ ;
	wire _w15606_ ;
	wire _w15605_ ;
	wire _w15604_ ;
	wire _w15603_ ;
	wire _w15602_ ;
	wire _w15601_ ;
	wire _w15600_ ;
	wire _w15599_ ;
	wire _w15598_ ;
	wire _w15597_ ;
	wire _w15596_ ;
	wire _w15595_ ;
	wire _w15594_ ;
	wire _w15593_ ;
	wire _w15592_ ;
	wire _w15591_ ;
	wire _w15590_ ;
	wire _w15589_ ;
	wire _w15588_ ;
	wire _w15587_ ;
	wire _w15586_ ;
	wire _w15585_ ;
	wire _w15584_ ;
	wire _w15583_ ;
	wire _w15582_ ;
	wire _w15581_ ;
	wire _w15580_ ;
	wire _w15579_ ;
	wire _w15578_ ;
	wire _w15577_ ;
	wire _w15576_ ;
	wire _w15575_ ;
	wire _w15574_ ;
	wire _w15573_ ;
	wire _w15572_ ;
	wire _w15571_ ;
	wire _w15570_ ;
	wire _w15569_ ;
	wire _w15568_ ;
	wire _w15567_ ;
	wire _w15566_ ;
	wire _w15565_ ;
	wire _w15564_ ;
	wire _w15563_ ;
	wire _w15562_ ;
	wire _w15561_ ;
	wire _w15560_ ;
	wire _w15559_ ;
	wire _w15558_ ;
	wire _w15557_ ;
	wire _w15556_ ;
	wire _w15555_ ;
	wire _w15554_ ;
	wire _w15553_ ;
	wire _w15552_ ;
	wire _w15551_ ;
	wire _w15550_ ;
	wire _w15549_ ;
	wire _w15548_ ;
	wire _w15547_ ;
	wire _w15546_ ;
	wire _w15545_ ;
	wire _w15544_ ;
	wire _w15543_ ;
	wire _w15542_ ;
	wire _w15541_ ;
	wire _w15540_ ;
	wire _w15539_ ;
	wire _w15538_ ;
	wire _w15537_ ;
	wire _w15536_ ;
	wire _w15535_ ;
	wire _w15534_ ;
	wire _w15533_ ;
	wire _w15532_ ;
	wire _w15531_ ;
	wire _w15530_ ;
	wire _w15529_ ;
	wire _w15528_ ;
	wire _w15527_ ;
	wire _w15526_ ;
	wire _w15525_ ;
	wire _w15524_ ;
	wire _w15523_ ;
	wire _w15522_ ;
	wire _w15521_ ;
	wire _w15520_ ;
	wire _w15519_ ;
	wire _w15518_ ;
	wire _w15517_ ;
	wire _w15516_ ;
	wire _w15515_ ;
	wire _w15514_ ;
	wire _w15513_ ;
	wire _w15512_ ;
	wire _w15511_ ;
	wire _w15510_ ;
	wire _w15509_ ;
	wire _w15508_ ;
	wire _w15507_ ;
	wire _w15506_ ;
	wire _w15505_ ;
	wire _w15504_ ;
	wire _w15503_ ;
	wire _w15502_ ;
	wire _w15501_ ;
	wire _w15500_ ;
	wire _w15499_ ;
	wire _w15498_ ;
	wire _w15497_ ;
	wire _w15496_ ;
	wire _w15495_ ;
	wire _w15494_ ;
	wire _w15493_ ;
	wire _w15492_ ;
	wire _w15491_ ;
	wire _w15490_ ;
	wire _w15489_ ;
	wire _w15488_ ;
	wire _w15487_ ;
	wire _w15486_ ;
	wire _w15485_ ;
	wire _w15484_ ;
	wire _w15483_ ;
	wire _w15482_ ;
	wire _w15481_ ;
	wire _w15480_ ;
	wire _w15479_ ;
	wire _w15478_ ;
	wire _w15477_ ;
	wire _w15476_ ;
	wire _w15475_ ;
	wire _w15474_ ;
	wire _w15473_ ;
	wire _w15472_ ;
	wire _w15471_ ;
	wire _w15470_ ;
	wire _w15469_ ;
	wire _w15468_ ;
	wire _w15467_ ;
	wire _w15466_ ;
	wire _w15465_ ;
	wire _w15464_ ;
	wire _w15463_ ;
	wire _w15462_ ;
	wire _w15461_ ;
	wire _w15460_ ;
	wire _w15459_ ;
	wire _w15458_ ;
	wire _w15457_ ;
	wire _w15456_ ;
	wire _w15455_ ;
	wire _w15454_ ;
	wire _w15453_ ;
	wire _w15452_ ;
	wire _w15451_ ;
	wire _w15450_ ;
	wire _w15449_ ;
	wire _w15448_ ;
	wire _w15447_ ;
	wire _w15446_ ;
	wire _w15445_ ;
	wire _w15444_ ;
	wire _w15443_ ;
	wire _w15442_ ;
	wire _w15441_ ;
	wire _w15440_ ;
	wire _w15439_ ;
	wire _w15438_ ;
	wire _w15437_ ;
	wire _w15436_ ;
	wire _w15435_ ;
	wire _w15434_ ;
	wire _w15433_ ;
	wire _w15432_ ;
	wire _w15431_ ;
	wire _w15430_ ;
	wire _w15429_ ;
	wire _w15428_ ;
	wire _w15427_ ;
	wire _w15426_ ;
	wire _w15425_ ;
	wire _w15424_ ;
	wire _w15423_ ;
	wire _w15422_ ;
	wire _w15421_ ;
	wire _w15420_ ;
	wire _w15419_ ;
	wire _w15418_ ;
	wire _w15417_ ;
	wire _w15416_ ;
	wire _w15415_ ;
	wire _w15414_ ;
	wire _w15413_ ;
	wire _w15412_ ;
	wire _w15411_ ;
	wire _w15410_ ;
	wire _w15409_ ;
	wire _w15408_ ;
	wire _w15407_ ;
	wire _w15406_ ;
	wire _w15405_ ;
	wire _w15404_ ;
	wire _w15403_ ;
	wire _w15402_ ;
	wire _w15401_ ;
	wire _w15400_ ;
	wire _w15399_ ;
	wire _w15398_ ;
	wire _w15397_ ;
	wire _w15396_ ;
	wire _w15395_ ;
	wire _w15394_ ;
	wire _w15393_ ;
	wire _w15392_ ;
	wire _w15391_ ;
	wire _w15390_ ;
	wire _w15389_ ;
	wire _w15388_ ;
	wire _w15387_ ;
	wire _w15386_ ;
	wire _w15385_ ;
	wire _w15384_ ;
	wire _w15383_ ;
	wire _w15382_ ;
	wire _w15381_ ;
	wire _w15380_ ;
	wire _w15379_ ;
	wire _w15378_ ;
	wire _w15377_ ;
	wire _w15376_ ;
	wire _w15375_ ;
	wire _w15374_ ;
	wire _w15373_ ;
	wire _w15372_ ;
	wire _w15371_ ;
	wire _w15370_ ;
	wire _w15369_ ;
	wire _w15368_ ;
	wire _w15367_ ;
	wire _w15366_ ;
	wire _w15365_ ;
	wire _w15364_ ;
	wire _w15363_ ;
	wire _w15362_ ;
	wire _w15361_ ;
	wire _w15360_ ;
	wire _w15359_ ;
	wire _w15358_ ;
	wire _w15357_ ;
	wire _w15356_ ;
	wire _w15355_ ;
	wire _w15354_ ;
	wire _w15353_ ;
	wire _w15352_ ;
	wire _w15351_ ;
	wire _w15350_ ;
	wire _w15349_ ;
	wire _w15348_ ;
	wire _w15347_ ;
	wire _w15346_ ;
	wire _w15345_ ;
	wire _w15344_ ;
	wire _w15343_ ;
	wire _w15342_ ;
	wire _w15341_ ;
	wire _w15340_ ;
	wire _w15339_ ;
	wire _w15338_ ;
	wire _w15337_ ;
	wire _w15336_ ;
	wire _w15335_ ;
	wire _w15334_ ;
	wire _w15333_ ;
	wire _w15332_ ;
	wire _w15331_ ;
	wire _w15330_ ;
	wire _w15329_ ;
	wire _w15328_ ;
	wire _w15327_ ;
	wire _w15326_ ;
	wire _w15325_ ;
	wire _w15324_ ;
	wire _w15323_ ;
	wire _w15322_ ;
	wire _w15321_ ;
	wire _w15320_ ;
	wire _w15319_ ;
	wire _w15318_ ;
	wire _w15317_ ;
	wire _w15316_ ;
	wire _w15315_ ;
	wire _w15314_ ;
	wire _w15313_ ;
	wire _w15312_ ;
	wire _w15311_ ;
	wire _w15310_ ;
	wire _w15309_ ;
	wire _w15308_ ;
	wire _w15307_ ;
	wire _w15306_ ;
	wire _w15305_ ;
	wire _w15304_ ;
	wire _w15303_ ;
	wire _w15302_ ;
	wire _w15301_ ;
	wire _w15300_ ;
	wire _w15299_ ;
	wire _w15298_ ;
	wire _w15297_ ;
	wire _w15296_ ;
	wire _w15295_ ;
	wire _w15294_ ;
	wire _w15293_ ;
	wire _w15292_ ;
	wire _w15291_ ;
	wire _w15290_ ;
	wire _w15289_ ;
	wire _w15288_ ;
	wire _w15287_ ;
	wire _w15286_ ;
	wire _w15285_ ;
	wire _w15284_ ;
	wire _w15283_ ;
	wire _w15282_ ;
	wire _w15281_ ;
	wire _w15280_ ;
	wire _w15279_ ;
	wire _w15278_ ;
	wire _w15277_ ;
	wire _w15276_ ;
	wire _w15275_ ;
	wire _w15274_ ;
	wire _w15273_ ;
	wire _w15272_ ;
	wire _w15271_ ;
	wire _w15270_ ;
	wire _w15269_ ;
	wire _w15268_ ;
	wire _w15267_ ;
	wire _w15266_ ;
	wire _w15265_ ;
	wire _w15264_ ;
	wire _w15263_ ;
	wire _w15262_ ;
	wire _w15261_ ;
	wire _w15260_ ;
	wire _w15259_ ;
	wire _w15258_ ;
	wire _w15257_ ;
	wire _w15256_ ;
	wire _w15255_ ;
	wire _w15254_ ;
	wire _w15253_ ;
	wire _w15252_ ;
	wire _w15251_ ;
	wire _w15250_ ;
	wire _w15249_ ;
	wire _w15248_ ;
	wire _w15247_ ;
	wire _w15246_ ;
	wire _w15245_ ;
	wire _w15244_ ;
	wire _w15243_ ;
	wire _w15242_ ;
	wire _w15241_ ;
	wire _w15240_ ;
	wire _w15239_ ;
	wire _w15238_ ;
	wire _w15237_ ;
	wire _w15236_ ;
	wire _w15235_ ;
	wire _w15234_ ;
	wire _w15233_ ;
	wire _w15232_ ;
	wire _w15231_ ;
	wire _w15230_ ;
	wire _w15229_ ;
	wire _w15228_ ;
	wire _w15227_ ;
	wire _w15226_ ;
	wire _w15225_ ;
	wire _w15224_ ;
	wire _w15223_ ;
	wire _w15222_ ;
	wire _w15221_ ;
	wire _w15220_ ;
	wire _w15219_ ;
	wire _w15218_ ;
	wire _w15217_ ;
	wire _w15216_ ;
	wire _w15215_ ;
	wire _w15214_ ;
	wire _w15213_ ;
	wire _w15212_ ;
	wire _w15211_ ;
	wire _w15210_ ;
	wire _w15209_ ;
	wire _w15208_ ;
	wire _w15207_ ;
	wire _w15206_ ;
	wire _w15205_ ;
	wire _w15204_ ;
	wire _w15203_ ;
	wire _w15202_ ;
	wire _w15201_ ;
	wire _w15200_ ;
	wire _w15199_ ;
	wire _w15198_ ;
	wire _w15197_ ;
	wire _w15196_ ;
	wire _w15195_ ;
	wire _w15194_ ;
	wire _w15193_ ;
	wire _w15192_ ;
	wire _w15191_ ;
	wire _w15190_ ;
	wire _w15189_ ;
	wire _w15188_ ;
	wire _w15187_ ;
	wire _w15186_ ;
	wire _w15185_ ;
	wire _w15184_ ;
	wire _w15183_ ;
	wire _w15182_ ;
	wire _w15181_ ;
	wire _w15180_ ;
	wire _w15179_ ;
	wire _w15178_ ;
	wire _w15177_ ;
	wire _w15176_ ;
	wire _w15175_ ;
	wire _w15174_ ;
	wire _w15173_ ;
	wire _w15172_ ;
	wire _w15171_ ;
	wire _w15170_ ;
	wire _w15169_ ;
	wire _w15168_ ;
	wire _w15167_ ;
	wire _w15166_ ;
	wire _w15165_ ;
	wire _w15164_ ;
	wire _w15163_ ;
	wire _w15162_ ;
	wire _w15161_ ;
	wire _w15160_ ;
	wire _w15159_ ;
	wire _w15158_ ;
	wire _w15157_ ;
	wire _w15156_ ;
	wire _w15155_ ;
	wire _w15154_ ;
	wire _w15153_ ;
	wire _w15152_ ;
	wire _w15151_ ;
	wire _w15150_ ;
	wire _w15149_ ;
	wire _w15148_ ;
	wire _w15147_ ;
	wire _w15146_ ;
	wire _w15145_ ;
	wire _w15144_ ;
	wire _w15143_ ;
	wire _w15142_ ;
	wire _w15141_ ;
	wire _w15140_ ;
	wire _w15139_ ;
	wire _w15138_ ;
	wire _w15137_ ;
	wire _w15136_ ;
	wire _w15135_ ;
	wire _w15134_ ;
	wire _w15133_ ;
	wire _w15132_ ;
	wire _w15131_ ;
	wire _w15130_ ;
	wire _w15129_ ;
	wire _w15128_ ;
	wire _w15127_ ;
	wire _w15126_ ;
	wire _w15125_ ;
	wire _w15124_ ;
	wire _w15123_ ;
	wire _w15122_ ;
	wire _w15121_ ;
	wire _w15120_ ;
	wire _w15119_ ;
	wire _w15118_ ;
	wire _w15117_ ;
	wire _w15116_ ;
	wire _w15115_ ;
	wire _w15114_ ;
	wire _w15113_ ;
	wire _w15112_ ;
	wire _w15111_ ;
	wire _w15110_ ;
	wire _w15109_ ;
	wire _w15108_ ;
	wire _w15107_ ;
	wire _w15106_ ;
	wire _w15105_ ;
	wire _w15104_ ;
	wire _w15103_ ;
	wire _w15102_ ;
	wire _w15101_ ;
	wire _w15100_ ;
	wire _w15099_ ;
	wire _w15098_ ;
	wire _w15097_ ;
	wire _w15096_ ;
	wire _w15095_ ;
	wire _w15094_ ;
	wire _w15093_ ;
	wire _w15092_ ;
	wire _w15091_ ;
	wire _w15090_ ;
	wire _w15089_ ;
	wire _w15088_ ;
	wire _w15087_ ;
	wire _w15086_ ;
	wire _w15085_ ;
	wire _w15084_ ;
	wire _w15083_ ;
	wire _w15082_ ;
	wire _w15081_ ;
	wire _w15080_ ;
	wire _w15079_ ;
	wire _w15078_ ;
	wire _w15077_ ;
	wire _w15076_ ;
	wire _w15075_ ;
	wire _w15074_ ;
	wire _w15073_ ;
	wire _w15072_ ;
	wire _w15071_ ;
	wire _w15070_ ;
	wire _w15069_ ;
	wire _w15068_ ;
	wire _w15067_ ;
	wire _w15066_ ;
	wire _w15065_ ;
	wire _w15064_ ;
	wire _w15063_ ;
	wire _w15062_ ;
	wire _w15061_ ;
	wire _w15060_ ;
	wire _w15059_ ;
	wire _w15058_ ;
	wire _w15057_ ;
	wire _w15056_ ;
	wire _w15055_ ;
	wire _w15054_ ;
	wire _w15053_ ;
	wire _w15052_ ;
	wire _w15051_ ;
	wire _w15050_ ;
	wire _w15049_ ;
	wire _w15048_ ;
	wire _w15047_ ;
	wire _w15046_ ;
	wire _w15045_ ;
	wire _w15044_ ;
	wire _w15043_ ;
	wire _w15042_ ;
	wire _w15041_ ;
	wire _w15040_ ;
	wire _w15039_ ;
	wire _w15038_ ;
	wire _w15037_ ;
	wire _w15036_ ;
	wire _w15035_ ;
	wire _w15034_ ;
	wire _w15033_ ;
	wire _w15032_ ;
	wire _w15031_ ;
	wire _w15030_ ;
	wire _w15029_ ;
	wire _w15028_ ;
	wire _w15027_ ;
	wire _w15026_ ;
	wire _w15025_ ;
	wire _w15024_ ;
	wire _w15023_ ;
	wire _w15022_ ;
	wire _w15021_ ;
	wire _w15020_ ;
	wire _w15019_ ;
	wire _w15018_ ;
	wire _w15017_ ;
	wire _w15016_ ;
	wire _w15015_ ;
	wire _w15014_ ;
	wire _w15013_ ;
	wire _w15012_ ;
	wire _w15011_ ;
	wire _w15010_ ;
	wire _w15009_ ;
	wire _w15008_ ;
	wire _w15007_ ;
	wire _w15006_ ;
	wire _w15005_ ;
	wire _w15004_ ;
	wire _w15003_ ;
	wire _w15002_ ;
	wire _w15001_ ;
	wire _w15000_ ;
	wire _w14999_ ;
	wire _w14998_ ;
	wire _w14997_ ;
	wire _w14996_ ;
	wire _w14995_ ;
	wire _w14994_ ;
	wire _w14993_ ;
	wire _w14992_ ;
	wire _w14991_ ;
	wire _w14990_ ;
	wire _w14989_ ;
	wire _w14988_ ;
	wire _w14987_ ;
	wire _w14986_ ;
	wire _w14985_ ;
	wire _w14984_ ;
	wire _w14983_ ;
	wire _w14982_ ;
	wire _w14981_ ;
	wire _w14980_ ;
	wire _w14979_ ;
	wire _w14978_ ;
	wire _w14977_ ;
	wire _w14976_ ;
	wire _w14975_ ;
	wire _w14974_ ;
	wire _w14973_ ;
	wire _w14972_ ;
	wire _w14971_ ;
	wire _w14970_ ;
	wire _w14969_ ;
	wire _w14968_ ;
	wire _w14967_ ;
	wire _w14966_ ;
	wire _w14965_ ;
	wire _w14964_ ;
	wire _w14963_ ;
	wire _w14962_ ;
	wire _w14961_ ;
	wire _w14960_ ;
	wire _w14959_ ;
	wire _w14958_ ;
	wire _w14957_ ;
	wire _w14956_ ;
	wire _w14955_ ;
	wire _w14954_ ;
	wire _w14953_ ;
	wire _w14952_ ;
	wire _w14951_ ;
	wire _w14950_ ;
	wire _w14949_ ;
	wire _w14948_ ;
	wire _w14947_ ;
	wire _w14946_ ;
	wire _w14945_ ;
	wire _w14944_ ;
	wire _w14943_ ;
	wire _w14942_ ;
	wire _w14941_ ;
	wire _w14940_ ;
	wire _w14939_ ;
	wire _w14938_ ;
	wire _w14937_ ;
	wire _w14936_ ;
	wire _w14935_ ;
	wire _w14934_ ;
	wire _w14933_ ;
	wire _w14932_ ;
	wire _w14931_ ;
	wire _w14930_ ;
	wire _w14929_ ;
	wire _w14928_ ;
	wire _w14927_ ;
	wire _w14926_ ;
	wire _w14925_ ;
	wire _w14924_ ;
	wire _w14923_ ;
	wire _w14922_ ;
	wire _w14921_ ;
	wire _w14920_ ;
	wire _w14919_ ;
	wire _w14918_ ;
	wire _w14917_ ;
	wire _w14916_ ;
	wire _w14915_ ;
	wire _w14914_ ;
	wire _w14913_ ;
	wire _w14912_ ;
	wire _w14911_ ;
	wire _w14910_ ;
	wire _w14909_ ;
	wire _w14908_ ;
	wire _w14907_ ;
	wire _w14906_ ;
	wire _w14905_ ;
	wire _w14904_ ;
	wire _w14903_ ;
	wire _w14902_ ;
	wire _w14901_ ;
	wire _w14900_ ;
	wire _w14899_ ;
	wire _w14898_ ;
	wire _w14897_ ;
	wire _w14896_ ;
	wire _w14895_ ;
	wire _w14894_ ;
	wire _w14893_ ;
	wire _w14892_ ;
	wire _w14891_ ;
	wire _w14890_ ;
	wire _w14889_ ;
	wire _w14888_ ;
	wire _w14887_ ;
	wire _w14886_ ;
	wire _w14885_ ;
	wire _w14884_ ;
	wire _w14883_ ;
	wire _w14882_ ;
	wire _w14881_ ;
	wire _w14880_ ;
	wire _w14879_ ;
	wire _w14878_ ;
	wire _w14877_ ;
	wire _w14876_ ;
	wire _w14875_ ;
	wire _w14874_ ;
	wire _w14873_ ;
	wire _w14872_ ;
	wire _w14871_ ;
	wire _w14870_ ;
	wire _w14869_ ;
	wire _w14868_ ;
	wire _w14867_ ;
	wire _w14866_ ;
	wire _w14865_ ;
	wire _w14864_ ;
	wire _w14863_ ;
	wire _w14862_ ;
	wire _w14861_ ;
	wire _w14860_ ;
	wire _w14859_ ;
	wire _w14858_ ;
	wire _w14857_ ;
	wire _w14856_ ;
	wire _w14855_ ;
	wire _w14854_ ;
	wire _w14853_ ;
	wire _w14852_ ;
	wire _w14851_ ;
	wire _w14850_ ;
	wire _w14849_ ;
	wire _w14848_ ;
	wire _w14847_ ;
	wire _w14846_ ;
	wire _w14845_ ;
	wire _w14844_ ;
	wire _w14843_ ;
	wire _w14842_ ;
	wire _w14841_ ;
	wire _w14840_ ;
	wire _w14839_ ;
	wire _w14838_ ;
	wire _w14837_ ;
	wire _w14836_ ;
	wire _w14835_ ;
	wire _w14834_ ;
	wire _w14833_ ;
	wire _w14832_ ;
	wire _w14831_ ;
	wire _w14830_ ;
	wire _w14829_ ;
	wire _w14828_ ;
	wire _w14827_ ;
	wire _w14826_ ;
	wire _w14825_ ;
	wire _w14824_ ;
	wire _w14823_ ;
	wire _w14822_ ;
	wire _w14821_ ;
	wire _w14820_ ;
	wire _w14819_ ;
	wire _w14818_ ;
	wire _w14817_ ;
	wire _w14816_ ;
	wire _w14815_ ;
	wire _w14814_ ;
	wire _w14813_ ;
	wire _w14812_ ;
	wire _w14811_ ;
	wire _w14810_ ;
	wire _w14809_ ;
	wire _w14808_ ;
	wire _w14807_ ;
	wire _w14806_ ;
	wire _w14805_ ;
	wire _w14804_ ;
	wire _w14803_ ;
	wire _w14802_ ;
	wire _w14801_ ;
	wire _w14800_ ;
	wire _w14799_ ;
	wire _w14798_ ;
	wire _w14797_ ;
	wire _w14796_ ;
	wire _w14795_ ;
	wire _w14794_ ;
	wire _w14793_ ;
	wire _w14792_ ;
	wire _w14791_ ;
	wire _w14790_ ;
	wire _w14789_ ;
	wire _w14788_ ;
	wire _w14787_ ;
	wire _w14786_ ;
	wire _w14785_ ;
	wire _w14784_ ;
	wire _w14783_ ;
	wire _w14782_ ;
	wire _w14781_ ;
	wire _w14780_ ;
	wire _w14779_ ;
	wire _w14778_ ;
	wire _w14777_ ;
	wire _w14776_ ;
	wire _w14775_ ;
	wire _w14774_ ;
	wire _w14773_ ;
	wire _w14772_ ;
	wire _w14771_ ;
	wire _w14770_ ;
	wire _w14769_ ;
	wire _w14768_ ;
	wire _w14767_ ;
	wire _w14766_ ;
	wire _w14765_ ;
	wire _w14764_ ;
	wire _w14763_ ;
	wire _w14762_ ;
	wire _w14761_ ;
	wire _w14760_ ;
	wire _w14759_ ;
	wire _w14758_ ;
	wire _w14757_ ;
	wire _w14756_ ;
	wire _w14755_ ;
	wire _w14754_ ;
	wire _w14753_ ;
	wire _w14752_ ;
	wire _w14751_ ;
	wire _w14750_ ;
	wire _w14749_ ;
	wire _w14748_ ;
	wire _w14747_ ;
	wire _w14746_ ;
	wire _w14745_ ;
	wire _w14744_ ;
	wire _w14743_ ;
	wire _w14742_ ;
	wire _w14741_ ;
	wire _w14740_ ;
	wire _w14739_ ;
	wire _w14738_ ;
	wire _w14737_ ;
	wire _w14736_ ;
	wire _w14735_ ;
	wire _w14734_ ;
	wire _w14733_ ;
	wire _w14732_ ;
	wire _w14731_ ;
	wire _w14730_ ;
	wire _w14729_ ;
	wire _w14728_ ;
	wire _w14727_ ;
	wire _w14726_ ;
	wire _w14725_ ;
	wire _w14724_ ;
	wire _w14723_ ;
	wire _w14722_ ;
	wire _w14721_ ;
	wire _w14720_ ;
	wire _w14719_ ;
	wire _w14718_ ;
	wire _w14717_ ;
	wire _w14716_ ;
	wire _w14715_ ;
	wire _w14714_ ;
	wire _w14713_ ;
	wire _w14712_ ;
	wire _w14711_ ;
	wire _w14710_ ;
	wire _w14709_ ;
	wire _w14708_ ;
	wire _w14707_ ;
	wire _w14706_ ;
	wire _w14705_ ;
	wire _w14704_ ;
	wire _w14703_ ;
	wire _w14702_ ;
	wire _w14701_ ;
	wire _w14700_ ;
	wire _w14699_ ;
	wire _w14698_ ;
	wire _w14697_ ;
	wire _w14696_ ;
	wire _w14695_ ;
	wire _w14694_ ;
	wire _w14693_ ;
	wire _w14692_ ;
	wire _w14691_ ;
	wire _w14690_ ;
	wire _w14689_ ;
	wire _w14688_ ;
	wire _w14687_ ;
	wire _w14686_ ;
	wire _w14685_ ;
	wire _w14684_ ;
	wire _w14683_ ;
	wire _w14682_ ;
	wire _w14681_ ;
	wire _w14680_ ;
	wire _w14679_ ;
	wire _w14678_ ;
	wire _w14677_ ;
	wire _w14676_ ;
	wire _w14675_ ;
	wire _w14674_ ;
	wire _w14673_ ;
	wire _w14672_ ;
	wire _w14671_ ;
	wire _w14670_ ;
	wire _w14669_ ;
	wire _w14668_ ;
	wire _w14667_ ;
	wire _w14666_ ;
	wire _w14665_ ;
	wire _w14664_ ;
	wire _w14663_ ;
	wire _w14662_ ;
	wire _w14661_ ;
	wire _w14660_ ;
	wire _w14659_ ;
	wire _w14658_ ;
	wire _w14657_ ;
	wire _w14656_ ;
	wire _w14655_ ;
	wire _w14654_ ;
	wire _w14653_ ;
	wire _w14652_ ;
	wire _w14651_ ;
	wire _w14650_ ;
	wire _w14649_ ;
	wire _w14648_ ;
	wire _w14647_ ;
	wire _w14646_ ;
	wire _w14645_ ;
	wire _w14644_ ;
	wire _w14643_ ;
	wire _w14642_ ;
	wire _w14641_ ;
	wire _w14640_ ;
	wire _w14639_ ;
	wire _w14638_ ;
	wire _w14637_ ;
	wire _w14636_ ;
	wire _w14635_ ;
	wire _w14634_ ;
	wire _w14633_ ;
	wire _w14632_ ;
	wire _w14631_ ;
	wire _w14630_ ;
	wire _w14629_ ;
	wire _w14628_ ;
	wire _w14627_ ;
	wire _w14626_ ;
	wire _w14625_ ;
	wire _w14624_ ;
	wire _w14623_ ;
	wire _w14622_ ;
	wire _w14621_ ;
	wire _w14620_ ;
	wire _w14619_ ;
	wire _w14618_ ;
	wire _w14617_ ;
	wire _w14616_ ;
	wire _w14615_ ;
	wire _w14614_ ;
	wire _w14613_ ;
	wire _w14612_ ;
	wire _w14611_ ;
	wire _w14610_ ;
	wire _w14609_ ;
	wire _w14608_ ;
	wire _w14607_ ;
	wire _w14606_ ;
	wire _w14605_ ;
	wire _w14604_ ;
	wire _w14603_ ;
	wire _w14602_ ;
	wire _w14601_ ;
	wire _w14600_ ;
	wire _w14599_ ;
	wire _w14598_ ;
	wire _w14597_ ;
	wire _w14596_ ;
	wire _w14595_ ;
	wire _w14594_ ;
	wire _w14593_ ;
	wire _w14592_ ;
	wire _w14591_ ;
	wire _w14590_ ;
	wire _w14589_ ;
	wire _w14588_ ;
	wire _w14587_ ;
	wire _w14586_ ;
	wire _w14585_ ;
	wire _w14584_ ;
	wire _w14583_ ;
	wire _w14582_ ;
	wire _w14581_ ;
	wire _w14580_ ;
	wire _w14579_ ;
	wire _w14578_ ;
	wire _w14577_ ;
	wire _w14576_ ;
	wire _w14575_ ;
	wire _w14574_ ;
	wire _w14573_ ;
	wire _w14572_ ;
	wire _w14571_ ;
	wire _w14570_ ;
	wire _w14569_ ;
	wire _w14568_ ;
	wire _w14567_ ;
	wire _w14566_ ;
	wire _w14565_ ;
	wire _w14564_ ;
	wire _w14563_ ;
	wire _w14562_ ;
	wire _w14561_ ;
	wire _w14560_ ;
	wire _w14559_ ;
	wire _w14558_ ;
	wire _w14557_ ;
	wire _w14556_ ;
	wire _w14555_ ;
	wire _w14554_ ;
	wire _w14553_ ;
	wire _w14552_ ;
	wire _w14551_ ;
	wire _w14550_ ;
	wire _w14549_ ;
	wire _w14548_ ;
	wire _w14547_ ;
	wire _w14546_ ;
	wire _w14545_ ;
	wire _w14544_ ;
	wire _w14543_ ;
	wire _w14542_ ;
	wire _w14541_ ;
	wire _w14540_ ;
	wire _w14539_ ;
	wire _w14538_ ;
	wire _w14537_ ;
	wire _w14536_ ;
	wire _w14535_ ;
	wire _w14534_ ;
	wire _w14533_ ;
	wire _w14532_ ;
	wire _w14531_ ;
	wire _w14530_ ;
	wire _w14529_ ;
	wire _w14528_ ;
	wire _w14527_ ;
	wire _w14526_ ;
	wire _w14525_ ;
	wire _w14524_ ;
	wire _w14523_ ;
	wire _w14522_ ;
	wire _w14521_ ;
	wire _w14520_ ;
	wire _w14519_ ;
	wire _w14518_ ;
	wire _w14517_ ;
	wire _w14516_ ;
	wire _w14515_ ;
	wire _w14514_ ;
	wire _w14513_ ;
	wire _w14512_ ;
	wire _w14511_ ;
	wire _w14510_ ;
	wire _w14509_ ;
	wire _w14508_ ;
	wire _w14507_ ;
	wire _w14506_ ;
	wire _w14505_ ;
	wire _w14504_ ;
	wire _w14503_ ;
	wire _w14502_ ;
	wire _w14501_ ;
	wire _w14500_ ;
	wire _w14499_ ;
	wire _w14498_ ;
	wire _w14497_ ;
	wire _w14496_ ;
	wire _w14495_ ;
	wire _w14494_ ;
	wire _w14493_ ;
	wire _w14492_ ;
	wire _w14491_ ;
	wire _w14490_ ;
	wire _w14489_ ;
	wire _w14488_ ;
	wire _w14487_ ;
	wire _w14486_ ;
	wire _w14485_ ;
	wire _w14484_ ;
	wire _w14483_ ;
	wire _w14482_ ;
	wire _w14481_ ;
	wire _w14480_ ;
	wire _w14479_ ;
	wire _w14478_ ;
	wire _w14477_ ;
	wire _w14476_ ;
	wire _w14475_ ;
	wire _w14474_ ;
	wire _w14473_ ;
	wire _w14472_ ;
	wire _w14471_ ;
	wire _w14470_ ;
	wire _w14469_ ;
	wire _w14468_ ;
	wire _w14467_ ;
	wire _w14466_ ;
	wire _w14465_ ;
	wire _w14464_ ;
	wire _w14463_ ;
	wire _w14462_ ;
	wire _w14461_ ;
	wire _w14460_ ;
	wire _w14459_ ;
	wire _w14458_ ;
	wire _w14457_ ;
	wire _w14456_ ;
	wire _w14455_ ;
	wire _w14454_ ;
	wire _w14453_ ;
	wire _w14452_ ;
	wire _w14451_ ;
	wire _w14450_ ;
	wire _w14449_ ;
	wire _w14448_ ;
	wire _w14447_ ;
	wire _w14446_ ;
	wire _w14445_ ;
	wire _w14444_ ;
	wire _w14443_ ;
	wire _w14442_ ;
	wire _w14441_ ;
	wire _w14440_ ;
	wire _w14439_ ;
	wire _w14438_ ;
	wire _w14437_ ;
	wire _w14436_ ;
	wire _w14435_ ;
	wire _w14434_ ;
	wire _w14433_ ;
	wire _w14432_ ;
	wire _w14431_ ;
	wire _w14430_ ;
	wire _w14429_ ;
	wire _w14428_ ;
	wire _w14427_ ;
	wire _w14426_ ;
	wire _w14425_ ;
	wire _w14424_ ;
	wire _w14423_ ;
	wire _w14422_ ;
	wire _w14421_ ;
	wire _w14420_ ;
	wire _w14419_ ;
	wire _w14418_ ;
	wire _w14417_ ;
	wire _w14416_ ;
	wire _w14415_ ;
	wire _w14414_ ;
	wire _w14413_ ;
	wire _w14412_ ;
	wire _w14411_ ;
	wire _w14410_ ;
	wire _w14409_ ;
	wire _w14408_ ;
	wire _w14407_ ;
	wire _w14406_ ;
	wire _w14405_ ;
	wire _w14404_ ;
	wire _w14403_ ;
	wire _w14402_ ;
	wire _w14401_ ;
	wire _w14400_ ;
	wire _w14399_ ;
	wire _w14398_ ;
	wire _w14397_ ;
	wire _w14396_ ;
	wire _w14395_ ;
	wire _w14394_ ;
	wire _w14393_ ;
	wire _w14392_ ;
	wire _w14391_ ;
	wire _w14390_ ;
	wire _w14389_ ;
	wire _w14388_ ;
	wire _w14387_ ;
	wire _w14386_ ;
	wire _w14385_ ;
	wire _w14384_ ;
	wire _w14383_ ;
	wire _w14382_ ;
	wire _w14381_ ;
	wire _w14380_ ;
	wire _w14379_ ;
	wire _w14378_ ;
	wire _w14377_ ;
	wire _w14376_ ;
	wire _w14375_ ;
	wire _w14374_ ;
	wire _w14373_ ;
	wire _w14372_ ;
	wire _w14371_ ;
	wire _w14370_ ;
	wire _w14369_ ;
	wire _w14368_ ;
	wire _w14367_ ;
	wire _w14366_ ;
	wire _w14365_ ;
	wire _w14364_ ;
	wire _w14363_ ;
	wire _w14362_ ;
	wire _w14361_ ;
	wire _w14360_ ;
	wire _w14359_ ;
	wire _w14358_ ;
	wire _w14357_ ;
	wire _w14356_ ;
	wire _w14355_ ;
	wire _w14354_ ;
	wire _w14353_ ;
	wire _w14352_ ;
	wire _w14351_ ;
	wire _w14350_ ;
	wire _w14349_ ;
	wire _w14348_ ;
	wire _w14347_ ;
	wire _w14346_ ;
	wire _w14345_ ;
	wire _w14344_ ;
	wire _w14343_ ;
	wire _w14342_ ;
	wire _w14341_ ;
	wire _w14340_ ;
	wire _w14339_ ;
	wire _w14338_ ;
	wire _w14337_ ;
	wire _w14336_ ;
	wire _w14335_ ;
	wire _w14334_ ;
	wire _w14333_ ;
	wire _w14332_ ;
	wire _w14331_ ;
	wire _w14330_ ;
	wire _w14329_ ;
	wire _w14328_ ;
	wire _w14327_ ;
	wire _w14326_ ;
	wire _w14325_ ;
	wire _w14324_ ;
	wire _w14323_ ;
	wire _w14322_ ;
	wire _w14321_ ;
	wire _w14320_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	wire _w10735_ ;
	wire _w10736_ ;
	wire _w10737_ ;
	wire _w10738_ ;
	wire _w10739_ ;
	wire _w10740_ ;
	wire _w10741_ ;
	wire _w10742_ ;
	wire _w10743_ ;
	wire _w10744_ ;
	wire _w10745_ ;
	wire _w10746_ ;
	wire _w10747_ ;
	wire _w10748_ ;
	wire _w10749_ ;
	wire _w10750_ ;
	wire _w10751_ ;
	wire _w10752_ ;
	wire _w10753_ ;
	wire _w10754_ ;
	wire _w10755_ ;
	wire _w10756_ ;
	wire _w10757_ ;
	wire _w10758_ ;
	wire _w10759_ ;
	wire _w10760_ ;
	wire _w10761_ ;
	wire _w10762_ ;
	wire _w10763_ ;
	wire _w10764_ ;
	wire _w10765_ ;
	wire _w10766_ ;
	wire _w10767_ ;
	wire _w10768_ ;
	wire _w10769_ ;
	wire _w10770_ ;
	wire _w10771_ ;
	wire _w10772_ ;
	wire _w10773_ ;
	wire _w10774_ ;
	wire _w10775_ ;
	wire _w10776_ ;
	wire _w10777_ ;
	wire _w10778_ ;
	wire _w10779_ ;
	wire _w10780_ ;
	wire _w10781_ ;
	wire _w10782_ ;
	wire _w10783_ ;
	wire _w10784_ ;
	wire _w10785_ ;
	wire _w10786_ ;
	wire _w10787_ ;
	wire _w10788_ ;
	wire _w10789_ ;
	wire _w10790_ ;
	wire _w10791_ ;
	wire _w10792_ ;
	wire _w10793_ ;
	wire _w10794_ ;
	wire _w10795_ ;
	wire _w10796_ ;
	wire _w10797_ ;
	wire _w10798_ ;
	wire _w10799_ ;
	wire _w10800_ ;
	wire _w10801_ ;
	wire _w10802_ ;
	wire _w10803_ ;
	wire _w10804_ ;
	wire _w10805_ ;
	wire _w10806_ ;
	wire _w10807_ ;
	wire _w10808_ ;
	wire _w10809_ ;
	wire _w10810_ ;
	wire _w10811_ ;
	wire _w10812_ ;
	wire _w10813_ ;
	wire _w10814_ ;
	wire _w10815_ ;
	wire _w10816_ ;
	wire _w10817_ ;
	wire _w10818_ ;
	wire _w10819_ ;
	wire _w10820_ ;
	wire _w10821_ ;
	wire _w10822_ ;
	wire _w10823_ ;
	wire _w10824_ ;
	wire _w10825_ ;
	wire _w10826_ ;
	wire _w10827_ ;
	wire _w10828_ ;
	wire _w10829_ ;
	wire _w10830_ ;
	wire _w10831_ ;
	wire _w10832_ ;
	wire _w10833_ ;
	wire _w10834_ ;
	wire _w10835_ ;
	wire _w10836_ ;
	wire _w10837_ ;
	wire _w10838_ ;
	wire _w10839_ ;
	wire _w10840_ ;
	wire _w10841_ ;
	wire _w10842_ ;
	wire _w10843_ ;
	wire _w10844_ ;
	wire _w10845_ ;
	wire _w10846_ ;
	wire _w10847_ ;
	wire _w10848_ ;
	wire _w10849_ ;
	wire _w10850_ ;
	wire _w10851_ ;
	wire _w10852_ ;
	wire _w10853_ ;
	wire _w10854_ ;
	wire _w10855_ ;
	wire _w10856_ ;
	wire _w10857_ ;
	wire _w10858_ ;
	wire _w10859_ ;
	wire _w10860_ ;
	wire _w10861_ ;
	wire _w10862_ ;
	wire _w10863_ ;
	wire _w10864_ ;
	wire _w10865_ ;
	wire _w10866_ ;
	wire _w10867_ ;
	wire _w10868_ ;
	wire _w10869_ ;
	wire _w10870_ ;
	wire _w10871_ ;
	wire _w10872_ ;
	wire _w10873_ ;
	wire _w10874_ ;
	wire _w10875_ ;
	wire _w10876_ ;
	wire _w10877_ ;
	wire _w10878_ ;
	wire _w10879_ ;
	wire _w10880_ ;
	wire _w10881_ ;
	wire _w10882_ ;
	wire _w10883_ ;
	wire _w10884_ ;
	wire _w10885_ ;
	wire _w10886_ ;
	wire _w10887_ ;
	wire _w10888_ ;
	wire _w10889_ ;
	wire _w10890_ ;
	wire _w10891_ ;
	wire _w10892_ ;
	wire _w10893_ ;
	wire _w10894_ ;
	wire _w10895_ ;
	wire _w10896_ ;
	wire _w10897_ ;
	wire _w10898_ ;
	wire _w10899_ ;
	wire _w10900_ ;
	wire _w10901_ ;
	wire _w10902_ ;
	wire _w10903_ ;
	wire _w10904_ ;
	wire _w10905_ ;
	wire _w10906_ ;
	wire _w10907_ ;
	wire _w10908_ ;
	wire _w10909_ ;
	wire _w10910_ ;
	wire _w10911_ ;
	wire _w10912_ ;
	wire _w10913_ ;
	wire _w10914_ ;
	wire _w10915_ ;
	wire _w10916_ ;
	wire _w10917_ ;
	wire _w10918_ ;
	wire _w10919_ ;
	wire _w10920_ ;
	wire _w10921_ ;
	wire _w10922_ ;
	wire _w10923_ ;
	wire _w10924_ ;
	wire _w10925_ ;
	wire _w10926_ ;
	wire _w10927_ ;
	wire _w10928_ ;
	wire _w10929_ ;
	wire _w10930_ ;
	wire _w10931_ ;
	wire _w10932_ ;
	wire _w10933_ ;
	wire _w10934_ ;
	wire _w10935_ ;
	wire _w10936_ ;
	wire _w10937_ ;
	wire _w10938_ ;
	wire _w10939_ ;
	wire _w10940_ ;
	wire _w10941_ ;
	wire _w10942_ ;
	wire _w10943_ ;
	wire _w10944_ ;
	wire _w10945_ ;
	wire _w10946_ ;
	wire _w10947_ ;
	wire _w10948_ ;
	wire _w10949_ ;
	wire _w10950_ ;
	wire _w10951_ ;
	wire _w10952_ ;
	wire _w10953_ ;
	wire _w10954_ ;
	wire _w10955_ ;
	wire _w10956_ ;
	wire _w10957_ ;
	wire _w10958_ ;
	wire _w10959_ ;
	wire _w10960_ ;
	wire _w10961_ ;
	wire _w10962_ ;
	wire _w10963_ ;
	wire _w10964_ ;
	wire _w10965_ ;
	wire _w10966_ ;
	wire _w10967_ ;
	wire _w10968_ ;
	wire _w10969_ ;
	wire _w10970_ ;
	wire _w10971_ ;
	wire _w10972_ ;
	wire _w10973_ ;
	wire _w10974_ ;
	wire _w10975_ ;
	wire _w10976_ ;
	wire _w10977_ ;
	wire _w10978_ ;
	wire _w10979_ ;
	wire _w10980_ ;
	wire _w10981_ ;
	wire _w10982_ ;
	wire _w10983_ ;
	wire _w10984_ ;
	wire _w10985_ ;
	wire _w10986_ ;
	wire _w10987_ ;
	wire _w10988_ ;
	wire _w10989_ ;
	wire _w10990_ ;
	wire _w10991_ ;
	wire _w10992_ ;
	wire _w10993_ ;
	wire _w10994_ ;
	wire _w10995_ ;
	wire _w10996_ ;
	wire _w10997_ ;
	wire _w10998_ ;
	wire _w10999_ ;
	wire _w11000_ ;
	wire _w11001_ ;
	wire _w11002_ ;
	wire _w11003_ ;
	wire _w11004_ ;
	wire _w11005_ ;
	wire _w11006_ ;
	wire _w11007_ ;
	wire _w11008_ ;
	wire _w11009_ ;
	wire _w11010_ ;
	wire _w11011_ ;
	wire _w11012_ ;
	wire _w11013_ ;
	wire _w11014_ ;
	wire _w11015_ ;
	wire _w11016_ ;
	wire _w11017_ ;
	wire _w11018_ ;
	wire _w11019_ ;
	wire _w11020_ ;
	wire _w11021_ ;
	wire _w11022_ ;
	wire _w11023_ ;
	wire _w11024_ ;
	wire _w11025_ ;
	wire _w11026_ ;
	wire _w11027_ ;
	wire _w11028_ ;
	wire _w11029_ ;
	wire _w11030_ ;
	wire _w11031_ ;
	wire _w11032_ ;
	wire _w11033_ ;
	wire _w11034_ ;
	wire _w11035_ ;
	wire _w11036_ ;
	wire _w11037_ ;
	wire _w11038_ ;
	wire _w11039_ ;
	wire _w11040_ ;
	wire _w11041_ ;
	wire _w11042_ ;
	wire _w11043_ ;
	wire _w11044_ ;
	wire _w11045_ ;
	wire _w11046_ ;
	wire _w11047_ ;
	wire _w11048_ ;
	wire _w11049_ ;
	wire _w11050_ ;
	wire _w11051_ ;
	wire _w11052_ ;
	wire _w11053_ ;
	wire _w11054_ ;
	wire _w11055_ ;
	wire _w11056_ ;
	wire _w11057_ ;
	wire _w11058_ ;
	wire _w11059_ ;
	wire _w11060_ ;
	wire _w11061_ ;
	wire _w11062_ ;
	wire _w11063_ ;
	wire _w11064_ ;
	wire _w11065_ ;
	wire _w11066_ ;
	wire _w11067_ ;
	wire _w11068_ ;
	wire _w11069_ ;
	wire _w11070_ ;
	wire _w11071_ ;
	wire _w11072_ ;
	wire _w11073_ ;
	wire _w11074_ ;
	wire _w11075_ ;
	wire _w11076_ ;
	wire _w11077_ ;
	wire _w11078_ ;
	wire _w11079_ ;
	wire _w11080_ ;
	wire _w11081_ ;
	wire _w11082_ ;
	wire _w11083_ ;
	wire _w11084_ ;
	wire _w11085_ ;
	wire _w11086_ ;
	wire _w11087_ ;
	wire _w11088_ ;
	wire _w11089_ ;
	wire _w11090_ ;
	wire _w11091_ ;
	wire _w11092_ ;
	wire _w11093_ ;
	wire _w11094_ ;
	wire _w11095_ ;
	wire _w11096_ ;
	wire _w11097_ ;
	wire _w11098_ ;
	wire _w11099_ ;
	wire _w11100_ ;
	wire _w11101_ ;
	wire _w11102_ ;
	wire _w11103_ ;
	wire _w11104_ ;
	wire _w11105_ ;
	wire _w11106_ ;
	wire _w11107_ ;
	wire _w11108_ ;
	wire _w11109_ ;
	wire _w11110_ ;
	wire _w11111_ ;
	wire _w11112_ ;
	wire _w11113_ ;
	wire _w11114_ ;
	wire _w11115_ ;
	wire _w11116_ ;
	wire _w11117_ ;
	wire _w11118_ ;
	wire _w11119_ ;
	wire _w11120_ ;
	wire _w11121_ ;
	wire _w11122_ ;
	wire _w11123_ ;
	wire _w11124_ ;
	wire _w11125_ ;
	wire _w11126_ ;
	wire _w11127_ ;
	wire _w11128_ ;
	wire _w11129_ ;
	wire _w11130_ ;
	wire _w11131_ ;
	wire _w11132_ ;
	wire _w11133_ ;
	wire _w11134_ ;
	wire _w11135_ ;
	wire _w11136_ ;
	wire _w11137_ ;
	wire _w11138_ ;
	wire _w11139_ ;
	wire _w11140_ ;
	wire _w11141_ ;
	wire _w11142_ ;
	wire _w11143_ ;
	wire _w11144_ ;
	wire _w11145_ ;
	wire _w11146_ ;
	wire _w11147_ ;
	wire _w11148_ ;
	wire _w11149_ ;
	wire _w11150_ ;
	wire _w11151_ ;
	wire _w11152_ ;
	wire _w11153_ ;
	wire _w11154_ ;
	wire _w11155_ ;
	wire _w11156_ ;
	wire _w11157_ ;
	wire _w11158_ ;
	wire _w11159_ ;
	wire _w11160_ ;
	wire _w11161_ ;
	wire _w11162_ ;
	wire _w11163_ ;
	wire _w11164_ ;
	wire _w11165_ ;
	wire _w11166_ ;
	wire _w11167_ ;
	wire _w11168_ ;
	wire _w11169_ ;
	wire _w11170_ ;
	wire _w11171_ ;
	wire _w11172_ ;
	wire _w11173_ ;
	wire _w11174_ ;
	wire _w11175_ ;
	wire _w11176_ ;
	wire _w11177_ ;
	wire _w11178_ ;
	wire _w11179_ ;
	wire _w11180_ ;
	wire _w11181_ ;
	wire _w11182_ ;
	wire _w11183_ ;
	wire _w11184_ ;
	wire _w11185_ ;
	wire _w11186_ ;
	wire _w11187_ ;
	wire _w11188_ ;
	wire _w11189_ ;
	wire _w11190_ ;
	wire _w11191_ ;
	wire _w11192_ ;
	wire _w11193_ ;
	wire _w11194_ ;
	wire _w11195_ ;
	wire _w11196_ ;
	wire _w11197_ ;
	wire _w11198_ ;
	wire _w11199_ ;
	wire _w11200_ ;
	wire _w11201_ ;
	wire _w11202_ ;
	wire _w11203_ ;
	wire _w11204_ ;
	wire _w11205_ ;
	wire _w11206_ ;
	wire _w11207_ ;
	wire _w11208_ ;
	wire _w11209_ ;
	wire _w11210_ ;
	wire _w11211_ ;
	wire _w11212_ ;
	wire _w11213_ ;
	wire _w11214_ ;
	wire _w11215_ ;
	wire _w11216_ ;
	wire _w11217_ ;
	wire _w11218_ ;
	wire _w11219_ ;
	wire _w11220_ ;
	wire _w11221_ ;
	wire _w11222_ ;
	wire _w11223_ ;
	wire _w11224_ ;
	wire _w11225_ ;
	wire _w11226_ ;
	wire _w11227_ ;
	wire _w11228_ ;
	wire _w11229_ ;
	wire _w11230_ ;
	wire _w11231_ ;
	wire _w11232_ ;
	wire _w11233_ ;
	wire _w11234_ ;
	wire _w11235_ ;
	wire _w11236_ ;
	wire _w11237_ ;
	wire _w11238_ ;
	wire _w11239_ ;
	wire _w11240_ ;
	wire _w11241_ ;
	wire _w11242_ ;
	wire _w11243_ ;
	wire _w11244_ ;
	wire _w11245_ ;
	wire _w11246_ ;
	wire _w11247_ ;
	wire _w11248_ ;
	wire _w11249_ ;
	wire _w11250_ ;
	wire _w11251_ ;
	wire _w11252_ ;
	wire _w11253_ ;
	wire _w11254_ ;
	wire _w11255_ ;
	wire _w11256_ ;
	wire _w11257_ ;
	wire _w11258_ ;
	wire _w11259_ ;
	wire _w11260_ ;
	wire _w11261_ ;
	wire _w11262_ ;
	wire _w11263_ ;
	wire _w11264_ ;
	wire _w11265_ ;
	wire _w11266_ ;
	wire _w11267_ ;
	wire _w11268_ ;
	wire _w11269_ ;
	wire _w11270_ ;
	wire _w11271_ ;
	wire _w11272_ ;
	wire _w11273_ ;
	wire _w11274_ ;
	wire _w11275_ ;
	wire _w11276_ ;
	wire _w11277_ ;
	wire _w11278_ ;
	wire _w11279_ ;
	wire _w11280_ ;
	wire _w11281_ ;
	wire _w11282_ ;
	wire _w11283_ ;
	wire _w11284_ ;
	wire _w11285_ ;
	wire _w11286_ ;
	wire _w11287_ ;
	wire _w11288_ ;
	wire _w11289_ ;
	wire _w11290_ ;
	wire _w11291_ ;
	wire _w11292_ ;
	wire _w11293_ ;
	wire _w11294_ ;
	wire _w11295_ ;
	wire _w11296_ ;
	wire _w11297_ ;
	wire _w11298_ ;
	wire _w11299_ ;
	wire _w11300_ ;
	wire _w11301_ ;
	wire _w11302_ ;
	wire _w11303_ ;
	wire _w11304_ ;
	wire _w11305_ ;
	wire _w11306_ ;
	wire _w11307_ ;
	wire _w11308_ ;
	wire _w11309_ ;
	wire _w11310_ ;
	wire _w11311_ ;
	wire _w11312_ ;
	wire _w11313_ ;
	wire _w11314_ ;
	wire _w11315_ ;
	wire _w11316_ ;
	wire _w11317_ ;
	wire _w11318_ ;
	wire _w11319_ ;
	wire _w11320_ ;
	wire _w11321_ ;
	wire _w11322_ ;
	wire _w11323_ ;
	wire _w11324_ ;
	wire _w11325_ ;
	wire _w11326_ ;
	wire _w11327_ ;
	wire _w11328_ ;
	wire _w11329_ ;
	wire _w11330_ ;
	wire _w11331_ ;
	wire _w11332_ ;
	wire _w11333_ ;
	wire _w11334_ ;
	wire _w11335_ ;
	wire _w11336_ ;
	wire _w11337_ ;
	wire _w11338_ ;
	wire _w11339_ ;
	wire _w11340_ ;
	wire _w11341_ ;
	wire _w11342_ ;
	wire _w11343_ ;
	wire _w11344_ ;
	wire _w11345_ ;
	wire _w11346_ ;
	wire _w11347_ ;
	wire _w11348_ ;
	wire _w11349_ ;
	wire _w11350_ ;
	wire _w11351_ ;
	wire _w11352_ ;
	wire _w11353_ ;
	wire _w11354_ ;
	wire _w11355_ ;
	wire _w11356_ ;
	wire _w11357_ ;
	wire _w11358_ ;
	wire _w11359_ ;
	wire _w11360_ ;
	wire _w11361_ ;
	wire _w11362_ ;
	wire _w11363_ ;
	wire _w11364_ ;
	wire _w11365_ ;
	wire _w11366_ ;
	wire _w11367_ ;
	wire _w11368_ ;
	wire _w11369_ ;
	wire _w11370_ ;
	wire _w11371_ ;
	wire _w11372_ ;
	wire _w11373_ ;
	wire _w11374_ ;
	wire _w11375_ ;
	wire _w11376_ ;
	wire _w11377_ ;
	wire _w11378_ ;
	wire _w11379_ ;
	wire _w11380_ ;
	wire _w11381_ ;
	wire _w11382_ ;
	wire _w11383_ ;
	wire _w11384_ ;
	wire _w11385_ ;
	wire _w11386_ ;
	wire _w11387_ ;
	wire _w11388_ ;
	wire _w11389_ ;
	wire _w11390_ ;
	wire _w11391_ ;
	wire _w11392_ ;
	wire _w11393_ ;
	wire _w11394_ ;
	wire _w11395_ ;
	wire _w11396_ ;
	wire _w11397_ ;
	wire _w11398_ ;
	wire _w11399_ ;
	wire _w11400_ ;
	wire _w11401_ ;
	wire _w11402_ ;
	wire _w11403_ ;
	wire _w11404_ ;
	wire _w11405_ ;
	wire _w11406_ ;
	wire _w11407_ ;
	wire _w11408_ ;
	wire _w11409_ ;
	wire _w11410_ ;
	wire _w11411_ ;
	wire _w11412_ ;
	wire _w11413_ ;
	wire _w11414_ ;
	wire _w11415_ ;
	wire _w11416_ ;
	wire _w11417_ ;
	wire _w11418_ ;
	wire _w11419_ ;
	wire _w11420_ ;
	wire _w11421_ ;
	wire _w11422_ ;
	wire _w11423_ ;
	wire _w11424_ ;
	wire _w11425_ ;
	wire _w11426_ ;
	wire _w11427_ ;
	wire _w11428_ ;
	wire _w11429_ ;
	wire _w11430_ ;
	wire _w11431_ ;
	wire _w11432_ ;
	wire _w11433_ ;
	wire _w11434_ ;
	wire _w11435_ ;
	wire _w11436_ ;
	wire _w11437_ ;
	wire _w11438_ ;
	wire _w11439_ ;
	wire _w11440_ ;
	wire _w11441_ ;
	wire _w11442_ ;
	wire _w11443_ ;
	wire _w11444_ ;
	wire _w11445_ ;
	wire _w11446_ ;
	wire _w11447_ ;
	wire _w11448_ ;
	wire _w11449_ ;
	wire _w11450_ ;
	wire _w11451_ ;
	wire _w11452_ ;
	wire _w11453_ ;
	wire _w11454_ ;
	wire _w11455_ ;
	wire _w11456_ ;
	wire _w11457_ ;
	wire _w11458_ ;
	wire _w11459_ ;
	wire _w11460_ ;
	wire _w11461_ ;
	wire _w11462_ ;
	wire _w11463_ ;
	wire _w11464_ ;
	wire _w11465_ ;
	wire _w11466_ ;
	wire _w11467_ ;
	wire _w11468_ ;
	wire _w11469_ ;
	wire _w11470_ ;
	wire _w11471_ ;
	wire _w11472_ ;
	wire _w11473_ ;
	wire _w11474_ ;
	wire _w11475_ ;
	wire _w11476_ ;
	wire _w11477_ ;
	wire _w11478_ ;
	wire _w11479_ ;
	wire _w11480_ ;
	wire _w11481_ ;
	wire _w11482_ ;
	wire _w11483_ ;
	wire _w11484_ ;
	wire _w11485_ ;
	wire _w11486_ ;
	wire _w11487_ ;
	wire _w11488_ ;
	wire _w11489_ ;
	wire _w11490_ ;
	wire _w11491_ ;
	wire _w11492_ ;
	wire _w11493_ ;
	wire _w11494_ ;
	wire _w11495_ ;
	wire _w11496_ ;
	wire _w11497_ ;
	wire _w11498_ ;
	wire _w11499_ ;
	wire _w11500_ ;
	wire _w11501_ ;
	wire _w11502_ ;
	wire _w11503_ ;
	wire _w11504_ ;
	wire _w11505_ ;
	wire _w11506_ ;
	wire _w11507_ ;
	wire _w11508_ ;
	wire _w11509_ ;
	wire _w11510_ ;
	wire _w11511_ ;
	wire _w11512_ ;
	wire _w11513_ ;
	wire _w11514_ ;
	wire _w11515_ ;
	wire _w11516_ ;
	wire _w11517_ ;
	wire _w11518_ ;
	wire _w11519_ ;
	wire _w11520_ ;
	wire _w11521_ ;
	wire _w11522_ ;
	wire _w11523_ ;
	wire _w11524_ ;
	wire _w11525_ ;
	wire _w11526_ ;
	wire _w11527_ ;
	wire _w11528_ ;
	wire _w11529_ ;
	wire _w11530_ ;
	wire _w11531_ ;
	wire _w11532_ ;
	wire _w11533_ ;
	wire _w11534_ ;
	wire _w11535_ ;
	wire _w11536_ ;
	wire _w11537_ ;
	wire _w11538_ ;
	wire _w11539_ ;
	wire _w11540_ ;
	wire _w11541_ ;
	wire _w11542_ ;
	wire _w11543_ ;
	wire _w11544_ ;
	wire _w11545_ ;
	wire _w11546_ ;
	wire _w11547_ ;
	wire _w11548_ ;
	wire _w11549_ ;
	wire _w11550_ ;
	wire _w11551_ ;
	wire _w11552_ ;
	wire _w11553_ ;
	wire _w11554_ ;
	wire _w11555_ ;
	wire _w11556_ ;
	wire _w11557_ ;
	wire _w11558_ ;
	wire _w11559_ ;
	wire _w11560_ ;
	wire _w11561_ ;
	wire _w11562_ ;
	wire _w11563_ ;
	wire _w11564_ ;
	wire _w11565_ ;
	wire _w11566_ ;
	wire _w11567_ ;
	wire _w11568_ ;
	wire _w11569_ ;
	wire _w11570_ ;
	wire _w11571_ ;
	wire _w11572_ ;
	wire _w11573_ ;
	wire _w11574_ ;
	wire _w11575_ ;
	wire _w11576_ ;
	wire _w11577_ ;
	wire _w11578_ ;
	wire _w11579_ ;
	wire _w11580_ ;
	wire _w11581_ ;
	wire _w11582_ ;
	wire _w11583_ ;
	wire _w11584_ ;
	wire _w11585_ ;
	wire _w11586_ ;
	wire _w11587_ ;
	wire _w11588_ ;
	wire _w11589_ ;
	wire _w11590_ ;
	wire _w11591_ ;
	wire _w11592_ ;
	wire _w11593_ ;
	wire _w11594_ ;
	wire _w11595_ ;
	wire _w11596_ ;
	wire _w11597_ ;
	wire _w11598_ ;
	wire _w11599_ ;
	wire _w11600_ ;
	wire _w11601_ ;
	wire _w11602_ ;
	wire _w11603_ ;
	wire _w11604_ ;
	wire _w11605_ ;
	wire _w11606_ ;
	wire _w11607_ ;
	wire _w11608_ ;
	wire _w11609_ ;
	wire _w11610_ ;
	wire _w11611_ ;
	wire _w11612_ ;
	wire _w11613_ ;
	wire _w11614_ ;
	wire _w11615_ ;
	wire _w11616_ ;
	wire _w11617_ ;
	wire _w11618_ ;
	wire _w11619_ ;
	wire _w11620_ ;
	wire _w11621_ ;
	wire _w11622_ ;
	LUT4 #(
		.INIT('hccc8)
	) name0 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[0]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1350_
	);
	LUT4 #(
		.INIT('h0010)
	) name1 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[0]/NET0131 ,
		\datao[30]_pad ,
		_w1351_
	);
	LUT2 #(
		.INIT('he)
	) name2 (
		_w1350_,
		_w1351_,
		_w1352_
	);
	LUT4 #(
		.INIT('hccc8)
	) name3 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[10]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1353_
	);
	LUT4 #(
		.INIT('h0010)
	) name4 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[10]/NET0131 ,
		\datao[30]_pad ,
		_w1354_
	);
	LUT2 #(
		.INIT('he)
	) name5 (
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('hccc8)
	) name6 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[11]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1356_
	);
	LUT4 #(
		.INIT('h0010)
	) name7 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[11]/NET0131 ,
		\datao[30]_pad ,
		_w1357_
	);
	LUT2 #(
		.INIT('he)
	) name8 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[12]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1359_
	);
	LUT4 #(
		.INIT('h0010)
	) name10 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[12]/NET0131 ,
		\datao[30]_pad ,
		_w1360_
	);
	LUT2 #(
		.INIT('he)
	) name11 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('hccc8)
	) name12 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[13]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1362_
	);
	LUT4 #(
		.INIT('h0010)
	) name13 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[13]/NET0131 ,
		\datao[30]_pad ,
		_w1363_
	);
	LUT2 #(
		.INIT('he)
	) name14 (
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('hccc8)
	) name15 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[14]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1365_
	);
	LUT4 #(
		.INIT('h0010)
	) name16 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[14]/NET0131 ,
		\datao[30]_pad ,
		_w1366_
	);
	LUT2 #(
		.INIT('he)
	) name17 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT4 #(
		.INIT('hccc8)
	) name18 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[15]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1368_
	);
	LUT4 #(
		.INIT('h0010)
	) name19 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[15]/NET0131 ,
		\datao[30]_pad ,
		_w1369_
	);
	LUT2 #(
		.INIT('he)
	) name20 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT4 #(
		.INIT('hccc8)
	) name21 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[16]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1371_
	);
	LUT4 #(
		.INIT('h0010)
	) name22 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[16]/NET0131 ,
		\datao[30]_pad ,
		_w1372_
	);
	LUT2 #(
		.INIT('he)
	) name23 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('hccc8)
	) name24 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[17]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1374_
	);
	LUT4 #(
		.INIT('h0010)
	) name25 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[17]/NET0131 ,
		\datao[30]_pad ,
		_w1375_
	);
	LUT2 #(
		.INIT('he)
	) name26 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('hccc8)
	) name27 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[18]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1377_
	);
	LUT4 #(
		.INIT('h0010)
	) name28 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[18]/NET0131 ,
		\datao[30]_pad ,
		_w1378_
	);
	LUT2 #(
		.INIT('he)
	) name29 (
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('hccc8)
	) name30 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[19]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1380_
	);
	LUT4 #(
		.INIT('h0010)
	) name31 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[19]/NET0131 ,
		\datao[30]_pad ,
		_w1381_
	);
	LUT2 #(
		.INIT('he)
	) name32 (
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('hccc8)
	) name33 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[1]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1383_
	);
	LUT4 #(
		.INIT('h0010)
	) name34 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[1]/NET0131 ,
		\datao[30]_pad ,
		_w1384_
	);
	LUT2 #(
		.INIT('he)
	) name35 (
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT4 #(
		.INIT('hccc8)
	) name36 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[20]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1386_
	);
	LUT4 #(
		.INIT('h0010)
	) name37 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[20]/NET0131 ,
		\datao[30]_pad ,
		_w1387_
	);
	LUT2 #(
		.INIT('he)
	) name38 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('hccc8)
	) name39 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[21]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1389_
	);
	LUT4 #(
		.INIT('h0010)
	) name40 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[21]/NET0131 ,
		\datao[30]_pad ,
		_w1390_
	);
	LUT2 #(
		.INIT('he)
	) name41 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT4 #(
		.INIT('hccc8)
	) name42 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[22]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1392_
	);
	LUT4 #(
		.INIT('h0010)
	) name43 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[22]/NET0131 ,
		\datao[30]_pad ,
		_w1393_
	);
	LUT2 #(
		.INIT('he)
	) name44 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('hccc8)
	) name45 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[23]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1395_
	);
	LUT4 #(
		.INIT('h0010)
	) name46 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[23]/NET0131 ,
		\datao[30]_pad ,
		_w1396_
	);
	LUT2 #(
		.INIT('he)
	) name47 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('hccc8)
	) name48 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[24]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1398_
	);
	LUT4 #(
		.INIT('h0010)
	) name49 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[24]/NET0131 ,
		\datao[30]_pad ,
		_w1399_
	);
	LUT2 #(
		.INIT('he)
	) name50 (
		_w1398_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('hccc8)
	) name51 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[25]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1401_
	);
	LUT4 #(
		.INIT('h0010)
	) name52 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[25]/NET0131 ,
		\datao[30]_pad ,
		_w1402_
	);
	LUT2 #(
		.INIT('he)
	) name53 (
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('hccc8)
	) name54 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[26]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1404_
	);
	LUT4 #(
		.INIT('h0010)
	) name55 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[26]/NET0131 ,
		\datao[30]_pad ,
		_w1405_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT4 #(
		.INIT('hccc8)
	) name57 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[27]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1407_
	);
	LUT4 #(
		.INIT('h0010)
	) name58 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[27]/NET0131 ,
		\datao[30]_pad ,
		_w1408_
	);
	LUT2 #(
		.INIT('he)
	) name59 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('hccc8)
	) name60 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[28]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1410_
	);
	LUT4 #(
		.INIT('h0010)
	) name61 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[28]/NET0131 ,
		\datao[30]_pad ,
		_w1411_
	);
	LUT2 #(
		.INIT('he)
	) name62 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('hccc8)
	) name63 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[29]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1413_
	);
	LUT4 #(
		.INIT('h0010)
	) name64 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[29]/NET0131 ,
		\datao[30]_pad ,
		_w1414_
	);
	LUT2 #(
		.INIT('he)
	) name65 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('hccc8)
	) name66 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[2]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1416_
	);
	LUT4 #(
		.INIT('h0010)
	) name67 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[2]/NET0131 ,
		\datao[30]_pad ,
		_w1417_
	);
	LUT2 #(
		.INIT('he)
	) name68 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('hccc8)
	) name69 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[3]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1419_
	);
	LUT4 #(
		.INIT('h0010)
	) name70 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[3]/NET0131 ,
		\datao[30]_pad ,
		_w1420_
	);
	LUT2 #(
		.INIT('he)
	) name71 (
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('hccc8)
	) name72 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[4]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1422_
	);
	LUT4 #(
		.INIT('h0010)
	) name73 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[4]/NET0131 ,
		\datao[30]_pad ,
		_w1423_
	);
	LUT2 #(
		.INIT('he)
	) name74 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('hccc8)
	) name75 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[5]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1425_
	);
	LUT4 #(
		.INIT('h0010)
	) name76 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[5]/NET0131 ,
		\datao[30]_pad ,
		_w1426_
	);
	LUT2 #(
		.INIT('he)
	) name77 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT4 #(
		.INIT('hccc8)
	) name78 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[6]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1428_
	);
	LUT4 #(
		.INIT('h0010)
	) name79 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[6]/NET0131 ,
		\datao[30]_pad ,
		_w1429_
	);
	LUT2 #(
		.INIT('he)
	) name80 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('hccc8)
	) name81 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[7]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1431_
	);
	LUT4 #(
		.INIT('h0010)
	) name82 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[7]/NET0131 ,
		\datao[30]_pad ,
		_w1432_
	);
	LUT2 #(
		.INIT('he)
	) name83 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT4 #(
		.INIT('hccc8)
	) name84 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[8]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1434_
	);
	LUT4 #(
		.INIT('h0010)
	) name85 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[8]/NET0131 ,
		\datao[30]_pad ,
		_w1435_
	);
	LUT2 #(
		.INIT('he)
	) name86 (
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('hccc8)
	) name87 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Address_reg[9]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\datao[30]_pad ,
		_w1437_
	);
	LUT4 #(
		.INIT('h0010)
	) name88 (
		\P1_Datao_reg[30]/NET0131 ,
		\P2_Datao_reg[30]/NET0131 ,
		\P3_Address_reg[9]/NET0131 ,
		\datao[30]_pad ,
		_w1438_
	);
	LUT2 #(
		.INIT('he)
	) name89 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1440_
	);
	LUT3 #(
		.INIT('h07)
	) name91 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1441_
	);
	LUT3 #(
		.INIT('h78)
	) name92 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1442_
	);
	LUT4 #(
		.INIT('h0400)
	) name93 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1443_
	);
	LUT4 #(
		.INIT('h0080)
	) name94 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1444_
	);
	LUT4 #(
		.INIT('h135f)
	) name95 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('h0001)
	) name96 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1446_
	);
	LUT4 #(
		.INIT('h1000)
	) name97 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1447_
	);
	LUT4 #(
		.INIT('h135f)
	) name98 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0020)
	) name99 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1449_
	);
	LUT4 #(
		.INIT('h0008)
	) name100 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1450_
	);
	LUT4 #(
		.INIT('h153f)
	) name101 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT4 #(
		.INIT('h0200)
	) name102 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1452_
	);
	LUT4 #(
		.INIT('h8000)
	) name103 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1453_
	);
	LUT4 #(
		.INIT('h153f)
	) name104 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h8000)
	) name105 (
		_w1451_,
		_w1454_,
		_w1445_,
		_w1448_,
		_w1455_
	);
	LUT4 #(
		.INIT('h0040)
	) name106 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1456_
	);
	LUT4 #(
		.INIT('h4000)
	) name107 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1457_
	);
	LUT4 #(
		.INIT('h153f)
	) name108 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT4 #(
		.INIT('h0800)
	) name109 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1459_
	);
	LUT4 #(
		.INIT('h2000)
	) name110 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1460_
	);
	LUT4 #(
		.INIT('h135f)
	) name111 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('h0002)
	) name112 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1462_
	);
	LUT4 #(
		.INIT('h0004)
	) name113 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1463_
	);
	LUT4 #(
		.INIT('h135f)
	) name114 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('h0100)
	) name115 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1465_
	);
	LUT4 #(
		.INIT('h0010)
	) name116 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1466_
	);
	LUT4 #(
		.INIT('h153f)
	) name117 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT4 #(
		.INIT('h8000)
	) name118 (
		_w1464_,
		_w1467_,
		_w1458_,
		_w1461_,
		_w1468_
	);
	LUT4 #(
		.INIT('h153f)
	) name119 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1452_,
		_w1444_,
		_w1469_
	);
	LUT4 #(
		.INIT('h153f)
	) name120 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1466_,
		_w1460_,
		_w1470_
	);
	LUT4 #(
		.INIT('h153f)
	) name121 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1450_,
		_w1443_,
		_w1471_
	);
	LUT4 #(
		.INIT('h135f)
	) name122 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1447_,
		_w1456_,
		_w1472_
	);
	LUT4 #(
		.INIT('h8000)
	) name123 (
		_w1471_,
		_w1472_,
		_w1469_,
		_w1470_,
		_w1473_
	);
	LUT4 #(
		.INIT('h135f)
	) name124 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1446_,
		_w1463_,
		_w1474_
	);
	LUT4 #(
		.INIT('h153f)
	) name125 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1453_,
		_w1457_,
		_w1475_
	);
	LUT4 #(
		.INIT('h153f)
	) name126 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w1462_,
		_w1459_,
		_w1476_
	);
	LUT4 #(
		.INIT('h135f)
	) name127 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1449_,
		_w1465_,
		_w1477_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		_w1476_,
		_w1477_,
		_w1474_,
		_w1475_,
		_w1478_
	);
	LUT4 #(
		.INIT('h0777)
	) name129 (
		_w1455_,
		_w1468_,
		_w1473_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h153f)
	) name130 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1450_,
		_w1457_,
		_w1480_
	);
	LUT4 #(
		.INIT('h153f)
	) name131 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1466_,
		_w1460_,
		_w1481_
	);
	LUT4 #(
		.INIT('h153f)
	) name132 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1456_,
		_w1459_,
		_w1482_
	);
	LUT4 #(
		.INIT('h135f)
	) name133 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1443_,
		_w1465_,
		_w1483_
	);
	LUT4 #(
		.INIT('h8000)
	) name134 (
		_w1482_,
		_w1483_,
		_w1480_,
		_w1481_,
		_w1484_
	);
	LUT4 #(
		.INIT('h135f)
	) name135 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1453_,
		_w1463_,
		_w1485_
	);
	LUT4 #(
		.INIT('h135f)
	) name136 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w1446_,
		_w1447_,
		_w1486_
	);
	LUT4 #(
		.INIT('h153f)
	) name137 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1452_,
		_w1444_,
		_w1487_
	);
	LUT4 #(
		.INIT('h153f)
	) name138 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1449_,
		_w1462_,
		_w1488_
	);
	LUT4 #(
		.INIT('h8000)
	) name139 (
		_w1487_,
		_w1488_,
		_w1485_,
		_w1486_,
		_w1489_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w1484_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h153f)
	) name141 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1444_,
		_w1459_,
		_w1491_
	);
	LUT4 #(
		.INIT('h153f)
	) name142 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w1443_,
		_w1446_,
		_w1492_
	);
	LUT4 #(
		.INIT('h153f)
	) name143 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1449_,
		_w1453_,
		_w1493_
	);
	LUT4 #(
		.INIT('h135f)
	) name144 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w1447_,
		_w1460_,
		_w1494_
	);
	LUT4 #(
		.INIT('h8000)
	) name145 (
		_w1493_,
		_w1494_,
		_w1491_,
		_w1492_,
		_w1495_
	);
	LUT4 #(
		.INIT('h135f)
	) name146 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1466_,
		_w1456_,
		_w1496_
	);
	LUT4 #(
		.INIT('h153f)
	) name147 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1465_,
		_w1457_,
		_w1497_
	);
	LUT4 #(
		.INIT('h135f)
	) name148 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1450_,
		_w1452_,
		_w1498_
	);
	LUT4 #(
		.INIT('h135f)
	) name149 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1462_,
		_w1463_,
		_w1499_
	);
	LUT4 #(
		.INIT('h8000)
	) name150 (
		_w1498_,
		_w1499_,
		_w1496_,
		_w1497_,
		_w1500_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w1495_,
		_w1500_,
		_w1501_
	);
	LUT4 #(
		.INIT('h0888)
	) name152 (
		_w1484_,
		_w1489_,
		_w1495_,
		_w1500_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w1479_,
		_w1502_,
		_w1503_
	);
	LUT4 #(
		.INIT('h135f)
	) name154 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1463_,
		_w1466_,
		_w1504_
	);
	LUT4 #(
		.INIT('h135f)
	) name155 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1453_,
		_w1462_,
		_w1505_
	);
	LUT4 #(
		.INIT('h135f)
	) name156 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w1446_,
		_w1459_,
		_w1506_
	);
	LUT4 #(
		.INIT('h135f)
	) name157 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1443_,
		_w1444_,
		_w1507_
	);
	LUT4 #(
		.INIT('h8000)
	) name158 (
		_w1506_,
		_w1507_,
		_w1504_,
		_w1505_,
		_w1508_
	);
	LUT4 #(
		.INIT('h153f)
	) name159 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1452_,
		_w1456_,
		_w1509_
	);
	LUT4 #(
		.INIT('h135f)
	) name160 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w1447_,
		_w1460_,
		_w1510_
	);
	LUT4 #(
		.INIT('h153f)
	) name161 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1465_,
		_w1457_,
		_w1511_
	);
	LUT4 #(
		.INIT('h153f)
	) name162 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1449_,
		_w1450_,
		_w1512_
	);
	LUT4 #(
		.INIT('h8000)
	) name163 (
		_w1511_,
		_w1512_,
		_w1509_,
		_w1510_,
		_w1513_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w1508_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('h135f)
	) name165 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1453_,
		_w1463_,
		_w1515_
	);
	LUT4 #(
		.INIT('h153f)
	) name166 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1452_,
		_w1443_,
		_w1516_
	);
	LUT4 #(
		.INIT('h135f)
	) name167 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w1446_,
		_w1459_,
		_w1517_
	);
	LUT4 #(
		.INIT('h153f)
	) name168 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1450_,
		_w1447_,
		_w1518_
	);
	LUT4 #(
		.INIT('h8000)
	) name169 (
		_w1517_,
		_w1518_,
		_w1515_,
		_w1516_,
		_w1519_
	);
	LUT4 #(
		.INIT('h135f)
	) name170 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1462_,
		_w1456_,
		_w1520_
	);
	LUT4 #(
		.INIT('h153f)
	) name171 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1466_,
		_w1460_,
		_w1521_
	);
	LUT4 #(
		.INIT('h153f)
	) name172 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1465_,
		_w1457_,
		_w1522_
	);
	LUT4 #(
		.INIT('h135f)
	) name173 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1449_,
		_w1444_,
		_w1523_
	);
	LUT4 #(
		.INIT('h8000)
	) name174 (
		_w1522_,
		_w1523_,
		_w1520_,
		_w1521_,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w1519_,
		_w1524_,
		_w1525_
	);
	LUT4 #(
		.INIT('h0888)
	) name176 (
		_w1508_,
		_w1513_,
		_w1519_,
		_w1524_,
		_w1526_
	);
	LUT4 #(
		.INIT('h135f)
	) name177 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1449_,
		_w1452_,
		_w1527_
	);
	LUT4 #(
		.INIT('h153f)
	) name178 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w1443_,
		_w1446_,
		_w1528_
	);
	LUT4 #(
		.INIT('h153f)
	) name179 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1463_,
		_w1460_,
		_w1529_
	);
	LUT4 #(
		.INIT('h153f)
	) name180 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1444_,
		_w1457_,
		_w1530_
	);
	LUT4 #(
		.INIT('h8000)
	) name181 (
		_w1529_,
		_w1530_,
		_w1527_,
		_w1528_,
		_w1531_
	);
	LUT4 #(
		.INIT('h135f)
	) name182 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1447_,
		_w1466_,
		_w1532_
	);
	LUT4 #(
		.INIT('h153f)
	) name183 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1465_,
		_w1456_,
		_w1533_
	);
	LUT4 #(
		.INIT('h153f)
	) name184 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1450_,
		_w1462_,
		_w1534_
	);
	LUT4 #(
		.INIT('h153f)
	) name185 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1453_,
		_w1459_,
		_w1535_
	);
	LUT4 #(
		.INIT('h8000)
	) name186 (
		_w1534_,
		_w1535_,
		_w1532_,
		_w1533_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w1531_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('h135f)
	) name188 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1462_,
		_w1466_,
		_w1538_
	);
	LUT4 #(
		.INIT('h135f)
	) name189 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1463_,
		_w1465_,
		_w1539_
	);
	LUT4 #(
		.INIT('h153f)
	) name190 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1449_,
		_w1447_,
		_w1540_
	);
	LUT4 #(
		.INIT('h153f)
	) name191 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1450_,
		_w1446_,
		_w1541_
	);
	LUT4 #(
		.INIT('h8000)
	) name192 (
		_w1540_,
		_w1541_,
		_w1538_,
		_w1539_,
		_w1542_
	);
	LUT4 #(
		.INIT('h153f)
	) name193 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w1457_,
		_w1459_,
		_w1543_
	);
	LUT4 #(
		.INIT('h153f)
	) name194 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1456_,
		_w1460_,
		_w1544_
	);
	LUT4 #(
		.INIT('h153f)
	) name195 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1452_,
		_w1444_,
		_w1545_
	);
	LUT4 #(
		.INIT('h153f)
	) name196 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1453_,
		_w1443_,
		_w1546_
	);
	LUT4 #(
		.INIT('h8000)
	) name197 (
		_w1545_,
		_w1546_,
		_w1543_,
		_w1544_,
		_w1547_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w1542_,
		_w1547_,
		_w1548_
	);
	LUT3 #(
		.INIT('h02)
	) name199 (
		_w1526_,
		_w1537_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w1503_,
		_w1549_,
		_w1550_
	);
	LUT4 #(
		.INIT('h0888)
	) name201 (
		_w1455_,
		_w1468_,
		_w1473_,
		_w1478_,
		_w1551_
	);
	LUT4 #(
		.INIT('h8000)
	) name202 (
		_w1484_,
		_w1489_,
		_w1495_,
		_w1500_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w1549_,
		_w1553_,
		_w1554_
	);
	LUT3 #(
		.INIT('h37)
	) name205 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w1555_
	);
	LUT4 #(
		.INIT('h0777)
	) name206 (
		_w1508_,
		_w1513_,
		_w1519_,
		_w1524_,
		_w1556_
	);
	LUT4 #(
		.INIT('h0888)
	) name207 (
		_w1531_,
		_w1536_,
		_w1542_,
		_w1547_,
		_w1557_
	);
	LUT4 #(
		.INIT('h8000)
	) name208 (
		_w1479_,
		_w1552_,
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h8000)
	) name209 (
		_w1479_,
		_w1502_,
		_w1556_,
		_w1557_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h8000)
	) name211 (
		_w1455_,
		_w1468_,
		_w1473_,
		_w1478_,
		_w1561_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w1552_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('h8000)
	) name213 (
		_w1548_,
		_w1552_,
		_w1556_,
		_w1561_,
		_w1563_
	);
	LUT4 #(
		.INIT('h8000)
	) name214 (
		_w1531_,
		_w1536_,
		_w1542_,
		_w1547_,
		_w1564_
	);
	LUT4 #(
		.INIT('h8000)
	) name215 (
		_w1479_,
		_w1502_,
		_w1526_,
		_w1564_,
		_w1565_
	);
	LUT4 #(
		.INIT('h8000)
	) name216 (
		_w1479_,
		_w1526_,
		_w1552_,
		_w1564_,
		_w1566_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w1490_,
		_w1561_,
		_w1567_
	);
	LUT4 #(
		.INIT('h4000)
	) name218 (
		_w1490_,
		_w1556_,
		_w1557_,
		_w1561_,
		_w1568_
	);
	LUT3 #(
		.INIT('h01)
	) name219 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('h0001)
	) name220 (
		_w1563_,
		_w1565_,
		_w1566_,
		_w1568_,
		_w1570_
	);
	LUT3 #(
		.INIT('h80)
	) name221 (
		_w1555_,
		_w1560_,
		_w1570_,
		_w1571_
	);
	LUT4 #(
		.INIT('h7000)
	) name222 (
		_w1508_,
		_w1513_,
		_w1519_,
		_w1524_,
		_w1572_
	);
	LUT3 #(
		.INIT('h40)
	) name223 (
		_w1501_,
		_w1557_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('h8000)
	) name224 (
		_w1495_,
		_w1500_,
		_w1508_,
		_w1513_,
		_w1574_
	);
	LUT4 #(
		.INIT('h0888)
	) name225 (
		_w1473_,
		_w1478_,
		_w1484_,
		_w1489_,
		_w1575_
	);
	LUT4 #(
		.INIT('h8000)
	) name226 (
		_w1525_,
		_w1564_,
		_w1575_,
		_w1574_,
		_w1576_
	);
	LUT4 #(
		.INIT('h7000)
	) name227 (
		_w1455_,
		_w1468_,
		_w1473_,
		_w1478_,
		_w1577_
	);
	LUT4 #(
		.INIT('h8000)
	) name228 (
		_w1502_,
		_w1564_,
		_w1572_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('h0007)
	) name229 (
		_w1567_,
		_w1573_,
		_w1576_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name230 (
		_w1514_,
		_w1525_,
		_w1537_,
		_w1564_,
		_w1580_
	);
	LUT4 #(
		.INIT('h8000)
	) name231 (
		_w1502_,
		_w1551_,
		_w1556_,
		_w1557_,
		_w1581_
	);
	LUT3 #(
		.INIT('h0d)
	) name232 (
		_w1562_,
		_w1580_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w1579_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1584_
	);
	LUT4 #(
		.INIT('h08ce)
	) name235 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1585_
	);
	LUT3 #(
		.INIT('hb2)
	) name236 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1585_,
		_w1586_
	);
	LUT4 #(
		.INIT('h40d0)
	) name237 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1584_,
		_w1585_,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1588_
	);
	LUT4 #(
		.INIT('h004d)
	) name239 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1585_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h9)
	) name240 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1590_
	);
	LUT2 #(
		.INIT('h9)
	) name241 (
		_w1585_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name242 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1586_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h9)
	) name243 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1593_
	);
	LUT4 #(
		.INIT('h8421)
	) name244 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1594_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w1587_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w1592_,
		_w1595_,
		_w1596_
	);
	LUT4 #(
		.INIT('haaa9)
	) name247 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1440_,
		_w1592_,
		_w1595_,
		_w1597_
	);
	LUT4 #(
		.INIT('hc800)
	) name248 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('h0075)
	) name249 (
		_w1442_,
		_w1571_,
		_w1583_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('hc639)
	) name250 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1600_
	);
	LUT3 #(
		.INIT('h0e)
	) name251 (
		_w1584_,
		_w1589_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		_w1592_,
		_w1601_,
		_w1602_
	);
	LUT4 #(
		.INIT('hdc00)
	) name253 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1602_,
		_w1603_
	);
	LUT3 #(
		.INIT('h13)
	) name254 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w1605_
	);
	LUT3 #(
		.INIT('h31)
	) name256 (
		_w1592_,
		_w1605_,
		_w1601_,
		_w1606_
	);
	LUT4 #(
		.INIT('h00ec)
	) name257 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w1608_
	);
	LUT3 #(
		.INIT('h04)
	) name259 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1609_
	);
	LUT3 #(
		.INIT('h10)
	) name260 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1610_
	);
	LUT3 #(
		.INIT('heb)
	) name261 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w1611_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w1605_,
		_w1611_,
		_w1612_
	);
	LUT4 #(
		.INIT('h00dc)
	) name263 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h01)
	) name264 (
		_w1607_,
		_w1613_,
		_w1603_,
		_w1614_
	);
	LUT4 #(
		.INIT('h0002)
	) name265 (
		_w1560_,
		_w1607_,
		_w1613_,
		_w1603_,
		_w1615_
	);
	LUT4 #(
		.INIT('h00dc)
	) name266 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1611_,
		_w1616_
	);
	LUT4 #(
		.INIT('h0545)
	) name267 (
		_w1563_,
		_w1604_,
		_w1606_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1618_
	);
	LUT4 #(
		.INIT('hf391)
	) name269 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1615_,
		_w1617_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w1599_,
		_w1619_,
		_w1620_
	);
	LUT3 #(
		.INIT('h80)
	) name271 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1599_,
		_w1619_,
		_w1621_
	);
	LUT4 #(
		.INIT('h007f)
	) name272 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1622_
	);
	LUT4 #(
		.INIT('h7f80)
	) name273 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1623_
	);
	LUT3 #(
		.INIT('hb0)
	) name274 (
		_w1571_,
		_w1583_,
		_w1623_,
		_w1624_
	);
	LUT4 #(
		.INIT('hdc00)
	) name275 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1611_,
		_w1625_
	);
	LUT4 #(
		.INIT('hfe00)
	) name276 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1602_,
		_w1626_
	);
	LUT3 #(
		.INIT('h78)
	) name277 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1627_
	);
	LUT3 #(
		.INIT('h65)
	) name278 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1605_,
		_w1618_,
		_w1628_
	);
	LUT4 #(
		.INIT('h00dc)
	) name279 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('h0002)
	) name280 (
		_w1560_,
		_w1625_,
		_w1626_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h0031)
	) name281 (
		_w1604_,
		_w1602_,
		_w1616_,
		_w1628_,
		_w1631_
	);
	LUT4 #(
		.INIT('h0002)
	) name282 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1441_,
		_w1592_,
		_w1595_,
		_w1632_
	);
	LUT4 #(
		.INIT('h5554)
	) name283 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1441_,
		_w1592_,
		_w1595_,
		_w1633_
	);
	LUT4 #(
		.INIT('h00c8)
	) name284 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w1563_,
		_w1627_,
		_w1635_
	);
	LUT3 #(
		.INIT('h0b)
	) name286 (
		_w1632_,
		_w1634_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h3100)
	) name287 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1631_,
		_w1630_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		_w1624_,
		_w1637_,
		_w1638_
	);
	LUT3 #(
		.INIT('h20)
	) name289 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1624_,
		_w1637_,
		_w1639_
	);
	LUT4 #(
		.INIT('hc800)
	) name290 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w1596_,
		_w1640_
	);
	LUT4 #(
		.INIT('h0010)
	) name291 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1571_,
		_w1583_,
		_w1640_,
		_w1641_
	);
	LUT3 #(
		.INIT('h08)
	) name292 (
		_w1549_,
		_w1553_,
		_w1596_,
		_w1642_
	);
	LUT4 #(
		.INIT('hff37)
	) name293 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w1596_,
		_w1643_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1560_,
		_w1570_,
		_w1643_,
		_w1644_
	);
	LUT3 #(
		.INIT('ha8)
	) name295 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1641_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h9)
	) name296 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1646_
	);
	LUT4 #(
		.INIT('h00fb)
	) name297 (
		_w1571_,
		_w1583_,
		_w1640_,
		_w1646_,
		_w1647_
	);
	LUT3 #(
		.INIT('h51)
	) name298 (
		_w1569_,
		_w1606_,
		_w1625_,
		_w1648_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w1560_,
		_w1643_,
		_w1649_
	);
	LUT4 #(
		.INIT('h4e44)
	) name300 (
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1617_,
		_w1648_,
		_w1649_,
		_w1650_
	);
	LUT3 #(
		.INIT('h20)
	) name301 (
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1647_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('h0001)
	) name302 (
		_w1621_,
		_w1639_,
		_w1645_,
		_w1651_,
		_w1652_
	);
	LUT3 #(
		.INIT('h45)
	) name303 (
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1647_,
		_w1650_,
		_w1653_
	);
	LUT4 #(
		.INIT('h0701)
	) name304 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1620_,
		_w1639_,
		_w1653_,
		_w1654_
	);
	LUT3 #(
		.INIT('h80)
	) name305 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1599_,
		_w1619_,
		_w1655_
	);
	LUT4 #(
		.INIT('h00ec)
	) name306 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1602_,
		_w1656_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w1602_,
		_w1613_,
		_w1657_
	);
	LUT4 #(
		.INIT('hf0fb)
	) name308 (
		_w1604_,
		_w1605_,
		_w1602_,
		_w1613_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w1558_,
		_w1596_,
		_w1659_
	);
	LUT4 #(
		.INIT('h000e)
	) name310 (
		_w1584_,
		_w1589_,
		_w1593_,
		_w1600_,
		_w1660_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		_w1592_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h5f13)
	) name312 (
		_w1558_,
		_w1559_,
		_w1596_,
		_w1661_,
		_w1662_
	);
	LUT3 #(
		.INIT('hd0)
	) name313 (
		\P2_Flush_reg/NET0131 ,
		_w1658_,
		_w1662_,
		_w1663_
	);
	LUT3 #(
		.INIT('h51)
	) name314 (
		\P2_More_reg/NET0131 ,
		_w1592_,
		_w1601_,
		_w1664_
	);
	LUT4 #(
		.INIT('h00fe)
	) name315 (
		_w1607_,
		_w1613_,
		_w1603_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w1559_,
		_w1661_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name317 (
		_w1558_,
		_w1596_,
		_w1667_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w1643_,
		_w1667_,
		_w1668_
	);
	LUT3 #(
		.INIT('h02)
	) name319 (
		_w1643_,
		_w1666_,
		_w1667_,
		_w1669_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w1665_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w1663_,
		_w1670_,
		_w1671_
	);
	LUT3 #(
		.INIT('he0)
	) name322 (
		_w1638_,
		_w1655_,
		_w1671_,
		_w1672_
	);
	LUT3 #(
		.INIT('h15)
	) name323 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w1673_
	);
	LUT3 #(
		.INIT('h0d)
	) name324 (
		_w1592_,
		_w1601_,
		_w1611_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w1566_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('h80)
	) name326 (
		_w1566_,
		_w1673_,
		_w1674_,
		_w1676_
	);
	LUT4 #(
		.INIT('h0010)
	) name327 (
		_w1654_,
		_w1652_,
		_w1672_,
		_w1676_,
		_w1677_
	);
	LUT4 #(
		.INIT('h0020)
	) name328 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1678_
	);
	LUT4 #(
		.INIT('h0004)
	) name329 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1679_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('h02)
	) name331 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1681_
	);
	LUT4 #(
		.INIT('h0002)
	) name332 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1683_
	);
	LUT3 #(
		.INIT('hf9)
	) name334 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w1684_
	);
	LUT4 #(
		.INIT('h1098)
	) name335 (
		\P2_State2_reg[1]/NET0131 ,
		_w1605_,
		_w1681_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w1680_,
		_w1685_,
		_w1686_
	);
	LUT3 #(
		.INIT('h4f)
	) name337 (
		_w1677_,
		_w1678_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('h0001)
	) name338 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1688_
	);
	LUT4 #(
		.INIT('h0010)
	) name339 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1689_
	);
	LUT4 #(
		.INIT('h135f)
	) name340 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1688_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h0020)
	) name341 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1691_
	);
	LUT4 #(
		.INIT('h0002)
	) name342 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1692_
	);
	LUT4 #(
		.INIT('h153f)
	) name343 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h0400)
	) name344 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1695_
	);
	LUT4 #(
		.INIT('h0800)
	) name346 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1696_
	);
	LUT4 #(
		.INIT('h135f)
	) name347 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w1694_,
		_w1696_,
		_w1697_
	);
	LUT4 #(
		.INIT('h1000)
	) name348 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1698_
	);
	LUT4 #(
		.INIT('h4000)
	) name349 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1699_
	);
	LUT4 #(
		.INIT('h135f)
	) name350 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h8000)
	) name351 (
		_w1697_,
		_w1700_,
		_w1690_,
		_w1693_,
		_w1701_
	);
	LUT4 #(
		.INIT('h0008)
	) name352 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1702_
	);
	LUT4 #(
		.INIT('h0200)
	) name353 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1703_
	);
	LUT4 #(
		.INIT('h135f)
	) name354 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h2000)
	) name355 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1705_
	);
	LUT4 #(
		.INIT('h8000)
	) name356 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1706_
	);
	LUT4 #(
		.INIT('h135f)
	) name357 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT4 #(
		.INIT('h0080)
	) name358 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1708_
	);
	LUT4 #(
		.INIT('h0004)
	) name359 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1709_
	);
	LUT4 #(
		.INIT('h153f)
	) name360 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h0040)
	) name361 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1711_
	);
	LUT4 #(
		.INIT('h0100)
	) name362 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1712_
	);
	LUT4 #(
		.INIT('h135f)
	) name363 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h8000)
	) name364 (
		_w1710_,
		_w1713_,
		_w1704_,
		_w1707_,
		_w1714_
	);
	LUT4 #(
		.INIT('h135f)
	) name365 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1696_,
		_w1703_,
		_w1715_
	);
	LUT4 #(
		.INIT('h153f)
	) name366 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1702_,
		_w1706_,
		_w1716_
	);
	LUT4 #(
		.INIT('h153f)
	) name367 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w1699_,
		_w1688_,
		_w1717_
	);
	LUT4 #(
		.INIT('h135f)
	) name368 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1698_,
		_w1711_,
		_w1718_
	);
	LUT4 #(
		.INIT('h8000)
	) name369 (
		_w1717_,
		_w1718_,
		_w1715_,
		_w1716_,
		_w1719_
	);
	LUT4 #(
		.INIT('h135f)
	) name370 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1692_,
		_w1709_,
		_w1720_
	);
	LUT4 #(
		.INIT('h135f)
	) name371 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1708_,
		_w1712_,
		_w1721_
	);
	LUT4 #(
		.INIT('h135f)
	) name372 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1694_,
		_w1691_,
		_w1722_
	);
	LUT4 #(
		.INIT('h153f)
	) name373 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1689_,
		_w1705_,
		_w1723_
	);
	LUT4 #(
		.INIT('h8000)
	) name374 (
		_w1722_,
		_w1723_,
		_w1720_,
		_w1721_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w1719_,
		_w1724_,
		_w1725_
	);
	LUT4 #(
		.INIT('h0888)
	) name376 (
		_w1701_,
		_w1714_,
		_w1719_,
		_w1724_,
		_w1726_
	);
	LUT4 #(
		.INIT('h135f)
	) name377 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1689_,
		_w1691_,
		_w1727_
	);
	LUT4 #(
		.INIT('h135f)
	) name378 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w1705_,
		_w1706_,
		_w1728_
	);
	LUT4 #(
		.INIT('h135f)
	) name379 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1699_,
		_w1708_,
		_w1729_
	);
	LUT4 #(
		.INIT('h135f)
	) name380 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1712_,
		_w1703_,
		_w1730_
	);
	LUT4 #(
		.INIT('h8000)
	) name381 (
		_w1729_,
		_w1730_,
		_w1727_,
		_w1728_,
		_w1731_
	);
	LUT4 #(
		.INIT('h153f)
	) name382 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w1696_,
		_w1688_,
		_w1732_
	);
	LUT4 #(
		.INIT('h135f)
	) name383 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w1698_,
		_w1709_,
		_w1733_
	);
	LUT4 #(
		.INIT('h135f)
	) name384 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1694_,
		_w1702_,
		_w1734_
	);
	LUT4 #(
		.INIT('h135f)
	) name385 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1692_,
		_w1711_,
		_w1735_
	);
	LUT4 #(
		.INIT('h8000)
	) name386 (
		_w1734_,
		_w1735_,
		_w1732_,
		_w1733_,
		_w1736_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w1731_,
		_w1736_,
		_w1737_
	);
	LUT4 #(
		.INIT('h135f)
	) name388 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1708_,
		_w1703_,
		_w1738_
	);
	LUT4 #(
		.INIT('h135f)
	) name389 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1699_,
		_w1689_,
		_w1739_
	);
	LUT4 #(
		.INIT('h135f)
	) name390 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1694_,
		_w1691_,
		_w1740_
	);
	LUT4 #(
		.INIT('h135f)
	) name391 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1696_,
		_w1709_,
		_w1741_
	);
	LUT4 #(
		.INIT('h8000)
	) name392 (
		_w1740_,
		_w1741_,
		_w1738_,
		_w1739_,
		_w1742_
	);
	LUT4 #(
		.INIT('h135f)
	) name393 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1698_,
		_w1692_,
		_w1743_
	);
	LUT4 #(
		.INIT('h135f)
	) name394 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1688_,
		_w1705_,
		_w1744_
	);
	LUT4 #(
		.INIT('h135f)
	) name395 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1711_,
		_w1712_,
		_w1745_
	);
	LUT4 #(
		.INIT('h153f)
	) name396 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1702_,
		_w1706_,
		_w1746_
	);
	LUT4 #(
		.INIT('h8000)
	) name397 (
		_w1745_,
		_w1746_,
		_w1743_,
		_w1744_,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w1742_,
		_w1747_,
		_w1748_
	);
	LUT4 #(
		.INIT('h0777)
	) name399 (
		_w1731_,
		_w1736_,
		_w1742_,
		_w1747_,
		_w1749_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w1726_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h135f)
	) name401 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1688_,
		_w1689_,
		_w1751_
	);
	LUT4 #(
		.INIT('h153f)
	) name402 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1691_,
		_w1692_,
		_w1752_
	);
	LUT4 #(
		.INIT('h135f)
	) name403 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w1694_,
		_w1696_,
		_w1753_
	);
	LUT4 #(
		.INIT('h135f)
	) name404 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1698_,
		_w1699_,
		_w1754_
	);
	LUT4 #(
		.INIT('h8000)
	) name405 (
		_w1753_,
		_w1754_,
		_w1751_,
		_w1752_,
		_w1755_
	);
	LUT4 #(
		.INIT('h135f)
	) name406 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1702_,
		_w1703_,
		_w1756_
	);
	LUT4 #(
		.INIT('h135f)
	) name407 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1705_,
		_w1706_,
		_w1757_
	);
	LUT4 #(
		.INIT('h153f)
	) name408 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1708_,
		_w1709_,
		_w1758_
	);
	LUT4 #(
		.INIT('h135f)
	) name409 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1711_,
		_w1712_,
		_w1759_
	);
	LUT4 #(
		.INIT('h8000)
	) name410 (
		_w1758_,
		_w1759_,
		_w1756_,
		_w1757_,
		_w1760_
	);
	LUT4 #(
		.INIT('h135f)
	) name411 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1688_,
		_w1689_,
		_w1761_
	);
	LUT4 #(
		.INIT('h153f)
	) name412 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1691_,
		_w1692_,
		_w1762_
	);
	LUT4 #(
		.INIT('h135f)
	) name413 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w1694_,
		_w1696_,
		_w1763_
	);
	LUT4 #(
		.INIT('h135f)
	) name414 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1698_,
		_w1699_,
		_w1764_
	);
	LUT4 #(
		.INIT('h8000)
	) name415 (
		_w1763_,
		_w1764_,
		_w1761_,
		_w1762_,
		_w1765_
	);
	LUT4 #(
		.INIT('h135f)
	) name416 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1702_,
		_w1703_,
		_w1766_
	);
	LUT4 #(
		.INIT('h135f)
	) name417 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w1705_,
		_w1706_,
		_w1767_
	);
	LUT4 #(
		.INIT('h153f)
	) name418 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1708_,
		_w1709_,
		_w1768_
	);
	LUT4 #(
		.INIT('h135f)
	) name419 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1711_,
		_w1712_,
		_w1769_
	);
	LUT4 #(
		.INIT('h8000)
	) name420 (
		_w1768_,
		_w1769_,
		_w1766_,
		_w1767_,
		_w1770_
	);
	LUT4 #(
		.INIT('h0888)
	) name421 (
		_w1755_,
		_w1760_,
		_w1765_,
		_w1770_,
		_w1771_
	);
	LUT4 #(
		.INIT('h135f)
	) name422 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1688_,
		_w1708_,
		_w1772_
	);
	LUT4 #(
		.INIT('h135f)
	) name423 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1699_,
		_w1692_,
		_w1773_
	);
	LUT4 #(
		.INIT('h135f)
	) name424 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1694_,
		_w1691_,
		_w1774_
	);
	LUT4 #(
		.INIT('h135f)
	) name425 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1696_,
		_w1698_,
		_w1775_
	);
	LUT4 #(
		.INIT('h8000)
	) name426 (
		_w1774_,
		_w1775_,
		_w1772_,
		_w1773_,
		_w1776_
	);
	LUT4 #(
		.INIT('h153f)
	) name427 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1689_,
		_w1702_,
		_w1777_
	);
	LUT4 #(
		.INIT('h153f)
	) name428 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1703_,
		_w1705_,
		_w1778_
	);
	LUT4 #(
		.INIT('h153f)
	) name429 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1711_,
		_w1706_,
		_w1779_
	);
	LUT4 #(
		.INIT('h135f)
	) name430 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1709_,
		_w1712_,
		_w1780_
	);
	LUT4 #(
		.INIT('h8000)
	) name431 (
		_w1779_,
		_w1780_,
		_w1777_,
		_w1778_,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w1776_,
		_w1781_,
		_w1782_
	);
	LUT4 #(
		.INIT('h135f)
	) name433 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1688_,
		_w1708_,
		_w1783_
	);
	LUT4 #(
		.INIT('h135f)
	) name434 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1699_,
		_w1692_,
		_w1784_
	);
	LUT4 #(
		.INIT('h135f)
	) name435 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1694_,
		_w1691_,
		_w1785_
	);
	LUT4 #(
		.INIT('h135f)
	) name436 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1696_,
		_w1698_,
		_w1786_
	);
	LUT4 #(
		.INIT('h8000)
	) name437 (
		_w1785_,
		_w1786_,
		_w1783_,
		_w1784_,
		_w1787_
	);
	LUT4 #(
		.INIT('h135f)
	) name438 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1702_,
		_w1703_,
		_w1788_
	);
	LUT4 #(
		.INIT('h153f)
	) name439 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1689_,
		_w1705_,
		_w1789_
	);
	LUT4 #(
		.INIT('h153f)
	) name440 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1711_,
		_w1706_,
		_w1790_
	);
	LUT4 #(
		.INIT('h135f)
	) name441 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1709_,
		_w1712_,
		_w1791_
	);
	LUT4 #(
		.INIT('h8000)
	) name442 (
		_w1790_,
		_w1791_,
		_w1788_,
		_w1789_,
		_w1792_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w1787_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h8000)
	) name444 (
		_w1776_,
		_w1781_,
		_w1787_,
		_w1792_,
		_w1794_
	);
	LUT4 #(
		.INIT('h8000)
	) name445 (
		_w1726_,
		_w1749_,
		_w1771_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h8000)
	) name446 (
		_w1701_,
		_w1714_,
		_w1719_,
		_w1724_,
		_w1796_
	);
	LUT4 #(
		.INIT('h8000)
	) name447 (
		_w1749_,
		_w1771_,
		_w1794_,
		_w1796_,
		_w1797_
	);
	LUT4 #(
		.INIT('h0777)
	) name448 (
		_w1755_,
		_w1760_,
		_w1765_,
		_w1770_,
		_w1798_
	);
	LUT4 #(
		.INIT('h0888)
	) name449 (
		_w1776_,
		_w1781_,
		_w1787_,
		_w1792_,
		_w1799_
	);
	LUT4 #(
		.INIT('h7000)
	) name450 (
		_w1701_,
		_w1714_,
		_w1731_,
		_w1736_,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w1748_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h8000)
	) name452 (
		_w1748_,
		_w1798_,
		_w1799_,
		_w1800_,
		_w1802_
	);
	LUT3 #(
		.INIT('h01)
	) name453 (
		_w1795_,
		_w1797_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		_w1748_,
		_w1796_,
		_w1804_
	);
	LUT3 #(
		.INIT('h80)
	) name455 (
		_w1737_,
		_w1748_,
		_w1796_,
		_w1805_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w1793_,
		_w1798_,
		_w1806_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w1805_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		_w1803_,
		_w1807_,
		_w1808_
	);
	LUT4 #(
		.INIT('h8000)
	) name459 (
		_w1749_,
		_w1796_,
		_w1798_,
		_w1799_,
		_w1809_
	);
	LUT4 #(
		.INIT('h8000)
	) name460 (
		_w1726_,
		_w1749_,
		_w1798_,
		_w1799_,
		_w1810_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w1809_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w1771_,
		_w1782_,
		_w1812_
	);
	LUT3 #(
		.INIT('h02)
	) name463 (
		_w1771_,
		_w1782_,
		_w1793_,
		_w1813_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w1750_,
		_w1813_,
		_w1814_
	);
	LUT3 #(
		.INIT('h1f)
	) name465 (
		_w1750_,
		_w1804_,
		_w1813_,
		_w1815_
	);
	LUT4 #(
		.INIT('h2000)
	) name466 (
		_w1803_,
		_w1807_,
		_w1811_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h7000)
	) name467 (
		_w1731_,
		_w1736_,
		_w1742_,
		_w1747_,
		_w1817_
	);
	LUT4 #(
		.INIT('h8000)
	) name468 (
		_w1726_,
		_w1798_,
		_w1799_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h7000)
	) name469 (
		_w1701_,
		_w1714_,
		_w1719_,
		_w1724_,
		_w1819_
	);
	LUT4 #(
		.INIT('h8000)
	) name470 (
		_w1755_,
		_w1760_,
		_w1765_,
		_w1770_,
		_w1820_
	);
	LUT4 #(
		.INIT('h8000)
	) name471 (
		_w1737_,
		_w1794_,
		_w1819_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h0007)
	) name472 (
		_w1805_,
		_w1812_,
		_w1818_,
		_w1821_,
		_w1822_
	);
	LUT4 #(
		.INIT('h7000)
	) name473 (
		_w1755_,
		_w1760_,
		_w1765_,
		_w1770_,
		_w1823_
	);
	LUT3 #(
		.INIT('h40)
	) name474 (
		_w1725_,
		_w1799_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w1801_,
		_w1824_,
		_w1825_
	);
	LUT3 #(
		.INIT('h80)
	) name476 (
		_w1737_,
		_w1794_,
		_w1823_,
		_w1826_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w1804_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w1726_,
		_w1748_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w1826_,
		_w1828_,
		_w1829_
	);
	LUT3 #(
		.INIT('h37)
	) name480 (
		_w1804_,
		_w1826_,
		_w1828_,
		_w1830_
	);
	LUT3 #(
		.INIT('h40)
	) name481 (
		_w1825_,
		_w1822_,
		_w1830_,
		_w1831_
	);
	LUT3 #(
		.INIT('h40)
	) name482 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w1832_
	);
	LUT4 #(
		.INIT('h23ff)
	) name483 (
		_w1737_,
		_w1750_,
		_w1804_,
		_w1813_,
		_w1833_
	);
	LUT2 #(
		.INIT('h4)
	) name484 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1834_
	);
	LUT4 #(
		.INIT('h08ce)
	) name485 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1835_
	);
	LUT3 #(
		.INIT('hb2)
	) name486 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('h40d0)
	) name487 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1834_,
		_w1835_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1838_
	);
	LUT4 #(
		.INIT('h004d)
	) name489 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1835_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h9)
	) name490 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1840_
	);
	LUT2 #(
		.INIT('h9)
	) name491 (
		_w1835_,
		_w1840_,
		_w1841_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name492 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1836_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h9)
	) name493 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1843_
	);
	LUT4 #(
		.INIT('h8421)
	) name494 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1844_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w1837_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1842_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h4)
	) name497 (
		_w1833_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h9)
	) name498 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1848_
	);
	LUT4 #(
		.INIT('h00fb)
	) name499 (
		_w1816_,
		_w1831_,
		_w1847_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('hc639)
	) name500 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1850_
	);
	LUT3 #(
		.INIT('h0e)
	) name501 (
		_w1834_,
		_w1839_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w1842_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w1725_,
		_w1802_,
		_w1853_
	);
	LUT3 #(
		.INIT('h13)
	) name504 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w1854_
	);
	LUT4 #(
		.INIT('h00ec)
	) name505 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w1852_,
		_w1855_
	);
	LUT3 #(
		.INIT('h04)
	) name506 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1856_
	);
	LUT3 #(
		.INIT('h10)
	) name507 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1857_
	);
	LUT3 #(
		.INIT('heb)
	) name508 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w1858_
	);
	LUT3 #(
		.INIT('h0d)
	) name509 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w1859_
	);
	LUT4 #(
		.INIT('hdc00)
	) name510 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1861_
	);
	LUT4 #(
		.INIT('h5501)
	) name512 (
		_w1807_,
		_w1855_,
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT3 #(
		.INIT('h08)
	) name513 (
		_w1750_,
		_w1813_,
		_w1846_,
		_w1863_
	);
	LUT4 #(
		.INIT('h0040)
	) name514 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w1846_,
		_w1864_
	);
	LUT3 #(
		.INIT('h02)
	) name515 (
		_w1811_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT4 #(
		.INIT('hdc00)
	) name516 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w1858_,
		_w1866_
	);
	LUT3 #(
		.INIT('h0d)
	) name517 (
		_w1842_,
		_w1851_,
		_w1861_,
		_w1867_
	);
	LUT3 #(
		.INIT('h45)
	) name518 (
		_w1803_,
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h8daf)
	) name519 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1868_,
		_w1862_,
		_w1865_,
		_w1869_
	);
	LUT3 #(
		.INIT('h54)
	) name520 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1849_,
		_w1869_,
		_w1870_
	);
	LUT4 #(
		.INIT('h0010)
	) name521 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1816_,
		_w1831_,
		_w1847_,
		_w1871_
	);
	LUT3 #(
		.INIT('h08)
	) name522 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1803_,
		_w1807_,
		_w1872_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w1865_,
		_w1872_,
		_w1873_
	);
	LUT3 #(
		.INIT('ha8)
	) name524 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w1871_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		_w1870_,
		_w1874_,
		_w1875_
	);
	LUT3 #(
		.INIT('h02)
	) name526 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1849_,
		_w1869_,
		_w1876_
	);
	LUT4 #(
		.INIT('hfe00)
	) name527 (
		_w1795_,
		_w1797_,
		_w1802_,
		_w1852_,
		_w1877_
	);
	LUT3 #(
		.INIT('h02)
	) name528 (
		_w1811_,
		_w1877_,
		_w1866_,
		_w1878_
	);
	LUT3 #(
		.INIT('h07)
	) name529 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1879_
	);
	LUT3 #(
		.INIT('h01)
	) name530 (
		_w1879_,
		_w1842_,
		_w1845_,
		_w1880_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w1833_,
		_w1880_,
		_w1881_
	);
	LUT3 #(
		.INIT('ha2)
	) name532 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1878_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h807f)
	) name533 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1883_
	);
	LUT3 #(
		.INIT('h0b)
	) name534 (
		_w1816_,
		_w1831_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1885_
	);
	LUT3 #(
		.INIT('h78)
	) name536 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1886_
	);
	LUT3 #(
		.INIT('h9a)
	) name537 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1861_,
		_w1885_,
		_w1887_
	);
	LUT3 #(
		.INIT('he0)
	) name538 (
		_w1855_,
		_w1860_,
		_w1887_,
		_w1888_
	);
	LUT3 #(
		.INIT('h80)
	) name539 (
		_w1805_,
		_w1806_,
		_w1886_,
		_w1889_
	);
	LUT4 #(
		.INIT('h0001)
	) name540 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1879_,
		_w1842_,
		_w1845_,
		_w1890_
	);
	LUT3 #(
		.INIT('h23)
	) name541 (
		_w1833_,
		_w1889_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w1888_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h10)
	) name543 (
		_w1884_,
		_w1882_,
		_w1892_,
		_w1893_
	);
	LUT4 #(
		.INIT('h0200)
	) name544 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1884_,
		_w1882_,
		_w1892_,
		_w1894_
	);
	LUT3 #(
		.INIT('h78)
	) name545 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1895_
	);
	LUT2 #(
		.INIT('h6)
	) name546 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1896_
	);
	LUT3 #(
		.INIT('h80)
	) name547 (
		_w1805_,
		_w1806_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('haaa9)
	) name548 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1695_,
		_w1842_,
		_w1845_,
		_w1898_
	);
	LUT3 #(
		.INIT('h45)
	) name549 (
		_w1897_,
		_w1833_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('h4f00)
	) name550 (
		_w1816_,
		_w1831_,
		_w1895_,
		_w1899_,
		_w1900_
	);
	LUT3 #(
		.INIT('ha8)
	) name551 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1797_,
		_w1802_,
		_w1901_
	);
	LUT4 #(
		.INIT('hc666)
	) name552 (
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1902_
	);
	LUT4 #(
		.INIT('hfe00)
	) name553 (
		_w1855_,
		_w1860_,
		_w1901_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('haaa2)
	) name554 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1811_,
		_w1877_,
		_w1866_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('h80)
	) name556 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1900_,
		_w1905_,
		_w1906_
	);
	LUT3 #(
		.INIT('h01)
	) name557 (
		_w1894_,
		_w1876_,
		_w1906_,
		_w1907_
	);
	LUT3 #(
		.INIT('h15)
	) name558 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1900_,
		_w1905_,
		_w1908_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w1894_,
		_w1908_,
		_w1909_
	);
	LUT3 #(
		.INIT('h80)
	) name560 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w1900_,
		_w1905_,
		_w1910_
	);
	LUT3 #(
		.INIT('h51)
	) name561 (
		\P1_More_reg/NET0131 ,
		_w1842_,
		_w1851_,
		_w1911_
	);
	LUT4 #(
		.INIT('h0045)
	) name562 (
		_w1803_,
		_w1866_,
		_w1867_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w1809_,
		_w1846_,
		_w1913_
	);
	LUT3 #(
		.INIT('h01)
	) name564 (
		_w1913_,
		_w1863_,
		_w1864_,
		_w1914_
	);
	LUT4 #(
		.INIT('h000e)
	) name565 (
		_w1834_,
		_w1839_,
		_w1850_,
		_w1843_,
		_w1915_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		_w1842_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w1810_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h0001)
	) name568 (
		_w1913_,
		_w1863_,
		_w1864_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		_w1912_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w1858_,
		_w1861_,
		_w1920_
	);
	LUT4 #(
		.INIT('h00dc)
	) name571 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w1920_,
		_w1921_
	);
	LUT4 #(
		.INIT('haaef)
	) name572 (
		_w1852_,
		_w1854_,
		_w1861_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		_w1810_,
		_w1916_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		_w1809_,
		_w1846_,
		_w1924_
	);
	LUT4 #(
		.INIT('h5f13)
	) name575 (
		_w1809_,
		_w1810_,
		_w1846_,
		_w1916_,
		_w1925_
	);
	LUT3 #(
		.INIT('hd0)
	) name576 (
		\P1_Flush_reg/NET0131 ,
		_w1922_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w1919_,
		_w1926_,
		_w1927_
	);
	LUT3 #(
		.INIT('he0)
	) name578 (
		_w1910_,
		_w1893_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h4500)
	) name579 (
		_w1909_,
		_w1875_,
		_w1907_,
		_w1928_,
		_w1929_
	);
	LUT3 #(
		.INIT('h15)
	) name580 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w1797_,
		_w1859_,
		_w1931_
	);
	LUT4 #(
		.INIT('h1555)
	) name582 (
		\P1_State2_reg[1]/NET0131 ,
		_w1797_,
		_w1859_,
		_w1930_,
		_w1932_
	);
	LUT4 #(
		.INIT('h0020)
	) name583 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		_w1934_
	);
	LUT4 #(
		.INIT('h0040)
	) name585 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1935_
	);
	LUT4 #(
		.INIT('h0008)
	) name586 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1936_
	);
	LUT4 #(
		.INIT('hffb7)
	) name587 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1937_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		_w1861_,
		_w1937_,
		_w1938_
	);
	LUT4 #(
		.INIT('h0004)
	) name589 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1939_
	);
	LUT3 #(
		.INIT('h02)
	) name590 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1940_
	);
	LUT4 #(
		.INIT('h0002)
	) name591 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w1941_
	);
	LUT4 #(
		.INIT('h8caf)
	) name592 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1861_,
		_w1939_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w1938_,
		_w1942_,
		_w1943_
	);
	LUT4 #(
		.INIT('h70ff)
	) name594 (
		_w1929_,
		_w1932_,
		_w1933_,
		_w1943_,
		_w1944_
	);
	LUT4 #(
		.INIT('h0020)
	) name595 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w1945_
	);
	LUT4 #(
		.INIT('h0010)
	) name596 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1946_
	);
	LUT4 #(
		.INIT('h1000)
	) name597 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1947_
	);
	LUT4 #(
		.INIT('h153f)
	) name598 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w1946_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h0040)
	) name599 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1949_
	);
	LUT4 #(
		.INIT('h0100)
	) name600 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1950_
	);
	LUT4 #(
		.INIT('h135f)
	) name601 (
		\P3_InstQueue_reg[6][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT4 #(
		.INIT('h0002)
	) name602 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w1953_
	);
	LUT4 #(
		.INIT('h0080)
	) name604 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1954_
	);
	LUT4 #(
		.INIT('h135f)
	) name605 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1952_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('h0400)
	) name606 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1956_
	);
	LUT4 #(
		.INIT('h0004)
	) name607 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1957_
	);
	LUT4 #(
		.INIT('h135f)
	) name608 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT4 #(
		.INIT('h8000)
	) name609 (
		_w1955_,
		_w1958_,
		_w1948_,
		_w1951_,
		_w1959_
	);
	LUT4 #(
		.INIT('h0800)
	) name610 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1960_
	);
	LUT4 #(
		.INIT('h4000)
	) name611 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1961_
	);
	LUT4 #(
		.INIT('h135f)
	) name612 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h0200)
	) name613 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1963_
	);
	LUT4 #(
		.INIT('h0020)
	) name614 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1964_
	);
	LUT4 #(
		.INIT('h153f)
	) name615 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1963_,
		_w1964_,
		_w1965_
	);
	LUT4 #(
		.INIT('h2000)
	) name616 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1966_
	);
	LUT4 #(
		.INIT('h0008)
	) name617 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1967_
	);
	LUT4 #(
		.INIT('h135f)
	) name618 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h0001)
	) name619 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1969_
	);
	LUT4 #(
		.INIT('h8000)
	) name620 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1970_
	);
	LUT4 #(
		.INIT('h135f)
	) name621 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h8000)
	) name622 (
		_w1968_,
		_w1971_,
		_w1962_,
		_w1965_,
		_w1972_
	);
	LUT4 #(
		.INIT('h135f)
	) name623 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w1956_,
		_w1966_,
		_w1973_
	);
	LUT4 #(
		.INIT('h135f)
	) name624 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1946_,
		_w1950_,
		_w1974_
	);
	LUT4 #(
		.INIT('h153f)
	) name625 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w1952_,
		_w1960_,
		_w1975_
	);
	LUT4 #(
		.INIT('h153f)
	) name626 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1949_,
		_w1970_,
		_w1976_
	);
	LUT4 #(
		.INIT('h8000)
	) name627 (
		_w1975_,
		_w1976_,
		_w1973_,
		_w1974_,
		_w1977_
	);
	LUT4 #(
		.INIT('h135f)
	) name628 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1967_,
		_w1963_,
		_w1978_
	);
	LUT4 #(
		.INIT('h153f)
	) name629 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1954_,
		_w1964_,
		_w1979_
	);
	LUT4 #(
		.INIT('h153f)
	) name630 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1957_,
		_w1961_,
		_w1980_
	);
	LUT4 #(
		.INIT('h153f)
	) name631 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w1947_,
		_w1969_,
		_w1981_
	);
	LUT4 #(
		.INIT('h8000)
	) name632 (
		_w1980_,
		_w1981_,
		_w1978_,
		_w1979_,
		_w1982_
	);
	LUT4 #(
		.INIT('h0777)
	) name633 (
		_w1959_,
		_w1972_,
		_w1977_,
		_w1982_,
		_w1983_
	);
	LUT4 #(
		.INIT('h135f)
	) name634 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w1969_,
		_w1960_,
		_w1984_
	);
	LUT4 #(
		.INIT('h135f)
	) name635 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1952_,
		_w1957_,
		_w1985_
	);
	LUT4 #(
		.INIT('h153f)
	) name636 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1954_,
		_w1966_,
		_w1986_
	);
	LUT4 #(
		.INIT('h135f)
	) name637 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1970_,
		_w1964_,
		_w1987_
	);
	LUT4 #(
		.INIT('h8000)
	) name638 (
		_w1986_,
		_w1987_,
		_w1984_,
		_w1985_,
		_w1988_
	);
	LUT4 #(
		.INIT('h153f)
	) name639 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1949_,
		_w1961_,
		_w1989_
	);
	LUT4 #(
		.INIT('h135f)
	) name640 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1956_,
		_w1950_,
		_w1990_
	);
	LUT4 #(
		.INIT('h135f)
	) name641 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w1947_,
		_w1967_,
		_w1991_
	);
	LUT4 #(
		.INIT('h135f)
	) name642 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1946_,
		_w1963_,
		_w1992_
	);
	LUT4 #(
		.INIT('h8000)
	) name643 (
		_w1991_,
		_w1992_,
		_w1989_,
		_w1990_,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		_w1988_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h153f)
	) name645 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1950_,
		_w1969_,
		_w1995_
	);
	LUT4 #(
		.INIT('h153f)
	) name646 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1952_,
		_w1966_,
		_w1996_
	);
	LUT4 #(
		.INIT('h135f)
	) name647 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1960_,
		_w1964_,
		_w1997_
	);
	LUT4 #(
		.INIT('h135f)
	) name648 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1956_,
		_w1963_,
		_w1998_
	);
	LUT4 #(
		.INIT('h8000)
	) name649 (
		_w1997_,
		_w1998_,
		_w1995_,
		_w1996_,
		_w1999_
	);
	LUT4 #(
		.INIT('h153f)
	) name650 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1954_,
		_w1967_,
		_w2000_
	);
	LUT4 #(
		.INIT('h135f)
	) name651 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1957_,
		_w1949_,
		_w2001_
	);
	LUT4 #(
		.INIT('h153f)
	) name652 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w1946_,
		_w1961_,
		_w2002_
	);
	LUT4 #(
		.INIT('h135f)
	) name653 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w1947_,
		_w1970_,
		_w2003_
	);
	LUT4 #(
		.INIT('h8000)
	) name654 (
		_w2002_,
		_w2003_,
		_w2000_,
		_w2001_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		_w1999_,
		_w2004_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0888)
	) name656 (
		_w1988_,
		_w1993_,
		_w1999_,
		_w2004_,
		_w2006_
	);
	LUT4 #(
		.INIT('h153f)
	) name657 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1954_,
		_w1946_,
		_w2007_
	);
	LUT4 #(
		.INIT('h153f)
	) name658 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w1967_,
		_w1969_,
		_w2008_
	);
	LUT4 #(
		.INIT('h153f)
	) name659 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w1952_,
		_w1956_,
		_w2009_
	);
	LUT4 #(
		.INIT('h153f)
	) name660 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1949_,
		_w1960_,
		_w2010_
	);
	LUT4 #(
		.INIT('h8000)
	) name661 (
		_w2009_,
		_w2010_,
		_w2007_,
		_w2008_,
		_w2011_
	);
	LUT4 #(
		.INIT('h135f)
	) name662 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1957_,
		_w1964_,
		_w2012_
	);
	LUT4 #(
		.INIT('h135f)
	) name663 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1966_,
		_w1963_,
		_w2013_
	);
	LUT4 #(
		.INIT('h135f)
	) name664 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1947_,
		_w1961_,
		_w2014_
	);
	LUT4 #(
		.INIT('h153f)
	) name665 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1950_,
		_w1970_,
		_w2015_
	);
	LUT4 #(
		.INIT('h8000)
	) name666 (
		_w2014_,
		_w2015_,
		_w2012_,
		_w2013_,
		_w2016_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w2011_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h153f)
	) name668 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w1946_,
		_w1947_,
		_w2018_
	);
	LUT4 #(
		.INIT('h153f)
	) name669 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1967_,
		_w1969_,
		_w2019_
	);
	LUT4 #(
		.INIT('h153f)
	) name670 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w1952_,
		_w1970_,
		_w2020_
	);
	LUT4 #(
		.INIT('h135f)
	) name671 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1954_,
		_w1963_,
		_w2021_
	);
	LUT4 #(
		.INIT('h8000)
	) name672 (
		_w2020_,
		_w2021_,
		_w2018_,
		_w2019_,
		_w2022_
	);
	LUT4 #(
		.INIT('h153f)
	) name673 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1957_,
		_w1966_,
		_w2023_
	);
	LUT4 #(
		.INIT('h135f)
	) name674 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w1956_,
		_w1960_,
		_w2024_
	);
	LUT4 #(
		.INIT('h153f)
	) name675 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1950_,
		_w1964_,
		_w2025_
	);
	LUT4 #(
		.INIT('h153f)
	) name676 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1949_,
		_w1961_,
		_w2026_
	);
	LUT4 #(
		.INIT('h8000)
	) name677 (
		_w2025_,
		_w2026_,
		_w2023_,
		_w2024_,
		_w2027_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		_w2022_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h135f)
	) name679 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1960_,
		_w1964_,
		_w2029_
	);
	LUT4 #(
		.INIT('h153f)
	) name680 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1954_,
		_w1961_,
		_w2030_
	);
	LUT4 #(
		.INIT('h153f)
	) name681 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1946_,
		_w1966_,
		_w2031_
	);
	LUT4 #(
		.INIT('h135f)
	) name682 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1947_,
		_w1949_,
		_w2032_
	);
	LUT4 #(
		.INIT('h8000)
	) name683 (
		_w2031_,
		_w2032_,
		_w2029_,
		_w2030_,
		_w2033_
	);
	LUT4 #(
		.INIT('h135f)
	) name684 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1969_,
		_w1963_,
		_w2034_
	);
	LUT4 #(
		.INIT('h135f)
	) name685 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1956_,
		_w1970_,
		_w2035_
	);
	LUT4 #(
		.INIT('h135f)
	) name686 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1957_,
		_w1950_,
		_w2036_
	);
	LUT4 #(
		.INIT('h135f)
	) name687 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1952_,
		_w1967_,
		_w2037_
	);
	LUT4 #(
		.INIT('h8000)
	) name688 (
		_w2036_,
		_w2037_,
		_w2034_,
		_w2035_,
		_w2038_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		_w2033_,
		_w2038_,
		_w2039_
	);
	LUT4 #(
		.INIT('h0777)
	) name690 (
		_w2022_,
		_w2027_,
		_w2033_,
		_w2038_,
		_w2040_
	);
	LUT4 #(
		.INIT('h8000)
	) name691 (
		_w2017_,
		_w1983_,
		_w2006_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('h7000)
	) name692 (
		_w2011_,
		_w2016_,
		_w2022_,
		_w2027_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		_w2039_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h8000)
	) name694 (
		_w2039_,
		_w2042_,
		_w1983_,
		_w2006_,
		_w2044_
	);
	LUT4 #(
		.INIT('h0888)
	) name695 (
		_w1959_,
		_w1972_,
		_w1977_,
		_w1982_,
		_w2045_
	);
	LUT4 #(
		.INIT('h8000)
	) name696 (
		_w1988_,
		_w1993_,
		_w1999_,
		_w2004_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8000)
	) name697 (
		_w2045_,
		_w2017_,
		_w2046_,
		_w2040_,
		_w2047_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w2044_,
		_w2047_,
		_w2048_
	);
	LUT4 #(
		.INIT('h8000)
	) name699 (
		_w2011_,
		_w2016_,
		_w2022_,
		_w2027_,
		_w2049_
	);
	LUT4 #(
		.INIT('h135f)
	) name700 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1956_,
		_w1967_,
		_w2050_
	);
	LUT4 #(
		.INIT('h135f)
	) name701 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1947_,
		_w1950_,
		_w2051_
	);
	LUT4 #(
		.INIT('h153f)
	) name702 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w1952_,
		_w1960_,
		_w2052_
	);
	LUT4 #(
		.INIT('h153f)
	) name703 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1946_,
		_w1961_,
		_w2053_
	);
	LUT4 #(
		.INIT('h8000)
	) name704 (
		_w2052_,
		_w2053_,
		_w2050_,
		_w2051_,
		_w2054_
	);
	LUT4 #(
		.INIT('h153f)
	) name705 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1949_,
		_w1964_,
		_w2055_
	);
	LUT4 #(
		.INIT('h135f)
	) name706 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1966_,
		_w1970_,
		_w2056_
	);
	LUT4 #(
		.INIT('h135f)
	) name707 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1957_,
		_w1963_,
		_w2057_
	);
	LUT4 #(
		.INIT('h153f)
	) name708 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1954_,
		_w1969_,
		_w2058_
	);
	LUT4 #(
		.INIT('h8000)
	) name709 (
		_w2057_,
		_w2058_,
		_w2055_,
		_w2056_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name710 (
		_w2054_,
		_w2059_,
		_w2060_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		_w2049_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h8000)
	) name712 (
		_w1999_,
		_w2004_,
		_w2033_,
		_w2038_,
		_w2062_
	);
	LUT3 #(
		.INIT('h80)
	) name713 (
		_w2049_,
		_w2060_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h8000)
	) name714 (
		_w2049_,
		_w2060_,
		_w2062_,
		_w1983_,
		_w2064_
	);
	LUT3 #(
		.INIT('h01)
	) name715 (
		_w2044_,
		_w2047_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h0001)
	) name716 (
		_w2041_,
		_w2044_,
		_w2047_,
		_w2064_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name717 (
		_w2045_,
		_w1994_,
		_w2067_
	);
	LUT3 #(
		.INIT('h02)
	) name718 (
		_w2045_,
		_w1994_,
		_w2005_,
		_w2068_
	);
	LUT4 #(
		.INIT('h0888)
	) name719 (
		_w2011_,
		_w2016_,
		_w2054_,
		_w2059_,
		_w2069_
	);
	LUT4 #(
		.INIT('h0200)
	) name720 (
		_w2045_,
		_w1994_,
		_w2005_,
		_w2040_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT4 #(
		.INIT('h5777)
	) name722 (
		_w2068_,
		_w2061_,
		_w2069_,
		_w2040_,
		_w2072_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		_w2066_,
		_w2072_,
		_w2073_
	);
	LUT4 #(
		.INIT('h7000)
	) name724 (
		_w1959_,
		_w1972_,
		_w1977_,
		_w1982_,
		_w2074_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		_w1994_,
		_w2074_,
		_w2075_
	);
	LUT3 #(
		.INIT('h20)
	) name726 (
		_w1994_,
		_w2005_,
		_w2074_,
		_w2076_
	);
	LUT4 #(
		.INIT('h2000)
	) name727 (
		_w2049_,
		_w2039_,
		_w1983_,
		_w2006_,
		_w2077_
	);
	LUT4 #(
		.INIT('h5540)
	) name728 (
		_w2060_,
		_w2043_,
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT4 #(
		.INIT('h8000)
	) name729 (
		_w1959_,
		_w1972_,
		_w1977_,
		_w1982_,
		_w2079_
	);
	LUT4 #(
		.INIT('h7000)
	) name730 (
		_w2011_,
		_w2016_,
		_w2054_,
		_w2059_,
		_w2080_
	);
	LUT3 #(
		.INIT('h80)
	) name731 (
		_w2046_,
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('hf800)
	) name732 (
		_w2068_,
		_w2061_,
		_w2081_,
		_w2039_,
		_w2082_
	);
	LUT3 #(
		.INIT('h40)
	) name733 (
		_w2028_,
		_w2062_,
		_w2069_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		_w2075_,
		_w2083_,
		_w2084_
	);
	LUT4 #(
		.INIT('h0737)
	) name735 (
		_w2067_,
		_w2063_,
		_w2075_,
		_w2083_,
		_w2085_
	);
	LUT3 #(
		.INIT('h10)
	) name736 (
		_w2082_,
		_w2078_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('h08)
	) name737 (
		_w2068_,
		_w2061_,
		_w2039_,
		_w2087_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2088_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2089_
	);
	LUT4 #(
		.INIT('h08ce)
	) name740 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2090_
	);
	LUT3 #(
		.INIT('hb2)
	) name741 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('h040d)
	) name742 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2089_,
		_w2090_,
		_w2092_
	);
	LUT2 #(
		.INIT('h9)
	) name743 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2093_
	);
	LUT2 #(
		.INIT('h9)
	) name744 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2094_
	);
	LUT2 #(
		.INIT('h9)
	) name745 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2095_
	);
	LUT4 #(
		.INIT('h8421)
	) name746 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2096_
	);
	LUT3 #(
		.INIT('h09)
	) name747 (
		_w2090_,
		_w2094_,
		_w2096_,
		_w2097_
	);
	LUT4 #(
		.INIT('h4d04)
	) name748 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2091_,
		_w2097_,
		_w2098_
	);
	LUT3 #(
		.INIT('he0)
	) name749 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h6)
	) name750 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2100_
	);
	LUT4 #(
		.INIT('hfb00)
	) name751 (
		_w2073_,
		_w2086_,
		_w2099_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h4290)
	) name752 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2093_,
		_w2090_,
		_w2102_
	);
	LUT3 #(
		.INIT('h32)
	) name753 (
		_w2088_,
		_w2102_,
		_w2092_,
		_w2103_
	);
	LUT4 #(
		.INIT('h39c6)
	) name754 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2104_
	);
	LUT4 #(
		.INIT('h05cd)
	) name755 (
		_w2088_,
		_w2102_,
		_w2092_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w2060_,
		_w2047_,
		_w2106_
	);
	LUT3 #(
		.INIT('h27)
	) name757 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2107_
	);
	LUT4 #(
		.INIT('h00d8)
	) name758 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w2108_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w2109_
	);
	LUT3 #(
		.INIT('h04)
	) name760 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w2110_
	);
	LUT3 #(
		.INIT('heb)
	) name761 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w2111_,
		_w2105_,
		_w2112_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w2060_,
		_w2047_,
		_w2113_
	);
	LUT3 #(
		.INIT('h1b)
	) name764 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2114_
	);
	LUT4 #(
		.INIT('he400)
	) name765 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2112_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2116_
	);
	LUT4 #(
		.INIT('h5501)
	) name767 (
		_w2064_,
		_w2108_,
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w2105_,
		_w2116_,
		_w2119_
	);
	LUT3 #(
		.INIT('h04)
	) name770 (
		_w2060_,
		_w2047_,
		_w2119_,
		_w2120_
	);
	LUT3 #(
		.INIT('h08)
	) name771 (
		_w2060_,
		_w2044_,
		_w2119_,
		_w2121_
	);
	LUT4 #(
		.INIT('hff27)
	) name772 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2119_,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w2111_,
		_w2116_,
		_w2123_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w2105_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('h00e4)
	) name775 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name776 (
		_w2122_,
		_w2125_,
		_w2126_
	);
	LUT3 #(
		.INIT('h0e)
	) name777 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2127_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2041_,
		_w2128_
	);
	LUT3 #(
		.INIT('h20)
	) name779 (
		_w2126_,
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT4 #(
		.INIT('h4445)
	) name780 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2101_,
		_w2118_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h0010)
	) name781 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2073_,
		_w2086_,
		_w2099_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2066_,
		_w2132_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w2127_,
		_w2132_,
		_w2133_
	);
	LUT3 #(
		.INIT('ha8)
	) name784 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2131_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h4)
	) name785 (
		_w2130_,
		_w2134_,
		_w2135_
	);
	LUT4 #(
		.INIT('hd800)
	) name786 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w2136_
	);
	LUT4 #(
		.INIT('h031b)
	) name787 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w2137_
	);
	LUT4 #(
		.INIT('h888a)
	) name788 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2041_,
		_w2112_,
		_w2137_,
		_w2138_
	);
	LUT3 #(
		.INIT('h07)
	) name789 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2139_
	);
	LUT3 #(
		.INIT('h78)
	) name790 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2140_
	);
	LUT3 #(
		.INIT('hb0)
	) name791 (
		_w2073_,
		_w2086_,
		_w2140_,
		_w2141_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2142_
	);
	LUT2 #(
		.INIT('h6)
	) name793 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2143_
	);
	LUT4 #(
		.INIT('hc666)
	) name794 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2144_
	);
	LUT3 #(
		.INIT('he0)
	) name795 (
		_w2108_,
		_w2115_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w2064_,
		_w2143_,
		_w2146_
	);
	LUT3 #(
		.INIT('h9a)
	) name797 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1953_,
		_w2098_,
		_w2147_
	);
	LUT4 #(
		.INIT('h0133)
	) name798 (
		_w2071_,
		_w2146_,
		_w2087_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name799 (
		_w2145_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h0200)
	) name800 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2141_,
		_w2138_,
		_w2149_,
		_w2150_
	);
	LUT4 #(
		.INIT('h88c8)
	) name801 (
		_w2064_,
		_w2142_,
		_w2108_,
		_w2116_,
		_w2151_
	);
	LUT4 #(
		.INIT('h0027)
	) name802 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2064_,
		_w2152_
	);
	LUT3 #(
		.INIT('h80)
	) name803 (
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2153_
	);
	LUT4 #(
		.INIT('h5444)
	) name804 (
		_w2041_,
		_w2152_,
		_w2122_,
		_w2153_,
		_w2154_
	);
	LUT3 #(
		.INIT('h0e)
	) name805 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2151_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('h807f)
	) name806 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2156_
	);
	LUT4 #(
		.INIT('h6555)
	) name807 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2105_,
		_w2142_,
		_w2123_,
		_w2157_
	);
	LUT4 #(
		.INIT('h00e4)
	) name808 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2157_,
		_w2158_
	);
	LUT3 #(
		.INIT('h9a)
	) name809 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2139_,
		_w2098_,
		_w2159_
	);
	LUT4 #(
		.INIT('h010f)
	) name810 (
		_w2071_,
		_w2087_,
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('hf400)
	) name811 (
		_w2073_,
		_w2086_,
		_w2156_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w2155_,
		_w2161_,
		_w2162_
	);
	LUT3 #(
		.INIT('h20)
	) name813 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2155_,
		_w2161_,
		_w2163_
	);
	LUT4 #(
		.INIT('h2220)
	) name814 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2101_,
		_w2118_,
		_w2129_,
		_w2164_
	);
	LUT3 #(
		.INIT('h01)
	) name815 (
		_w2163_,
		_w2164_,
		_w2150_,
		_w2165_
	);
	LUT4 #(
		.INIT('h5455)
	) name816 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2141_,
		_w2138_,
		_w2149_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w2163_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('h0200)
	) name818 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2141_,
		_w2138_,
		_w2149_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		\P3_More_reg/NET0131 ,
		_w2105_,
		_w2169_
	);
	LUT3 #(
		.INIT('h0d)
	) name820 (
		_w2122_,
		_w2125_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w2060_,
		_w2041_,
		_w2171_
	);
	LUT4 #(
		.INIT('h00e0)
	) name822 (
		_w2088_,
		_w2092_,
		_w2104_,
		_w2095_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w2103_,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('h40)
	) name824 (
		_w2060_,
		_w2041_,
		_w2173_,
		_w2174_
	);
	LUT3 #(
		.INIT('h08)
	) name825 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w2175_
	);
	LUT4 #(
		.INIT('h00f1)
	) name826 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('he400)
	) name827 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2111_,
		_w2177_
	);
	LUT3 #(
		.INIT('hf1)
	) name828 (
		_w2044_,
		_w2047_,
		_w2105_,
		_w2178_
	);
	LUT4 #(
		.INIT('h00a8)
	) name829 (
		\P3_Flush_reg/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w2179_
	);
	LUT3 #(
		.INIT('h04)
	) name830 (
		_w2060_,
		_w2041_,
		_w2173_,
		_w2180_
	);
	LUT3 #(
		.INIT('h80)
	) name831 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w2181_
	);
	LUT4 #(
		.INIT('h7f3b)
	) name832 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w2173_,
		_w2182_
	);
	LUT4 #(
		.INIT('h1f00)
	) name833 (
		_w2116_,
		_w2177_,
		_w2179_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h1000)
	) name834 (
		_w2170_,
		_w2174_,
		_w2176_,
		_w2183_,
		_w2184_
	);
	LUT3 #(
		.INIT('he0)
	) name835 (
		_w2168_,
		_w2162_,
		_w2184_,
		_w2185_
	);
	LUT4 #(
		.INIT('h4500)
	) name836 (
		_w2167_,
		_w2135_,
		_w2165_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('h15)
	) name837 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2187_
	);
	LUT3 #(
		.INIT('h10)
	) name838 (
		_w2111_,
		_w2105_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h80)
	) name839 (
		_w2060_,
		_w2047_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2190_
	);
	LUT3 #(
		.INIT('h02)
	) name841 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2191_
	);
	LUT4 #(
		.INIT('h0048)
	) name842 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		_w2116_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h0004)
	) name844 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2194_
	);
	LUT4 #(
		.INIT('h0002)
	) name845 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2195_
	);
	LUT4 #(
		.INIT('h8caf)
	) name846 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2116_,
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		_w2193_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name848 (
		_w1945_,
		_w2186_,
		_w2189_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w2199_
	);
	LUT4 #(
		.INIT('h0008)
	) name850 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2200_
	);
	LUT4 #(
		.INIT('hff8f)
	) name851 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2201_
	);
	LUT3 #(
		.INIT('hb0)
	) name852 (
		_w2116_,
		_w2200_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('hb)
	) name853 (
		_w2199_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h1000)
	) name854 (
		_w1654_,
		_w1652_,
		_w1672_,
		_w1676_,
		_w2204_
	);
	LUT4 #(
		.INIT('h0080)
	) name855 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2205_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2206_
	);
	LUT3 #(
		.INIT('he0)
	) name857 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2207_
	);
	LUT3 #(
		.INIT('h2a)
	) name858 (
		_w2205_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name859 (
		_w1605_,
		_w1681_,
		_w2209_
	);
	LUT4 #(
		.INIT('h8000)
	) name860 (
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w2210_
	);
	LUT4 #(
		.INIT('h0200)
	) name861 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2211_
	);
	LUT3 #(
		.INIT('h0d)
	) name862 (
		_w1683_,
		_w2210_,
		_w2211_,
		_w2212_
	);
	LUT3 #(
		.INIT('h10)
	) name863 (
		_w2208_,
		_w2209_,
		_w2212_,
		_w2213_
	);
	LUT3 #(
		.INIT('h2f)
	) name864 (
		_w1678_,
		_w2204_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h0100)
	) name865 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2215_
	);
	LUT4 #(
		.INIT('h0080)
	) name866 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2216_
	);
	LUT4 #(
		.INIT('h0180)
	) name867 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2217_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name868 (
		\P3_State2_reg[0]/NET0131 ,
		_w2111_,
		_w2105_,
		_w2187_,
		_w2218_
	);
	LUT3 #(
		.INIT('h08)
	) name869 (
		_w2060_,
		_w2047_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2220_
	);
	LUT3 #(
		.INIT('he0)
	) name871 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2221_
	);
	LUT3 #(
		.INIT('h2a)
	) name872 (
		_w2216_,
		_w2220_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h8000)
	) name873 (
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w2190_,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('h0200)
	) name875 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w2225_
	);
	LUT3 #(
		.INIT('h07)
	) name876 (
		_w2116_,
		_w2191_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h10)
	) name877 (
		_w2224_,
		_w2222_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('h2aff)
	) name878 (
		_w1945_,
		_w2186_,
		_w2219_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h7f00)
	) name879 (
		_w1797_,
		_w1859_,
		_w1930_,
		_w1933_,
		_w2229_
	);
	LUT4 #(
		.INIT('h0080)
	) name880 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2230_
	);
	LUT2 #(
		.INIT('h4)
	) name881 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2231_
	);
	LUT3 #(
		.INIT('he0)
	) name882 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2232_
	);
	LUT3 #(
		.INIT('h2a)
	) name883 (
		_w2230_,
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT4 #(
		.INIT('h0200)
	) name884 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2234_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2235_
	);
	LUT4 #(
		.INIT('h085f)
	) name886 (
		_w1861_,
		_w1934_,
		_w1940_,
		_w2235_,
		_w2236_
	);
	LUT3 #(
		.INIT('h10)
	) name887 (
		_w2233_,
		_w2234_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		_w2229_,
		_w2237_,
		_w2238_
	);
	LUT3 #(
		.INIT('h4f)
	) name889 (
		_w1929_,
		_w1933_,
		_w2238_,
		_w2239_
	);
	LUT4 #(
		.INIT('h0008)
	) name890 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2240_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		_w1605_,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2242_
	);
	LUT4 #(
		.INIT('hff8f)
	) name893 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2243_
	);
	LUT3 #(
		.INIT('h70)
	) name894 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('hb)
	) name895 (
		_w2241_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('h0100)
	) name896 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2246_
	);
	LUT4 #(
		.INIT('h0180)
	) name897 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2247_
	);
	LUT4 #(
		.INIT('h0100)
	) name898 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2248_
	);
	LUT4 #(
		.INIT('h0180)
	) name899 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2249_
	);
	LUT4 #(
		.INIT('h0100)
	) name900 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2250_
	);
	LUT4 #(
		.INIT('h0001)
	) name901 (
		\P2_Address_reg[26]/NET0131 ,
		\P2_Address_reg[27]/NET0131 ,
		\P2_Address_reg[28]/NET0131 ,
		\P2_Address_reg[2]/NET0131 ,
		_w2251_
	);
	LUT4 #(
		.INIT('h0001)
	) name902 (
		\P2_Address_reg[22]/NET0131 ,
		\P2_Address_reg[23]/NET0131 ,
		\P2_Address_reg[24]/NET0131 ,
		\P2_Address_reg[25]/NET0131 ,
		_w2252_
	);
	LUT3 #(
		.INIT('h01)
	) name903 (
		\P2_Address_reg[7]/NET0131 ,
		\P2_Address_reg[8]/NET0131 ,
		\P2_Address_reg[9]/NET0131 ,
		_w2253_
	);
	LUT4 #(
		.INIT('h0001)
	) name904 (
		\P2_Address_reg[3]/NET0131 ,
		\P2_Address_reg[4]/NET0131 ,
		\P2_Address_reg[5]/NET0131 ,
		\P2_Address_reg[6]/NET0131 ,
		_w2254_
	);
	LUT4 #(
		.INIT('h8000)
	) name905 (
		_w2253_,
		_w2254_,
		_w2251_,
		_w2252_,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		\P2_Address_reg[0]/NET0131 ,
		\P2_Address_reg[10]/NET0131 ,
		_w2256_
	);
	LUT4 #(
		.INIT('h0001)
	) name907 (
		\P2_Address_reg[11]/NET0131 ,
		\P2_Address_reg[12]/NET0131 ,
		\P2_Address_reg[13]/NET0131 ,
		\P2_Address_reg[14]/NET0131 ,
		_w2257_
	);
	LUT4 #(
		.INIT('h0001)
	) name908 (
		\P2_Address_reg[19]/NET0131 ,
		\P2_Address_reg[1]/NET0131 ,
		\P2_Address_reg[20]/NET0131 ,
		\P2_Address_reg[21]/NET0131 ,
		_w2258_
	);
	LUT4 #(
		.INIT('h0001)
	) name909 (
		\P2_Address_reg[15]/NET0131 ,
		\P2_Address_reg[16]/NET0131 ,
		\P2_Address_reg[17]/NET0131 ,
		\P2_Address_reg[18]/NET0131 ,
		_w2259_
	);
	LUT4 #(
		.INIT('h8000)
	) name910 (
		_w2256_,
		_w2258_,
		_w2259_,
		_w2257_,
		_w2260_
	);
	LUT4 #(
		.INIT('hc444)
	) name911 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h0888)
	) name912 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[28]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2262_
	);
	LUT3 #(
		.INIT('ha8)
	) name913 (
		_w2250_,
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h0200)
	) name914 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2264_
	);
	LUT4 #(
		.INIT('hc444)
	) name915 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[20]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2265_
	);
	LUT4 #(
		.INIT('h0888)
	) name916 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[20]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT3 #(
		.INIT('ha8)
	) name918 (
		_w2264_,
		_w2265_,
		_w2266_,
		_w2268_
	);
	LUT3 #(
		.INIT('ha8)
	) name919 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2263_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2270_
	);
	LUT4 #(
		.INIT('h0400)
	) name921 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2271_
	);
	LUT4 #(
		.INIT('h0800)
	) name922 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2272_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name923 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2273_
	);
	LUT4 #(
		.INIT('hc444)
	) name924 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2274_
	);
	LUT4 #(
		.INIT('h0888)
	) name925 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[4]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT3 #(
		.INIT('h02)
	) name927 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w2271_,
		_w2272_,
		_w2277_
	);
	LUT4 #(
		.INIT('h00ab)
	) name928 (
		_w2273_,
		_w2274_,
		_w2275_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('hfcff)
	) name929 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w2278_,
		_w2280_,
		_w2281_
	);
	LUT3 #(
		.INIT('ha8)
	) name932 (
		_w1679_,
		_w2269_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('h0010)
	) name933 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2283_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		_w2278_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('hc055)
	) name935 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2272_,
		_w2285_
	);
	LUT4 #(
		.INIT('h0001)
	) name936 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2286_
	);
	LUT4 #(
		.INIT('hfffc)
	) name937 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2287_
	);
	LUT4 #(
		.INIT('hfd14)
	) name938 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2288_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		_w2288_,
		_w2289_
	);
	LUT3 #(
		.INIT('h0d)
	) name940 (
		_w2246_,
		_w2285_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w2284_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('hb)
	) name942 (
		_w2282_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('hc444)
	) name943 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2293_
	);
	LUT4 #(
		.INIT('h0888)
	) name944 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[7]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2294_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT3 #(
		.INIT('h02)
	) name946 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w2271_,
		_w2272_,
		_w2296_
	);
	LUT4 #(
		.INIT('h00ab)
	) name947 (
		_w2273_,
		_w2293_,
		_w2294_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('hffeb)
	) name948 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w2298_
	);
	LUT4 #(
		.INIT('h00fd)
	) name949 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2279_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w2297_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('hc055)
	) name951 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2272_,
		_w2301_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		_w2288_,
		_w2302_
	);
	LUT4 #(
		.INIT('hc444)
	) name953 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2303_
	);
	LUT4 #(
		.INIT('h0888)
	) name954 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[23]/NET0131 ,
		_w2255_,
		_w2260_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT3 #(
		.INIT('h80)
	) name956 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2264_,
		_w2306_
	);
	LUT4 #(
		.INIT('h0155)
	) name957 (
		_w2302_,
		_w2303_,
		_w2304_,
		_w2306_,
		_w2307_
	);
	LUT3 #(
		.INIT('hd0)
	) name958 (
		_w2246_,
		_w2301_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('hb)
	) name959 (
		_w2300_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w2310_
	);
	LUT4 #(
		.INIT('hff8f)
	) name961 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w2311_
	);
	LUT3 #(
		.INIT('hb0)
	) name962 (
		_w1861_,
		_w1936_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w2310_,
		_w2312_,
		_w2313_
	);
	LUT3 #(
		.INIT('h4f)
	) name964 (
		_w1929_,
		_w1933_,
		_w2313_,
		_w2314_
	);
	LUT4 #(
		.INIT('h2000)
	) name965 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2315_
	);
	LUT3 #(
		.INIT('he0)
	) name966 (
		_w2261_,
		_w2262_,
		_w2315_,
		_w2316_
	);
	LUT4 #(
		.INIT('h4000)
	) name967 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2317_
	);
	LUT3 #(
		.INIT('he0)
	) name968 (
		_w2265_,
		_w2266_,
		_w2317_,
		_w2318_
	);
	LUT3 #(
		.INIT('ha8)
	) name969 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2316_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('h0001)
	) name970 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2320_
	);
	LUT3 #(
		.INIT('h80)
	) name971 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2321_
	);
	LUT4 #(
		.INIT('h8000)
	) name972 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2322_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name973 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2323_
	);
	LUT3 #(
		.INIT('h02)
	) name974 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w2320_,
		_w2322_,
		_w2324_
	);
	LUT4 #(
		.INIT('h00f1)
	) name975 (
		_w2274_,
		_w2275_,
		_w2323_,
		_w2324_,
		_w2325_
	);
	LUT4 #(
		.INIT('h9fff)
	) name976 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2326_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w2325_,
		_w2327_,
		_w2328_
	);
	LUT3 #(
		.INIT('ha8)
	) name979 (
		_w1679_,
		_w2319_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		_w2283_,
		_w2325_,
		_w2330_
	);
	LUT4 #(
		.INIT('hc055)
	) name981 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2320_,
		_w2331_
	);
	LUT2 #(
		.INIT('h2)
	) name982 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		_w2288_,
		_w2332_
	);
	LUT3 #(
		.INIT('h0d)
	) name983 (
		_w2246_,
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h4)
	) name984 (
		_w2330_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('hb)
	) name985 (
		_w2329_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('h02)
	) name986 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w2320_,
		_w2322_,
		_w2336_
	);
	LUT4 #(
		.INIT('h00f1)
	) name987 (
		_w2293_,
		_w2294_,
		_w2323_,
		_w2336_,
		_w2337_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name988 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2326_,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT4 #(
		.INIT('hc055)
	) name990 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2320_,
		_w2340_
	);
	LUT2 #(
		.INIT('h2)
	) name991 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		_w2288_,
		_w2341_
	);
	LUT3 #(
		.INIT('h80)
	) name992 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2317_,
		_w2342_
	);
	LUT4 #(
		.INIT('h010f)
	) name993 (
		_w2303_,
		_w2304_,
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT3 #(
		.INIT('hd0)
	) name994 (
		_w2246_,
		_w2340_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('hb)
	) name995 (
		_w2339_,
		_w2344_,
		_w2345_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name996 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2346_
	);
	LUT3 #(
		.INIT('h02)
	) name997 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w2271_,
		_w2264_,
		_w2347_
	);
	LUT4 #(
		.INIT('h00f1)
	) name998 (
		_w2293_,
		_w2294_,
		_w2346_,
		_w2347_,
		_w2348_
	);
	LUT4 #(
		.INIT('h0080)
	) name999 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2349_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name1000 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2350_
	);
	LUT2 #(
		.INIT('h2)
	) name1001 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2350_,
		_w2351_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1002 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2350_,
		_w2352_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w2348_,
		_w2352_,
		_w2353_
	);
	LUT4 #(
		.INIT('hc055)
	) name1004 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2271_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w2288_,
		_w2355_
	);
	LUT3 #(
		.INIT('h80)
	) name1006 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2250_,
		_w2356_
	);
	LUT4 #(
		.INIT('h010f)
	) name1007 (
		_w2303_,
		_w2304_,
		_w2355_,
		_w2356_,
		_w2357_
	);
	LUT3 #(
		.INIT('hd0)
	) name1008 (
		_w2246_,
		_w2354_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('hb)
	) name1009 (
		_w2353_,
		_w2358_,
		_w2359_
	);
	LUT3 #(
		.INIT('ha8)
	) name1010 (
		_w2250_,
		_w2265_,
		_w2266_,
		_w2360_
	);
	LUT3 #(
		.INIT('he0)
	) name1011 (
		_w2261_,
		_w2262_,
		_w2349_,
		_w2361_
	);
	LUT3 #(
		.INIT('ha8)
	) name1012 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2360_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('h02)
	) name1013 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w2271_,
		_w2264_,
		_w2363_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1014 (
		_w2274_,
		_w2275_,
		_w2346_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w2351_,
		_w2364_,
		_w2365_
	);
	LUT3 #(
		.INIT('ha8)
	) name1016 (
		_w1679_,
		_w2362_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		_w2283_,
		_w2364_,
		_w2367_
	);
	LUT4 #(
		.INIT('hc055)
	) name1018 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2271_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1019 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		_w2288_,
		_w2369_
	);
	LUT3 #(
		.INIT('h0d)
	) name1020 (
		_w2246_,
		_w2368_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h4)
	) name1021 (
		_w2367_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('hb)
	) name1022 (
		_w2366_,
		_w2371_,
		_w2372_
	);
	LUT3 #(
		.INIT('he0)
	) name1023 (
		_w2261_,
		_w2262_,
		_w2264_,
		_w2373_
	);
	LUT3 #(
		.INIT('ha8)
	) name1024 (
		_w2271_,
		_w2265_,
		_w2266_,
		_w2374_
	);
	LUT3 #(
		.INIT('ha8)
	) name1025 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2373_,
		_w2374_,
		_w2375_
	);
	LUT4 #(
		.INIT('h1000)
	) name1026 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2376_
	);
	LUT4 #(
		.INIT('he7ff)
	) name1027 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2377_
	);
	LUT3 #(
		.INIT('h02)
	) name1028 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w2272_,
		_w2376_,
		_w2378_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1029 (
		_w2274_,
		_w2275_,
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2346_,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT3 #(
		.INIT('ha8)
	) name1032 (
		_w1679_,
		_w2375_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		_w2283_,
		_w2379_,
		_w2383_
	);
	LUT4 #(
		.INIT('hc055)
	) name1034 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2376_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1035 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w2288_,
		_w2385_
	);
	LUT3 #(
		.INIT('h0d)
	) name1036 (
		_w2246_,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		_w2383_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('hb)
	) name1038 (
		_w2382_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h02)
	) name1039 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w2272_,
		_w2376_,
		_w2389_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1040 (
		_w2293_,
		_w2294_,
		_w2377_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1041 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2346_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('hc055)
	) name1043 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2376_,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		_w2288_,
		_w2394_
	);
	LUT3 #(
		.INIT('h80)
	) name1045 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2271_,
		_w2395_
	);
	LUT4 #(
		.INIT('h010f)
	) name1046 (
		_w2303_,
		_w2304_,
		_w2394_,
		_w2395_,
		_w2396_
	);
	LUT3 #(
		.INIT('hd0)
	) name1047 (
		_w2246_,
		_w2393_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('hb)
	) name1048 (
		_w2392_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('ha8)
	) name1049 (
		_w2271_,
		_w2261_,
		_w2262_,
		_w2399_
	);
	LUT3 #(
		.INIT('ha8)
	) name1050 (
		_w2272_,
		_w2265_,
		_w2266_,
		_w2400_
	);
	LUT3 #(
		.INIT('ha8)
	) name1051 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2399_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('hcfff)
	) name1052 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2402_
	);
	LUT3 #(
		.INIT('h02)
	) name1053 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w2315_,
		_w2376_,
		_w2403_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1054 (
		_w2274_,
		_w2275_,
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2273_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w2404_,
		_w2405_,
		_w2406_
	);
	LUT3 #(
		.INIT('ha8)
	) name1057 (
		_w1679_,
		_w2401_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name1058 (
		_w2283_,
		_w2404_,
		_w2408_
	);
	LUT4 #(
		.INIT('hc055)
	) name1059 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2315_,
		_w2409_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w2288_,
		_w2410_
	);
	LUT3 #(
		.INIT('h0d)
	) name1061 (
		_w2246_,
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w2408_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('hb)
	) name1063 (
		_w2407_,
		_w2412_,
		_w2413_
	);
	LUT3 #(
		.INIT('h02)
	) name1064 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w2315_,
		_w2376_,
		_w2414_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1065 (
		_w2293_,
		_w2294_,
		_w2402_,
		_w2414_,
		_w2415_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1066 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2273_,
		_w2283_,
		_w2298_,
		_w2416_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w2415_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('hc055)
	) name1068 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2315_,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name1069 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		_w2288_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name1070 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2272_,
		_w2420_
	);
	LUT4 #(
		.INIT('h010f)
	) name1071 (
		_w2303_,
		_w2304_,
		_w2419_,
		_w2420_,
		_w2421_
	);
	LUT3 #(
		.INIT('hd0)
	) name1072 (
		_w2246_,
		_w2418_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('hb)
	) name1073 (
		_w2417_,
		_w2422_,
		_w2423_
	);
	LUT3 #(
		.INIT('ha8)
	) name1074 (
		_w2272_,
		_w2261_,
		_w2262_,
		_w2424_
	);
	LUT3 #(
		.INIT('he0)
	) name1075 (
		_w2265_,
		_w2266_,
		_w2376_,
		_w2425_
	);
	LUT3 #(
		.INIT('ha8)
	) name1076 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2424_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('h02)
	) name1077 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w2315_,
		_w2317_,
		_w2427_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1078 (
		_w2274_,
		_w2275_,
		_w2326_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h2)
	) name1079 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2377_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT3 #(
		.INIT('ha8)
	) name1081 (
		_w1679_,
		_w2426_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name1082 (
		_w2283_,
		_w2428_,
		_w2432_
	);
	LUT4 #(
		.INIT('hc055)
	) name1083 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2317_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name1084 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w2288_,
		_w2434_
	);
	LUT3 #(
		.INIT('h0d)
	) name1085 (
		_w2246_,
		_w2433_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w2432_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('hb)
	) name1087 (
		_w2431_,
		_w2436_,
		_w2437_
	);
	LUT3 #(
		.INIT('h02)
	) name1088 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w2315_,
		_w2317_,
		_w2438_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1089 (
		_w2293_,
		_w2294_,
		_w2326_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1090 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2377_,
		_w2440_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w2439_,
		_w2440_,
		_w2441_
	);
	LUT4 #(
		.INIT('hc055)
	) name1092 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2317_,
		_w2442_
	);
	LUT2 #(
		.INIT('h2)
	) name1093 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w2288_,
		_w2443_
	);
	LUT3 #(
		.INIT('h80)
	) name1094 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2376_,
		_w2444_
	);
	LUT4 #(
		.INIT('h010f)
	) name1095 (
		_w2303_,
		_w2304_,
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT3 #(
		.INIT('hd0)
	) name1096 (
		_w2246_,
		_w2442_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('hb)
	) name1097 (
		_w2441_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('he0)
	) name1098 (
		_w2261_,
		_w2262_,
		_w2376_,
		_w2448_
	);
	LUT3 #(
		.INIT('he0)
	) name1099 (
		_w2265_,
		_w2266_,
		_w2315_,
		_w2449_
	);
	LUT3 #(
		.INIT('ha8)
	) name1100 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT4 #(
		.INIT('h3fff)
	) name1101 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2451_
	);
	LUT3 #(
		.INIT('h02)
	) name1102 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w2322_,
		_w2317_,
		_w2452_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1103 (
		_w2274_,
		_w2275_,
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name1104 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2402_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT3 #(
		.INIT('ha8)
	) name1106 (
		_w1679_,
		_w2450_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		_w2283_,
		_w2453_,
		_w2457_
	);
	LUT4 #(
		.INIT('hc055)
	) name1108 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2322_,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w2288_,
		_w2459_
	);
	LUT3 #(
		.INIT('h0d)
	) name1110 (
		_w2246_,
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name1111 (
		_w2457_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('hb)
	) name1112 (
		_w2456_,
		_w2461_,
		_w2462_
	);
	LUT3 #(
		.INIT('h02)
	) name1113 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w2322_,
		_w2317_,
		_w2463_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1114 (
		_w2293_,
		_w2294_,
		_w2451_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1115 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2402_,
		_w2465_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT4 #(
		.INIT('hc055)
	) name1117 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2322_,
		_w2467_
	);
	LUT2 #(
		.INIT('h2)
	) name1118 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w2288_,
		_w2468_
	);
	LUT3 #(
		.INIT('h80)
	) name1119 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2315_,
		_w2469_
	);
	LUT4 #(
		.INIT('h010f)
	) name1120 (
		_w2303_,
		_w2304_,
		_w2468_,
		_w2469_,
		_w2470_
	);
	LUT3 #(
		.INIT('hd0)
	) name1121 (
		_w2246_,
		_w2467_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('hb)
	) name1122 (
		_w2466_,
		_w2471_,
		_w2472_
	);
	LUT4 #(
		.INIT('h0002)
	) name1123 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2473_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1124 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2474_
	);
	LUT3 #(
		.INIT('h02)
	) name1125 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w2320_,
		_w2473_,
		_w2475_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1126 (
		_w2293_,
		_w2294_,
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2451_,
		_w2477_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1128 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2451_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		_w2476_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('hc055)
	) name1130 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2473_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name1131 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w2288_,
		_w2481_
	);
	LUT3 #(
		.INIT('h80)
	) name1132 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2322_,
		_w2482_
	);
	LUT4 #(
		.INIT('h010f)
	) name1133 (
		_w2303_,
		_w2304_,
		_w2481_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('hd0)
	) name1134 (
		_w2246_,
		_w2480_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('hb)
	) name1135 (
		_w2479_,
		_w2484_,
		_w2485_
	);
	LUT3 #(
		.INIT('he0)
	) name1136 (
		_w2261_,
		_w2262_,
		_w2317_,
		_w2486_
	);
	LUT3 #(
		.INIT('he0)
	) name1137 (
		_w2265_,
		_w2266_,
		_w2322_,
		_w2487_
	);
	LUT3 #(
		.INIT('ha8)
	) name1138 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2486_,
		_w2487_,
		_w2488_
	);
	LUT3 #(
		.INIT('h02)
	) name1139 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w2320_,
		_w2473_,
		_w2489_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1140 (
		_w2274_,
		_w2275_,
		_w2474_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w2477_,
		_w2490_,
		_w2491_
	);
	LUT3 #(
		.INIT('ha8)
	) name1142 (
		_w1679_,
		_w2488_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h2)
	) name1143 (
		_w2283_,
		_w2490_,
		_w2493_
	);
	LUT4 #(
		.INIT('hc055)
	) name1144 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2473_,
		_w2494_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w2288_,
		_w2495_
	);
	LUT3 #(
		.INIT('h0d)
	) name1146 (
		_w2246_,
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w2493_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('hb)
	) name1148 (
		_w2492_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('he0)
	) name1149 (
		_w2265_,
		_w2266_,
		_w2320_,
		_w2499_
	);
	LUT3 #(
		.INIT('he0)
	) name1150 (
		_w2261_,
		_w2262_,
		_w2322_,
		_w2500_
	);
	LUT3 #(
		.INIT('ha8)
	) name1151 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h0004)
	) name1152 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2502_
	);
	LUT4 #(
		.INIT('hfff9)
	) name1153 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2503_
	);
	LUT3 #(
		.INIT('h02)
	) name1154 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w2473_,
		_w2502_,
		_w2504_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1155 (
		_w2274_,
		_w2275_,
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2323_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT3 #(
		.INIT('ha8)
	) name1158 (
		_w1679_,
		_w2501_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w2283_,
		_w2505_,
		_w2509_
	);
	LUT4 #(
		.INIT('hc055)
	) name1160 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2502_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w2288_,
		_w2511_
	);
	LUT3 #(
		.INIT('h0d)
	) name1162 (
		_w2246_,
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w2509_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('hb)
	) name1164 (
		_w2508_,
		_w2513_,
		_w2514_
	);
	LUT3 #(
		.INIT('h02)
	) name1165 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w2473_,
		_w2502_,
		_w2515_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1166 (
		_w2293_,
		_w2294_,
		_w2503_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1167 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2323_,
		_w2517_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('hc055)
	) name1169 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2502_,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name1170 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w2288_,
		_w2520_
	);
	LUT3 #(
		.INIT('h80)
	) name1171 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2320_,
		_w2521_
	);
	LUT4 #(
		.INIT('h010f)
	) name1172 (
		_w2303_,
		_w2304_,
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT3 #(
		.INIT('hd0)
	) name1173 (
		_w2246_,
		_w2519_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('hb)
	) name1174 (
		_w2518_,
		_w2523_,
		_w2524_
	);
	LUT3 #(
		.INIT('he0)
	) name1175 (
		_w2261_,
		_w2262_,
		_w2320_,
		_w2525_
	);
	LUT3 #(
		.INIT('he0)
	) name1176 (
		_w2265_,
		_w2266_,
		_w2473_,
		_w2526_
	);
	LUT3 #(
		.INIT('ha8)
	) name1177 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h0008)
	) name1178 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2528_
	);
	LUT4 #(
		.INIT('hfff3)
	) name1179 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2529_
	);
	LUT3 #(
		.INIT('h02)
	) name1180 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w2502_,
		_w2528_,
		_w2530_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1181 (
		_w2274_,
		_w2275_,
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2474_,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('ha8)
	) name1184 (
		_w1679_,
		_w2527_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		_w2283_,
		_w2531_,
		_w2535_
	);
	LUT4 #(
		.INIT('hc055)
	) name1186 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2528_,
		_w2536_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w2288_,
		_w2537_
	);
	LUT3 #(
		.INIT('h0d)
	) name1188 (
		_w2246_,
		_w2536_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h4)
	) name1189 (
		_w2535_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('hb)
	) name1190 (
		_w2534_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h02)
	) name1191 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w2502_,
		_w2528_,
		_w2541_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1192 (
		_w2293_,
		_w2294_,
		_w2529_,
		_w2541_,
		_w2542_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1193 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2474_,
		_w2543_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT4 #(
		.INIT('hc055)
	) name1195 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2528_,
		_w2545_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w2288_,
		_w2546_
	);
	LUT3 #(
		.INIT('h80)
	) name1197 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2473_,
		_w2547_
	);
	LUT4 #(
		.INIT('h010f)
	) name1198 (
		_w2303_,
		_w2304_,
		_w2546_,
		_w2547_,
		_w2548_
	);
	LUT3 #(
		.INIT('hd0)
	) name1199 (
		_w2246_,
		_w2545_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('hb)
	) name1200 (
		_w2544_,
		_w2549_,
		_w2550_
	);
	LUT3 #(
		.INIT('he0)
	) name1201 (
		_w2261_,
		_w2262_,
		_w2473_,
		_w2551_
	);
	LUT3 #(
		.INIT('he0)
	) name1202 (
		_w2265_,
		_w2266_,
		_w2502_,
		_w2552_
	);
	LUT3 #(
		.INIT('ha8)
	) name1203 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2551_,
		_w2552_,
		_w2553_
	);
	LUT4 #(
		.INIT('h0010)
	) name1204 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2554_
	);
	LUT4 #(
		.INIT('hffe7)
	) name1205 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2555_
	);
	LUT3 #(
		.INIT('h02)
	) name1206 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w2528_,
		_w2554_,
		_w2556_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1207 (
		_w2274_,
		_w2275_,
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name1208 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2503_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT3 #(
		.INIT('ha8)
	) name1210 (
		_w1679_,
		_w2553_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name1211 (
		_w2283_,
		_w2557_,
		_w2561_
	);
	LUT4 #(
		.INIT('hc055)
	) name1212 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2554_,
		_w2562_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w2288_,
		_w2563_
	);
	LUT3 #(
		.INIT('h0d)
	) name1214 (
		_w2246_,
		_w2562_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h4)
	) name1215 (
		_w2561_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('hb)
	) name1216 (
		_w2560_,
		_w2565_,
		_w2566_
	);
	LUT3 #(
		.INIT('h02)
	) name1217 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w2528_,
		_w2554_,
		_w2567_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1218 (
		_w2293_,
		_w2294_,
		_w2555_,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1219 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2503_,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		_w2568_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('hc055)
	) name1221 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2554_,
		_w2571_
	);
	LUT2 #(
		.INIT('h2)
	) name1222 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w2288_,
		_w2572_
	);
	LUT3 #(
		.INIT('h80)
	) name1223 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2502_,
		_w2573_
	);
	LUT4 #(
		.INIT('h010f)
	) name1224 (
		_w2303_,
		_w2304_,
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('hd0)
	) name1225 (
		_w2246_,
		_w2571_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('hb)
	) name1226 (
		_w2570_,
		_w2575_,
		_w2576_
	);
	LUT3 #(
		.INIT('he0)
	) name1227 (
		_w2261_,
		_w2262_,
		_w2502_,
		_w2577_
	);
	LUT3 #(
		.INIT('he0)
	) name1228 (
		_w2265_,
		_w2266_,
		_w2528_,
		_w2578_
	);
	LUT3 #(
		.INIT('ha8)
	) name1229 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT4 #(
		.INIT('h0020)
	) name1230 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2580_
	);
	LUT4 #(
		.INIT('hffcf)
	) name1231 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2581_
	);
	LUT3 #(
		.INIT('h02)
	) name1232 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w2554_,
		_w2580_,
		_w2582_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1233 (
		_w2274_,
		_w2275_,
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2529_,
		_w2584_
	);
	LUT2 #(
		.INIT('h1)
	) name1235 (
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT3 #(
		.INIT('ha8)
	) name1236 (
		_w1679_,
		_w2579_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		_w2283_,
		_w2583_,
		_w2587_
	);
	LUT4 #(
		.INIT('hc055)
	) name1238 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2580_,
		_w2588_
	);
	LUT2 #(
		.INIT('h2)
	) name1239 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w2288_,
		_w2589_
	);
	LUT3 #(
		.INIT('h0d)
	) name1240 (
		_w2246_,
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		_w2587_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('hb)
	) name1242 (
		_w2586_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('h02)
	) name1243 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w2554_,
		_w2580_,
		_w2593_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1244 (
		_w2293_,
		_w2294_,
		_w2581_,
		_w2593_,
		_w2594_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1245 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2529_,
		_w2595_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT4 #(
		.INIT('hc055)
	) name1247 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2580_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name1248 (
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w2288_,
		_w2598_
	);
	LUT3 #(
		.INIT('h80)
	) name1249 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2528_,
		_w2599_
	);
	LUT4 #(
		.INIT('h010f)
	) name1250 (
		_w2303_,
		_w2304_,
		_w2598_,
		_w2599_,
		_w2600_
	);
	LUT3 #(
		.INIT('hd0)
	) name1251 (
		_w2246_,
		_w2597_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('hb)
	) name1252 (
		_w2596_,
		_w2601_,
		_w2602_
	);
	LUT3 #(
		.INIT('he0)
	) name1253 (
		_w2261_,
		_w2262_,
		_w2528_,
		_w2603_
	);
	LUT3 #(
		.INIT('he0)
	) name1254 (
		_w2265_,
		_w2266_,
		_w2554_,
		_w2604_
	);
	LUT3 #(
		.INIT('ha8)
	) name1255 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2603_,
		_w2604_,
		_w2605_
	);
	LUT4 #(
		.INIT('h0040)
	) name1256 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2606_
	);
	LUT4 #(
		.INIT('hff9f)
	) name1257 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2607_
	);
	LUT3 #(
		.INIT('h02)
	) name1258 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w2580_,
		_w2606_,
		_w2608_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1259 (
		_w2274_,
		_w2275_,
		_w2607_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h2)
	) name1260 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2555_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name1261 (
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT3 #(
		.INIT('ha8)
	) name1262 (
		_w1679_,
		_w2605_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h2)
	) name1263 (
		_w2283_,
		_w2609_,
		_w2613_
	);
	LUT4 #(
		.INIT('hc055)
	) name1264 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2606_,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w2288_,
		_w2615_
	);
	LUT3 #(
		.INIT('h0d)
	) name1266 (
		_w2246_,
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w2613_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('hb)
	) name1268 (
		_w2612_,
		_w2617_,
		_w2618_
	);
	LUT3 #(
		.INIT('h02)
	) name1269 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w2580_,
		_w2606_,
		_w2619_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1270 (
		_w2293_,
		_w2294_,
		_w2607_,
		_w2619_,
		_w2620_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1271 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2555_,
		_w2621_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT4 #(
		.INIT('hc055)
	) name1273 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2606_,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name1274 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w2288_,
		_w2624_
	);
	LUT3 #(
		.INIT('h80)
	) name1275 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2554_,
		_w2625_
	);
	LUT4 #(
		.INIT('h010f)
	) name1276 (
		_w2303_,
		_w2304_,
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT3 #(
		.INIT('hd0)
	) name1277 (
		_w2246_,
		_w2623_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('hb)
	) name1278 (
		_w2622_,
		_w2627_,
		_w2628_
	);
	LUT3 #(
		.INIT('he0)
	) name1279 (
		_w2261_,
		_w2262_,
		_w2554_,
		_w2629_
	);
	LUT3 #(
		.INIT('he0)
	) name1280 (
		_w2265_,
		_w2266_,
		_w2580_,
		_w2630_
	);
	LUT3 #(
		.INIT('ha8)
	) name1281 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('hff3f)
	) name1282 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2632_
	);
	LUT3 #(
		.INIT('h02)
	) name1283 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w2349_,
		_w2606_,
		_w2633_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1284 (
		_w2274_,
		_w2275_,
		_w2632_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2581_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w2634_,
		_w2635_,
		_w2636_
	);
	LUT3 #(
		.INIT('ha8)
	) name1287 (
		_w1679_,
		_w2631_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w2283_,
		_w2634_,
		_w2638_
	);
	LUT4 #(
		.INIT('hc055)
	) name1289 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2349_,
		_w2639_
	);
	LUT2 #(
		.INIT('h2)
	) name1290 (
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w2288_,
		_w2640_
	);
	LUT3 #(
		.INIT('h0d)
	) name1291 (
		_w2246_,
		_w2639_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name1292 (
		_w2638_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('hb)
	) name1293 (
		_w2637_,
		_w2642_,
		_w2643_
	);
	LUT3 #(
		.INIT('h02)
	) name1294 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w2349_,
		_w2606_,
		_w2644_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1295 (
		_w2293_,
		_w2294_,
		_w2632_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1296 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2581_,
		_w2646_
	);
	LUT2 #(
		.INIT('h4)
	) name1297 (
		_w2645_,
		_w2646_,
		_w2647_
	);
	LUT4 #(
		.INIT('hc055)
	) name1298 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2349_,
		_w2648_
	);
	LUT2 #(
		.INIT('h2)
	) name1299 (
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w2288_,
		_w2649_
	);
	LUT3 #(
		.INIT('h80)
	) name1300 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2580_,
		_w2650_
	);
	LUT4 #(
		.INIT('h010f)
	) name1301 (
		_w2303_,
		_w2304_,
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT3 #(
		.INIT('hd0)
	) name1302 (
		_w2246_,
		_w2648_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('hb)
	) name1303 (
		_w2647_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('he0)
	) name1304 (
		_w2261_,
		_w2262_,
		_w2580_,
		_w2654_
	);
	LUT3 #(
		.INIT('he0)
	) name1305 (
		_w2265_,
		_w2266_,
		_w2606_,
		_w2655_
	);
	LUT3 #(
		.INIT('ha8)
	) name1306 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT3 #(
		.INIT('h02)
	) name1307 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w2250_,
		_w2349_,
		_w2657_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1308 (
		_w2274_,
		_w2275_,
		_w2350_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2607_,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT3 #(
		.INIT('ha8)
	) name1311 (
		_w1679_,
		_w2656_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		_w2283_,
		_w2658_,
		_w2662_
	);
	LUT4 #(
		.INIT('hc055)
	) name1313 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2250_,
		_w2663_
	);
	LUT2 #(
		.INIT('h2)
	) name1314 (
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w2288_,
		_w2664_
	);
	LUT3 #(
		.INIT('h0d)
	) name1315 (
		_w2246_,
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w2662_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('hb)
	) name1317 (
		_w2661_,
		_w2666_,
		_w2667_
	);
	LUT3 #(
		.INIT('h02)
	) name1318 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w2250_,
		_w2349_,
		_w2668_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1319 (
		_w2293_,
		_w2294_,
		_w2350_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1320 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2607_,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w2669_,
		_w2670_,
		_w2671_
	);
	LUT4 #(
		.INIT('hc055)
	) name1322 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2250_,
		_w2672_
	);
	LUT2 #(
		.INIT('h2)
	) name1323 (
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w2288_,
		_w2673_
	);
	LUT3 #(
		.INIT('h80)
	) name1324 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2606_,
		_w2674_
	);
	LUT4 #(
		.INIT('h010f)
	) name1325 (
		_w2303_,
		_w2304_,
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT3 #(
		.INIT('hd0)
	) name1326 (
		_w2246_,
		_w2672_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('hb)
	) name1327 (
		_w2671_,
		_w2676_,
		_w2677_
	);
	LUT3 #(
		.INIT('he0)
	) name1328 (
		_w2261_,
		_w2262_,
		_w2606_,
		_w2678_
	);
	LUT3 #(
		.INIT('he0)
	) name1329 (
		_w2265_,
		_w2266_,
		_w2349_,
		_w2679_
	);
	LUT3 #(
		.INIT('ha8)
	) name1330 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h02)
	) name1331 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w2250_,
		_w2264_,
		_w2681_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1332 (
		_w2274_,
		_w2275_,
		_w2279_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h2)
	) name1333 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2632_,
		_w2683_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('ha8)
	) name1335 (
		_w1679_,
		_w2680_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		_w2283_,
		_w2682_,
		_w2686_
	);
	LUT4 #(
		.INIT('hc055)
	) name1337 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1531_,
		_w1536_,
		_w2264_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w2288_,
		_w2688_
	);
	LUT3 #(
		.INIT('h0d)
	) name1339 (
		_w2246_,
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		_w2686_,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('hb)
	) name1341 (
		_w2685_,
		_w2690_,
		_w2691_
	);
	LUT3 #(
		.INIT('h02)
	) name1342 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w2250_,
		_w2264_,
		_w2692_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1343 (
		_w2279_,
		_w2293_,
		_w2294_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1344 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w2632_,
		_w2694_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		_w2693_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('hc055)
	) name1346 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1519_,
		_w1524_,
		_w2264_,
		_w2696_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w2288_,
		_w2697_
	);
	LUT3 #(
		.INIT('h80)
	) name1348 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2349_,
		_w2698_
	);
	LUT4 #(
		.INIT('h010f)
	) name1349 (
		_w2303_,
		_w2304_,
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT3 #(
		.INIT('hd0)
	) name1350 (
		_w2246_,
		_w2696_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('hb)
	) name1351 (
		_w2695_,
		_w2700_,
		_w2701_
	);
	LUT3 #(
		.INIT('h02)
	) name1352 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2103_,
		_w2172_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2703_
	);
	LUT3 #(
		.INIT('h80)
	) name1354 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2704_
	);
	LUT4 #(
		.INIT('h8000)
	) name1355 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2705_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2706_
	);
	LUT3 #(
		.INIT('h80)
	) name1357 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2708_
	);
	LUT3 #(
		.INIT('h80)
	) name1359 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2710_
	);
	LUT3 #(
		.INIT('h80)
	) name1361 (
		_w2709_,
		_w2707_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h8000)
	) name1362 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2709_,
		_w2707_,
		_w2710_,
		_w2712_
	);
	LUT3 #(
		.INIT('h80)
	) name1363 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2713_
	);
	LUT4 #(
		.INIT('h8000)
	) name1364 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2714_
	);
	LUT4 #(
		.INIT('h8000)
	) name1365 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2716_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2717_
	);
	LUT3 #(
		.INIT('h80)
	) name1368 (
		_w2715_,
		_w2716_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h8)
	) name1369 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2719_
	);
	LUT4 #(
		.INIT('h8000)
	) name1370 (
		_w2715_,
		_w2716_,
		_w2717_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2721_
	);
	LUT3 #(
		.INIT('h80)
	) name1372 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2722_
	);
	LUT4 #(
		.INIT('h8000)
	) name1373 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2723_
	);
	LUT3 #(
		.INIT('h80)
	) name1374 (
		_w2712_,
		_w2720_,
		_w2723_,
		_w2724_
	);
	LUT4 #(
		.INIT('h8000)
	) name1375 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2723_,
		_w2725_
	);
	LUT4 #(
		.INIT('h8000)
	) name1376 (
		_w2712_,
		_w2720_,
		_w2723_,
		_w2705_,
		_w2726_
	);
	LUT4 #(
		.INIT('h9333)
	) name1377 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2724_,
		_w2705_,
		_w2727_
	);
	LUT2 #(
		.INIT('h6)
	) name1378 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2725_,
		_w2728_
	);
	LUT3 #(
		.INIT('h6c)
	) name1379 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2725_,
		_w2729_
	);
	LUT3 #(
		.INIT('h81)
	) name1380 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2725_,
		_w2730_
	);
	LUT3 #(
		.INIT('h6a)
	) name1381 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2703_,
		_w2725_,
		_w2731_
	);
	LUT4 #(
		.INIT('h8001)
	) name1382 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2725_,
		_w2732_
	);
	LUT2 #(
		.INIT('h8)
	) name1383 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2733_
	);
	LUT3 #(
		.INIT('h80)
	) name1384 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2734_
	);
	LUT4 #(
		.INIT('h8000)
	) name1385 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2735_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2735_,
		_w2736_
	);
	LUT3 #(
		.INIT('h80)
	) name1387 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2715_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h8000)
	) name1388 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2711_,
		_w2715_,
		_w2736_,
		_w2738_
	);
	LUT4 #(
		.INIT('h8000)
	) name1389 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2738_,
		_w2722_,
		_w2739_
	);
	LUT3 #(
		.INIT('h80)
	) name1390 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2705_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h8000)
	) name1391 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2738_,
		_w2722_,
		_w2741_
	);
	LUT4 #(
		.INIT('h1333)
	) name1392 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2741_,
		_w2704_,
		_w2742_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w2740_,
		_w2742_,
		_w2743_
	);
	LUT3 #(
		.INIT('ha8)
	) name1394 (
		_w2732_,
		_w2740_,
		_w2742_,
		_w2744_
	);
	LUT4 #(
		.INIT('h153f)
	) name1395 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1966_,
		_w1970_,
		_w2745_
	);
	LUT4 #(
		.INIT('h135f)
	) name1396 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1957_,
		_w1946_,
		_w2746_
	);
	LUT4 #(
		.INIT('h153f)
	) name1397 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1954_,
		_w1960_,
		_w2747_
	);
	LUT4 #(
		.INIT('h153f)
	) name1398 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1952_,
		_w1969_,
		_w2748_
	);
	LUT4 #(
		.INIT('h8000)
	) name1399 (
		_w2747_,
		_w2748_,
		_w2745_,
		_w2746_,
		_w2749_
	);
	LUT4 #(
		.INIT('h153f)
	) name1400 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1949_,
		_w1967_,
		_w2750_
	);
	LUT4 #(
		.INIT('h135f)
	) name1401 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1947_,
		_w1964_,
		_w2751_
	);
	LUT4 #(
		.INIT('h135f)
	) name1402 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1956_,
		_w1950_,
		_w2752_
	);
	LUT4 #(
		.INIT('h153f)
	) name1403 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w1961_,
		_w1963_,
		_w2753_
	);
	LUT4 #(
		.INIT('h8000)
	) name1404 (
		_w2752_,
		_w2753_,
		_w2750_,
		_w2751_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name1405 (
		_w2749_,
		_w2754_,
		_w2755_
	);
	LUT4 #(
		.INIT('h8000)
	) name1406 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2714_,
		_w2756_
	);
	LUT2 #(
		.INIT('h6)
	) name1407 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2756_,
		_w2757_
	);
	LUT3 #(
		.INIT('h08)
	) name1408 (
		_w2749_,
		_w2754_,
		_w2757_,
		_w2758_
	);
	LUT4 #(
		.INIT('h153f)
	) name1409 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1954_,
		_w1956_,
		_w2759_
	);
	LUT4 #(
		.INIT('h153f)
	) name1410 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1946_,
		_w1963_,
		_w2760_
	);
	LUT4 #(
		.INIT('h135f)
	) name1411 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w1966_,
		_w1961_,
		_w2761_
	);
	LUT4 #(
		.INIT('h135f)
	) name1412 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1957_,
		_w1950_,
		_w2762_
	);
	LUT4 #(
		.INIT('h8000)
	) name1413 (
		_w2761_,
		_w2762_,
		_w2759_,
		_w2760_,
		_w2763_
	);
	LUT4 #(
		.INIT('h153f)
	) name1414 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1949_,
		_w1969_,
		_w2764_
	);
	LUT4 #(
		.INIT('h135f)
	) name1415 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1960_,
		_w1964_,
		_w2765_
	);
	LUT4 #(
		.INIT('h135f)
	) name1416 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w1947_,
		_w1967_,
		_w2766_
	);
	LUT4 #(
		.INIT('h153f)
	) name1417 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1952_,
		_w1970_,
		_w2767_
	);
	LUT4 #(
		.INIT('h8000)
	) name1418 (
		_w2766_,
		_w2767_,
		_w2764_,
		_w2765_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		_w2763_,
		_w2768_,
		_w2769_
	);
	LUT3 #(
		.INIT('h07)
	) name1420 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2770_
	);
	LUT3 #(
		.INIT('h78)
	) name1421 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2771_
	);
	LUT3 #(
		.INIT('h70)
	) name1422 (
		_w2763_,
		_w2768_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h153f)
	) name1423 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1957_,
		_w1963_,
		_w2773_
	);
	LUT4 #(
		.INIT('h153f)
	) name1424 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1954_,
		_w1960_,
		_w2774_
	);
	LUT4 #(
		.INIT('h153f)
	) name1425 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1949_,
		_w1964_,
		_w2775_
	);
	LUT4 #(
		.INIT('h135f)
	) name1426 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1952_,
		_w1950_,
		_w2776_
	);
	LUT4 #(
		.INIT('h8000)
	) name1427 (
		_w2775_,
		_w2776_,
		_w2773_,
		_w2774_,
		_w2777_
	);
	LUT4 #(
		.INIT('h153f)
	) name1428 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w1946_,
		_w1970_,
		_w2778_
	);
	LUT4 #(
		.INIT('h135f)
	) name1429 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w1956_,
		_w1969_,
		_w2779_
	);
	LUT4 #(
		.INIT('h135f)
	) name1430 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1947_,
		_w1967_,
		_w2780_
	);
	LUT4 #(
		.INIT('h135f)
	) name1431 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1966_,
		_w1961_,
		_w2781_
	);
	LUT4 #(
		.INIT('h8000)
	) name1432 (
		_w2780_,
		_w2781_,
		_w2778_,
		_w2779_,
		_w2782_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		_w2777_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h135f)
	) name1434 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1952_,
		_w1949_,
		_w2784_
	);
	LUT4 #(
		.INIT('h153f)
	) name1435 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w1969_,
		_w1970_,
		_w2785_
	);
	LUT4 #(
		.INIT('h153f)
	) name1436 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1954_,
		_w1966_,
		_w2786_
	);
	LUT4 #(
		.INIT('h135f)
	) name1437 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1957_,
		_w1946_,
		_w2787_
	);
	LUT4 #(
		.INIT('h8000)
	) name1438 (
		_w2786_,
		_w2787_,
		_w2784_,
		_w2785_,
		_w2788_
	);
	LUT4 #(
		.INIT('h135f)
	) name1439 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w1956_,
		_w1947_,
		_w2789_
	);
	LUT4 #(
		.INIT('h153f)
	) name1440 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1950_,
		_w1964_,
		_w2790_
	);
	LUT4 #(
		.INIT('h153f)
	) name1441 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w1967_,
		_w1960_,
		_w2791_
	);
	LUT4 #(
		.INIT('h153f)
	) name1442 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w1961_,
		_w1963_,
		_w2792_
	);
	LUT4 #(
		.INIT('h8000)
	) name1443 (
		_w2791_,
		_w2792_,
		_w2789_,
		_w2790_,
		_w2793_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		_w2788_,
		_w2793_,
		_w2794_
	);
	LUT3 #(
		.INIT('h2a)
	) name1445 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2788_,
		_w2793_,
		_w2795_
	);
	LUT3 #(
		.INIT('h8e)
	) name1446 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2783_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('hb890)
	) name1447 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2783_,
		_w2794_,
		_w2797_
	);
	LUT3 #(
		.INIT('h08)
	) name1448 (
		_w2763_,
		_w2768_,
		_w2771_,
		_w2798_
	);
	LUT4 #(
		.INIT('h135f)
	) name1449 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w1956_,
		_w1947_,
		_w2799_
	);
	LUT4 #(
		.INIT('h153f)
	) name1450 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w1969_,
		_w1960_,
		_w2800_
	);
	LUT4 #(
		.INIT('h153f)
	) name1451 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1946_,
		_w1961_,
		_w2801_
	);
	LUT4 #(
		.INIT('h135f)
	) name1452 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1963_,
		_w1964_,
		_w2802_
	);
	LUT4 #(
		.INIT('h8000)
	) name1453 (
		_w2801_,
		_w2802_,
		_w2799_,
		_w2800_,
		_w2803_
	);
	LUT4 #(
		.INIT('h135f)
	) name1454 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1954_,
		_w1950_,
		_w2804_
	);
	LUT4 #(
		.INIT('h153f)
	) name1455 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1949_,
		_w1966_,
		_w2805_
	);
	LUT4 #(
		.INIT('h135f)
	) name1456 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1952_,
		_w1967_,
		_w2806_
	);
	LUT4 #(
		.INIT('h153f)
	) name1457 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1957_,
		_w1970_,
		_w2807_
	);
	LUT4 #(
		.INIT('h8000)
	) name1458 (
		_w2806_,
		_w2807_,
		_w2804_,
		_w2805_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		_w2803_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('h8000)
	) name1460 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2810_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1461 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2811_
	);
	LUT3 #(
		.INIT('h08)
	) name1462 (
		_w2803_,
		_w2808_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h1)
	) name1463 (
		_w2798_,
		_w2812_,
		_w2813_
	);
	LUT4 #(
		.INIT('h135f)
	) name1464 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1956_,
		_w1964_,
		_w2814_
	);
	LUT4 #(
		.INIT('h135f)
	) name1465 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1952_,
		_w1950_,
		_w2815_
	);
	LUT4 #(
		.INIT('h153f)
	) name1466 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w1947_,
		_w1963_,
		_w2816_
	);
	LUT4 #(
		.INIT('h153f)
	) name1467 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1949_,
		_w1961_,
		_w2817_
	);
	LUT4 #(
		.INIT('h8000)
	) name1468 (
		_w2816_,
		_w2817_,
		_w2814_,
		_w2815_,
		_w2818_
	);
	LUT4 #(
		.INIT('h135f)
	) name1469 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1957_,
		_w1946_,
		_w2819_
	);
	LUT4 #(
		.INIT('h153f)
	) name1470 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1954_,
		_w1967_,
		_w2820_
	);
	LUT4 #(
		.INIT('h135f)
	) name1471 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w1970_,
		_w1960_,
		_w2821_
	);
	LUT4 #(
		.INIT('h135f)
	) name1472 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w1966_,
		_w1969_,
		_w2822_
	);
	LUT4 #(
		.INIT('h8000)
	) name1473 (
		_w2821_,
		_w2822_,
		_w2819_,
		_w2820_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		_w2818_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name1475 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2713_,
		_w2810_,
		_w2825_
	);
	LUT3 #(
		.INIT('h08)
	) name1476 (
		_w2818_,
		_w2823_,
		_w2825_,
		_w2826_
	);
	LUT3 #(
		.INIT('h01)
	) name1477 (
		_w2798_,
		_w2812_,
		_w2826_,
		_w2827_
	);
	LUT3 #(
		.INIT('h70)
	) name1478 (
		_w2818_,
		_w2823_,
		_w2825_,
		_w2828_
	);
	LUT3 #(
		.INIT('h70)
	) name1479 (
		_w2803_,
		_w2808_,
		_w2811_,
		_w2829_
	);
	LUT3 #(
		.INIT('h54)
	) name1480 (
		_w2826_,
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('h004f)
	) name1481 (
		_w2772_,
		_w2797_,
		_w2827_,
		_w2830_,
		_w2831_
	);
	LUT4 #(
		.INIT('h153f)
	) name1482 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1949_,
		_w1967_,
		_w2832_
	);
	LUT4 #(
		.INIT('h135f)
	) name1483 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w1956_,
		_w1960_,
		_w2833_
	);
	LUT4 #(
		.INIT('h135f)
	) name1484 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1952_,
		_w1950_,
		_w2834_
	);
	LUT4 #(
		.INIT('h153f)
	) name1485 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1957_,
		_w1961_,
		_w2835_
	);
	LUT4 #(
		.INIT('h8000)
	) name1486 (
		_w2834_,
		_w2835_,
		_w2832_,
		_w2833_,
		_w2836_
	);
	LUT4 #(
		.INIT('h153f)
	) name1487 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1946_,
		_w1970_,
		_w2837_
	);
	LUT4 #(
		.INIT('h153f)
	) name1488 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1966_,
		_w1963_,
		_w2838_
	);
	LUT4 #(
		.INIT('h153f)
	) name1489 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1954_,
		_w1969_,
		_w2839_
	);
	LUT4 #(
		.INIT('h135f)
	) name1490 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1947_,
		_w1964_,
		_w2840_
	);
	LUT4 #(
		.INIT('h8000)
	) name1491 (
		_w2839_,
		_w2840_,
		_w2837_,
		_w2838_,
		_w2841_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		_w2836_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1493 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2714_,
		_w2843_
	);
	LUT3 #(
		.INIT('h08)
	) name1494 (
		_w2836_,
		_w2841_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('h135f)
	) name1495 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1967_,
		_w1964_,
		_w2845_
	);
	LUT4 #(
		.INIT('h135f)
	) name1496 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w1956_,
		_w1960_,
		_w2846_
	);
	LUT4 #(
		.INIT('h135f)
	) name1497 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w1952_,
		_w1957_,
		_w2847_
	);
	LUT4 #(
		.INIT('h153f)
	) name1498 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w1969_,
		_w1961_,
		_w2848_
	);
	LUT4 #(
		.INIT('h8000)
	) name1499 (
		_w2847_,
		_w2848_,
		_w2845_,
		_w2846_,
		_w2849_
	);
	LUT4 #(
		.INIT('h153f)
	) name1500 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1946_,
		_w1970_,
		_w2850_
	);
	LUT4 #(
		.INIT('h135f)
	) name1501 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1947_,
		_w1966_,
		_w2851_
	);
	LUT4 #(
		.INIT('h153f)
	) name1502 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1954_,
		_w1963_,
		_w2852_
	);
	LUT4 #(
		.INIT('h135f)
	) name1503 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1949_,
		_w1950_,
		_w2853_
	);
	LUT4 #(
		.INIT('h8000)
	) name1504 (
		_w2852_,
		_w2853_,
		_w2850_,
		_w2851_,
		_w2854_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w2849_,
		_w2854_,
		_w2855_
	);
	LUT3 #(
		.INIT('h6c)
	) name1506 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w2714_,
		_w2856_
	);
	LUT3 #(
		.INIT('h08)
	) name1507 (
		_w2849_,
		_w2854_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w2844_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w2758_,
		_w2844_,
		_w2859_
	);
	LUT3 #(
		.INIT('h70)
	) name1510 (
		_w2836_,
		_w2841_,
		_w2843_,
		_w2860_
	);
	LUT3 #(
		.INIT('h70)
	) name1511 (
		_w2849_,
		_w2854_,
		_w2856_,
		_w2861_
	);
	LUT4 #(
		.INIT('h3110)
	) name1512 (
		_w2842_,
		_w2758_,
		_w2843_,
		_w2861_,
		_w2862_
	);
	LUT3 #(
		.INIT('h70)
	) name1513 (
		_w2749_,
		_w2754_,
		_w2757_,
		_w2863_
	);
	LUT3 #(
		.INIT('h6c)
	) name1514 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2756_,
		_w2864_
	);
	LUT4 #(
		.INIT('h008f)
	) name1515 (
		_w2749_,
		_w2754_,
		_w2757_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h4)
	) name1516 (
		_w2862_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h8000)
	) name1517 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2867_
	);
	LUT3 #(
		.INIT('h80)
	) name1518 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2868_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1519 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2869_
	);
	LUT4 #(
		.INIT('h070f)
	) name1520 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2756_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w2868_,
		_w2870_,
		_w2871_
	);
	LUT3 #(
		.INIT('h32)
	) name1522 (
		_w2868_,
		_w2869_,
		_w2870_,
		_w2872_
	);
	LUT3 #(
		.INIT('h40)
	) name1523 (
		_w2862_,
		_w2865_,
		_w2872_,
		_w2873_
	);
	LUT4 #(
		.INIT('hef00)
	) name1524 (
		_w2758_,
		_w2831_,
		_w2858_,
		_w2873_,
		_w2874_
	);
	LUT4 #(
		.INIT('h8000)
	) name1525 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2717_,
		_w2875_
	);
	LUT3 #(
		.INIT('h0e)
	) name1526 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2867_,
		_w2875_,
		_w2876_
	);
	LUT4 #(
		.INIT('h8000)
	) name1527 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2735_,
		_w2756_,
		_w2877_
	);
	LUT3 #(
		.INIT('h0e)
	) name1528 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w2876_,
		_w2878_,
		_w2879_
	);
	LUT4 #(
		.INIT('h8000)
	) name1530 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2715_,
		_w2736_,
		_w2880_
	);
	LUT3 #(
		.INIT('h6c)
	) name1531 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2737_,
		_w2881_
	);
	LUT4 #(
		.INIT('h8000)
	) name1532 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2717_,
		_w2882_
	);
	LUT4 #(
		.INIT('h4e4c)
	) name1533 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2737_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h0001)
	) name1534 (
		_w2876_,
		_w2878_,
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2885_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1536 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2885_,
		_w2875_,
		_w2886_
	);
	LUT4 #(
		.INIT('h1555)
	) name1537 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2706_,
		_w2885_,
		_w2875_,
		_w2887_
	);
	LUT3 #(
		.INIT('h80)
	) name1538 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2707_,
		_w2880_,
		_w2888_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w2887_,
		_w2888_,
		_w2889_
	);
	LUT3 #(
		.INIT('h54)
	) name1540 (
		_w2886_,
		_w2887_,
		_w2888_,
		_w2890_
	);
	LUT3 #(
		.INIT('h6a)
	) name1541 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2885_,
		_w2875_,
		_w2891_
	);
	LUT4 #(
		.INIT('h0054)
	) name1542 (
		_w2886_,
		_w2887_,
		_w2888_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('h8000)
	) name1543 (
		_w2715_,
		_w2716_,
		_w2717_,
		_w2885_,
		_w2893_
	);
	LUT2 #(
		.INIT('h8)
	) name1544 (
		_w2707_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h8000)
	) name1545 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2707_,
		_w2893_,
		_w2895_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1546 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2707_,
		_w2893_,
		_w2896_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		_w2892_,
		_w2896_,
		_w2897_
	);
	LUT3 #(
		.INIT('h80)
	) name1548 (
		_w2708_,
		_w2707_,
		_w2893_,
		_w2898_
	);
	LUT4 #(
		.INIT('h8000)
	) name1549 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2708_,
		_w2707_,
		_w2893_,
		_w2899_
	);
	LUT2 #(
		.INIT('h6)
	) name1550 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2899_,
		_w2900_
	);
	LUT3 #(
		.INIT('h6c)
	) name1551 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2899_,
		_w2901_
	);
	LUT3 #(
		.INIT('h81)
	) name1552 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2899_,
		_w2902_
	);
	LUT4 #(
		.INIT('h8000)
	) name1553 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2903_
	);
	LUT4 #(
		.INIT('h8000)
	) name1554 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2721_,
		_w2712_,
		_w2720_,
		_w2904_
	);
	LUT3 #(
		.INIT('h0e)
	) name1555 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1556 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2906_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1557 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2711_,
		_w2737_,
		_w2907_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		_w2906_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h9)
	) name1559 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2904_,
		_w2909_
	);
	LUT3 #(
		.INIT('h40)
	) name1560 (
		_w2905_,
		_w2908_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h6)
	) name1561 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2739_,
		_w2911_
	);
	LUT4 #(
		.INIT('h0040)
	) name1562 (
		_w2905_,
		_w2908_,
		_w2909_,
		_w2911_,
		_w2912_
	);
	LUT3 #(
		.INIT('h0e)
	) name1563 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2895_,
		_w2899_,
		_w2913_
	);
	LUT3 #(
		.INIT('h08)
	) name1564 (
		_w2902_,
		_w2912_,
		_w2913_,
		_w2914_
	);
	LUT4 #(
		.INIT('h8000)
	) name1565 (
		_w2874_,
		_w2884_,
		_w2897_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('h1444)
	) name1566 (
		_w2755_,
		_w2727_,
		_w2744_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h6)
	) name1567 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w2917_
	);
	LUT3 #(
		.INIT('h70)
	) name1568 (
		_w2763_,
		_w2768_,
		_w2917_,
		_w2918_
	);
	LUT4 #(
		.INIT('h2032)
	) name1569 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2918_,
		_w2783_,
		_w2795_,
		_w2919_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1570 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2920_
	);
	LUT3 #(
		.INIT('h40)
	) name1571 (
		_w2920_,
		_w2818_,
		_w2823_,
		_w2921_
	);
	LUT3 #(
		.INIT('h78)
	) name1572 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2922_
	);
	LUT3 #(
		.INIT('h08)
	) name1573 (
		_w2803_,
		_w2808_,
		_w2922_,
		_w2923_
	);
	LUT3 #(
		.INIT('h08)
	) name1574 (
		_w2763_,
		_w2768_,
		_w2917_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w2923_,
		_w2924_,
		_w2925_
	);
	LUT3 #(
		.INIT('h01)
	) name1576 (
		_w2921_,
		_w2923_,
		_w2924_,
		_w2926_
	);
	LUT3 #(
		.INIT('h2a)
	) name1577 (
		_w2920_,
		_w2818_,
		_w2823_,
		_w2927_
	);
	LUT3 #(
		.INIT('h70)
	) name1578 (
		_w2803_,
		_w2808_,
		_w2922_,
		_w2928_
	);
	LUT3 #(
		.INIT('h23)
	) name1579 (
		_w2921_,
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h6)
	) name1580 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w2714_,
		_w2930_
	);
	LUT3 #(
		.INIT('h40)
	) name1581 (
		_w2930_,
		_w2849_,
		_w2854_,
		_w2931_
	);
	LUT3 #(
		.INIT('h6c)
	) name1582 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2714_,
		_w2932_
	);
	LUT3 #(
		.INIT('h40)
	) name1583 (
		_w2932_,
		_w2836_,
		_w2841_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w2931_,
		_w2933_,
		_w2934_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1585 (
		_w2919_,
		_w2926_,
		_w2929_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1586 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2714_,
		_w2936_
	);
	LUT3 #(
		.INIT('h70)
	) name1587 (
		_w2749_,
		_w2754_,
		_w2936_,
		_w2937_
	);
	LUT3 #(
		.INIT('h2a)
	) name1588 (
		_w2932_,
		_w2836_,
		_w2841_,
		_w2938_
	);
	LUT3 #(
		.INIT('h2a)
	) name1589 (
		_w2930_,
		_w2849_,
		_w2854_,
		_w2939_
	);
	LUT3 #(
		.INIT('h23)
	) name1590 (
		_w2933_,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h040d)
	) name1591 (
		_w2932_,
		_w2842_,
		_w2937_,
		_w2939_,
		_w2941_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1592 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2717_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h6)
	) name1594 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2715_,
		_w2944_
	);
	LUT3 #(
		.INIT('h48)
	) name1595 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2715_,
		_w2945_
	);
	LUT4 #(
		.INIT('h2080)
	) name1596 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2715_,
		_w2946_
	);
	LUT3 #(
		.INIT('h08)
	) name1597 (
		_w2749_,
		_w2754_,
		_w2936_,
		_w2947_
	);
	LUT4 #(
		.INIT('hf700)
	) name1598 (
		_w2749_,
		_w2754_,
		_w2936_,
		_w2946_,
		_w2948_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1599 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2715_,
		_w2736_,
		_w2949_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1600 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2715_,
		_w2716_,
		_w2950_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		_w2949_,
		_w2950_,
		_w2951_
	);
	LUT3 #(
		.INIT('h80)
	) name1602 (
		_w2943_,
		_w2948_,
		_w2951_,
		_w2952_
	);
	LUT3 #(
		.INIT('hb0)
	) name1603 (
		_w2935_,
		_w2941_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2893_,
		_w2954_
	);
	LUT3 #(
		.INIT('h6c)
	) name1605 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2893_,
		_w2955_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1606 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2893_,
		_w2956_
	);
	LUT2 #(
		.INIT('h6)
	) name1607 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2893_,
		_w2957_
	);
	LUT3 #(
		.INIT('h48)
	) name1608 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2893_,
		_w2958_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w2956_,
		_w2958_,
		_w2959_
	);
	LUT4 #(
		.INIT('hb000)
	) name1610 (
		_w2935_,
		_w2941_,
		_w2952_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h6)
	) name1611 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2738_,
		_w2961_
	);
	LUT4 #(
		.INIT('h8000)
	) name1612 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2707_,
		_w2893_,
		_w2962_
	);
	LUT2 #(
		.INIT('h6)
	) name1613 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2962_,
		_w2963_
	);
	LUT3 #(
		.INIT('h48)
	) name1614 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2961_,
		_w2962_,
		_w2964_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1615 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2708_,
		_w2707_,
		_w2893_,
		_w2965_
	);
	LUT4 #(
		.INIT('h4080)
	) name1616 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2961_,
		_w2898_,
		_w2966_
	);
	LUT4 #(
		.INIT('h9333)
	) name1617 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2707_,
		_w2893_,
		_w2967_
	);
	LUT2 #(
		.INIT('h2)
	) name1618 (
		_w2966_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1619 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2738_,
		_w2722_,
		_w2969_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1620 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2721_,
		_w2712_,
		_w2720_,
		_w2970_
	);
	LUT3 #(
		.INIT('h6a)
	) name1621 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2971_
	);
	LUT4 #(
		.INIT('h4888)
	) name1622 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2972_
	);
	LUT3 #(
		.INIT('h80)
	) name1623 (
		_w2969_,
		_w2970_,
		_w2972_,
		_w2973_
	);
	LUT3 #(
		.INIT('h80)
	) name1624 (
		_w2960_,
		_w2968_,
		_w2973_,
		_w2974_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1625 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2712_,
		_w2720_,
		_w2723_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2975_,
		_w2976_
	);
	LUT3 #(
		.INIT('h80)
	) name1627 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2975_,
		_w2977_
	);
	LUT3 #(
		.INIT('h95)
	) name1628 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2741_,
		_w2704_,
		_w2978_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT4 #(
		.INIT('h8000)
	) name1630 (
		_w2960_,
		_w2968_,
		_w2973_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h9)
	) name1631 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2726_,
		_w2981_
	);
	LUT4 #(
		.INIT('h5115)
	) name1632 (
		_w2173_,
		_w2755_,
		_w2980_,
		_w2981_,
		_w2982_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1633 (
		_w2171_,
		_w2702_,
		_w2916_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('hf800)
	) name1634 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2984_
	);
	LUT4 #(
		.INIT('h8000)
	) name1635 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h8000)
	) name1636 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2716_,
		_w2985_,
		_w2986_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1637 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2716_,
		_w2985_,
		_w2987_
	);
	LUT3 #(
		.INIT('h6c)
	) name1638 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2985_,
		_w2988_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1639 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2734_,
		_w2985_,
		_w2989_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		_w2987_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('h80)
	) name1641 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2987_,
		_w2989_,
		_w2991_
	);
	LUT2 #(
		.INIT('h6)
	) name1642 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2985_,
		_w2992_
	);
	LUT3 #(
		.INIT('h70)
	) name1643 (
		_w2749_,
		_w2754_,
		_w2992_,
		_w2993_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1644 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w2984_,
		_w2994_
	);
	LUT3 #(
		.INIT('h08)
	) name1645 (
		_w2836_,
		_w2841_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h6)
	) name1646 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2984_,
		_w2996_
	);
	LUT3 #(
		.INIT('h08)
	) name1647 (
		_w2818_,
		_w2823_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('h6c)
	) name1648 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w2984_,
		_w2998_
	);
	LUT3 #(
		.INIT('h08)
	) name1649 (
		_w2849_,
		_w2854_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		_w2997_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('h07)
	) name1651 (
		_w2763_,
		_w2768_,
		_w2771_,
		_w3001_
	);
	LUT2 #(
		.INIT('h9)
	) name1652 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w3002_
	);
	LUT3 #(
		.INIT('h07)
	) name1653 (
		_w2777_,
		_w2782_,
		_w3002_,
		_w3003_
	);
	LUT3 #(
		.INIT('h80)
	) name1654 (
		_w2777_,
		_w2782_,
		_w3002_,
		_w3004_
	);
	LUT3 #(
		.INIT('h15)
	) name1655 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2788_,
		_w2793_,
		_w3005_
	);
	LUT4 #(
		.INIT('h2032)
	) name1656 (
		_w2783_,
		_w3001_,
		_w3002_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('h80)
	) name1657 (
		_w2763_,
		_w2768_,
		_w2771_,
		_w3007_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1658 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w3008_
	);
	LUT3 #(
		.INIT('h08)
	) name1659 (
		_w2803_,
		_w2808_,
		_w3008_,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name1660 (
		_w3007_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('h70)
	) name1661 (
		_w2803_,
		_w2808_,
		_w3008_,
		_w3011_
	);
	LUT3 #(
		.INIT('h70)
	) name1662 (
		_w2818_,
		_w2823_,
		_w2996_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1664 (
		_w3000_,
		_w3006_,
		_w3010_,
		_w3013_,
		_w3014_
	);
	LUT3 #(
		.INIT('h70)
	) name1665 (
		_w2836_,
		_w2841_,
		_w2994_,
		_w3015_
	);
	LUT3 #(
		.INIT('h70)
	) name1666 (
		_w2849_,
		_w2854_,
		_w2998_,
		_w3016_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT3 #(
		.INIT('h45)
	) name1668 (
		_w2995_,
		_w3014_,
		_w3017_,
		_w3018_
	);
	LUT3 #(
		.INIT('h08)
	) name1669 (
		_w2749_,
		_w2754_,
		_w2992_,
		_w3019_
	);
	LUT4 #(
		.INIT('h0045)
	) name1670 (
		_w2995_,
		_w3014_,
		_w3017_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('h80)
	) name1671 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2733_,
		_w2986_,
		_w3021_
	);
	LUT4 #(
		.INIT('h8000)
	) name1672 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2733_,
		_w2986_,
		_w3022_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1673 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2733_,
		_w2986_,
		_w3023_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w2706_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('ha800)
	) name1675 (
		_w2991_,
		_w2993_,
		_w3020_,
		_w3024_,
		_w3025_
	);
	LUT3 #(
		.INIT('h80)
	) name1676 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2706_,
		_w3022_,
		_w3026_
	);
	LUT3 #(
		.INIT('h6a)
	) name1677 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2706_,
		_w3022_,
		_w3027_
	);
	LUT4 #(
		.INIT('h4888)
	) name1678 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2709_,
		_w2706_,
		_w3022_,
		_w3028_
	);
	LUT4 #(
		.INIT('h8000)
	) name1679 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2706_,
		_w3022_,
		_w3029_
	);
	LUT4 #(
		.INIT('h070f)
	) name1680 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h8000)
	) name1681 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2711_,
		_w2733_,
		_w2986_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w3030_,
		_w3031_,
		_w3032_
	);
	LUT4 #(
		.INIT('h8000)
	) name1683 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2733_,
		_w2712_,
		_w2986_,
		_w3033_
	);
	LUT3 #(
		.INIT('h6a)
	) name1684 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2711_,
		_w3021_,
		_w3034_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1685 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2721_,
		_w3031_,
		_w3033_,
		_w3035_
	);
	LUT3 #(
		.INIT('h10)
	) name1686 (
		_w3030_,
		_w3031_,
		_w3035_,
		_w3036_
	);
	LUT3 #(
		.INIT('h80)
	) name1687 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h8000)
	) name1688 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3033_,
		_w3038_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1689 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w3033_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3039_,
		_w3040_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1691 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2704_,
		_w3038_,
		_w3041_
	);
	LUT3 #(
		.INIT('h6c)
	) name1692 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w3038_,
		_w3042_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1693 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3038_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h8000)
	) name1695 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w3040_,
		_w3041_,
		_w3043_,
		_w3045_
	);
	LUT4 #(
		.INIT('h8000)
	) name1696 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1697 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2705_,
		_w3038_,
		_w3047_
	);
	LUT4 #(
		.INIT('he000)
	) name1698 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w2117_,
		_w2981_,
		_w3049_
	);
	LUT3 #(
		.INIT('h0b)
	) name1700 (
		_w2073_,
		_w2086_,
		_w2727_,
		_w3050_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1701 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w3051_
	);
	LUT4 #(
		.INIT('h0001)
	) name1702 (
		_w3050_,
		_w3051_,
		_w3049_,
		_w3048_,
		_w3052_
	);
	LUT4 #(
		.INIT('hd700)
	) name1703 (
		_w2181_,
		_w3046_,
		_w3047_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h0001)
	) name1704 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3054_
	);
	LUT4 #(
		.INIT('h0010)
	) name1705 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3055_
	);
	LUT4 #(
		.INIT('hfc21)
	) name1706 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w3056_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1707 (
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w3054_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1708 (
		_w1945_,
		_w2983_,
		_w3053_,
		_w3057_,
		_w3058_
	);
	LUT3 #(
		.INIT('h08)
	) name1709 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1842_,
		_w1915_,
		_w3059_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3060_
	);
	LUT3 #(
		.INIT('h80)
	) name1711 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3061_
	);
	LUT4 #(
		.INIT('h8000)
	) name1712 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w3062_
	);
	LUT3 #(
		.INIT('h80)
	) name1713 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3064_
	);
	LUT2 #(
		.INIT('h8)
	) name1715 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3065_
	);
	LUT3 #(
		.INIT('h80)
	) name1716 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		_w3064_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name1718 (
		_w3063_,
		_w3067_,
		_w3068_
	);
	LUT3 #(
		.INIT('h80)
	) name1719 (
		_w3060_,
		_w3063_,
		_w3067_,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w3070_
	);
	LUT3 #(
		.INIT('h80)
	) name1721 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3071_
	);
	LUT4 #(
		.INIT('h8000)
	) name1722 (
		_w3060_,
		_w3063_,
		_w3067_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w3073_
	);
	LUT3 #(
		.INIT('h80)
	) name1724 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3074_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3075_
	);
	LUT4 #(
		.INIT('h8000)
	) name1726 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w3076_
	);
	LUT3 #(
		.INIT('h80)
	) name1727 (
		_w3072_,
		_w3074_,
		_w3076_,
		_w3077_
	);
	LUT4 #(
		.INIT('h8000)
	) name1728 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3076_,
		_w3078_
	);
	LUT3 #(
		.INIT('h80)
	) name1729 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('h8000)
	) name1730 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3078_,
		_w3080_
	);
	LUT4 #(
		.INIT('h8000)
	) name1731 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h6)
	) name1732 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name1733 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3083_
	);
	LUT4 #(
		.INIT('h8000)
	) name1734 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3084_
	);
	LUT4 #(
		.INIT('h8000)
	) name1735 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3084_,
		_w3085_
	);
	LUT3 #(
		.INIT('h80)
	) name1736 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('h8000)
	) name1737 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3085_,
		_w3087_
	);
	LUT4 #(
		.INIT('h8000)
	) name1738 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3062_,
		_w3064_,
		_w3088_
	);
	LUT4 #(
		.INIT('h8000)
	) name1739 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3088_,
		_w3089_
	);
	LUT3 #(
		.INIT('h0e)
	) name1740 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w3087_,
		_w3089_,
		_w3090_
	);
	LUT4 #(
		.INIT('h135f)
	) name1741 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1694_,
		_w1711_,
		_w3091_
	);
	LUT4 #(
		.INIT('h135f)
	) name1742 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1703_,
		_w1705_,
		_w3092_
	);
	LUT4 #(
		.INIT('h135f)
	) name1743 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1688_,
		_w1708_,
		_w3093_
	);
	LUT4 #(
		.INIT('h135f)
	) name1744 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w1696_,
		_w1698_,
		_w3094_
	);
	LUT4 #(
		.INIT('h8000)
	) name1745 (
		_w3093_,
		_w3094_,
		_w3091_,
		_w3092_,
		_w3095_
	);
	LUT4 #(
		.INIT('h153f)
	) name1746 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1692_,
		_w1706_,
		_w3096_
	);
	LUT4 #(
		.INIT('h135f)
	) name1747 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1709_,
		_w1702_,
		_w3097_
	);
	LUT4 #(
		.INIT('h135f)
	) name1748 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1691_,
		_w1712_,
		_w3098_
	);
	LUT4 #(
		.INIT('h135f)
	) name1749 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1699_,
		_w1689_,
		_w3099_
	);
	LUT4 #(
		.INIT('h8000)
	) name1750 (
		_w3098_,
		_w3099_,
		_w3096_,
		_w3097_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		_w3095_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h6)
	) name1752 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w3085_,
		_w3102_
	);
	LUT3 #(
		.INIT('h08)
	) name1753 (
		_w3095_,
		_w3100_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h135f)
	) name1754 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1698_,
		_w1702_,
		_w3104_
	);
	LUT4 #(
		.INIT('h135f)
	) name1755 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1696_,
		_w1712_,
		_w3105_
	);
	LUT4 #(
		.INIT('h153f)
	) name1756 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1688_,
		_w1705_,
		_w3106_
	);
	LUT4 #(
		.INIT('h153f)
	) name1757 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1709_,
		_w1703_,
		_w3107_
	);
	LUT4 #(
		.INIT('h8000)
	) name1758 (
		_w3106_,
		_w3107_,
		_w3104_,
		_w3105_,
		_w3108_
	);
	LUT4 #(
		.INIT('h135f)
	) name1759 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1699_,
		_w1691_,
		_w3109_
	);
	LUT4 #(
		.INIT('h135f)
	) name1760 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1689_,
		_w1711_,
		_w3110_
	);
	LUT4 #(
		.INIT('h153f)
	) name1761 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1708_,
		_w1706_,
		_w3111_
	);
	LUT4 #(
		.INIT('h135f)
	) name1762 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1694_,
		_w1692_,
		_w3112_
	);
	LUT4 #(
		.INIT('h8000)
	) name1763 (
		_w3111_,
		_w3112_,
		_w3109_,
		_w3110_,
		_w3113_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		_w3108_,
		_w3113_,
		_w3114_
	);
	LUT3 #(
		.INIT('h6c)
	) name1765 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w3084_,
		_w3115_
	);
	LUT3 #(
		.INIT('h08)
	) name1766 (
		_w3108_,
		_w3113_,
		_w3115_,
		_w3116_
	);
	LUT4 #(
		.INIT('h153f)
	) name1767 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1699_,
		_w1705_,
		_w3117_
	);
	LUT4 #(
		.INIT('h135f)
	) name1768 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1688_,
		_w1708_,
		_w3118_
	);
	LUT4 #(
		.INIT('h135f)
	) name1769 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1692_,
		_w1709_,
		_w3119_
	);
	LUT4 #(
		.INIT('h135f)
	) name1770 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1689_,
		_w1711_,
		_w3120_
	);
	LUT4 #(
		.INIT('h8000)
	) name1771 (
		_w3119_,
		_w3120_,
		_w3117_,
		_w3118_,
		_w3121_
	);
	LUT4 #(
		.INIT('h135f)
	) name1772 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1691_,
		_w1712_,
		_w3122_
	);
	LUT4 #(
		.INIT('h153f)
	) name1773 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1702_,
		_w1706_,
		_w3123_
	);
	LUT4 #(
		.INIT('h135f)
	) name1774 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w1694_,
		_w1696_,
		_w3124_
	);
	LUT4 #(
		.INIT('h153f)
	) name1775 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w1698_,
		_w1703_,
		_w3125_
	);
	LUT4 #(
		.INIT('h8000)
	) name1776 (
		_w3124_,
		_w3125_,
		_w3122_,
		_w3123_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w3121_,
		_w3126_,
		_w3127_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1778 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3084_,
		_w3128_
	);
	LUT3 #(
		.INIT('h08)
	) name1779 (
		_w3121_,
		_w3126_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name1780 (
		_w3116_,
		_w3129_,
		_w3130_
	);
	LUT3 #(
		.INIT('h01)
	) name1781 (
		_w3103_,
		_w3116_,
		_w3129_,
		_w3131_
	);
	LUT4 #(
		.INIT('h135f)
	) name1782 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w1694_,
		_w1692_,
		_w3132_
	);
	LUT4 #(
		.INIT('h153f)
	) name1783 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1712_,
		_w1705_,
		_w3133_
	);
	LUT4 #(
		.INIT('h153f)
	) name1784 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w1698_,
		_w1706_,
		_w3134_
	);
	LUT4 #(
		.INIT('h153f)
	) name1785 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1688_,
		_w1703_,
		_w3135_
	);
	LUT4 #(
		.INIT('h8000)
	) name1786 (
		_w3134_,
		_w3135_,
		_w3132_,
		_w3133_,
		_w3136_
	);
	LUT4 #(
		.INIT('h153f)
	) name1787 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1708_,
		_w1702_,
		_w3137_
	);
	LUT4 #(
		.INIT('h135f)
	) name1788 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1709_,
		_w1711_,
		_w3138_
	);
	LUT4 #(
		.INIT('h135f)
	) name1789 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1696_,
		_w1691_,
		_w3139_
	);
	LUT4 #(
		.INIT('h135f)
	) name1790 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1699_,
		_w1689_,
		_w3140_
	);
	LUT4 #(
		.INIT('h8000)
	) name1791 (
		_w3139_,
		_w3140_,
		_w3137_,
		_w3138_,
		_w3141_
	);
	LUT2 #(
		.INIT('h6)
	) name1792 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w3084_,
		_w3142_
	);
	LUT3 #(
		.INIT('h08)
	) name1793 (
		_w3136_,
		_w3141_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('h135f)
	) name1794 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1696_,
		_w1688_,
		_w3144_
	);
	LUT4 #(
		.INIT('h153f)
	) name1795 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1689_,
		_w1709_,
		_w3145_
	);
	LUT4 #(
		.INIT('h153f)
	) name1796 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1691_,
		_w1705_,
		_w3146_
	);
	LUT4 #(
		.INIT('h153f)
	) name1797 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1708_,
		_w1702_,
		_w3147_
	);
	LUT4 #(
		.INIT('h8000)
	) name1798 (
		_w3146_,
		_w3147_,
		_w3144_,
		_w3145_,
		_w3148_
	);
	LUT4 #(
		.INIT('h153f)
	) name1799 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w1694_,
		_w1703_,
		_w3149_
	);
	LUT4 #(
		.INIT('h135f)
	) name1800 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1692_,
		_w1712_,
		_w3150_
	);
	LUT4 #(
		.INIT('h153f)
	) name1801 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w1698_,
		_w1706_,
		_w3151_
	);
	LUT4 #(
		.INIT('h135f)
	) name1802 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1699_,
		_w1711_,
		_w3152_
	);
	LUT4 #(
		.INIT('h8000)
	) name1803 (
		_w3151_,
		_w3152_,
		_w3149_,
		_w3150_,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		_w3148_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h6)
	) name1805 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3155_
	);
	LUT3 #(
		.INIT('h08)
	) name1806 (
		_w3148_,
		_w3153_,
		_w3155_,
		_w3156_
	);
	LUT3 #(
		.INIT('h15)
	) name1807 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3148_,
		_w3153_,
		_w3157_
	);
	LUT4 #(
		.INIT('h153f)
	) name1808 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1708_,
		_w1711_,
		_w3158_
	);
	LUT4 #(
		.INIT('h135f)
	) name1809 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1696_,
		_w1712_,
		_w3159_
	);
	LUT4 #(
		.INIT('h135f)
	) name1810 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1698_,
		_w1688_,
		_w3160_
	);
	LUT4 #(
		.INIT('h153f)
	) name1811 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1709_,
		_w1705_,
		_w3161_
	);
	LUT4 #(
		.INIT('h8000)
	) name1812 (
		_w3160_,
		_w3161_,
		_w3158_,
		_w3159_,
		_w3162_
	);
	LUT4 #(
		.INIT('h135f)
	) name1813 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1694_,
		_w1692_,
		_w3163_
	);
	LUT4 #(
		.INIT('h153f)
	) name1814 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1691_,
		_w1703_,
		_w3164_
	);
	LUT4 #(
		.INIT('h153f)
	) name1815 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1689_,
		_w1706_,
		_w3165_
	);
	LUT4 #(
		.INIT('h135f)
	) name1816 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1699_,
		_w1702_,
		_w3166_
	);
	LUT4 #(
		.INIT('h8000)
	) name1817 (
		_w3165_,
		_w3166_,
		_w3163_,
		_w3164_,
		_w3167_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w3162_,
		_w3167_,
		_w3168_
	);
	LUT3 #(
		.INIT('h80)
	) name1819 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3162_,
		_w3167_,
		_w3169_
	);
	LUT3 #(
		.INIT('h23)
	) name1820 (
		_w3157_,
		_w3156_,
		_w3169_,
		_w3170_
	);
	LUT4 #(
		.INIT('h153f)
	) name1821 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1691_,
		_w1692_,
		_w3171_
	);
	LUT4 #(
		.INIT('h135f)
	) name1822 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1708_,
		_w1712_,
		_w3172_
	);
	LUT4 #(
		.INIT('h153f)
	) name1823 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1711_,
		_w1706_,
		_w3173_
	);
	LUT4 #(
		.INIT('h135f)
	) name1824 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w1696_,
		_w1705_,
		_w3174_
	);
	LUT4 #(
		.INIT('h8000)
	) name1825 (
		_w3173_,
		_w3174_,
		_w3171_,
		_w3172_,
		_w3175_
	);
	LUT4 #(
		.INIT('h135f)
	) name1826 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1698_,
		_w1689_,
		_w3176_
	);
	LUT4 #(
		.INIT('h135f)
	) name1827 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1694_,
		_w1709_,
		_w3177_
	);
	LUT4 #(
		.INIT('h153f)
	) name1828 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w1699_,
		_w1703_,
		_w3178_
	);
	LUT4 #(
		.INIT('h135f)
	) name1829 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1688_,
		_w1702_,
		_w3179_
	);
	LUT4 #(
		.INIT('h8000)
	) name1830 (
		_w3178_,
		_w3179_,
		_w3176_,
		_w3177_,
		_w3180_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1831 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3181_
	);
	LUT3 #(
		.INIT('h08)
	) name1832 (
		_w3175_,
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT4 #(
		.INIT('h153f)
	) name1833 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1691_,
		_w1703_,
		_w3183_
	);
	LUT4 #(
		.INIT('h135f)
	) name1834 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1698_,
		_w1689_,
		_w3184_
	);
	LUT4 #(
		.INIT('h135f)
	) name1835 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1694_,
		_w1709_,
		_w3185_
	);
	LUT4 #(
		.INIT('h153f)
	) name1836 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1708_,
		_w1705_,
		_w3186_
	);
	LUT4 #(
		.INIT('h8000)
	) name1837 (
		_w3185_,
		_w3186_,
		_w3183_,
		_w3184_,
		_w3187_
	);
	LUT4 #(
		.INIT('h0200)
	) name1838 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name1839 (
		_w1883_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h8)
	) name1840 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1702_,
		_w3190_
	);
	LUT4 #(
		.INIT('h135f)
	) name1841 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1688_,
		_w1711_,
		_w3191_
	);
	LUT4 #(
		.INIT('h153f)
	) name1842 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w1696_,
		_w1706_,
		_w3192_
	);
	LUT4 #(
		.INIT('h135f)
	) name1843 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1699_,
		_w1712_,
		_w3193_
	);
	LUT4 #(
		.INIT('h4000)
	) name1844 (
		_w3190_,
		_w3192_,
		_w3193_,
		_w3191_,
		_w3194_
	);
	LUT3 #(
		.INIT('h40)
	) name1845 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3195_
	);
	LUT3 #(
		.INIT('h78)
	) name1846 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w3196_
	);
	LUT4 #(
		.INIT('h0040)
	) name1847 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name1848 (
		_w3182_,
		_w3197_,
		_w3198_
	);
	LUT3 #(
		.INIT('h70)
	) name1849 (
		_w3175_,
		_w3180_,
		_w3181_,
		_w3199_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1850 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3196_,
		_w3200_
	);
	LUT3 #(
		.INIT('h23)
	) name1851 (
		_w3182_,
		_w3199_,
		_w3200_,
		_w3201_
	);
	LUT3 #(
		.INIT('h70)
	) name1852 (
		_w3170_,
		_w3198_,
		_w3201_,
		_w3202_
	);
	LUT4 #(
		.INIT('h4055)
	) name1853 (
		_w3143_,
		_w3170_,
		_w3198_,
		_w3201_,
		_w3203_
	);
	LUT3 #(
		.INIT('h70)
	) name1854 (
		_w3136_,
		_w3141_,
		_w3142_,
		_w3204_
	);
	LUT3 #(
		.INIT('h70)
	) name1855 (
		_w3108_,
		_w3113_,
		_w3115_,
		_w3205_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w3204_,
		_w3205_,
		_w3206_
	);
	LUT3 #(
		.INIT('h70)
	) name1857 (
		_w3095_,
		_w3100_,
		_w3102_,
		_w3207_
	);
	LUT3 #(
		.INIT('h70)
	) name1858 (
		_w3121_,
		_w3126_,
		_w3128_,
		_w3208_
	);
	LUT3 #(
		.INIT('h54)
	) name1859 (
		_w3103_,
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT3 #(
		.INIT('h6c)
	) name1860 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3085_,
		_w3210_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1861 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3085_,
		_w3211_
	);
	LUT4 #(
		.INIT('h8103)
	) name1862 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3085_,
		_w3212_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1863 (
		_w3101_,
		_w3102_,
		_w3208_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('h7500)
	) name1864 (
		_w3131_,
		_w3203_,
		_w3206_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h8)
	) name1865 (
		_w3067_,
		_w3085_,
		_w3215_
	);
	LUT3 #(
		.INIT('h0e)
	) name1866 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w3089_,
		_w3215_,
		_w3216_
	);
	LUT4 #(
		.INIT('h8000)
	) name1867 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3063_,
		_w3067_,
		_w3217_
	);
	LUT3 #(
		.INIT('h80)
	) name1868 (
		_w3060_,
		_w3067_,
		_w3085_,
		_w3218_
	);
	LUT3 #(
		.INIT('h0e)
	) name1869 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3217_,
		_w3218_,
		_w3219_
	);
	LUT3 #(
		.INIT('h15)
	) name1870 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3067_,
		_w3085_,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name1871 (
		_w3217_,
		_w3220_,
		_w3221_
	);
	LUT4 #(
		.INIT('h8001)
	) name1872 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3215_,
		_w3217_,
		_w3222_
	);
	LUT2 #(
		.INIT('h4)
	) name1873 (
		_w3216_,
		_w3222_,
		_w3223_
	);
	LUT3 #(
		.INIT('h40)
	) name1874 (
		_w3090_,
		_w3214_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('h8000)
	) name1875 (
		_w3060_,
		_w3067_,
		_w3071_,
		_w3085_,
		_w3225_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w3074_,
		_w3225_,
		_w3226_
	);
	LUT3 #(
		.INIT('h80)
	) name1877 (
		_w3074_,
		_w3076_,
		_w3225_,
		_w3227_
	);
	LUT4 #(
		.INIT('h1555)
	) name1878 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3074_,
		_w3076_,
		_w3225_,
		_w3228_
	);
	LUT3 #(
		.INIT('h07)
	) name1879 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3078_,
		_w3228_,
		_w3229_
	);
	LUT3 #(
		.INIT('h80)
	) name1880 (
		_w3072_,
		_w3074_,
		_w3075_,
		_w3230_
	);
	LUT4 #(
		.INIT('h8000)
	) name1881 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3075_,
		_w3231_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1882 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w3231_,
		_w3227_,
		_w3232_
	);
	LUT4 #(
		.INIT('h8000)
	) name1883 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3233_
	);
	LUT3 #(
		.INIT('h80)
	) name1884 (
		_w3074_,
		_w3075_,
		_w3225_,
		_w3234_
	);
	LUT3 #(
		.INIT('h0e)
	) name1885 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3233_,
		_w3234_,
		_w3235_
	);
	LUT4 #(
		.INIT('h1555)
	) name1886 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3074_,
		_w3075_,
		_w3225_,
		_w3236_
	);
	LUT3 #(
		.INIT('h07)
	) name1887 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3231_,
		_w3236_,
		_w3237_
	);
	LUT3 #(
		.INIT('h01)
	) name1888 (
		_w3232_,
		_w3235_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('h0001)
	) name1889 (
		_w3229_,
		_w3232_,
		_w3235_,
		_w3237_,
		_w3239_
	);
	LUT3 #(
		.INIT('h6c)
	) name1890 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3078_,
		_w3240_
	);
	LUT4 #(
		.INIT('h8000)
	) name1891 (
		_w3060_,
		_w3063_,
		_w3067_,
		_w3070_,
		_w3241_
	);
	LUT4 #(
		.INIT('h8000)
	) name1892 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3060_,
		_w3067_,
		_w3085_,
		_w3242_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name1893 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1894 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w3072_,
		_w3244_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name1895 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3072_,
		_w3225_,
		_w3245_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1896 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3241_,
		_w3225_,
		_w3246_
	);
	LUT3 #(
		.INIT('h01)
	) name1897 (
		_w3245_,
		_w3246_,
		_w3244_,
		_w3247_
	);
	LUT4 #(
		.INIT('h0001)
	) name1898 (
		_w3243_,
		_w3245_,
		_w3246_,
		_w3244_,
		_w3248_
	);
	LUT4 #(
		.INIT('h1333)
	) name1899 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3072_,
		_w3073_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w3226_,
		_w3249_,
		_w3250_
	);
	LUT3 #(
		.INIT('h15)
	) name1901 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3074_,
		_w3225_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w3233_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('hf1c0)
	) name1903 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3226_,
		_w3233_,
		_w3249_,
		_w3253_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1904 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3060_,
		_w3067_,
		_w3085_,
		_w3254_
	);
	LUT3 #(
		.INIT('h08)
	) name1905 (
		_w3248_,
		_w3253_,
		_w3254_,
		_w3255_
	);
	LUT3 #(
		.INIT('h20)
	) name1906 (
		_w3239_,
		_w3240_,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('h4000)
	) name1907 (
		_w3090_,
		_w3214_,
		_w3223_,
		_w3256_,
		_w3257_
	);
	LUT3 #(
		.INIT('h6c)
	) name1908 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3080_,
		_w3258_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1909 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3078_,
		_w3259_
	);
	LUT3 #(
		.INIT('h6c)
	) name1910 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3079_,
		_w3260_
	);
	LUT4 #(
		.INIT('h0093)
	) name1911 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3079_,
		_w3259_,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w3258_,
		_w3261_,
		_w3262_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1913 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3080_,
		_w3263_
	);
	LUT3 #(
		.INIT('h04)
	) name1914 (
		_w3258_,
		_w3261_,
		_w3263_,
		_w3264_
	);
	LUT3 #(
		.INIT('h40)
	) name1915 (
		_w3082_,
		_w3257_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('h4111)
	) name1916 (
		_w3101_,
		_w3082_,
		_w3257_,
		_w3264_,
		_w3266_
	);
	LUT2 #(
		.INIT('h6)
	) name1917 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3088_,
		_w3267_
	);
	LUT3 #(
		.INIT('h6c)
	) name1918 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3063_,
		_w3268_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1919 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w3062_,
		_w3269_
	);
	LUT3 #(
		.INIT('h08)
	) name1920 (
		_w3095_,
		_w3100_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('hf070)
	) name1921 (
		_w3095_,
		_w3100_,
		_w3268_,
		_w3269_,
		_w3271_
	);
	LUT2 #(
		.INIT('h6)
	) name1922 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w3272_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1923 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('h0040)
	) name1924 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3272_,
		_w3274_
	);
	LUT3 #(
		.INIT('h2a)
	) name1925 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3162_,
		_w3167_,
		_w3275_
	);
	LUT4 #(
		.INIT('h1301)
	) name1926 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3274_,
		_w3154_,
		_w3275_,
		_w3276_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1927 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w3277_
	);
	LUT3 #(
		.INIT('h40)
	) name1928 (
		_w3277_,
		_w3136_,
		_w3141_,
		_w3278_
	);
	LUT3 #(
		.INIT('h78)
	) name1929 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3279_
	);
	LUT3 #(
		.INIT('h08)
	) name1930 (
		_w3175_,
		_w3180_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w3278_,
		_w3280_,
		_w3281_
	);
	LUT3 #(
		.INIT('h2a)
	) name1932 (
		_w3277_,
		_w3136_,
		_w3141_,
		_w3282_
	);
	LUT3 #(
		.INIT('h70)
	) name1933 (
		_w3175_,
		_w3180_,
		_w3279_,
		_w3283_
	);
	LUT3 #(
		.INIT('h23)
	) name1934 (
		_w3278_,
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1935 (
		_w3273_,
		_w3276_,
		_w3281_,
		_w3284_,
		_w3285_
	);
	LUT3 #(
		.INIT('h6c)
	) name1936 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3062_,
		_w3286_
	);
	LUT3 #(
		.INIT('h40)
	) name1937 (
		_w3286_,
		_w3121_,
		_w3126_,
		_w3287_
	);
	LUT2 #(
		.INIT('h6)
	) name1938 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w3062_,
		_w3288_
	);
	LUT3 #(
		.INIT('h40)
	) name1939 (
		_w3288_,
		_w3108_,
		_w3113_,
		_w3289_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w3287_,
		_w3289_,
		_w3290_
	);
	LUT3 #(
		.INIT('h70)
	) name1941 (
		_w3095_,
		_w3100_,
		_w3269_,
		_w3291_
	);
	LUT3 #(
		.INIT('h2a)
	) name1942 (
		_w3286_,
		_w3121_,
		_w3126_,
		_w3292_
	);
	LUT3 #(
		.INIT('h2a)
	) name1943 (
		_w3288_,
		_w3108_,
		_w3113_,
		_w3293_
	);
	LUT3 #(
		.INIT('h23)
	) name1944 (
		_w3287_,
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT4 #(
		.INIT('h040d)
	) name1945 (
		_w3286_,
		_w3127_,
		_w3291_,
		_w3293_,
		_w3295_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1946 (
		_w3271_,
		_w3285_,
		_w3290_,
		_w3295_,
		_w3296_
	);
	LUT3 #(
		.INIT('h32)
	) name1947 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3072_,
		_w3241_,
		_w3297_
	);
	LUT4 #(
		.INIT('h4888)
	) name1948 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3069_,
		_w3070_,
		_w3298_
	);
	LUT4 #(
		.INIT('h1333)
	) name1949 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3088_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w3068_,
		_w3299_,
		_w3300_
	);
	LUT3 #(
		.INIT('h02)
	) name1951 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3068_,
		_w3299_,
		_w3301_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1952 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3063_,
		_w3067_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name1953 (
		_w3070_,
		_w3302_,
		_w3303_
	);
	LUT3 #(
		.INIT('h80)
	) name1954 (
		_w3301_,
		_w3298_,
		_w3303_,
		_w3304_
	);
	LUT3 #(
		.INIT('h6c)
	) name1955 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w3072_,
		_w3305_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1956 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3072_,
		_w3306_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3306_,
		_w3307_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1958 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3308_
	);
	LUT3 #(
		.INIT('h6a)
	) name1959 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3088_,
		_w3309_
	);
	LUT4 #(
		.INIT('h8000)
	) name1960 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3308_,
		_w3309_,
		_w3306_,
		_w3310_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		_w3304_,
		_w3310_,
		_w3311_
	);
	LUT3 #(
		.INIT('h80)
	) name1962 (
		_w3267_,
		_w3296_,
		_w3311_,
		_w3312_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1963 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3075_,
		_w3313_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1964 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3078_,
		_w3314_
	);
	LUT3 #(
		.INIT('h0e)
	) name1965 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w3231_,
		_w3077_,
		_w3315_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1966 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3231_,
		_w3077_,
		_w3316_
	);
	LUT2 #(
		.INIT('h6)
	) name1967 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3078_,
		_w3317_
	);
	LUT3 #(
		.INIT('h48)
	) name1968 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3078_,
		_w3318_
	);
	LUT4 #(
		.INIT('h8000)
	) name1969 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3316_,
		_w3318_,
		_w3314_,
		_w3319_
	);
	LUT3 #(
		.INIT('h80)
	) name1970 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3313_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h8000)
	) name1971 (
		_w3267_,
		_w3296_,
		_w3311_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3322_
	);
	LUT3 #(
		.INIT('h6a)
	) name1973 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3080_,
		_w3322_,
		_w3323_
	);
	LUT4 #(
		.INIT('h1551)
	) name1974 (
		_w1916_,
		_w3101_,
		_w3321_,
		_w3323_,
		_w3324_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1975 (
		_w1810_,
		_w3059_,
		_w3266_,
		_w3324_,
		_w3325_
	);
	LUT4 #(
		.INIT('hf800)
	) name1976 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3326_
	);
	LUT3 #(
		.INIT('h6c)
	) name1977 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w3326_,
		_w3327_
	);
	LUT3 #(
		.INIT('h08)
	) name1978 (
		_w3108_,
		_w3113_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h6)
	) name1979 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w3326_,
		_w3329_
	);
	LUT3 #(
		.INIT('h08)
	) name1980 (
		_w3136_,
		_w3141_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name1981 (
		_w3328_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1982 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w3332_
	);
	LUT3 #(
		.INIT('h08)
	) name1983 (
		_w3175_,
		_w3180_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('h4000)
	) name1984 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3196_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name1985 (
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('h70)
	) name1986 (
		_w3148_,
		_w3153_,
		_w3155_,
		_w3336_
	);
	LUT3 #(
		.INIT('h15)
	) name1987 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3162_,
		_w3167_,
		_w3337_
	);
	LUT3 #(
		.INIT('h54)
	) name1988 (
		_w3156_,
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT3 #(
		.INIT('h70)
	) name1989 (
		_w3175_,
		_w3180_,
		_w3332_,
		_w3339_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1990 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3196_,
		_w3340_
	);
	LUT3 #(
		.INIT('h23)
	) name1991 (
		_w3333_,
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT3 #(
		.INIT('h70)
	) name1992 (
		_w3335_,
		_w3338_,
		_w3341_,
		_w3342_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1993 (
		_w3331_,
		_w3335_,
		_w3338_,
		_w3341_,
		_w3343_
	);
	LUT3 #(
		.INIT('h70)
	) name1994 (
		_w3108_,
		_w3113_,
		_w3327_,
		_w3344_
	);
	LUT3 #(
		.INIT('h70)
	) name1995 (
		_w3136_,
		_w3141_,
		_w3329_,
		_w3345_
	);
	LUT3 #(
		.INIT('h23)
	) name1996 (
		_w3328_,
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT4 #(
		.INIT('h8000)
	) name1997 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3326_,
		_w3347_
	);
	LUT2 #(
		.INIT('h6)
	) name1998 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w3347_,
		_w3348_
	);
	LUT3 #(
		.INIT('h08)
	) name1999 (
		_w3095_,
		_w3100_,
		_w3348_,
		_w3349_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2000 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w3326_,
		_w3350_
	);
	LUT3 #(
		.INIT('h08)
	) name2001 (
		_w3121_,
		_w3126_,
		_w3350_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w3349_,
		_w3351_,
		_w3352_
	);
	LUT3 #(
		.INIT('h70)
	) name2003 (
		_w3095_,
		_w3100_,
		_w3348_,
		_w3353_
	);
	LUT3 #(
		.INIT('h70)
	) name2004 (
		_w3121_,
		_w3126_,
		_w3350_,
		_w3354_
	);
	LUT3 #(
		.INIT('h23)
	) name2005 (
		_w3349_,
		_w3353_,
		_w3354_,
		_w3355_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2006 (
		_w3343_,
		_w3346_,
		_w3352_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h8)
	) name2007 (
		_w3064_,
		_w3347_,
		_w3357_
	);
	LUT3 #(
		.INIT('h6c)
	) name2008 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3347_,
		_w3358_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2009 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3347_,
		_w3359_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2010 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3064_,
		_w3347_,
		_w3360_
	);
	LUT4 #(
		.INIT('h8000)
	) name2011 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w3065_,
		_w3064_,
		_w3347_,
		_w3361_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2012 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w3065_,
		_w3064_,
		_w3347_,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		_w3060_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h4000)
	) name2014 (
		_w3356_,
		_w3359_,
		_w3360_,
		_w3363_,
		_w3364_
	);
	LUT3 #(
		.INIT('h80)
	) name2015 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3361_,
		_w3365_
	);
	LUT4 #(
		.INIT('h8000)
	) name2016 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3071_,
		_w3361_,
		_w3366_
	);
	LUT4 #(
		.INIT('h8000)
	) name2017 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3361_,
		_w3367_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2018 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w3365_,
		_w3368_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2019 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3361_,
		_w3369_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3370_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w3368_,
		_w3371_,
		_w3372_
	);
	LUT3 #(
		.INIT('h6c)
	) name2023 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w3366_,
		_w3373_
	);
	LUT3 #(
		.INIT('h6a)
	) name2024 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3073_,
		_w3366_,
		_w3374_
	);
	LUT4 #(
		.INIT('h60a0)
	) name2025 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3073_,
		_w3075_,
		_w3366_,
		_w3375_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w3373_,
		_w3375_,
		_w3376_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		_w3364_,
		_w3372_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h80)
	) name2028 (
		_w3074_,
		_w3076_,
		_w3366_,
		_w3378_
	);
	LUT4 #(
		.INIT('h8000)
	) name2029 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3074_,
		_w3076_,
		_w3366_,
		_w3379_
	);
	LUT2 #(
		.INIT('h6)
	) name2030 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h8000)
	) name2031 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3074_,
		_w3075_,
		_w3366_,
		_w3381_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2032 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3074_,
		_w3075_,
		_w3366_,
		_w3382_
	);
	LUT3 #(
		.INIT('h80)
	) name2033 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2034 (
		_w3380_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('h8000)
	) name2035 (
		_w3364_,
		_w3372_,
		_w3376_,
		_w3384_,
		_w3385_
	);
	LUT3 #(
		.INIT('h6c)
	) name2036 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3379_,
		_w3386_
	);
	LUT4 #(
		.INIT('h8000)
	) name2037 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3379_,
		_w3387_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2038 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3379_,
		_w3388_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		_w3322_,
		_w3388_,
		_w3389_
	);
	LUT3 #(
		.INIT('h6a)
	) name2040 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3322_,
		_w3387_,
		_w3390_
	);
	LUT4 #(
		.INIT('h007f)
	) name2041 (
		_w3385_,
		_w3386_,
		_w3389_,
		_w3390_,
		_w3391_
	);
	LUT3 #(
		.INIT('h80)
	) name2042 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3322_,
		_w3388_,
		_w3392_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2043 (
		_w1924_,
		_w3385_,
		_w3386_,
		_w3392_,
		_w3393_
	);
	LUT4 #(
		.INIT('h8444)
	) name2044 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1846_,
		_w3322_,
		_w3387_,
		_w3394_
	);
	LUT3 #(
		.INIT('h54)
	) name2045 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1842_,
		_w1845_,
		_w3395_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		_w1833_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w3394_,
		_w3396_,
		_w3397_
	);
	LUT4 #(
		.INIT('h8444)
	) name2048 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1867_,
		_w3080_,
		_w3322_,
		_w3398_
	);
	LUT4 #(
		.INIT('h0203)
	) name2049 (
		_w1725_,
		_w1795_,
		_w1797_,
		_w1802_,
		_w3399_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name2050 (
		_w1852_,
		_w1853_,
		_w3398_,
		_w3399_,
		_w3400_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2051 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w1913_,
		_w1922_,
		_w3400_,
		_w3401_
	);
	LUT3 #(
		.INIT('hb0)
	) name2052 (
		_w1816_,
		_w1831_,
		_w3082_,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name2053 (
		_w1862_,
		_w3323_,
		_w3403_
	);
	LUT4 #(
		.INIT('h0001)
	) name2054 (
		_w3402_,
		_w3397_,
		_w3403_,
		_w3401_,
		_w3404_
	);
	LUT4 #(
		.INIT('h4500)
	) name2055 (
		_w3325_,
		_w3391_,
		_w3393_,
		_w3404_,
		_w3405_
	);
	LUT4 #(
		.INIT('h0001)
	) name2056 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3406_
	);
	LUT4 #(
		.INIT('h0010)
	) name2057 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3407_
	);
	LUT4 #(
		.INIT('hfc21)
	) name2058 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3408_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2059 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w3406_,
		_w3408_,
		_w3409_
	);
	LUT3 #(
		.INIT('h2f)
	) name2060 (
		_w1933_,
		_w3405_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h0100)
	) name2061 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3411_
	);
	LUT4 #(
		.INIT('h0200)
	) name2062 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3412_
	);
	LUT4 #(
		.INIT('hfcff)
	) name2063 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3413_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('h0001)
	) name2065 (
		\address1[26]_pad ,
		\address1[27]_pad ,
		\address1[28]_pad ,
		\address1[2]_pad ,
		_w3415_
	);
	LUT4 #(
		.INIT('h0001)
	) name2066 (
		\address1[22]_pad ,
		\address1[23]_pad ,
		\address1[24]_pad ,
		\address1[25]_pad ,
		_w3416_
	);
	LUT3 #(
		.INIT('h01)
	) name2067 (
		\address1[7]_pad ,
		\address1[8]_pad ,
		\address1[9]_pad ,
		_w3417_
	);
	LUT4 #(
		.INIT('h0001)
	) name2068 (
		\address1[3]_pad ,
		\address1[4]_pad ,
		\address1[5]_pad ,
		\address1[6]_pad ,
		_w3418_
	);
	LUT4 #(
		.INIT('h8000)
	) name2069 (
		_w3417_,
		_w3418_,
		_w3415_,
		_w3416_,
		_w3419_
	);
	LUT2 #(
		.INIT('h1)
	) name2070 (
		\address1[0]_pad ,
		\address1[10]_pad ,
		_w3420_
	);
	LUT4 #(
		.INIT('h0001)
	) name2071 (
		\address1[11]_pad ,
		\address1[12]_pad ,
		\address1[13]_pad ,
		\address1[14]_pad ,
		_w3421_
	);
	LUT4 #(
		.INIT('h0001)
	) name2072 (
		\address1[19]_pad ,
		\address1[1]_pad ,
		\address1[20]_pad ,
		\address1[21]_pad ,
		_w3422_
	);
	LUT4 #(
		.INIT('h0001)
	) name2073 (
		\address1[15]_pad ,
		\address1[16]_pad ,
		\address1[17]_pad ,
		\address1[18]_pad ,
		_w3423_
	);
	LUT4 #(
		.INIT('h8000)
	) name2074 (
		_w3420_,
		_w3422_,
		_w3423_,
		_w3421_,
		_w3424_
	);
	LUT4 #(
		.INIT('hc444)
	) name2075 (
		\address1[29]_pad ,
		\datai[31]_pad ,
		_w3419_,
		_w3424_,
		_w3425_
	);
	LUT4 #(
		.INIT('hc444)
	) name2076 (
		\address1[29]_pad ,
		\datai[3]_pad ,
		_w3419_,
		_w3424_,
		_w3426_
	);
	LUT4 #(
		.INIT('h0888)
	) name2077 (
		\address1[29]_pad ,
		\buf1_reg[3]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3427_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('hc444)
	) name2079 (
		\address1[29]_pad ,
		\datai[11]_pad ,
		_w3419_,
		_w3424_,
		_w3429_
	);
	LUT4 #(
		.INIT('h0888)
	) name2080 (
		\address1[29]_pad ,
		\buf1_reg[11]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('h0001)
	) name2082 (
		_w3426_,
		_w3427_,
		_w3429_,
		_w3430_,
		_w3432_
	);
	LUT4 #(
		.INIT('hc444)
	) name2083 (
		\address1[29]_pad ,
		\datai[8]_pad ,
		_w3419_,
		_w3424_,
		_w3433_
	);
	LUT4 #(
		.INIT('h0888)
	) name2084 (
		\address1[29]_pad ,
		\buf1_reg[8]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3434_
	);
	LUT2 #(
		.INIT('h1)
	) name2085 (
		_w3433_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('hc444)
	) name2086 (
		\address1[29]_pad ,
		\datai[7]_pad ,
		_w3419_,
		_w3424_,
		_w3436_
	);
	LUT4 #(
		.INIT('h0888)
	) name2087 (
		\address1[29]_pad ,
		\buf1_reg[7]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w3436_,
		_w3437_,
		_w3438_
	);
	LUT4 #(
		.INIT('h0001)
	) name2089 (
		_w3433_,
		_w3434_,
		_w3436_,
		_w3437_,
		_w3439_
	);
	LUT4 #(
		.INIT('hc444)
	) name2090 (
		\address1[29]_pad ,
		\datai[4]_pad ,
		_w3419_,
		_w3424_,
		_w3440_
	);
	LUT4 #(
		.INIT('h0888)
	) name2091 (
		\address1[29]_pad ,
		\buf1_reg[4]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3441_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w3440_,
		_w3441_,
		_w3442_
	);
	LUT4 #(
		.INIT('hc444)
	) name2093 (
		\address1[29]_pad ,
		\datai[9]_pad ,
		_w3419_,
		_w3424_,
		_w3443_
	);
	LUT4 #(
		.INIT('h0888)
	) name2094 (
		\address1[29]_pad ,
		\buf1_reg[9]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		_w3443_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h0001)
	) name2096 (
		_w3440_,
		_w3441_,
		_w3443_,
		_w3444_,
		_w3446_
	);
	LUT4 #(
		.INIT('hc444)
	) name2097 (
		\address1[29]_pad ,
		\datai[10]_pad ,
		_w3419_,
		_w3424_,
		_w3447_
	);
	LUT4 #(
		.INIT('h0888)
	) name2098 (
		\address1[29]_pad ,
		\buf1_reg[10]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name2099 (
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('hc444)
	) name2100 (
		\address1[29]_pad ,
		\datai[5]_pad ,
		_w3419_,
		_w3424_,
		_w3450_
	);
	LUT4 #(
		.INIT('h0888)
	) name2101 (
		\address1[29]_pad ,
		\buf1_reg[5]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2102 (
		_w3450_,
		_w3451_,
		_w3452_
	);
	LUT4 #(
		.INIT('h0001)
	) name2103 (
		_w3447_,
		_w3448_,
		_w3450_,
		_w3451_,
		_w3453_
	);
	LUT4 #(
		.INIT('h8000)
	) name2104 (
		_w3446_,
		_w3453_,
		_w3432_,
		_w3439_,
		_w3454_
	);
	LUT4 #(
		.INIT('hc444)
	) name2105 (
		\address1[29]_pad ,
		\datai[14]_pad ,
		_w3419_,
		_w3424_,
		_w3455_
	);
	LUT4 #(
		.INIT('h0888)
	) name2106 (
		\address1[29]_pad ,
		\buf1_reg[14]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3456_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w3455_,
		_w3456_,
		_w3457_
	);
	LUT4 #(
		.INIT('hc444)
	) name2108 (
		\address1[29]_pad ,
		\datai[15]_pad ,
		_w3419_,
		_w3424_,
		_w3458_
	);
	LUT4 #(
		.INIT('h0888)
	) name2109 (
		\address1[29]_pad ,
		\buf1_reg[15]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3459_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h0001)
	) name2111 (
		_w3455_,
		_w3456_,
		_w3458_,
		_w3459_,
		_w3461_
	);
	LUT4 #(
		.INIT('hc444)
	) name2112 (
		\address1[29]_pad ,
		\datai[12]_pad ,
		_w3419_,
		_w3424_,
		_w3462_
	);
	LUT4 #(
		.INIT('h0888)
	) name2113 (
		\address1[29]_pad ,
		\buf1_reg[12]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3463_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('hc444)
	) name2115 (
		\address1[29]_pad ,
		\datai[13]_pad ,
		_w3419_,
		_w3424_,
		_w3465_
	);
	LUT4 #(
		.INIT('h0888)
	) name2116 (
		\address1[29]_pad ,
		\buf1_reg[13]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT4 #(
		.INIT('h0001)
	) name2118 (
		_w3462_,
		_w3463_,
		_w3465_,
		_w3466_,
		_w3468_
	);
	LUT4 #(
		.INIT('hc444)
	) name2119 (
		\address1[29]_pad ,
		\datai[0]_pad ,
		_w3419_,
		_w3424_,
		_w3469_
	);
	LUT4 #(
		.INIT('h0888)
	) name2120 (
		\address1[29]_pad ,
		\buf1_reg[0]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3470_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		_w3469_,
		_w3470_,
		_w3471_
	);
	LUT4 #(
		.INIT('hc444)
	) name2122 (
		\address1[29]_pad ,
		\datai[6]_pad ,
		_w3419_,
		_w3424_,
		_w3472_
	);
	LUT4 #(
		.INIT('h0888)
	) name2123 (
		\address1[29]_pad ,
		\buf1_reg[6]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3473_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w3472_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h0001)
	) name2125 (
		_w3469_,
		_w3470_,
		_w3472_,
		_w3473_,
		_w3475_
	);
	LUT4 #(
		.INIT('hc444)
	) name2126 (
		\address1[29]_pad ,
		\datai[1]_pad ,
		_w3419_,
		_w3424_,
		_w3476_
	);
	LUT4 #(
		.INIT('h0888)
	) name2127 (
		\address1[29]_pad ,
		\buf1_reg[1]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w3476_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('hc444)
	) name2129 (
		\address1[29]_pad ,
		\datai[2]_pad ,
		_w3419_,
		_w3424_,
		_w3479_
	);
	LUT4 #(
		.INIT('h0888)
	) name2130 (
		\address1[29]_pad ,
		\buf1_reg[2]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3480_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h0001)
	) name2132 (
		_w3476_,
		_w3477_,
		_w3479_,
		_w3480_,
		_w3482_
	);
	LUT4 #(
		.INIT('h8000)
	) name2133 (
		_w3475_,
		_w3482_,
		_w3461_,
		_w3468_,
		_w3483_
	);
	LUT4 #(
		.INIT('hc444)
	) name2134 (
		\address1[29]_pad ,
		\datai[19]_pad ,
		_w3419_,
		_w3424_,
		_w3484_
	);
	LUT4 #(
		.INIT('h0888)
	) name2135 (
		\address1[29]_pad ,
		\buf1_reg[19]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w3484_,
		_w3485_,
		_w3486_
	);
	LUT4 #(
		.INIT('hc444)
	) name2137 (
		\address1[29]_pad ,
		\datai[18]_pad ,
		_w3419_,
		_w3424_,
		_w3487_
	);
	LUT4 #(
		.INIT('h0888)
	) name2138 (
		\address1[29]_pad ,
		\buf1_reg[18]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w3487_,
		_w3488_,
		_w3489_
	);
	LUT4 #(
		.INIT('h0001)
	) name2140 (
		_w3484_,
		_w3485_,
		_w3487_,
		_w3488_,
		_w3490_
	);
	LUT4 #(
		.INIT('hc444)
	) name2141 (
		\address1[29]_pad ,
		\datai[17]_pad ,
		_w3419_,
		_w3424_,
		_w3491_
	);
	LUT4 #(
		.INIT('h0888)
	) name2142 (
		\address1[29]_pad ,
		\buf1_reg[17]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3492_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT4 #(
		.INIT('hc444)
	) name2144 (
		\address1[29]_pad ,
		\datai[20]_pad ,
		_w3419_,
		_w3424_,
		_w3494_
	);
	LUT4 #(
		.INIT('h0888)
	) name2145 (
		\address1[29]_pad ,
		\buf1_reg[20]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3495_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w3494_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('h0001)
	) name2147 (
		_w3491_,
		_w3492_,
		_w3494_,
		_w3495_,
		_w3497_
	);
	LUT4 #(
		.INIT('hc444)
	) name2148 (
		\address1[29]_pad ,
		\datai[16]_pad ,
		_w3419_,
		_w3424_,
		_w3498_
	);
	LUT4 #(
		.INIT('h0888)
	) name2149 (
		\address1[29]_pad ,
		\buf1_reg[16]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3499_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT4 #(
		.INIT('hc444)
	) name2151 (
		\address1[29]_pad ,
		\datai[22]_pad ,
		_w3419_,
		_w3424_,
		_w3501_
	);
	LUT4 #(
		.INIT('h0888)
	) name2152 (
		\address1[29]_pad ,
		\buf1_reg[22]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3502_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		_w3501_,
		_w3502_,
		_w3503_
	);
	LUT4 #(
		.INIT('h0001)
	) name2154 (
		_w3498_,
		_w3499_,
		_w3501_,
		_w3502_,
		_w3504_
	);
	LUT4 #(
		.INIT('hc444)
	) name2155 (
		\address1[29]_pad ,
		\datai[23]_pad ,
		_w3419_,
		_w3424_,
		_w3505_
	);
	LUT4 #(
		.INIT('h0888)
	) name2156 (
		\address1[29]_pad ,
		\buf1_reg[23]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3506_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT4 #(
		.INIT('hc444)
	) name2158 (
		\address1[29]_pad ,
		\datai[21]_pad ,
		_w3419_,
		_w3424_,
		_w3508_
	);
	LUT4 #(
		.INIT('h0888)
	) name2159 (
		\address1[29]_pad ,
		\buf1_reg[21]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3509_
	);
	LUT2 #(
		.INIT('h1)
	) name2160 (
		_w3508_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('h0001)
	) name2161 (
		_w3505_,
		_w3506_,
		_w3508_,
		_w3509_,
		_w3511_
	);
	LUT4 #(
		.INIT('h8000)
	) name2162 (
		_w3504_,
		_w3511_,
		_w3490_,
		_w3497_,
		_w3512_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2163 (
		_w3425_,
		_w3454_,
		_w3483_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('hc444)
	) name2164 (
		\address1[29]_pad ,
		\datai[24]_pad ,
		_w3419_,
		_w3424_,
		_w3514_
	);
	LUT4 #(
		.INIT('h0888)
	) name2165 (
		\address1[29]_pad ,
		\buf1_reg[24]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3515_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT4 #(
		.INIT('hc444)
	) name2167 (
		\address1[29]_pad ,
		\datai[25]_pad ,
		_w3419_,
		_w3424_,
		_w3517_
	);
	LUT4 #(
		.INIT('h0888)
	) name2168 (
		\address1[29]_pad ,
		\buf1_reg[25]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name2169 (
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('hc444)
	) name2170 (
		\address1[29]_pad ,
		\datai[26]_pad ,
		_w3419_,
		_w3424_,
		_w3520_
	);
	LUT4 #(
		.INIT('h0888)
	) name2171 (
		\address1[29]_pad ,
		\buf1_reg[26]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3521_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w3520_,
		_w3521_,
		_w3522_
	);
	LUT4 #(
		.INIT('h0002)
	) name2173 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3522_,
		_w3523_
	);
	LUT4 #(
		.INIT('hc444)
	) name2174 (
		\address1[29]_pad ,
		\datai[27]_pad ,
		_w3419_,
		_w3424_,
		_w3524_
	);
	LUT4 #(
		.INIT('h0888)
	) name2175 (
		\address1[29]_pad ,
		\buf1_reg[27]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('hc444)
	) name2177 (
		\address1[29]_pad ,
		\datai[28]_pad ,
		_w3419_,
		_w3424_,
		_w3527_
	);
	LUT4 #(
		.INIT('h0888)
	) name2178 (
		\address1[29]_pad ,
		\buf1_reg[28]/NET0131 ,
		_w3419_,
		_w3424_,
		_w3528_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w3527_,
		_w3528_,
		_w3529_
	);
	LUT4 #(
		.INIT('ha208)
	) name2180 (
		_w3411_,
		_w3523_,
		_w3526_,
		_w3529_,
		_w3530_
	);
	LUT4 #(
		.INIT('h002a)
	) name2181 (
		_w3425_,
		_w3454_,
		_w3483_,
		_w3500_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0100)
	) name2182 (
		_w3486_,
		_w3489_,
		_w3493_,
		_w3531_,
		_w3532_
	);
	LUT3 #(
		.INIT('h14)
	) name2183 (
		_w3411_,
		_w3496_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h0800)
	) name2184 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3534_
	);
	LUT2 #(
		.INIT('h4)
	) name2185 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w3535_
	);
	LUT4 #(
		.INIT('h0400)
	) name2186 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3536_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name2187 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3537_
	);
	LUT3 #(
		.INIT('h02)
	) name2188 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		_w3534_,
		_w3536_,
		_w3538_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2189 (
		_w3537_,
		_w3440_,
		_w3441_,
		_w3538_,
		_w3539_
	);
	LUT3 #(
		.INIT('ha2)
	) name2190 (
		_w1939_,
		_w3539_,
		_w3414_,
		_w3540_
	);
	LUT4 #(
		.INIT('h5700)
	) name2191 (
		_w3414_,
		_w3530_,
		_w3533_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w3407_,
		_w3539_,
		_w3542_
	);
	LUT4 #(
		.INIT('hc055)
	) name2193 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3534_,
		_w3543_
	);
	LUT4 #(
		.INIT('hfff4)
	) name2194 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3544_
	);
	LUT4 #(
		.INIT('hfd14)
	) name2195 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w3545_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		_w3545_,
		_w3546_
	);
	LUT3 #(
		.INIT('h0d)
	) name2197 (
		_w2248_,
		_w3543_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h4)
	) name2198 (
		_w3542_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('hb)
	) name2199 (
		_w3541_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('hc444)
	) name2200 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3550_
	);
	LUT4 #(
		.INIT('h0888)
	) name2201 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[27]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3551_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		_w3550_,
		_w3551_,
		_w3552_
	);
	LUT3 #(
		.INIT('ha8)
	) name2203 (
		_w2250_,
		_w3550_,
		_w3551_,
		_w3553_
	);
	LUT4 #(
		.INIT('hc444)
	) name2204 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[19]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3554_
	);
	LUT4 #(
		.INIT('h0888)
	) name2205 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[19]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3555_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w3554_,
		_w3555_,
		_w3556_
	);
	LUT3 #(
		.INIT('ha8)
	) name2207 (
		_w2264_,
		_w3554_,
		_w3555_,
		_w3557_
	);
	LUT3 #(
		.INIT('ha8)
	) name2208 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3553_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('hc444)
	) name2209 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3559_
	);
	LUT4 #(
		.INIT('h0888)
	) name2210 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[3]/NET0131 ,
		_w2255_,
		_w2260_,
		_w3560_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w3559_,
		_w3560_,
		_w3561_
	);
	LUT3 #(
		.INIT('h02)
	) name2212 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w2271_,
		_w2272_,
		_w3562_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2213 (
		_w2273_,
		_w3559_,
		_w3560_,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		_w2280_,
		_w3563_,
		_w3564_
	);
	LUT3 #(
		.INIT('ha8)
	) name2215 (
		_w1679_,
		_w3558_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		_w2283_,
		_w3563_,
		_w3566_
	);
	LUT4 #(
		.INIT('hc055)
	) name2217 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2272_,
		_w3567_
	);
	LUT2 #(
		.INIT('h2)
	) name2218 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		_w2288_,
		_w3568_
	);
	LUT3 #(
		.INIT('h0d)
	) name2219 (
		_w2246_,
		_w3567_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h4)
	) name2220 (
		_w3566_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('hb)
	) name2221 (
		_w3565_,
		_w3570_,
		_w3571_
	);
	LUT4 #(
		.INIT('h2000)
	) name2222 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3572_
	);
	LUT4 #(
		.INIT('h4000)
	) name2223 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3573_
	);
	LUT4 #(
		.INIT('h9fff)
	) name2224 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3574_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('hd200)
	) name2226 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3572_,
		_w3576_
	);
	LUT3 #(
		.INIT('h06)
	) name2227 (
		_w3496_,
		_w3532_,
		_w3572_,
		_w3577_
	);
	LUT4 #(
		.INIT('h0001)
	) name2228 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3578_
	);
	LUT3 #(
		.INIT('h80)
	) name2229 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3579_
	);
	LUT4 #(
		.INIT('h8000)
	) name2230 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3580_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name2231 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3581_
	);
	LUT3 #(
		.INIT('h02)
	) name2232 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w3578_,
		_w3580_,
		_w3582_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2233 (
		_w3440_,
		_w3441_,
		_w3581_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('ha2)
	) name2234 (
		_w1939_,
		_w3583_,
		_w3575_,
		_w3584_
	);
	LUT4 #(
		.INIT('h5700)
	) name2235 (
		_w3575_,
		_w3576_,
		_w3577_,
		_w3584_,
		_w3585_
	);
	LUT2 #(
		.INIT('h2)
	) name2236 (
		_w3407_,
		_w3583_,
		_w3586_
	);
	LUT4 #(
		.INIT('hc055)
	) name2237 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3578_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		_w3545_,
		_w3588_
	);
	LUT3 #(
		.INIT('h0d)
	) name2239 (
		_w2248_,
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name2240 (
		_w3586_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('hb)
	) name2241 (
		_w3585_,
		_w3590_,
		_w3591_
	);
	LUT4 #(
		.INIT('h0080)
	) name2242 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3592_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name2243 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3593_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3593_,
		_w3594_
	);
	LUT4 #(
		.INIT('hd200)
	) name2245 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3592_,
		_w3595_
	);
	LUT3 #(
		.INIT('h06)
	) name2246 (
		_w3496_,
		_w3532_,
		_w3592_,
		_w3596_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name2247 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3597_
	);
	LUT3 #(
		.INIT('h02)
	) name2248 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w3536_,
		_w3412_,
		_w3598_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2249 (
		_w3440_,
		_w3441_,
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT3 #(
		.INIT('ha2)
	) name2250 (
		_w1939_,
		_w3599_,
		_w3594_,
		_w3600_
	);
	LUT4 #(
		.INIT('h5700)
	) name2251 (
		_w3594_,
		_w3595_,
		_w3596_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		_w3407_,
		_w3599_,
		_w3602_
	);
	LUT4 #(
		.INIT('hc055)
	) name2253 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3536_,
		_w3603_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		_w3545_,
		_w3604_
	);
	LUT3 #(
		.INIT('h0d)
	) name2255 (
		_w2248_,
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h4)
	) name2256 (
		_w3602_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('hb)
	) name2257 (
		_w3601_,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3597_,
		_w3608_
	);
	LUT4 #(
		.INIT('ha208)
	) name2259 (
		_w3412_,
		_w3523_,
		_w3526_,
		_w3529_,
		_w3609_
	);
	LUT3 #(
		.INIT('h14)
	) name2260 (
		_w3412_,
		_w3496_,
		_w3532_,
		_w3610_
	);
	LUT4 #(
		.INIT('h1000)
	) name2261 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3611_
	);
	LUT4 #(
		.INIT('he7ff)
	) name2262 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3612_
	);
	LUT3 #(
		.INIT('h02)
	) name2263 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w3534_,
		_w3611_,
		_w3613_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2264 (
		_w3440_,
		_w3441_,
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT3 #(
		.INIT('ha2)
	) name2265 (
		_w1939_,
		_w3614_,
		_w3608_,
		_w3615_
	);
	LUT4 #(
		.INIT('h5700)
	) name2266 (
		_w3608_,
		_w3609_,
		_w3610_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h2)
	) name2267 (
		_w3407_,
		_w3614_,
		_w3617_
	);
	LUT4 #(
		.INIT('hc055)
	) name2268 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3611_,
		_w3618_
	);
	LUT2 #(
		.INIT('h2)
	) name2269 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w3545_,
		_w3619_
	);
	LUT3 #(
		.INIT('h0d)
	) name2270 (
		_w2248_,
		_w3618_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h4)
	) name2271 (
		_w3617_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('hb)
	) name2272 (
		_w3616_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h2)
	) name2273 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3537_,
		_w3623_
	);
	LUT4 #(
		.INIT('ha208)
	) name2274 (
		_w3536_,
		_w3523_,
		_w3526_,
		_w3529_,
		_w3624_
	);
	LUT3 #(
		.INIT('h14)
	) name2275 (
		_w3536_,
		_w3496_,
		_w3532_,
		_w3625_
	);
	LUT4 #(
		.INIT('hcfff)
	) name2276 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3626_
	);
	LUT3 #(
		.INIT('h02)
	) name2277 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w3572_,
		_w3611_,
		_w3627_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2278 (
		_w3440_,
		_w3441_,
		_w3626_,
		_w3627_,
		_w3628_
	);
	LUT3 #(
		.INIT('ha2)
	) name2279 (
		_w1939_,
		_w3628_,
		_w3623_,
		_w3629_
	);
	LUT4 #(
		.INIT('h5700)
	) name2280 (
		_w3623_,
		_w3624_,
		_w3625_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('h2)
	) name2281 (
		_w3407_,
		_w3628_,
		_w3631_
	);
	LUT4 #(
		.INIT('hc055)
	) name2282 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3572_,
		_w3632_
	);
	LUT2 #(
		.INIT('h2)
	) name2283 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		_w3545_,
		_w3633_
	);
	LUT3 #(
		.INIT('h0d)
	) name2284 (
		_w2248_,
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h4)
	) name2285 (
		_w3631_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('hb)
	) name2286 (
		_w3630_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name2287 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3612_,
		_w3637_
	);
	LUT4 #(
		.INIT('ha208)
	) name2288 (
		_w3534_,
		_w3523_,
		_w3526_,
		_w3529_,
		_w3638_
	);
	LUT3 #(
		.INIT('h14)
	) name2289 (
		_w3534_,
		_w3496_,
		_w3532_,
		_w3639_
	);
	LUT3 #(
		.INIT('h02)
	) name2290 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w3572_,
		_w3573_,
		_w3640_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2291 (
		_w3440_,
		_w3441_,
		_w3574_,
		_w3640_,
		_w3641_
	);
	LUT3 #(
		.INIT('ha2)
	) name2292 (
		_w1939_,
		_w3641_,
		_w3637_,
		_w3642_
	);
	LUT4 #(
		.INIT('h5700)
	) name2293 (
		_w3637_,
		_w3638_,
		_w3639_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w3407_,
		_w3641_,
		_w3644_
	);
	LUT4 #(
		.INIT('hc055)
	) name2295 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3573_,
		_w3645_
	);
	LUT2 #(
		.INIT('h2)
	) name2296 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w3545_,
		_w3646_
	);
	LUT3 #(
		.INIT('h0d)
	) name2297 (
		_w2248_,
		_w3645_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h4)
	) name2298 (
		_w3644_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('hb)
	) name2299 (
		_w3643_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3626_,
		_w3650_
	);
	LUT4 #(
		.INIT('hd200)
	) name2301 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3611_,
		_w3651_
	);
	LUT3 #(
		.INIT('h06)
	) name2302 (
		_w3496_,
		_w3532_,
		_w3611_,
		_w3652_
	);
	LUT4 #(
		.INIT('h3fff)
	) name2303 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3653_
	);
	LUT3 #(
		.INIT('h02)
	) name2304 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w3580_,
		_w3573_,
		_w3654_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2305 (
		_w3440_,
		_w3441_,
		_w3653_,
		_w3654_,
		_w3655_
	);
	LUT3 #(
		.INIT('ha2)
	) name2306 (
		_w1939_,
		_w3655_,
		_w3650_,
		_w3656_
	);
	LUT4 #(
		.INIT('h5700)
	) name2307 (
		_w3650_,
		_w3651_,
		_w3652_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h2)
	) name2308 (
		_w3407_,
		_w3655_,
		_w3658_
	);
	LUT4 #(
		.INIT('hc055)
	) name2309 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3580_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w3545_,
		_w3660_
	);
	LUT3 #(
		.INIT('h0d)
	) name2311 (
		_w2248_,
		_w3659_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h4)
	) name2312 (
		_w3658_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('hb)
	) name2313 (
		_w3657_,
		_w3662_,
		_w3663_
	);
	LUT2 #(
		.INIT('h2)
	) name2314 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3653_,
		_w3664_
	);
	LUT4 #(
		.INIT('hd200)
	) name2315 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3573_,
		_w3665_
	);
	LUT3 #(
		.INIT('h06)
	) name2316 (
		_w3496_,
		_w3532_,
		_w3573_,
		_w3666_
	);
	LUT4 #(
		.INIT('h0002)
	) name2317 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3667_
	);
	LUT4 #(
		.INIT('hfffc)
	) name2318 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3668_
	);
	LUT3 #(
		.INIT('h02)
	) name2319 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w3578_,
		_w3667_,
		_w3669_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2320 (
		_w3440_,
		_w3441_,
		_w3668_,
		_w3669_,
		_w3670_
	);
	LUT3 #(
		.INIT('ha2)
	) name2321 (
		_w1939_,
		_w3670_,
		_w3664_,
		_w3671_
	);
	LUT4 #(
		.INIT('h5700)
	) name2322 (
		_w3664_,
		_w3665_,
		_w3666_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h2)
	) name2323 (
		_w3407_,
		_w3670_,
		_w3673_
	);
	LUT4 #(
		.INIT('hc055)
	) name2324 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3667_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w3545_,
		_w3675_
	);
	LUT3 #(
		.INIT('h0d)
	) name2326 (
		_w2248_,
		_w3674_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h4)
	) name2327 (
		_w3673_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('hb)
	) name2328 (
		_w3672_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h2)
	) name2329 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3668_,
		_w3679_
	);
	LUT4 #(
		.INIT('hd200)
	) name2330 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3578_,
		_w3680_
	);
	LUT3 #(
		.INIT('h06)
	) name2331 (
		_w3496_,
		_w3532_,
		_w3578_,
		_w3681_
	);
	LUT4 #(
		.INIT('h0008)
	) name2332 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3682_
	);
	LUT4 #(
		.INIT('h0004)
	) name2333 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3683_
	);
	LUT4 #(
		.INIT('hfff3)
	) name2334 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3684_
	);
	LUT3 #(
		.INIT('h02)
	) name2335 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w3682_,
		_w3683_,
		_w3685_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2336 (
		_w3440_,
		_w3441_,
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT3 #(
		.INIT('ha2)
	) name2337 (
		_w1939_,
		_w3686_,
		_w3679_,
		_w3687_
	);
	LUT4 #(
		.INIT('h5700)
	) name2338 (
		_w3679_,
		_w3680_,
		_w3681_,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name2339 (
		_w3407_,
		_w3686_,
		_w3689_
	);
	LUT4 #(
		.INIT('hc055)
	) name2340 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3682_,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name2341 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w3545_,
		_w3691_
	);
	LUT3 #(
		.INIT('h0d)
	) name2342 (
		_w2248_,
		_w3690_,
		_w3691_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name2343 (
		_w3689_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('hb)
	) name2344 (
		_w3688_,
		_w3693_,
		_w3694_
	);
	LUT2 #(
		.INIT('h2)
	) name2345 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3581_,
		_w3695_
	);
	LUT4 #(
		.INIT('hd200)
	) name2346 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3580_,
		_w3696_
	);
	LUT3 #(
		.INIT('h06)
	) name2347 (
		_w3496_,
		_w3532_,
		_w3580_,
		_w3697_
	);
	LUT4 #(
		.INIT('hfff9)
	) name2348 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3698_
	);
	LUT3 #(
		.INIT('h02)
	) name2349 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w3667_,
		_w3683_,
		_w3699_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2350 (
		_w3440_,
		_w3441_,
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT3 #(
		.INIT('ha2)
	) name2351 (
		_w1939_,
		_w3700_,
		_w3695_,
		_w3701_
	);
	LUT4 #(
		.INIT('h5700)
	) name2352 (
		_w3695_,
		_w3696_,
		_w3697_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		_w3407_,
		_w3700_,
		_w3703_
	);
	LUT4 #(
		.INIT('hc055)
	) name2354 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3683_,
		_w3704_
	);
	LUT2 #(
		.INIT('h2)
	) name2355 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w3545_,
		_w3705_
	);
	LUT3 #(
		.INIT('h0d)
	) name2356 (
		_w2248_,
		_w3704_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h4)
	) name2357 (
		_w3703_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('hb)
	) name2358 (
		_w3702_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h2)
	) name2359 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3698_,
		_w3709_
	);
	LUT4 #(
		.INIT('hd200)
	) name2360 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3667_,
		_w3710_
	);
	LUT3 #(
		.INIT('h06)
	) name2361 (
		_w3496_,
		_w3532_,
		_w3667_,
		_w3711_
	);
	LUT4 #(
		.INIT('h0010)
	) name2362 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3712_
	);
	LUT4 #(
		.INIT('hffe7)
	) name2363 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3713_
	);
	LUT3 #(
		.INIT('h02)
	) name2364 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w3682_,
		_w3712_,
		_w3714_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2365 (
		_w3440_,
		_w3441_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT3 #(
		.INIT('ha2)
	) name2366 (
		_w1939_,
		_w3715_,
		_w3709_,
		_w3716_
	);
	LUT4 #(
		.INIT('h5700)
	) name2367 (
		_w3709_,
		_w3710_,
		_w3711_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name2368 (
		_w3407_,
		_w3715_,
		_w3718_
	);
	LUT4 #(
		.INIT('hc055)
	) name2369 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3712_,
		_w3719_
	);
	LUT2 #(
		.INIT('h2)
	) name2370 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w3545_,
		_w3720_
	);
	LUT3 #(
		.INIT('h0d)
	) name2371 (
		_w2248_,
		_w3719_,
		_w3720_,
		_w3721_
	);
	LUT2 #(
		.INIT('h4)
	) name2372 (
		_w3718_,
		_w3721_,
		_w3722_
	);
	LUT2 #(
		.INIT('hb)
	) name2373 (
		_w3717_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h2)
	) name2374 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3684_,
		_w3724_
	);
	LUT4 #(
		.INIT('hd200)
	) name2375 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3683_,
		_w3725_
	);
	LUT3 #(
		.INIT('h06)
	) name2376 (
		_w3496_,
		_w3532_,
		_w3683_,
		_w3726_
	);
	LUT4 #(
		.INIT('h0020)
	) name2377 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3727_
	);
	LUT4 #(
		.INIT('hffcf)
	) name2378 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3728_
	);
	LUT3 #(
		.INIT('h02)
	) name2379 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w3712_,
		_w3727_,
		_w3729_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2380 (
		_w3440_,
		_w3441_,
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('ha2)
	) name2381 (
		_w1939_,
		_w3730_,
		_w3724_,
		_w3731_
	);
	LUT4 #(
		.INIT('h5700)
	) name2382 (
		_w3724_,
		_w3725_,
		_w3726_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h2)
	) name2383 (
		_w3407_,
		_w3730_,
		_w3733_
	);
	LUT4 #(
		.INIT('hc055)
	) name2384 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3727_,
		_w3734_
	);
	LUT2 #(
		.INIT('h2)
	) name2385 (
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w3545_,
		_w3735_
	);
	LUT3 #(
		.INIT('h0d)
	) name2386 (
		_w2248_,
		_w3734_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h4)
	) name2387 (
		_w3733_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('hb)
	) name2388 (
		_w3732_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name2389 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3713_,
		_w3739_
	);
	LUT4 #(
		.INIT('hd200)
	) name2390 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3682_,
		_w3740_
	);
	LUT3 #(
		.INIT('h06)
	) name2391 (
		_w3496_,
		_w3532_,
		_w3682_,
		_w3741_
	);
	LUT4 #(
		.INIT('h0040)
	) name2392 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3742_
	);
	LUT4 #(
		.INIT('hff9f)
	) name2393 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3743_
	);
	LUT3 #(
		.INIT('h02)
	) name2394 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w3727_,
		_w3742_,
		_w3744_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2395 (
		_w3440_,
		_w3441_,
		_w3743_,
		_w3744_,
		_w3745_
	);
	LUT3 #(
		.INIT('ha2)
	) name2396 (
		_w1939_,
		_w3745_,
		_w3739_,
		_w3746_
	);
	LUT4 #(
		.INIT('h5700)
	) name2397 (
		_w3739_,
		_w3740_,
		_w3741_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h2)
	) name2398 (
		_w3407_,
		_w3745_,
		_w3748_
	);
	LUT4 #(
		.INIT('hc055)
	) name2399 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3742_,
		_w3749_
	);
	LUT2 #(
		.INIT('h2)
	) name2400 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w3545_,
		_w3750_
	);
	LUT3 #(
		.INIT('h0d)
	) name2401 (
		_w2248_,
		_w3749_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h4)
	) name2402 (
		_w3748_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('hb)
	) name2403 (
		_w3747_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name2404 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3728_,
		_w3754_
	);
	LUT4 #(
		.INIT('hd200)
	) name2405 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3712_,
		_w3755_
	);
	LUT3 #(
		.INIT('h06)
	) name2406 (
		_w3496_,
		_w3532_,
		_w3712_,
		_w3756_
	);
	LUT4 #(
		.INIT('hff3f)
	) name2407 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3757_
	);
	LUT3 #(
		.INIT('h02)
	) name2408 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w3592_,
		_w3742_,
		_w3758_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2409 (
		_w3440_,
		_w3441_,
		_w3757_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('ha2)
	) name2410 (
		_w1939_,
		_w3759_,
		_w3754_,
		_w3760_
	);
	LUT4 #(
		.INIT('h5700)
	) name2411 (
		_w3754_,
		_w3755_,
		_w3756_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h2)
	) name2412 (
		_w3407_,
		_w3759_,
		_w3762_
	);
	LUT4 #(
		.INIT('hc055)
	) name2413 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3592_,
		_w3763_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w3545_,
		_w3764_
	);
	LUT3 #(
		.INIT('h0d)
	) name2415 (
		_w2248_,
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h4)
	) name2416 (
		_w3762_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('hb)
	) name2417 (
		_w3761_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h2)
	) name2418 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3743_,
		_w3768_
	);
	LUT4 #(
		.INIT('hd200)
	) name2419 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3727_,
		_w3769_
	);
	LUT3 #(
		.INIT('h06)
	) name2420 (
		_w3496_,
		_w3532_,
		_w3727_,
		_w3770_
	);
	LUT3 #(
		.INIT('h02)
	) name2421 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w3411_,
		_w3592_,
		_w3771_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2422 (
		_w3440_,
		_w3441_,
		_w3593_,
		_w3771_,
		_w3772_
	);
	LUT3 #(
		.INIT('ha2)
	) name2423 (
		_w1939_,
		_w3772_,
		_w3768_,
		_w3773_
	);
	LUT4 #(
		.INIT('h5700)
	) name2424 (
		_w3768_,
		_w3769_,
		_w3770_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h2)
	) name2425 (
		_w3407_,
		_w3772_,
		_w3775_
	);
	LUT4 #(
		.INIT('hc055)
	) name2426 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3411_,
		_w3776_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w3545_,
		_w3777_
	);
	LUT3 #(
		.INIT('h0d)
	) name2428 (
		_w2248_,
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h4)
	) name2429 (
		_w3775_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('hb)
	) name2430 (
		_w3774_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3757_,
		_w3781_
	);
	LUT4 #(
		.INIT('hd200)
	) name2432 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w3742_,
		_w3782_
	);
	LUT3 #(
		.INIT('h06)
	) name2433 (
		_w3496_,
		_w3532_,
		_w3742_,
		_w3783_
	);
	LUT3 #(
		.INIT('h02)
	) name2434 (
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w3411_,
		_w3412_,
		_w3784_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2435 (
		_w3440_,
		_w3441_,
		_w3413_,
		_w3784_,
		_w3785_
	);
	LUT3 #(
		.INIT('ha2)
	) name2436 (
		_w1939_,
		_w3785_,
		_w3781_,
		_w3786_
	);
	LUT4 #(
		.INIT('h5700)
	) name2437 (
		_w3781_,
		_w3782_,
		_w3783_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h2)
	) name2438 (
		_w3407_,
		_w3785_,
		_w3788_
	);
	LUT4 #(
		.INIT('hc055)
	) name2439 (
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1776_,
		_w1781_,
		_w3412_,
		_w3789_
	);
	LUT2 #(
		.INIT('h2)
	) name2440 (
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w3545_,
		_w3790_
	);
	LUT3 #(
		.INIT('h0d)
	) name2441 (
		_w2248_,
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w3788_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('hb)
	) name2443 (
		_w3787_,
		_w3792_,
		_w3793_
	);
	LUT3 #(
		.INIT('ha8)
	) name2444 (
		_w2315_,
		_w3550_,
		_w3551_,
		_w3794_
	);
	LUT3 #(
		.INIT('ha8)
	) name2445 (
		_w2317_,
		_w3554_,
		_w3555_,
		_w3795_
	);
	LUT3 #(
		.INIT('ha8)
	) name2446 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT3 #(
		.INIT('h02)
	) name2447 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w2320_,
		_w2322_,
		_w3797_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2448 (
		_w2323_,
		_w3559_,
		_w3560_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w2327_,
		_w3798_,
		_w3799_
	);
	LUT3 #(
		.INIT('ha8)
	) name2450 (
		_w1679_,
		_w3796_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h2)
	) name2451 (
		_w2283_,
		_w3798_,
		_w3801_
	);
	LUT4 #(
		.INIT('hc055)
	) name2452 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2320_,
		_w3802_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		_w2288_,
		_w3803_
	);
	LUT3 #(
		.INIT('h0d)
	) name2454 (
		_w2246_,
		_w3802_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('h4)
	) name2455 (
		_w3801_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('hb)
	) name2456 (
		_w3800_,
		_w3805_,
		_w3806_
	);
	LUT3 #(
		.INIT('ha8)
	) name2457 (
		_w2250_,
		_w3554_,
		_w3555_,
		_w3807_
	);
	LUT3 #(
		.INIT('ha8)
	) name2458 (
		_w2349_,
		_w3550_,
		_w3551_,
		_w3808_
	);
	LUT3 #(
		.INIT('ha8)
	) name2459 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT3 #(
		.INIT('h02)
	) name2460 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w2271_,
		_w2264_,
		_w3810_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2461 (
		_w2346_,
		_w3559_,
		_w3560_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w2351_,
		_w3811_,
		_w3812_
	);
	LUT3 #(
		.INIT('ha8)
	) name2463 (
		_w1679_,
		_w3809_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		_w2283_,
		_w3811_,
		_w3814_
	);
	LUT4 #(
		.INIT('hc055)
	) name2465 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2271_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		_w2288_,
		_w3816_
	);
	LUT3 #(
		.INIT('h0d)
	) name2467 (
		_w2246_,
		_w3815_,
		_w3816_,
		_w3817_
	);
	LUT2 #(
		.INIT('h4)
	) name2468 (
		_w3814_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('hb)
	) name2469 (
		_w3813_,
		_w3818_,
		_w3819_
	);
	LUT3 #(
		.INIT('ha8)
	) name2470 (
		_w2264_,
		_w3550_,
		_w3551_,
		_w3820_
	);
	LUT3 #(
		.INIT('ha8)
	) name2471 (
		_w2271_,
		_w3554_,
		_w3555_,
		_w3821_
	);
	LUT3 #(
		.INIT('ha8)
	) name2472 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT3 #(
		.INIT('h02)
	) name2473 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w2272_,
		_w2376_,
		_w3823_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2474 (
		_w2377_,
		_w3559_,
		_w3560_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w2380_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('ha8)
	) name2476 (
		_w1679_,
		_w3822_,
		_w3825_,
		_w3826_
	);
	LUT2 #(
		.INIT('h2)
	) name2477 (
		_w2283_,
		_w3824_,
		_w3827_
	);
	LUT4 #(
		.INIT('hc055)
	) name2478 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2376_,
		_w3828_
	);
	LUT2 #(
		.INIT('h2)
	) name2479 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w2288_,
		_w3829_
	);
	LUT3 #(
		.INIT('h0d)
	) name2480 (
		_w2246_,
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w3827_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('hb)
	) name2482 (
		_w3826_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('ha8)
	) name2483 (
		_w2271_,
		_w3550_,
		_w3551_,
		_w3833_
	);
	LUT3 #(
		.INIT('ha8)
	) name2484 (
		_w2272_,
		_w3554_,
		_w3555_,
		_w3834_
	);
	LUT3 #(
		.INIT('ha8)
	) name2485 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT3 #(
		.INIT('h02)
	) name2486 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w2315_,
		_w2376_,
		_w3836_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2487 (
		_w2402_,
		_w3559_,
		_w3560_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name2488 (
		_w2405_,
		_w3837_,
		_w3838_
	);
	LUT3 #(
		.INIT('ha8)
	) name2489 (
		_w1679_,
		_w3835_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h2)
	) name2490 (
		_w2283_,
		_w3837_,
		_w3840_
	);
	LUT4 #(
		.INIT('hc055)
	) name2491 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2315_,
		_w3841_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w2288_,
		_w3842_
	);
	LUT3 #(
		.INIT('h0d)
	) name2493 (
		_w2246_,
		_w3841_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w3840_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('hb)
	) name2495 (
		_w3839_,
		_w3844_,
		_w3845_
	);
	LUT3 #(
		.INIT('ha8)
	) name2496 (
		_w2272_,
		_w3550_,
		_w3551_,
		_w3846_
	);
	LUT3 #(
		.INIT('ha8)
	) name2497 (
		_w2376_,
		_w3554_,
		_w3555_,
		_w3847_
	);
	LUT3 #(
		.INIT('ha8)
	) name2498 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3846_,
		_w3847_,
		_w3848_
	);
	LUT3 #(
		.INIT('h02)
	) name2499 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w2315_,
		_w2317_,
		_w3849_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2500 (
		_w2326_,
		_w3559_,
		_w3560_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('h1)
	) name2501 (
		_w2429_,
		_w3850_,
		_w3851_
	);
	LUT3 #(
		.INIT('ha8)
	) name2502 (
		_w1679_,
		_w3848_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h2)
	) name2503 (
		_w2283_,
		_w3850_,
		_w3853_
	);
	LUT4 #(
		.INIT('hc055)
	) name2504 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2317_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		_w2288_,
		_w3855_
	);
	LUT3 #(
		.INIT('h0d)
	) name2506 (
		_w2246_,
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h4)
	) name2507 (
		_w3853_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('hb)
	) name2508 (
		_w3852_,
		_w3857_,
		_w3858_
	);
	LUT3 #(
		.INIT('ha8)
	) name2509 (
		_w2376_,
		_w3550_,
		_w3551_,
		_w3859_
	);
	LUT3 #(
		.INIT('ha8)
	) name2510 (
		_w2315_,
		_w3554_,
		_w3555_,
		_w3860_
	);
	LUT3 #(
		.INIT('ha8)
	) name2511 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT3 #(
		.INIT('h02)
	) name2512 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w2322_,
		_w2317_,
		_w3862_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2513 (
		_w2451_,
		_w3559_,
		_w3560_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w2454_,
		_w3863_,
		_w3864_
	);
	LUT3 #(
		.INIT('ha8)
	) name2515 (
		_w1679_,
		_w3861_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h2)
	) name2516 (
		_w2283_,
		_w3863_,
		_w3866_
	);
	LUT4 #(
		.INIT('hc055)
	) name2517 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2322_,
		_w3867_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w2288_,
		_w3868_
	);
	LUT3 #(
		.INIT('h0d)
	) name2519 (
		_w2246_,
		_w3867_,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h4)
	) name2520 (
		_w3866_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('hb)
	) name2521 (
		_w3865_,
		_w3870_,
		_w3871_
	);
	LUT3 #(
		.INIT('ha8)
	) name2522 (
		_w2317_,
		_w3550_,
		_w3551_,
		_w3872_
	);
	LUT3 #(
		.INIT('ha8)
	) name2523 (
		_w2322_,
		_w3554_,
		_w3555_,
		_w3873_
	);
	LUT3 #(
		.INIT('ha8)
	) name2524 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3872_,
		_w3873_,
		_w3874_
	);
	LUT3 #(
		.INIT('h02)
	) name2525 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w2320_,
		_w2473_,
		_w3875_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2526 (
		_w2474_,
		_w3559_,
		_w3560_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w2477_,
		_w3876_,
		_w3877_
	);
	LUT3 #(
		.INIT('ha8)
	) name2528 (
		_w1679_,
		_w3874_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		_w2283_,
		_w3876_,
		_w3879_
	);
	LUT4 #(
		.INIT('hc055)
	) name2530 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2473_,
		_w3880_
	);
	LUT2 #(
		.INIT('h2)
	) name2531 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w2288_,
		_w3881_
	);
	LUT3 #(
		.INIT('h0d)
	) name2532 (
		_w2246_,
		_w3880_,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		_w3879_,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('hb)
	) name2534 (
		_w3878_,
		_w3883_,
		_w3884_
	);
	LUT3 #(
		.INIT('ha8)
	) name2535 (
		_w2320_,
		_w3554_,
		_w3555_,
		_w3885_
	);
	LUT3 #(
		.INIT('ha8)
	) name2536 (
		_w2322_,
		_w3550_,
		_w3551_,
		_w3886_
	);
	LUT3 #(
		.INIT('ha8)
	) name2537 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3885_,
		_w3886_,
		_w3887_
	);
	LUT3 #(
		.INIT('h02)
	) name2538 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w2473_,
		_w2502_,
		_w3888_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2539 (
		_w2503_,
		_w3559_,
		_w3560_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w2506_,
		_w3889_,
		_w3890_
	);
	LUT3 #(
		.INIT('ha8)
	) name2541 (
		_w1679_,
		_w3887_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h2)
	) name2542 (
		_w2283_,
		_w3889_,
		_w3892_
	);
	LUT4 #(
		.INIT('hc055)
	) name2543 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2502_,
		_w3893_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w2288_,
		_w3894_
	);
	LUT3 #(
		.INIT('h0d)
	) name2545 (
		_w2246_,
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w3892_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('hb)
	) name2547 (
		_w3891_,
		_w3896_,
		_w3897_
	);
	LUT3 #(
		.INIT('ha8)
	) name2548 (
		_w2320_,
		_w3550_,
		_w3551_,
		_w3898_
	);
	LUT3 #(
		.INIT('ha8)
	) name2549 (
		_w2473_,
		_w3554_,
		_w3555_,
		_w3899_
	);
	LUT3 #(
		.INIT('ha8)
	) name2550 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3898_,
		_w3899_,
		_w3900_
	);
	LUT3 #(
		.INIT('h02)
	) name2551 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w2502_,
		_w2528_,
		_w3901_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2552 (
		_w2529_,
		_w3559_,
		_w3560_,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		_w2532_,
		_w3902_,
		_w3903_
	);
	LUT3 #(
		.INIT('ha8)
	) name2554 (
		_w1679_,
		_w3900_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h2)
	) name2555 (
		_w2283_,
		_w3902_,
		_w3905_
	);
	LUT4 #(
		.INIT('hc055)
	) name2556 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2528_,
		_w3906_
	);
	LUT2 #(
		.INIT('h2)
	) name2557 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w2288_,
		_w3907_
	);
	LUT3 #(
		.INIT('h0d)
	) name2558 (
		_w2246_,
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h4)
	) name2559 (
		_w3905_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('hb)
	) name2560 (
		_w3904_,
		_w3909_,
		_w3910_
	);
	LUT3 #(
		.INIT('ha8)
	) name2561 (
		_w2473_,
		_w3550_,
		_w3551_,
		_w3911_
	);
	LUT3 #(
		.INIT('ha8)
	) name2562 (
		_w2502_,
		_w3554_,
		_w3555_,
		_w3912_
	);
	LUT3 #(
		.INIT('ha8)
	) name2563 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT3 #(
		.INIT('h02)
	) name2564 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w2528_,
		_w2554_,
		_w3914_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2565 (
		_w2555_,
		_w3559_,
		_w3560_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		_w2558_,
		_w3915_,
		_w3916_
	);
	LUT3 #(
		.INIT('ha8)
	) name2567 (
		_w1679_,
		_w3913_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h2)
	) name2568 (
		_w2283_,
		_w3915_,
		_w3918_
	);
	LUT4 #(
		.INIT('hc055)
	) name2569 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2554_,
		_w3919_
	);
	LUT2 #(
		.INIT('h2)
	) name2570 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w2288_,
		_w3920_
	);
	LUT3 #(
		.INIT('h0d)
	) name2571 (
		_w2246_,
		_w3919_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h4)
	) name2572 (
		_w3918_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('hb)
	) name2573 (
		_w3917_,
		_w3922_,
		_w3923_
	);
	LUT3 #(
		.INIT('ha8)
	) name2574 (
		_w2502_,
		_w3550_,
		_w3551_,
		_w3924_
	);
	LUT3 #(
		.INIT('ha8)
	) name2575 (
		_w2528_,
		_w3554_,
		_w3555_,
		_w3925_
	);
	LUT3 #(
		.INIT('ha8)
	) name2576 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3924_,
		_w3925_,
		_w3926_
	);
	LUT3 #(
		.INIT('h02)
	) name2577 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w2554_,
		_w2580_,
		_w3927_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2578 (
		_w2581_,
		_w3559_,
		_w3560_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w2584_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('ha8)
	) name2580 (
		_w1679_,
		_w3926_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		_w2283_,
		_w3928_,
		_w3931_
	);
	LUT4 #(
		.INIT('hc055)
	) name2582 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2580_,
		_w3932_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w2288_,
		_w3933_
	);
	LUT3 #(
		.INIT('h0d)
	) name2584 (
		_w2246_,
		_w3932_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name2585 (
		_w3931_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('hb)
	) name2586 (
		_w3930_,
		_w3935_,
		_w3936_
	);
	LUT3 #(
		.INIT('ha8)
	) name2587 (
		_w2528_,
		_w3550_,
		_w3551_,
		_w3937_
	);
	LUT3 #(
		.INIT('ha8)
	) name2588 (
		_w2554_,
		_w3554_,
		_w3555_,
		_w3938_
	);
	LUT3 #(
		.INIT('ha8)
	) name2589 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3937_,
		_w3938_,
		_w3939_
	);
	LUT3 #(
		.INIT('h02)
	) name2590 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w2580_,
		_w2606_,
		_w3940_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2591 (
		_w2607_,
		_w3559_,
		_w3560_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w2610_,
		_w3941_,
		_w3942_
	);
	LUT3 #(
		.INIT('ha8)
	) name2593 (
		_w1679_,
		_w3939_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		_w2283_,
		_w3941_,
		_w3944_
	);
	LUT4 #(
		.INIT('hc055)
	) name2595 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2606_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w2288_,
		_w3946_
	);
	LUT3 #(
		.INIT('h0d)
	) name2597 (
		_w2246_,
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h4)
	) name2598 (
		_w3944_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('hb)
	) name2599 (
		_w3943_,
		_w3948_,
		_w3949_
	);
	LUT3 #(
		.INIT('ha8)
	) name2600 (
		_w2554_,
		_w3550_,
		_w3551_,
		_w3950_
	);
	LUT3 #(
		.INIT('ha8)
	) name2601 (
		_w2580_,
		_w3554_,
		_w3555_,
		_w3951_
	);
	LUT3 #(
		.INIT('ha8)
	) name2602 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3950_,
		_w3951_,
		_w3952_
	);
	LUT3 #(
		.INIT('h02)
	) name2603 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w2349_,
		_w2606_,
		_w3953_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2604 (
		_w2632_,
		_w3559_,
		_w3560_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w2635_,
		_w3954_,
		_w3955_
	);
	LUT3 #(
		.INIT('ha8)
	) name2606 (
		_w1679_,
		_w3952_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		_w2283_,
		_w3954_,
		_w3957_
	);
	LUT4 #(
		.INIT('hc055)
	) name2608 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2349_,
		_w3958_
	);
	LUT2 #(
		.INIT('h2)
	) name2609 (
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w2288_,
		_w3959_
	);
	LUT3 #(
		.INIT('h0d)
	) name2610 (
		_w2246_,
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h4)
	) name2611 (
		_w3957_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('hb)
	) name2612 (
		_w3956_,
		_w3961_,
		_w3962_
	);
	LUT3 #(
		.INIT('ha8)
	) name2613 (
		_w2580_,
		_w3550_,
		_w3551_,
		_w3963_
	);
	LUT3 #(
		.INIT('ha8)
	) name2614 (
		_w2606_,
		_w3554_,
		_w3555_,
		_w3964_
	);
	LUT3 #(
		.INIT('ha8)
	) name2615 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3963_,
		_w3964_,
		_w3965_
	);
	LUT3 #(
		.INIT('h02)
	) name2616 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w2250_,
		_w2349_,
		_w3966_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2617 (
		_w2350_,
		_w3559_,
		_w3560_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h1)
	) name2618 (
		_w2659_,
		_w3967_,
		_w3968_
	);
	LUT3 #(
		.INIT('ha8)
	) name2619 (
		_w1679_,
		_w3965_,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		_w2283_,
		_w3967_,
		_w3970_
	);
	LUT4 #(
		.INIT('hc055)
	) name2621 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2250_,
		_w3971_
	);
	LUT2 #(
		.INIT('h2)
	) name2622 (
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w2288_,
		_w3972_
	);
	LUT3 #(
		.INIT('h0d)
	) name2623 (
		_w2246_,
		_w3971_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h4)
	) name2624 (
		_w3970_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('hb)
	) name2625 (
		_w3969_,
		_w3974_,
		_w3975_
	);
	LUT3 #(
		.INIT('ha8)
	) name2626 (
		_w2606_,
		_w3550_,
		_w3551_,
		_w3976_
	);
	LUT3 #(
		.INIT('ha8)
	) name2627 (
		_w2349_,
		_w3554_,
		_w3555_,
		_w3977_
	);
	LUT3 #(
		.INIT('ha8)
	) name2628 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w3976_,
		_w3977_,
		_w3978_
	);
	LUT3 #(
		.INIT('h02)
	) name2629 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w2250_,
		_w2264_,
		_w3979_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2630 (
		_w2279_,
		_w3559_,
		_w3560_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w2683_,
		_w3980_,
		_w3981_
	);
	LUT3 #(
		.INIT('ha8)
	) name2632 (
		_w1679_,
		_w3978_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		_w2283_,
		_w3980_,
		_w3983_
	);
	LUT4 #(
		.INIT('hc055)
	) name2634 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1473_,
		_w1478_,
		_w2264_,
		_w3984_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w2288_,
		_w3985_
	);
	LUT3 #(
		.INIT('h0d)
	) name2636 (
		_w2246_,
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h4)
	) name2637 (
		_w3983_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('hb)
	) name2638 (
		_w3982_,
		_w3987_,
		_w3988_
	);
	LUT3 #(
		.INIT('h08)
	) name2639 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w1842_,
		_w1915_,
		_w3989_
	);
	LUT3 #(
		.INIT('h6c)
	) name2640 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3080_,
		_w3990_
	);
	LUT2 #(
		.INIT('h6)
	) name2641 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3072_,
		_w3991_
	);
	LUT3 #(
		.INIT('h28)
	) name2642 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3088_,
		_w3992_
	);
	LUT4 #(
		.INIT('h0200)
	) name2643 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3068_,
		_w3299_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		_w3071_,
		_w3302_,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		_w3993_,
		_w3994_,
		_w3995_
	);
	LUT4 #(
		.INIT('h8000)
	) name2646 (
		_w3296_,
		_w3307_,
		_w3991_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3308_,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		_w3319_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('h8222)
	) name2649 (
		_w3101_,
		_w3990_,
		_w3996_,
		_w3998_,
		_w3999_
	);
	LUT4 #(
		.INIT('h00dc)
	) name2650 (
		_w3157_,
		_w3156_,
		_w3169_,
		_w3200_,
		_w4000_
	);
	LUT3 #(
		.INIT('h01)
	) name2651 (
		_w3143_,
		_w3182_,
		_w3197_,
		_w4001_
	);
	LUT3 #(
		.INIT('h0b)
	) name2652 (
		_w3143_,
		_w3199_,
		_w3204_,
		_w4002_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2653 (
		_w3131_,
		_w4000_,
		_w4001_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('h008f)
	) name2654 (
		_w3095_,
		_w3100_,
		_w3102_,
		_w3210_,
		_w4004_
	);
	LUT3 #(
		.INIT('h0b)
	) name2655 (
		_w3129_,
		_w3205_,
		_w3208_,
		_w4005_
	);
	LUT4 #(
		.INIT('h3110)
	) name2656 (
		_w3127_,
		_w3103_,
		_w3128_,
		_w3205_,
		_w4006_
	);
	LUT2 #(
		.INIT('h2)
	) name2657 (
		_w4004_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('hc301)
	) name2658 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3086_,
		_w3089_,
		_w4008_
	);
	LUT3 #(
		.INIT('h10)
	) name2659 (
		_w3216_,
		_w3221_,
		_w4008_,
		_w4009_
	);
	LUT3 #(
		.INIT('h40)
	) name2660 (
		_w4003_,
		_w4007_,
		_w4009_,
		_w4010_
	);
	LUT4 #(
		.INIT('h1000)
	) name2661 (
		_w3219_,
		_w4003_,
		_w4007_,
		_w4009_,
		_w4011_
	);
	LUT3 #(
		.INIT('h80)
	) name2662 (
		_w3256_,
		_w3262_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h4554)
	) name2663 (
		_w1916_,
		_w3101_,
		_w3263_,
		_w4012_,
		_w4013_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2664 (
		_w1810_,
		_w3989_,
		_w3999_,
		_w4013_,
		_w4014_
	);
	LUT3 #(
		.INIT('h6c)
	) name2665 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w3387_,
		_w4015_
	);
	LUT3 #(
		.INIT('h6a)
	) name2666 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3074_,
		_w3366_,
		_w4016_
	);
	LUT4 #(
		.INIT('h4888)
	) name2667 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3074_,
		_w3366_,
		_w4017_
	);
	LUT4 #(
		.INIT('h002b)
	) name2668 (
		_w3154_,
		_w3155_,
		_w3337_,
		_w3340_,
		_w4018_
	);
	LUT2 #(
		.INIT('h1)
	) name2669 (
		_w3339_,
		_w3345_,
		_w4019_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2670 (
		_w3331_,
		_w3335_,
		_w4018_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w3344_,
		_w3354_,
		_w4021_
	);
	LUT3 #(
		.INIT('h45)
	) name2672 (
		_w3351_,
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT4 #(
		.INIT('h2322)
	) name2673 (
		_w3351_,
		_w3353_,
		_w4020_,
		_w4021_,
		_w4023_
	);
	LUT4 #(
		.INIT('hf070)
	) name2674 (
		_w3095_,
		_w3100_,
		_w3358_,
		_w3348_,
		_w4024_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		_w3065_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h6)
	) name2676 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w3367_,
		_w4026_
	);
	LUT3 #(
		.INIT('h80)
	) name2677 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3060_,
		_w3362_,
		_w4027_
	);
	LUT3 #(
		.INIT('h60)
	) name2678 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w3367_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h8)
	) name2679 (
		_w3074_,
		_w3368_,
		_w4029_
	);
	LUT4 #(
		.INIT('h4000)
	) name2680 (
		_w4023_,
		_w4025_,
		_w4028_,
		_w4029_,
		_w4030_
	);
	LUT4 #(
		.INIT('h4080)
	) name2681 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w3379_,
		_w4031_
	);
	LUT2 #(
		.INIT('h6)
	) name2682 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3387_,
		_w4032_
	);
	LUT3 #(
		.INIT('h60)
	) name2683 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3387_,
		_w4031_,
		_w4033_
	);
	LUT4 #(
		.INIT('h8000)
	) name2684 (
		_w3383_,
		_w4017_,
		_w4030_,
		_w4033_,
		_w4034_
	);
	LUT2 #(
		.INIT('h8)
	) name2685 (
		_w1847_,
		_w4015_,
		_w4035_
	);
	LUT3 #(
		.INIT('hb0)
	) name2686 (
		_w1816_,
		_w1831_,
		_w3263_,
		_w4036_
	);
	LUT4 #(
		.INIT('h0001)
	) name2687 (
		_w1877_,
		_w1913_,
		_w1863_,
		_w1864_,
		_w4037_
	);
	LUT3 #(
		.INIT('h2a)
	) name2688 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		_w1922_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h4)
	) name2689 (
		_w1862_,
		_w3990_,
		_w4039_
	);
	LUT4 #(
		.INIT('h0001)
	) name2690 (
		_w4036_,
		_w4038_,
		_w4039_,
		_w4035_,
		_w4040_
	);
	LUT4 #(
		.INIT('hd700)
	) name2691 (
		_w1924_,
		_w4015_,
		_w4034_,
		_w4040_,
		_w4041_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2692 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w3406_,
		_w3408_,
		_w4042_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2693 (
		_w1933_,
		_w4014_,
		_w4041_,
		_w4042_,
		_w4043_
	);
	LUT3 #(
		.INIT('h02)
	) name2694 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2103_,
		_w2172_,
		_w4044_
	);
	LUT3 #(
		.INIT('h32)
	) name2695 (
		_w2918_,
		_w2923_,
		_w2928_,
		_w4045_
	);
	LUT2 #(
		.INIT('h1)
	) name2696 (
		_w2931_,
		_w2921_,
		_w4046_
	);
	LUT4 #(
		.INIT('hf400)
	) name2697 (
		_w2796_,
		_w2925_,
		_w4045_,
		_w4046_,
		_w4047_
	);
	LUT3 #(
		.INIT('h0b)
	) name2698 (
		_w2931_,
		_w2927_,
		_w2939_,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w2933_,
		_w2947_,
		_w4049_
	);
	LUT3 #(
		.INIT('h0e)
	) name2700 (
		_w2937_,
		_w2938_,
		_w2947_,
		_w4050_
	);
	LUT4 #(
		.INIT('h004f)
	) name2701 (
		_w4047_,
		_w4048_,
		_w4049_,
		_w4050_,
		_w4051_
	);
	LUT3 #(
		.INIT('h6a)
	) name2702 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2715_,
		_w2716_,
		_w4052_
	);
	LUT4 #(
		.INIT('h4888)
	) name2703 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2715_,
		_w2716_,
		_w4053_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w2945_,
		_w4053_,
		_w4054_
	);
	LUT3 #(
		.INIT('h60)
	) name2705 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2893_,
		_w2949_,
		_w4055_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		_w2943_,
		_w4055_,
		_w4056_
	);
	LUT4 #(
		.INIT('h8000)
	) name2707 (
		_w2708_,
		_w2943_,
		_w2956_,
		_w4055_,
		_w4057_
	);
	LUT3 #(
		.INIT('h40)
	) name2708 (
		_w4051_,
		_w4054_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w2966_,
		_w2971_,
		_w4059_
	);
	LUT4 #(
		.INIT('h4000)
	) name2710 (
		_w4051_,
		_w4054_,
		_w4057_,
		_w4059_,
		_w4060_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2711 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2712_,
		_w2720_,
		_w4061_
	);
	LUT3 #(
		.INIT('h80)
	) name2712 (
		_w2969_,
		_w2970_,
		_w2975_,
		_w4062_
	);
	LUT3 #(
		.INIT('h80)
	) name2713 (
		_w4060_,
		_w4061_,
		_w4062_,
		_w4063_
	);
	LUT3 #(
		.INIT('h6c)
	) name2714 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2724_,
		_w4064_
	);
	LUT3 #(
		.INIT('h01)
	) name2715 (
		_w2881_,
		_w2883_,
		_w2891_,
		_w4065_
	);
	LUT3 #(
		.INIT('h0e)
	) name2716 (
		_w2868_,
		_w2870_,
		_w2864_,
		_w4066_
	);
	LUT4 #(
		.INIT('h0032)
	) name2717 (
		_w2868_,
		_w2869_,
		_w2870_,
		_w2864_,
		_w4067_
	);
	LUT3 #(
		.INIT('h10)
	) name2718 (
		_w2876_,
		_w2878_,
		_w4067_,
		_w4068_
	);
	LUT3 #(
		.INIT('h0d)
	) name2719 (
		_w2772_,
		_w2812_,
		_w2829_,
		_w4069_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w2857_,
		_w2826_,
		_w4070_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2721 (
		_w2797_,
		_w2813_,
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT3 #(
		.INIT('h0b)
	) name2722 (
		_w2857_,
		_w2828_,
		_w2861_,
		_w4072_
	);
	LUT3 #(
		.INIT('h23)
	) name2723 (
		_w2758_,
		_w2863_,
		_w2860_,
		_w4073_
	);
	LUT4 #(
		.INIT('h7500)
	) name2724 (
		_w2859_,
		_w4071_,
		_w4072_,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('h8103)
	) name2725 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2894_,
		_w4075_
	);
	LUT3 #(
		.INIT('h40)
	) name2726 (
		_w2728_,
		_w2890_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('h80)
	) name2727 (
		_w2902_,
		_w2912_,
		_w4076_,
		_w4077_
	);
	LUT4 #(
		.INIT('h8000)
	) name2728 (
		_w4065_,
		_w4068_,
		_w4074_,
		_w4077_,
		_w4078_
	);
	LUT4 #(
		.INIT('h4554)
	) name2729 (
		_w2173_,
		_w2755_,
		_w2729_,
		_w4078_,
		_w4079_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2730 (
		_w2755_,
		_w4063_,
		_w4064_,
		_w4079_,
		_w4080_
	);
	LUT3 #(
		.INIT('ha8)
	) name2731 (
		_w2171_,
		_w4044_,
		_w4080_,
		_w4081_
	);
	LUT3 #(
		.INIT('h80)
	) name2732 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2703_,
		_w3038_,
		_w4082_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2733 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w3038_,
		_w4083_
	);
	LUT4 #(
		.INIT('haa20)
	) name2734 (
		_w3000_,
		_w3006_,
		_w3010_,
		_w3011_,
		_w4084_
	);
	LUT3 #(
		.INIT('h0b)
	) name2735 (
		_w2999_,
		_w3012_,
		_w3016_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w2995_,
		_w3019_,
		_w4086_
	);
	LUT3 #(
		.INIT('h51)
	) name2737 (
		_w2993_,
		_w3015_,
		_w3019_,
		_w4087_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2738 (
		_w4084_,
		_w4085_,
		_w4086_,
		_w4087_,
		_w4088_
	);
	LUT4 #(
		.INIT('h0080)
	) name2739 (
		_w2991_,
		_w3024_,
		_w3028_,
		_w4088_,
		_w4089_
	);
	LUT4 #(
		.INIT('h8000)
	) name2740 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3036_,
		_w3039_,
		_w4089_,
		_w4090_
	);
	LUT3 #(
		.INIT('h13)
	) name2741 (
		_w3042_,
		_w4083_,
		_w4090_,
		_w4091_
	);
	LUT3 #(
		.INIT('h2a)
	) name2742 (
		_w2181_,
		_w3043_,
		_w4090_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2098_,
		_w4093_
	);
	LUT4 #(
		.INIT('h00e0)
	) name2744 (
		_w2071_,
		_w2087_,
		_w4083_,
		_w4093_,
		_w4094_
	);
	LUT3 #(
		.INIT('h0e)
	) name2745 (
		_w2044_,
		_w2047_,
		_w2119_,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w2177_,
		_w4095_,
		_w4096_
	);
	LUT3 #(
		.INIT('h2a)
	) name2747 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		_w2176_,
		_w4096_,
		_w4097_
	);
	LUT3 #(
		.INIT('hb0)
	) name2748 (
		_w2073_,
		_w2086_,
		_w2729_,
		_w4098_
	);
	LUT2 #(
		.INIT('h4)
	) name2749 (
		_w2117_,
		_w4064_,
		_w4099_
	);
	LUT4 #(
		.INIT('h0001)
	) name2750 (
		_w4098_,
		_w4094_,
		_w4099_,
		_w4097_,
		_w4100_
	);
	LUT3 #(
		.INIT('hb0)
	) name2751 (
		_w4091_,
		_w4092_,
		_w4100_,
		_w4101_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2752 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w3054_,
		_w3056_,
		_w4102_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2753 (
		_w1945_,
		_w4081_,
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT3 #(
		.INIT('h08)
	) name2754 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w1592_,
		_w1660_,
		_w4104_
	);
	LUT4 #(
		.INIT('h153f)
	) name2755 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1466_,
		_w1457_,
		_w4105_
	);
	LUT4 #(
		.INIT('h135f)
	) name2756 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1447_,
		_w1462_,
		_w4106_
	);
	LUT4 #(
		.INIT('h153f)
	) name2757 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1450_,
		_w1453_,
		_w4107_
	);
	LUT4 #(
		.INIT('h135f)
	) name2758 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1446_,
		_w1465_,
		_w4108_
	);
	LUT4 #(
		.INIT('h8000)
	) name2759 (
		_w4107_,
		_w4108_,
		_w4105_,
		_w4106_,
		_w4109_
	);
	LUT4 #(
		.INIT('h135f)
	) name2760 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1452_,
		_w1463_,
		_w4110_
	);
	LUT4 #(
		.INIT('h135f)
	) name2761 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1443_,
		_w1456_,
		_w4111_
	);
	LUT4 #(
		.INIT('h135f)
	) name2762 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1449_,
		_w1444_,
		_w4112_
	);
	LUT4 #(
		.INIT('h135f)
	) name2763 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1459_,
		_w1460_,
		_w4113_
	);
	LUT4 #(
		.INIT('h8000)
	) name2764 (
		_w4112_,
		_w4113_,
		_w4110_,
		_w4111_,
		_w4114_
	);
	LUT2 #(
		.INIT('h6)
	) name2765 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4115_
	);
	LUT3 #(
		.INIT('h70)
	) name2766 (
		_w4109_,
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h135f)
	) name2767 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1446_,
		_w1466_,
		_w4117_
	);
	LUT4 #(
		.INIT('h135f)
	) name2768 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1452_,
		_w1463_,
		_w4118_
	);
	LUT4 #(
		.INIT('h153f)
	) name2769 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1465_,
		_w1457_,
		_w4119_
	);
	LUT4 #(
		.INIT('h135f)
	) name2770 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1453_,
		_w1456_,
		_w4120_
	);
	LUT4 #(
		.INIT('h8000)
	) name2771 (
		_w4119_,
		_w4120_,
		_w4117_,
		_w4118_,
		_w4121_
	);
	LUT4 #(
		.INIT('h153f)
	) name2772 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1462_,
		_w1459_,
		_w4122_
	);
	LUT4 #(
		.INIT('h135f)
	) name2773 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1443_,
		_w1460_,
		_w4123_
	);
	LUT4 #(
		.INIT('h153f)
	) name2774 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1450_,
		_w1447_,
		_w4124_
	);
	LUT4 #(
		.INIT('h135f)
	) name2775 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1449_,
		_w1444_,
		_w4125_
	);
	LUT4 #(
		.INIT('h8000)
	) name2776 (
		_w4124_,
		_w4125_,
		_w4122_,
		_w4123_,
		_w4126_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		_w4121_,
		_w4126_,
		_w4127_
	);
	LUT3 #(
		.INIT('h15)
	) name2778 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4121_,
		_w4126_,
		_w4128_
	);
	LUT4 #(
		.INIT('h153f)
	) name2779 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w1446_,
		_w1460_,
		_w4129_
	);
	LUT4 #(
		.INIT('h153f)
	) name2780 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1462_,
		_w1459_,
		_w4130_
	);
	LUT4 #(
		.INIT('h153f)
	) name2781 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1449_,
		_w1466_,
		_w4131_
	);
	LUT4 #(
		.INIT('h135f)
	) name2782 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1443_,
		_w1463_,
		_w4132_
	);
	LUT4 #(
		.INIT('h8000)
	) name2783 (
		_w4131_,
		_w4132_,
		_w4129_,
		_w4130_,
		_w4133_
	);
	LUT4 #(
		.INIT('h135f)
	) name2784 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1447_,
		_w1456_,
		_w4134_
	);
	LUT4 #(
		.INIT('h153f)
	) name2785 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1465_,
		_w1457_,
		_w4135_
	);
	LUT4 #(
		.INIT('h135f)
	) name2786 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1453_,
		_w1444_,
		_w4136_
	);
	LUT4 #(
		.INIT('h153f)
	) name2787 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1450_,
		_w1452_,
		_w4137_
	);
	LUT4 #(
		.INIT('h8000)
	) name2788 (
		_w4136_,
		_w4137_,
		_w4134_,
		_w4135_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		_w4133_,
		_w4138_,
		_w4139_
	);
	LUT3 #(
		.INIT('h2a)
	) name2790 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4133_,
		_w4138_,
		_w4140_
	);
	LUT3 #(
		.INIT('h8e)
	) name2791 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4127_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h080e)
	) name2792 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4127_,
		_w4116_,
		_w4140_,
		_w4142_
	);
	LUT4 #(
		.INIT('h135f)
	) name2793 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[13][4]/NET0131 ,
		_w1443_,
		_w1447_,
		_w4143_
	);
	LUT4 #(
		.INIT('h135f)
	) name2794 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1462_,
		_w1465_,
		_w4144_
	);
	LUT4 #(
		.INIT('h153f)
	) name2795 (
		\P2_InstQueue_reg[5][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1449_,
		_w1466_,
		_w4145_
	);
	LUT4 #(
		.INIT('h135f)
	) name2796 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[12][4]/NET0131 ,
		_w1453_,
		_w1459_,
		_w4146_
	);
	LUT4 #(
		.INIT('h8000)
	) name2797 (
		_w4145_,
		_w4146_,
		_w4143_,
		_w4144_,
		_w4147_
	);
	LUT4 #(
		.INIT('h135f)
	) name2798 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1463_,
		_w1456_,
		_w4148_
	);
	LUT4 #(
		.INIT('h135f)
	) name2799 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1452_,
		_w1446_,
		_w4149_
	);
	LUT4 #(
		.INIT('h153f)
	) name2800 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1450_,
		_w1460_,
		_w4150_
	);
	LUT4 #(
		.INIT('h153f)
	) name2801 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1444_,
		_w1457_,
		_w4151_
	);
	LUT4 #(
		.INIT('h8000)
	) name2802 (
		_w4150_,
		_w4151_,
		_w4148_,
		_w4149_,
		_w4152_
	);
	LUT4 #(
		.INIT('h8000)
	) name2803 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4153_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2804 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4154_
	);
	LUT3 #(
		.INIT('h08)
	) name2805 (
		_w4147_,
		_w4152_,
		_w4154_,
		_w4155_
	);
	LUT4 #(
		.INIT('h135f)
	) name2806 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[12][3]/NET0131 ,
		_w1452_,
		_w1459_,
		_w4156_
	);
	LUT4 #(
		.INIT('h135f)
	) name2807 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w1443_,
		_w1447_,
		_w4157_
	);
	LUT4 #(
		.INIT('h135f)
	) name2808 (
		\P2_InstQueue_reg[4][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1450_,
		_w1465_,
		_w4158_
	);
	LUT4 #(
		.INIT('h153f)
	) name2809 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1463_,
		_w1460_,
		_w4159_
	);
	LUT4 #(
		.INIT('h8000)
	) name2810 (
		_w4158_,
		_w4159_,
		_w4156_,
		_w4157_,
		_w4160_
	);
	LUT4 #(
		.INIT('h153f)
	) name2811 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1449_,
		_w1457_,
		_w4161_
	);
	LUT4 #(
		.INIT('h135f)
	) name2812 (
		\P2_InstQueue_reg[5][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1466_,
		_w1456_,
		_w4162_
	);
	LUT4 #(
		.INIT('h135f)
	) name2813 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1453_,
		_w1444_,
		_w4163_
	);
	LUT4 #(
		.INIT('h135f)
	) name2814 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1446_,
		_w1462_,
		_w4164_
	);
	LUT4 #(
		.INIT('h8000)
	) name2815 (
		_w4163_,
		_w4164_,
		_w4161_,
		_w4162_,
		_w4165_
	);
	LUT3 #(
		.INIT('h78)
	) name2816 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4166_
	);
	LUT3 #(
		.INIT('h08)
	) name2817 (
		_w4160_,
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT3 #(
		.INIT('h08)
	) name2818 (
		_w4109_,
		_w4114_,
		_w4115_,
		_w4168_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT3 #(
		.INIT('h01)
	) name2820 (
		_w4155_,
		_w4167_,
		_w4168_,
		_w4170_
	);
	LUT3 #(
		.INIT('h70)
	) name2821 (
		_w4147_,
		_w4152_,
		_w4154_,
		_w4171_
	);
	LUT3 #(
		.INIT('h70)
	) name2822 (
		_w4160_,
		_w4165_,
		_w4166_,
		_w4172_
	);
	LUT3 #(
		.INIT('h23)
	) name2823 (
		_w4155_,
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('h153f)
	) name2824 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1449_,
		_w1459_,
		_w4174_
	);
	LUT4 #(
		.INIT('h135f)
	) name2825 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1462_,
		_w1456_,
		_w4175_
	);
	LUT4 #(
		.INIT('h135f)
	) name2826 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1453_,
		_w1466_,
		_w4176_
	);
	LUT4 #(
		.INIT('h135f)
	) name2827 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1443_,
		_w1465_,
		_w4177_
	);
	LUT4 #(
		.INIT('h8000)
	) name2828 (
		_w4176_,
		_w4177_,
		_w4174_,
		_w4175_,
		_w4178_
	);
	LUT4 #(
		.INIT('h153f)
	) name2829 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1457_,
		_w1460_,
		_w4179_
	);
	LUT4 #(
		.INIT('h135f)
	) name2830 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1452_,
		_w1463_,
		_w4180_
	);
	LUT4 #(
		.INIT('h153f)
	) name2831 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1450_,
		_w1446_,
		_w4181_
	);
	LUT4 #(
		.INIT('h153f)
	) name2832 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1444_,
		_w1447_,
		_w4182_
	);
	LUT4 #(
		.INIT('h8000)
	) name2833 (
		_w4181_,
		_w4182_,
		_w4179_,
		_w4180_,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		_w4178_,
		_w4183_,
		_w4184_
	);
	LUT3 #(
		.INIT('h80)
	) name2835 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4153_,
		_w4185_
	);
	LUT3 #(
		.INIT('h6c)
	) name2836 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4153_,
		_w4186_
	);
	LUT3 #(
		.INIT('h08)
	) name2837 (
		_w4178_,
		_w4183_,
		_w4186_,
		_w4187_
	);
	LUT4 #(
		.INIT('h135f)
	) name2838 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1447_,
		_w1463_,
		_w4188_
	);
	LUT4 #(
		.INIT('h135f)
	) name2839 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1453_,
		_w1446_,
		_w4189_
	);
	LUT4 #(
		.INIT('h135f)
	) name2840 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1443_,
		_w1456_,
		_w4190_
	);
	LUT4 #(
		.INIT('h153f)
	) name2841 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1465_,
		_w1459_,
		_w4191_
	);
	LUT4 #(
		.INIT('h8000)
	) name2842 (
		_w4190_,
		_w4191_,
		_w4188_,
		_w4189_,
		_w4192_
	);
	LUT4 #(
		.INIT('h135f)
	) name2843 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1452_,
		_w1457_,
		_w4193_
	);
	LUT4 #(
		.INIT('h153f)
	) name2844 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1466_,
		_w1460_,
		_w4194_
	);
	LUT4 #(
		.INIT('h135f)
	) name2845 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1449_,
		_w1444_,
		_w4195_
	);
	LUT4 #(
		.INIT('h153f)
	) name2846 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1450_,
		_w1462_,
		_w4196_
	);
	LUT4 #(
		.INIT('h8000)
	) name2847 (
		_w4195_,
		_w4196_,
		_w4193_,
		_w4194_,
		_w4197_
	);
	LUT2 #(
		.INIT('h6)
	) name2848 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4153_,
		_w4198_
	);
	LUT3 #(
		.INIT('h08)
	) name2849 (
		_w4192_,
		_w4197_,
		_w4198_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name2850 (
		_w4187_,
		_w4199_,
		_w4200_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2851 (
		_w4142_,
		_w4170_,
		_w4173_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('h153f)
	) name2852 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1462_,
		_w1459_,
		_w4202_
	);
	LUT4 #(
		.INIT('h135f)
	) name2853 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1449_,
		_w1456_,
		_w4203_
	);
	LUT4 #(
		.INIT('h153f)
	) name2854 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1465_,
		_w1460_,
		_w4204_
	);
	LUT4 #(
		.INIT('h153f)
	) name2855 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[10][7]/NET0131 ,
		_w1452_,
		_w1453_,
		_w4205_
	);
	LUT4 #(
		.INIT('h8000)
	) name2856 (
		_w4204_,
		_w4205_,
		_w4202_,
		_w4203_,
		_w4206_
	);
	LUT4 #(
		.INIT('h1000)
	) name2857 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		_w1622_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1450_,
		_w4209_
	);
	LUT4 #(
		.INIT('h153f)
	) name2860 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w1446_,
		_w1447_,
		_w4210_
	);
	LUT4 #(
		.INIT('h135f)
	) name2861 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1443_,
		_w1444_,
		_w4211_
	);
	LUT4 #(
		.INIT('h153f)
	) name2862 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1463_,
		_w1457_,
		_w4212_
	);
	LUT4 #(
		.INIT('h4000)
	) name2863 (
		_w4209_,
		_w4211_,
		_w4212_,
		_w4210_,
		_w4213_
	);
	LUT3 #(
		.INIT('h40)
	) name2864 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4214_
	);
	LUT4 #(
		.INIT('h8000)
	) name2865 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4153_,
		_w4215_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2866 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4153_,
		_w4216_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2867 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4216_,
		_w4217_
	);
	LUT3 #(
		.INIT('h70)
	) name2868 (
		_w4178_,
		_w4183_,
		_w4186_,
		_w4218_
	);
	LUT3 #(
		.INIT('h70)
	) name2869 (
		_w4192_,
		_w4197_,
		_w4198_,
		_w4219_
	);
	LUT3 #(
		.INIT('h23)
	) name2870 (
		_w4187_,
		_w4218_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h020b)
	) name2871 (
		_w4184_,
		_w4186_,
		_w4217_,
		_w4219_,
		_w4221_
	);
	LUT4 #(
		.INIT('h0040)
	) name2872 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4216_,
		_w4222_
	);
	LUT2 #(
		.INIT('h6)
	) name2873 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4215_,
		_w4223_
	);
	LUT2 #(
		.INIT('h4)
	) name2874 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4225_
	);
	LUT3 #(
		.INIT('h80)
	) name2876 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4226_
	);
	LUT4 #(
		.INIT('h8000)
	) name2877 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4153_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2878 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4185_,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT3 #(
		.INIT('h80)
	) name2880 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4225_,
		_w4228_,
		_w4230_
	);
	LUT4 #(
		.INIT('hb000)
	) name2881 (
		_w4201_,
		_w4221_,
		_w4224_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w4225_,
		_w4227_,
		_w4232_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4233_
	);
	LUT3 #(
		.INIT('h80)
	) name2884 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4234_
	);
	LUT3 #(
		.INIT('h80)
	) name2885 (
		_w4225_,
		_w4227_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4236_
	);
	LUT3 #(
		.INIT('h80)
	) name2887 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4215_,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4238_
	);
	LUT4 #(
		.INIT('h8000)
	) name2889 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4215_,
		_w4238_,
		_w4239_
	);
	LUT4 #(
		.INIT('h00ec)
	) name2890 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4239_,
		_w4235_,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h6)
	) name2892 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4239_,
		_w4242_
	);
	LUT3 #(
		.INIT('h48)
	) name2893 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4239_,
		_w4243_
	);
	LUT3 #(
		.INIT('h80)
	) name2894 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4240_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w4234_,
		_w4245_,
		_w4246_
	);
	LUT3 #(
		.INIT('h80)
	) name2897 (
		_w4225_,
		_w4227_,
		_w4246_,
		_w4247_
	);
	LUT4 #(
		.INIT('h8000)
	) name2898 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4225_,
		_w4227_,
		_w4246_,
		_w4248_
	);
	LUT2 #(
		.INIT('h6)
	) name2899 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4248_,
		_w4249_
	);
	LUT3 #(
		.INIT('h48)
	) name2900 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4248_,
		_w4250_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2901 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4225_,
		_w4227_,
		_w4246_,
		_w4251_
	);
	LUT3 #(
		.INIT('h80)
	) name2902 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h8000)
	) name2905 (
		_w4225_,
		_w4227_,
		_w4234_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h6)
	) name2906 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4255_,
		_w4256_
	);
	LUT3 #(
		.INIT('h60)
	) name2907 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4255_,
		_w4251_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		_w4250_,
		_w4257_,
		_w4258_
	);
	LUT3 #(
		.INIT('h80)
	) name2909 (
		_w4231_,
		_w4244_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4260_
	);
	LUT3 #(
		.INIT('h6c)
	) name2911 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4255_,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4262_
	);
	LUT3 #(
		.INIT('h80)
	) name2913 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4263_
	);
	LUT3 #(
		.INIT('h6a)
	) name2914 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4255_,
		_w4260_,
		_w4264_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2915 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4255_,
		_w4260_,
		_w4262_,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		_w4261_,
		_w4265_,
		_w4266_
	);
	LUT4 #(
		.INIT('h8000)
	) name2917 (
		_w4231_,
		_w4244_,
		_w4258_,
		_w4266_,
		_w4267_
	);
	LUT3 #(
		.INIT('h80)
	) name2918 (
		_w4255_,
		_w4263_,
		_w4262_,
		_w4268_
	);
	LUT4 #(
		.INIT('h8000)
	) name2919 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4262_,
		_w4269_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2920 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4262_,
		_w4270_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h8)
	) name2922 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4272_
	);
	LUT2 #(
		.INIT('h8)
	) name2923 (
		_w4269_,
		_w4272_,
		_w4273_
	);
	LUT3 #(
		.INIT('h6c)
	) name2924 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4269_,
		_w4274_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2925 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name2926 (
		_w4271_,
		_w4275_,
		_w4276_
	);
	LUT3 #(
		.INIT('h80)
	) name2927 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4272_,
		_w4277_
	);
	LUT4 #(
		.INIT('h8000)
	) name2928 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4269_,
		_w4272_,
		_w4278_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2929 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4269_,
		_w4272_,
		_w4279_
	);
	LUT4 #(
		.INIT('h802a)
	) name2930 (
		_w4214_,
		_w4267_,
		_w4276_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('h8000)
	) name2931 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4281_
	);
	LUT4 #(
		.INIT('h8000)
	) name2932 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h6)
	) name2933 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('h0040)
	) name2934 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4283_,
		_w4284_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2935 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4281_,
		_w4285_
	);
	LUT3 #(
		.INIT('h40)
	) name2936 (
		_w4285_,
		_w4178_,
		_w4183_,
		_w4286_
	);
	LUT3 #(
		.INIT('h6c)
	) name2937 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4281_,
		_w4287_
	);
	LUT3 #(
		.INIT('h40)
	) name2938 (
		_w4287_,
		_w4192_,
		_w4197_,
		_w4288_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		_w4286_,
		_w4288_,
		_w4289_
	);
	LUT3 #(
		.INIT('h01)
	) name2940 (
		_w4284_,
		_w4286_,
		_w4288_,
		_w4290_
	);
	LUT3 #(
		.INIT('h78)
	) name2941 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w4291_
	);
	LUT3 #(
		.INIT('h70)
	) name2942 (
		_w4109_,
		_w4114_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h6)
	) name2943 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4293_
	);
	LUT3 #(
		.INIT('h08)
	) name2944 (
		_w4121_,
		_w4126_,
		_w4293_,
		_w4294_
	);
	LUT3 #(
		.INIT('h80)
	) name2945 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4133_,
		_w4138_,
		_w4295_
	);
	LUT3 #(
		.INIT('h45)
	) name2946 (
		_w4294_,
		_w4128_,
		_w4295_,
		_w4296_
	);
	LUT4 #(
		.INIT('h4544)
	) name2947 (
		_w4292_,
		_w4294_,
		_w4128_,
		_w4295_,
		_w4297_
	);
	LUT2 #(
		.INIT('h6)
	) name2948 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4281_,
		_w4298_
	);
	LUT3 #(
		.INIT('h40)
	) name2949 (
		_w4298_,
		_w4147_,
		_w4152_,
		_w4299_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2950 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4300_
	);
	LUT3 #(
		.INIT('h08)
	) name2951 (
		_w4160_,
		_w4165_,
		_w4300_,
		_w4301_
	);
	LUT3 #(
		.INIT('h08)
	) name2952 (
		_w4109_,
		_w4114_,
		_w4291_,
		_w4302_
	);
	LUT2 #(
		.INIT('h1)
	) name2953 (
		_w4301_,
		_w4302_,
		_w4303_
	);
	LUT3 #(
		.INIT('h01)
	) name2954 (
		_w4299_,
		_w4301_,
		_w4302_,
		_w4304_
	);
	LUT3 #(
		.INIT('h2a)
	) name2955 (
		_w4298_,
		_w4147_,
		_w4152_,
		_w4305_
	);
	LUT3 #(
		.INIT('h70)
	) name2956 (
		_w4160_,
		_w4165_,
		_w4300_,
		_w4306_
	);
	LUT3 #(
		.INIT('h23)
	) name2957 (
		_w4299_,
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2958 (
		_w4290_,
		_w4297_,
		_w4304_,
		_w4307_,
		_w4308_
	);
	LUT3 #(
		.INIT('h2a)
	) name2959 (
		_w4285_,
		_w4178_,
		_w4183_,
		_w4309_
	);
	LUT3 #(
		.INIT('h2a)
	) name2960 (
		_w4287_,
		_w4192_,
		_w4197_,
		_w4310_
	);
	LUT3 #(
		.INIT('h23)
	) name2961 (
		_w4286_,
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('h4504)
	) name2962 (
		_w4284_,
		_w4285_,
		_w4184_,
		_w4310_,
		_w4312_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2963 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4283_,
		_w4313_
	);
	LUT3 #(
		.INIT('h80)
	) name2964 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4282_,
		_w4314_
	);
	LUT3 #(
		.INIT('h6c)
	) name2965 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4282_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		_w4313_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		_w4312_,
		_w4316_,
		_w4317_
	);
	LUT4 #(
		.INIT('h8000)
	) name2968 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4215_,
		_w4318_
	);
	LUT3 #(
		.INIT('h6c)
	) name2969 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h8000)
	) name2970 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4282_,
		_w4320_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2971 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4282_,
		_w4321_
	);
	LUT3 #(
		.INIT('h32)
	) name2972 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4318_,
		_w4320_,
		_w4322_
	);
	LUT4 #(
		.INIT('hc301)
	) name2973 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4314_,
		_w4318_,
		_w4323_
	);
	LUT2 #(
		.INIT('h6)
	) name2974 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4318_,
		_w4324_
	);
	LUT3 #(
		.INIT('h04)
	) name2975 (
		_w4319_,
		_w4323_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h070f)
	) name2976 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4239_,
		_w4326_
	);
	LUT4 #(
		.INIT('h8000)
	) name2977 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4225_,
		_w4227_,
		_w4234_,
		_w4327_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w4326_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4327_,
		_w4329_
	);
	LUT4 #(
		.INIT('h8000)
	) name2980 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4330_
	);
	LUT3 #(
		.INIT('h80)
	) name2981 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4318_,
		_w4330_,
		_w4331_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		_w4329_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('hfc04)
	) name2983 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4326_,
		_w4327_,
		_w4331_,
		_w4333_
	);
	LUT4 #(
		.INIT('h820a)
	) name2984 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4234_,
		_w4334_
	);
	LUT3 #(
		.INIT('h80)
	) name2985 (
		_w4225_,
		_w4227_,
		_w4334_,
		_w4335_
	);
	LUT4 #(
		.INIT('h00ec)
	) name2986 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4318_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2987 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4237_,
		_w4238_,
		_w4337_
	);
	LUT3 #(
		.INIT('h02)
	) name2988 (
		_w4333_,
		_w4336_,
		_w4337_,
		_w4338_
	);
	LUT4 #(
		.INIT('h4000)
	) name2989 (
		_w4308_,
		_w4317_,
		_w4325_,
		_w4338_,
		_w4339_
	);
	LUT3 #(
		.INIT('h6a)
	) name2990 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4327_,
		_w4245_,
		_w4340_
	);
	LUT4 #(
		.INIT('h8000)
	) name2991 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4327_,
		_w4245_,
		_w4341_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2992 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4327_,
		_w4245_,
		_w4342_
	);
	LUT4 #(
		.INIT('h8111)
	) name2993 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4327_,
		_w4245_,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name2994 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4255_,
		_w4344_
	);
	LUT3 #(
		.INIT('h6c)
	) name2995 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4255_,
		_w4345_
	);
	LUT3 #(
		.INIT('h0e)
	) name2996 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4341_,
		_w4344_,
		_w4346_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2997 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4341_,
		_w4344_,
		_w4345_,
		_w4347_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		_w4343_,
		_w4347_,
		_w4348_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2999 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4255_,
		_w4349_
	);
	LUT3 #(
		.INIT('h80)
	) name3000 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4350_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3001 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4255_,
		_w4260_,
		_w4351_
	);
	LUT2 #(
		.INIT('h1)
	) name3002 (
		_w4349_,
		_w4351_,
		_w4352_
	);
	LUT4 #(
		.INIT('h8000)
	) name3003 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4353_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3004 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4354_
	);
	LUT4 #(
		.INIT('h8000)
	) name3005 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4255_,
		_w4263_,
		_w4262_,
		_w4355_
	);
	LUT3 #(
		.INIT('h0e)
	) name3006 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4353_,
		_w4355_,
		_w4356_
	);
	LUT4 #(
		.INIT('ha501)
	) name3007 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4350_,
		_w4355_,
		_w4357_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		_w4352_,
		_w4357_,
		_w4358_
	);
	LUT3 #(
		.INIT('h80)
	) name3009 (
		_w4339_,
		_w4348_,
		_w4358_,
		_w4359_
	);
	LUT3 #(
		.INIT('h6c)
	) name3010 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4269_,
		_w4360_
	);
	LUT3 #(
		.INIT('h6c)
	) name3011 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4268_,
		_w4361_
	);
	LUT4 #(
		.INIT('h8103)
	) name3012 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4268_,
		_w4362_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3013 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4269_,
		_w4363_
	);
	LUT4 #(
		.INIT('h8000)
	) name3014 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4272_,
		_w4364_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3015 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4272_,
		_w4365_
	);
	LUT2 #(
		.INIT('h1)
	) name3016 (
		_w4363_,
		_w4365_,
		_w4366_
	);
	LUT3 #(
		.INIT('h02)
	) name3017 (
		_w4362_,
		_w4363_,
		_w4365_,
		_w4367_
	);
	LUT4 #(
		.INIT('h8000)
	) name3018 (
		_w4339_,
		_w4348_,
		_w4358_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h74fc)
	) name3019 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4364_,
		_w4277_,
		_w4369_
	);
	LUT4 #(
		.INIT('h4554)
	) name3020 (
		_w1661_,
		_w4214_,
		_w4368_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3021 (
		_w1559_,
		_w4104_,
		_w4280_,
		_w4370_,
		_w4371_
	);
	LUT4 #(
		.INIT('hf800)
	) name3022 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4372_,
		_w4373_
	);
	LUT4 #(
		.INIT('h8000)
	) name3024 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4372_,
		_w4374_
	);
	LUT2 #(
		.INIT('h6)
	) name3025 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w4374_,
		_w4375_
	);
	LUT4 #(
		.INIT('hbf00)
	) name3026 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4375_,
		_w4376_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3027 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w4372_,
		_w4377_
	);
	LUT3 #(
		.INIT('h08)
	) name3028 (
		_w4178_,
		_w4183_,
		_w4377_,
		_w4378_
	);
	LUT3 #(
		.INIT('h6c)
	) name3029 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w4372_,
		_w4379_
	);
	LUT3 #(
		.INIT('h08)
	) name3030 (
		_w4192_,
		_w4197_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name3031 (
		_w4378_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h6)
	) name3032 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w4372_,
		_w4382_
	);
	LUT3 #(
		.INIT('h08)
	) name3033 (
		_w4147_,
		_w4152_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('h07f8)
	) name3034 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w4384_
	);
	LUT3 #(
		.INIT('h08)
	) name3035 (
		_w4160_,
		_w4165_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w4383_,
		_w4385_,
		_w4386_
	);
	LUT3 #(
		.INIT('h80)
	) name3037 (
		_w4109_,
		_w4114_,
		_w4291_,
		_w4387_
	);
	LUT3 #(
		.INIT('h07)
	) name3038 (
		_w4109_,
		_w4114_,
		_w4291_,
		_w4388_
	);
	LUT3 #(
		.INIT('h70)
	) name3039 (
		_w4121_,
		_w4126_,
		_w4293_,
		_w4389_
	);
	LUT3 #(
		.INIT('h15)
	) name3040 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4133_,
		_w4138_,
		_w4390_
	);
	LUT4 #(
		.INIT('h020b)
	) name3041 (
		_w4127_,
		_w4293_,
		_w4388_,
		_w4390_,
		_w4391_
	);
	LUT3 #(
		.INIT('h70)
	) name3042 (
		_w4147_,
		_w4152_,
		_w4382_,
		_w4392_
	);
	LUT3 #(
		.INIT('h70)
	) name3043 (
		_w4160_,
		_w4165_,
		_w4384_,
		_w4393_
	);
	LUT3 #(
		.INIT('h23)
	) name3044 (
		_w4383_,
		_w4392_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3045 (
		_w4386_,
		_w4387_,
		_w4391_,
		_w4394_,
		_w4395_
	);
	LUT3 #(
		.INIT('h70)
	) name3046 (
		_w4178_,
		_w4183_,
		_w4377_,
		_w4396_
	);
	LUT3 #(
		.INIT('h70)
	) name3047 (
		_w4192_,
		_w4197_,
		_w4379_,
		_w4397_
	);
	LUT3 #(
		.INIT('h23)
	) name3048 (
		_w4378_,
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT3 #(
		.INIT('hd0)
	) name3049 (
		_w4381_,
		_w4395_,
		_w4398_,
		_w4399_
	);
	LUT4 #(
		.INIT('h5100)
	) name3050 (
		_w4376_,
		_w4381_,
		_w4395_,
		_w4398_,
		_w4400_
	);
	LUT4 #(
		.INIT('h0040)
	) name3051 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4375_,
		_w4401_
	);
	LUT3 #(
		.INIT('h80)
	) name3052 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4374_,
		_w4402_
	);
	LUT3 #(
		.INIT('h6c)
	) name3053 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4374_,
		_w4403_
	);
	LUT2 #(
		.INIT('h4)
	) name3054 (
		_w4401_,
		_w4403_,
		_w4404_
	);
	LUT3 #(
		.INIT('h20)
	) name3055 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4401_,
		_w4403_,
		_w4405_
	);
	LUT4 #(
		.INIT('h8000)
	) name3056 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4374_,
		_w4406_
	);
	LUT3 #(
		.INIT('h6a)
	) name3057 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4402_,
		_w4407_
	);
	LUT4 #(
		.INIT('h60a0)
	) name3058 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4238_,
		_w4402_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('h8000)
	) name3060 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4238_,
		_w4406_,
		_w4410_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3061 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4238_,
		_w4406_,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name3062 (
		_w4245_,
		_w4411_,
		_w4412_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3063 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4410_,
		_w4413_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		_w4253_,
		_w4413_,
		_w4414_
	);
	LUT3 #(
		.INIT('h80)
	) name3065 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4253_,
		_w4413_,
		_w4415_
	);
	LUT4 #(
		.INIT('h8000)
	) name3066 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4253_,
		_w4412_,
		_w4413_,
		_w4416_
	);
	LUT4 #(
		.INIT('h4000)
	) name3067 (
		_w4400_,
		_w4405_,
		_w4409_,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3068 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4254_,
		_w4410_,
		_w4418_
	);
	LUT4 #(
		.INIT('h8000)
	) name3069 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4254_,
		_w4260_,
		_w4410_,
		_w4419_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3070 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w4254_,
		_w4260_,
		_w4410_,
		_w4420_
	);
	LUT2 #(
		.INIT('h8)
	) name3071 (
		_w4262_,
		_w4420_,
		_w4421_
	);
	LUT3 #(
		.INIT('h80)
	) name3072 (
		_w4417_,
		_w4418_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h8)
	) name3073 (
		_w4262_,
		_w4419_,
		_w4423_
	);
	LUT3 #(
		.INIT('h80)
	) name3074 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4262_,
		_w4419_,
		_w4424_
	);
	LUT4 #(
		.INIT('h8000)
	) name3075 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4262_,
		_w4272_,
		_w4419_,
		_w4425_
	);
	LUT3 #(
		.INIT('h6c)
	) name3076 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4424_,
		_w4426_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3077 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4424_,
		_w4427_
	);
	LUT3 #(
		.INIT('h6a)
	) name3078 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4262_,
		_w4419_,
		_w4428_
	);
	LUT4 #(
		.INIT('h4888)
	) name3079 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4262_,
		_w4419_,
		_w4429_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		_w4427_,
		_w4429_,
		_w4430_
	);
	LUT4 #(
		.INIT('h8000)
	) name3081 (
		_w4417_,
		_w4418_,
		_w4421_,
		_w4430_,
		_w4431_
	);
	LUT3 #(
		.INIT('h6c)
	) name3082 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4425_,
		_w4432_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3083 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w1640_,
		_w4425_,
		_w4433_
	);
	LUT3 #(
		.INIT('hb0)
	) name3084 (
		_w1571_,
		_w1583_,
		_w4369_,
		_w4434_
	);
	LUT4 #(
		.INIT('h0c04)
	) name3085 (
		_w1604_,
		_w1605_,
		_w1602_,
		_w1616_,
		_w4435_
	);
	LUT4 #(
		.INIT('h0010)
	) name3086 (
		_w1625_,
		_w1626_,
		_w1643_,
		_w1667_,
		_w4436_
	);
	LUT3 #(
		.INIT('h8a)
	) name3087 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name3088 (
		_w1617_,
		_w4279_,
		_w4438_
	);
	LUT4 #(
		.INIT('h0001)
	) name3089 (
		_w4433_,
		_w4437_,
		_w4434_,
		_w4438_,
		_w4439_
	);
	LUT4 #(
		.INIT('hd700)
	) name3090 (
		_w1659_,
		_w4431_,
		_w4432_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('hfc21)
	) name3091 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w4441_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3092 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2286_,
		_w4441_,
		_w4442_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3093 (
		_w1678_,
		_w4371_,
		_w4440_,
		_w4442_,
		_w4443_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3094 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w3063_,
		_w3065_,
		_w4444_
	);
	LUT4 #(
		.INIT('h7000)
	) name3095 (
		_w3095_,
		_w3100_,
		_w3269_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h8)
	) name3096 (
		_w3271_,
		_w3992_,
		_w4446_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3097 (
		_w3285_,
		_w3290_,
		_w3294_,
		_w4446_,
		_w4447_
	);
	LUT3 #(
		.INIT('h6a)
	) name3098 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w3072_,
		_w3074_,
		_w4448_
	);
	LUT3 #(
		.INIT('h80)
	) name3099 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3308_,
		_w4448_,
		_w4449_
	);
	LUT3 #(
		.INIT('h6a)
	) name3100 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w3072_,
		_w3073_,
		_w4450_
	);
	LUT4 #(
		.INIT('h8000)
	) name3101 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w3308_,
		_w4448_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h8000)
	) name3102 (
		_w3305_,
		_w3301_,
		_w3298_,
		_w3303_,
		_w4452_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		_w4451_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('h0155)
	) name3104 (
		_w3315_,
		_w4445_,
		_w4447_,
		_w4453_,
		_w4454_
	);
	LUT4 #(
		.INIT('h5554)
	) name3105 (
		_w3280_,
		_w3273_,
		_w3276_,
		_w3283_,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name3106 (
		_w3289_,
		_w3278_,
		_w4456_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w3270_,
		_w3287_,
		_w4457_
	);
	LUT4 #(
		.INIT('h0001)
	) name3108 (
		_w3270_,
		_w3287_,
		_w3289_,
		_w3278_,
		_w4458_
	);
	LUT3 #(
		.INIT('h0b)
	) name3109 (
		_w3289_,
		_w3282_,
		_w3293_,
		_w4459_
	);
	LUT4 #(
		.INIT('h004d)
	) name3110 (
		_w3288_,
		_w3114_,
		_w3282_,
		_w3292_,
		_w4460_
	);
	LUT3 #(
		.INIT('h51)
	) name3111 (
		_w3291_,
		_w4457_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h8)
	) name3112 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w4444_,
		_w4462_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3113 (
		_w4455_,
		_w4458_,
		_w4461_,
		_w4462_,
		_w4463_
	);
	LUT3 #(
		.INIT('h6a)
	) name3114 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3063_,
		_w3067_,
		_w4464_
	);
	LUT3 #(
		.INIT('h80)
	) name3115 (
		_w3070_,
		_w3302_,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h8)
	) name3116 (
		_w4463_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		_w3306_,
		_w3298_,
		_w4467_
	);
	LUT3 #(
		.INIT('h80)
	) name3118 (
		_w4463_,
		_w4465_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h8)
	) name3119 (
		_w3315_,
		_w4449_,
		_w4469_
	);
	LUT4 #(
		.INIT('h8000)
	) name3120 (
		_w4463_,
		_w4465_,
		_w4467_,
		_w4469_,
		_w4470_
	);
	LUT3 #(
		.INIT('h02)
	) name3121 (
		_w3101_,
		_w4470_,
		_w4454_,
		_w4471_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3122 (
		_w3130_,
		_w4000_,
		_w4001_,
		_w4002_,
		_w4472_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		_w4008_,
		_w4004_,
		_w4473_
	);
	LUT4 #(
		.INIT('hae00)
	) name3124 (
		_w3103_,
		_w4005_,
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT3 #(
		.INIT('h04)
	) name3125 (
		_w3216_,
		_w3222_,
		_w3254_,
		_w4475_
	);
	LUT2 #(
		.INIT('h4)
	) name3126 (
		_w3235_,
		_w3253_,
		_w4476_
	);
	LUT3 #(
		.INIT('h10)
	) name3127 (
		_w3235_,
		_w3237_,
		_w3253_,
		_w4477_
	);
	LUT4 #(
		.INIT('h8000)
	) name3128 (
		_w3248_,
		_w4474_,
		_w4475_,
		_w4477_,
		_w4478_
	);
	LUT3 #(
		.INIT('h14)
	) name3129 (
		_w3101_,
		_w3232_,
		_w4478_,
		_w4479_
	);
	LUT4 #(
		.INIT('h4447)
	) name3130 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1916_,
		_w4471_,
		_w4479_,
		_w4480_
	);
	LUT3 #(
		.INIT('h32)
	) name3131 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w3378_,
		_w3381_,
		_w4481_
	);
	LUT4 #(
		.INIT('h8000)
	) name3132 (
		_w3073_,
		_w3375_,
		_w3368_,
		_w3382_,
		_w4482_
	);
	LUT4 #(
		.INIT('h4000)
	) name3133 (
		_w4023_,
		_w4025_,
		_w4028_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('h28)
	) name3134 (
		_w1924_,
		_w4481_,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name3135 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1846_,
		_w3378_,
		_w3381_,
		_w4485_
	);
	LUT3 #(
		.INIT('h54)
	) name3136 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1842_,
		_w1845_,
		_w4486_
	);
	LUT3 #(
		.INIT('h01)
	) name3137 (
		_w1833_,
		_w4486_,
		_w4485_,
		_w4487_
	);
	LUT4 #(
		.INIT('h0e00)
	) name3138 (
		_w1855_,
		_w1860_,
		_w1861_,
		_w3231_,
		_w4488_
	);
	LUT4 #(
		.INIT('hfe00)
	) name3139 (
		_w1795_,
		_w1797_,
		_w1802_,
		_w3315_,
		_w4489_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w1913_,
		_w4489_,
		_w4490_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name3141 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w1868_,
		_w4488_,
		_w4490_,
		_w4491_
	);
	LUT3 #(
		.INIT('h80)
	) name3142 (
		_w1805_,
		_w1806_,
		_w3315_,
		_w4492_
	);
	LUT4 #(
		.INIT('h004f)
	) name3143 (
		_w1816_,
		_w1831_,
		_w3232_,
		_w4492_,
		_w4493_
	);
	LUT3 #(
		.INIT('h10)
	) name3144 (
		_w4491_,
		_w4487_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		_w4484_,
		_w4494_,
		_w4495_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3146 (
		_w1810_,
		_w1933_,
		_w4480_,
		_w4495_,
		_w4496_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w3406_,
		_w4497_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3148 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w3406_,
		_w3408_,
		_w4498_
	);
	LUT2 #(
		.INIT('hb)
	) name3149 (
		_w4496_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('hc444)
	) name3150 (
		\address1[29]_pad ,
		\datai[29]_pad ,
		_w3419_,
		_w3424_,
		_w4500_
	);
	LUT4 #(
		.INIT('h0888)
	) name3151 (
		\address1[29]_pad ,
		\buf1_reg[29]/NET0131 ,
		_w3419_,
		_w3424_,
		_w4501_
	);
	LUT2 #(
		.INIT('h1)
	) name3152 (
		_w4500_,
		_w4501_,
		_w4502_
	);
	LUT4 #(
		.INIT('h0002)
	) name3153 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w4502_,
		_w4503_
	);
	LUT4 #(
		.INIT('hc444)
	) name3154 (
		\address1[29]_pad ,
		\datai[30]_pad ,
		_w3419_,
		_w3424_,
		_w4504_
	);
	LUT4 #(
		.INIT('h0888)
	) name3155 (
		\address1[29]_pad ,
		\buf1_reg[30]/NET0131 ,
		_w3419_,
		_w3424_,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name3156 (
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT4 #(
		.INIT('h8828)
	) name3157 (
		_w3411_,
		_w3425_,
		_w4503_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('h0100)
	) name3158 (
		_w3503_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w4508_
	);
	LUT3 #(
		.INIT('h82)
	) name3159 (
		_w3412_,
		_w3507_,
		_w4508_,
		_w4509_
	);
	LUT3 #(
		.INIT('h02)
	) name3160 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w3534_,
		_w3536_,
		_w4510_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3161 (
		_w3537_,
		_w3436_,
		_w3437_,
		_w4510_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w3414_,
		_w4511_,
		_w4512_
	);
	LUT4 #(
		.INIT('h0057)
	) name3163 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4507_,
		_w4509_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h2)
	) name3164 (
		_w3407_,
		_w4511_,
		_w4514_
	);
	LUT4 #(
		.INIT('hc055)
	) name3165 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3534_,
		_w4515_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		_w3545_,
		_w4516_
	);
	LUT3 #(
		.INIT('h0d)
	) name3167 (
		_w2248_,
		_w4515_,
		_w4516_,
		_w4517_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		_w4514_,
		_w4517_,
		_w4518_
	);
	LUT3 #(
		.INIT('h2f)
	) name3169 (
		_w1939_,
		_w4513_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('h8848)
	) name3170 (
		_w3425_,
		_w3572_,
		_w4503_,
		_w4506_,
		_w4520_
	);
	LUT3 #(
		.INIT('h84)
	) name3171 (
		_w3507_,
		_w3573_,
		_w4508_,
		_w4521_
	);
	LUT3 #(
		.INIT('h02)
	) name3172 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w3578_,
		_w3580_,
		_w4522_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3173 (
		_w3436_,
		_w3437_,
		_w3581_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h1)
	) name3174 (
		_w3575_,
		_w4523_,
		_w4524_
	);
	LUT4 #(
		.INIT('h0057)
	) name3175 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4520_,
		_w4521_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h2)
	) name3176 (
		_w3407_,
		_w4523_,
		_w4526_
	);
	LUT4 #(
		.INIT('hc055)
	) name3177 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3578_,
		_w4527_
	);
	LUT2 #(
		.INIT('h2)
	) name3178 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		_w3545_,
		_w4528_
	);
	LUT3 #(
		.INIT('h0d)
	) name3179 (
		_w2248_,
		_w4527_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h4)
	) name3180 (
		_w4526_,
		_w4529_,
		_w4530_
	);
	LUT3 #(
		.INIT('h2f)
	) name3181 (
		_w1939_,
		_w4525_,
		_w4530_,
		_w4531_
	);
	LUT4 #(
		.INIT('h8848)
	) name3182 (
		_w3425_,
		_w3592_,
		_w4503_,
		_w4506_,
		_w4532_
	);
	LUT3 #(
		.INIT('h82)
	) name3183 (
		_w3411_,
		_w3507_,
		_w4508_,
		_w4533_
	);
	LUT3 #(
		.INIT('h02)
	) name3184 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		_w3536_,
		_w3412_,
		_w4534_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3185 (
		_w3436_,
		_w3437_,
		_w3597_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h1)
	) name3186 (
		_w3594_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h0057)
	) name3187 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4532_,
		_w4533_,
		_w4536_,
		_w4537_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		_w3407_,
		_w4535_,
		_w4538_
	);
	LUT4 #(
		.INIT('hc055)
	) name3189 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3536_,
		_w4539_
	);
	LUT2 #(
		.INIT('h2)
	) name3190 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		_w3545_,
		_w4540_
	);
	LUT3 #(
		.INIT('h0d)
	) name3191 (
		_w2248_,
		_w4539_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h4)
	) name3192 (
		_w4538_,
		_w4541_,
		_w4542_
	);
	LUT3 #(
		.INIT('h2f)
	) name3193 (
		_w1939_,
		_w4537_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('h8828)
	) name3194 (
		_w3412_,
		_w3425_,
		_w4503_,
		_w4506_,
		_w4544_
	);
	LUT3 #(
		.INIT('h82)
	) name3195 (
		_w3536_,
		_w3507_,
		_w4508_,
		_w4545_
	);
	LUT3 #(
		.INIT('h02)
	) name3196 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w3534_,
		_w3611_,
		_w4546_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3197 (
		_w3436_,
		_w3437_,
		_w3612_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h1)
	) name3198 (
		_w3608_,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h0057)
	) name3199 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4544_,
		_w4545_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h2)
	) name3200 (
		_w3407_,
		_w4547_,
		_w4550_
	);
	LUT4 #(
		.INIT('hc055)
	) name3201 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3611_,
		_w4551_
	);
	LUT2 #(
		.INIT('h2)
	) name3202 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w3545_,
		_w4552_
	);
	LUT3 #(
		.INIT('h0d)
	) name3203 (
		_w2248_,
		_w4551_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h4)
	) name3204 (
		_w4550_,
		_w4553_,
		_w4554_
	);
	LUT3 #(
		.INIT('h2f)
	) name3205 (
		_w1939_,
		_w4549_,
		_w4554_,
		_w4555_
	);
	LUT4 #(
		.INIT('h8828)
	) name3206 (
		_w3536_,
		_w3425_,
		_w4503_,
		_w4506_,
		_w4556_
	);
	LUT3 #(
		.INIT('h82)
	) name3207 (
		_w3534_,
		_w3507_,
		_w4508_,
		_w4557_
	);
	LUT3 #(
		.INIT('h02)
	) name3208 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w3572_,
		_w3611_,
		_w4558_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3209 (
		_w3436_,
		_w3437_,
		_w3626_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w3623_,
		_w4559_,
		_w4560_
	);
	LUT4 #(
		.INIT('h0057)
	) name3211 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4556_,
		_w4557_,
		_w4560_,
		_w4561_
	);
	LUT2 #(
		.INIT('h2)
	) name3212 (
		_w3407_,
		_w4559_,
		_w4562_
	);
	LUT4 #(
		.INIT('hc055)
	) name3213 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3572_,
		_w4563_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w3545_,
		_w4564_
	);
	LUT3 #(
		.INIT('h0d)
	) name3215 (
		_w2248_,
		_w4563_,
		_w4564_,
		_w4565_
	);
	LUT2 #(
		.INIT('h4)
	) name3216 (
		_w4562_,
		_w4565_,
		_w4566_
	);
	LUT3 #(
		.INIT('h2f)
	) name3217 (
		_w1939_,
		_w4561_,
		_w4566_,
		_w4567_
	);
	LUT4 #(
		.INIT('h8828)
	) name3218 (
		_w3534_,
		_w3425_,
		_w4503_,
		_w4506_,
		_w4568_
	);
	LUT3 #(
		.INIT('h84)
	) name3219 (
		_w3507_,
		_w3611_,
		_w4508_,
		_w4569_
	);
	LUT3 #(
		.INIT('h02)
	) name3220 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w3572_,
		_w3573_,
		_w4570_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3221 (
		_w3436_,
		_w3437_,
		_w3574_,
		_w4570_,
		_w4571_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w3637_,
		_w4571_,
		_w4572_
	);
	LUT4 #(
		.INIT('h0057)
	) name3223 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4568_,
		_w4569_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h2)
	) name3224 (
		_w3407_,
		_w4571_,
		_w4574_
	);
	LUT4 #(
		.INIT('hc055)
	) name3225 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3573_,
		_w4575_
	);
	LUT2 #(
		.INIT('h2)
	) name3226 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w3545_,
		_w4576_
	);
	LUT3 #(
		.INIT('h0d)
	) name3227 (
		_w2248_,
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h4)
	) name3228 (
		_w4574_,
		_w4577_,
		_w4578_
	);
	LUT3 #(
		.INIT('h2f)
	) name3229 (
		_w1939_,
		_w4573_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('h8848)
	) name3230 (
		_w3425_,
		_w3611_,
		_w4503_,
		_w4506_,
		_w4580_
	);
	LUT3 #(
		.INIT('h84)
	) name3231 (
		_w3507_,
		_w3572_,
		_w4508_,
		_w4581_
	);
	LUT3 #(
		.INIT('h02)
	) name3232 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w3580_,
		_w3573_,
		_w4582_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3233 (
		_w3436_,
		_w3437_,
		_w3653_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h1)
	) name3234 (
		_w3650_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('h0057)
	) name3235 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4580_,
		_w4581_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name3236 (
		_w3407_,
		_w4583_,
		_w4586_
	);
	LUT4 #(
		.INIT('hc055)
	) name3237 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3580_,
		_w4587_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w3545_,
		_w4588_
	);
	LUT3 #(
		.INIT('h0d)
	) name3239 (
		_w2248_,
		_w4587_,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h4)
	) name3240 (
		_w4586_,
		_w4589_,
		_w4590_
	);
	LUT3 #(
		.INIT('h2f)
	) name3241 (
		_w1939_,
		_w4585_,
		_w4590_,
		_w4591_
	);
	LUT4 #(
		.INIT('h8848)
	) name3242 (
		_w3425_,
		_w3573_,
		_w4503_,
		_w4506_,
		_w4592_
	);
	LUT3 #(
		.INIT('h84)
	) name3243 (
		_w3507_,
		_w3580_,
		_w4508_,
		_w4593_
	);
	LUT3 #(
		.INIT('h02)
	) name3244 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w3578_,
		_w3667_,
		_w4594_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3245 (
		_w3436_,
		_w3437_,
		_w3668_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name3246 (
		_w3664_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h0057)
	) name3247 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4592_,
		_w4593_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3248 (
		_w3407_,
		_w4595_,
		_w4598_
	);
	LUT4 #(
		.INIT('hc055)
	) name3249 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3667_,
		_w4599_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w3545_,
		_w4600_
	);
	LUT3 #(
		.INIT('h0d)
	) name3251 (
		_w2248_,
		_w4599_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h4)
	) name3252 (
		_w4598_,
		_w4601_,
		_w4602_
	);
	LUT3 #(
		.INIT('h2f)
	) name3253 (
		_w1939_,
		_w4597_,
		_w4602_,
		_w4603_
	);
	LUT4 #(
		.INIT('h8848)
	) name3254 (
		_w3425_,
		_w3580_,
		_w4503_,
		_w4506_,
		_w4604_
	);
	LUT3 #(
		.INIT('h84)
	) name3255 (
		_w3507_,
		_w3578_,
		_w4508_,
		_w4605_
	);
	LUT3 #(
		.INIT('h02)
	) name3256 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w3667_,
		_w3683_,
		_w4606_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3257 (
		_w3436_,
		_w3437_,
		_w3698_,
		_w4606_,
		_w4607_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w3695_,
		_w4607_,
		_w4608_
	);
	LUT4 #(
		.INIT('h0057)
	) name3259 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4604_,
		_w4605_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		_w3407_,
		_w4607_,
		_w4610_
	);
	LUT4 #(
		.INIT('hc055)
	) name3261 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3683_,
		_w4611_
	);
	LUT2 #(
		.INIT('h2)
	) name3262 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w3545_,
		_w4612_
	);
	LUT3 #(
		.INIT('h0d)
	) name3263 (
		_w2248_,
		_w4611_,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h4)
	) name3264 (
		_w4610_,
		_w4613_,
		_w4614_
	);
	LUT3 #(
		.INIT('h2f)
	) name3265 (
		_w1939_,
		_w4609_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('h8848)
	) name3266 (
		_w3425_,
		_w3578_,
		_w4503_,
		_w4506_,
		_w4616_
	);
	LUT3 #(
		.INIT('h84)
	) name3267 (
		_w3507_,
		_w3667_,
		_w4508_,
		_w4617_
	);
	LUT3 #(
		.INIT('h02)
	) name3268 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w3682_,
		_w3683_,
		_w4618_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3269 (
		_w3436_,
		_w3437_,
		_w3684_,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w3679_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h0057)
	) name3271 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4616_,
		_w4617_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		_w3407_,
		_w4619_,
		_w4622_
	);
	LUT4 #(
		.INIT('hc055)
	) name3273 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3682_,
		_w4623_
	);
	LUT2 #(
		.INIT('h2)
	) name3274 (
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w3545_,
		_w4624_
	);
	LUT3 #(
		.INIT('h0d)
	) name3275 (
		_w2248_,
		_w4623_,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h4)
	) name3276 (
		_w4622_,
		_w4625_,
		_w4626_
	);
	LUT3 #(
		.INIT('h2f)
	) name3277 (
		_w1939_,
		_w4621_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('h8848)
	) name3278 (
		_w3425_,
		_w3667_,
		_w4503_,
		_w4506_,
		_w4628_
	);
	LUT3 #(
		.INIT('h84)
	) name3279 (
		_w3507_,
		_w3683_,
		_w4508_,
		_w4629_
	);
	LUT3 #(
		.INIT('h02)
	) name3280 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w3682_,
		_w3712_,
		_w4630_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3281 (
		_w3436_,
		_w3437_,
		_w3713_,
		_w4630_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w3709_,
		_w4631_,
		_w4632_
	);
	LUT4 #(
		.INIT('h0057)
	) name3283 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4628_,
		_w4629_,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h2)
	) name3284 (
		_w3407_,
		_w4631_,
		_w4634_
	);
	LUT4 #(
		.INIT('hc055)
	) name3285 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3712_,
		_w4635_
	);
	LUT2 #(
		.INIT('h2)
	) name3286 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w3545_,
		_w4636_
	);
	LUT3 #(
		.INIT('h0d)
	) name3287 (
		_w2248_,
		_w4635_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h4)
	) name3288 (
		_w4634_,
		_w4637_,
		_w4638_
	);
	LUT3 #(
		.INIT('h2f)
	) name3289 (
		_w1939_,
		_w4633_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h8848)
	) name3290 (
		_w3425_,
		_w3683_,
		_w4503_,
		_w4506_,
		_w4640_
	);
	LUT3 #(
		.INIT('h84)
	) name3291 (
		_w3507_,
		_w3682_,
		_w4508_,
		_w4641_
	);
	LUT3 #(
		.INIT('h02)
	) name3292 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w3712_,
		_w3727_,
		_w4642_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3293 (
		_w3436_,
		_w3437_,
		_w3728_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w3724_,
		_w4643_,
		_w4644_
	);
	LUT4 #(
		.INIT('h0057)
	) name3295 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4640_,
		_w4641_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h2)
	) name3296 (
		_w3407_,
		_w4643_,
		_w4646_
	);
	LUT4 #(
		.INIT('hc055)
	) name3297 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3727_,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name3298 (
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w3545_,
		_w4648_
	);
	LUT3 #(
		.INIT('h0d)
	) name3299 (
		_w2248_,
		_w4647_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h4)
	) name3300 (
		_w4646_,
		_w4649_,
		_w4650_
	);
	LUT3 #(
		.INIT('h2f)
	) name3301 (
		_w1939_,
		_w4645_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('h8848)
	) name3302 (
		_w3425_,
		_w3682_,
		_w4503_,
		_w4506_,
		_w4652_
	);
	LUT3 #(
		.INIT('h84)
	) name3303 (
		_w3507_,
		_w3712_,
		_w4508_,
		_w4653_
	);
	LUT3 #(
		.INIT('h02)
	) name3304 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w3727_,
		_w3742_,
		_w4654_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3305 (
		_w3436_,
		_w3437_,
		_w3743_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w3739_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h0057)
	) name3307 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4652_,
		_w4653_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h2)
	) name3308 (
		_w3407_,
		_w4655_,
		_w4658_
	);
	LUT4 #(
		.INIT('hc055)
	) name3309 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3742_,
		_w4659_
	);
	LUT2 #(
		.INIT('h2)
	) name3310 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w3545_,
		_w4660_
	);
	LUT3 #(
		.INIT('h0d)
	) name3311 (
		_w2248_,
		_w4659_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h4)
	) name3312 (
		_w4658_,
		_w4661_,
		_w4662_
	);
	LUT3 #(
		.INIT('h2f)
	) name3313 (
		_w1939_,
		_w4657_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h8848)
	) name3314 (
		_w3425_,
		_w3712_,
		_w4503_,
		_w4506_,
		_w4664_
	);
	LUT3 #(
		.INIT('h84)
	) name3315 (
		_w3507_,
		_w3727_,
		_w4508_,
		_w4665_
	);
	LUT3 #(
		.INIT('h02)
	) name3316 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w3592_,
		_w3742_,
		_w4666_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3317 (
		_w3436_,
		_w3437_,
		_w3757_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h1)
	) name3318 (
		_w3754_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h0057)
	) name3319 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4664_,
		_w4665_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h2)
	) name3320 (
		_w3407_,
		_w4667_,
		_w4670_
	);
	LUT4 #(
		.INIT('hc055)
	) name3321 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3592_,
		_w4671_
	);
	LUT2 #(
		.INIT('h2)
	) name3322 (
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w3545_,
		_w4672_
	);
	LUT3 #(
		.INIT('h0d)
	) name3323 (
		_w2248_,
		_w4671_,
		_w4672_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		_w4670_,
		_w4673_,
		_w4674_
	);
	LUT3 #(
		.INIT('h2f)
	) name3325 (
		_w1939_,
		_w4669_,
		_w4674_,
		_w4675_
	);
	LUT4 #(
		.INIT('h8848)
	) name3326 (
		_w3425_,
		_w3727_,
		_w4503_,
		_w4506_,
		_w4676_
	);
	LUT3 #(
		.INIT('h84)
	) name3327 (
		_w3507_,
		_w3742_,
		_w4508_,
		_w4677_
	);
	LUT3 #(
		.INIT('h02)
	) name3328 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w3411_,
		_w3592_,
		_w4678_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3329 (
		_w3436_,
		_w3437_,
		_w3593_,
		_w4678_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		_w3768_,
		_w4679_,
		_w4680_
	);
	LUT4 #(
		.INIT('h0057)
	) name3331 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4676_,
		_w4677_,
		_w4680_,
		_w4681_
	);
	LUT2 #(
		.INIT('h2)
	) name3332 (
		_w3407_,
		_w4679_,
		_w4682_
	);
	LUT4 #(
		.INIT('hc055)
	) name3333 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3411_,
		_w4683_
	);
	LUT2 #(
		.INIT('h2)
	) name3334 (
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w3545_,
		_w4684_
	);
	LUT3 #(
		.INIT('h0d)
	) name3335 (
		_w2248_,
		_w4683_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h4)
	) name3336 (
		_w4682_,
		_w4685_,
		_w4686_
	);
	LUT3 #(
		.INIT('h2f)
	) name3337 (
		_w1939_,
		_w4681_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h8848)
	) name3338 (
		_w3425_,
		_w3742_,
		_w4503_,
		_w4506_,
		_w4688_
	);
	LUT3 #(
		.INIT('h84)
	) name3339 (
		_w3507_,
		_w3592_,
		_w4508_,
		_w4689_
	);
	LUT3 #(
		.INIT('h02)
	) name3340 (
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w3411_,
		_w3412_,
		_w4690_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3341 (
		_w3413_,
		_w3436_,
		_w3437_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w3781_,
		_w4691_,
		_w4692_
	);
	LUT4 #(
		.INIT('h0057)
	) name3343 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w4688_,
		_w4689_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name3344 (
		_w3407_,
		_w4691_,
		_w4694_
	);
	LUT4 #(
		.INIT('hc055)
	) name3345 (
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1765_,
		_w1770_,
		_w3412_,
		_w4695_
	);
	LUT2 #(
		.INIT('h2)
	) name3346 (
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w3545_,
		_w4696_
	);
	LUT3 #(
		.INIT('h0d)
	) name3347 (
		_w2248_,
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT2 #(
		.INIT('h4)
	) name3348 (
		_w4694_,
		_w4697_,
		_w4698_
	);
	LUT3 #(
		.INIT('h2f)
	) name3349 (
		_w1939_,
		_w4693_,
		_w4698_,
		_w4699_
	);
	LUT3 #(
		.INIT('h08)
	) name3350 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w1842_,
		_w1915_,
		_w4700_
	);
	LUT3 #(
		.INIT('h6c)
	) name3351 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3078_,
		_w4701_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w3316_,
		_w3997_,
		_w4702_
	);
	LUT3 #(
		.INIT('h80)
	) name3353 (
		_w3316_,
		_w3317_,
		_w3997_,
		_w4703_
	);
	LUT4 #(
		.INIT('h820a)
	) name3354 (
		_w3101_,
		_w3996_,
		_w4701_,
		_w4703_,
		_w4704_
	);
	LUT4 #(
		.INIT('h4554)
	) name3355 (
		_w1916_,
		_w3101_,
		_w3257_,
		_w3259_,
		_w4705_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3356 (
		_w1810_,
		_w4700_,
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT3 #(
		.INIT('h20)
	) name3357 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w1846_,
		_w3379_,
		_w4707_
	);
	LUT3 #(
		.INIT('h04)
	) name3358 (
		_w1833_,
		_w3386_,
		_w4707_,
		_w4708_
	);
	LUT2 #(
		.INIT('h2)
	) name3359 (
		_w1795_,
		_w1852_,
		_w4709_
	);
	LUT4 #(
		.INIT('h5f13)
	) name3360 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w1852_,
		_w4710_
	);
	LUT4 #(
		.INIT('haf23)
	) name3361 (
		_w1852_,
		_w1861_,
		_w1921_,
		_w4710_,
		_w4711_
	);
	LUT3 #(
		.INIT('h2a)
	) name3362 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w4037_,
		_w4711_,
		_w4712_
	);
	LUT3 #(
		.INIT('hb0)
	) name3363 (
		_w1816_,
		_w1831_,
		_w3259_,
		_w4713_
	);
	LUT2 #(
		.INIT('h4)
	) name3364 (
		_w1862_,
		_w4701_,
		_w4714_
	);
	LUT4 #(
		.INIT('h0001)
	) name3365 (
		_w4712_,
		_w4713_,
		_w4714_,
		_w4708_,
		_w4715_
	);
	LUT4 #(
		.INIT('hd700)
	) name3366 (
		_w1924_,
		_w3385_,
		_w3386_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name3367 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w3406_,
		_w4717_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3368 (
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w3406_,
		_w3408_,
		_w4718_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3369 (
		_w1933_,
		_w4706_,
		_w4716_,
		_w4718_,
		_w4719_
	);
	LUT3 #(
		.INIT('h08)
	) name3370 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w1842_,
		_w1915_,
		_w4720_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3371 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3072_,
		_w3074_,
		_w3076_,
		_w4721_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name3372 (
		_w3996_,
		_w4470_,
		_w4702_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h2)
	) name3373 (
		_w3101_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h0075)
	) name3374 (
		_w3131_,
		_w3203_,
		_w3206_,
		_w3209_,
		_w4724_
	);
	LUT3 #(
		.INIT('h10)
	) name3375 (
		_w3210_,
		_w3216_,
		_w4008_,
		_w4725_
	);
	LUT2 #(
		.INIT('h1)
	) name3376 (
		_w3243_,
		_w3254_,
		_w4726_
	);
	LUT3 #(
		.INIT('h02)
	) name3377 (
		_w3222_,
		_w3243_,
		_w3254_,
		_w4727_
	);
	LUT2 #(
		.INIT('h2)
	) name3378 (
		_w3247_,
		_w3250_,
		_w4728_
	);
	LUT4 #(
		.INIT('h8000)
	) name3379 (
		_w4724_,
		_w4725_,
		_w4727_,
		_w4728_,
		_w4729_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name3380 (
		_w3229_,
		_w3238_,
		_w3252_,
		_w4729_,
		_w4730_
	);
	LUT4 #(
		.INIT('h1555)
	) name3381 (
		_w3101_,
		_w3239_,
		_w3255_,
		_w4011_,
		_w4731_
	);
	LUT3 #(
		.INIT('h45)
	) name3382 (
		_w1916_,
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3383 (
		_w1810_,
		_w4720_,
		_w4723_,
		_w4732_,
		_w4733_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3384 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w3074_,
		_w3076_,
		_w3366_,
		_w4734_
	);
	LUT4 #(
		.INIT('h2000)
	) name3385 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w3356_,
		_w3359_,
		_w4028_,
		_w4735_
	);
	LUT3 #(
		.INIT('h80)
	) name3386 (
		\P1_InstAddrPointer_reg[23]/NET0131 ,
		_w3382_,
		_w4017_,
		_w4736_
	);
	LUT3 #(
		.INIT('h80)
	) name3387 (
		_w4029_,
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT4 #(
		.INIT('h8000)
	) name3388 (
		_w4029_,
		_w4734_,
		_w4735_,
		_w4736_,
		_w4738_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3389 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w1852_,
		_w4739_
	);
	LUT4 #(
		.INIT('h0103)
	) name3390 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w1855_,
		_w1860_,
		_w4739_,
		_w4740_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w1858_,
		_w4739_,
		_w4741_
	);
	LUT4 #(
		.INIT('h00c4)
	) name3392 (
		_w1861_,
		_w4037_,
		_w4740_,
		_w4741_,
		_w4742_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name3393 (
		_w1807_,
		_w1861_,
		_w4721_,
		_w4740_,
		_w4743_
	);
	LUT3 #(
		.INIT('h40)
	) name3394 (
		_w1833_,
		_w1846_,
		_w4734_,
		_w4744_
	);
	LUT4 #(
		.INIT('h004f)
	) name3395 (
		_w1816_,
		_w1831_,
		_w3229_,
		_w4744_,
		_w4745_
	);
	LUT4 #(
		.INIT('h3100)
	) name3396 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		_w4743_,
		_w4742_,
		_w4745_,
		_w4746_
	);
	LUT4 #(
		.INIT('hd700)
	) name3397 (
		_w1924_,
		_w4734_,
		_w4737_,
		_w4746_,
		_w4747_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3398 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w3406_,
		_w3408_,
		_w4748_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3399 (
		_w1933_,
		_w4733_,
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT3 #(
		.INIT('h02)
	) name3400 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2103_,
		_w2172_,
		_w4750_
	);
	LUT3 #(
		.INIT('h08)
	) name3401 (
		_w2874_,
		_w2884_,
		_w2891_,
		_w4751_
	);
	LUT4 #(
		.INIT('h4015)
	) name3402 (
		_w2755_,
		_w2874_,
		_w2884_,
		_w2891_,
		_w4752_
	);
	LUT4 #(
		.INIT('h004f)
	) name3403 (
		_w2935_,
		_w2941_,
		_w2952_,
		_w2957_,
		_w4753_
	);
	LUT4 #(
		.INIT('h00bf)
	) name3404 (
		_w4051_,
		_w4054_,
		_w4056_,
		_w4753_,
		_w4754_
	);
	LUT4 #(
		.INIT('h0051)
	) name3405 (
		_w2173_,
		_w2755_,
		_w4754_,
		_w4752_,
		_w4755_
	);
	LUT3 #(
		.INIT('ha8)
	) name3406 (
		_w2171_,
		_w4750_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h6)
	) name3407 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w3022_,
		_w4757_
	);
	LUT4 #(
		.INIT('ha800)
	) name3408 (
		_w2991_,
		_w2993_,
		_w3020_,
		_w3023_,
		_w4758_
	);
	LUT4 #(
		.INIT('h4448)
	) name3409 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2181_,
		_w3022_,
		_w4758_,
		_w4759_
	);
	LUT4 #(
		.INIT('h5155)
	) name3410 (
		_w2065_,
		_w2122_,
		_w2125_,
		_w2954_,
		_w4760_
	);
	LUT4 #(
		.INIT('hba00)
	) name3411 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2117_,
		_w2893_,
		_w4760_,
		_w4761_
	);
	LUT3 #(
		.INIT('hb0)
	) name3412 (
		_w2073_,
		_w2086_,
		_w2891_,
		_w4762_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2098_,
		_w4763_
	);
	LUT3 #(
		.INIT('he0)
	) name3414 (
		_w2071_,
		_w2087_,
		_w4757_,
		_w4764_
	);
	LUT3 #(
		.INIT('h31)
	) name3415 (
		_w2176_,
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT3 #(
		.INIT('h01)
	) name3416 (
		_w4762_,
		_w4765_,
		_w4761_,
		_w4766_
	);
	LUT2 #(
		.INIT('h4)
	) name3417 (
		_w4759_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h8)
	) name3418 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w3054_,
		_w4768_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3419 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w3054_,
		_w3056_,
		_w4769_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3420 (
		_w1945_,
		_w4756_,
		_w4767_,
		_w4769_,
		_w4770_
	);
	LUT3 #(
		.INIT('h02)
	) name3421 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2103_,
		_w2172_,
		_w4771_
	);
	LUT4 #(
		.INIT('h2000)
	) name3422 (
		_w2956_,
		_w4051_,
		_w4054_,
		_w4056_,
		_w4772_
	);
	LUT4 #(
		.INIT('h4888)
	) name3423 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w2707_,
		_w2893_,
		_w4773_
	);
	LUT4 #(
		.INIT('h4800)
	) name3424 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2898_,
		_w4773_,
		_w4774_
	);
	LUT4 #(
		.INIT('h8222)
	) name3425 (
		_w2755_,
		_w2961_,
		_w4772_,
		_w4774_,
		_w4775_
	);
	LUT2 #(
		.INIT('h4)
	) name3426 (
		_w2881_,
		_w2892_,
		_w4776_
	);
	LUT4 #(
		.INIT('h0100)
	) name3427 (
		_w2876_,
		_w2878_,
		_w2883_,
		_w4067_,
		_w4777_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		_w2902_,
		_w4075_,
		_w4778_
	);
	LUT4 #(
		.INIT('h8000)
	) name3429 (
		_w4074_,
		_w4776_,
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT4 #(
		.INIT('h4554)
	) name3430 (
		_w2173_,
		_w2755_,
		_w2907_,
		_w4779_,
		_w4780_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3431 (
		_w2171_,
		_w4771_,
		_w4775_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('h13)
	) name3432 (
		_w3032_,
		_w3034_,
		_w4089_,
		_w4782_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3433 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2181_,
		_w3032_,
		_w4089_,
		_w4783_
	);
	LUT3 #(
		.INIT('he0)
	) name3434 (
		_w2108_,
		_w2115_,
		_w2116_,
		_w4784_
	);
	LUT3 #(
		.INIT('h0e)
	) name3435 (
		_w2112_,
		_w2137_,
		_w2175_,
		_w4785_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3436 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w2127_,
		_w4784_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h4)
	) name3437 (
		_w2117_,
		_w2961_,
		_w4787_
	);
	LUT4 #(
		.INIT('he000)
	) name3438 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3034_,
		_w4788_
	);
	LUT4 #(
		.INIT('h004f)
	) name3439 (
		_w2073_,
		_w2086_,
		_w2907_,
		_w4788_,
		_w4789_
	);
	LUT3 #(
		.INIT('h10)
	) name3440 (
		_w4787_,
		_w4786_,
		_w4789_,
		_w4790_
	);
	LUT3 #(
		.INIT('hb0)
	) name3441 (
		_w4782_,
		_w4783_,
		_w4790_,
		_w4791_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3442 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w3054_,
		_w3056_,
		_w4792_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3443 (
		_w1945_,
		_w4781_,
		_w4791_,
		_w4792_,
		_w4793_
	);
	LUT4 #(
		.INIT('h8000)
	) name3444 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4225_,
		_w4227_,
		_w4234_,
		_w4794_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3445 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4225_,
		_w4227_,
		_w4234_,
		_w4795_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3446 (
		_w4236_,
		_w4201_,
		_w4221_,
		_w4224_,
		_w4796_
	);
	LUT4 #(
		.INIT('h1555)
	) name3447 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4215_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w4232_,
		_w4797_,
		_w4798_
	);
	LUT3 #(
		.INIT('h04)
	) name3449 (
		_w4232_,
		_w4234_,
		_w4797_,
		_w4799_
	);
	LUT3 #(
		.INIT('h15)
	) name3450 (
		_w4795_,
		_w4796_,
		_w4799_,
		_w4800_
	);
	LUT3 #(
		.INIT('h0d)
	) name3451 (
		_w4116_,
		_w4167_,
		_w4172_,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name3452 (
		_w4199_,
		_w4155_,
		_w4802_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3453 (
		_w4141_,
		_w4169_,
		_w4801_,
		_w4802_,
		_w4803_
	);
	LUT3 #(
		.INIT('h0b)
	) name3454 (
		_w4199_,
		_w4171_,
		_w4219_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name3455 (
		_w4222_,
		_w4187_,
		_w4805_
	);
	LUT3 #(
		.INIT('h54)
	) name3456 (
		_w4222_,
		_w4217_,
		_w4218_,
		_w4806_
	);
	LUT4 #(
		.INIT('h004f)
	) name3457 (
		_w4803_,
		_w4804_,
		_w4805_,
		_w4806_,
		_w4807_
	);
	LUT3 #(
		.INIT('h04)
	) name3458 (
		_w4232_,
		_w4233_,
		_w4797_,
		_w4808_
	);
	LUT3 #(
		.INIT('h48)
	) name3459 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4236_,
		_w4215_,
		_w4809_
	);
	LUT4 #(
		.INIT('h0400)
	) name3460 (
		_w4232_,
		_w4233_,
		_w4797_,
		_w4809_,
		_w4810_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name3461 (
		_w4214_,
		_w4241_,
		_w4807_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h4)
	) name3462 (
		_w4800_,
		_w4811_,
		_w4812_
	);
	LUT3 #(
		.INIT('h0d)
	) name3463 (
		_w4292_,
		_w4301_,
		_w4306_,
		_w4813_
	);
	LUT3 #(
		.INIT('h70)
	) name3464 (
		_w4296_,
		_w4303_,
		_w4813_,
		_w4814_
	);
	LUT4 #(
		.INIT('h2033)
	) name3465 (
		_w4296_,
		_w4299_,
		_w4303_,
		_w4813_,
		_w4815_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		_w4305_,
		_w4310_,
		_w4816_
	);
	LUT3 #(
		.INIT('h0b)
	) name3467 (
		_w4284_,
		_w4309_,
		_w4313_,
		_w4817_
	);
	LUT4 #(
		.INIT('h7500)
	) name3468 (
		_w4290_,
		_w4815_,
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name3469 (
		_w4319_,
		_w4337_,
		_w4819_
	);
	LUT3 #(
		.INIT('h54)
	) name3470 (
		_w4324_,
		_w4326_,
		_w4327_,
		_w4820_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT3 #(
		.INIT('h40)
	) name3472 (
		_w4214_,
		_w4819_,
		_w4820_,
		_w4822_
	);
	LUT4 #(
		.INIT('h4000)
	) name3473 (
		_w4315_,
		_w4323_,
		_w4818_,
		_w4822_,
		_w4823_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3474 (
		_w4289_,
		_w4297_,
		_w4304_,
		_w4307_,
		_w4824_
	);
	LUT3 #(
		.INIT('h10)
	) name3475 (
		_w4313_,
		_w4315_,
		_w4323_,
		_w4825_
	);
	LUT4 #(
		.INIT('hae00)
	) name3476 (
		_w4284_,
		_w4311_,
		_w4824_,
		_w4825_,
		_w4826_
	);
	LUT3 #(
		.INIT('h01)
	) name3477 (
		_w4214_,
		_w4329_,
		_w4331_,
		_w4827_
	);
	LUT3 #(
		.INIT('h70)
	) name3478 (
		_w4821_,
		_w4826_,
		_w4827_,
		_w4828_
	);
	LUT3 #(
		.INIT('h0b)
	) name3479 (
		_w4332_,
		_w4823_,
		_w4828_,
		_w4829_
	);
	LUT4 #(
		.INIT('h4744)
	) name3480 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w1661_,
		_w4812_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h6)
	) name3481 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4410_,
		_w4831_
	);
	LUT3 #(
		.INIT('h20)
	) name3482 (
		_w4236_,
		_w4401_,
		_w4403_,
		_w4832_
	);
	LUT3 #(
		.INIT('h6a)
	) name3483 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w4238_,
		_w4406_,
		_w4833_
	);
	LUT4 #(
		.INIT('h4888)
	) name3484 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w4238_,
		_w4406_,
		_w4834_
	);
	LUT2 #(
		.INIT('h8)
	) name3485 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4406_,
		_w4835_
	);
	LUT2 #(
		.INIT('h6)
	) name3486 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w4406_,
		_w4836_
	);
	LUT3 #(
		.INIT('h48)
	) name3487 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4406_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		_w4834_,
		_w4837_,
		_w4838_
	);
	LUT3 #(
		.INIT('h40)
	) name3489 (
		_w4400_,
		_w4832_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h4000)
	) name3490 (
		_w4400_,
		_w4831_,
		_w4832_,
		_w4838_,
		_w4840_
	);
	LUT4 #(
		.INIT('h2333)
	) name3491 (
		_w4400_,
		_w4831_,
		_w4832_,
		_w4838_,
		_w4841_
	);
	LUT3 #(
		.INIT('h02)
	) name3492 (
		_w1659_,
		_w4841_,
		_w4840_,
		_w4842_
	);
	LUT4 #(
		.INIT('h00c8)
	) name3493 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w4410_,
		_w4843_
	);
	LUT3 #(
		.INIT('h04)
	) name3494 (
		_w1626_,
		_w1643_,
		_w1667_,
		_w4844_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name3495 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w1658_,
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT3 #(
		.INIT('hb0)
	) name3496 (
		_w1571_,
		_w1583_,
		_w4332_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		_w1640_,
		_w4831_,
		_w4847_
	);
	LUT3 #(
		.INIT('h0b)
	) name3498 (
		_w1617_,
		_w4795_,
		_w4847_,
		_w4848_
	);
	LUT3 #(
		.INIT('h10)
	) name3499 (
		_w4845_,
		_w4846_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h4)
	) name3500 (
		_w4842_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3501 (
		_w1559_,
		_w1678_,
		_w4830_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3502 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w2286_,
		_w4441_,
		_w4852_
	);
	LUT2 #(
		.INIT('hb)
	) name3503 (
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT3 #(
		.INIT('h08)
	) name3504 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1592_,
		_w1660_,
		_w4854_
	);
	LUT4 #(
		.INIT('h4000)
	) name3505 (
		_w4315_,
		_w4325_,
		_w4338_,
		_w4818_,
		_w4855_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name3506 (
		_w4348_,
		_w4349_,
		_w4351_,
		_w4855_,
		_w4856_
	);
	LUT4 #(
		.INIT('h1555)
	) name3507 (
		_w4214_,
		_w4348_,
		_w4352_,
		_w4855_,
		_w4857_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		_w4252_,
		_w4240_,
		_w4858_
	);
	LUT3 #(
		.INIT('h80)
	) name3509 (
		_w4252_,
		_w4240_,
		_w4250_,
		_w4859_
	);
	LUT3 #(
		.INIT('h40)
	) name3510 (
		_w4807_,
		_w4810_,
		_w4859_,
		_w4860_
	);
	LUT3 #(
		.INIT('h48)
	) name3511 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w4255_,
		_w4861_
	);
	LUT4 #(
		.INIT('h4000)
	) name3512 (
		_w4807_,
		_w4810_,
		_w4859_,
		_w4861_,
		_w4862_
	);
	LUT4 #(
		.INIT('h1551)
	) name3513 (
		_w1661_,
		_w4214_,
		_w4264_,
		_w4862_,
		_w4863_
	);
	LUT4 #(
		.INIT('h1055)
	) name3514 (
		_w4854_,
		_w4856_,
		_w4857_,
		_w4863_,
		_w4864_
	);
	LUT3 #(
		.INIT('h6a)
	) name3515 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4252_,
		_w4410_,
		_w4865_
	);
	LUT4 #(
		.INIT('haa02)
	) name3516 (
		_w4386_,
		_w4387_,
		_w4391_,
		_w4393_,
		_w4866_
	);
	LUT2 #(
		.INIT('h1)
	) name3517 (
		_w4392_,
		_w4397_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w4376_,
		_w4396_,
		_w4868_
	);
	LUT4 #(
		.INIT('h7500)
	) name3519 (
		_w4381_,
		_w4866_,
		_w4867_,
		_w4868_,
		_w4869_
	);
	LUT3 #(
		.INIT('h08)
	) name3520 (
		_w4405_,
		_w4409_,
		_w4869_,
		_w4870_
	);
	LUT3 #(
		.INIT('h80)
	) name3521 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w4245_,
		_w4411_,
		_w4871_
	);
	LUT4 #(
		.INIT('h0800)
	) name3522 (
		_w4405_,
		_w4409_,
		_w4869_,
		_w4871_,
		_w4872_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3523 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4252_,
		_w4410_,
		_w4873_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		_w4260_,
		_w4873_,
		_w4874_
	);
	LUT4 #(
		.INIT('h1555)
	) name3525 (
		_w4420_,
		_w4865_,
		_w4872_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h8)
	) name3526 (
		_w4263_,
		_w4873_,
		_w4876_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3527 (
		_w1659_,
		_w4865_,
		_w4872_,
		_w4876_,
		_w4877_
	);
	LUT4 #(
		.INIT('h1222)
	) name3528 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1605_,
		_w4255_,
		_w4260_,
		_w4878_
	);
	LUT4 #(
		.INIT('h6555)
	) name3529 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1605_,
		_w4255_,
		_w4260_,
		_w4879_
	);
	LUT4 #(
		.INIT('h00ec)
	) name3530 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w4879_,
		_w4880_
	);
	LUT3 #(
		.INIT('ha8)
	) name3531 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1605_,
		_w1611_,
		_w4881_
	);
	LUT3 #(
		.INIT('h0b)
	) name3532 (
		_w1611_,
		_w4878_,
		_w4881_,
		_w4882_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3533 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w4882_,
		_w4883_
	);
	LUT3 #(
		.INIT('h54)
	) name3534 (
		_w1602_,
		_w4880_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		_w1640_,
		_w4420_,
		_w4885_
	);
	LUT3 #(
		.INIT('hb0)
	) name3536 (
		_w1571_,
		_w1583_,
		_w4351_,
		_w4886_
	);
	LUT4 #(
		.INIT('haa8a)
	) name3537 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		_w1626_,
		_w1643_,
		_w1667_,
		_w4887_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		_w1563_,
		_w4264_,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w4887_,
		_w4888_,
		_w4889_
	);
	LUT4 #(
		.INIT('h0100)
	) name3540 (
		_w4886_,
		_w4884_,
		_w4885_,
		_w4889_,
		_w4890_
	);
	LUT3 #(
		.INIT('hb0)
	) name3541 (
		_w4875_,
		_w4877_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3542 (
		_w1559_,
		_w1678_,
		_w4864_,
		_w4891_,
		_w4892_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3543 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2286_,
		_w4441_,
		_w4893_
	);
	LUT2 #(
		.INIT('hb)
	) name3544 (
		_w4892_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('h6)
	) name3545 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4269_,
		_w4895_
	);
	LUT4 #(
		.INIT('h8000)
	) name3546 (
		_w4252_,
		_w4240_,
		_w4249_,
		_w4808_,
		_w4896_
	);
	LUT2 #(
		.INIT('h8)
	) name3547 (
		_w4796_,
		_w4896_,
		_w4897_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name3548 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w4255_,
		_w4248_,
		_w4898_
	);
	LUT3 #(
		.INIT('h80)
	) name3549 (
		_w4260_,
		_w4265_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name3550 (
		_w4271_,
		_w4899_,
		_w4900_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3551 (
		_w4214_,
		_w4796_,
		_w4896_,
		_w4900_,
		_w4901_
	);
	LUT4 #(
		.INIT('hf800)
	) name3552 (
		_w4267_,
		_w4270_,
		_w4895_,
		_w4901_,
		_w4902_
	);
	LUT3 #(
		.INIT('h04)
	) name3553 (
		_w4315_,
		_w4323_,
		_w4324_,
		_w4903_
	);
	LUT3 #(
		.INIT('h02)
	) name3554 (
		_w4333_,
		_w4336_,
		_w4361_,
		_w4904_
	);
	LUT3 #(
		.INIT('h80)
	) name3555 (
		_w4348_,
		_w4358_,
		_w4904_,
		_w4905_
	);
	LUT4 #(
		.INIT('h8000)
	) name3556 (
		_w4818_,
		_w4819_,
		_w4903_,
		_w4905_,
		_w4906_
	);
	LUT3 #(
		.INIT('h14)
	) name3557 (
		_w4214_,
		_w4360_,
		_w4906_,
		_w4907_
	);
	LUT4 #(
		.INIT('h4447)
	) name3558 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1661_,
		_w4902_,
		_w4907_,
		_w4908_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3559 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4262_,
		_w4419_,
		_w4909_
	);
	LUT3 #(
		.INIT('h80)
	) name3560 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4262_,
		_w4420_,
		_w4910_
	);
	LUT4 #(
		.INIT('h8000)
	) name3561 (
		_w4865_,
		_w4872_,
		_w4874_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h6)
	) name3562 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4419_,
		_w4912_
	);
	LUT3 #(
		.INIT('h6c)
	) name3563 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4419_,
		_w4913_
	);
	LUT2 #(
		.INIT('h8)
	) name3564 (
		_w4429_,
		_w4913_,
		_w4914_
	);
	LUT3 #(
		.INIT('h80)
	) name3565 (
		_w4429_,
		_w4912_,
		_w4913_,
		_w4915_
	);
	LUT4 #(
		.INIT('h8000)
	) name3566 (
		_w4865_,
		_w4872_,
		_w4876_,
		_w4915_,
		_w4916_
	);
	LUT4 #(
		.INIT('h00a8)
	) name3567 (
		_w1659_,
		_w4909_,
		_w4911_,
		_w4916_,
		_w4917_
	);
	LUT3 #(
		.INIT('h54)
	) name3568 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1592_,
		_w1595_,
		_w4918_
	);
	LUT4 #(
		.INIT('h00c8)
	) name3569 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w4918_,
		_w4919_
	);
	LUT3 #(
		.INIT('hd0)
	) name3570 (
		_w1596_,
		_w4909_,
		_w4919_,
		_w4920_
	);
	LUT3 #(
		.INIT('h21)
	) name3571 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1605_,
		_w4269_,
		_w4921_
	);
	LUT3 #(
		.INIT('h40)
	) name3572 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w4922_
	);
	LUT4 #(
		.INIT('h0031)
	) name3573 (
		_w1604_,
		_w1602_,
		_w1616_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h4)
	) name3574 (
		_w4921_,
		_w4923_,
		_w4924_
	);
	LUT3 #(
		.INIT('hb0)
	) name3575 (
		_w1571_,
		_w1583_,
		_w4360_,
		_w4925_
	);
	LUT4 #(
		.INIT('h008b)
	) name3576 (
		_w1569_,
		_w1602_,
		_w1613_,
		_w1667_,
		_w4926_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3577 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w1602_,
		_w4927_
	);
	LUT4 #(
		.INIT('h4a48)
	) name3578 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w1563_,
		_w4269_,
		_w4927_,
		_w4928_
	);
	LUT3 #(
		.INIT('h0d)
	) name3579 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		_w4926_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('h0100)
	) name3580 (
		_w4925_,
		_w4920_,
		_w4924_,
		_w4929_,
		_w4930_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3581 (
		_w1559_,
		_w4908_,
		_w4917_,
		_w4930_,
		_w4931_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3582 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2286_,
		_w4441_,
		_w4932_
	);
	LUT3 #(
		.INIT('h2f)
	) name3583 (
		_w1678_,
		_w4931_,
		_w4932_,
		_w4933_
	);
	LUT3 #(
		.INIT('h08)
	) name3584 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w1842_,
		_w1915_,
		_w4934_
	);
	LUT3 #(
		.INIT('h41)
	) name3585 (
		_w3101_,
		_w3252_,
		_w4729_,
		_w4935_
	);
	LUT4 #(
		.INIT('h007f)
	) name3586 (
		_w4463_,
		_w4465_,
		_w4467_,
		_w4448_,
		_w4936_
	);
	LUT4 #(
		.INIT('h1115)
	) name3587 (
		_w1916_,
		_w3101_,
		_w3996_,
		_w4936_,
		_w4937_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3588 (
		_w1810_,
		_w4934_,
		_w4935_,
		_w4937_,
		_w4938_
	);
	LUT4 #(
		.INIT('h2888)
	) name3589 (
		_w1924_,
		_w4016_,
		_w4029_,
		_w4735_,
		_w4939_
	);
	LUT4 #(
		.INIT('h8444)
	) name3590 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w1920_,
		_w3072_,
		_w3074_,
		_w4940_
	);
	LUT2 #(
		.INIT('h2)
	) name3591 (
		_w4739_,
		_w4940_,
		_w4941_
	);
	LUT3 #(
		.INIT('ha2)
	) name3592 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w4037_,
		_w4941_,
		_w4942_
	);
	LUT3 #(
		.INIT('h40)
	) name3593 (
		_w1846_,
		_w3074_,
		_w3366_,
		_w4943_
	);
	LUT3 #(
		.INIT('h04)
	) name3594 (
		_w1833_,
		_w4016_,
		_w4943_,
		_w4944_
	);
	LUT3 #(
		.INIT('h80)
	) name3595 (
		_w1805_,
		_w1806_,
		_w4448_,
		_w4945_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name3596 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		_w1861_,
		_w3072_,
		_w3074_,
		_w4946_
	);
	LUT4 #(
		.INIT('h010f)
	) name3597 (
		_w1855_,
		_w1860_,
		_w4945_,
		_w4946_,
		_w4947_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3598 (
		_w1816_,
		_w1831_,
		_w3252_,
		_w4947_,
		_w4948_
	);
	LUT3 #(
		.INIT('h10)
	) name3599 (
		_w4942_,
		_w4944_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h4)
	) name3600 (
		_w4939_,
		_w4949_,
		_w4950_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3601 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w3406_,
		_w3408_,
		_w4951_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3602 (
		_w1933_,
		_w4938_,
		_w4950_,
		_w4951_,
		_w4952_
	);
	LUT4 #(
		.INIT('hffeb)
	) name3603 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w4953_
	);
	LUT3 #(
		.INIT('h02)
	) name3604 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w3534_,
		_w3536_,
		_w4954_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3605 (
		_w3537_,
		_w3426_,
		_w3427_,
		_w4954_,
		_w4955_
	);
	LUT3 #(
		.INIT('h08)
	) name3606 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3413_,
		_w4956_
	);
	LUT3 #(
		.INIT('h0e)
	) name3607 (
		_w4953_,
		_w4955_,
		_w4956_,
		_w4957_
	);
	LUT3 #(
		.INIT('h82)
	) name3608 (
		_w3411_,
		_w3523_,
		_w3526_,
		_w4958_
	);
	LUT4 #(
		.INIT('h5655)
	) name3609 (
		_w3486_,
		_w3489_,
		_w3493_,
		_w3531_,
		_w4959_
	);
	LUT3 #(
		.INIT('hc4)
	) name3610 (
		_w3407_,
		_w3414_,
		_w4955_,
		_w4960_
	);
	LUT3 #(
		.INIT('hb0)
	) name3611 (
		_w3411_,
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h2)
	) name3612 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w3545_,
		_w4962_
	);
	LUT4 #(
		.INIT('hc055)
	) name3613 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3534_,
		_w4963_
	);
	LUT3 #(
		.INIT('h31)
	) name3614 (
		_w2248_,
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3615 (
		_w4957_,
		_w4958_,
		_w4961_,
		_w4964_,
		_w4965_
	);
	LUT4 #(
		.INIT('hc444)
	) name3616 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4966_
	);
	LUT4 #(
		.INIT('h0888)
	) name3617 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[30]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name3618 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT3 #(
		.INIT('ha8)
	) name3619 (
		_w2250_,
		_w4966_,
		_w4967_,
		_w4969_
	);
	LUT4 #(
		.INIT('hc444)
	) name3620 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[22]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4970_
	);
	LUT4 #(
		.INIT('h0888)
	) name3621 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[22]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4971_
	);
	LUT2 #(
		.INIT('h1)
	) name3622 (
		_w4970_,
		_w4971_,
		_w4972_
	);
	LUT3 #(
		.INIT('ha8)
	) name3623 (
		_w2264_,
		_w4970_,
		_w4971_,
		_w4973_
	);
	LUT3 #(
		.INIT('ha8)
	) name3624 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w4969_,
		_w4973_,
		_w4974_
	);
	LUT4 #(
		.INIT('hc444)
	) name3625 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4975_
	);
	LUT4 #(
		.INIT('h0888)
	) name3626 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[6]/NET0131 ,
		_w2255_,
		_w2260_,
		_w4976_
	);
	LUT2 #(
		.INIT('h1)
	) name3627 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT3 #(
		.INIT('h02)
	) name3628 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w2271_,
		_w2272_,
		_w4978_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3629 (
		_w2273_,
		_w4975_,
		_w4976_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		_w2280_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('ha8)
	) name3631 (
		_w1679_,
		_w4974_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h2)
	) name3632 (
		_w2283_,
		_w4979_,
		_w4982_
	);
	LUT4 #(
		.INIT('hc055)
	) name3633 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2272_,
		_w4983_
	);
	LUT2 #(
		.INIT('h2)
	) name3634 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		_w2288_,
		_w4984_
	);
	LUT3 #(
		.INIT('h0d)
	) name3635 (
		_w2246_,
		_w4983_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h4)
	) name3636 (
		_w4982_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('hb)
	) name3637 (
		_w4981_,
		_w4986_,
		_w4987_
	);
	LUT3 #(
		.INIT('h02)
	) name3638 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w3578_,
		_w3580_,
		_w4988_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3639 (
		_w3426_,
		_w3427_,
		_w3581_,
		_w4988_,
		_w4989_
	);
	LUT3 #(
		.INIT('h08)
	) name3640 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3574_,
		_w4990_
	);
	LUT3 #(
		.INIT('h0e)
	) name3641 (
		_w4953_,
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT3 #(
		.INIT('h90)
	) name3642 (
		_w3523_,
		_w3526_,
		_w3572_,
		_w4992_
	);
	LUT3 #(
		.INIT('hc4)
	) name3643 (
		_w3407_,
		_w3575_,
		_w4989_,
		_w4993_
	);
	LUT3 #(
		.INIT('hb0)
	) name3644 (
		_w3572_,
		_w4959_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h2)
	) name3645 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w3545_,
		_w4995_
	);
	LUT4 #(
		.INIT('hc055)
	) name3646 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3578_,
		_w4996_
	);
	LUT3 #(
		.INIT('h31)
	) name3647 (
		_w2248_,
		_w4995_,
		_w4996_,
		_w4997_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3648 (
		_w4991_,
		_w4992_,
		_w4994_,
		_w4997_,
		_w4998_
	);
	LUT3 #(
		.INIT('h02)
	) name3649 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		_w3536_,
		_w3412_,
		_w4999_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3650 (
		_w3426_,
		_w3427_,
		_w3597_,
		_w4999_,
		_w5000_
	);
	LUT3 #(
		.INIT('h08)
	) name3651 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3593_,
		_w5001_
	);
	LUT3 #(
		.INIT('h0e)
	) name3652 (
		_w4953_,
		_w5000_,
		_w5001_,
		_w5002_
	);
	LUT3 #(
		.INIT('h90)
	) name3653 (
		_w3523_,
		_w3526_,
		_w3592_,
		_w5003_
	);
	LUT3 #(
		.INIT('hc4)
	) name3654 (
		_w3407_,
		_w3594_,
		_w5000_,
		_w5004_
	);
	LUT3 #(
		.INIT('hb0)
	) name3655 (
		_w3592_,
		_w4959_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h2)
	) name3656 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		_w3545_,
		_w5006_
	);
	LUT4 #(
		.INIT('hc055)
	) name3657 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3536_,
		_w5007_
	);
	LUT3 #(
		.INIT('h31)
	) name3658 (
		_w2248_,
		_w5006_,
		_w5007_,
		_w5008_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3659 (
		_w5002_,
		_w5003_,
		_w5005_,
		_w5008_,
		_w5009_
	);
	LUT3 #(
		.INIT('h02)
	) name3660 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w3534_,
		_w3611_,
		_w5010_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3661 (
		_w3426_,
		_w3427_,
		_w3612_,
		_w5010_,
		_w5011_
	);
	LUT3 #(
		.INIT('h08)
	) name3662 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3597_,
		_w5012_
	);
	LUT3 #(
		.INIT('h0e)
	) name3663 (
		_w4953_,
		_w5011_,
		_w5012_,
		_w5013_
	);
	LUT3 #(
		.INIT('h82)
	) name3664 (
		_w3412_,
		_w3523_,
		_w3526_,
		_w5014_
	);
	LUT3 #(
		.INIT('hc4)
	) name3665 (
		_w3407_,
		_w3608_,
		_w5011_,
		_w5015_
	);
	LUT3 #(
		.INIT('hb0)
	) name3666 (
		_w3412_,
		_w4959_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h2)
	) name3667 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w3545_,
		_w5017_
	);
	LUT4 #(
		.INIT('hc055)
	) name3668 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3611_,
		_w5018_
	);
	LUT3 #(
		.INIT('h31)
	) name3669 (
		_w2248_,
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3670 (
		_w5013_,
		_w5014_,
		_w5016_,
		_w5019_,
		_w5020_
	);
	LUT3 #(
		.INIT('h02)
	) name3671 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w3572_,
		_w3611_,
		_w5021_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3672 (
		_w3426_,
		_w3427_,
		_w3626_,
		_w5021_,
		_w5022_
	);
	LUT3 #(
		.INIT('h08)
	) name3673 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3537_,
		_w5023_
	);
	LUT3 #(
		.INIT('h0e)
	) name3674 (
		_w4953_,
		_w5022_,
		_w5023_,
		_w5024_
	);
	LUT3 #(
		.INIT('h82)
	) name3675 (
		_w3536_,
		_w3523_,
		_w3526_,
		_w5025_
	);
	LUT3 #(
		.INIT('hc4)
	) name3676 (
		_w3407_,
		_w3623_,
		_w5022_,
		_w5026_
	);
	LUT3 #(
		.INIT('hb0)
	) name3677 (
		_w3536_,
		_w4959_,
		_w5026_,
		_w5027_
	);
	LUT2 #(
		.INIT('h2)
	) name3678 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w3545_,
		_w5028_
	);
	LUT4 #(
		.INIT('hc055)
	) name3679 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3572_,
		_w5029_
	);
	LUT3 #(
		.INIT('h31)
	) name3680 (
		_w2248_,
		_w5028_,
		_w5029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3681 (
		_w5024_,
		_w5025_,
		_w5027_,
		_w5030_,
		_w5031_
	);
	LUT3 #(
		.INIT('h02)
	) name3682 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w3572_,
		_w3573_,
		_w5032_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3683 (
		_w3426_,
		_w3427_,
		_w3574_,
		_w5032_,
		_w5033_
	);
	LUT3 #(
		.INIT('h08)
	) name3684 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3612_,
		_w5034_
	);
	LUT3 #(
		.INIT('h0e)
	) name3685 (
		_w4953_,
		_w5033_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('h82)
	) name3686 (
		_w3534_,
		_w3523_,
		_w3526_,
		_w5036_
	);
	LUT3 #(
		.INIT('hc4)
	) name3687 (
		_w3407_,
		_w3637_,
		_w5033_,
		_w5037_
	);
	LUT3 #(
		.INIT('hb0)
	) name3688 (
		_w3534_,
		_w4959_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h2)
	) name3689 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w3545_,
		_w5039_
	);
	LUT4 #(
		.INIT('hc055)
	) name3690 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3573_,
		_w5040_
	);
	LUT3 #(
		.INIT('h31)
	) name3691 (
		_w2248_,
		_w5039_,
		_w5040_,
		_w5041_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3692 (
		_w5035_,
		_w5036_,
		_w5038_,
		_w5041_,
		_w5042_
	);
	LUT3 #(
		.INIT('h02)
	) name3693 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w3580_,
		_w3573_,
		_w5043_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3694 (
		_w3426_,
		_w3427_,
		_w3653_,
		_w5043_,
		_w5044_
	);
	LUT3 #(
		.INIT('h08)
	) name3695 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3626_,
		_w5045_
	);
	LUT3 #(
		.INIT('h0e)
	) name3696 (
		_w4953_,
		_w5044_,
		_w5045_,
		_w5046_
	);
	LUT3 #(
		.INIT('h90)
	) name3697 (
		_w3523_,
		_w3526_,
		_w3611_,
		_w5047_
	);
	LUT3 #(
		.INIT('hc4)
	) name3698 (
		_w3407_,
		_w3650_,
		_w5044_,
		_w5048_
	);
	LUT3 #(
		.INIT('hb0)
	) name3699 (
		_w3611_,
		_w4959_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h2)
	) name3700 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w3545_,
		_w5050_
	);
	LUT4 #(
		.INIT('hc055)
	) name3701 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3580_,
		_w5051_
	);
	LUT3 #(
		.INIT('h31)
	) name3702 (
		_w2248_,
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3703 (
		_w5046_,
		_w5047_,
		_w5049_,
		_w5052_,
		_w5053_
	);
	LUT3 #(
		.INIT('h02)
	) name3704 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w3578_,
		_w3667_,
		_w5054_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3705 (
		_w3426_,
		_w3427_,
		_w3668_,
		_w5054_,
		_w5055_
	);
	LUT3 #(
		.INIT('h08)
	) name3706 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3653_,
		_w5056_
	);
	LUT3 #(
		.INIT('h0e)
	) name3707 (
		_w4953_,
		_w5055_,
		_w5056_,
		_w5057_
	);
	LUT3 #(
		.INIT('h90)
	) name3708 (
		_w3523_,
		_w3526_,
		_w3573_,
		_w5058_
	);
	LUT3 #(
		.INIT('hc4)
	) name3709 (
		_w3407_,
		_w3664_,
		_w5055_,
		_w5059_
	);
	LUT3 #(
		.INIT('hb0)
	) name3710 (
		_w3573_,
		_w4959_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w3545_,
		_w5061_
	);
	LUT4 #(
		.INIT('hc055)
	) name3712 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3667_,
		_w5062_
	);
	LUT3 #(
		.INIT('h31)
	) name3713 (
		_w2248_,
		_w5061_,
		_w5062_,
		_w5063_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3714 (
		_w5057_,
		_w5058_,
		_w5060_,
		_w5063_,
		_w5064_
	);
	LUT3 #(
		.INIT('h02)
	) name3715 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w3667_,
		_w3683_,
		_w5065_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3716 (
		_w3426_,
		_w3427_,
		_w3698_,
		_w5065_,
		_w5066_
	);
	LUT3 #(
		.INIT('h08)
	) name3717 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3581_,
		_w5067_
	);
	LUT3 #(
		.INIT('h0e)
	) name3718 (
		_w4953_,
		_w5066_,
		_w5067_,
		_w5068_
	);
	LUT3 #(
		.INIT('h90)
	) name3719 (
		_w3523_,
		_w3526_,
		_w3580_,
		_w5069_
	);
	LUT3 #(
		.INIT('hc4)
	) name3720 (
		_w3407_,
		_w3695_,
		_w5066_,
		_w5070_
	);
	LUT3 #(
		.INIT('hb0)
	) name3721 (
		_w3580_,
		_w4959_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h2)
	) name3722 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w3545_,
		_w5072_
	);
	LUT4 #(
		.INIT('hc055)
	) name3723 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3683_,
		_w5073_
	);
	LUT3 #(
		.INIT('h31)
	) name3724 (
		_w2248_,
		_w5072_,
		_w5073_,
		_w5074_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3725 (
		_w5068_,
		_w5069_,
		_w5071_,
		_w5074_,
		_w5075_
	);
	LUT3 #(
		.INIT('h02)
	) name3726 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w3682_,
		_w3683_,
		_w5076_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3727 (
		_w3426_,
		_w3427_,
		_w3684_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h08)
	) name3728 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3668_,
		_w5078_
	);
	LUT3 #(
		.INIT('h0e)
	) name3729 (
		_w4953_,
		_w5077_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('h90)
	) name3730 (
		_w3523_,
		_w3526_,
		_w3578_,
		_w5080_
	);
	LUT3 #(
		.INIT('hc4)
	) name3731 (
		_w3407_,
		_w3679_,
		_w5077_,
		_w5081_
	);
	LUT3 #(
		.INIT('hb0)
	) name3732 (
		_w3578_,
		_w4959_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h2)
	) name3733 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w3545_,
		_w5083_
	);
	LUT4 #(
		.INIT('hc055)
	) name3734 (
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3682_,
		_w5084_
	);
	LUT3 #(
		.INIT('h31)
	) name3735 (
		_w2248_,
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3736 (
		_w5079_,
		_w5080_,
		_w5082_,
		_w5085_,
		_w5086_
	);
	LUT3 #(
		.INIT('h02)
	) name3737 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w3682_,
		_w3712_,
		_w5087_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3738 (
		_w3426_,
		_w3427_,
		_w3713_,
		_w5087_,
		_w5088_
	);
	LUT3 #(
		.INIT('h08)
	) name3739 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3698_,
		_w5089_
	);
	LUT3 #(
		.INIT('h0e)
	) name3740 (
		_w4953_,
		_w5088_,
		_w5089_,
		_w5090_
	);
	LUT3 #(
		.INIT('h90)
	) name3741 (
		_w3523_,
		_w3526_,
		_w3667_,
		_w5091_
	);
	LUT3 #(
		.INIT('hc4)
	) name3742 (
		_w3407_,
		_w3709_,
		_w5088_,
		_w5092_
	);
	LUT3 #(
		.INIT('hb0)
	) name3743 (
		_w3667_,
		_w4959_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h2)
	) name3744 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w3545_,
		_w5094_
	);
	LUT4 #(
		.INIT('hc055)
	) name3745 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3712_,
		_w5095_
	);
	LUT3 #(
		.INIT('h31)
	) name3746 (
		_w2248_,
		_w5094_,
		_w5095_,
		_w5096_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3747 (
		_w5090_,
		_w5091_,
		_w5093_,
		_w5096_,
		_w5097_
	);
	LUT3 #(
		.INIT('h02)
	) name3748 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w3712_,
		_w3727_,
		_w5098_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3749 (
		_w3426_,
		_w3427_,
		_w3728_,
		_w5098_,
		_w5099_
	);
	LUT3 #(
		.INIT('h08)
	) name3750 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3684_,
		_w5100_
	);
	LUT3 #(
		.INIT('h0e)
	) name3751 (
		_w4953_,
		_w5099_,
		_w5100_,
		_w5101_
	);
	LUT3 #(
		.INIT('h90)
	) name3752 (
		_w3523_,
		_w3526_,
		_w3683_,
		_w5102_
	);
	LUT3 #(
		.INIT('hc4)
	) name3753 (
		_w3407_,
		_w3724_,
		_w5099_,
		_w5103_
	);
	LUT3 #(
		.INIT('hb0)
	) name3754 (
		_w3683_,
		_w4959_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h2)
	) name3755 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w3545_,
		_w5105_
	);
	LUT4 #(
		.INIT('hc055)
	) name3756 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3727_,
		_w5106_
	);
	LUT3 #(
		.INIT('h31)
	) name3757 (
		_w2248_,
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3758 (
		_w5101_,
		_w5102_,
		_w5104_,
		_w5107_,
		_w5108_
	);
	LUT3 #(
		.INIT('h02)
	) name3759 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w3727_,
		_w3742_,
		_w5109_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3760 (
		_w3426_,
		_w3427_,
		_w3743_,
		_w5109_,
		_w5110_
	);
	LUT3 #(
		.INIT('h08)
	) name3761 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3713_,
		_w5111_
	);
	LUT3 #(
		.INIT('h0e)
	) name3762 (
		_w4953_,
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT3 #(
		.INIT('h90)
	) name3763 (
		_w3523_,
		_w3526_,
		_w3682_,
		_w5113_
	);
	LUT3 #(
		.INIT('hc4)
	) name3764 (
		_w3407_,
		_w3739_,
		_w5110_,
		_w5114_
	);
	LUT3 #(
		.INIT('hb0)
	) name3765 (
		_w3682_,
		_w4959_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h2)
	) name3766 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w3545_,
		_w5116_
	);
	LUT4 #(
		.INIT('hc055)
	) name3767 (
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3742_,
		_w5117_
	);
	LUT3 #(
		.INIT('h31)
	) name3768 (
		_w2248_,
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3769 (
		_w5112_,
		_w5113_,
		_w5115_,
		_w5118_,
		_w5119_
	);
	LUT3 #(
		.INIT('h02)
	) name3770 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w3592_,
		_w3742_,
		_w5120_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3771 (
		_w3426_,
		_w3427_,
		_w3757_,
		_w5120_,
		_w5121_
	);
	LUT3 #(
		.INIT('h08)
	) name3772 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3728_,
		_w5122_
	);
	LUT3 #(
		.INIT('h0e)
	) name3773 (
		_w4953_,
		_w5121_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h90)
	) name3774 (
		_w3523_,
		_w3526_,
		_w3712_,
		_w5124_
	);
	LUT3 #(
		.INIT('hc4)
	) name3775 (
		_w3407_,
		_w3754_,
		_w5121_,
		_w5125_
	);
	LUT3 #(
		.INIT('hb0)
	) name3776 (
		_w3712_,
		_w4959_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h2)
	) name3777 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w3545_,
		_w5127_
	);
	LUT4 #(
		.INIT('hc055)
	) name3778 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3592_,
		_w5128_
	);
	LUT3 #(
		.INIT('h31)
	) name3779 (
		_w2248_,
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3780 (
		_w5123_,
		_w5124_,
		_w5126_,
		_w5129_,
		_w5130_
	);
	LUT3 #(
		.INIT('h02)
	) name3781 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w3411_,
		_w3592_,
		_w5131_
	);
	LUT4 #(
		.INIT('h00f1)
	) name3782 (
		_w3426_,
		_w3427_,
		_w3593_,
		_w5131_,
		_w5132_
	);
	LUT3 #(
		.INIT('h08)
	) name3783 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3743_,
		_w5133_
	);
	LUT3 #(
		.INIT('h0e)
	) name3784 (
		_w4953_,
		_w5132_,
		_w5133_,
		_w5134_
	);
	LUT3 #(
		.INIT('h90)
	) name3785 (
		_w3523_,
		_w3526_,
		_w3727_,
		_w5135_
	);
	LUT3 #(
		.INIT('hc4)
	) name3786 (
		_w3407_,
		_w3768_,
		_w5132_,
		_w5136_
	);
	LUT3 #(
		.INIT('hb0)
	) name3787 (
		_w3727_,
		_w4959_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h2)
	) name3788 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w3545_,
		_w5138_
	);
	LUT4 #(
		.INIT('hc055)
	) name3789 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3411_,
		_w5139_
	);
	LUT3 #(
		.INIT('h31)
	) name3790 (
		_w2248_,
		_w5138_,
		_w5139_,
		_w5140_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3791 (
		_w5134_,
		_w5135_,
		_w5137_,
		_w5140_,
		_w5141_
	);
	LUT3 #(
		.INIT('h02)
	) name3792 (
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w3411_,
		_w3412_,
		_w5142_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3793 (
		_w3413_,
		_w3426_,
		_w3427_,
		_w5142_,
		_w5143_
	);
	LUT3 #(
		.INIT('h08)
	) name3794 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3757_,
		_w5144_
	);
	LUT3 #(
		.INIT('h0e)
	) name3795 (
		_w4953_,
		_w5143_,
		_w5144_,
		_w5145_
	);
	LUT3 #(
		.INIT('h90)
	) name3796 (
		_w3523_,
		_w3526_,
		_w3742_,
		_w5146_
	);
	LUT3 #(
		.INIT('hc4)
	) name3797 (
		_w3407_,
		_w3781_,
		_w5143_,
		_w5147_
	);
	LUT3 #(
		.INIT('hb0)
	) name3798 (
		_w3742_,
		_w4959_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h2)
	) name3799 (
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w3545_,
		_w5149_
	);
	LUT4 #(
		.INIT('hc055)
	) name3800 (
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1731_,
		_w1736_,
		_w3412_,
		_w5150_
	);
	LUT3 #(
		.INIT('h31)
	) name3801 (
		_w2248_,
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3802 (
		_w5145_,
		_w5146_,
		_w5148_,
		_w5151_,
		_w5152_
	);
	LUT3 #(
		.INIT('ha8)
	) name3803 (
		_w2315_,
		_w4966_,
		_w4967_,
		_w5153_
	);
	LUT3 #(
		.INIT('ha8)
	) name3804 (
		_w2317_,
		_w4970_,
		_w4971_,
		_w5154_
	);
	LUT3 #(
		.INIT('ha8)
	) name3805 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5153_,
		_w5154_,
		_w5155_
	);
	LUT3 #(
		.INIT('h02)
	) name3806 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w2320_,
		_w2322_,
		_w5156_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3807 (
		_w2323_,
		_w4975_,
		_w4976_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		_w2327_,
		_w5157_,
		_w5158_
	);
	LUT3 #(
		.INIT('ha8)
	) name3809 (
		_w1679_,
		_w5155_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		_w2283_,
		_w5157_,
		_w5160_
	);
	LUT4 #(
		.INIT('hc055)
	) name3811 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2320_,
		_w5161_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		_w2288_,
		_w5162_
	);
	LUT3 #(
		.INIT('h0d)
	) name3813 (
		_w2246_,
		_w5161_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h4)
	) name3814 (
		_w5160_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('hb)
	) name3815 (
		_w5159_,
		_w5164_,
		_w5165_
	);
	LUT3 #(
		.INIT('ha8)
	) name3816 (
		_w2250_,
		_w4970_,
		_w4971_,
		_w5166_
	);
	LUT3 #(
		.INIT('ha8)
	) name3817 (
		_w2349_,
		_w4966_,
		_w4967_,
		_w5167_
	);
	LUT3 #(
		.INIT('ha8)
	) name3818 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5166_,
		_w5167_,
		_w5168_
	);
	LUT3 #(
		.INIT('h02)
	) name3819 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w2271_,
		_w2264_,
		_w5169_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3820 (
		_w2346_,
		_w4975_,
		_w4976_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name3821 (
		_w2351_,
		_w5170_,
		_w5171_
	);
	LUT3 #(
		.INIT('ha8)
	) name3822 (
		_w1679_,
		_w5168_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h2)
	) name3823 (
		_w2283_,
		_w5170_,
		_w5173_
	);
	LUT4 #(
		.INIT('hc055)
	) name3824 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2271_,
		_w5174_
	);
	LUT2 #(
		.INIT('h2)
	) name3825 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		_w2288_,
		_w5175_
	);
	LUT3 #(
		.INIT('h0d)
	) name3826 (
		_w2246_,
		_w5174_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		_w5173_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('hb)
	) name3828 (
		_w5172_,
		_w5177_,
		_w5178_
	);
	LUT3 #(
		.INIT('ha8)
	) name3829 (
		_w2264_,
		_w4966_,
		_w4967_,
		_w5179_
	);
	LUT3 #(
		.INIT('ha8)
	) name3830 (
		_w2271_,
		_w4970_,
		_w4971_,
		_w5180_
	);
	LUT3 #(
		.INIT('ha8)
	) name3831 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT3 #(
		.INIT('h02)
	) name3832 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w2272_,
		_w2376_,
		_w5182_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3833 (
		_w2377_,
		_w4975_,
		_w4976_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h1)
	) name3834 (
		_w2380_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('ha8)
	) name3835 (
		_w1679_,
		_w5181_,
		_w5184_,
		_w5185_
	);
	LUT2 #(
		.INIT('h2)
	) name3836 (
		_w2283_,
		_w5183_,
		_w5186_
	);
	LUT4 #(
		.INIT('hc055)
	) name3837 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2376_,
		_w5187_
	);
	LUT2 #(
		.INIT('h2)
	) name3838 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		_w2288_,
		_w5188_
	);
	LUT3 #(
		.INIT('h0d)
	) name3839 (
		_w2246_,
		_w5187_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name3840 (
		_w5186_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('hb)
	) name3841 (
		_w5185_,
		_w5190_,
		_w5191_
	);
	LUT3 #(
		.INIT('ha8)
	) name3842 (
		_w2271_,
		_w4966_,
		_w4967_,
		_w5192_
	);
	LUT3 #(
		.INIT('ha8)
	) name3843 (
		_w2272_,
		_w4970_,
		_w4971_,
		_w5193_
	);
	LUT3 #(
		.INIT('ha8)
	) name3844 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5192_,
		_w5193_,
		_w5194_
	);
	LUT3 #(
		.INIT('h02)
	) name3845 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w2315_,
		_w2376_,
		_w5195_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3846 (
		_w2402_,
		_w4975_,
		_w4976_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name3847 (
		_w2405_,
		_w5196_,
		_w5197_
	);
	LUT3 #(
		.INIT('ha8)
	) name3848 (
		_w1679_,
		_w5194_,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name3849 (
		_w2283_,
		_w5196_,
		_w5199_
	);
	LUT4 #(
		.INIT('hc055)
	) name3850 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2315_,
		_w5200_
	);
	LUT2 #(
		.INIT('h2)
	) name3851 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w2288_,
		_w5201_
	);
	LUT3 #(
		.INIT('h0d)
	) name3852 (
		_w2246_,
		_w5200_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h4)
	) name3853 (
		_w5199_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('hb)
	) name3854 (
		_w5198_,
		_w5203_,
		_w5204_
	);
	LUT3 #(
		.INIT('ha8)
	) name3855 (
		_w2272_,
		_w4966_,
		_w4967_,
		_w5205_
	);
	LUT3 #(
		.INIT('ha8)
	) name3856 (
		_w2376_,
		_w4970_,
		_w4971_,
		_w5206_
	);
	LUT3 #(
		.INIT('ha8)
	) name3857 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5205_,
		_w5206_,
		_w5207_
	);
	LUT3 #(
		.INIT('h02)
	) name3858 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w2315_,
		_w2317_,
		_w5208_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3859 (
		_w2326_,
		_w4975_,
		_w4976_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		_w2429_,
		_w5209_,
		_w5210_
	);
	LUT3 #(
		.INIT('ha8)
	) name3861 (
		_w1679_,
		_w5207_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		_w2283_,
		_w5209_,
		_w5212_
	);
	LUT4 #(
		.INIT('hc055)
	) name3863 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2317_,
		_w5213_
	);
	LUT2 #(
		.INIT('h2)
	) name3864 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		_w2288_,
		_w5214_
	);
	LUT3 #(
		.INIT('h0d)
	) name3865 (
		_w2246_,
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h4)
	) name3866 (
		_w5212_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('hb)
	) name3867 (
		_w5211_,
		_w5216_,
		_w5217_
	);
	LUT3 #(
		.INIT('ha8)
	) name3868 (
		_w2376_,
		_w4966_,
		_w4967_,
		_w5218_
	);
	LUT3 #(
		.INIT('ha8)
	) name3869 (
		_w2315_,
		_w4970_,
		_w4971_,
		_w5219_
	);
	LUT3 #(
		.INIT('ha8)
	) name3870 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5218_,
		_w5219_,
		_w5220_
	);
	LUT3 #(
		.INIT('h02)
	) name3871 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w2322_,
		_w2317_,
		_w5221_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3872 (
		_w2451_,
		_w4975_,
		_w4976_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w2454_,
		_w5222_,
		_w5223_
	);
	LUT3 #(
		.INIT('ha8)
	) name3874 (
		_w1679_,
		_w5220_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h2)
	) name3875 (
		_w2283_,
		_w5222_,
		_w5225_
	);
	LUT4 #(
		.INIT('hc055)
	) name3876 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2322_,
		_w5226_
	);
	LUT2 #(
		.INIT('h2)
	) name3877 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w2288_,
		_w5227_
	);
	LUT3 #(
		.INIT('h0d)
	) name3878 (
		_w2246_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		_w5225_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('hb)
	) name3880 (
		_w5224_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('ha8)
	) name3881 (
		_w2317_,
		_w4966_,
		_w4967_,
		_w5231_
	);
	LUT3 #(
		.INIT('ha8)
	) name3882 (
		_w2322_,
		_w4970_,
		_w4971_,
		_w5232_
	);
	LUT3 #(
		.INIT('ha8)
	) name3883 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5231_,
		_w5232_,
		_w5233_
	);
	LUT3 #(
		.INIT('h02)
	) name3884 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w2320_,
		_w2473_,
		_w5234_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3885 (
		_w2474_,
		_w4975_,
		_w4976_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h1)
	) name3886 (
		_w2477_,
		_w5235_,
		_w5236_
	);
	LUT3 #(
		.INIT('ha8)
	) name3887 (
		_w1679_,
		_w5233_,
		_w5236_,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name3888 (
		_w2283_,
		_w5235_,
		_w5238_
	);
	LUT4 #(
		.INIT('hc055)
	) name3889 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2473_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name3890 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w2288_,
		_w5240_
	);
	LUT3 #(
		.INIT('h0d)
	) name3891 (
		_w2246_,
		_w5239_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h4)
	) name3892 (
		_w5238_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('hb)
	) name3893 (
		_w5237_,
		_w5242_,
		_w5243_
	);
	LUT3 #(
		.INIT('ha8)
	) name3894 (
		_w2320_,
		_w4970_,
		_w4971_,
		_w5244_
	);
	LUT3 #(
		.INIT('ha8)
	) name3895 (
		_w2322_,
		_w4966_,
		_w4967_,
		_w5245_
	);
	LUT3 #(
		.INIT('ha8)
	) name3896 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5244_,
		_w5245_,
		_w5246_
	);
	LUT3 #(
		.INIT('h02)
	) name3897 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w2473_,
		_w2502_,
		_w5247_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3898 (
		_w2503_,
		_w4975_,
		_w4976_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name3899 (
		_w2506_,
		_w5248_,
		_w5249_
	);
	LUT3 #(
		.INIT('ha8)
	) name3900 (
		_w1679_,
		_w5246_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		_w2283_,
		_w5248_,
		_w5251_
	);
	LUT4 #(
		.INIT('hc055)
	) name3902 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2502_,
		_w5252_
	);
	LUT2 #(
		.INIT('h2)
	) name3903 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w2288_,
		_w5253_
	);
	LUT3 #(
		.INIT('h0d)
	) name3904 (
		_w2246_,
		_w5252_,
		_w5253_,
		_w5254_
	);
	LUT2 #(
		.INIT('h4)
	) name3905 (
		_w5251_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('hb)
	) name3906 (
		_w5250_,
		_w5255_,
		_w5256_
	);
	LUT3 #(
		.INIT('ha8)
	) name3907 (
		_w2320_,
		_w4966_,
		_w4967_,
		_w5257_
	);
	LUT3 #(
		.INIT('ha8)
	) name3908 (
		_w2473_,
		_w4970_,
		_w4971_,
		_w5258_
	);
	LUT3 #(
		.INIT('ha8)
	) name3909 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5257_,
		_w5258_,
		_w5259_
	);
	LUT3 #(
		.INIT('h02)
	) name3910 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w2502_,
		_w2528_,
		_w5260_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3911 (
		_w2529_,
		_w4975_,
		_w4976_,
		_w5260_,
		_w5261_
	);
	LUT2 #(
		.INIT('h1)
	) name3912 (
		_w2532_,
		_w5261_,
		_w5262_
	);
	LUT3 #(
		.INIT('ha8)
	) name3913 (
		_w1679_,
		_w5259_,
		_w5262_,
		_w5263_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		_w2283_,
		_w5261_,
		_w5264_
	);
	LUT4 #(
		.INIT('hc055)
	) name3915 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2528_,
		_w5265_
	);
	LUT2 #(
		.INIT('h2)
	) name3916 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w2288_,
		_w5266_
	);
	LUT3 #(
		.INIT('h0d)
	) name3917 (
		_w2246_,
		_w5265_,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name3918 (
		_w5264_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('hb)
	) name3919 (
		_w5263_,
		_w5268_,
		_w5269_
	);
	LUT3 #(
		.INIT('ha8)
	) name3920 (
		_w2473_,
		_w4966_,
		_w4967_,
		_w5270_
	);
	LUT3 #(
		.INIT('ha8)
	) name3921 (
		_w2502_,
		_w4970_,
		_w4971_,
		_w5271_
	);
	LUT3 #(
		.INIT('ha8)
	) name3922 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5270_,
		_w5271_,
		_w5272_
	);
	LUT3 #(
		.INIT('h02)
	) name3923 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w2528_,
		_w2554_,
		_w5273_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3924 (
		_w2555_,
		_w4975_,
		_w4976_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name3925 (
		_w2558_,
		_w5274_,
		_w5275_
	);
	LUT3 #(
		.INIT('ha8)
	) name3926 (
		_w1679_,
		_w5272_,
		_w5275_,
		_w5276_
	);
	LUT2 #(
		.INIT('h2)
	) name3927 (
		_w2283_,
		_w5274_,
		_w5277_
	);
	LUT4 #(
		.INIT('hc055)
	) name3928 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2554_,
		_w5278_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w2288_,
		_w5279_
	);
	LUT3 #(
		.INIT('h0d)
	) name3930 (
		_w2246_,
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h4)
	) name3931 (
		_w5277_,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('hb)
	) name3932 (
		_w5276_,
		_w5281_,
		_w5282_
	);
	LUT3 #(
		.INIT('ha8)
	) name3933 (
		_w2502_,
		_w4966_,
		_w4967_,
		_w5283_
	);
	LUT3 #(
		.INIT('ha8)
	) name3934 (
		_w2528_,
		_w4970_,
		_w4971_,
		_w5284_
	);
	LUT3 #(
		.INIT('ha8)
	) name3935 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5283_,
		_w5284_,
		_w5285_
	);
	LUT3 #(
		.INIT('h02)
	) name3936 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w2554_,
		_w2580_,
		_w5286_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3937 (
		_w2581_,
		_w4975_,
		_w4976_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name3938 (
		_w2584_,
		_w5287_,
		_w5288_
	);
	LUT3 #(
		.INIT('ha8)
	) name3939 (
		_w1679_,
		_w5285_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h2)
	) name3940 (
		_w2283_,
		_w5287_,
		_w5290_
	);
	LUT4 #(
		.INIT('hc055)
	) name3941 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2580_,
		_w5291_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w2288_,
		_w5292_
	);
	LUT3 #(
		.INIT('h0d)
	) name3943 (
		_w2246_,
		_w5291_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h4)
	) name3944 (
		_w5290_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('hb)
	) name3945 (
		_w5289_,
		_w5294_,
		_w5295_
	);
	LUT3 #(
		.INIT('ha8)
	) name3946 (
		_w2528_,
		_w4966_,
		_w4967_,
		_w5296_
	);
	LUT3 #(
		.INIT('ha8)
	) name3947 (
		_w2554_,
		_w4970_,
		_w4971_,
		_w5297_
	);
	LUT3 #(
		.INIT('ha8)
	) name3948 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5298_
	);
	LUT3 #(
		.INIT('h02)
	) name3949 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w2580_,
		_w2606_,
		_w5299_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3950 (
		_w2607_,
		_w4975_,
		_w4976_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w2610_,
		_w5300_,
		_w5301_
	);
	LUT3 #(
		.INIT('ha8)
	) name3952 (
		_w1679_,
		_w5298_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h2)
	) name3953 (
		_w2283_,
		_w5300_,
		_w5303_
	);
	LUT4 #(
		.INIT('hc055)
	) name3954 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2606_,
		_w5304_
	);
	LUT2 #(
		.INIT('h2)
	) name3955 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w2288_,
		_w5305_
	);
	LUT3 #(
		.INIT('h0d)
	) name3956 (
		_w2246_,
		_w5304_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w5303_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('hb)
	) name3958 (
		_w5302_,
		_w5307_,
		_w5308_
	);
	LUT3 #(
		.INIT('ha8)
	) name3959 (
		_w2554_,
		_w4966_,
		_w4967_,
		_w5309_
	);
	LUT3 #(
		.INIT('ha8)
	) name3960 (
		_w2580_,
		_w4970_,
		_w4971_,
		_w5310_
	);
	LUT3 #(
		.INIT('ha8)
	) name3961 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5309_,
		_w5310_,
		_w5311_
	);
	LUT3 #(
		.INIT('h02)
	) name3962 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w2349_,
		_w2606_,
		_w5312_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3963 (
		_w2632_,
		_w4975_,
		_w4976_,
		_w5312_,
		_w5313_
	);
	LUT2 #(
		.INIT('h1)
	) name3964 (
		_w2635_,
		_w5313_,
		_w5314_
	);
	LUT3 #(
		.INIT('ha8)
	) name3965 (
		_w1679_,
		_w5311_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h2)
	) name3966 (
		_w2283_,
		_w5313_,
		_w5316_
	);
	LUT4 #(
		.INIT('hc055)
	) name3967 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2349_,
		_w5317_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w2288_,
		_w5318_
	);
	LUT3 #(
		.INIT('h0d)
	) name3969 (
		_w2246_,
		_w5317_,
		_w5318_,
		_w5319_
	);
	LUT2 #(
		.INIT('h4)
	) name3970 (
		_w5316_,
		_w5319_,
		_w5320_
	);
	LUT2 #(
		.INIT('hb)
	) name3971 (
		_w5315_,
		_w5320_,
		_w5321_
	);
	LUT3 #(
		.INIT('ha8)
	) name3972 (
		_w2580_,
		_w4966_,
		_w4967_,
		_w5322_
	);
	LUT3 #(
		.INIT('ha8)
	) name3973 (
		_w2606_,
		_w4970_,
		_w4971_,
		_w5323_
	);
	LUT3 #(
		.INIT('ha8)
	) name3974 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5322_,
		_w5323_,
		_w5324_
	);
	LUT3 #(
		.INIT('h02)
	) name3975 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w2250_,
		_w2349_,
		_w5325_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3976 (
		_w2350_,
		_w4975_,
		_w4976_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		_w2659_,
		_w5326_,
		_w5327_
	);
	LUT3 #(
		.INIT('ha8)
	) name3978 (
		_w1679_,
		_w5324_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h2)
	) name3979 (
		_w2283_,
		_w5326_,
		_w5329_
	);
	LUT4 #(
		.INIT('hc055)
	) name3980 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2250_,
		_w5330_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w2288_,
		_w5331_
	);
	LUT3 #(
		.INIT('h0d)
	) name3982 (
		_w2246_,
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h4)
	) name3983 (
		_w5329_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('hb)
	) name3984 (
		_w5328_,
		_w5333_,
		_w5334_
	);
	LUT3 #(
		.INIT('ha8)
	) name3985 (
		_w2606_,
		_w4966_,
		_w4967_,
		_w5335_
	);
	LUT3 #(
		.INIT('ha8)
	) name3986 (
		_w2349_,
		_w4970_,
		_w4971_,
		_w5336_
	);
	LUT3 #(
		.INIT('ha8)
	) name3987 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5335_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('h02)
	) name3988 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w2250_,
		_w2264_,
		_w5338_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3989 (
		_w2279_,
		_w4975_,
		_w4976_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w2683_,
		_w5339_,
		_w5340_
	);
	LUT3 #(
		.INIT('ha8)
	) name3991 (
		_w1679_,
		_w5337_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		_w2283_,
		_w5339_,
		_w5342_
	);
	LUT4 #(
		.INIT('hc055)
	) name3993 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1508_,
		_w1513_,
		_w2264_,
		_w5343_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w2288_,
		_w5344_
	);
	LUT3 #(
		.INIT('h0d)
	) name3995 (
		_w2246_,
		_w5343_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name3996 (
		_w5342_,
		_w5345_,
		_w5346_
	);
	LUT2 #(
		.INIT('hb)
	) name3997 (
		_w5341_,
		_w5346_,
		_w5347_
	);
	LUT3 #(
		.INIT('h80)
	) name3998 (
		_w2890_,
		_w4065_,
		_w4075_,
		_w5348_
	);
	LUT4 #(
		.INIT('h2000)
	) name3999 (
		_w2890_,
		_w2900_,
		_w4065_,
		_w4075_,
		_w5349_
	);
	LUT4 #(
		.INIT('h0800)
	) name4000 (
		_w2879_,
		_w2874_,
		_w2901_,
		_w5349_,
		_w5350_
	);
	LUT4 #(
		.INIT('h870f)
	) name4001 (
		_w2879_,
		_w2874_,
		_w2901_,
		_w5349_,
		_w5351_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w2755_,
		_w5351_,
		_w5352_
	);
	LUT4 #(
		.INIT('hf700)
	) name4003 (
		_w2749_,
		_w2754_,
		_w2936_,
		_w2944_,
		_w5353_
	);
	LUT3 #(
		.INIT('h6c)
	) name4004 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2715_,
		_w5354_
	);
	LUT4 #(
		.INIT('h28a0)
	) name4005 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2715_,
		_w5355_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w4053_,
		_w5355_,
		_w5356_
	);
	LUT4 #(
		.INIT('hb000)
	) name4007 (
		_w2935_,
		_w2941_,
		_w5353_,
		_w5356_,
		_w5357_
	);
	LUT3 #(
		.INIT('h6c)
	) name4008 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2718_,
		_w5358_
	);
	LUT3 #(
		.INIT('h80)
	) name4009 (
		_w2955_,
		_w4055_,
		_w5358_,
		_w5359_
	);
	LUT3 #(
		.INIT('h6a)
	) name4010 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2706_,
		_w2893_,
		_w5360_
	);
	LUT3 #(
		.INIT('h80)
	) name4011 (
		_w2965_,
		_w4773_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h1555)
	) name4012 (
		_w2963_,
		_w5357_,
		_w5359_,
		_w5361_,
		_w5362_
	);
	LUT4 #(
		.INIT('h2000)
	) name4013 (
		_w2965_,
		_w4051_,
		_w4054_,
		_w4057_,
		_w5363_
	);
	LUT4 #(
		.INIT('h002a)
	) name4014 (
		_w2755_,
		_w2963_,
		_w5363_,
		_w5362_,
		_w5364_
	);
	LUT4 #(
		.INIT('h4447)
	) name4015 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2173_,
		_w5352_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('h2a80)
	) name4016 (
		_w2181_,
		_w3025_,
		_w3028_,
		_w3032_,
		_w5366_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2098_,
		_w5367_
	);
	LUT3 #(
		.INIT('h0e)
	) name4018 (
		_w2071_,
		_w2087_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w3032_,
		_w5368_,
		_w5369_
	);
	LUT4 #(
		.INIT('he400)
	) name4020 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2963_,
		_w5370_
	);
	LUT4 #(
		.INIT('h001f)
	) name4021 (
		_w2108_,
		_w2115_,
		_w2116_,
		_w2125_,
		_w5371_
	);
	LUT4 #(
		.INIT('h0400)
	) name4022 (
		_w2136_,
		_w2176_,
		_w5370_,
		_w5371_,
		_w5372_
	);
	LUT3 #(
		.INIT('hb0)
	) name4023 (
		_w2073_,
		_w2086_,
		_w2901_,
		_w5373_
	);
	LUT2 #(
		.INIT('h4)
	) name4024 (
		_w2117_,
		_w2963_,
		_w5374_
	);
	LUT4 #(
		.INIT('h0031)
	) name4025 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w5373_,
		_w5372_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h10)
	) name4026 (
		_w5366_,
		_w5369_,
		_w5375_,
		_w5376_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4027 (
		_w1945_,
		_w2171_,
		_w5365_,
		_w5376_,
		_w5377_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4028 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w3054_,
		_w3056_,
		_w5378_
	);
	LUT2 #(
		.INIT('hb)
	) name4029 (
		_w5377_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h8)
	) name4030 (
		_w2902_,
		_w2908_,
		_w5380_
	);
	LUT4 #(
		.INIT('h8000)
	) name4031 (
		_w4068_,
		_w4074_,
		_w5348_,
		_w5380_,
		_w5381_
	);
	LUT3 #(
		.INIT('h8c)
	) name4032 (
		_w2905_,
		_w2909_,
		_w5381_,
		_w5382_
	);
	LUT3 #(
		.INIT('h04)
	) name4033 (
		_w2905_,
		_w2908_,
		_w2909_,
		_w5383_
	);
	LUT3 #(
		.INIT('h15)
	) name4034 (
		_w2755_,
		_w5350_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('h4800)
	) name4035 (
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2961_,
		_w2962_,
		_w2972_,
		_w5385_
	);
	LUT4 #(
		.INIT('h8000)
	) name4036 (
		_w5357_,
		_w5359_,
		_w5361_,
		_w5385_,
		_w5386_
	);
	LUT3 #(
		.INIT('h28)
	) name4037 (
		_w2755_,
		_w2970_,
		_w5386_,
		_w5387_
	);
	LUT4 #(
		.INIT('h5510)
	) name4038 (
		_w2173_,
		_w5382_,
		_w5384_,
		_w5387_,
		_w5388_
	);
	LUT3 #(
		.INIT('h02)
	) name4039 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w2103_,
		_w2172_,
		_w5389_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w2116_,
		_w2970_,
		_w5390_
	);
	LUT3 #(
		.INIT('h08)
	) name4041 (
		_w2060_,
		_w2044_,
		_w5390_,
		_w5391_
	);
	LUT4 #(
		.INIT('h0010)
	) name4042 (
		_w2127_,
		_w4784_,
		_w4785_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h4)
	) name4043 (
		_w2117_,
		_w2970_,
		_w5393_
	);
	LUT4 #(
		.INIT('he000)
	) name4044 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3039_,
		_w5394_
	);
	LUT4 #(
		.INIT('h00f4)
	) name4045 (
		_w2073_,
		_w2086_,
		_w2909_,
		_w5394_,
		_w5395_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4046 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		_w5392_,
		_w5393_,
		_w5395_,
		_w5396_
	);
	LUT4 #(
		.INIT('hd700)
	) name4047 (
		_w2181_,
		_w3037_,
		_w3039_,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('h5700)
	) name4048 (
		_w2171_,
		_w5388_,
		_w5389_,
		_w5397_,
		_w5398_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4049 (
		\P3_InstAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w3054_,
		_w3056_,
		_w5399_
	);
	LUT3 #(
		.INIT('h2f)
	) name4050 (
		_w1945_,
		_w5398_,
		_w5399_,
		_w5400_
	);
	LUT3 #(
		.INIT('h08)
	) name4051 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5401_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		_w4798_,
		_w4796_,
		_w5402_
	);
	LUT3 #(
		.INIT('h08)
	) name4053 (
		_w4223_,
		_w4229_,
		_w4807_,
		_w5403_
	);
	LUT4 #(
		.INIT('h4554)
	) name4054 (
		_w1661_,
		_w4214_,
		_w4324_,
		_w4826_,
		_w5404_
	);
	LUT4 #(
		.INIT('h5700)
	) name4055 (
		_w4214_,
		_w5402_,
		_w5403_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4056 (
		_w1659_,
		_w4400_,
		_w4832_,
		_w4836_,
		_w5406_
	);
	LUT4 #(
		.INIT('h01aa)
	) name4057 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w1592_,
		_w1595_,
		_w4406_,
		_w5407_
	);
	LUT4 #(
		.INIT('hc800)
	) name4058 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w5407_,
		_w5408_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4059 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		_w1658_,
		_w4844_,
		_w5408_,
		_w5409_
	);
	LUT3 #(
		.INIT('hb0)
	) name4060 (
		_w1571_,
		_w1583_,
		_w4324_,
		_w5410_
	);
	LUT2 #(
		.INIT('h4)
	) name4061 (
		_w1617_,
		_w4798_,
		_w5411_
	);
	LUT4 #(
		.INIT('h0100)
	) name4062 (
		_w5406_,
		_w5410_,
		_w5411_,
		_w5409_,
		_w5412_
	);
	LUT4 #(
		.INIT('h5700)
	) name4063 (
		_w1559_,
		_w5401_,
		_w5405_,
		_w5412_,
		_w5413_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4064 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5414_
	);
	LUT3 #(
		.INIT('h2f)
	) name4065 (
		_w1678_,
		_w5413_,
		_w5414_,
		_w5415_
	);
	LUT3 #(
		.INIT('h08)
	) name4066 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5416_
	);
	LUT4 #(
		.INIT('h1405)
	) name4067 (
		_w4214_,
		_w4340_,
		_w4342_,
		_w4855_,
		_w5417_
	);
	LUT4 #(
		.INIT('h4555)
	) name4068 (
		_w4249_,
		_w4807_,
		_w4810_,
		_w4858_,
		_w5418_
	);
	LUT4 #(
		.INIT('h1115)
	) name4069 (
		_w1661_,
		_w4214_,
		_w4897_,
		_w5418_,
		_w5419_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4070 (
		_w1559_,
		_w5416_,
		_w5417_,
		_w5419_,
		_w5420_
	);
	LUT3 #(
		.INIT('h28)
	) name4071 (
		_w1659_,
		_w4865_,
		_w4872_,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w1656_,
		_w5422_
	);
	LUT3 #(
		.INIT('hc4)
	) name4073 (
		_w1617_,
		_w4249_,
		_w5422_,
		_w5423_
	);
	LUT4 #(
		.INIT('h0800)
	) name4074 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1596_,
		_w4410_,
		_w5424_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w5424_,
		_w5425_
	);
	LUT4 #(
		.INIT('hc800)
	) name4076 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w4865_,
		_w5426_
	);
	LUT2 #(
		.INIT('h4)
	) name4077 (
		_w5425_,
		_w5426_,
		_w5427_
	);
	LUT3 #(
		.INIT('hb0)
	) name4078 (
		_w1571_,
		_w1583_,
		_w4342_,
		_w5428_
	);
	LUT3 #(
		.INIT('h13)
	) name4079 (
		_w1605_,
		_w1613_,
		_w1656_,
		_w5429_
	);
	LUT3 #(
		.INIT('h2a)
	) name4080 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w4844_,
		_w5429_,
		_w5430_
	);
	LUT4 #(
		.INIT('h0001)
	) name4081 (
		_w5428_,
		_w5423_,
		_w5430_,
		_w5427_,
		_w5431_
	);
	LUT2 #(
		.INIT('h4)
	) name4082 (
		_w5421_,
		_w5431_,
		_w5432_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4083 (
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5433_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4084 (
		_w1678_,
		_w5420_,
		_w5432_,
		_w5433_,
		_w5434_
	);
	LUT3 #(
		.INIT('h08)
	) name4085 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5435_
	);
	LUT3 #(
		.INIT('h82)
	) name4086 (
		_w4214_,
		_w4267_,
		_w4270_,
		_w5436_
	);
	LUT4 #(
		.INIT('h4554)
	) name4087 (
		_w1661_,
		_w4214_,
		_w4359_,
		_w4361_,
		_w5437_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4088 (
		_w1559_,
		_w5435_,
		_w5436_,
		_w5437_,
		_w5438_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		_w1640_,
		_w4428_,
		_w5439_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		_w1555_,
		_w4423_,
		_w5440_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4091 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1605_,
		_w5441_
	);
	LUT3 #(
		.INIT('h54)
	) name4092 (
		_w1602_,
		_w1625_,
		_w5441_,
		_w5442_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4093 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		_w4844_,
		_w5440_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		_w1617_,
		_w4270_,
		_w5444_
	);
	LUT3 #(
		.INIT('hb0)
	) name4095 (
		_w1571_,
		_w1583_,
		_w4361_,
		_w5445_
	);
	LUT4 #(
		.INIT('h0001)
	) name4096 (
		_w5444_,
		_w5443_,
		_w5445_,
		_w5439_,
		_w5446_
	);
	LUT4 #(
		.INIT('hd700)
	) name4097 (
		_w1659_,
		_w4422_,
		_w4428_,
		_w5446_,
		_w5447_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4098 (
		\P2_InstAddrPointer_reg[25]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5448_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4099 (
		_w1678_,
		_w5438_,
		_w5447_,
		_w5448_,
		_w5449_
	);
	LUT3 #(
		.INIT('h08)
	) name4100 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1842_,
		_w1915_,
		_w5450_
	);
	LUT3 #(
		.INIT('h01)
	) name4101 (
		_w3243_,
		_w3246_,
		_w3254_,
		_w5451_
	);
	LUT4 #(
		.INIT('h0001)
	) name4102 (
		_w3243_,
		_w3245_,
		_w3246_,
		_w3254_,
		_w5452_
	);
	LUT4 #(
		.INIT('h4000)
	) name4103 (
		_w3090_,
		_w3214_,
		_w3223_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h2)
	) name4104 (
		_w3244_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h4000)
	) name4105 (
		_w3090_,
		_w3214_,
		_w3223_,
		_w4726_,
		_w5455_
	);
	LUT3 #(
		.INIT('h15)
	) name4106 (
		_w3101_,
		_w3247_,
		_w5455_,
		_w5456_
	);
	LUT4 #(
		.INIT('h1333)
	) name4107 (
		_w3296_,
		_w3305_,
		_w3991_,
		_w3995_,
		_w5457_
	);
	LUT4 #(
		.INIT('h8000)
	) name4108 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w3296_,
		_w3991_,
		_w3995_,
		_w5458_
	);
	LUT4 #(
		.INIT('h1115)
	) name4109 (
		_w1916_,
		_w3101_,
		_w5457_,
		_w5458_,
		_w5459_
	);
	LUT4 #(
		.INIT('h1055)
	) name4110 (
		_w5450_,
		_w5454_,
		_w5456_,
		_w5459_,
		_w5460_
	);
	LUT4 #(
		.INIT('h2888)
	) name4111 (
		_w1924_,
		_w3373_,
		_w3364_,
		_w3372_,
		_w5461_
	);
	LUT4 #(
		.INIT('h9030)
	) name4112 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1920_,
		_w3072_,
		_w5462_
	);
	LUT2 #(
		.INIT('h2)
	) name4113 (
		_w4739_,
		_w5462_,
		_w5463_
	);
	LUT3 #(
		.INIT('ha2)
	) name4114 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w4037_,
		_w5463_,
		_w5464_
	);
	LUT3 #(
		.INIT('h54)
	) name4115 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1842_,
		_w1845_,
		_w5465_
	);
	LUT3 #(
		.INIT('h04)
	) name4116 (
		_w1833_,
		_w3373_,
		_w5465_,
		_w5466_
	);
	LUT3 #(
		.INIT('h80)
	) name4117 (
		_w1805_,
		_w1806_,
		_w3305_,
		_w5467_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name4118 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		_w1861_,
		_w3072_,
		_w5468_
	);
	LUT4 #(
		.INIT('h010f)
	) name4119 (
		_w1855_,
		_w1860_,
		_w5467_,
		_w5468_,
		_w5469_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4120 (
		_w1816_,
		_w1831_,
		_w3244_,
		_w5469_,
		_w5470_
	);
	LUT3 #(
		.INIT('h10)
	) name4121 (
		_w5464_,
		_w5466_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h4)
	) name4122 (
		_w5461_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4123 (
		_w1810_,
		_w1933_,
		_w5460_,
		_w5472_,
		_w5473_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4124 (
		\P1_InstAddrPointer_reg[18]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w3406_,
		_w3408_,
		_w5474_
	);
	LUT2 #(
		.INIT('hb)
	) name4125 (
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT4 #(
		.INIT('hc444)
	) name4126 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5476_
	);
	LUT4 #(
		.INIT('h0888)
	) name4127 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[26]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5477_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		_w5476_,
		_w5477_,
		_w5478_
	);
	LUT3 #(
		.INIT('ha8)
	) name4129 (
		_w2250_,
		_w5476_,
		_w5477_,
		_w5479_
	);
	LUT4 #(
		.INIT('hc444)
	) name4130 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[18]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5480_
	);
	LUT4 #(
		.INIT('h0888)
	) name4131 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[18]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w5480_,
		_w5481_,
		_w5482_
	);
	LUT3 #(
		.INIT('ha8)
	) name4133 (
		_w2264_,
		_w5480_,
		_w5481_,
		_w5483_
	);
	LUT3 #(
		.INIT('ha8)
	) name4134 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5479_,
		_w5483_,
		_w5484_
	);
	LUT4 #(
		.INIT('hc444)
	) name4135 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5485_
	);
	LUT4 #(
		.INIT('h0888)
	) name4136 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[2]/NET0131 ,
		_w2255_,
		_w2260_,
		_w5486_
	);
	LUT2 #(
		.INIT('h1)
	) name4137 (
		_w5485_,
		_w5486_,
		_w5487_
	);
	LUT3 #(
		.INIT('h02)
	) name4138 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w2271_,
		_w2272_,
		_w5488_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4139 (
		_w2273_,
		_w5485_,
		_w5486_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		_w2280_,
		_w5489_,
		_w5490_
	);
	LUT3 #(
		.INIT('ha8)
	) name4141 (
		_w1679_,
		_w5484_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h2)
	) name4142 (
		_w2283_,
		_w5489_,
		_w5492_
	);
	LUT4 #(
		.INIT('hc055)
	) name4143 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2272_,
		_w5493_
	);
	LUT2 #(
		.INIT('h2)
	) name4144 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		_w2288_,
		_w5494_
	);
	LUT3 #(
		.INIT('h0d)
	) name4145 (
		_w2246_,
		_w5493_,
		_w5494_,
		_w5495_
	);
	LUT2 #(
		.INIT('h4)
	) name4146 (
		_w5492_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('hb)
	) name4147 (
		_w5491_,
		_w5496_,
		_w5497_
	);
	LUT3 #(
		.INIT('ha8)
	) name4148 (
		_w2315_,
		_w5476_,
		_w5477_,
		_w5498_
	);
	LUT3 #(
		.INIT('ha8)
	) name4149 (
		_w2317_,
		_w5480_,
		_w5481_,
		_w5499_
	);
	LUT3 #(
		.INIT('ha8)
	) name4150 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5498_,
		_w5499_,
		_w5500_
	);
	LUT3 #(
		.INIT('h02)
	) name4151 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w2320_,
		_w2322_,
		_w5501_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4152 (
		_w2323_,
		_w5485_,
		_w5486_,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		_w2327_,
		_w5502_,
		_w5503_
	);
	LUT3 #(
		.INIT('ha8)
	) name4154 (
		_w1679_,
		_w5500_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h2)
	) name4155 (
		_w2283_,
		_w5502_,
		_w5505_
	);
	LUT4 #(
		.INIT('hc055)
	) name4156 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2320_,
		_w5506_
	);
	LUT2 #(
		.INIT('h2)
	) name4157 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		_w2288_,
		_w5507_
	);
	LUT3 #(
		.INIT('h0d)
	) name4158 (
		_w2246_,
		_w5506_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h4)
	) name4159 (
		_w5505_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('hb)
	) name4160 (
		_w5504_,
		_w5509_,
		_w5510_
	);
	LUT3 #(
		.INIT('ha8)
	) name4161 (
		_w2250_,
		_w5480_,
		_w5481_,
		_w5511_
	);
	LUT3 #(
		.INIT('ha8)
	) name4162 (
		_w2349_,
		_w5476_,
		_w5477_,
		_w5512_
	);
	LUT3 #(
		.INIT('ha8)
	) name4163 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5511_,
		_w5512_,
		_w5513_
	);
	LUT3 #(
		.INIT('h02)
	) name4164 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w2271_,
		_w2264_,
		_w5514_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4165 (
		_w2346_,
		_w5485_,
		_w5486_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		_w2351_,
		_w5515_,
		_w5516_
	);
	LUT3 #(
		.INIT('ha8)
	) name4167 (
		_w1679_,
		_w5513_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h2)
	) name4168 (
		_w2283_,
		_w5515_,
		_w5518_
	);
	LUT4 #(
		.INIT('hc055)
	) name4169 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2271_,
		_w5519_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		_w2288_,
		_w5520_
	);
	LUT3 #(
		.INIT('h0d)
	) name4171 (
		_w2246_,
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h4)
	) name4172 (
		_w5518_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('hb)
	) name4173 (
		_w5517_,
		_w5522_,
		_w5523_
	);
	LUT3 #(
		.INIT('ha8)
	) name4174 (
		_w2264_,
		_w5476_,
		_w5477_,
		_w5524_
	);
	LUT3 #(
		.INIT('ha8)
	) name4175 (
		_w2271_,
		_w5480_,
		_w5481_,
		_w5525_
	);
	LUT3 #(
		.INIT('ha8)
	) name4176 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5524_,
		_w5525_,
		_w5526_
	);
	LUT3 #(
		.INIT('h02)
	) name4177 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w2272_,
		_w2376_,
		_w5527_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4178 (
		_w2377_,
		_w5485_,
		_w5486_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name4179 (
		_w2380_,
		_w5528_,
		_w5529_
	);
	LUT3 #(
		.INIT('ha8)
	) name4180 (
		_w1679_,
		_w5526_,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h2)
	) name4181 (
		_w2283_,
		_w5528_,
		_w5531_
	);
	LUT4 #(
		.INIT('hc055)
	) name4182 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2376_,
		_w5532_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		_w2288_,
		_w5533_
	);
	LUT3 #(
		.INIT('h0d)
	) name4184 (
		_w2246_,
		_w5532_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h4)
	) name4185 (
		_w5531_,
		_w5534_,
		_w5535_
	);
	LUT2 #(
		.INIT('hb)
	) name4186 (
		_w5530_,
		_w5535_,
		_w5536_
	);
	LUT3 #(
		.INIT('ha8)
	) name4187 (
		_w2271_,
		_w5476_,
		_w5477_,
		_w5537_
	);
	LUT3 #(
		.INIT('ha8)
	) name4188 (
		_w2272_,
		_w5480_,
		_w5481_,
		_w5538_
	);
	LUT3 #(
		.INIT('ha8)
	) name4189 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5537_,
		_w5538_,
		_w5539_
	);
	LUT3 #(
		.INIT('h02)
	) name4190 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w2315_,
		_w2376_,
		_w5540_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4191 (
		_w2402_,
		_w5485_,
		_w5486_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name4192 (
		_w2405_,
		_w5541_,
		_w5542_
	);
	LUT3 #(
		.INIT('ha8)
	) name4193 (
		_w1679_,
		_w5539_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		_w2283_,
		_w5541_,
		_w5544_
	);
	LUT4 #(
		.INIT('hc055)
	) name4195 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2315_,
		_w5545_
	);
	LUT2 #(
		.INIT('h2)
	) name4196 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w2288_,
		_w5546_
	);
	LUT3 #(
		.INIT('h0d)
	) name4197 (
		_w2246_,
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		_w5544_,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('hb)
	) name4199 (
		_w5543_,
		_w5548_,
		_w5549_
	);
	LUT3 #(
		.INIT('ha8)
	) name4200 (
		_w2272_,
		_w5476_,
		_w5477_,
		_w5550_
	);
	LUT3 #(
		.INIT('ha8)
	) name4201 (
		_w2376_,
		_w5480_,
		_w5481_,
		_w5551_
	);
	LUT3 #(
		.INIT('ha8)
	) name4202 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5550_,
		_w5551_,
		_w5552_
	);
	LUT3 #(
		.INIT('h02)
	) name4203 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w2315_,
		_w2317_,
		_w5553_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4204 (
		_w2326_,
		_w5485_,
		_w5486_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w2429_,
		_w5554_,
		_w5555_
	);
	LUT3 #(
		.INIT('ha8)
	) name4206 (
		_w1679_,
		_w5552_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		_w2283_,
		_w5554_,
		_w5557_
	);
	LUT4 #(
		.INIT('hc055)
	) name4208 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2317_,
		_w5558_
	);
	LUT2 #(
		.INIT('h2)
	) name4209 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		_w2288_,
		_w5559_
	);
	LUT3 #(
		.INIT('h0d)
	) name4210 (
		_w2246_,
		_w5558_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h4)
	) name4211 (
		_w5557_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('hb)
	) name4212 (
		_w5556_,
		_w5561_,
		_w5562_
	);
	LUT3 #(
		.INIT('ha8)
	) name4213 (
		_w2376_,
		_w5476_,
		_w5477_,
		_w5563_
	);
	LUT3 #(
		.INIT('ha8)
	) name4214 (
		_w2315_,
		_w5480_,
		_w5481_,
		_w5564_
	);
	LUT3 #(
		.INIT('ha8)
	) name4215 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5563_,
		_w5564_,
		_w5565_
	);
	LUT3 #(
		.INIT('h02)
	) name4216 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w2322_,
		_w2317_,
		_w5566_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4217 (
		_w2451_,
		_w5485_,
		_w5486_,
		_w5566_,
		_w5567_
	);
	LUT2 #(
		.INIT('h1)
	) name4218 (
		_w2454_,
		_w5567_,
		_w5568_
	);
	LUT3 #(
		.INIT('ha8)
	) name4219 (
		_w1679_,
		_w5565_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('h2)
	) name4220 (
		_w2283_,
		_w5567_,
		_w5570_
	);
	LUT4 #(
		.INIT('hc055)
	) name4221 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2322_,
		_w5571_
	);
	LUT2 #(
		.INIT('h2)
	) name4222 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w2288_,
		_w5572_
	);
	LUT3 #(
		.INIT('h0d)
	) name4223 (
		_w2246_,
		_w5571_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h4)
	) name4224 (
		_w5570_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('hb)
	) name4225 (
		_w5569_,
		_w5574_,
		_w5575_
	);
	LUT3 #(
		.INIT('ha8)
	) name4226 (
		_w2317_,
		_w5476_,
		_w5477_,
		_w5576_
	);
	LUT3 #(
		.INIT('ha8)
	) name4227 (
		_w2322_,
		_w5480_,
		_w5481_,
		_w5577_
	);
	LUT3 #(
		.INIT('ha8)
	) name4228 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5576_,
		_w5577_,
		_w5578_
	);
	LUT3 #(
		.INIT('h02)
	) name4229 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w2320_,
		_w2473_,
		_w5579_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4230 (
		_w2474_,
		_w5485_,
		_w5486_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w2477_,
		_w5580_,
		_w5581_
	);
	LUT3 #(
		.INIT('ha8)
	) name4232 (
		_w1679_,
		_w5578_,
		_w5581_,
		_w5582_
	);
	LUT2 #(
		.INIT('h2)
	) name4233 (
		_w2283_,
		_w5580_,
		_w5583_
	);
	LUT4 #(
		.INIT('hc055)
	) name4234 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2473_,
		_w5584_
	);
	LUT2 #(
		.INIT('h2)
	) name4235 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w2288_,
		_w5585_
	);
	LUT3 #(
		.INIT('h0d)
	) name4236 (
		_w2246_,
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h4)
	) name4237 (
		_w5583_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('hb)
	) name4238 (
		_w5582_,
		_w5587_,
		_w5588_
	);
	LUT3 #(
		.INIT('ha8)
	) name4239 (
		_w2320_,
		_w5480_,
		_w5481_,
		_w5589_
	);
	LUT3 #(
		.INIT('ha8)
	) name4240 (
		_w2322_,
		_w5476_,
		_w5477_,
		_w5590_
	);
	LUT3 #(
		.INIT('ha8)
	) name4241 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5589_,
		_w5590_,
		_w5591_
	);
	LUT3 #(
		.INIT('h02)
	) name4242 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w2473_,
		_w2502_,
		_w5592_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4243 (
		_w2503_,
		_w5485_,
		_w5486_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h1)
	) name4244 (
		_w2506_,
		_w5593_,
		_w5594_
	);
	LUT3 #(
		.INIT('ha8)
	) name4245 (
		_w1679_,
		_w5591_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name4246 (
		_w2283_,
		_w5593_,
		_w5596_
	);
	LUT4 #(
		.INIT('hc055)
	) name4247 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2502_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name4248 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w2288_,
		_w5598_
	);
	LUT3 #(
		.INIT('h0d)
	) name4249 (
		_w2246_,
		_w5597_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h4)
	) name4250 (
		_w5596_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('hb)
	) name4251 (
		_w5595_,
		_w5600_,
		_w5601_
	);
	LUT3 #(
		.INIT('ha8)
	) name4252 (
		_w2320_,
		_w5476_,
		_w5477_,
		_w5602_
	);
	LUT3 #(
		.INIT('ha8)
	) name4253 (
		_w2473_,
		_w5480_,
		_w5481_,
		_w5603_
	);
	LUT3 #(
		.INIT('ha8)
	) name4254 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5602_,
		_w5603_,
		_w5604_
	);
	LUT3 #(
		.INIT('h02)
	) name4255 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w2502_,
		_w2528_,
		_w5605_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4256 (
		_w2529_,
		_w5485_,
		_w5486_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name4257 (
		_w2532_,
		_w5606_,
		_w5607_
	);
	LUT3 #(
		.INIT('ha8)
	) name4258 (
		_w1679_,
		_w5604_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h2)
	) name4259 (
		_w2283_,
		_w5606_,
		_w5609_
	);
	LUT4 #(
		.INIT('hc055)
	) name4260 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2528_,
		_w5610_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w2288_,
		_w5611_
	);
	LUT3 #(
		.INIT('h0d)
	) name4262 (
		_w2246_,
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT2 #(
		.INIT('h4)
	) name4263 (
		_w5609_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('hb)
	) name4264 (
		_w5608_,
		_w5613_,
		_w5614_
	);
	LUT3 #(
		.INIT('ha8)
	) name4265 (
		_w2473_,
		_w5476_,
		_w5477_,
		_w5615_
	);
	LUT3 #(
		.INIT('ha8)
	) name4266 (
		_w2502_,
		_w5480_,
		_w5481_,
		_w5616_
	);
	LUT3 #(
		.INIT('ha8)
	) name4267 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5615_,
		_w5616_,
		_w5617_
	);
	LUT3 #(
		.INIT('h02)
	) name4268 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w2528_,
		_w2554_,
		_w5618_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4269 (
		_w2555_,
		_w5485_,
		_w5486_,
		_w5618_,
		_w5619_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w2558_,
		_w5619_,
		_w5620_
	);
	LUT3 #(
		.INIT('ha8)
	) name4271 (
		_w1679_,
		_w5617_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		_w2283_,
		_w5619_,
		_w5622_
	);
	LUT4 #(
		.INIT('hc055)
	) name4273 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2554_,
		_w5623_
	);
	LUT2 #(
		.INIT('h2)
	) name4274 (
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w2288_,
		_w5624_
	);
	LUT3 #(
		.INIT('h0d)
	) name4275 (
		_w2246_,
		_w5623_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h4)
	) name4276 (
		_w5622_,
		_w5625_,
		_w5626_
	);
	LUT2 #(
		.INIT('hb)
	) name4277 (
		_w5621_,
		_w5626_,
		_w5627_
	);
	LUT3 #(
		.INIT('ha8)
	) name4278 (
		_w2502_,
		_w5476_,
		_w5477_,
		_w5628_
	);
	LUT3 #(
		.INIT('ha8)
	) name4279 (
		_w2528_,
		_w5480_,
		_w5481_,
		_w5629_
	);
	LUT3 #(
		.INIT('ha8)
	) name4280 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5628_,
		_w5629_,
		_w5630_
	);
	LUT3 #(
		.INIT('h02)
	) name4281 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w2554_,
		_w2580_,
		_w5631_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4282 (
		_w2581_,
		_w5485_,
		_w5486_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		_w2584_,
		_w5632_,
		_w5633_
	);
	LUT3 #(
		.INIT('ha8)
	) name4284 (
		_w1679_,
		_w5630_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h2)
	) name4285 (
		_w2283_,
		_w5632_,
		_w5635_
	);
	LUT4 #(
		.INIT('hc055)
	) name4286 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2580_,
		_w5636_
	);
	LUT2 #(
		.INIT('h2)
	) name4287 (
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w2288_,
		_w5637_
	);
	LUT3 #(
		.INIT('h0d)
	) name4288 (
		_w2246_,
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h4)
	) name4289 (
		_w5635_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('hb)
	) name4290 (
		_w5634_,
		_w5639_,
		_w5640_
	);
	LUT3 #(
		.INIT('ha8)
	) name4291 (
		_w2528_,
		_w5476_,
		_w5477_,
		_w5641_
	);
	LUT3 #(
		.INIT('ha8)
	) name4292 (
		_w2554_,
		_w5480_,
		_w5481_,
		_w5642_
	);
	LUT3 #(
		.INIT('ha8)
	) name4293 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5641_,
		_w5642_,
		_w5643_
	);
	LUT3 #(
		.INIT('h02)
	) name4294 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w2580_,
		_w2606_,
		_w5644_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4295 (
		_w2607_,
		_w5485_,
		_w5486_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name4296 (
		_w2610_,
		_w5645_,
		_w5646_
	);
	LUT3 #(
		.INIT('ha8)
	) name4297 (
		_w1679_,
		_w5643_,
		_w5646_,
		_w5647_
	);
	LUT2 #(
		.INIT('h2)
	) name4298 (
		_w2283_,
		_w5645_,
		_w5648_
	);
	LUT4 #(
		.INIT('hc055)
	) name4299 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2606_,
		_w5649_
	);
	LUT2 #(
		.INIT('h2)
	) name4300 (
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w2288_,
		_w5650_
	);
	LUT3 #(
		.INIT('h0d)
	) name4301 (
		_w2246_,
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w5648_,
		_w5651_,
		_w5652_
	);
	LUT2 #(
		.INIT('hb)
	) name4303 (
		_w5647_,
		_w5652_,
		_w5653_
	);
	LUT3 #(
		.INIT('ha8)
	) name4304 (
		_w2554_,
		_w5476_,
		_w5477_,
		_w5654_
	);
	LUT3 #(
		.INIT('ha8)
	) name4305 (
		_w2580_,
		_w5480_,
		_w5481_,
		_w5655_
	);
	LUT3 #(
		.INIT('ha8)
	) name4306 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5654_,
		_w5655_,
		_w5656_
	);
	LUT3 #(
		.INIT('h02)
	) name4307 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w2349_,
		_w2606_,
		_w5657_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4308 (
		_w2632_,
		_w5485_,
		_w5486_,
		_w5657_,
		_w5658_
	);
	LUT2 #(
		.INIT('h1)
	) name4309 (
		_w2635_,
		_w5658_,
		_w5659_
	);
	LUT3 #(
		.INIT('ha8)
	) name4310 (
		_w1679_,
		_w5656_,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h2)
	) name4311 (
		_w2283_,
		_w5658_,
		_w5661_
	);
	LUT4 #(
		.INIT('hc055)
	) name4312 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2349_,
		_w5662_
	);
	LUT2 #(
		.INIT('h2)
	) name4313 (
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w2288_,
		_w5663_
	);
	LUT3 #(
		.INIT('h0d)
	) name4314 (
		_w2246_,
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h4)
	) name4315 (
		_w5661_,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('hb)
	) name4316 (
		_w5660_,
		_w5665_,
		_w5666_
	);
	LUT3 #(
		.INIT('ha8)
	) name4317 (
		_w2580_,
		_w5476_,
		_w5477_,
		_w5667_
	);
	LUT3 #(
		.INIT('ha8)
	) name4318 (
		_w2606_,
		_w5480_,
		_w5481_,
		_w5668_
	);
	LUT3 #(
		.INIT('ha8)
	) name4319 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5667_,
		_w5668_,
		_w5669_
	);
	LUT3 #(
		.INIT('h02)
	) name4320 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w2250_,
		_w2349_,
		_w5670_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4321 (
		_w2350_,
		_w5485_,
		_w5486_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h1)
	) name4322 (
		_w2659_,
		_w5671_,
		_w5672_
	);
	LUT3 #(
		.INIT('ha8)
	) name4323 (
		_w1679_,
		_w5669_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h2)
	) name4324 (
		_w2283_,
		_w5671_,
		_w5674_
	);
	LUT4 #(
		.INIT('hc055)
	) name4325 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2250_,
		_w5675_
	);
	LUT2 #(
		.INIT('h2)
	) name4326 (
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w2288_,
		_w5676_
	);
	LUT3 #(
		.INIT('h0d)
	) name4327 (
		_w2246_,
		_w5675_,
		_w5676_,
		_w5677_
	);
	LUT2 #(
		.INIT('h4)
	) name4328 (
		_w5674_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('hb)
	) name4329 (
		_w5673_,
		_w5678_,
		_w5679_
	);
	LUT3 #(
		.INIT('ha8)
	) name4330 (
		_w2606_,
		_w5476_,
		_w5477_,
		_w5680_
	);
	LUT3 #(
		.INIT('ha8)
	) name4331 (
		_w2349_,
		_w5480_,
		_w5481_,
		_w5681_
	);
	LUT3 #(
		.INIT('ha8)
	) name4332 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5680_,
		_w5681_,
		_w5682_
	);
	LUT3 #(
		.INIT('h02)
	) name4333 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w2250_,
		_w2264_,
		_w5683_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4334 (
		_w2279_,
		_w5485_,
		_w5486_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h1)
	) name4335 (
		_w2683_,
		_w5684_,
		_w5685_
	);
	LUT3 #(
		.INIT('ha8)
	) name4336 (
		_w1679_,
		_w5682_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h2)
	) name4337 (
		_w2283_,
		_w5684_,
		_w5687_
	);
	LUT4 #(
		.INIT('hc055)
	) name4338 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1484_,
		_w1489_,
		_w2264_,
		_w5688_
	);
	LUT2 #(
		.INIT('h2)
	) name4339 (
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w2288_,
		_w5689_
	);
	LUT3 #(
		.INIT('h0d)
	) name4340 (
		_w2246_,
		_w5688_,
		_w5689_,
		_w5690_
	);
	LUT2 #(
		.INIT('h4)
	) name4341 (
		_w5687_,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('hb)
	) name4342 (
		_w5686_,
		_w5691_,
		_w5692_
	);
	LUT3 #(
		.INIT('h08)
	) name4343 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5693_
	);
	LUT2 #(
		.INIT('h4)
	) name4344 (
		_w4336_,
		_w4343_,
		_w5694_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4345 (
		_w4329_,
		_w4331_,
		_w4336_,
		_w4343_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name4346 (
		_w4347_,
		_w4352_,
		_w5696_
	);
	LUT4 #(
		.INIT('h8000)
	) name4347 (
		_w4821_,
		_w4826_,
		_w5695_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h2)
	) name4348 (
		_w4366_,
		_w4369_,
		_w5698_
	);
	LUT3 #(
		.INIT('h6c)
	) name4349 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4278_,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name4350 (
		_w4357_,
		_w4362_,
		_w5700_
	);
	LUT4 #(
		.INIT('h0200)
	) name4351 (
		_w4366_,
		_w4369_,
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT4 #(
		.INIT('h870f)
	) name4352 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w4278_,
		_w5702_
	);
	LUT4 #(
		.INIT('h1540)
	) name4353 (
		_w4214_,
		_w5697_,
		_w5701_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w5704_
	);
	LUT2 #(
		.INIT('h8)
	) name4355 (
		_w4275_,
		_w5704_,
		_w5705_
	);
	LUT4 #(
		.INIT('h8000)
	) name4356 (
		_w4796_,
		_w4896_,
		_w4900_,
		_w5705_,
		_w5706_
	);
	LUT4 #(
		.INIT('h8000)
	) name4357 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4272_,
		_w5704_,
		_w5707_
	);
	LUT2 #(
		.INIT('h6)
	) name4358 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w5707_,
		_w5708_
	);
	LUT4 #(
		.INIT('h1551)
	) name4359 (
		_w1661_,
		_w4214_,
		_w5706_,
		_w5708_,
		_w5709_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4360 (
		_w1559_,
		_w5693_,
		_w5703_,
		_w5709_,
		_w5710_
	);
	LUT4 #(
		.INIT('h028a)
	) name4361 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w5711_
	);
	LUT2 #(
		.INIT('h8)
	) name4362 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_InstAddrPointer_reg[18]/NET0131 ,
		_w5712_
	);
	LUT3 #(
		.INIT('h60)
	) name4363 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4410_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h8)
	) name4364 (
		_w4413_,
		_w5713_,
		_w5714_
	);
	LUT4 #(
		.INIT('h4000)
	) name4365 (
		_w4400_,
		_w4832_,
		_w4838_,
		_w5714_,
		_w5715_
	);
	LUT3 #(
		.INIT('h80)
	) name4366 (
		_w4876_,
		_w4915_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h8)
	) name4367 (
		_w4427_,
		_w5704_,
		_w5717_
	);
	LUT4 #(
		.INIT('h8000)
	) name4368 (
		_w4876_,
		_w4915_,
		_w5715_,
		_w5717_,
		_w5718_
	);
	LUT4 #(
		.INIT('h9333)
	) name4369 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w4425_,
		_w5704_,
		_w5719_
	);
	LUT4 #(
		.INIT('h1331)
	) name4370 (
		_w1659_,
		_w5711_,
		_w5718_,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w5721_
	);
	LUT3 #(
		.INIT('h80)
	) name4372 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w5722_
	);
	LUT4 #(
		.INIT('h8000)
	) name4373 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5723_
	);
	LUT3 #(
		.INIT('h80)
	) name4374 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5723_,
		_w5724_
	);
	LUT4 #(
		.INIT('h8000)
	) name4375 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w5723_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name4376 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w5726_
	);
	LUT3 #(
		.INIT('h80)
	) name4377 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h8)
	) name4378 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w5728_
	);
	LUT3 #(
		.INIT('h80)
	) name4379 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w5729_
	);
	LUT4 #(
		.INIT('h8000)
	) name4380 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w5729_,
		_w5730_
	);
	LUT3 #(
		.INIT('h80)
	) name4381 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w5731_
	);
	LUT3 #(
		.INIT('h80)
	) name4382 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w5730_,
		_w5731_,
		_w5732_
	);
	LUT4 #(
		.INIT('h8000)
	) name4383 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w5730_,
		_w5731_,
		_w5733_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w5734_
	);
	LUT3 #(
		.INIT('h80)
	) name4385 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w5734_,
		_w5735_
	);
	LUT4 #(
		.INIT('h8000)
	) name4386 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w5733_,
		_w5734_,
		_w5736_
	);
	LUT3 #(
		.INIT('h80)
	) name4387 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5736_,
		_w5737_
	);
	LUT4 #(
		.INIT('h8000)
	) name4388 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w5736_,
		_w5738_
	);
	LUT4 #(
		.INIT('h8000)
	) name4389 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5738_,
		_w5739_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4390 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w2242_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name4391 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5741_
	);
	LUT2 #(
		.INIT('h8)
	) name4392 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5742_
	);
	LUT4 #(
		.INIT('h8000)
	) name4393 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5736_,
		_w5741_,
		_w5742_,
		_w5743_
	);
	LUT3 #(
		.INIT('h80)
	) name4394 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5743_,
		_w5744_
	);
	LUT4 #(
		.INIT('h8000)
	) name4395 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w5743_,
		_w5745_
	);
	LUT3 #(
		.INIT('h0d)
	) name4396 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w2283_,
		_w2298_,
		_w5746_
	);
	LUT4 #(
		.INIT('hfc35)
	) name4397 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w5747_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4398 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2286_,
		_w5747_,
		_w5748_
	);
	LUT4 #(
		.INIT('h9f00)
	) name4399 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w5746_,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h4)
	) name4400 (
		_w5740_,
		_w5749_,
		_w5750_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4401 (
		_w1678_,
		_w5710_,
		_w5720_,
		_w5750_,
		_w5751_
	);
	LUT3 #(
		.INIT('h02)
	) name4402 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w2103_,
		_w2172_,
		_w5752_
	);
	LUT4 #(
		.INIT('haa20)
	) name4403 (
		_w2171_,
		_w2916_,
		_w2982_,
		_w5752_,
		_w5753_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4404 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w5754_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4405 (
		_w2181_,
		_w3046_,
		_w3047_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h8)
	) name4406 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5756_
	);
	LUT3 #(
		.INIT('h80)
	) name4407 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w5757_
	);
	LUT4 #(
		.INIT('h8000)
	) name4408 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w5758_
	);
	LUT3 #(
		.INIT('h80)
	) name4409 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5758_,
		_w5759_
	);
	LUT4 #(
		.INIT('h8000)
	) name4410 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w5758_,
		_w5760_
	);
	LUT3 #(
		.INIT('h80)
	) name4411 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w5761_
	);
	LUT4 #(
		.INIT('h8000)
	) name4412 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w5762_
	);
	LUT3 #(
		.INIT('h80)
	) name4413 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h8)
	) name4414 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w5764_
	);
	LUT3 #(
		.INIT('h80)
	) name4415 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w5765_
	);
	LUT4 #(
		.INIT('h8000)
	) name4416 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5762_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h8)
	) name4417 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h8)
	) name4418 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w5768_
	);
	LUT3 #(
		.INIT('h80)
	) name4419 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w5769_
	);
	LUT3 #(
		.INIT('h80)
	) name4420 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5766_,
		_w5769_,
		_w5770_
	);
	LUT4 #(
		.INIT('h8000)
	) name4421 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w5766_,
		_w5769_,
		_w5771_
	);
	LUT2 #(
		.INIT('h8)
	) name4422 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5772_
	);
	LUT3 #(
		.INIT('h80)
	) name4423 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w5773_
	);
	LUT4 #(
		.INIT('h8000)
	) name4424 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5774_
	);
	LUT4 #(
		.INIT('h8000)
	) name4425 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w5774_,
		_w5775_
	);
	LUT4 #(
		.INIT('h8000)
	) name4426 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w5756_,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('h8000)
	) name4427 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w5771_,
		_w5774_,
		_w5777_
	);
	LUT3 #(
		.INIT('h80)
	) name4428 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w5756_,
		_w5777_,
		_w5778_
	);
	LUT4 #(
		.INIT('hd1f3)
	) name4429 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5776_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w5780_
	);
	LUT4 #(
		.INIT('h9333)
	) name4431 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		_w5756_,
		_w5777_,
		_w5781_
	);
	LUT4 #(
		.INIT('h048c)
	) name4432 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w5779_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('hfc35)
	) name4433 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w5783_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4434 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w3054_,
		_w5783_,
		_w5784_
	);
	LUT3 #(
		.INIT('hd0)
	) name4435 (
		_w3055_,
		_w5779_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h4)
	) name4436 (
		_w5782_,
		_w5785_,
		_w5786_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4437 (
		_w1945_,
		_w5753_,
		_w5755_,
		_w5786_,
		_w5787_
	);
	LUT3 #(
		.INIT('h08)
	) name4438 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2988_,
		_w4088_,
		_w5788_
	);
	LUT4 #(
		.INIT('h0080)
	) name4439 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2987_,
		_w2988_,
		_w4088_,
		_w5789_
	);
	LUT3 #(
		.INIT('h80)
	) name4440 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w5789_,
		_w5790_
	);
	LUT3 #(
		.INIT('h6c)
	) name4441 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2986_,
		_w5791_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name4442 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2181_,
		_w5791_,
		_w5789_,
		_w5792_
	);
	LUT2 #(
		.INIT('h4)
	) name4443 (
		_w5790_,
		_w5792_,
		_w5793_
	);
	LUT3 #(
		.INIT('h02)
	) name4444 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2103_,
		_w2172_,
		_w5794_
	);
	LUT4 #(
		.INIT('h2822)
	) name4445 (
		_w2755_,
		_w2942_,
		_w4051_,
		_w4054_,
		_w5795_
	);
	LUT2 #(
		.INIT('h4)
	) name4446 (
		_w2876_,
		_w4067_,
		_w5796_
	);
	LUT3 #(
		.INIT('h2a)
	) name4447 (
		_w2878_,
		_w4074_,
		_w5796_,
		_w5797_
	);
	LUT3 #(
		.INIT('h15)
	) name4448 (
		_w2755_,
		_w4068_,
		_w4074_,
		_w5798_
	);
	LUT4 #(
		.INIT('h0045)
	) name4449 (
		_w2173_,
		_w5797_,
		_w5798_,
		_w5795_,
		_w5799_
	);
	LUT3 #(
		.INIT('h80)
	) name4450 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2060_,
		_w2044_,
		_w5800_
	);
	LUT4 #(
		.INIT('h000c)
	) name4451 (
		_w2112_,
		_w2114_,
		_w2108_,
		_w5800_,
		_w5801_
	);
	LUT4 #(
		.INIT('h00e4)
	) name4452 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2112_,
		_w5802_
	);
	LUT2 #(
		.INIT('h1)
	) name4453 (
		_w2116_,
		_w2942_,
		_w5803_
	);
	LUT2 #(
		.INIT('h4)
	) name4454 (
		_w5802_,
		_w5803_,
		_w5804_
	);
	LUT4 #(
		.INIT('h4440)
	) name4455 (
		_w2136_,
		_w2176_,
		_w5801_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name4456 (
		_w2108_,
		_w2115_,
		_w2116_,
		_w5800_,
		_w5806_
	);
	LUT3 #(
		.INIT('hc8)
	) name4457 (
		_w2064_,
		_w2942_,
		_w5806_,
		_w5807_
	);
	LUT4 #(
		.INIT('h64cc)
	) name4458 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w2098_,
		_w2986_,
		_w5808_
	);
	LUT3 #(
		.INIT('he0)
	) name4459 (
		_w2071_,
		_w2087_,
		_w5808_,
		_w5809_
	);
	LUT4 #(
		.INIT('h004f)
	) name4460 (
		_w2073_,
		_w2086_,
		_w2878_,
		_w5809_,
		_w5810_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4461 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		_w5805_,
		_w5807_,
		_w5810_,
		_w5811_
	);
	LUT4 #(
		.INIT('h5700)
	) name4462 (
		_w2171_,
		_w5794_,
		_w5799_,
		_w5811_,
		_w5812_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4463 (
		\P3_InstAddrPointer_reg[12]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w3054_,
		_w3056_,
		_w5813_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4464 (
		_w1945_,
		_w5793_,
		_w5812_,
		_w5813_,
		_w5814_
	);
	LUT3 #(
		.INIT('h82)
	) name4465 (
		_w2755_,
		_w2944_,
		_w4051_,
		_w5815_
	);
	LUT3 #(
		.INIT('h54)
	) name4466 (
		_w2844_,
		_w2860_,
		_w2861_,
		_w5816_
	);
	LUT3 #(
		.INIT('h07)
	) name4467 (
		_w2749_,
		_w2754_,
		_w2757_,
		_w5817_
	);
	LUT4 #(
		.INIT('h0b00)
	) name4468 (
		_w2831_,
		_w2858_,
		_w5816_,
		_w5817_,
		_w5818_
	);
	LUT4 #(
		.INIT('hc8fb)
	) name4469 (
		_w2755_,
		_w2864_,
		_w4074_,
		_w5818_,
		_w5819_
	);
	LUT4 #(
		.INIT('h4744)
	) name4470 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2173_,
		_w5815_,
		_w5819_,
		_w5820_
	);
	LUT3 #(
		.INIT('h82)
	) name4471 (
		_w2181_,
		_w2988_,
		_w4088_,
		_w5821_
	);
	LUT3 #(
		.INIT('h21)
	) name4472 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2116_,
		_w2715_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w2137_,
		_w5822_,
		_w5823_
	);
	LUT4 #(
		.INIT('h0010)
	) name4474 (
		_w2127_,
		_w4784_,
		_w4785_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h4)
	) name4475 (
		_w2117_,
		_w2944_,
		_w5825_
	);
	LUT3 #(
		.INIT('he0)
	) name4476 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w2098_,
		_w2988_,
		_w5826_
	);
	LUT3 #(
		.INIT('he0)
	) name4477 (
		_w2071_,
		_w2087_,
		_w5826_,
		_w5827_
	);
	LUT4 #(
		.INIT('h004f)
	) name4478 (
		_w2073_,
		_w2086_,
		_w2864_,
		_w5827_,
		_w5828_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4479 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		_w5824_,
		_w5825_,
		_w5828_,
		_w5829_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4480 (
		_w2171_,
		_w5820_,
		_w5821_,
		_w5829_,
		_w5830_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4481 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w3054_,
		_w3056_,
		_w5831_
	);
	LUT3 #(
		.INIT('h2f)
	) name4482 (
		_w1945_,
		_w5830_,
		_w5831_,
		_w5832_
	);
	LUT3 #(
		.INIT('h08)
	) name4483 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5833_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4484 (
		_w4216_,
		_w4201_,
		_w4220_,
		_w4809_,
		_w5834_
	);
	LUT2 #(
		.INIT('h1)
	) name4485 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w4227_,
		_w5835_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		_w4237_,
		_w5835_,
		_w5836_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4487 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4223_,
		_w4807_,
		_w5836_,
		_w5837_
	);
	LUT3 #(
		.INIT('ha8)
	) name4488 (
		_w4214_,
		_w5834_,
		_w5837_,
		_w5838_
	);
	LUT4 #(
		.INIT('he0f0)
	) name4489 (
		_w4315_,
		_w4321_,
		_w4322_,
		_w4818_,
		_w5839_
	);
	LUT4 #(
		.INIT('h4555)
	) name4490 (
		_w4214_,
		_w4315_,
		_w4323_,
		_w4818_,
		_w5840_
	);
	LUT3 #(
		.INIT('h45)
	) name4491 (
		_w1661_,
		_w5839_,
		_w5840_,
		_w5841_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4492 (
		_w1559_,
		_w5833_,
		_w5838_,
		_w5841_,
		_w5842_
	);
	LUT4 #(
		.INIT('ha028)
	) name4493 (
		_w1659_,
		_w4405_,
		_w4407_,
		_w4869_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		_w1640_,
		_w4407_,
		_w5844_
	);
	LUT4 #(
		.INIT('h004f)
	) name4495 (
		_w1571_,
		_w1583_,
		_w4322_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h4)
	) name4496 (
		_w1617_,
		_w5836_,
		_w5846_
	);
	LUT3 #(
		.INIT('h2a)
	) name4497 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		_w1658_,
		_w4844_,
		_w5847_
	);
	LUT4 #(
		.INIT('h0100)
	) name4498 (
		_w5843_,
		_w5846_,
		_w5847_,
		_w5845_,
		_w5848_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4499 (
		\P2_InstAddrPointer_reg[10]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5849_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4500 (
		_w1678_,
		_w5842_,
		_w5848_,
		_w5849_,
		_w5850_
	);
	LUT3 #(
		.INIT('h08)
	) name4501 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w1842_,
		_w1915_,
		_w5851_
	);
	LUT4 #(
		.INIT('h00f8)
	) name4502 (
		_w3267_,
		_w3296_,
		_w3309_,
		_w4447_,
		_w5852_
	);
	LUT4 #(
		.INIT('h4554)
	) name4503 (
		_w1916_,
		_w3101_,
		_w3090_,
		_w3214_,
		_w5853_
	);
	LUT4 #(
		.INIT('h0233)
	) name4504 (
		_w3101_,
		_w5851_,
		_w5852_,
		_w5853_,
		_w5854_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4505 (
		_w1924_,
		_w3356_,
		_w3359_,
		_w3360_,
		_w5855_
	);
	LUT3 #(
		.INIT('h2a)
	) name4506 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w1922_,
		_w4037_,
		_w5856_
	);
	LUT2 #(
		.INIT('h4)
	) name4507 (
		_w1862_,
		_w3309_,
		_w5857_
	);
	LUT3 #(
		.INIT('h40)
	) name4508 (
		_w1833_,
		_w1846_,
		_w3360_,
		_w5858_
	);
	LUT4 #(
		.INIT('h004f)
	) name4509 (
		_w1816_,
		_w1831_,
		_w3090_,
		_w5858_,
		_w5859_
	);
	LUT4 #(
		.INIT('h0100)
	) name4510 (
		_w5855_,
		_w5857_,
		_w5856_,
		_w5859_,
		_w5860_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4511 (
		_w1810_,
		_w1933_,
		_w5854_,
		_w5860_,
		_w5861_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4512 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w3406_,
		_w3408_,
		_w5862_
	);
	LUT2 #(
		.INIT('hb)
	) name4513 (
		_w5861_,
		_w5862_,
		_w5863_
	);
	LUT3 #(
		.INIT('h08)
	) name4514 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5864_
	);
	LUT3 #(
		.INIT('h15)
	) name4515 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4225_,
		_w4227_,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name4516 (
		_w4239_,
		_w5865_,
		_w5866_
	);
	LUT4 #(
		.INIT('hf700)
	) name4517 (
		_w4223_,
		_w4229_,
		_w4807_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h0008)
	) name4518 (
		_w4223_,
		_w4229_,
		_w4807_,
		_w5866_,
		_w5868_
	);
	LUT3 #(
		.INIT('h02)
	) name4519 (
		_w4214_,
		_w5868_,
		_w5867_,
		_w5869_
	);
	LUT3 #(
		.INIT('h2a)
	) name4520 (
		_w4319_,
		_w4818_,
		_w4903_,
		_w5870_
	);
	LUT4 #(
		.INIT('h4555)
	) name4521 (
		_w4214_,
		_w4315_,
		_w4325_,
		_w4818_,
		_w5871_
	);
	LUT3 #(
		.INIT('h45)
	) name4522 (
		_w1661_,
		_w5870_,
		_w5871_,
		_w5872_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4523 (
		_w1559_,
		_w5864_,
		_w5869_,
		_w5872_,
		_w5873_
	);
	LUT3 #(
		.INIT('h6c)
	) name4524 (
		\P2_InstAddrPointer_reg[11]/NET0131 ,
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w4406_,
		_w5874_
	);
	LUT4 #(
		.INIT('h2000)
	) name4525 (
		_w4236_,
		_w4401_,
		_w4403_,
		_w4836_,
		_w5875_
	);
	LUT4 #(
		.INIT('h82a0)
	) name4526 (
		_w1659_,
		_w4869_,
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4527 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w4835_,
		_w5877_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4528 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		_w1658_,
		_w4844_,
		_w5877_,
		_w5878_
	);
	LUT3 #(
		.INIT('hb0)
	) name4529 (
		_w1571_,
		_w1583_,
		_w4319_,
		_w5879_
	);
	LUT2 #(
		.INIT('h8)
	) name4530 (
		_w1640_,
		_w5874_,
		_w5880_
	);
	LUT3 #(
		.INIT('h0b)
	) name4531 (
		_w1617_,
		_w5866_,
		_w5880_,
		_w5881_
	);
	LUT4 #(
		.INIT('h0100)
	) name4532 (
		_w5876_,
		_w5878_,
		_w5879_,
		_w5881_,
		_w5882_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4533 (
		\P2_InstAddrPointer_reg[12]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5883_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4534 (
		_w1678_,
		_w5873_,
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT3 #(
		.INIT('h08)
	) name4535 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w1592_,
		_w1660_,
		_w5885_
	);
	LUT4 #(
		.INIT('he0ee)
	) name4536 (
		_w4231_,
		_w4242_,
		_w4807_,
		_w4810_,
		_w5886_
	);
	LUT2 #(
		.INIT('h2)
	) name4537 (
		_w4214_,
		_w5886_,
		_w5887_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4538 (
		_w4308_,
		_w4317_,
		_w4325_,
		_w4337_,
		_w5888_
	);
	LUT4 #(
		.INIT('h1555)
	) name4539 (
		_w4214_,
		_w4818_,
		_w4819_,
		_w4903_,
		_w5889_
	);
	LUT3 #(
		.INIT('h45)
	) name4540 (
		_w1661_,
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4541 (
		_w1559_,
		_w5885_,
		_w5887_,
		_w5890_,
		_w5891_
	);
	LUT4 #(
		.INIT('h00bf)
	) name4542 (
		_w4400_,
		_w4405_,
		_w4408_,
		_w4833_,
		_w5892_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4543 (
		_w1659_,
		_w4400_,
		_w4405_,
		_w4409_,
		_w5893_
	);
	LUT2 #(
		.INIT('h4)
	) name4544 (
		_w5892_,
		_w5893_,
		_w5894_
	);
	LUT4 #(
		.INIT('he000)
	) name4545 (
		_w1592_,
		_w1595_,
		_w4238_,
		_w4406_,
		_w5895_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4546 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w5895_,
		_w5896_
	);
	LUT2 #(
		.INIT('h8)
	) name4547 (
		_w4833_,
		_w5896_,
		_w5897_
	);
	LUT3 #(
		.INIT('h0b)
	) name4548 (
		_w1617_,
		_w4242_,
		_w5897_,
		_w5898_
	);
	LUT3 #(
		.INIT('hb0)
	) name4549 (
		_w1571_,
		_w1583_,
		_w4337_,
		_w5899_
	);
	LUT3 #(
		.INIT('h2a)
	) name4550 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		_w1658_,
		_w4844_,
		_w5900_
	);
	LUT3 #(
		.INIT('h10)
	) name4551 (
		_w5899_,
		_w5900_,
		_w5898_,
		_w5901_
	);
	LUT2 #(
		.INIT('h4)
	) name4552 (
		_w5894_,
		_w5901_,
		_w5902_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4553 (
		\P2_InstAddrPointer_reg[13]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w2286_,
		_w4441_,
		_w5903_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4554 (
		_w1678_,
		_w5891_,
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT3 #(
		.INIT('h82)
	) name4555 (
		_w3101_,
		_w4463_,
		_w4464_,
		_w5905_
	);
	LUT4 #(
		.INIT('h4111)
	) name4556 (
		_w3101_,
		_w3221_,
		_w4724_,
		_w4725_,
		_w5906_
	);
	LUT4 #(
		.INIT('h7774)
	) name4557 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1916_,
		_w5906_,
		_w5905_,
		_w5907_
	);
	LUT4 #(
		.INIT('h2000)
	) name4558 (
		\P1_InstAddrPointer_reg[10]/NET0131 ,
		_w3356_,
		_w3359_,
		_w3362_,
		_w5908_
	);
	LUT4 #(
		.INIT('h4448)
	) name4559 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1924_,
		_w3361_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h4)
	) name4560 (
		_w1862_,
		_w4464_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w1877_,
		_w1913_,
		_w5911_
	);
	LUT3 #(
		.INIT('h2a)
	) name4562 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1922_,
		_w5911_,
		_w5912_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name4563 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w1842_,
		_w1845_,
		_w3361_,
		_w5913_
	);
	LUT2 #(
		.INIT('h4)
	) name4564 (
		_w1833_,
		_w5913_,
		_w5914_
	);
	LUT4 #(
		.INIT('h004f)
	) name4565 (
		_w1816_,
		_w1831_,
		_w3221_,
		_w5914_,
		_w5915_
	);
	LUT3 #(
		.INIT('h10)
	) name4566 (
		_w5912_,
		_w5910_,
		_w5915_,
		_w5916_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4567 (
		_w1810_,
		_w5907_,
		_w5909_,
		_w5916_,
		_w5917_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4568 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w3406_,
		_w3408_,
		_w5918_
	);
	LUT3 #(
		.INIT('h2f)
	) name4569 (
		_w1933_,
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT4 #(
		.INIT('h1444)
	) name4570 (
		_w3101_,
		_w3245_,
		_w4011_,
		_w5451_,
		_w5920_
	);
	LUT4 #(
		.INIT('h28a0)
	) name4571 (
		_w3101_,
		_w3296_,
		_w3991_,
		_w3995_,
		_w5921_
	);
	LUT4 #(
		.INIT('h4447)
	) name4572 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1916_,
		_w5920_,
		_w5921_,
		_w5922_
	);
	LUT2 #(
		.INIT('h6)
	) name4573 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w3366_,
		_w5923_
	);
	LUT4 #(
		.INIT('h2000)
	) name4574 (
		_w3368_,
		_w4023_,
		_w4025_,
		_w4028_,
		_w5924_
	);
	LUT4 #(
		.INIT('h4448)
	) name4575 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1924_,
		_w3366_,
		_w5924_,
		_w5925_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		_w1833_,
		_w3366_,
		_w5926_
	);
	LUT3 #(
		.INIT('ha2)
	) name4577 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w4037_,
		_w5926_,
		_w5927_
	);
	LUT3 #(
		.INIT('h65)
	) name4578 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1861_,
		_w3072_,
		_w5928_
	);
	LUT4 #(
		.INIT('h00ec)
	) name4579 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w5928_,
		_w5929_
	);
	LUT4 #(
		.INIT('h5655)
	) name4580 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		_w1858_,
		_w1861_,
		_w3072_,
		_w5930_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4581 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w5930_,
		_w5931_
	);
	LUT3 #(
		.INIT('h54)
	) name4582 (
		_w1852_,
		_w5929_,
		_w5931_,
		_w5932_
	);
	LUT3 #(
		.INIT('h80)
	) name4583 (
		_w1805_,
		_w1806_,
		_w3991_,
		_w5933_
	);
	LUT4 #(
		.INIT('h00bf)
	) name4584 (
		_w1833_,
		_w1846_,
		_w5923_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4585 (
		_w1816_,
		_w1831_,
		_w3245_,
		_w5934_,
		_w5935_
	);
	LUT3 #(
		.INIT('h10)
	) name4586 (
		_w5927_,
		_w5932_,
		_w5935_,
		_w5936_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4587 (
		_w1810_,
		_w5922_,
		_w5925_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4588 (
		\P1_InstAddrPointer_reg[17]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w3406_,
		_w3408_,
		_w5938_
	);
	LUT3 #(
		.INIT('h2f)
	) name4589 (
		_w1933_,
		_w5937_,
		_w5938_,
		_w5939_
	);
	LUT4 #(
		.INIT('h02fd)
	) name4590 (
		_w3523_,
		_w3526_,
		_w3529_,
		_w4502_,
		_w5940_
	);
	LUT4 #(
		.INIT('h2822)
	) name4591 (
		_w3412_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w5941_
	);
	LUT4 #(
		.INIT('haa80)
	) name4592 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3411_,
		_w5940_,
		_w5941_,
		_w5942_
	);
	LUT3 #(
		.INIT('h02)
	) name4593 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w3534_,
		_w3536_,
		_w5943_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4594 (
		_w3537_,
		_w3450_,
		_w3451_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h1)
	) name4595 (
		_w3414_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w3407_,
		_w5944_,
		_w5946_
	);
	LUT4 #(
		.INIT('hc055)
	) name4597 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3534_,
		_w5947_
	);
	LUT2 #(
		.INIT('h2)
	) name4598 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		_w3545_,
		_w5948_
	);
	LUT3 #(
		.INIT('h0d)
	) name4599 (
		_w2248_,
		_w5947_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h4)
	) name4600 (
		_w5946_,
		_w5949_,
		_w5950_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4601 (
		_w1939_,
		_w5942_,
		_w5945_,
		_w5950_,
		_w5951_
	);
	LUT3 #(
		.INIT('h82)
	) name4602 (
		_w3411_,
		_w4503_,
		_w4506_,
		_w5952_
	);
	LUT4 #(
		.INIT('h5655)
	) name4603 (
		_w3503_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w5953_
	);
	LUT2 #(
		.INIT('h8)
	) name4604 (
		_w3412_,
		_w5953_,
		_w5954_
	);
	LUT3 #(
		.INIT('h02)
	) name4605 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w3534_,
		_w3536_,
		_w5955_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4606 (
		_w3537_,
		_w3472_,
		_w3473_,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h1)
	) name4607 (
		_w3414_,
		_w5956_,
		_w5957_
	);
	LUT4 #(
		.INIT('h0057)
	) name4608 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5952_,
		_w5954_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h2)
	) name4609 (
		_w3407_,
		_w5956_,
		_w5959_
	);
	LUT4 #(
		.INIT('hc055)
	) name4610 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3534_,
		_w5960_
	);
	LUT2 #(
		.INIT('h2)
	) name4611 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w3545_,
		_w5961_
	);
	LUT3 #(
		.INIT('h0d)
	) name4612 (
		_w2248_,
		_w5960_,
		_w5961_,
		_w5962_
	);
	LUT2 #(
		.INIT('h4)
	) name4613 (
		_w5959_,
		_w5962_,
		_w5963_
	);
	LUT3 #(
		.INIT('h2f)
	) name4614 (
		_w1939_,
		_w5958_,
		_w5963_,
		_w5964_
	);
	LUT4 #(
		.INIT('h6500)
	) name4615 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3573_,
		_w5965_
	);
	LUT4 #(
		.INIT('haa80)
	) name4616 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3572_,
		_w5940_,
		_w5965_,
		_w5966_
	);
	LUT3 #(
		.INIT('h02)
	) name4617 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w3578_,
		_w3580_,
		_w5967_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4618 (
		_w3450_,
		_w3451_,
		_w3581_,
		_w5967_,
		_w5968_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w3575_,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		_w3407_,
		_w5968_,
		_w5970_
	);
	LUT4 #(
		.INIT('hc055)
	) name4621 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3578_,
		_w5971_
	);
	LUT2 #(
		.INIT('h2)
	) name4622 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		_w3545_,
		_w5972_
	);
	LUT3 #(
		.INIT('h0d)
	) name4623 (
		_w2248_,
		_w5971_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h4)
	) name4624 (
		_w5970_,
		_w5973_,
		_w5974_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4625 (
		_w1939_,
		_w5966_,
		_w5969_,
		_w5974_,
		_w5975_
	);
	LUT3 #(
		.INIT('h82)
	) name4626 (
		_w3572_,
		_w4503_,
		_w4506_,
		_w5976_
	);
	LUT2 #(
		.INIT('h8)
	) name4627 (
		_w3573_,
		_w5953_,
		_w5977_
	);
	LUT3 #(
		.INIT('h02)
	) name4628 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w3578_,
		_w3580_,
		_w5978_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4629 (
		_w3472_,
		_w3473_,
		_w3581_,
		_w5978_,
		_w5979_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w3575_,
		_w5979_,
		_w5980_
	);
	LUT4 #(
		.INIT('h0057)
	) name4631 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5976_,
		_w5977_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h2)
	) name4632 (
		_w3407_,
		_w5979_,
		_w5982_
	);
	LUT4 #(
		.INIT('hc055)
	) name4633 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3578_,
		_w5983_
	);
	LUT2 #(
		.INIT('h2)
	) name4634 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		_w3545_,
		_w5984_
	);
	LUT3 #(
		.INIT('h0d)
	) name4635 (
		_w2248_,
		_w5983_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h4)
	) name4636 (
		_w5982_,
		_w5985_,
		_w5986_
	);
	LUT3 #(
		.INIT('h2f)
	) name4637 (
		_w1939_,
		_w5981_,
		_w5986_,
		_w5987_
	);
	LUT4 #(
		.INIT('h2822)
	) name4638 (
		_w3411_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w5988_
	);
	LUT4 #(
		.INIT('haa80)
	) name4639 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3592_,
		_w5940_,
		_w5988_,
		_w5989_
	);
	LUT3 #(
		.INIT('h02)
	) name4640 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		_w3536_,
		_w3412_,
		_w5990_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4641 (
		_w3450_,
		_w3451_,
		_w3597_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w3594_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		_w3407_,
		_w5991_,
		_w5993_
	);
	LUT4 #(
		.INIT('hc055)
	) name4644 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3536_,
		_w5994_
	);
	LUT2 #(
		.INIT('h2)
	) name4645 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		_w3545_,
		_w5995_
	);
	LUT3 #(
		.INIT('h0d)
	) name4646 (
		_w2248_,
		_w5994_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h4)
	) name4647 (
		_w5993_,
		_w5996_,
		_w5997_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4648 (
		_w1939_,
		_w5989_,
		_w5992_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h8)
	) name4649 (
		_w3411_,
		_w5953_,
		_w5999_
	);
	LUT3 #(
		.INIT('h82)
	) name4650 (
		_w3592_,
		_w4503_,
		_w4506_,
		_w6000_
	);
	LUT3 #(
		.INIT('h02)
	) name4651 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		_w3536_,
		_w3412_,
		_w6001_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4652 (
		_w3472_,
		_w3473_,
		_w3597_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h1)
	) name4653 (
		_w3594_,
		_w6002_,
		_w6003_
	);
	LUT4 #(
		.INIT('h0057)
	) name4654 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w5999_,
		_w6000_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		_w3407_,
		_w6002_,
		_w6005_
	);
	LUT4 #(
		.INIT('hc055)
	) name4656 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3536_,
		_w6006_
	);
	LUT2 #(
		.INIT('h2)
	) name4657 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		_w3545_,
		_w6007_
	);
	LUT3 #(
		.INIT('h0d)
	) name4658 (
		_w2248_,
		_w6006_,
		_w6007_,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name4659 (
		_w6005_,
		_w6008_,
		_w6009_
	);
	LUT3 #(
		.INIT('h2f)
	) name4660 (
		_w1939_,
		_w6004_,
		_w6009_,
		_w6010_
	);
	LUT4 #(
		.INIT('h2822)
	) name4661 (
		_w3536_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w6011_
	);
	LUT4 #(
		.INIT('haa80)
	) name4662 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3412_,
		_w5940_,
		_w6011_,
		_w6012_
	);
	LUT3 #(
		.INIT('h02)
	) name4663 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w3534_,
		_w3611_,
		_w6013_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4664 (
		_w3450_,
		_w3451_,
		_w3612_,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w3608_,
		_w6014_,
		_w6015_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w3407_,
		_w6014_,
		_w6016_
	);
	LUT4 #(
		.INIT('hc055)
	) name4667 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3611_,
		_w6017_
	);
	LUT2 #(
		.INIT('h2)
	) name4668 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w3545_,
		_w6018_
	);
	LUT3 #(
		.INIT('h0d)
	) name4669 (
		_w2248_,
		_w6017_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h4)
	) name4670 (
		_w6016_,
		_w6019_,
		_w6020_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4671 (
		_w1939_,
		_w6012_,
		_w6015_,
		_w6020_,
		_w6021_
	);
	LUT3 #(
		.INIT('h82)
	) name4672 (
		_w3412_,
		_w4503_,
		_w4506_,
		_w6022_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		_w3536_,
		_w5953_,
		_w6023_
	);
	LUT3 #(
		.INIT('h02)
	) name4674 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w3534_,
		_w3611_,
		_w6024_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4675 (
		_w3472_,
		_w3473_,
		_w3612_,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name4676 (
		_w3608_,
		_w6025_,
		_w6026_
	);
	LUT4 #(
		.INIT('h0057)
	) name4677 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6022_,
		_w6023_,
		_w6026_,
		_w6027_
	);
	LUT2 #(
		.INIT('h2)
	) name4678 (
		_w3407_,
		_w6025_,
		_w6028_
	);
	LUT4 #(
		.INIT('hc055)
	) name4679 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3611_,
		_w6029_
	);
	LUT2 #(
		.INIT('h2)
	) name4680 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w3545_,
		_w6030_
	);
	LUT3 #(
		.INIT('h0d)
	) name4681 (
		_w2248_,
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h4)
	) name4682 (
		_w6028_,
		_w6031_,
		_w6032_
	);
	LUT3 #(
		.INIT('h2f)
	) name4683 (
		_w1939_,
		_w6027_,
		_w6032_,
		_w6033_
	);
	LUT4 #(
		.INIT('h2822)
	) name4684 (
		_w3534_,
		_w3510_,
		_w3496_,
		_w3532_,
		_w6034_
	);
	LUT4 #(
		.INIT('haa80)
	) name4685 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3536_,
		_w5940_,
		_w6034_,
		_w6035_
	);
	LUT3 #(
		.INIT('h02)
	) name4686 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w3572_,
		_w3611_,
		_w6036_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4687 (
		_w3450_,
		_w3451_,
		_w3626_,
		_w6036_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name4688 (
		_w3623_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h2)
	) name4689 (
		_w3407_,
		_w6037_,
		_w6039_
	);
	LUT4 #(
		.INIT('hc055)
	) name4690 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3572_,
		_w6040_
	);
	LUT2 #(
		.INIT('h2)
	) name4691 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		_w3545_,
		_w6041_
	);
	LUT3 #(
		.INIT('h0d)
	) name4692 (
		_w2248_,
		_w6040_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h4)
	) name4693 (
		_w6039_,
		_w6042_,
		_w6043_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4694 (
		_w1939_,
		_w6035_,
		_w6038_,
		_w6043_,
		_w6044_
	);
	LUT3 #(
		.INIT('h82)
	) name4695 (
		_w3536_,
		_w4503_,
		_w4506_,
		_w6045_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		_w3534_,
		_w5953_,
		_w6046_
	);
	LUT3 #(
		.INIT('h02)
	) name4697 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w3572_,
		_w3611_,
		_w6047_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4698 (
		_w3472_,
		_w3473_,
		_w3626_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name4699 (
		_w3623_,
		_w6048_,
		_w6049_
	);
	LUT4 #(
		.INIT('h0057)
	) name4700 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6045_,
		_w6046_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h2)
	) name4701 (
		_w3407_,
		_w6048_,
		_w6051_
	);
	LUT4 #(
		.INIT('hc055)
	) name4702 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3572_,
		_w6052_
	);
	LUT2 #(
		.INIT('h2)
	) name4703 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w3545_,
		_w6053_
	);
	LUT3 #(
		.INIT('h0d)
	) name4704 (
		_w2248_,
		_w6052_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h4)
	) name4705 (
		_w6051_,
		_w6054_,
		_w6055_
	);
	LUT3 #(
		.INIT('h2f)
	) name4706 (
		_w1939_,
		_w6050_,
		_w6055_,
		_w6056_
	);
	LUT4 #(
		.INIT('h6500)
	) name4707 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3611_,
		_w6057_
	);
	LUT4 #(
		.INIT('haa80)
	) name4708 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3534_,
		_w5940_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('h02)
	) name4709 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w3572_,
		_w3573_,
		_w6059_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4710 (
		_w3450_,
		_w3451_,
		_w3574_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name4711 (
		_w3637_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h2)
	) name4712 (
		_w3407_,
		_w6060_,
		_w6062_
	);
	LUT4 #(
		.INIT('hc055)
	) name4713 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3573_,
		_w6063_
	);
	LUT2 #(
		.INIT('h2)
	) name4714 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w3545_,
		_w6064_
	);
	LUT3 #(
		.INIT('h0d)
	) name4715 (
		_w2248_,
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h4)
	) name4716 (
		_w6062_,
		_w6065_,
		_w6066_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4717 (
		_w1939_,
		_w6058_,
		_w6061_,
		_w6066_,
		_w6067_
	);
	LUT3 #(
		.INIT('h82)
	) name4718 (
		_w3534_,
		_w4503_,
		_w4506_,
		_w6068_
	);
	LUT2 #(
		.INIT('h8)
	) name4719 (
		_w3611_,
		_w5953_,
		_w6069_
	);
	LUT3 #(
		.INIT('h02)
	) name4720 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w3572_,
		_w3573_,
		_w6070_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4721 (
		_w3472_,
		_w3473_,
		_w3574_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h1)
	) name4722 (
		_w3637_,
		_w6071_,
		_w6072_
	);
	LUT4 #(
		.INIT('h0057)
	) name4723 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6068_,
		_w6069_,
		_w6072_,
		_w6073_
	);
	LUT2 #(
		.INIT('h2)
	) name4724 (
		_w3407_,
		_w6071_,
		_w6074_
	);
	LUT4 #(
		.INIT('hc055)
	) name4725 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3573_,
		_w6075_
	);
	LUT2 #(
		.INIT('h2)
	) name4726 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w3545_,
		_w6076_
	);
	LUT3 #(
		.INIT('h0d)
	) name4727 (
		_w2248_,
		_w6075_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h4)
	) name4728 (
		_w6074_,
		_w6077_,
		_w6078_
	);
	LUT3 #(
		.INIT('h2f)
	) name4729 (
		_w1939_,
		_w6073_,
		_w6078_,
		_w6079_
	);
	LUT4 #(
		.INIT('h6500)
	) name4730 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3572_,
		_w6080_
	);
	LUT4 #(
		.INIT('haa80)
	) name4731 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3611_,
		_w5940_,
		_w6080_,
		_w6081_
	);
	LUT3 #(
		.INIT('h02)
	) name4732 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w3580_,
		_w3573_,
		_w6082_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4733 (
		_w3450_,
		_w3451_,
		_w3653_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w3650_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h2)
	) name4735 (
		_w3407_,
		_w6083_,
		_w6085_
	);
	LUT4 #(
		.INIT('hc055)
	) name4736 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3580_,
		_w6086_
	);
	LUT2 #(
		.INIT('h2)
	) name4737 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		_w3545_,
		_w6087_
	);
	LUT3 #(
		.INIT('h0d)
	) name4738 (
		_w2248_,
		_w6086_,
		_w6087_,
		_w6088_
	);
	LUT2 #(
		.INIT('h4)
	) name4739 (
		_w6085_,
		_w6088_,
		_w6089_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4740 (
		_w1939_,
		_w6081_,
		_w6084_,
		_w6089_,
		_w6090_
	);
	LUT3 #(
		.INIT('h82)
	) name4741 (
		_w3611_,
		_w4503_,
		_w4506_,
		_w6091_
	);
	LUT2 #(
		.INIT('h8)
	) name4742 (
		_w3572_,
		_w5953_,
		_w6092_
	);
	LUT3 #(
		.INIT('h02)
	) name4743 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w3580_,
		_w3573_,
		_w6093_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4744 (
		_w3472_,
		_w3473_,
		_w3653_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name4745 (
		_w3650_,
		_w6094_,
		_w6095_
	);
	LUT4 #(
		.INIT('h0057)
	) name4746 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6091_,
		_w6092_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h2)
	) name4747 (
		_w3407_,
		_w6094_,
		_w6097_
	);
	LUT4 #(
		.INIT('hc055)
	) name4748 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3580_,
		_w6098_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		_w3545_,
		_w6099_
	);
	LUT3 #(
		.INIT('h0d)
	) name4750 (
		_w2248_,
		_w6098_,
		_w6099_,
		_w6100_
	);
	LUT2 #(
		.INIT('h4)
	) name4751 (
		_w6097_,
		_w6100_,
		_w6101_
	);
	LUT3 #(
		.INIT('h2f)
	) name4752 (
		_w1939_,
		_w6096_,
		_w6101_,
		_w6102_
	);
	LUT4 #(
		.INIT('h6500)
	) name4753 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3580_,
		_w6103_
	);
	LUT4 #(
		.INIT('haa80)
	) name4754 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3573_,
		_w5940_,
		_w6103_,
		_w6104_
	);
	LUT3 #(
		.INIT('h02)
	) name4755 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w3578_,
		_w3667_,
		_w6105_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4756 (
		_w3450_,
		_w3451_,
		_w3668_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name4757 (
		_w3664_,
		_w6106_,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name4758 (
		_w3407_,
		_w6106_,
		_w6108_
	);
	LUT4 #(
		.INIT('hc055)
	) name4759 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3667_,
		_w6109_
	);
	LUT2 #(
		.INIT('h2)
	) name4760 (
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w3545_,
		_w6110_
	);
	LUT3 #(
		.INIT('h0d)
	) name4761 (
		_w2248_,
		_w6109_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h4)
	) name4762 (
		_w6108_,
		_w6111_,
		_w6112_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4763 (
		_w1939_,
		_w6104_,
		_w6107_,
		_w6112_,
		_w6113_
	);
	LUT3 #(
		.INIT('h82)
	) name4764 (
		_w3573_,
		_w4503_,
		_w4506_,
		_w6114_
	);
	LUT2 #(
		.INIT('h8)
	) name4765 (
		_w3580_,
		_w5953_,
		_w6115_
	);
	LUT3 #(
		.INIT('h02)
	) name4766 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w3578_,
		_w3667_,
		_w6116_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4767 (
		_w3472_,
		_w3473_,
		_w3668_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h1)
	) name4768 (
		_w3664_,
		_w6117_,
		_w6118_
	);
	LUT4 #(
		.INIT('h0057)
	) name4769 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6114_,
		_w6115_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h2)
	) name4770 (
		_w3407_,
		_w6117_,
		_w6120_
	);
	LUT4 #(
		.INIT('hc055)
	) name4771 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3667_,
		_w6121_
	);
	LUT2 #(
		.INIT('h2)
	) name4772 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w3545_,
		_w6122_
	);
	LUT3 #(
		.INIT('h0d)
	) name4773 (
		_w2248_,
		_w6121_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name4774 (
		_w6120_,
		_w6123_,
		_w6124_
	);
	LUT3 #(
		.INIT('h2f)
	) name4775 (
		_w1939_,
		_w6119_,
		_w6124_,
		_w6125_
	);
	LUT4 #(
		.INIT('h6500)
	) name4776 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3578_,
		_w6126_
	);
	LUT4 #(
		.INIT('haa80)
	) name4777 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3580_,
		_w5940_,
		_w6126_,
		_w6127_
	);
	LUT3 #(
		.INIT('h02)
	) name4778 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w3667_,
		_w3683_,
		_w6128_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4779 (
		_w3450_,
		_w3451_,
		_w3698_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		_w3695_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('h2)
	) name4781 (
		_w3407_,
		_w6129_,
		_w6131_
	);
	LUT4 #(
		.INIT('hc055)
	) name4782 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3683_,
		_w6132_
	);
	LUT2 #(
		.INIT('h2)
	) name4783 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w3545_,
		_w6133_
	);
	LUT3 #(
		.INIT('h0d)
	) name4784 (
		_w2248_,
		_w6132_,
		_w6133_,
		_w6134_
	);
	LUT2 #(
		.INIT('h4)
	) name4785 (
		_w6131_,
		_w6134_,
		_w6135_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4786 (
		_w1939_,
		_w6127_,
		_w6130_,
		_w6135_,
		_w6136_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		_w3578_,
		_w5953_,
		_w6137_
	);
	LUT3 #(
		.INIT('h82)
	) name4788 (
		_w3580_,
		_w4503_,
		_w4506_,
		_w6138_
	);
	LUT3 #(
		.INIT('h02)
	) name4789 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w3667_,
		_w3683_,
		_w6139_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4790 (
		_w3472_,
		_w3473_,
		_w3698_,
		_w6139_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name4791 (
		_w3695_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h0057)
	) name4792 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6137_,
		_w6138_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h2)
	) name4793 (
		_w3407_,
		_w6140_,
		_w6143_
	);
	LUT4 #(
		.INIT('hc055)
	) name4794 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3683_,
		_w6144_
	);
	LUT2 #(
		.INIT('h2)
	) name4795 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w3545_,
		_w6145_
	);
	LUT3 #(
		.INIT('h0d)
	) name4796 (
		_w2248_,
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h4)
	) name4797 (
		_w6143_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h2f)
	) name4798 (
		_w1939_,
		_w6142_,
		_w6147_,
		_w6148_
	);
	LUT4 #(
		.INIT('h6500)
	) name4799 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3667_,
		_w6149_
	);
	LUT4 #(
		.INIT('haa80)
	) name4800 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3578_,
		_w5940_,
		_w6149_,
		_w6150_
	);
	LUT3 #(
		.INIT('h02)
	) name4801 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w3682_,
		_w3683_,
		_w6151_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4802 (
		_w3450_,
		_w3451_,
		_w3684_,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h1)
	) name4803 (
		_w3679_,
		_w6152_,
		_w6153_
	);
	LUT2 #(
		.INIT('h2)
	) name4804 (
		_w3407_,
		_w6152_,
		_w6154_
	);
	LUT4 #(
		.INIT('hc055)
	) name4805 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3682_,
		_w6155_
	);
	LUT2 #(
		.INIT('h2)
	) name4806 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w3545_,
		_w6156_
	);
	LUT3 #(
		.INIT('h0d)
	) name4807 (
		_w2248_,
		_w6155_,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h4)
	) name4808 (
		_w6154_,
		_w6157_,
		_w6158_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4809 (
		_w1939_,
		_w6150_,
		_w6153_,
		_w6158_,
		_w6159_
	);
	LUT3 #(
		.INIT('h82)
	) name4810 (
		_w3578_,
		_w4503_,
		_w4506_,
		_w6160_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		_w3667_,
		_w5953_,
		_w6161_
	);
	LUT3 #(
		.INIT('h02)
	) name4812 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w3682_,
		_w3683_,
		_w6162_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4813 (
		_w3472_,
		_w3473_,
		_w3684_,
		_w6162_,
		_w6163_
	);
	LUT2 #(
		.INIT('h1)
	) name4814 (
		_w3679_,
		_w6163_,
		_w6164_
	);
	LUT4 #(
		.INIT('h0057)
	) name4815 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6160_,
		_w6161_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h2)
	) name4816 (
		_w3407_,
		_w6163_,
		_w6166_
	);
	LUT4 #(
		.INIT('hc055)
	) name4817 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3682_,
		_w6167_
	);
	LUT2 #(
		.INIT('h2)
	) name4818 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w3545_,
		_w6168_
	);
	LUT3 #(
		.INIT('h0d)
	) name4819 (
		_w2248_,
		_w6167_,
		_w6168_,
		_w6169_
	);
	LUT2 #(
		.INIT('h4)
	) name4820 (
		_w6166_,
		_w6169_,
		_w6170_
	);
	LUT3 #(
		.INIT('h2f)
	) name4821 (
		_w1939_,
		_w6165_,
		_w6170_,
		_w6171_
	);
	LUT4 #(
		.INIT('h6500)
	) name4822 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3683_,
		_w6172_
	);
	LUT4 #(
		.INIT('haa80)
	) name4823 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3667_,
		_w5940_,
		_w6172_,
		_w6173_
	);
	LUT3 #(
		.INIT('h02)
	) name4824 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w3682_,
		_w3712_,
		_w6174_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4825 (
		_w3450_,
		_w3451_,
		_w3713_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h1)
	) name4826 (
		_w3709_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('h2)
	) name4827 (
		_w3407_,
		_w6175_,
		_w6177_
	);
	LUT4 #(
		.INIT('hc055)
	) name4828 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3712_,
		_w6178_
	);
	LUT2 #(
		.INIT('h2)
	) name4829 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w3545_,
		_w6179_
	);
	LUT3 #(
		.INIT('h0d)
	) name4830 (
		_w2248_,
		_w6178_,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('h4)
	) name4831 (
		_w6177_,
		_w6180_,
		_w6181_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4832 (
		_w1939_,
		_w6173_,
		_w6176_,
		_w6181_,
		_w6182_
	);
	LUT3 #(
		.INIT('h82)
	) name4833 (
		_w3667_,
		_w4503_,
		_w4506_,
		_w6183_
	);
	LUT2 #(
		.INIT('h8)
	) name4834 (
		_w3683_,
		_w5953_,
		_w6184_
	);
	LUT3 #(
		.INIT('h02)
	) name4835 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w3682_,
		_w3712_,
		_w6185_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4836 (
		_w3472_,
		_w3473_,
		_w3713_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w3709_,
		_w6186_,
		_w6187_
	);
	LUT4 #(
		.INIT('h0057)
	) name4838 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6183_,
		_w6184_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h2)
	) name4839 (
		_w3407_,
		_w6186_,
		_w6189_
	);
	LUT4 #(
		.INIT('hc055)
	) name4840 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3712_,
		_w6190_
	);
	LUT2 #(
		.INIT('h2)
	) name4841 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w3545_,
		_w6191_
	);
	LUT3 #(
		.INIT('h0d)
	) name4842 (
		_w2248_,
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h4)
	) name4843 (
		_w6189_,
		_w6192_,
		_w6193_
	);
	LUT3 #(
		.INIT('h2f)
	) name4844 (
		_w1939_,
		_w6188_,
		_w6193_,
		_w6194_
	);
	LUT4 #(
		.INIT('h6500)
	) name4845 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3682_,
		_w6195_
	);
	LUT4 #(
		.INIT('haa80)
	) name4846 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3683_,
		_w5940_,
		_w6195_,
		_w6196_
	);
	LUT3 #(
		.INIT('h02)
	) name4847 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w3712_,
		_w3727_,
		_w6197_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4848 (
		_w3450_,
		_w3451_,
		_w3728_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w3724_,
		_w6198_,
		_w6199_
	);
	LUT2 #(
		.INIT('h2)
	) name4850 (
		_w3407_,
		_w6198_,
		_w6200_
	);
	LUT4 #(
		.INIT('hc055)
	) name4851 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3727_,
		_w6201_
	);
	LUT2 #(
		.INIT('h2)
	) name4852 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w3545_,
		_w6202_
	);
	LUT3 #(
		.INIT('h0d)
	) name4853 (
		_w2248_,
		_w6201_,
		_w6202_,
		_w6203_
	);
	LUT2 #(
		.INIT('h4)
	) name4854 (
		_w6200_,
		_w6203_,
		_w6204_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4855 (
		_w1939_,
		_w6196_,
		_w6199_,
		_w6204_,
		_w6205_
	);
	LUT3 #(
		.INIT('h82)
	) name4856 (
		_w3683_,
		_w4503_,
		_w4506_,
		_w6206_
	);
	LUT2 #(
		.INIT('h8)
	) name4857 (
		_w3682_,
		_w5953_,
		_w6207_
	);
	LUT3 #(
		.INIT('h02)
	) name4858 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w3712_,
		_w3727_,
		_w6208_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4859 (
		_w3472_,
		_w3473_,
		_w3728_,
		_w6208_,
		_w6209_
	);
	LUT2 #(
		.INIT('h1)
	) name4860 (
		_w3724_,
		_w6209_,
		_w6210_
	);
	LUT4 #(
		.INIT('h0057)
	) name4861 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6206_,
		_w6207_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h2)
	) name4862 (
		_w3407_,
		_w6209_,
		_w6212_
	);
	LUT4 #(
		.INIT('hc055)
	) name4863 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3727_,
		_w6213_
	);
	LUT2 #(
		.INIT('h2)
	) name4864 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w3545_,
		_w6214_
	);
	LUT3 #(
		.INIT('h0d)
	) name4865 (
		_w2248_,
		_w6213_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h4)
	) name4866 (
		_w6212_,
		_w6215_,
		_w6216_
	);
	LUT3 #(
		.INIT('h2f)
	) name4867 (
		_w1939_,
		_w6211_,
		_w6216_,
		_w6217_
	);
	LUT4 #(
		.INIT('h6500)
	) name4868 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3712_,
		_w6218_
	);
	LUT4 #(
		.INIT('haa80)
	) name4869 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3682_,
		_w5940_,
		_w6218_,
		_w6219_
	);
	LUT3 #(
		.INIT('h02)
	) name4870 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w3727_,
		_w3742_,
		_w6220_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4871 (
		_w3450_,
		_w3451_,
		_w3743_,
		_w6220_,
		_w6221_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		_w3739_,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h2)
	) name4873 (
		_w3407_,
		_w6221_,
		_w6223_
	);
	LUT4 #(
		.INIT('hc055)
	) name4874 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3742_,
		_w6224_
	);
	LUT2 #(
		.INIT('h2)
	) name4875 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w3545_,
		_w6225_
	);
	LUT3 #(
		.INIT('h0d)
	) name4876 (
		_w2248_,
		_w6224_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h4)
	) name4877 (
		_w6223_,
		_w6226_,
		_w6227_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4878 (
		_w1939_,
		_w6219_,
		_w6222_,
		_w6227_,
		_w6228_
	);
	LUT3 #(
		.INIT('h82)
	) name4879 (
		_w3682_,
		_w4503_,
		_w4506_,
		_w6229_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		_w3712_,
		_w5953_,
		_w6230_
	);
	LUT3 #(
		.INIT('h02)
	) name4881 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w3727_,
		_w3742_,
		_w6231_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4882 (
		_w3472_,
		_w3473_,
		_w3743_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name4883 (
		_w3739_,
		_w6232_,
		_w6233_
	);
	LUT4 #(
		.INIT('h0057)
	) name4884 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6229_,
		_w6230_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name4885 (
		_w3407_,
		_w6232_,
		_w6235_
	);
	LUT4 #(
		.INIT('hc055)
	) name4886 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3742_,
		_w6236_
	);
	LUT2 #(
		.INIT('h2)
	) name4887 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w3545_,
		_w6237_
	);
	LUT3 #(
		.INIT('h0d)
	) name4888 (
		_w2248_,
		_w6236_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		_w6235_,
		_w6238_,
		_w6239_
	);
	LUT3 #(
		.INIT('h2f)
	) name4890 (
		_w1939_,
		_w6234_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h6500)
	) name4891 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3727_,
		_w6241_
	);
	LUT4 #(
		.INIT('haa80)
	) name4892 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3712_,
		_w5940_,
		_w6241_,
		_w6242_
	);
	LUT3 #(
		.INIT('h02)
	) name4893 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w3592_,
		_w3742_,
		_w6243_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4894 (
		_w3450_,
		_w3451_,
		_w3757_,
		_w6243_,
		_w6244_
	);
	LUT2 #(
		.INIT('h1)
	) name4895 (
		_w3754_,
		_w6244_,
		_w6245_
	);
	LUT2 #(
		.INIT('h2)
	) name4896 (
		_w3407_,
		_w6244_,
		_w6246_
	);
	LUT4 #(
		.INIT('hc055)
	) name4897 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3592_,
		_w6247_
	);
	LUT2 #(
		.INIT('h2)
	) name4898 (
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w3545_,
		_w6248_
	);
	LUT3 #(
		.INIT('h0d)
	) name4899 (
		_w2248_,
		_w6247_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h4)
	) name4900 (
		_w6246_,
		_w6249_,
		_w6250_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4901 (
		_w1939_,
		_w6242_,
		_w6245_,
		_w6250_,
		_w6251_
	);
	LUT3 #(
		.INIT('h82)
	) name4902 (
		_w3712_,
		_w4503_,
		_w4506_,
		_w6252_
	);
	LUT2 #(
		.INIT('h8)
	) name4903 (
		_w3727_,
		_w5953_,
		_w6253_
	);
	LUT3 #(
		.INIT('h02)
	) name4904 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w3592_,
		_w3742_,
		_w6254_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4905 (
		_w3472_,
		_w3473_,
		_w3757_,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h1)
	) name4906 (
		_w3754_,
		_w6255_,
		_w6256_
	);
	LUT4 #(
		.INIT('h0057)
	) name4907 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6252_,
		_w6253_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h2)
	) name4908 (
		_w3407_,
		_w6255_,
		_w6258_
	);
	LUT4 #(
		.INIT('hc055)
	) name4909 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3592_,
		_w6259_
	);
	LUT2 #(
		.INIT('h2)
	) name4910 (
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w3545_,
		_w6260_
	);
	LUT3 #(
		.INIT('h0d)
	) name4911 (
		_w2248_,
		_w6259_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h4)
	) name4912 (
		_w6258_,
		_w6261_,
		_w6262_
	);
	LUT3 #(
		.INIT('h2f)
	) name4913 (
		_w1939_,
		_w6257_,
		_w6262_,
		_w6263_
	);
	LUT4 #(
		.INIT('h6500)
	) name4914 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3742_,
		_w6264_
	);
	LUT4 #(
		.INIT('haa80)
	) name4915 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3727_,
		_w5940_,
		_w6264_,
		_w6265_
	);
	LUT3 #(
		.INIT('h02)
	) name4916 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w3411_,
		_w3592_,
		_w6266_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4917 (
		_w3450_,
		_w3451_,
		_w3593_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		_w3768_,
		_w6267_,
		_w6268_
	);
	LUT2 #(
		.INIT('h2)
	) name4919 (
		_w3407_,
		_w6267_,
		_w6269_
	);
	LUT4 #(
		.INIT('hc055)
	) name4920 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3411_,
		_w6270_
	);
	LUT2 #(
		.INIT('h2)
	) name4921 (
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w3545_,
		_w6271_
	);
	LUT3 #(
		.INIT('h0d)
	) name4922 (
		_w2248_,
		_w6270_,
		_w6271_,
		_w6272_
	);
	LUT2 #(
		.INIT('h4)
	) name4923 (
		_w6269_,
		_w6272_,
		_w6273_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4924 (
		_w1939_,
		_w6265_,
		_w6268_,
		_w6273_,
		_w6274_
	);
	LUT3 #(
		.INIT('h82)
	) name4925 (
		_w3727_,
		_w4503_,
		_w4506_,
		_w6275_
	);
	LUT2 #(
		.INIT('h8)
	) name4926 (
		_w3742_,
		_w5953_,
		_w6276_
	);
	LUT3 #(
		.INIT('h02)
	) name4927 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w3411_,
		_w3592_,
		_w6277_
	);
	LUT4 #(
		.INIT('h00f1)
	) name4928 (
		_w3472_,
		_w3473_,
		_w3593_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w3768_,
		_w6278_,
		_w6279_
	);
	LUT4 #(
		.INIT('h0057)
	) name4930 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6275_,
		_w6276_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h2)
	) name4931 (
		_w3407_,
		_w6278_,
		_w6281_
	);
	LUT4 #(
		.INIT('hc055)
	) name4932 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3411_,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name4933 (
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w3545_,
		_w6283_
	);
	LUT3 #(
		.INIT('h0d)
	) name4934 (
		_w2248_,
		_w6282_,
		_w6283_,
		_w6284_
	);
	LUT2 #(
		.INIT('h4)
	) name4935 (
		_w6281_,
		_w6284_,
		_w6285_
	);
	LUT3 #(
		.INIT('h2f)
	) name4936 (
		_w1939_,
		_w6280_,
		_w6285_,
		_w6286_
	);
	LUT4 #(
		.INIT('h6500)
	) name4937 (
		_w3510_,
		_w3496_,
		_w3532_,
		_w3592_,
		_w6287_
	);
	LUT4 #(
		.INIT('haa80)
	) name4938 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3742_,
		_w5940_,
		_w6287_,
		_w6288_
	);
	LUT3 #(
		.INIT('h02)
	) name4939 (
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w3411_,
		_w3412_,
		_w6289_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4940 (
		_w3413_,
		_w3450_,
		_w3451_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w3781_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h2)
	) name4942 (
		_w3407_,
		_w6290_,
		_w6292_
	);
	LUT4 #(
		.INIT('hc055)
	) name4943 (
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1787_,
		_w1792_,
		_w3412_,
		_w6293_
	);
	LUT2 #(
		.INIT('h2)
	) name4944 (
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w3545_,
		_w6294_
	);
	LUT3 #(
		.INIT('h0d)
	) name4945 (
		_w2248_,
		_w6293_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h4)
	) name4946 (
		_w6292_,
		_w6295_,
		_w6296_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4947 (
		_w1939_,
		_w6288_,
		_w6291_,
		_w6296_,
		_w6297_
	);
	LUT3 #(
		.INIT('h82)
	) name4948 (
		_w3742_,
		_w4503_,
		_w4506_,
		_w6298_
	);
	LUT2 #(
		.INIT('h8)
	) name4949 (
		_w3592_,
		_w5953_,
		_w6299_
	);
	LUT3 #(
		.INIT('h02)
	) name4950 (
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w3411_,
		_w3412_,
		_w6300_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4951 (
		_w3413_,
		_w3472_,
		_w3473_,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w3781_,
		_w6301_,
		_w6302_
	);
	LUT4 #(
		.INIT('h0057)
	) name4953 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6298_,
		_w6299_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h2)
	) name4954 (
		_w3407_,
		_w6301_,
		_w6304_
	);
	LUT4 #(
		.INIT('hc055)
	) name4955 (
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1755_,
		_w1760_,
		_w3412_,
		_w6305_
	);
	LUT2 #(
		.INIT('h2)
	) name4956 (
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w3545_,
		_w6306_
	);
	LUT3 #(
		.INIT('h0d)
	) name4957 (
		_w2248_,
		_w6305_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h4)
	) name4958 (
		_w6304_,
		_w6307_,
		_w6308_
	);
	LUT3 #(
		.INIT('h2f)
	) name4959 (
		_w1939_,
		_w6303_,
		_w6308_,
		_w6309_
	);
	LUT3 #(
		.INIT('h08)
	) name4960 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w1592_,
		_w1660_,
		_w6310_
	);
	LUT4 #(
		.INIT('h0400)
	) name4961 (
		_w4360_,
		_w4906_,
		_w5699_,
		_w5698_,
		_w6311_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name4962 (
		_w4360_,
		_w4906_,
		_w5699_,
		_w5698_,
		_w6312_
	);
	LUT3 #(
		.INIT('h01)
	) name4963 (
		_w4214_,
		_w6312_,
		_w6311_,
		_w6313_
	);
	LUT3 #(
		.INIT('h6c)
	) name4964 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4277_,
		_w6314_
	);
	LUT2 #(
		.INIT('h8)
	) name4965 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4265_,
		_w6315_
	);
	LUT3 #(
		.INIT('h80)
	) name4966 (
		_w4271_,
		_w4275_,
		_w6315_,
		_w6316_
	);
	LUT4 #(
		.INIT('h820a)
	) name4967 (
		_w4214_,
		_w4862_,
		_w6314_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h1)
	) name4968 (
		_w1661_,
		_w6317_,
		_w6318_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4969 (
		_w1559_,
		_w6310_,
		_w6313_,
		_w6318_,
		_w6319_
	);
	LUT4 #(
		.INIT('h028a)
	) name4970 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w6320_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4971 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w4425_,
		_w6321_
	);
	LUT2 #(
		.INIT('h8)
	) name4972 (
		\P2_InstAddrPointer_reg[29]/NET0131 ,
		_w4427_,
		_w6322_
	);
	LUT3 #(
		.INIT('h13)
	) name4973 (
		_w4916_,
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT3 #(
		.INIT('h2a)
	) name4974 (
		_w1659_,
		_w4916_,
		_w5717_,
		_w6324_
	);
	LUT3 #(
		.INIT('h45)
	) name4975 (
		_w6320_,
		_w6323_,
		_w6324_,
		_w6325_
	);
	LUT3 #(
		.INIT('h48)
	) name4976 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w2242_,
		_w5739_,
		_w6326_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4977 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		_w5743_,
		_w6327_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4978 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2286_,
		_w5747_,
		_w6328_
	);
	LUT3 #(
		.INIT('h70)
	) name4979 (
		_w5746_,
		_w6327_,
		_w6328_,
		_w6329_
	);
	LUT2 #(
		.INIT('h4)
	) name4980 (
		_w6326_,
		_w6329_,
		_w6330_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4981 (
		_w1678_,
		_w6319_,
		_w6325_,
		_w6330_,
		_w6331_
	);
	LUT3 #(
		.INIT('h02)
	) name4982 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6332_
	);
	LUT3 #(
		.INIT('h80)
	) name4983 (
		_w2965_,
		_w2970_,
		_w4773_,
		_w6333_
	);
	LUT2 #(
		.INIT('h8)
	) name4984 (
		_w5385_,
		_w6333_,
		_w6334_
	);
	LUT4 #(
		.INIT('h8000)
	) name4985 (
		\P3_InstAddrPointer_reg[28]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2969_,
		_w2975_,
		_w6335_
	);
	LUT4 #(
		.INIT('h8000)
	) name4986 (
		_w2978_,
		_w4772_,
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT4 #(
		.INIT('h1555)
	) name4987 (
		_w2978_,
		_w4772_,
		_w6334_,
		_w6335_,
		_w6337_
	);
	LUT3 #(
		.INIT('h02)
	) name4988 (
		_w2755_,
		_w6337_,
		_w6336_,
		_w6338_
	);
	LUT3 #(
		.INIT('h80)
	) name4989 (
		_w2910_,
		_w4776_,
		_w4778_,
		_w6339_
	);
	LUT3 #(
		.INIT('h80)
	) name4990 (
		_w4074_,
		_w4777_,
		_w6339_,
		_w6340_
	);
	LUT4 #(
		.INIT('h4000)
	) name4991 (
		_w2911_,
		_w4074_,
		_w4777_,
		_w6339_,
		_w6341_
	);
	LUT4 #(
		.INIT('h4105)
	) name4992 (
		_w2755_,
		_w2732_,
		_w2743_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w2173_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4994 (
		_w2171_,
		_w6332_,
		_w6338_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4995 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w6345_
	);
	LUT4 #(
		.INIT('h2888)
	) name4996 (
		_w2181_,
		_w3041_,
		_w3044_,
		_w4090_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w6345_,
		_w6346_,
		_w6347_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name4998 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w5756_,
		_w5775_,
		_w6348_
	);
	LUT4 #(
		.INIT('hffeb)
	) name4999 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w6349_
	);
	LUT3 #(
		.INIT('h0d)
	) name5000 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w3055_,
		_w6349_,
		_w6350_
	);
	LUT4 #(
		.INIT('h4888)
	) name5001 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		_w2199_,
		_w5756_,
		_w5777_,
		_w6351_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5002 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w3054_,
		_w5783_,
		_w6352_
	);
	LUT4 #(
		.INIT('h1500)
	) name5003 (
		_w6351_,
		_w6348_,
		_w6350_,
		_w6352_,
		_w6353_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5004 (
		_w1945_,
		_w6344_,
		_w6347_,
		_w6353_,
		_w6354_
	);
	LUT3 #(
		.INIT('h08)
	) name5005 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w1842_,
		_w1915_,
		_w6355_
	);
	LUT4 #(
		.INIT('haa20)
	) name5006 (
		_w1810_,
		_w3266_,
		_w3324_,
		_w6355_,
		_w6356_
	);
	LUT3 #(
		.INIT('he4)
	) name5007 (
		_w1809_,
		_w1810_,
		_w1846_,
		_w6357_
	);
	LUT4 #(
		.INIT('h028a)
	) name5008 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w6358_
	);
	LUT4 #(
		.INIT('h000b)
	) name5009 (
		_w3391_,
		_w3393_,
		_w6356_,
		_w6358_,
		_w6359_
	);
	LUT3 #(
		.INIT('h80)
	) name5010 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w6360_
	);
	LUT2 #(
		.INIT('h8)
	) name5011 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6361_
	);
	LUT4 #(
		.INIT('h8000)
	) name5012 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w6362_
	);
	LUT4 #(
		.INIT('h8000)
	) name5013 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w6363_
	);
	LUT3 #(
		.INIT('h80)
	) name5014 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w6364_
	);
	LUT4 #(
		.INIT('h8000)
	) name5015 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w6365_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w6365_,
		_w6366_
	);
	LUT4 #(
		.INIT('h8000)
	) name5017 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w6365_,
		_w6367_
	);
	LUT4 #(
		.INIT('h8000)
	) name5018 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w6367_,
		_w6368_
	);
	LUT3 #(
		.INIT('h80)
	) name5019 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w6368_,
		_w6369_
	);
	LUT4 #(
		.INIT('h8000)
	) name5020 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w6368_,
		_w6370_
	);
	LUT3 #(
		.INIT('h80)
	) name5021 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w6370_,
		_w6371_
	);
	LUT4 #(
		.INIT('h8000)
	) name5022 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w6370_,
		_w6372_
	);
	LUT3 #(
		.INIT('h80)
	) name5023 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6363_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('h8000)
	) name5024 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6363_,
		_w6362_,
		_w6372_,
		_w6374_
	);
	LUT3 #(
		.INIT('h80)
	) name5025 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6360_,
		_w6374_,
		_w6375_
	);
	LUT4 #(
		.INIT('h8000)
	) name5026 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w6360_,
		_w6374_,
		_w6376_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name5027 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w6360_,
		_w6374_,
		_w6377_
	);
	LUT3 #(
		.INIT('h0d)
	) name5028 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w4953_,
		_w6378_
	);
	LUT4 #(
		.INIT('h8000)
	) name5029 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6370_,
		_w6379_
	);
	LUT4 #(
		.INIT('h8000)
	) name5030 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6379_,
		_w6363_,
		_w6362_,
		_w6380_
	);
	LUT3 #(
		.INIT('h80)
	) name5031 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w6380_,
		_w6360_,
		_w6381_
	);
	LUT4 #(
		.INIT('h4888)
	) name5032 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		_w2310_,
		_w6380_,
		_w6360_,
		_w6382_
	);
	LUT4 #(
		.INIT('hfc35)
	) name5033 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w6383_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5034 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w3406_,
		_w6383_,
		_w6384_
	);
	LUT4 #(
		.INIT('h1500)
	) name5035 (
		_w6382_,
		_w6377_,
		_w6378_,
		_w6384_,
		_w6385_
	);
	LUT3 #(
		.INIT('h2f)
	) name5036 (
		_w1933_,
		_w6359_,
		_w6385_,
		_w6386_
	);
	LUT3 #(
		.INIT('h02)
	) name5037 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6387_
	);
	LUT4 #(
		.INIT('h280a)
	) name5038 (
		_w2755_,
		_w2935_,
		_w2936_,
		_w2940_,
		_w6388_
	);
	LUT4 #(
		.INIT('hf040)
	) name5039 (
		_w2831_,
		_w2858_,
		_w2863_,
		_w5816_,
		_w6389_
	);
	LUT4 #(
		.INIT('h5554)
	) name5040 (
		_w2173_,
		_w5818_,
		_w6389_,
		_w6388_,
		_w6390_
	);
	LUT3 #(
		.INIT('ha8)
	) name5041 (
		_w2171_,
		_w6387_,
		_w6390_,
		_w6391_
	);
	LUT3 #(
		.INIT('h87)
	) name5042 (
		_w2749_,
		_w2754_,
		_w2992_,
		_w6392_
	);
	LUT4 #(
		.INIT('h4500)
	) name5043 (
		_w2995_,
		_w3014_,
		_w3017_,
		_w6392_,
		_w6393_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5044 (
		_w2995_,
		_w3014_,
		_w3017_,
		_w6392_,
		_w6394_
	);
	LUT3 #(
		.INIT('h02)
	) name5045 (
		_w2181_,
		_w6394_,
		_w6393_,
		_w6395_
	);
	LUT4 #(
		.INIT('he000)
	) name5046 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2992_,
		_w6396_
	);
	LUT4 #(
		.INIT('h004f)
	) name5047 (
		_w2073_,
		_w2086_,
		_w2757_,
		_w6396_,
		_w6397_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5048 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w6398_
	);
	LUT2 #(
		.INIT('h4)
	) name5049 (
		_w2117_,
		_w2936_,
		_w6399_
	);
	LUT4 #(
		.INIT('h0100)
	) name5050 (
		_w6398_,
		_w6399_,
		_w6395_,
		_w6397_,
		_w6400_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5051 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w3054_,
		_w3056_,
		_w6401_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5052 (
		_w1945_,
		_w6391_,
		_w6400_,
		_w6401_,
		_w6402_
	);
	LUT3 #(
		.INIT('h02)
	) name5053 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6403_
	);
	LUT2 #(
		.INIT('h8)
	) name5054 (
		_w4066_,
		_w4074_,
		_w6404_
	);
	LUT4 #(
		.INIT('hef00)
	) name5055 (
		_w2758_,
		_w2831_,
		_w2858_,
		_w2866_,
		_w6405_
	);
	LUT3 #(
		.INIT('h51)
	) name5056 (
		_w2755_,
		_w2871_,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h4)
	) name5057 (
		_w6404_,
		_w6406_,
		_w6407_
	);
	LUT4 #(
		.INIT('h004f)
	) name5058 (
		_w2935_,
		_w2941_,
		_w5353_,
		_w5354_,
		_w6408_
	);
	LUT4 #(
		.INIT('h00f7)
	) name5059 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2944_,
		_w4051_,
		_w6408_,
		_w6409_
	);
	LUT3 #(
		.INIT('h51)
	) name5060 (
		_w2173_,
		_w2755_,
		_w6409_,
		_w6410_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5061 (
		_w2171_,
		_w6403_,
		_w6407_,
		_w6410_,
		_w6411_
	);
	LUT4 #(
		.INIT('h8880)
	) name5062 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2988_,
		_w2993_,
		_w3020_,
		_w6412_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5063 (
		\P3_InstAddrPointer_reg[7]/NET0131 ,
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2985_,
		_w6413_
	);
	LUT4 #(
		.INIT('h0057)
	) name5064 (
		_w2988_,
		_w2993_,
		_w3020_,
		_w6413_,
		_w6414_
	);
	LUT3 #(
		.INIT('h02)
	) name5065 (
		_w2181_,
		_w6414_,
		_w6412_,
		_w6415_
	);
	LUT4 #(
		.INIT('h0903)
	) name5066 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2116_,
		_w2715_,
		_w6416_
	);
	LUT4 #(
		.INIT('h00e4)
	) name5067 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w6416_,
		_w6417_
	);
	LUT4 #(
		.INIT('h000e)
	) name5068 (
		_w2112_,
		_w2137_,
		_w2175_,
		_w6417_,
		_w6418_
	);
	LUT2 #(
		.INIT('h2)
	) name5069 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w6418_,
		_w6419_
	);
	LUT3 #(
		.INIT('hb0)
	) name5070 (
		_w2073_,
		_w2086_,
		_w2871_,
		_w6420_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name5071 (
		\P3_InstAddrPointer_reg[8]/NET0131 ,
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2116_,
		_w2715_,
		_w6421_
	);
	LUT3 #(
		.INIT('he0)
	) name5072 (
		_w2108_,
		_w2115_,
		_w6421_,
		_w6422_
	);
	LUT2 #(
		.INIT('h8)
	) name5073 (
		_w2064_,
		_w5354_,
		_w6423_
	);
	LUT3 #(
		.INIT('he2)
	) name5074 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2098_,
		_w6413_,
		_w6424_
	);
	LUT4 #(
		.INIT('h010f)
	) name5075 (
		_w2071_,
		_w2087_,
		_w6423_,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('h4)
	) name5076 (
		_w6422_,
		_w6425_,
		_w6426_
	);
	LUT3 #(
		.INIT('h10)
	) name5077 (
		_w6419_,
		_w6420_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h4)
	) name5078 (
		_w6415_,
		_w6427_,
		_w6428_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5079 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w3054_,
		_w3056_,
		_w6429_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5080 (
		_w1945_,
		_w6411_,
		_w6428_,
		_w6429_,
		_w6430_
	);
	LUT4 #(
		.INIT('h4414)
	) name5081 (
		_w4214_,
		_w4283_,
		_w4311_,
		_w4824_,
		_w6431_
	);
	LUT4 #(
		.INIT('h2822)
	) name5082 (
		_w4214_,
		_w4216_,
		_w4201_,
		_w4220_,
		_w6432_
	);
	LUT4 #(
		.INIT('h4447)
	) name5083 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w1661_,
		_w6431_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		_w1559_,
		_w6433_,
		_w6434_
	);
	LUT4 #(
		.INIT('h40bf)
	) name5085 (
		_w4208_,
		_w4206_,
		_w4213_,
		_w4375_,
		_w6435_
	);
	LUT4 #(
		.INIT('h2f00)
	) name5086 (
		_w4381_,
		_w4395_,
		_w4398_,
		_w6435_,
		_w6436_
	);
	LUT4 #(
		.INIT('h00d0)
	) name5087 (
		_w4381_,
		_w4395_,
		_w4398_,
		_w6435_,
		_w6437_
	);
	LUT3 #(
		.INIT('h02)
	) name5088 (
		_w1659_,
		_w6437_,
		_w6436_,
		_w6438_
	);
	LUT2 #(
		.INIT('h2)
	) name5089 (
		_w1565_,
		_w1602_,
		_w6439_
	);
	LUT4 #(
		.INIT('h5f13)
	) name5090 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1602_,
		_w6440_
	);
	LUT2 #(
		.INIT('h1)
	) name5091 (
		_w4185_,
		_w6440_,
		_w6441_
	);
	LUT3 #(
		.INIT('hc4)
	) name5092 (
		_w1617_,
		_w4216_,
		_w6441_,
		_w6442_
	);
	LUT3 #(
		.INIT('h01)
	) name5093 (
		_w1592_,
		_w1595_,
		_w4375_,
		_w6443_
	);
	LUT4 #(
		.INIT('h00c8)
	) name5094 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w6443_,
		_w6444_
	);
	LUT4 #(
		.INIT('h0203)
	) name5095 (
		_w1501_,
		_w1565_,
		_w1566_,
		_w1568_,
		_w6445_
	);
	LUT2 #(
		.INIT('h2)
	) name5096 (
		_w1602_,
		_w6445_,
		_w6446_
	);
	LUT3 #(
		.INIT('h32)
	) name5097 (
		_w1606_,
		_w1667_,
		_w6440_,
		_w6447_
	);
	LUT4 #(
		.INIT('h0100)
	) name5098 (
		_w1657_,
		_w6444_,
		_w6446_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h8)
	) name5099 (
		_w1596_,
		_w6444_,
		_w6449_
	);
	LUT4 #(
		.INIT('h004f)
	) name5100 (
		_w1571_,
		_w1583_,
		_w4283_,
		_w6449_,
		_w6450_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5101 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		_w6448_,
		_w6442_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5102 (
		_w1678_,
		_w6434_,
		_w6438_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5103 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w2286_,
		_w4441_,
		_w6453_
	);
	LUT2 #(
		.INIT('hb)
	) name5104 (
		_w6452_,
		_w6453_,
		_w6454_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5105 (
		_w4201_,
		_w4221_,
		_w4224_,
		_w4228_,
		_w6455_
	);
	LUT4 #(
		.INIT('h00b0)
	) name5106 (
		_w4201_,
		_w4221_,
		_w4224_,
		_w4228_,
		_w6456_
	);
	LUT3 #(
		.INIT('h02)
	) name5107 (
		_w4214_,
		_w6456_,
		_w6455_,
		_w6457_
	);
	LUT4 #(
		.INIT('h1055)
	) name5108 (
		_w4214_,
		_w4308_,
		_w4317_,
		_w4321_,
		_w6458_
	);
	LUT4 #(
		.INIT('hef00)
	) name5109 (
		_w4315_,
		_w4321_,
		_w4818_,
		_w6458_,
		_w6459_
	);
	LUT4 #(
		.INIT('h7774)
	) name5110 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1661_,
		_w6459_,
		_w6457_,
		_w6460_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5111 (
		\P2_InstAddrPointer_reg[7]/NET0131 ,
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w4374_,
		_w6461_
	);
	LUT3 #(
		.INIT('h0b)
	) name5112 (
		_w4400_,
		_w4404_,
		_w6461_,
		_w6462_
	);
	LUT3 #(
		.INIT('h8a)
	) name5113 (
		_w1659_,
		_w4400_,
		_w4405_,
		_w6463_
	);
	LUT3 #(
		.INIT('hb0)
	) name5114 (
		_w1571_,
		_w1583_,
		_w4321_,
		_w6464_
	);
	LUT3 #(
		.INIT('h47)
	) name5115 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1605_,
		_w4228_,
		_w6465_
	);
	LUT4 #(
		.INIT('h00ec)
	) name5116 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w6465_,
		_w6466_
	);
	LUT4 #(
		.INIT('h5457)
	) name5117 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1605_,
		_w1611_,
		_w4228_,
		_w6467_
	);
	LUT4 #(
		.INIT('h00dc)
	) name5118 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w6467_,
		_w6468_
	);
	LUT3 #(
		.INIT('h54)
	) name5119 (
		_w1602_,
		_w6466_,
		_w6468_,
		_w6469_
	);
	LUT3 #(
		.INIT('ha8)
	) name5120 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1626_,
		_w1667_,
		_w6470_
	);
	LUT2 #(
		.INIT('h8)
	) name5121 (
		_w1563_,
		_w4228_,
		_w6471_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5122 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		_w1592_,
		_w1595_,
		_w4402_,
		_w6472_
	);
	LUT4 #(
		.INIT('hc800)
	) name5123 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h1)
	) name5124 (
		_w6471_,
		_w6473_,
		_w6474_
	);
	LUT3 #(
		.INIT('h10)
	) name5125 (
		_w6470_,
		_w6469_,
		_w6474_,
		_w6475_
	);
	LUT4 #(
		.INIT('h0b00)
	) name5126 (
		_w6462_,
		_w6463_,
		_w6464_,
		_w6475_,
		_w6476_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5127 (
		_w1559_,
		_w1678_,
		_w6460_,
		_w6476_,
		_w6477_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5128 (
		\P2_InstAddrPointer_reg[9]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w2286_,
		_w4441_,
		_w6478_
	);
	LUT2 #(
		.INIT('hb)
	) name5129 (
		_w6477_,
		_w6478_,
		_w6479_
	);
	LUT3 #(
		.INIT('h02)
	) name5130 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w3534_,
		_w3536_,
		_w6480_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5131 (
		_w3537_,
		_w3479_,
		_w3480_,
		_w6480_,
		_w6481_
	);
	LUT3 #(
		.INIT('h32)
	) name5132 (
		_w4953_,
		_w4956_,
		_w6481_,
		_w6482_
	);
	LUT4 #(
		.INIT('h02fd)
	) name5133 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3522_,
		_w6483_
	);
	LUT3 #(
		.INIT('h65)
	) name5134 (
		_w3489_,
		_w3493_,
		_w3531_,
		_w6484_
	);
	LUT3 #(
		.INIT('hc4)
	) name5135 (
		_w3407_,
		_w3414_,
		_w6481_,
		_w6485_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5136 (
		_w3411_,
		_w6484_,
		_w6483_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h2)
	) name5137 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w3545_,
		_w6487_
	);
	LUT4 #(
		.INIT('hc055)
	) name5138 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3534_,
		_w6488_
	);
	LUT3 #(
		.INIT('h31)
	) name5139 (
		_w2248_,
		_w6487_,
		_w6488_,
		_w6489_
	);
	LUT3 #(
		.INIT('h1f)
	) name5140 (
		_w6482_,
		_w6486_,
		_w6489_,
		_w6490_
	);
	LUT4 #(
		.INIT('hc444)
	) name5141 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6491_
	);
	LUT4 #(
		.INIT('h0888)
	) name5142 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[29]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6492_
	);
	LUT2 #(
		.INIT('h1)
	) name5143 (
		_w6491_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('ha8)
	) name5144 (
		_w2250_,
		_w6491_,
		_w6492_,
		_w6494_
	);
	LUT4 #(
		.INIT('hc444)
	) name5145 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[21]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6495_
	);
	LUT4 #(
		.INIT('h0888)
	) name5146 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[21]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6496_
	);
	LUT2 #(
		.INIT('h1)
	) name5147 (
		_w6495_,
		_w6496_,
		_w6497_
	);
	LUT3 #(
		.INIT('ha8)
	) name5148 (
		_w2264_,
		_w6495_,
		_w6496_,
		_w6498_
	);
	LUT3 #(
		.INIT('ha8)
	) name5149 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6494_,
		_w6498_,
		_w6499_
	);
	LUT4 #(
		.INIT('hc444)
	) name5150 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6500_
	);
	LUT4 #(
		.INIT('h0888)
	) name5151 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[5]/NET0131 ,
		_w2255_,
		_w2260_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		_w6500_,
		_w6501_,
		_w6502_
	);
	LUT3 #(
		.INIT('h02)
	) name5153 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w2271_,
		_w2272_,
		_w6503_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5154 (
		_w2273_,
		_w6500_,
		_w6501_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name5155 (
		_w2280_,
		_w6504_,
		_w6505_
	);
	LUT3 #(
		.INIT('ha8)
	) name5156 (
		_w1679_,
		_w6499_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h2)
	) name5157 (
		_w2283_,
		_w6504_,
		_w6507_
	);
	LUT4 #(
		.INIT('hc055)
	) name5158 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2272_,
		_w6508_
	);
	LUT2 #(
		.INIT('h2)
	) name5159 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		_w2288_,
		_w6509_
	);
	LUT3 #(
		.INIT('h0d)
	) name5160 (
		_w2246_,
		_w6508_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h4)
	) name5161 (
		_w6507_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('hb)
	) name5162 (
		_w6506_,
		_w6511_,
		_w6512_
	);
	LUT3 #(
		.INIT('h02)
	) name5163 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w3578_,
		_w3580_,
		_w6513_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5164 (
		_w3479_,
		_w3480_,
		_w3581_,
		_w6513_,
		_w6514_
	);
	LUT3 #(
		.INIT('h32)
	) name5165 (
		_w4953_,
		_w4990_,
		_w6514_,
		_w6515_
	);
	LUT3 #(
		.INIT('hc4)
	) name5166 (
		_w3407_,
		_w3575_,
		_w6514_,
		_w6516_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5167 (
		_w3572_,
		_w6484_,
		_w6483_,
		_w6516_,
		_w6517_
	);
	LUT2 #(
		.INIT('h2)
	) name5168 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w3545_,
		_w6518_
	);
	LUT4 #(
		.INIT('hc055)
	) name5169 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3578_,
		_w6519_
	);
	LUT3 #(
		.INIT('h31)
	) name5170 (
		_w2248_,
		_w6518_,
		_w6519_,
		_w6520_
	);
	LUT3 #(
		.INIT('h1f)
	) name5171 (
		_w6515_,
		_w6517_,
		_w6520_,
		_w6521_
	);
	LUT3 #(
		.INIT('h02)
	) name5172 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		_w3536_,
		_w3412_,
		_w6522_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5173 (
		_w3479_,
		_w3480_,
		_w3597_,
		_w6522_,
		_w6523_
	);
	LUT3 #(
		.INIT('h32)
	) name5174 (
		_w4953_,
		_w5001_,
		_w6523_,
		_w6524_
	);
	LUT3 #(
		.INIT('hc4)
	) name5175 (
		_w3407_,
		_w3594_,
		_w6523_,
		_w6525_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5176 (
		_w3592_,
		_w6484_,
		_w6483_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h2)
	) name5177 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		_w3545_,
		_w6527_
	);
	LUT4 #(
		.INIT('hc055)
	) name5178 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3536_,
		_w6528_
	);
	LUT3 #(
		.INIT('h31)
	) name5179 (
		_w2248_,
		_w6527_,
		_w6528_,
		_w6529_
	);
	LUT3 #(
		.INIT('h1f)
	) name5180 (
		_w6524_,
		_w6526_,
		_w6529_,
		_w6530_
	);
	LUT3 #(
		.INIT('h02)
	) name5181 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w3534_,
		_w3611_,
		_w6531_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5182 (
		_w3479_,
		_w3480_,
		_w3612_,
		_w6531_,
		_w6532_
	);
	LUT3 #(
		.INIT('h32)
	) name5183 (
		_w4953_,
		_w5012_,
		_w6532_,
		_w6533_
	);
	LUT3 #(
		.INIT('hc4)
	) name5184 (
		_w3407_,
		_w3608_,
		_w6532_,
		_w6534_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5185 (
		_w3412_,
		_w6484_,
		_w6483_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h2)
	) name5186 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w3545_,
		_w6536_
	);
	LUT4 #(
		.INIT('hc055)
	) name5187 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3611_,
		_w6537_
	);
	LUT3 #(
		.INIT('h31)
	) name5188 (
		_w2248_,
		_w6536_,
		_w6537_,
		_w6538_
	);
	LUT3 #(
		.INIT('h1f)
	) name5189 (
		_w6533_,
		_w6535_,
		_w6538_,
		_w6539_
	);
	LUT3 #(
		.INIT('h02)
	) name5190 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w3572_,
		_w3611_,
		_w6540_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5191 (
		_w3479_,
		_w3480_,
		_w3626_,
		_w6540_,
		_w6541_
	);
	LUT3 #(
		.INIT('h32)
	) name5192 (
		_w4953_,
		_w5023_,
		_w6541_,
		_w6542_
	);
	LUT3 #(
		.INIT('hc4)
	) name5193 (
		_w3407_,
		_w3623_,
		_w6541_,
		_w6543_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5194 (
		_w3536_,
		_w6484_,
		_w6483_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h2)
	) name5195 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w3545_,
		_w6545_
	);
	LUT4 #(
		.INIT('hc055)
	) name5196 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3572_,
		_w6546_
	);
	LUT3 #(
		.INIT('h31)
	) name5197 (
		_w2248_,
		_w6545_,
		_w6546_,
		_w6547_
	);
	LUT3 #(
		.INIT('h1f)
	) name5198 (
		_w6542_,
		_w6544_,
		_w6547_,
		_w6548_
	);
	LUT3 #(
		.INIT('h02)
	) name5199 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w3572_,
		_w3573_,
		_w6549_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5200 (
		_w3479_,
		_w3480_,
		_w3574_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h32)
	) name5201 (
		_w4953_,
		_w5034_,
		_w6550_,
		_w6551_
	);
	LUT3 #(
		.INIT('hc4)
	) name5202 (
		_w3407_,
		_w3637_,
		_w6550_,
		_w6552_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5203 (
		_w3534_,
		_w6484_,
		_w6483_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h2)
	) name5204 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w3545_,
		_w6554_
	);
	LUT4 #(
		.INIT('hc055)
	) name5205 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3573_,
		_w6555_
	);
	LUT3 #(
		.INIT('h31)
	) name5206 (
		_w2248_,
		_w6554_,
		_w6555_,
		_w6556_
	);
	LUT3 #(
		.INIT('h1f)
	) name5207 (
		_w6551_,
		_w6553_,
		_w6556_,
		_w6557_
	);
	LUT3 #(
		.INIT('h02)
	) name5208 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w3580_,
		_w3573_,
		_w6558_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5209 (
		_w3479_,
		_w3480_,
		_w3653_,
		_w6558_,
		_w6559_
	);
	LUT3 #(
		.INIT('h32)
	) name5210 (
		_w4953_,
		_w5045_,
		_w6559_,
		_w6560_
	);
	LUT3 #(
		.INIT('hc4)
	) name5211 (
		_w3407_,
		_w3650_,
		_w6559_,
		_w6561_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5212 (
		_w3611_,
		_w6484_,
		_w6483_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h2)
	) name5213 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w3545_,
		_w6563_
	);
	LUT4 #(
		.INIT('hc055)
	) name5214 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3580_,
		_w6564_
	);
	LUT3 #(
		.INIT('h31)
	) name5215 (
		_w2248_,
		_w6563_,
		_w6564_,
		_w6565_
	);
	LUT3 #(
		.INIT('h1f)
	) name5216 (
		_w6560_,
		_w6562_,
		_w6565_,
		_w6566_
	);
	LUT3 #(
		.INIT('h02)
	) name5217 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w3578_,
		_w3667_,
		_w6567_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5218 (
		_w3479_,
		_w3480_,
		_w3668_,
		_w6567_,
		_w6568_
	);
	LUT3 #(
		.INIT('h32)
	) name5219 (
		_w4953_,
		_w5056_,
		_w6568_,
		_w6569_
	);
	LUT3 #(
		.INIT('hc4)
	) name5220 (
		_w3407_,
		_w3664_,
		_w6568_,
		_w6570_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5221 (
		_w3573_,
		_w6484_,
		_w6483_,
		_w6570_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name5222 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w3545_,
		_w6572_
	);
	LUT4 #(
		.INIT('hc055)
	) name5223 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3667_,
		_w6573_
	);
	LUT3 #(
		.INIT('h31)
	) name5224 (
		_w2248_,
		_w6572_,
		_w6573_,
		_w6574_
	);
	LUT3 #(
		.INIT('h1f)
	) name5225 (
		_w6569_,
		_w6571_,
		_w6574_,
		_w6575_
	);
	LUT3 #(
		.INIT('h02)
	) name5226 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w3667_,
		_w3683_,
		_w6576_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5227 (
		_w3479_,
		_w3480_,
		_w3698_,
		_w6576_,
		_w6577_
	);
	LUT3 #(
		.INIT('h32)
	) name5228 (
		_w4953_,
		_w5067_,
		_w6577_,
		_w6578_
	);
	LUT3 #(
		.INIT('hc4)
	) name5229 (
		_w3407_,
		_w3695_,
		_w6577_,
		_w6579_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5230 (
		_w3580_,
		_w6484_,
		_w6483_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h2)
	) name5231 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w3545_,
		_w6581_
	);
	LUT4 #(
		.INIT('hc055)
	) name5232 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3683_,
		_w6582_
	);
	LUT3 #(
		.INIT('h31)
	) name5233 (
		_w2248_,
		_w6581_,
		_w6582_,
		_w6583_
	);
	LUT3 #(
		.INIT('h1f)
	) name5234 (
		_w6578_,
		_w6580_,
		_w6583_,
		_w6584_
	);
	LUT3 #(
		.INIT('h02)
	) name5235 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w3682_,
		_w3683_,
		_w6585_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5236 (
		_w3479_,
		_w3480_,
		_w3684_,
		_w6585_,
		_w6586_
	);
	LUT3 #(
		.INIT('h32)
	) name5237 (
		_w4953_,
		_w5078_,
		_w6586_,
		_w6587_
	);
	LUT3 #(
		.INIT('hc4)
	) name5238 (
		_w3407_,
		_w3679_,
		_w6586_,
		_w6588_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5239 (
		_w3578_,
		_w6484_,
		_w6483_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name5240 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w3545_,
		_w6590_
	);
	LUT4 #(
		.INIT('hc055)
	) name5241 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3682_,
		_w6591_
	);
	LUT3 #(
		.INIT('h31)
	) name5242 (
		_w2248_,
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('h1f)
	) name5243 (
		_w6587_,
		_w6589_,
		_w6592_,
		_w6593_
	);
	LUT3 #(
		.INIT('h02)
	) name5244 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w3682_,
		_w3712_,
		_w6594_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5245 (
		_w3479_,
		_w3480_,
		_w3713_,
		_w6594_,
		_w6595_
	);
	LUT3 #(
		.INIT('h32)
	) name5246 (
		_w4953_,
		_w5089_,
		_w6595_,
		_w6596_
	);
	LUT3 #(
		.INIT('hc4)
	) name5247 (
		_w3407_,
		_w3709_,
		_w6595_,
		_w6597_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5248 (
		_w3667_,
		_w6484_,
		_w6483_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name5249 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w3545_,
		_w6599_
	);
	LUT4 #(
		.INIT('hc055)
	) name5250 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3712_,
		_w6600_
	);
	LUT3 #(
		.INIT('h31)
	) name5251 (
		_w2248_,
		_w6599_,
		_w6600_,
		_w6601_
	);
	LUT3 #(
		.INIT('h1f)
	) name5252 (
		_w6596_,
		_w6598_,
		_w6601_,
		_w6602_
	);
	LUT3 #(
		.INIT('h02)
	) name5253 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w3712_,
		_w3727_,
		_w6603_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5254 (
		_w3479_,
		_w3480_,
		_w3728_,
		_w6603_,
		_w6604_
	);
	LUT3 #(
		.INIT('h32)
	) name5255 (
		_w4953_,
		_w5100_,
		_w6604_,
		_w6605_
	);
	LUT3 #(
		.INIT('hc4)
	) name5256 (
		_w3407_,
		_w3724_,
		_w6604_,
		_w6606_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5257 (
		_w3683_,
		_w6484_,
		_w6483_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h2)
	) name5258 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w3545_,
		_w6608_
	);
	LUT4 #(
		.INIT('hc055)
	) name5259 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3727_,
		_w6609_
	);
	LUT3 #(
		.INIT('h31)
	) name5260 (
		_w2248_,
		_w6608_,
		_w6609_,
		_w6610_
	);
	LUT3 #(
		.INIT('h1f)
	) name5261 (
		_w6605_,
		_w6607_,
		_w6610_,
		_w6611_
	);
	LUT3 #(
		.INIT('h02)
	) name5262 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w3727_,
		_w3742_,
		_w6612_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5263 (
		_w3479_,
		_w3480_,
		_w3743_,
		_w6612_,
		_w6613_
	);
	LUT3 #(
		.INIT('h32)
	) name5264 (
		_w4953_,
		_w5111_,
		_w6613_,
		_w6614_
	);
	LUT3 #(
		.INIT('hc4)
	) name5265 (
		_w3407_,
		_w3739_,
		_w6613_,
		_w6615_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5266 (
		_w3682_,
		_w6484_,
		_w6483_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h2)
	) name5267 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w3545_,
		_w6617_
	);
	LUT4 #(
		.INIT('hc055)
	) name5268 (
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3742_,
		_w6618_
	);
	LUT3 #(
		.INIT('h31)
	) name5269 (
		_w2248_,
		_w6617_,
		_w6618_,
		_w6619_
	);
	LUT3 #(
		.INIT('h1f)
	) name5270 (
		_w6614_,
		_w6616_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('h02)
	) name5271 (
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w3592_,
		_w3742_,
		_w6621_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5272 (
		_w3479_,
		_w3480_,
		_w3757_,
		_w6621_,
		_w6622_
	);
	LUT3 #(
		.INIT('h32)
	) name5273 (
		_w4953_,
		_w5122_,
		_w6622_,
		_w6623_
	);
	LUT3 #(
		.INIT('hc4)
	) name5274 (
		_w3407_,
		_w3754_,
		_w6622_,
		_w6624_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5275 (
		_w3712_,
		_w6484_,
		_w6483_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h2)
	) name5276 (
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w3545_,
		_w6626_
	);
	LUT4 #(
		.INIT('hc055)
	) name5277 (
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3592_,
		_w6627_
	);
	LUT3 #(
		.INIT('h31)
	) name5278 (
		_w2248_,
		_w6626_,
		_w6627_,
		_w6628_
	);
	LUT3 #(
		.INIT('h1f)
	) name5279 (
		_w6623_,
		_w6625_,
		_w6628_,
		_w6629_
	);
	LUT3 #(
		.INIT('h02)
	) name5280 (
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w3411_,
		_w3592_,
		_w6630_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5281 (
		_w3479_,
		_w3480_,
		_w3593_,
		_w6630_,
		_w6631_
	);
	LUT3 #(
		.INIT('h32)
	) name5282 (
		_w4953_,
		_w5133_,
		_w6631_,
		_w6632_
	);
	LUT3 #(
		.INIT('hc4)
	) name5283 (
		_w3407_,
		_w3768_,
		_w6631_,
		_w6633_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5284 (
		_w3727_,
		_w6484_,
		_w6483_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w3545_,
		_w6635_
	);
	LUT4 #(
		.INIT('hc055)
	) name5286 (
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3411_,
		_w6636_
	);
	LUT3 #(
		.INIT('h31)
	) name5287 (
		_w2248_,
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT3 #(
		.INIT('h1f)
	) name5288 (
		_w6632_,
		_w6634_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h02)
	) name5289 (
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w3411_,
		_w3412_,
		_w6639_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5290 (
		_w3413_,
		_w3479_,
		_w3480_,
		_w6639_,
		_w6640_
	);
	LUT3 #(
		.INIT('h32)
	) name5291 (
		_w4953_,
		_w5144_,
		_w6640_,
		_w6641_
	);
	LUT3 #(
		.INIT('hc4)
	) name5292 (
		_w3407_,
		_w3781_,
		_w6640_,
		_w6642_
	);
	LUT4 #(
		.INIT('h1b00)
	) name5293 (
		_w3742_,
		_w6484_,
		_w6483_,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h2)
	) name5294 (
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w3545_,
		_w6644_
	);
	LUT4 #(
		.INIT('hc055)
	) name5295 (
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1701_,
		_w1714_,
		_w3412_,
		_w6645_
	);
	LUT3 #(
		.INIT('h31)
	) name5296 (
		_w2248_,
		_w6644_,
		_w6645_,
		_w6646_
	);
	LUT3 #(
		.INIT('h1f)
	) name5297 (
		_w6641_,
		_w6643_,
		_w6646_,
		_w6647_
	);
	LUT3 #(
		.INIT('ha8)
	) name5298 (
		_w2315_,
		_w6491_,
		_w6492_,
		_w6648_
	);
	LUT3 #(
		.INIT('ha8)
	) name5299 (
		_w2317_,
		_w6495_,
		_w6496_,
		_w6649_
	);
	LUT3 #(
		.INIT('ha8)
	) name5300 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6648_,
		_w6649_,
		_w6650_
	);
	LUT3 #(
		.INIT('h02)
	) name5301 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w2320_,
		_w2322_,
		_w6651_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5302 (
		_w2323_,
		_w6500_,
		_w6501_,
		_w6651_,
		_w6652_
	);
	LUT2 #(
		.INIT('h1)
	) name5303 (
		_w2327_,
		_w6652_,
		_w6653_
	);
	LUT3 #(
		.INIT('ha8)
	) name5304 (
		_w1679_,
		_w6650_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h2)
	) name5305 (
		_w2283_,
		_w6652_,
		_w6655_
	);
	LUT4 #(
		.INIT('hc055)
	) name5306 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2320_,
		_w6656_
	);
	LUT2 #(
		.INIT('h2)
	) name5307 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		_w2288_,
		_w6657_
	);
	LUT3 #(
		.INIT('h0d)
	) name5308 (
		_w2246_,
		_w6656_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h4)
	) name5309 (
		_w6655_,
		_w6658_,
		_w6659_
	);
	LUT2 #(
		.INIT('hb)
	) name5310 (
		_w6654_,
		_w6659_,
		_w6660_
	);
	LUT3 #(
		.INIT('ha8)
	) name5311 (
		_w2250_,
		_w6495_,
		_w6496_,
		_w6661_
	);
	LUT3 #(
		.INIT('ha8)
	) name5312 (
		_w2349_,
		_w6491_,
		_w6492_,
		_w6662_
	);
	LUT3 #(
		.INIT('ha8)
	) name5313 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6661_,
		_w6662_,
		_w6663_
	);
	LUT3 #(
		.INIT('h02)
	) name5314 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w2271_,
		_w2264_,
		_w6664_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5315 (
		_w2346_,
		_w6500_,
		_w6501_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('h1)
	) name5316 (
		_w2351_,
		_w6665_,
		_w6666_
	);
	LUT3 #(
		.INIT('ha8)
	) name5317 (
		_w1679_,
		_w6663_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h2)
	) name5318 (
		_w2283_,
		_w6665_,
		_w6668_
	);
	LUT4 #(
		.INIT('hc055)
	) name5319 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2271_,
		_w6669_
	);
	LUT2 #(
		.INIT('h2)
	) name5320 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		_w2288_,
		_w6670_
	);
	LUT3 #(
		.INIT('h0d)
	) name5321 (
		_w2246_,
		_w6669_,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('h4)
	) name5322 (
		_w6668_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('hb)
	) name5323 (
		_w6667_,
		_w6672_,
		_w6673_
	);
	LUT3 #(
		.INIT('ha8)
	) name5324 (
		_w2264_,
		_w6491_,
		_w6492_,
		_w6674_
	);
	LUT3 #(
		.INIT('ha8)
	) name5325 (
		_w2271_,
		_w6495_,
		_w6496_,
		_w6675_
	);
	LUT3 #(
		.INIT('ha8)
	) name5326 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6674_,
		_w6675_,
		_w6676_
	);
	LUT3 #(
		.INIT('h02)
	) name5327 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w2272_,
		_w2376_,
		_w6677_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5328 (
		_w2377_,
		_w6500_,
		_w6501_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('h1)
	) name5329 (
		_w2380_,
		_w6678_,
		_w6679_
	);
	LUT3 #(
		.INIT('ha8)
	) name5330 (
		_w1679_,
		_w6676_,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h2)
	) name5331 (
		_w2283_,
		_w6678_,
		_w6681_
	);
	LUT4 #(
		.INIT('hc055)
	) name5332 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2376_,
		_w6682_
	);
	LUT2 #(
		.INIT('h2)
	) name5333 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		_w2288_,
		_w6683_
	);
	LUT3 #(
		.INIT('h0d)
	) name5334 (
		_w2246_,
		_w6682_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h4)
	) name5335 (
		_w6681_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('hb)
	) name5336 (
		_w6680_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('ha8)
	) name5337 (
		_w2271_,
		_w6491_,
		_w6492_,
		_w6687_
	);
	LUT3 #(
		.INIT('ha8)
	) name5338 (
		_w2272_,
		_w6495_,
		_w6496_,
		_w6688_
	);
	LUT3 #(
		.INIT('ha8)
	) name5339 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT3 #(
		.INIT('h02)
	) name5340 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w2315_,
		_w2376_,
		_w6690_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5341 (
		_w2402_,
		_w6500_,
		_w6501_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name5342 (
		_w2405_,
		_w6691_,
		_w6692_
	);
	LUT3 #(
		.INIT('ha8)
	) name5343 (
		_w1679_,
		_w6689_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h2)
	) name5344 (
		_w2283_,
		_w6691_,
		_w6694_
	);
	LUT4 #(
		.INIT('hc055)
	) name5345 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2315_,
		_w6695_
	);
	LUT2 #(
		.INIT('h2)
	) name5346 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w2288_,
		_w6696_
	);
	LUT3 #(
		.INIT('h0d)
	) name5347 (
		_w2246_,
		_w6695_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name5348 (
		_w6694_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('hb)
	) name5349 (
		_w6693_,
		_w6698_,
		_w6699_
	);
	LUT3 #(
		.INIT('ha8)
	) name5350 (
		_w2272_,
		_w6491_,
		_w6492_,
		_w6700_
	);
	LUT3 #(
		.INIT('ha8)
	) name5351 (
		_w2376_,
		_w6495_,
		_w6496_,
		_w6701_
	);
	LUT3 #(
		.INIT('ha8)
	) name5352 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6700_,
		_w6701_,
		_w6702_
	);
	LUT3 #(
		.INIT('h02)
	) name5353 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w2315_,
		_w2317_,
		_w6703_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5354 (
		_w2326_,
		_w6500_,
		_w6501_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h1)
	) name5355 (
		_w2429_,
		_w6704_,
		_w6705_
	);
	LUT3 #(
		.INIT('ha8)
	) name5356 (
		_w1679_,
		_w6702_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h2)
	) name5357 (
		_w2283_,
		_w6704_,
		_w6707_
	);
	LUT4 #(
		.INIT('hc055)
	) name5358 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2317_,
		_w6708_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		_w2288_,
		_w6709_
	);
	LUT3 #(
		.INIT('h0d)
	) name5360 (
		_w2246_,
		_w6708_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h4)
	) name5361 (
		_w6707_,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('hb)
	) name5362 (
		_w6706_,
		_w6711_,
		_w6712_
	);
	LUT3 #(
		.INIT('ha8)
	) name5363 (
		_w2376_,
		_w6491_,
		_w6492_,
		_w6713_
	);
	LUT3 #(
		.INIT('ha8)
	) name5364 (
		_w2315_,
		_w6495_,
		_w6496_,
		_w6714_
	);
	LUT3 #(
		.INIT('ha8)
	) name5365 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6713_,
		_w6714_,
		_w6715_
	);
	LUT3 #(
		.INIT('h02)
	) name5366 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w2322_,
		_w2317_,
		_w6716_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5367 (
		_w2451_,
		_w6500_,
		_w6501_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		_w2454_,
		_w6717_,
		_w6718_
	);
	LUT3 #(
		.INIT('ha8)
	) name5369 (
		_w1679_,
		_w6715_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h2)
	) name5370 (
		_w2283_,
		_w6717_,
		_w6720_
	);
	LUT4 #(
		.INIT('hc055)
	) name5371 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2322_,
		_w6721_
	);
	LUT2 #(
		.INIT('h2)
	) name5372 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w2288_,
		_w6722_
	);
	LUT3 #(
		.INIT('h0d)
	) name5373 (
		_w2246_,
		_w6721_,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h4)
	) name5374 (
		_w6720_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('hb)
	) name5375 (
		_w6719_,
		_w6724_,
		_w6725_
	);
	LUT3 #(
		.INIT('ha8)
	) name5376 (
		_w2317_,
		_w6491_,
		_w6492_,
		_w6726_
	);
	LUT3 #(
		.INIT('ha8)
	) name5377 (
		_w2322_,
		_w6495_,
		_w6496_,
		_w6727_
	);
	LUT3 #(
		.INIT('ha8)
	) name5378 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT3 #(
		.INIT('h02)
	) name5379 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w2320_,
		_w2473_,
		_w6729_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5380 (
		_w2474_,
		_w6500_,
		_w6501_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name5381 (
		_w2477_,
		_w6730_,
		_w6731_
	);
	LUT3 #(
		.INIT('ha8)
	) name5382 (
		_w1679_,
		_w6728_,
		_w6731_,
		_w6732_
	);
	LUT2 #(
		.INIT('h2)
	) name5383 (
		_w2283_,
		_w6730_,
		_w6733_
	);
	LUT4 #(
		.INIT('hc055)
	) name5384 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2473_,
		_w6734_
	);
	LUT2 #(
		.INIT('h2)
	) name5385 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w2288_,
		_w6735_
	);
	LUT3 #(
		.INIT('h0d)
	) name5386 (
		_w2246_,
		_w6734_,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h4)
	) name5387 (
		_w6733_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('hb)
	) name5388 (
		_w6732_,
		_w6737_,
		_w6738_
	);
	LUT3 #(
		.INIT('ha8)
	) name5389 (
		_w2320_,
		_w6495_,
		_w6496_,
		_w6739_
	);
	LUT3 #(
		.INIT('ha8)
	) name5390 (
		_w2322_,
		_w6491_,
		_w6492_,
		_w6740_
	);
	LUT3 #(
		.INIT('ha8)
	) name5391 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6739_,
		_w6740_,
		_w6741_
	);
	LUT3 #(
		.INIT('h02)
	) name5392 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w2473_,
		_w2502_,
		_w6742_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5393 (
		_w2503_,
		_w6500_,
		_w6501_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w2506_,
		_w6743_,
		_w6744_
	);
	LUT3 #(
		.INIT('ha8)
	) name5395 (
		_w1679_,
		_w6741_,
		_w6744_,
		_w6745_
	);
	LUT2 #(
		.INIT('h2)
	) name5396 (
		_w2283_,
		_w6743_,
		_w6746_
	);
	LUT4 #(
		.INIT('hc055)
	) name5397 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2502_,
		_w6747_
	);
	LUT2 #(
		.INIT('h2)
	) name5398 (
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w2288_,
		_w6748_
	);
	LUT3 #(
		.INIT('h0d)
	) name5399 (
		_w2246_,
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h4)
	) name5400 (
		_w6746_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('hb)
	) name5401 (
		_w6745_,
		_w6750_,
		_w6751_
	);
	LUT3 #(
		.INIT('ha8)
	) name5402 (
		_w2320_,
		_w6491_,
		_w6492_,
		_w6752_
	);
	LUT3 #(
		.INIT('ha8)
	) name5403 (
		_w2473_,
		_w6495_,
		_w6496_,
		_w6753_
	);
	LUT3 #(
		.INIT('ha8)
	) name5404 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6752_,
		_w6753_,
		_w6754_
	);
	LUT3 #(
		.INIT('h02)
	) name5405 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w2502_,
		_w2528_,
		_w6755_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5406 (
		_w2529_,
		_w6500_,
		_w6501_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h1)
	) name5407 (
		_w2532_,
		_w6756_,
		_w6757_
	);
	LUT3 #(
		.INIT('ha8)
	) name5408 (
		_w1679_,
		_w6754_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h2)
	) name5409 (
		_w2283_,
		_w6756_,
		_w6759_
	);
	LUT4 #(
		.INIT('hc055)
	) name5410 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2528_,
		_w6760_
	);
	LUT2 #(
		.INIT('h2)
	) name5411 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w2288_,
		_w6761_
	);
	LUT3 #(
		.INIT('h0d)
	) name5412 (
		_w2246_,
		_w6760_,
		_w6761_,
		_w6762_
	);
	LUT2 #(
		.INIT('h4)
	) name5413 (
		_w6759_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('hb)
	) name5414 (
		_w6758_,
		_w6763_,
		_w6764_
	);
	LUT3 #(
		.INIT('ha8)
	) name5415 (
		_w2473_,
		_w6491_,
		_w6492_,
		_w6765_
	);
	LUT3 #(
		.INIT('ha8)
	) name5416 (
		_w2502_,
		_w6495_,
		_w6496_,
		_w6766_
	);
	LUT3 #(
		.INIT('ha8)
	) name5417 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT3 #(
		.INIT('h02)
	) name5418 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w2528_,
		_w2554_,
		_w6768_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5419 (
		_w2555_,
		_w6500_,
		_w6501_,
		_w6768_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w2558_,
		_w6769_,
		_w6770_
	);
	LUT3 #(
		.INIT('ha8)
	) name5421 (
		_w1679_,
		_w6767_,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		_w2283_,
		_w6769_,
		_w6772_
	);
	LUT4 #(
		.INIT('hc055)
	) name5423 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2554_,
		_w6773_
	);
	LUT2 #(
		.INIT('h2)
	) name5424 (
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w2288_,
		_w6774_
	);
	LUT3 #(
		.INIT('h0d)
	) name5425 (
		_w2246_,
		_w6773_,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h4)
	) name5426 (
		_w6772_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('hb)
	) name5427 (
		_w6771_,
		_w6776_,
		_w6777_
	);
	LUT3 #(
		.INIT('ha8)
	) name5428 (
		_w2502_,
		_w6491_,
		_w6492_,
		_w6778_
	);
	LUT3 #(
		.INIT('ha8)
	) name5429 (
		_w2528_,
		_w6495_,
		_w6496_,
		_w6779_
	);
	LUT3 #(
		.INIT('ha8)
	) name5430 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6778_,
		_w6779_,
		_w6780_
	);
	LUT3 #(
		.INIT('h02)
	) name5431 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w2554_,
		_w2580_,
		_w6781_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5432 (
		_w2581_,
		_w6500_,
		_w6501_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h1)
	) name5433 (
		_w2584_,
		_w6782_,
		_w6783_
	);
	LUT3 #(
		.INIT('ha8)
	) name5434 (
		_w1679_,
		_w6780_,
		_w6783_,
		_w6784_
	);
	LUT2 #(
		.INIT('h2)
	) name5435 (
		_w2283_,
		_w6782_,
		_w6785_
	);
	LUT4 #(
		.INIT('hc055)
	) name5436 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2580_,
		_w6786_
	);
	LUT2 #(
		.INIT('h2)
	) name5437 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w2288_,
		_w6787_
	);
	LUT3 #(
		.INIT('h0d)
	) name5438 (
		_w2246_,
		_w6786_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h4)
	) name5439 (
		_w6785_,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('hb)
	) name5440 (
		_w6784_,
		_w6789_,
		_w6790_
	);
	LUT3 #(
		.INIT('ha8)
	) name5441 (
		_w2528_,
		_w6491_,
		_w6492_,
		_w6791_
	);
	LUT3 #(
		.INIT('ha8)
	) name5442 (
		_w2554_,
		_w6495_,
		_w6496_,
		_w6792_
	);
	LUT3 #(
		.INIT('ha8)
	) name5443 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6791_,
		_w6792_,
		_w6793_
	);
	LUT3 #(
		.INIT('h02)
	) name5444 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w2580_,
		_w2606_,
		_w6794_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5445 (
		_w2607_,
		_w6500_,
		_w6501_,
		_w6794_,
		_w6795_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w2610_,
		_w6795_,
		_w6796_
	);
	LUT3 #(
		.INIT('ha8)
	) name5447 (
		_w1679_,
		_w6793_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h2)
	) name5448 (
		_w2283_,
		_w6795_,
		_w6798_
	);
	LUT4 #(
		.INIT('hc055)
	) name5449 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2606_,
		_w6799_
	);
	LUT2 #(
		.INIT('h2)
	) name5450 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w2288_,
		_w6800_
	);
	LUT3 #(
		.INIT('h0d)
	) name5451 (
		_w2246_,
		_w6799_,
		_w6800_,
		_w6801_
	);
	LUT2 #(
		.INIT('h4)
	) name5452 (
		_w6798_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('hb)
	) name5453 (
		_w6797_,
		_w6802_,
		_w6803_
	);
	LUT3 #(
		.INIT('ha8)
	) name5454 (
		_w2554_,
		_w6491_,
		_w6492_,
		_w6804_
	);
	LUT3 #(
		.INIT('ha8)
	) name5455 (
		_w2580_,
		_w6495_,
		_w6496_,
		_w6805_
	);
	LUT3 #(
		.INIT('ha8)
	) name5456 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT3 #(
		.INIT('h02)
	) name5457 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w2349_,
		_w2606_,
		_w6807_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5458 (
		_w2632_,
		_w6500_,
		_w6501_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		_w2635_,
		_w6808_,
		_w6809_
	);
	LUT3 #(
		.INIT('ha8)
	) name5460 (
		_w1679_,
		_w6806_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h2)
	) name5461 (
		_w2283_,
		_w6808_,
		_w6811_
	);
	LUT4 #(
		.INIT('hc055)
	) name5462 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2349_,
		_w6812_
	);
	LUT2 #(
		.INIT('h2)
	) name5463 (
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w2288_,
		_w6813_
	);
	LUT3 #(
		.INIT('h0d)
	) name5464 (
		_w2246_,
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h4)
	) name5465 (
		_w6811_,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('hb)
	) name5466 (
		_w6810_,
		_w6815_,
		_w6816_
	);
	LUT3 #(
		.INIT('ha8)
	) name5467 (
		_w2580_,
		_w6491_,
		_w6492_,
		_w6817_
	);
	LUT3 #(
		.INIT('ha8)
	) name5468 (
		_w2606_,
		_w6495_,
		_w6496_,
		_w6818_
	);
	LUT3 #(
		.INIT('ha8)
	) name5469 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6817_,
		_w6818_,
		_w6819_
	);
	LUT3 #(
		.INIT('h02)
	) name5470 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w2250_,
		_w2349_,
		_w6820_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5471 (
		_w2350_,
		_w6500_,
		_w6501_,
		_w6820_,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w2659_,
		_w6821_,
		_w6822_
	);
	LUT3 #(
		.INIT('ha8)
	) name5473 (
		_w1679_,
		_w6819_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h2)
	) name5474 (
		_w2283_,
		_w6821_,
		_w6824_
	);
	LUT4 #(
		.INIT('hc055)
	) name5475 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2250_,
		_w6825_
	);
	LUT2 #(
		.INIT('h2)
	) name5476 (
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w2288_,
		_w6826_
	);
	LUT3 #(
		.INIT('h0d)
	) name5477 (
		_w2246_,
		_w6825_,
		_w6826_,
		_w6827_
	);
	LUT2 #(
		.INIT('h4)
	) name5478 (
		_w6824_,
		_w6827_,
		_w6828_
	);
	LUT2 #(
		.INIT('hb)
	) name5479 (
		_w6823_,
		_w6828_,
		_w6829_
	);
	LUT3 #(
		.INIT('ha8)
	) name5480 (
		_w2606_,
		_w6491_,
		_w6492_,
		_w6830_
	);
	LUT3 #(
		.INIT('ha8)
	) name5481 (
		_w2349_,
		_w6495_,
		_w6496_,
		_w6831_
	);
	LUT3 #(
		.INIT('ha8)
	) name5482 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT3 #(
		.INIT('h02)
	) name5483 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w2250_,
		_w2264_,
		_w6833_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5484 (
		_w2279_,
		_w6500_,
		_w6501_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w2683_,
		_w6834_,
		_w6835_
	);
	LUT3 #(
		.INIT('ha8)
	) name5486 (
		_w1679_,
		_w6832_,
		_w6835_,
		_w6836_
	);
	LUT2 #(
		.INIT('h2)
	) name5487 (
		_w2283_,
		_w6834_,
		_w6837_
	);
	LUT4 #(
		.INIT('hc055)
	) name5488 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1542_,
		_w1547_,
		_w2264_,
		_w6838_
	);
	LUT2 #(
		.INIT('h2)
	) name5489 (
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w2288_,
		_w6839_
	);
	LUT3 #(
		.INIT('h0d)
	) name5490 (
		_w2246_,
		_w6838_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h4)
	) name5491 (
		_w6837_,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('hb)
	) name5492 (
		_w6836_,
		_w6841_,
		_w6842_
	);
	LUT3 #(
		.INIT('h08)
	) name5493 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w1592_,
		_w1660_,
		_w6843_
	);
	LUT2 #(
		.INIT('h2)
	) name5494 (
		_w4354_,
		_w5697_,
		_w6844_
	);
	LUT4 #(
		.INIT('h4000)
	) name5495 (
		_w4346_,
		_w4821_,
		_w4826_,
		_w5695_,
		_w6845_
	);
	LUT4 #(
		.INIT('h0001)
	) name5496 (
		_w4345_,
		_w4349_,
		_w4351_,
		_w4354_,
		_w6846_
	);
	LUT3 #(
		.INIT('h15)
	) name5497 (
		_w4214_,
		_w6845_,
		_w6846_,
		_w6847_
	);
	LUT3 #(
		.INIT('h6a)
	) name5498 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4255_,
		_w4263_,
		_w6848_
	);
	LUT2 #(
		.INIT('h8)
	) name5499 (
		_w4263_,
		_w4898_,
		_w6849_
	);
	LUT3 #(
		.INIT('h80)
	) name5500 (
		_w4796_,
		_w4896_,
		_w6849_,
		_w6850_
	);
	LUT4 #(
		.INIT('h1551)
	) name5501 (
		_w1661_,
		_w4214_,
		_w6848_,
		_w6850_,
		_w6851_
	);
	LUT4 #(
		.INIT('h1055)
	) name5502 (
		_w6843_,
		_w6844_,
		_w6847_,
		_w6851_,
		_w6852_
	);
	LUT4 #(
		.INIT('h028a)
	) name5503 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w6853_
	);
	LUT4 #(
		.INIT('h28a0)
	) name5504 (
		_w1659_,
		_w4876_,
		_w4912_,
		_w5715_,
		_w6854_
	);
	LUT2 #(
		.INIT('h1)
	) name5505 (
		_w6853_,
		_w6854_,
		_w6855_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5506 (
		_w1559_,
		_w1678_,
		_w6852_,
		_w6855_,
		_w6856_
	);
	LUT2 #(
		.INIT('h1)
	) name5507 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w6857_
	);
	LUT4 #(
		.INIT('h0080)
	) name5508 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w5734_,
		_w6857_,
		_w6858_
	);
	LUT3 #(
		.INIT('h48)
	) name5509 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w1679_,
		_w6858_,
		_w6859_
	);
	LUT4 #(
		.INIT('h8000)
	) name5510 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w5734_,
		_w6860_
	);
	LUT3 #(
		.INIT('h6c)
	) name5511 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w5735_,
		_w6861_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5512 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		_w2283_,
		_w5735_,
		_w6862_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5513 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2286_,
		_w5747_,
		_w6863_
	);
	LUT3 #(
		.INIT('h10)
	) name5514 (
		_w6862_,
		_w6859_,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('hb)
	) name5515 (
		_w6856_,
		_w6864_,
		_w6865_
	);
	LUT3 #(
		.INIT('h08)
	) name5516 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w1592_,
		_w1660_,
		_w6866_
	);
	LUT3 #(
		.INIT('h40)
	) name5517 (
		_w4356_,
		_w4362_,
		_w4363_,
		_w6867_
	);
	LUT3 #(
		.INIT('h80)
	) name5518 (
		_w6845_,
		_w6846_,
		_w6867_,
		_w6868_
	);
	LUT4 #(
		.INIT('h5150)
	) name5519 (
		_w4214_,
		_w4360_,
		_w4363_,
		_w4906_,
		_w6869_
	);
	LUT4 #(
		.INIT('h8000)
	) name5520 (
		_w4274_,
		_w4796_,
		_w4896_,
		_w4900_,
		_w6870_
	);
	LUT4 #(
		.INIT('h1555)
	) name5521 (
		_w4274_,
		_w4796_,
		_w4896_,
		_w4900_,
		_w6871_
	);
	LUT3 #(
		.INIT('h02)
	) name5522 (
		_w4214_,
		_w6871_,
		_w6870_,
		_w6872_
	);
	LUT4 #(
		.INIT('h5510)
	) name5523 (
		_w1661_,
		_w6868_,
		_w6869_,
		_w6872_,
		_w6873_
	);
	LUT4 #(
		.INIT('h028a)
	) name5524 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w6874_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5525 (
		_w1659_,
		_w4426_,
		_w5716_,
		_w6874_,
		_w6875_
	);
	LUT4 #(
		.INIT('h5700)
	) name5526 (
		_w1559_,
		_w6866_,
		_w6873_,
		_w6875_,
		_w6876_
	);
	LUT4 #(
		.INIT('h00ec)
	) name5527 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w5738_,
		_w5743_,
		_w6877_
	);
	LUT4 #(
		.INIT('h8848)
	) name5528 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		_w1679_,
		_w5738_,
		_w6857_,
		_w6878_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5529 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2286_,
		_w5747_,
		_w6879_
	);
	LUT4 #(
		.INIT('h1300)
	) name5530 (
		_w2283_,
		_w6878_,
		_w6877_,
		_w6879_,
		_w6880_
	);
	LUT3 #(
		.INIT('h2f)
	) name5531 (
		_w1678_,
		_w6876_,
		_w6880_,
		_w6881_
	);
	LUT3 #(
		.INIT('h08)
	) name5532 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w1592_,
		_w1660_,
		_w6882_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		_w4333_,
		_w4819_,
		_w6883_
	);
	LUT2 #(
		.INIT('h4)
	) name5534 (
		_w4346_,
		_w5694_,
		_w6884_
	);
	LUT4 #(
		.INIT('h8000)
	) name5535 (
		_w4818_,
		_w4903_,
		_w6883_,
		_w6884_,
		_w6885_
	);
	LUT3 #(
		.INIT('h04)
	) name5536 (
		_w4356_,
		_w4362_,
		_w4363_,
		_w6886_
	);
	LUT4 #(
		.INIT('h4000)
	) name5537 (
		_w4365_,
		_w6846_,
		_w6885_,
		_w6886_,
		_w6887_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5538 (
		_w4365_,
		_w6846_,
		_w6885_,
		_w6886_,
		_w6888_
	);
	LUT3 #(
		.INIT('h01)
	) name5539 (
		_w4214_,
		_w6888_,
		_w6887_,
		_w6889_
	);
	LUT3 #(
		.INIT('h6a)
	) name5540 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4269_,
		_w4272_,
		_w6890_
	);
	LUT4 #(
		.INIT('h8884)
	) name5541 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4214_,
		_w4273_,
		_w6870_,
		_w6891_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		_w1661_,
		_w6891_,
		_w6892_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5543 (
		_w1559_,
		_w6882_,
		_w6889_,
		_w6892_,
		_w6893_
	);
	LUT4 #(
		.INIT('h028a)
	) name5544 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w6894_
	);
	LUT2 #(
		.INIT('h6)
	) name5545 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4425_,
		_w6895_
	);
	LUT2 #(
		.INIT('h8)
	) name5546 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		_w4834_,
		_w6896_
	);
	LUT4 #(
		.INIT('h4000)
	) name5547 (
		_w4869_,
		_w5874_,
		_w5875_,
		_w6896_,
		_w6897_
	);
	LUT3 #(
		.INIT('h6c)
	) name5548 (
		\P2_InstAddrPointer_reg[15]/NET0131 ,
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4410_,
		_w6898_
	);
	LUT3 #(
		.INIT('h6a)
	) name5549 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4254_,
		_w4410_,
		_w6899_
	);
	LUT2 #(
		.INIT('h8)
	) name5550 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w6900_
	);
	LUT4 #(
		.INIT('h6a00)
	) name5551 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w4254_,
		_w4410_,
		_w6900_,
		_w6901_
	);
	LUT2 #(
		.INIT('h8)
	) name5552 (
		_w4420_,
		_w6901_,
		_w6902_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5553 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w4424_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h8)
	) name5554 (
		_w4914_,
		_w6903_,
		_w6904_
	);
	LUT4 #(
		.INIT('h8000)
	) name5555 (
		_w4414_,
		_w6897_,
		_w6898_,
		_w6904_,
		_w6905_
	);
	LUT4 #(
		.INIT('h3113)
	) name5556 (
		_w1659_,
		_w6894_,
		_w6895_,
		_w6905_,
		_w6906_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5557 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w2242_,
		_w5738_,
		_w6907_
	);
	LUT2 #(
		.INIT('h6)
	) name5558 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5743_,
		_w6908_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5559 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w2286_,
		_w5747_,
		_w6909_
	);
	LUT4 #(
		.INIT('h9f00)
	) name5560 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5743_,
		_w5746_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		_w6907_,
		_w6910_,
		_w6911_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5562 (
		_w1678_,
		_w6893_,
		_w6906_,
		_w6911_,
		_w6912_
	);
	LUT3 #(
		.INIT('h08)
	) name5563 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w1592_,
		_w1660_,
		_w6913_
	);
	LUT4 #(
		.INIT('haa20)
	) name5564 (
		_w1559_,
		_w4280_,
		_w4370_,
		_w6913_,
		_w6914_
	);
	LUT4 #(
		.INIT('h028a)
	) name5565 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w6915_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5566 (
		_w1659_,
		_w4431_,
		_w4432_,
		_w6915_,
		_w6916_
	);
	LUT4 #(
		.INIT('h0080)
	) name5567 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		_w5738_,
		_w6857_,
		_w6917_
	);
	LUT3 #(
		.INIT('h48)
	) name5568 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w1679_,
		_w6917_,
		_w6918_
	);
	LUT3 #(
		.INIT('h6c)
	) name5569 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w5743_,
		_w6919_
	);
	LUT4 #(
		.INIT('h60c0)
	) name5570 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		_w2283_,
		_w5743_,
		_w6920_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5571 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2286_,
		_w5747_,
		_w6921_
	);
	LUT2 #(
		.INIT('h4)
	) name5572 (
		_w6920_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h4)
	) name5573 (
		_w6918_,
		_w6922_,
		_w6923_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5574 (
		_w1678_,
		_w6914_,
		_w6916_,
		_w6923_,
		_w6924_
	);
	LUT4 #(
		.INIT('h8000)
	) name5575 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		_w3025_,
		_w3028_,
		_w3032_,
		_w6925_
	);
	LUT2 #(
		.INIT('h6)
	) name5576 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3033_,
		_w6926_
	);
	LUT4 #(
		.INIT('h4448)
	) name5577 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2181_,
		_w3033_,
		_w6925_,
		_w6927_
	);
	LUT3 #(
		.INIT('h02)
	) name5578 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6928_
	);
	LUT4 #(
		.INIT('h0080)
	) name5579 (
		_w2874_,
		_w2884_,
		_w2897_,
		_w2913_,
		_w6929_
	);
	LUT4 #(
		.INIT('h0081)
	) name5580 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_InstAddrPointer_reg[21]/NET0131 ,
		_w2899_,
		_w2907_,
		_w6930_
	);
	LUT3 #(
		.INIT('h2a)
	) name5581 (
		_w2906_,
		_w6929_,
		_w6930_,
		_w6931_
	);
	LUT3 #(
		.INIT('h15)
	) name5582 (
		_w2755_,
		_w5380_,
		_w6929_,
		_w6932_
	);
	LUT4 #(
		.INIT('h802a)
	) name5583 (
		_w2755_,
		_w2960_,
		_w2968_,
		_w2971_,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w2173_,
		_w6933_,
		_w6934_
	);
	LUT4 #(
		.INIT('h1055)
	) name5585 (
		_w6928_,
		_w6931_,
		_w6932_,
		_w6934_,
		_w6935_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5586 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w6936_
	);
	LUT4 #(
		.INIT('h000d)
	) name5587 (
		_w2171_,
		_w6935_,
		_w6936_,
		_w6927_,
		_w6937_
	);
	LUT2 #(
		.INIT('h1)
	) name5588 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w6938_
	);
	LUT3 #(
		.INIT('h08)
	) name5589 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w6938_,
		_w6939_
	);
	LUT3 #(
		.INIT('h48)
	) name5590 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w2194_,
		_w6939_,
		_w6940_
	);
	LUT3 #(
		.INIT('h80)
	) name5591 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w6941_
	);
	LUT4 #(
		.INIT('h8000)
	) name5592 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5771_,
		_w6942_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5593 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5771_,
		_w6943_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5594 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w3054_,
		_w5783_,
		_w6944_
	);
	LUT3 #(
		.INIT('h70)
	) name5595 (
		_w3055_,
		_w6943_,
		_w6944_,
		_w6945_
	);
	LUT2 #(
		.INIT('h4)
	) name5596 (
		_w6940_,
		_w6945_,
		_w6946_
	);
	LUT3 #(
		.INIT('h2f)
	) name5597 (
		_w1945_,
		_w6937_,
		_w6946_,
		_w6947_
	);
	LUT4 #(
		.INIT('h8000)
	) name5598 (
		_w3025_,
		_w3028_,
		_w3036_,
		_w3040_,
		_w6948_
	);
	LUT3 #(
		.INIT('h28)
	) name5599 (
		_w2181_,
		_w3042_,
		_w6948_,
		_w6949_
	);
	LUT3 #(
		.INIT('h02)
	) name5600 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6950_
	);
	LUT3 #(
		.INIT('h41)
	) name5601 (
		_w2755_,
		_w2728_,
		_w2915_,
		_w6951_
	);
	LUT4 #(
		.INIT('h1551)
	) name5602 (
		_w2173_,
		_w2755_,
		_w2974_,
		_w2975_,
		_w6952_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5603 (
		_w2171_,
		_w6950_,
		_w6951_,
		_w6952_,
		_w6953_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5604 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w6954_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5605 (
		_w1945_,
		_w6953_,
		_w6954_,
		_w6949_,
		_w6955_
	);
	LUT2 #(
		.INIT('h6)
	) name5606 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w5775_,
		_w6956_
	);
	LUT3 #(
		.INIT('h48)
	) name5607 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w3055_,
		_w5775_,
		_w6957_
	);
	LUT4 #(
		.INIT('h0080)
	) name5608 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w5774_,
		_w6938_,
		_w6958_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5609 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w3054_,
		_w5783_,
		_w6959_
	);
	LUT4 #(
		.INIT('hb700)
	) name5610 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w2194_,
		_w6958_,
		_w6959_,
		_w6960_
	);
	LUT2 #(
		.INIT('h4)
	) name5611 (
		_w6957_,
		_w6960_,
		_w6961_
	);
	LUT2 #(
		.INIT('hb)
	) name5612 (
		_w6955_,
		_w6961_,
		_w6962_
	);
	LUT3 #(
		.INIT('h02)
	) name5613 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2103_,
		_w2172_,
		_w6963_
	);
	LUT3 #(
		.INIT('ha8)
	) name5614 (
		_w2171_,
		_w4080_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5615 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w6965_
	);
	LUT3 #(
		.INIT('h0b)
	) name5616 (
		_w4091_,
		_w4092_,
		_w6965_,
		_w6966_
	);
	LUT3 #(
		.INIT('h6c)
	) name5617 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5775_,
		_w6967_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5618 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5775_,
		_w6350_,
		_w6968_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5619 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w3054_,
		_w5783_,
		_w6969_
	);
	LUT4 #(
		.INIT('hb700)
	) name5620 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w2199_,
		_w5777_,
		_w6969_,
		_w6970_
	);
	LUT2 #(
		.INIT('h4)
	) name5621 (
		_w6968_,
		_w6970_,
		_w6971_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5622 (
		_w1945_,
		_w6964_,
		_w6966_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('h8)
	) name5623 (
		_w2730_,
		_w2912_,
		_w6973_
	);
	LUT4 #(
		.INIT('h4111)
	) name5624 (
		_w2755_,
		_w2731_,
		_w5350_,
		_w6973_,
		_w6974_
	);
	LUT3 #(
		.INIT('h6a)
	) name5625 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2724_,
		_w2703_,
		_w6975_
	);
	LUT3 #(
		.INIT('h80)
	) name5626 (
		_w2964_,
		_w2973_,
		_w2976_,
		_w6976_
	);
	LUT4 #(
		.INIT('h820a)
	) name5627 (
		_w2755_,
		_w5363_,
		_w6975_,
		_w6976_,
		_w6977_
	);
	LUT4 #(
		.INIT('h7774)
	) name5628 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w2173_,
		_w6977_,
		_w6974_,
		_w6978_
	);
	LUT2 #(
		.INIT('h2)
	) name5629 (
		_w2171_,
		_w6978_,
		_w6979_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5630 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w6980_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name5631 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2703_,
		_w3038_,
		_w6981_
	);
	LUT3 #(
		.INIT('h07)
	) name5632 (
		_w3043_,
		_w6948_,
		_w6981_,
		_w6982_
	);
	LUT3 #(
		.INIT('h2a)
	) name5633 (
		_w2181_,
		_w3044_,
		_w6948_,
		_w6983_
	);
	LUT3 #(
		.INIT('h45)
	) name5634 (
		_w6980_,
		_w6982_,
		_w6983_,
		_w6984_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5635 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5775_,
		_w6985_
	);
	LUT3 #(
		.INIT('h6c)
	) name5636 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		_w5777_,
		_w6986_
	);
	LUT4 #(
		.INIT('hc840)
	) name5637 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w6985_,
		_w6986_,
		_w6987_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5638 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w3054_,
		_w5783_,
		_w6988_
	);
	LUT3 #(
		.INIT('h70)
	) name5639 (
		_w3055_,
		_w6985_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h4)
	) name5640 (
		_w6987_,
		_w6989_,
		_w6990_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5641 (
		_w1945_,
		_w6979_,
		_w6984_,
		_w6990_,
		_w6991_
	);
	LUT4 #(
		.INIT('h4447)
	) name5642 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w1916_,
		_w4471_,
		_w4479_,
		_w6992_
	);
	LUT4 #(
		.INIT('h028a)
	) name5643 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w6993_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5644 (
		_w1924_,
		_w4481_,
		_w4483_,
		_w6993_,
		_w6994_
	);
	LUT4 #(
		.INIT('h08cc)
	) name5645 (
		_w1810_,
		_w1933_,
		_w6992_,
		_w6994_,
		_w6995_
	);
	LUT4 #(
		.INIT('h8000)
	) name5646 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w6363_,
		_w6372_,
		_w6996_
	);
	LUT4 #(
		.INIT('h8000)
	) name5647 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6363_,
		_w6361_,
		_w6372_,
		_w6997_
	);
	LUT3 #(
		.INIT('h6c)
	) name5648 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6373_,
		_w6998_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5649 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6373_,
		_w6378_,
		_w6999_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name5650 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w2310_,
		_w6379_,
		_w6363_,
		_w7000_
	);
	LUT3 #(
		.INIT('ha2)
	) name5651 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6383_,
		_w7000_,
		_w7001_
	);
	LUT3 #(
		.INIT('h20)
	) name5652 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w1939_,
		_w7002_
	);
	LUT4 #(
		.INIT('h8000)
	) name5653 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w6379_,
		_w6363_,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w4497_,
		_w7003_,
		_w7004_
	);
	LUT3 #(
		.INIT('h10)
	) name5655 (
		_w7001_,
		_w6999_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('hb)
	) name5656 (
		_w6995_,
		_w7005_,
		_w7006_
	);
	LUT3 #(
		.INIT('h08)
	) name5657 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7007_
	);
	LUT3 #(
		.INIT('h80)
	) name5658 (
		_w3316_,
		_w3318_,
		_w4451_,
		_w7008_
	);
	LUT3 #(
		.INIT('h15)
	) name5659 (
		_w3314_,
		_w5458_,
		_w7008_,
		_w7009_
	);
	LUT4 #(
		.INIT('h4080)
	) name5660 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3077_,
		_w7010_
	);
	LUT2 #(
		.INIT('h8)
	) name5661 (
		_w3314_,
		_w7010_,
		_w7011_
	);
	LUT3 #(
		.INIT('h2a)
	) name5662 (
		_w3101_,
		_w4470_,
		_w7011_,
		_w7012_
	);
	LUT2 #(
		.INIT('h1)
	) name5663 (
		_w3252_,
		_w3259_,
		_w7013_
	);
	LUT4 #(
		.INIT('h0200)
	) name5664 (
		_w3239_,
		_w3240_,
		_w3250_,
		_w7013_,
		_w7014_
	);
	LUT4 #(
		.INIT('h8000)
	) name5665 (
		_w3248_,
		_w4474_,
		_w4475_,
		_w7014_,
		_w7015_
	);
	LUT3 #(
		.INIT('h14)
	) name5666 (
		_w3101_,
		_w3260_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('h5510)
	) name5667 (
		_w1916_,
		_w7009_,
		_w7012_,
		_w7016_,
		_w7017_
	);
	LUT4 #(
		.INIT('h028a)
	) name5668 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7018_
	);
	LUT4 #(
		.INIT('h4080)
	) name5669 (
		\P1_InstAddrPointer_reg[24]/NET0131 ,
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_InstAddrPointer_reg[26]/NET0131 ,
		_w3378_,
		_w7019_
	);
	LUT3 #(
		.INIT('h80)
	) name5670 (
		_w4481_,
		_w4483_,
		_w7019_,
		_w7020_
	);
	LUT4 #(
		.INIT('h0d07)
	) name5671 (
		_w1924_,
		_w3388_,
		_w7018_,
		_w7020_,
		_w7021_
	);
	LUT4 #(
		.INIT('h5700)
	) name5672 (
		_w1810_,
		_w7007_,
		_w7017_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h13)
	) name5673 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w6374_,
		_w7023_
	);
	LUT3 #(
		.INIT('h80)
	) name5674 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w6380_,
		_w7024_
	);
	LUT2 #(
		.INIT('h1)
	) name5675 (
		_w7023_,
		_w7024_,
		_w7025_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5676 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7026_
	);
	LUT4 #(
		.INIT('hb700)
	) name5677 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w2310_,
		_w6380_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5678 (
		_w6378_,
		_w7023_,
		_w7024_,
		_w7027_,
		_w7028_
	);
	LUT3 #(
		.INIT('h2f)
	) name5679 (
		_w1933_,
		_w7022_,
		_w7028_,
		_w7029_
	);
	LUT2 #(
		.INIT('h6)
	) name5680 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w3080_,
		_w7030_
	);
	LUT4 #(
		.INIT('h802a)
	) name5681 (
		_w3101_,
		_w4470_,
		_w7011_,
		_w7030_,
		_w7031_
	);
	LUT4 #(
		.INIT('h0200)
	) name5682 (
		_w3239_,
		_w3240_,
		_w3260_,
		_w7013_,
		_w7032_
	);
	LUT4 #(
		.INIT('h4111)
	) name5683 (
		_w3101_,
		_w3258_,
		_w4729_,
		_w7032_,
		_w7033_
	);
	LUT4 #(
		.INIT('h7774)
	) name5684 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w1916_,
		_w7033_,
		_w7031_,
		_w7034_
	);
	LUT4 #(
		.INIT('h028a)
	) name5685 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7035_
	);
	LUT4 #(
		.INIT('h28a0)
	) name5686 (
		_w1924_,
		_w4031_,
		_w4032_,
		_w4738_,
		_w7036_
	);
	LUT4 #(
		.INIT('h000d)
	) name5687 (
		_w1810_,
		_w7034_,
		_w7035_,
		_w7036_,
		_w7037_
	);
	LUT4 #(
		.INIT('h8000)
	) name5688 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w6380_,
		_w7038_
	);
	LUT4 #(
		.INIT('h78f0)
	) name5689 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w6380_,
		_w7039_
	);
	LUT2 #(
		.INIT('h8)
	) name5690 (
		_w3407_,
		_w7039_,
		_w7040_
	);
	LUT2 #(
		.INIT('h1)
	) name5691 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w7041_
	);
	LUT3 #(
		.INIT('h08)
	) name5692 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w6380_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5693 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7043_
	);
	LUT4 #(
		.INIT('hb700)
	) name5694 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		_w1939_,
		_w7042_,
		_w7043_,
		_w7044_
	);
	LUT2 #(
		.INIT('h4)
	) name5695 (
		_w7040_,
		_w7044_,
		_w7045_
	);
	LUT3 #(
		.INIT('h2f)
	) name5696 (
		_w1933_,
		_w7037_,
		_w7045_,
		_w7046_
	);
	LUT3 #(
		.INIT('h08)
	) name5697 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7047_
	);
	LUT4 #(
		.INIT('haa20)
	) name5698 (
		_w1810_,
		_w3999_,
		_w4013_,
		_w7047_,
		_w7048_
	);
	LUT4 #(
		.INIT('h028a)
	) name5699 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7049_
	);
	LUT4 #(
		.INIT('h00d7)
	) name5700 (
		_w1924_,
		_w4015_,
		_w4034_,
		_w7049_,
		_w7050_
	);
	LUT3 #(
		.INIT('h32)
	) name5701 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w6375_,
		_w7038_,
		_w7051_
	);
	LUT4 #(
		.INIT('h3020)
	) name5702 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w6375_,
		_w6378_,
		_w7038_,
		_w7052_
	);
	LUT4 #(
		.INIT('h070f)
	) name5703 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w6380_,
		_w7053_
	);
	LUT3 #(
		.INIT('h2a)
	) name5704 (
		_w2310_,
		_w6380_,
		_w6360_,
		_w7054_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5705 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7055_
	);
	LUT3 #(
		.INIT('hb0)
	) name5706 (
		_w7053_,
		_w7054_,
		_w7055_,
		_w7056_
	);
	LUT2 #(
		.INIT('h4)
	) name5707 (
		_w7052_,
		_w7056_,
		_w7057_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5708 (
		_w1933_,
		_w7048_,
		_w7050_,
		_w7057_,
		_w7058_
	);
	LUT3 #(
		.INIT('h08)
	) name5709 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7059_
	);
	LUT3 #(
		.INIT('h95)
	) name5710 (
		_w3277_,
		_w3136_,
		_w3141_,
		_w7060_
	);
	LUT3 #(
		.INIT('h82)
	) name5711 (
		_w3101_,
		_w4455_,
		_w7060_,
		_w7061_
	);
	LUT3 #(
		.INIT('h87)
	) name5712 (
		_w3136_,
		_w3141_,
		_w3142_,
		_w7062_
	);
	LUT4 #(
		.INIT('h5445)
	) name5713 (
		_w1916_,
		_w3101_,
		_w3202_,
		_w7062_,
		_w7063_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5714 (
		_w1810_,
		_w7059_,
		_w7061_,
		_w7063_,
		_w7064_
	);
	LUT2 #(
		.INIT('h4)
	) name5715 (
		_w1862_,
		_w3277_,
		_w7065_
	);
	LUT4 #(
		.INIT('h00ec)
	) name5716 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w3061_,
		_w7066_
	);
	LUT2 #(
		.INIT('h1)
	) name5717 (
		_w1913_,
		_w7066_,
		_w7067_
	);
	LUT3 #(
		.INIT('h8a)
	) name5718 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1868_,
		_w7067_,
		_w7068_
	);
	LUT3 #(
		.INIT('hb0)
	) name5719 (
		_w1816_,
		_w1831_,
		_w3142_,
		_w7069_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name5720 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		_w1842_,
		_w1845_,
		_w3326_,
		_w7070_
	);
	LUT2 #(
		.INIT('h4)
	) name5721 (
		_w1833_,
		_w7070_,
		_w7071_
	);
	LUT3 #(
		.INIT('h87)
	) name5722 (
		_w3136_,
		_w3141_,
		_w3329_,
		_w7072_
	);
	LUT4 #(
		.INIT('h8f00)
	) name5723 (
		_w3335_,
		_w3338_,
		_w3341_,
		_w7072_,
		_w7073_
	);
	LUT4 #(
		.INIT('h0070)
	) name5724 (
		_w3335_,
		_w3338_,
		_w3341_,
		_w7072_,
		_w7074_
	);
	LUT3 #(
		.INIT('h02)
	) name5725 (
		_w1924_,
		_w7074_,
		_w7073_,
		_w7075_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		_w7071_,
		_w7075_,
		_w7076_
	);
	LUT4 #(
		.INIT('h0100)
	) name5727 (
		_w7068_,
		_w7065_,
		_w7069_,
		_w7076_,
		_w7077_
	);
	LUT2 #(
		.INIT('h8)
	) name5728 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w3406_,
		_w7078_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5729 (
		\P1_InstAddrPointer_reg[4]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w3406_,
		_w3408_,
		_w7079_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5730 (
		_w1933_,
		_w7064_,
		_w7077_,
		_w7079_,
		_w7080_
	);
	LUT3 #(
		.INIT('h87)
	) name5731 (
		_w3121_,
		_w3126_,
		_w3128_,
		_w7081_
	);
	LUT4 #(
		.INIT('hba45)
	) name5732 (
		_w3116_,
		_w3203_,
		_w3206_,
		_w7081_,
		_w7082_
	);
	LUT3 #(
		.INIT('h95)
	) name5733 (
		_w3286_,
		_w3121_,
		_w3126_,
		_w7083_
	);
	LUT3 #(
		.INIT('h70)
	) name5734 (
		_w4456_,
		_w4455_,
		_w4459_,
		_w7084_
	);
	LUT4 #(
		.INIT('he44e)
	) name5735 (
		_w3101_,
		_w7082_,
		_w7083_,
		_w7084_,
		_w7085_
	);
	LUT2 #(
		.INIT('h8)
	) name5736 (
		_w1923_,
		_w7085_,
		_w7086_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5737 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		_w1914_,
		_w1917_,
		_w1868_,
		_w7087_
	);
	LUT3 #(
		.INIT('h87)
	) name5738 (
		_w3121_,
		_w3126_,
		_w3350_,
		_w7088_
	);
	LUT4 #(
		.INIT('h208a)
	) name5739 (
		_w1924_,
		_w3343_,
		_w3346_,
		_w7088_,
		_w7089_
	);
	LUT2 #(
		.INIT('h4)
	) name5740 (
		_w1862_,
		_w3286_,
		_w7090_
	);
	LUT3 #(
		.INIT('h40)
	) name5741 (
		_w1833_,
		_w1846_,
		_w3350_,
		_w7091_
	);
	LUT4 #(
		.INIT('h004f)
	) name5742 (
		_w1816_,
		_w1831_,
		_w3128_,
		_w7091_,
		_w7092_
	);
	LUT4 #(
		.INIT('h0100)
	) name5743 (
		_w7090_,
		_w7087_,
		_w7089_,
		_w7092_,
		_w7093_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5744 (
		\P1_InstAddrPointer_reg[6]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w3406_,
		_w3408_,
		_w7094_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5745 (
		_w1933_,
		_w7086_,
		_w7093_,
		_w7094_,
		_w7095_
	);
	LUT3 #(
		.INIT('h95)
	) name5746 (
		_w2932_,
		_w2836_,
		_w2841_,
		_w7096_
	);
	LUT4 #(
		.INIT('h208a)
	) name5747 (
		_w2180_,
		_w4047_,
		_w4048_,
		_w7096_,
		_w7097_
	);
	LUT4 #(
		.INIT('he000)
	) name5748 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2994_,
		_w7098_
	);
	LUT2 #(
		.INIT('h1)
	) name5749 (
		_w7097_,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h4)
	) name5750 (
		_w2117_,
		_w2932_,
		_w7100_
	);
	LUT3 #(
		.INIT('hb0)
	) name5751 (
		_w2073_,
		_w2086_,
		_w2843_,
		_w7101_
	);
	LUT3 #(
		.INIT('h10)
	) name5752 (
		_w7100_,
		_w7101_,
		_w7099_,
		_w7102_
	);
	LUT4 #(
		.INIT('h0002)
	) name5753 (
		_w2126_,
		_w2174_,
		_w2127_,
		_w2175_,
		_w7103_
	);
	LUT3 #(
		.INIT('h87)
	) name5754 (
		_w2836_,
		_w2841_,
		_w2994_,
		_w7104_
	);
	LUT4 #(
		.INIT('h208a)
	) name5755 (
		_w2181_,
		_w4084_,
		_w4085_,
		_w7104_,
		_w7105_
	);
	LUT3 #(
		.INIT('h0d)
	) name5756 (
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		_w7103_,
		_w7105_,
		_w7106_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5757 (
		\P3_InstAddrPointer_reg[6]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w3054_,
		_w3056_,
		_w7107_
	);
	LUT4 #(
		.INIT('h2aff)
	) name5758 (
		_w1945_,
		_w7102_,
		_w7106_,
		_w7107_,
		_w7108_
	);
	LUT3 #(
		.INIT('h08)
	) name5759 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7109_
	);
	LUT3 #(
		.INIT('h87)
	) name5760 (
		_w4147_,
		_w4152_,
		_w4154_,
		_w7110_
	);
	LUT4 #(
		.INIT('hb04f)
	) name5761 (
		_w4141_,
		_w4169_,
		_w4801_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h2)
	) name5762 (
		_w4214_,
		_w7111_,
		_w7112_
	);
	LUT3 #(
		.INIT('h95)
	) name5763 (
		_w4298_,
		_w4147_,
		_w4152_,
		_w7113_
	);
	LUT4 #(
		.INIT('h5445)
	) name5764 (
		_w1661_,
		_w4214_,
		_w4814_,
		_w7113_,
		_w7114_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5765 (
		_w1559_,
		_w7109_,
		_w7112_,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h8)
	) name5766 (
		_w1640_,
		_w4382_,
		_w7116_
	);
	LUT4 #(
		.INIT('h00d5)
	) name5767 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		_w1658_,
		_w4844_,
		_w7116_,
		_w7117_
	);
	LUT2 #(
		.INIT('h4)
	) name5768 (
		_w1617_,
		_w4154_,
		_w7118_
	);
	LUT3 #(
		.INIT('h87)
	) name5769 (
		_w4147_,
		_w4152_,
		_w4382_,
		_w7119_
	);
	LUT4 #(
		.INIT('h5501)
	) name5770 (
		_w4385_,
		_w4387_,
		_w4391_,
		_w4393_,
		_w7120_
	);
	LUT3 #(
		.INIT('h28)
	) name5771 (
		_w1659_,
		_w7119_,
		_w7120_,
		_w7121_
	);
	LUT4 #(
		.INIT('h004f)
	) name5772 (
		_w1571_,
		_w1583_,
		_w4298_,
		_w7121_,
		_w7122_
	);
	LUT4 #(
		.INIT('h1000)
	) name5773 (
		_w7118_,
		_w7115_,
		_w7117_,
		_w7122_,
		_w7123_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5774 (
		\P2_InstAddrPointer_reg[4]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w2286_,
		_w4441_,
		_w7124_
	);
	LUT3 #(
		.INIT('h2f)
	) name5775 (
		_w1678_,
		_w7123_,
		_w7124_,
		_w7125_
	);
	LUT3 #(
		.INIT('h08)
	) name5776 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7126_
	);
	LUT3 #(
		.INIT('h95)
	) name5777 (
		_w4285_,
		_w4178_,
		_w4183_,
		_w7127_
	);
	LUT4 #(
		.INIT('hba45)
	) name5778 (
		_w4288_,
		_w4815_,
		_w4816_,
		_w7127_,
		_w7128_
	);
	LUT3 #(
		.INIT('h87)
	) name5779 (
		_w4178_,
		_w4183_,
		_w4186_,
		_w7129_
	);
	LUT4 #(
		.INIT('h8a20)
	) name5780 (
		_w4214_,
		_w4803_,
		_w4804_,
		_w7129_,
		_w7130_
	);
	LUT4 #(
		.INIT('h0504)
	) name5781 (
		_w1661_,
		_w4214_,
		_w7130_,
		_w7128_,
		_w7131_
	);
	LUT3 #(
		.INIT('ha8)
	) name5782 (
		_w1559_,
		_w7126_,
		_w7131_,
		_w7132_
	);
	LUT3 #(
		.INIT('h87)
	) name5783 (
		_w4178_,
		_w4183_,
		_w4377_,
		_w7133_
	);
	LUT3 #(
		.INIT('h45)
	) name5784 (
		_w4380_,
		_w4866_,
		_w4867_,
		_w7134_
	);
	LUT4 #(
		.INIT('h4500)
	) name5785 (
		_w4380_,
		_w4866_,
		_w4867_,
		_w7133_,
		_w7135_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5786 (
		_w4380_,
		_w4866_,
		_w4867_,
		_w7133_,
		_w7136_
	);
	LUT3 #(
		.INIT('h02)
	) name5787 (
		_w1659_,
		_w7136_,
		_w7135_,
		_w7137_
	);
	LUT2 #(
		.INIT('h8)
	) name5788 (
		_w1640_,
		_w4377_,
		_w7138_
	);
	LUT4 #(
		.INIT('h004f)
	) name5789 (
		_w1571_,
		_w1583_,
		_w4285_,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h4)
	) name5790 (
		_w1617_,
		_w4186_,
		_w7140_
	);
	LUT3 #(
		.INIT('h2a)
	) name5791 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		_w1658_,
		_w4844_,
		_w7141_
	);
	LUT4 #(
		.INIT('h0100)
	) name5792 (
		_w7140_,
		_w7141_,
		_w7137_,
		_w7139_,
		_w7142_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5793 (
		\P2_InstAddrPointer_reg[6]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w2286_,
		_w4441_,
		_w7143_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5794 (
		_w1678_,
		_w7132_,
		_w7142_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('hc444)
	) name5795 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7145_
	);
	LUT4 #(
		.INIT('h0888)
	) name5796 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[25]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7146_
	);
	LUT2 #(
		.INIT('h1)
	) name5797 (
		_w7145_,
		_w7146_,
		_w7147_
	);
	LUT3 #(
		.INIT('ha8)
	) name5798 (
		_w2250_,
		_w7145_,
		_w7146_,
		_w7148_
	);
	LUT4 #(
		.INIT('hc444)
	) name5799 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[17]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7149_
	);
	LUT4 #(
		.INIT('h0888)
	) name5800 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[17]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7150_
	);
	LUT2 #(
		.INIT('h1)
	) name5801 (
		_w7149_,
		_w7150_,
		_w7151_
	);
	LUT3 #(
		.INIT('ha8)
	) name5802 (
		_w2264_,
		_w7149_,
		_w7150_,
		_w7152_
	);
	LUT3 #(
		.INIT('ha8)
	) name5803 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7148_,
		_w7152_,
		_w7153_
	);
	LUT4 #(
		.INIT('hc444)
	) name5804 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7154_
	);
	LUT4 #(
		.INIT('h0888)
	) name5805 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[1]/NET0131 ,
		_w2255_,
		_w2260_,
		_w7155_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w7154_,
		_w7155_,
		_w7156_
	);
	LUT3 #(
		.INIT('h02)
	) name5807 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w2271_,
		_w2272_,
		_w7157_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5808 (
		_w2273_,
		_w7154_,
		_w7155_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h1)
	) name5809 (
		_w2280_,
		_w7158_,
		_w7159_
	);
	LUT3 #(
		.INIT('ha8)
	) name5810 (
		_w1679_,
		_w7153_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h2)
	) name5811 (
		_w2283_,
		_w7158_,
		_w7161_
	);
	LUT4 #(
		.INIT('hc055)
	) name5812 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2272_,
		_w7162_
	);
	LUT2 #(
		.INIT('h2)
	) name5813 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		_w2288_,
		_w7163_
	);
	LUT3 #(
		.INIT('h0d)
	) name5814 (
		_w2246_,
		_w7162_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h4)
	) name5815 (
		_w7161_,
		_w7164_,
		_w7165_
	);
	LUT2 #(
		.INIT('hb)
	) name5816 (
		_w7160_,
		_w7165_,
		_w7166_
	);
	LUT3 #(
		.INIT('ha8)
	) name5817 (
		_w2315_,
		_w7145_,
		_w7146_,
		_w7167_
	);
	LUT3 #(
		.INIT('ha8)
	) name5818 (
		_w2317_,
		_w7149_,
		_w7150_,
		_w7168_
	);
	LUT3 #(
		.INIT('ha8)
	) name5819 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7167_,
		_w7168_,
		_w7169_
	);
	LUT3 #(
		.INIT('h02)
	) name5820 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w2320_,
		_w2322_,
		_w7170_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5821 (
		_w2323_,
		_w7154_,
		_w7155_,
		_w7170_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name5822 (
		_w2327_,
		_w7171_,
		_w7172_
	);
	LUT3 #(
		.INIT('ha8)
	) name5823 (
		_w1679_,
		_w7169_,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h2)
	) name5824 (
		_w2283_,
		_w7171_,
		_w7174_
	);
	LUT4 #(
		.INIT('hc055)
	) name5825 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2320_,
		_w7175_
	);
	LUT2 #(
		.INIT('h2)
	) name5826 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		_w2288_,
		_w7176_
	);
	LUT3 #(
		.INIT('h0d)
	) name5827 (
		_w2246_,
		_w7175_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h4)
	) name5828 (
		_w7174_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('hb)
	) name5829 (
		_w7173_,
		_w7178_,
		_w7179_
	);
	LUT3 #(
		.INIT('ha8)
	) name5830 (
		_w2250_,
		_w7149_,
		_w7150_,
		_w7180_
	);
	LUT3 #(
		.INIT('ha8)
	) name5831 (
		_w2349_,
		_w7145_,
		_w7146_,
		_w7181_
	);
	LUT3 #(
		.INIT('ha8)
	) name5832 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7180_,
		_w7181_,
		_w7182_
	);
	LUT3 #(
		.INIT('h02)
	) name5833 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w2271_,
		_w2264_,
		_w7183_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5834 (
		_w2346_,
		_w7154_,
		_w7155_,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h1)
	) name5835 (
		_w2351_,
		_w7184_,
		_w7185_
	);
	LUT3 #(
		.INIT('ha8)
	) name5836 (
		_w1679_,
		_w7182_,
		_w7185_,
		_w7186_
	);
	LUT2 #(
		.INIT('h2)
	) name5837 (
		_w2283_,
		_w7184_,
		_w7187_
	);
	LUT4 #(
		.INIT('hc055)
	) name5838 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2271_,
		_w7188_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		_w2288_,
		_w7189_
	);
	LUT3 #(
		.INIT('h0d)
	) name5840 (
		_w2246_,
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h4)
	) name5841 (
		_w7187_,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('hb)
	) name5842 (
		_w7186_,
		_w7191_,
		_w7192_
	);
	LUT3 #(
		.INIT('ha8)
	) name5843 (
		_w2264_,
		_w7145_,
		_w7146_,
		_w7193_
	);
	LUT3 #(
		.INIT('ha8)
	) name5844 (
		_w2271_,
		_w7149_,
		_w7150_,
		_w7194_
	);
	LUT3 #(
		.INIT('ha8)
	) name5845 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7193_,
		_w7194_,
		_w7195_
	);
	LUT3 #(
		.INIT('h02)
	) name5846 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w2272_,
		_w2376_,
		_w7196_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5847 (
		_w2377_,
		_w7154_,
		_w7155_,
		_w7196_,
		_w7197_
	);
	LUT2 #(
		.INIT('h1)
	) name5848 (
		_w2380_,
		_w7197_,
		_w7198_
	);
	LUT3 #(
		.INIT('ha8)
	) name5849 (
		_w1679_,
		_w7195_,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h2)
	) name5850 (
		_w2283_,
		_w7197_,
		_w7200_
	);
	LUT4 #(
		.INIT('hc055)
	) name5851 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2376_,
		_w7201_
	);
	LUT2 #(
		.INIT('h2)
	) name5852 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		_w2288_,
		_w7202_
	);
	LUT3 #(
		.INIT('h0d)
	) name5853 (
		_w2246_,
		_w7201_,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h4)
	) name5854 (
		_w7200_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('hb)
	) name5855 (
		_w7199_,
		_w7204_,
		_w7205_
	);
	LUT3 #(
		.INIT('ha8)
	) name5856 (
		_w2271_,
		_w7145_,
		_w7146_,
		_w7206_
	);
	LUT3 #(
		.INIT('ha8)
	) name5857 (
		_w2272_,
		_w7149_,
		_w7150_,
		_w7207_
	);
	LUT3 #(
		.INIT('ha8)
	) name5858 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7206_,
		_w7207_,
		_w7208_
	);
	LUT3 #(
		.INIT('h02)
	) name5859 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w2315_,
		_w2376_,
		_w7209_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5860 (
		_w2402_,
		_w7154_,
		_w7155_,
		_w7209_,
		_w7210_
	);
	LUT2 #(
		.INIT('h1)
	) name5861 (
		_w2405_,
		_w7210_,
		_w7211_
	);
	LUT3 #(
		.INIT('ha8)
	) name5862 (
		_w1679_,
		_w7208_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h2)
	) name5863 (
		_w2283_,
		_w7210_,
		_w7213_
	);
	LUT4 #(
		.INIT('hc055)
	) name5864 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2315_,
		_w7214_
	);
	LUT2 #(
		.INIT('h2)
	) name5865 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		_w2288_,
		_w7215_
	);
	LUT3 #(
		.INIT('h0d)
	) name5866 (
		_w2246_,
		_w7214_,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('h4)
	) name5867 (
		_w7213_,
		_w7216_,
		_w7217_
	);
	LUT2 #(
		.INIT('hb)
	) name5868 (
		_w7212_,
		_w7217_,
		_w7218_
	);
	LUT3 #(
		.INIT('ha8)
	) name5869 (
		_w2272_,
		_w7145_,
		_w7146_,
		_w7219_
	);
	LUT3 #(
		.INIT('ha8)
	) name5870 (
		_w2376_,
		_w7149_,
		_w7150_,
		_w7220_
	);
	LUT3 #(
		.INIT('ha8)
	) name5871 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT3 #(
		.INIT('h02)
	) name5872 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w2315_,
		_w2317_,
		_w7222_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5873 (
		_w2326_,
		_w7154_,
		_w7155_,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name5874 (
		_w2429_,
		_w7223_,
		_w7224_
	);
	LUT3 #(
		.INIT('ha8)
	) name5875 (
		_w1679_,
		_w7221_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h2)
	) name5876 (
		_w2283_,
		_w7223_,
		_w7226_
	);
	LUT4 #(
		.INIT('hc055)
	) name5877 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2317_,
		_w7227_
	);
	LUT2 #(
		.INIT('h2)
	) name5878 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w2288_,
		_w7228_
	);
	LUT3 #(
		.INIT('h0d)
	) name5879 (
		_w2246_,
		_w7227_,
		_w7228_,
		_w7229_
	);
	LUT2 #(
		.INIT('h4)
	) name5880 (
		_w7226_,
		_w7229_,
		_w7230_
	);
	LUT2 #(
		.INIT('hb)
	) name5881 (
		_w7225_,
		_w7230_,
		_w7231_
	);
	LUT3 #(
		.INIT('ha8)
	) name5882 (
		_w2376_,
		_w7145_,
		_w7146_,
		_w7232_
	);
	LUT3 #(
		.INIT('ha8)
	) name5883 (
		_w2315_,
		_w7149_,
		_w7150_,
		_w7233_
	);
	LUT3 #(
		.INIT('ha8)
	) name5884 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7232_,
		_w7233_,
		_w7234_
	);
	LUT3 #(
		.INIT('h02)
	) name5885 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w2322_,
		_w2317_,
		_w7235_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5886 (
		_w2451_,
		_w7154_,
		_w7155_,
		_w7235_,
		_w7236_
	);
	LUT2 #(
		.INIT('h1)
	) name5887 (
		_w2454_,
		_w7236_,
		_w7237_
	);
	LUT3 #(
		.INIT('ha8)
	) name5888 (
		_w1679_,
		_w7234_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h2)
	) name5889 (
		_w2283_,
		_w7236_,
		_w7239_
	);
	LUT4 #(
		.INIT('hc055)
	) name5890 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2322_,
		_w7240_
	);
	LUT2 #(
		.INIT('h2)
	) name5891 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w2288_,
		_w7241_
	);
	LUT3 #(
		.INIT('h0d)
	) name5892 (
		_w2246_,
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT2 #(
		.INIT('h4)
	) name5893 (
		_w7239_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('hb)
	) name5894 (
		_w7238_,
		_w7243_,
		_w7244_
	);
	LUT3 #(
		.INIT('ha8)
	) name5895 (
		_w2317_,
		_w7145_,
		_w7146_,
		_w7245_
	);
	LUT3 #(
		.INIT('ha8)
	) name5896 (
		_w2322_,
		_w7149_,
		_w7150_,
		_w7246_
	);
	LUT3 #(
		.INIT('ha8)
	) name5897 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7245_,
		_w7246_,
		_w7247_
	);
	LUT3 #(
		.INIT('h02)
	) name5898 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w2320_,
		_w2473_,
		_w7248_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5899 (
		_w2474_,
		_w7154_,
		_w7155_,
		_w7248_,
		_w7249_
	);
	LUT2 #(
		.INIT('h1)
	) name5900 (
		_w2477_,
		_w7249_,
		_w7250_
	);
	LUT3 #(
		.INIT('ha8)
	) name5901 (
		_w1679_,
		_w7247_,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('h2)
	) name5902 (
		_w2283_,
		_w7249_,
		_w7252_
	);
	LUT4 #(
		.INIT('hc055)
	) name5903 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2473_,
		_w7253_
	);
	LUT2 #(
		.INIT('h2)
	) name5904 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w2288_,
		_w7254_
	);
	LUT3 #(
		.INIT('h0d)
	) name5905 (
		_w2246_,
		_w7253_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h4)
	) name5906 (
		_w7252_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('hb)
	) name5907 (
		_w7251_,
		_w7256_,
		_w7257_
	);
	LUT3 #(
		.INIT('ha8)
	) name5908 (
		_w2320_,
		_w7149_,
		_w7150_,
		_w7258_
	);
	LUT3 #(
		.INIT('ha8)
	) name5909 (
		_w2322_,
		_w7145_,
		_w7146_,
		_w7259_
	);
	LUT3 #(
		.INIT('ha8)
	) name5910 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7258_,
		_w7259_,
		_w7260_
	);
	LUT3 #(
		.INIT('h02)
	) name5911 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w2473_,
		_w2502_,
		_w7261_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5912 (
		_w2503_,
		_w7154_,
		_w7155_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h1)
	) name5913 (
		_w2506_,
		_w7262_,
		_w7263_
	);
	LUT3 #(
		.INIT('ha8)
	) name5914 (
		_w1679_,
		_w7260_,
		_w7263_,
		_w7264_
	);
	LUT2 #(
		.INIT('h2)
	) name5915 (
		_w2283_,
		_w7262_,
		_w7265_
	);
	LUT4 #(
		.INIT('hc055)
	) name5916 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2502_,
		_w7266_
	);
	LUT2 #(
		.INIT('h2)
	) name5917 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w2288_,
		_w7267_
	);
	LUT3 #(
		.INIT('h0d)
	) name5918 (
		_w2246_,
		_w7266_,
		_w7267_,
		_w7268_
	);
	LUT2 #(
		.INIT('h4)
	) name5919 (
		_w7265_,
		_w7268_,
		_w7269_
	);
	LUT2 #(
		.INIT('hb)
	) name5920 (
		_w7264_,
		_w7269_,
		_w7270_
	);
	LUT3 #(
		.INIT('ha8)
	) name5921 (
		_w2320_,
		_w7145_,
		_w7146_,
		_w7271_
	);
	LUT3 #(
		.INIT('ha8)
	) name5922 (
		_w2473_,
		_w7149_,
		_w7150_,
		_w7272_
	);
	LUT3 #(
		.INIT('ha8)
	) name5923 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7271_,
		_w7272_,
		_w7273_
	);
	LUT3 #(
		.INIT('h02)
	) name5924 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w2502_,
		_w2528_,
		_w7274_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5925 (
		_w2529_,
		_w7154_,
		_w7155_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w2532_,
		_w7275_,
		_w7276_
	);
	LUT3 #(
		.INIT('ha8)
	) name5927 (
		_w1679_,
		_w7273_,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('h2)
	) name5928 (
		_w2283_,
		_w7275_,
		_w7278_
	);
	LUT4 #(
		.INIT('hc055)
	) name5929 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2528_,
		_w7279_
	);
	LUT2 #(
		.INIT('h2)
	) name5930 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w2288_,
		_w7280_
	);
	LUT3 #(
		.INIT('h0d)
	) name5931 (
		_w2246_,
		_w7279_,
		_w7280_,
		_w7281_
	);
	LUT2 #(
		.INIT('h4)
	) name5932 (
		_w7278_,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('hb)
	) name5933 (
		_w7277_,
		_w7282_,
		_w7283_
	);
	LUT3 #(
		.INIT('ha8)
	) name5934 (
		_w2473_,
		_w7145_,
		_w7146_,
		_w7284_
	);
	LUT3 #(
		.INIT('ha8)
	) name5935 (
		_w2502_,
		_w7149_,
		_w7150_,
		_w7285_
	);
	LUT3 #(
		.INIT('ha8)
	) name5936 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT3 #(
		.INIT('h02)
	) name5937 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w2528_,
		_w2554_,
		_w7287_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5938 (
		_w2555_,
		_w7154_,
		_w7155_,
		_w7287_,
		_w7288_
	);
	LUT2 #(
		.INIT('h1)
	) name5939 (
		_w2558_,
		_w7288_,
		_w7289_
	);
	LUT3 #(
		.INIT('ha8)
	) name5940 (
		_w1679_,
		_w7286_,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h2)
	) name5941 (
		_w2283_,
		_w7288_,
		_w7291_
	);
	LUT4 #(
		.INIT('hc055)
	) name5942 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2554_,
		_w7292_
	);
	LUT2 #(
		.INIT('h2)
	) name5943 (
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w2288_,
		_w7293_
	);
	LUT3 #(
		.INIT('h0d)
	) name5944 (
		_w2246_,
		_w7292_,
		_w7293_,
		_w7294_
	);
	LUT2 #(
		.INIT('h4)
	) name5945 (
		_w7291_,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('hb)
	) name5946 (
		_w7290_,
		_w7295_,
		_w7296_
	);
	LUT3 #(
		.INIT('ha8)
	) name5947 (
		_w2502_,
		_w7145_,
		_w7146_,
		_w7297_
	);
	LUT3 #(
		.INIT('ha8)
	) name5948 (
		_w2528_,
		_w7149_,
		_w7150_,
		_w7298_
	);
	LUT3 #(
		.INIT('ha8)
	) name5949 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7297_,
		_w7298_,
		_w7299_
	);
	LUT3 #(
		.INIT('h02)
	) name5950 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w2554_,
		_w2580_,
		_w7300_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5951 (
		_w2581_,
		_w7154_,
		_w7155_,
		_w7300_,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name5952 (
		_w2584_,
		_w7301_,
		_w7302_
	);
	LUT3 #(
		.INIT('ha8)
	) name5953 (
		_w1679_,
		_w7299_,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h2)
	) name5954 (
		_w2283_,
		_w7301_,
		_w7304_
	);
	LUT4 #(
		.INIT('hc055)
	) name5955 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2580_,
		_w7305_
	);
	LUT2 #(
		.INIT('h2)
	) name5956 (
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w2288_,
		_w7306_
	);
	LUT3 #(
		.INIT('h0d)
	) name5957 (
		_w2246_,
		_w7305_,
		_w7306_,
		_w7307_
	);
	LUT2 #(
		.INIT('h4)
	) name5958 (
		_w7304_,
		_w7307_,
		_w7308_
	);
	LUT2 #(
		.INIT('hb)
	) name5959 (
		_w7303_,
		_w7308_,
		_w7309_
	);
	LUT3 #(
		.INIT('ha8)
	) name5960 (
		_w2528_,
		_w7145_,
		_w7146_,
		_w7310_
	);
	LUT3 #(
		.INIT('ha8)
	) name5961 (
		_w2554_,
		_w7149_,
		_w7150_,
		_w7311_
	);
	LUT3 #(
		.INIT('ha8)
	) name5962 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7310_,
		_w7311_,
		_w7312_
	);
	LUT3 #(
		.INIT('h02)
	) name5963 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w2580_,
		_w2606_,
		_w7313_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5964 (
		_w2607_,
		_w7154_,
		_w7155_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h1)
	) name5965 (
		_w2610_,
		_w7314_,
		_w7315_
	);
	LUT3 #(
		.INIT('ha8)
	) name5966 (
		_w1679_,
		_w7312_,
		_w7315_,
		_w7316_
	);
	LUT2 #(
		.INIT('h2)
	) name5967 (
		_w2283_,
		_w7314_,
		_w7317_
	);
	LUT4 #(
		.INIT('hc055)
	) name5968 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2606_,
		_w7318_
	);
	LUT2 #(
		.INIT('h2)
	) name5969 (
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w2288_,
		_w7319_
	);
	LUT3 #(
		.INIT('h0d)
	) name5970 (
		_w2246_,
		_w7318_,
		_w7319_,
		_w7320_
	);
	LUT2 #(
		.INIT('h4)
	) name5971 (
		_w7317_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('hb)
	) name5972 (
		_w7316_,
		_w7321_,
		_w7322_
	);
	LUT3 #(
		.INIT('ha8)
	) name5973 (
		_w2554_,
		_w7145_,
		_w7146_,
		_w7323_
	);
	LUT3 #(
		.INIT('ha8)
	) name5974 (
		_w2580_,
		_w7149_,
		_w7150_,
		_w7324_
	);
	LUT3 #(
		.INIT('ha8)
	) name5975 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7323_,
		_w7324_,
		_w7325_
	);
	LUT3 #(
		.INIT('h02)
	) name5976 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w2349_,
		_w2606_,
		_w7326_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5977 (
		_w2632_,
		_w7154_,
		_w7155_,
		_w7326_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name5978 (
		_w2635_,
		_w7327_,
		_w7328_
	);
	LUT3 #(
		.INIT('ha8)
	) name5979 (
		_w1679_,
		_w7325_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h2)
	) name5980 (
		_w2283_,
		_w7327_,
		_w7330_
	);
	LUT4 #(
		.INIT('hc055)
	) name5981 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2349_,
		_w7331_
	);
	LUT2 #(
		.INIT('h2)
	) name5982 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w2288_,
		_w7332_
	);
	LUT3 #(
		.INIT('h0d)
	) name5983 (
		_w2246_,
		_w7331_,
		_w7332_,
		_w7333_
	);
	LUT2 #(
		.INIT('h4)
	) name5984 (
		_w7330_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('hb)
	) name5985 (
		_w7329_,
		_w7334_,
		_w7335_
	);
	LUT3 #(
		.INIT('ha8)
	) name5986 (
		_w2580_,
		_w7145_,
		_w7146_,
		_w7336_
	);
	LUT3 #(
		.INIT('ha8)
	) name5987 (
		_w2606_,
		_w7149_,
		_w7150_,
		_w7337_
	);
	LUT3 #(
		.INIT('ha8)
	) name5988 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT3 #(
		.INIT('h02)
	) name5989 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w2250_,
		_w2349_,
		_w7339_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5990 (
		_w2350_,
		_w7154_,
		_w7155_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w2659_,
		_w7340_,
		_w7341_
	);
	LUT3 #(
		.INIT('ha8)
	) name5992 (
		_w1679_,
		_w7338_,
		_w7341_,
		_w7342_
	);
	LUT2 #(
		.INIT('h2)
	) name5993 (
		_w2283_,
		_w7340_,
		_w7343_
	);
	LUT4 #(
		.INIT('hc055)
	) name5994 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2250_,
		_w7344_
	);
	LUT2 #(
		.INIT('h2)
	) name5995 (
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w2288_,
		_w7345_
	);
	LUT3 #(
		.INIT('h0d)
	) name5996 (
		_w2246_,
		_w7344_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h4)
	) name5997 (
		_w7343_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('hb)
	) name5998 (
		_w7342_,
		_w7347_,
		_w7348_
	);
	LUT3 #(
		.INIT('ha8)
	) name5999 (
		_w2606_,
		_w7145_,
		_w7146_,
		_w7349_
	);
	LUT3 #(
		.INIT('ha8)
	) name6000 (
		_w2349_,
		_w7149_,
		_w7150_,
		_w7350_
	);
	LUT3 #(
		.INIT('ha8)
	) name6001 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7349_,
		_w7350_,
		_w7351_
	);
	LUT3 #(
		.INIT('h02)
	) name6002 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w2250_,
		_w2264_,
		_w7352_
	);
	LUT4 #(
		.INIT('h00ab)
	) name6003 (
		_w2279_,
		_w7154_,
		_w7155_,
		_w7352_,
		_w7353_
	);
	LUT2 #(
		.INIT('h1)
	) name6004 (
		_w2683_,
		_w7353_,
		_w7354_
	);
	LUT3 #(
		.INIT('ha8)
	) name6005 (
		_w1679_,
		_w7351_,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('h2)
	) name6006 (
		_w2283_,
		_w7353_,
		_w7356_
	);
	LUT4 #(
		.INIT('hc055)
	) name6007 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1495_,
		_w1500_,
		_w2264_,
		_w7357_
	);
	LUT2 #(
		.INIT('h2)
	) name6008 (
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w2288_,
		_w7358_
	);
	LUT3 #(
		.INIT('h0d)
	) name6009 (
		_w2246_,
		_w7357_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h4)
	) name6010 (
		_w7356_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('hb)
	) name6011 (
		_w7355_,
		_w7360_,
		_w7361_
	);
	LUT3 #(
		.INIT('h08)
	) name6012 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7362_
	);
	LUT2 #(
		.INIT('h2)
	) name6013 (
		_w4345_,
		_w6885_,
		_w7363_
	);
	LUT3 #(
		.INIT('h15)
	) name6014 (
		_w4214_,
		_w4348_,
		_w4855_,
		_w7364_
	);
	LUT4 #(
		.INIT('h4555)
	) name6015 (
		_w4256_,
		_w4807_,
		_w4810_,
		_w4859_,
		_w7365_
	);
	LUT4 #(
		.INIT('h1115)
	) name6016 (
		_w1661_,
		_w4214_,
		_w4259_,
		_w7365_,
		_w7366_
	);
	LUT4 #(
		.INIT('h1055)
	) name6017 (
		_w7362_,
		_w7363_,
		_w7364_,
		_w7366_,
		_w7367_
	);
	LUT4 #(
		.INIT('h028a)
	) name6018 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7368_
	);
	LUT4 #(
		.INIT('h007f)
	) name6019 (
		_w4414_,
		_w6897_,
		_w6898_,
		_w6899_,
		_w7369_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6020 (
		_w1659_,
		_w4415_,
		_w6897_,
		_w6898_,
		_w7370_
	);
	LUT3 #(
		.INIT('h45)
	) name6021 (
		_w7368_,
		_w7369_,
		_w7370_,
		_w7371_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6022 (
		_w1559_,
		_w1678_,
		_w7367_,
		_w7371_,
		_w7372_
	);
	LUT3 #(
		.INIT('h6c)
	) name6023 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w7373_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6024 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w5746_,
		_w7374_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6025 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7375_
	);
	LUT4 #(
		.INIT('hb700)
	) name6026 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w2242_,
		_w5733_,
		_w7375_,
		_w7376_
	);
	LUT2 #(
		.INIT('h4)
	) name6027 (
		_w7374_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('hb)
	) name6028 (
		_w7372_,
		_w7377_,
		_w7378_
	);
	LUT3 #(
		.INIT('h08)
	) name6029 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7379_
	);
	LUT4 #(
		.INIT('h004f)
	) name6030 (
		_w4856_,
		_w4857_,
		_w4863_,
		_w7379_,
		_w7380_
	);
	LUT4 #(
		.INIT('h028a)
	) name6031 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7381_
	);
	LUT3 #(
		.INIT('h0b)
	) name6032 (
		_w4875_,
		_w4877_,
		_w7381_,
		_w7382_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6033 (
		_w1559_,
		_w1678_,
		_w7380_,
		_w7382_,
		_w7383_
	);
	LUT4 #(
		.INIT('h8000)
	) name6034 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w5733_,
		_w7384_
	);
	LUT3 #(
		.INIT('h32)
	) name6035 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w6860_,
		_w7384_,
		_w7385_
	);
	LUT4 #(
		.INIT('h0c08)
	) name6036 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w5746_,
		_w6860_,
		_w7384_,
		_w7386_
	);
	LUT4 #(
		.INIT('h070f)
	) name6037 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		_w5733_,
		_w7387_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6038 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w2242_,
		_w5733_,
		_w5734_,
		_w7388_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6039 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7389_
	);
	LUT3 #(
		.INIT('hb0)
	) name6040 (
		_w7387_,
		_w7388_,
		_w7389_,
		_w7390_
	);
	LUT2 #(
		.INIT('h4)
	) name6041 (
		_w7386_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('hb)
	) name6042 (
		_w7383_,
		_w7391_,
		_w7392_
	);
	LUT3 #(
		.INIT('h08)
	) name6043 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7393_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6044 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w4255_,
		_w4263_,
		_w7394_
	);
	LUT4 #(
		.INIT('h4888)
	) name6045 (
		\P2_InstAddrPointer_reg[22]/NET0131 ,
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w4255_,
		_w4260_,
		_w7395_
	);
	LUT4 #(
		.INIT('h5450)
	) name6046 (
		_w4267_,
		_w4862_,
		_w7394_,
		_w7395_,
		_w7396_
	);
	LUT3 #(
		.INIT('h6a)
	) name6047 (
		_w4356_,
		_w6846_,
		_w6885_,
		_w7397_
	);
	LUT4 #(
		.INIT('h5410)
	) name6048 (
		_w1661_,
		_w4214_,
		_w7397_,
		_w7396_,
		_w7398_
	);
	LUT4 #(
		.INIT('h028a)
	) name6049 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7399_
	);
	LUT4 #(
		.INIT('h8000)
	) name6050 (
		_w4414_,
		_w6897_,
		_w6898_,
		_w6902_,
		_w7400_
	);
	LUT4 #(
		.INIT('h0d07)
	) name6051 (
		_w1659_,
		_w4913_,
		_w7399_,
		_w7400_,
		_w7401_
	);
	LUT4 #(
		.INIT('h5700)
	) name6052 (
		_w1559_,
		_w7393_,
		_w7398_,
		_w7401_,
		_w7402_
	);
	LUT3 #(
		.INIT('h6c)
	) name6053 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5736_,
		_w7403_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6054 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5736_,
		_w5746_,
		_w7404_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6055 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7405_
	);
	LUT4 #(
		.INIT('hb700)
	) name6056 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w2242_,
		_w5736_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h4)
	) name6057 (
		_w7404_,
		_w7406_,
		_w7407_
	);
	LUT3 #(
		.INIT('h2f)
	) name6058 (
		_w1678_,
		_w7402_,
		_w7407_,
		_w7408_
	);
	LUT4 #(
		.INIT('h4447)
	) name6059 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w1661_,
		_w4902_,
		_w4907_,
		_w7409_
	);
	LUT4 #(
		.INIT('h028a)
	) name6060 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7410_
	);
	LUT4 #(
		.INIT('h0031)
	) name6061 (
		_w1559_,
		_w4917_,
		_w7409_,
		_w7410_,
		_w7411_
	);
	LUT4 #(
		.INIT('h1333)
	) name6062 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w5736_,
		_w5742_,
		_w7412_
	);
	LUT3 #(
		.INIT('h07)
	) name6063 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5738_,
		_w7412_,
		_w7413_
	);
	LUT4 #(
		.INIT('h0070)
	) name6064 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5738_,
		_w5746_,
		_w7412_,
		_w7414_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6065 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7415_
	);
	LUT4 #(
		.INIT('hb700)
	) name6066 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		_w2242_,
		_w5737_,
		_w7415_,
		_w7416_
	);
	LUT2 #(
		.INIT('h4)
	) name6067 (
		_w7414_,
		_w7416_,
		_w7417_
	);
	LUT3 #(
		.INIT('h2f)
	) name6068 (
		_w1678_,
		_w7411_,
		_w7417_,
		_w7418_
	);
	LUT3 #(
		.INIT('h80)
	) name6069 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2987_,
		_w6412_,
		_w7419_
	);
	LUT2 #(
		.INIT('h6)
	) name6070 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2986_,
		_w7420_
	);
	LUT4 #(
		.INIT('haa80)
	) name6071 (
		_w2181_,
		_w2987_,
		_w6412_,
		_w7420_,
		_w7421_
	);
	LUT4 #(
		.INIT('h80c4)
	) name6072 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w2173_,
		_w7422_
	);
	LUT2 #(
		.INIT('h2)
	) name6073 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w7422_,
		_w7423_
	);
	LUT4 #(
		.INIT('h8c00)
	) name6074 (
		_w2935_,
		_w2936_,
		_w2940_,
		_w2946_,
		_w7424_
	);
	LUT4 #(
		.INIT('hcf8a)
	) name6075 (
		_w2950_,
		_w4051_,
		_w4054_,
		_w7424_,
		_w7425_
	);
	LUT4 #(
		.INIT('h4554)
	) name6076 (
		_w2173_,
		_w2755_,
		_w2876_,
		_w2874_,
		_w7426_
	);
	LUT4 #(
		.INIT('ha200)
	) name6077 (
		_w2171_,
		_w2755_,
		_w7425_,
		_w7426_,
		_w7427_
	);
	LUT4 #(
		.INIT('h1011)
	) name6078 (
		_w7423_,
		_w7427_,
		_w7419_,
		_w7421_,
		_w7428_
	);
	LUT3 #(
		.INIT('h6a)
	) name6079 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5761_,
		_w7429_
	);
	LUT4 #(
		.INIT('h4111)
	) name6080 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5761_,
		_w7430_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6081 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w7431_
	);
	LUT3 #(
		.INIT('hc4)
	) name6082 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w7431_,
		_w7432_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6083 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w3055_,
		_w5761_,
		_w7433_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6084 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7434_
	);
	LUT4 #(
		.INIT('h4500)
	) name6085 (
		_w7433_,
		_w7430_,
		_w7432_,
		_w7434_,
		_w7435_
	);
	LUT3 #(
		.INIT('h2f)
	) name6086 (
		_w1945_,
		_w7428_,
		_w7435_,
		_w7436_
	);
	LUT3 #(
		.INIT('h02)
	) name6087 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7437_
	);
	LUT3 #(
		.INIT('ha8)
	) name6088 (
		_w2171_,
		_w4755_,
		_w7437_,
		_w7438_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6089 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7439_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		_w4759_,
		_w7439_,
		_w7440_
	);
	LUT4 #(
		.INIT('h8000)
	) name6091 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5762_,
		_w7441_
	);
	LUT3 #(
		.INIT('h13)
	) name6092 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w7441_,
		_w7442_
	);
	LUT4 #(
		.INIT('h8000)
	) name6093 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5762_,
		_w5764_,
		_w7443_
	);
	LUT2 #(
		.INIT('h8)
	) name6094 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('h1)
	) name6095 (
		_w7442_,
		_w7444_,
		_w7445_
	);
	LUT3 #(
		.INIT('h02)
	) name6096 (
		_w3055_,
		_w7442_,
		_w7444_,
		_w7446_
	);
	LUT4 #(
		.INIT('h0080)
	) name6097 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5762_,
		_w6938_,
		_w7447_
	);
	LUT4 #(
		.INIT('hb030)
	) name6098 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2194_,
		_w5783_,
		_w7447_,
		_w7448_
	);
	LUT2 #(
		.INIT('h4)
	) name6099 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2194_,
		_w7449_
	);
	LUT4 #(
		.INIT('h1333)
	) name6100 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w4768_,
		_w7447_,
		_w7449_,
		_w7450_
	);
	LUT3 #(
		.INIT('hd0)
	) name6101 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w7448_,
		_w7450_,
		_w7451_
	);
	LUT2 #(
		.INIT('h4)
	) name6102 (
		_w7446_,
		_w7451_,
		_w7452_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6103 (
		_w1945_,
		_w7438_,
		_w7440_,
		_w7452_,
		_w7453_
	);
	LUT3 #(
		.INIT('h02)
	) name6104 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7454_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6105 (
		_w2900_,
		_w4068_,
		_w4074_,
		_w5348_,
		_w7455_
	);
	LUT4 #(
		.INIT('h1555)
	) name6106 (
		_w2755_,
		_w2879_,
		_w2874_,
		_w5349_,
		_w7456_
	);
	LUT2 #(
		.INIT('h4)
	) name6107 (
		_w7455_,
		_w7456_,
		_w7457_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name6108 (
		_w2965_,
		_w4051_,
		_w4054_,
		_w4057_,
		_w7458_
	);
	LUT3 #(
		.INIT('h51)
	) name6109 (
		_w2173_,
		_w2755_,
		_w7458_,
		_w7459_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6110 (
		_w2171_,
		_w7454_,
		_w7457_,
		_w7459_,
		_w7460_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6111 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7461_
	);
	LUT3 #(
		.INIT('h6c)
	) name6112 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w3029_,
		_w7462_
	);
	LUT4 #(
		.INIT('h0080)
	) name6113 (
		_w2991_,
		_w3024_,
		_w3027_,
		_w4088_,
		_w7463_
	);
	LUT3 #(
		.INIT('h13)
	) name6114 (
		_w2708_,
		_w7462_,
		_w7463_,
		_w7464_
	);
	LUT2 #(
		.INIT('h2)
	) name6115 (
		_w2181_,
		_w4089_,
		_w7465_
	);
	LUT3 #(
		.INIT('h45)
	) name6116 (
		_w7461_,
		_w7464_,
		_w7465_,
		_w7466_
	);
	LUT4 #(
		.INIT('h8000)
	) name6117 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5766_,
		_w5768_,
		_w7467_
	);
	LUT4 #(
		.INIT('h8000)
	) name6118 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5766_,
		_w5769_,
		_w7468_
	);
	LUT3 #(
		.INIT('h0e)
	) name6119 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w7467_,
		_w7468_,
		_w7469_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6120 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w6350_,
		_w7467_,
		_w7468_,
		_w7470_
	);
	LUT4 #(
		.INIT('h1333)
	) name6121 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		_w5766_,
		_w5768_,
		_w7471_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6122 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2199_,
		_w5766_,
		_w5769_,
		_w7472_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6123 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7473_
	);
	LUT3 #(
		.INIT('hb0)
	) name6124 (
		_w7471_,
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h4)
	) name6125 (
		_w7470_,
		_w7474_,
		_w7475_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6126 (
		_w1945_,
		_w7460_,
		_w7466_,
		_w7475_,
		_w7476_
	);
	LUT3 #(
		.INIT('h02)
	) name6127 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7477_
	);
	LUT4 #(
		.INIT('haa20)
	) name6128 (
		_w2171_,
		_w4775_,
		_w4780_,
		_w7477_,
		_w7478_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6129 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7479_
	);
	LUT3 #(
		.INIT('h0b)
	) name6130 (
		_w4782_,
		_w4783_,
		_w7479_,
		_w7480_
	);
	LUT3 #(
		.INIT('h6c)
	) name6131 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w7481_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6132 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w6350_,
		_w7482_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6133 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7483_
	);
	LUT4 #(
		.INIT('hb700)
	) name6134 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2199_,
		_w5771_,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('h4)
	) name6135 (
		_w7482_,
		_w7484_,
		_w7485_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6136 (
		_w1945_,
		_w7478_,
		_w7480_,
		_w7485_,
		_w7486_
	);
	LUT3 #(
		.INIT('h14)
	) name6137 (
		_w2755_,
		_w2905_,
		_w5381_,
		_w7487_
	);
	LUT3 #(
		.INIT('h28)
	) name6138 (
		_w2755_,
		_w4060_,
		_w4061_,
		_w7488_
	);
	LUT4 #(
		.INIT('h2220)
	) name6139 (
		_w2171_,
		_w2173_,
		_w7487_,
		_w7488_,
		_w7489_
	);
	LUT3 #(
		.INIT('h6c)
	) name6140 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w3033_,
		_w7490_
	);
	LUT4 #(
		.INIT('h8000)
	) name6141 (
		\P3_InstAddrPointer_reg[22]/NET0131 ,
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w3032_,
		_w4089_,
		_w7491_
	);
	LUT3 #(
		.INIT('h2a)
	) name6142 (
		_w2181_,
		_w3036_,
		_w4089_,
		_w7492_
	);
	LUT2 #(
		.INIT('h2)
	) name6143 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w7422_,
		_w7493_
	);
	LUT4 #(
		.INIT('h001f)
	) name6144 (
		_w7490_,
		_w7491_,
		_w7492_,
		_w7493_,
		_w7494_
	);
	LUT4 #(
		.INIT('h8000)
	) name6145 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w5772_,
		_w7495_
	);
	LUT3 #(
		.INIT('h0e)
	) name6146 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w6942_,
		_w7495_,
		_w7496_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6147 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w6350_,
		_w6942_,
		_w7495_,
		_w7497_
	);
	LUT4 #(
		.INIT('h070f)
	) name6148 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		_w5771_,
		_w7498_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6149 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2199_,
		_w5771_,
		_w5772_,
		_w7499_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6150 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7500_
	);
	LUT3 #(
		.INIT('hb0)
	) name6151 (
		_w7498_,
		_w7499_,
		_w7500_,
		_w7501_
	);
	LUT2 #(
		.INIT('h4)
	) name6152 (
		_w7497_,
		_w7501_,
		_w7502_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6153 (
		_w1945_,
		_w7489_,
		_w7494_,
		_w7502_,
		_w7503_
	);
	LUT3 #(
		.INIT('h02)
	) name6154 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7504_
	);
	LUT4 #(
		.INIT('h8222)
	) name6155 (
		_w2755_,
		_w2969_,
		_w4772_,
		_w6334_,
		_w7505_
	);
	LUT4 #(
		.INIT('h4554)
	) name6156 (
		_w2173_,
		_w2755_,
		_w2911_,
		_w6340_,
		_w7506_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6157 (
		_w2171_,
		_w7504_,
		_w7505_,
		_w7506_,
		_w7507_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6158 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7508_
	);
	LUT2 #(
		.INIT('h6)
	) name6159 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w3038_,
		_w7509_
	);
	LUT4 #(
		.INIT('h007f)
	) name6160 (
		_w3036_,
		_w3039_,
		_w4089_,
		_w7509_,
		_w7510_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name6161 (
		_w2181_,
		_w4090_,
		_w7508_,
		_w7510_,
		_w7511_
	);
	LUT4 #(
		.INIT('h8000)
	) name6162 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w5771_,
		_w5773_,
		_w7512_
	);
	LUT3 #(
		.INIT('h32)
	) name6163 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5775_,
		_w7512_,
		_w7513_
	);
	LUT4 #(
		.INIT('h3020)
	) name6164 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5775_,
		_w6350_,
		_w7512_,
		_w7514_
	);
	LUT4 #(
		.INIT('h1333)
	) name6165 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		_w5771_,
		_w5773_,
		_w7515_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6166 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2199_,
		_w5771_,
		_w5774_,
		_w7516_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6167 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7517_
	);
	LUT3 #(
		.INIT('hb0)
	) name6168 (
		_w7515_,
		_w7516_,
		_w7517_,
		_w7518_
	);
	LUT2 #(
		.INIT('h4)
	) name6169 (
		_w7514_,
		_w7518_,
		_w7519_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6170 (
		_w1945_,
		_w7507_,
		_w7511_,
		_w7519_,
		_w7520_
	);
	LUT3 #(
		.INIT('h08)
	) name6171 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7521_
	);
	LUT4 #(
		.INIT('h3332)
	) name6172 (
		_w3300_,
		_w4463_,
		_w4445_,
		_w4447_,
		_w7522_
	);
	LUT4 #(
		.INIT('h4554)
	) name6173 (
		_w1916_,
		_w3101_,
		_w3216_,
		_w4474_,
		_w7523_
	);
	LUT4 #(
		.INIT('h0233)
	) name6174 (
		_w3101_,
		_w7521_,
		_w7522_,
		_w7523_,
		_w7524_
	);
	LUT4 #(
		.INIT('h8288)
	) name6175 (
		_w1924_,
		_w3362_,
		_w4023_,
		_w4025_,
		_w7525_
	);
	LUT4 #(
		.INIT('h028a)
	) name6176 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7526_
	);
	LUT2 #(
		.INIT('h1)
	) name6177 (
		_w7525_,
		_w7526_,
		_w7527_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6178 (
		_w1810_,
		_w1933_,
		_w7524_,
		_w7527_,
		_w7528_
	);
	LUT4 #(
		.INIT('h8000)
	) name6179 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w6365_,
		_w7529_
	);
	LUT4 #(
		.INIT('h8000)
	) name6180 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w7529_,
		_w7530_
	);
	LUT2 #(
		.INIT('h6)
	) name6181 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w7530_,
		_w7531_
	);
	LUT3 #(
		.INIT('h41)
	) name6182 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w7530_,
		_w7532_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6183 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w6367_,
		_w7533_
	);
	LUT3 #(
		.INIT('hc4)
	) name6184 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w7533_,
		_w7534_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6185 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7535_
	);
	LUT4 #(
		.INIT('hb700)
	) name6186 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w3407_,
		_w7530_,
		_w7535_,
		_w7536_
	);
	LUT3 #(
		.INIT('hb0)
	) name6187 (
		_w7532_,
		_w7534_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('hb)
	) name6188 (
		_w7528_,
		_w7537_,
		_w7538_
	);
	LUT3 #(
		.INIT('h6c)
	) name6189 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w3069_,
		_w7539_
	);
	LUT4 #(
		.INIT('h8000)
	) name6190 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3296_,
		_w3302_,
		_w3993_,
		_w7540_
	);
	LUT4 #(
		.INIT('h888a)
	) name6191 (
		_w3101_,
		_w4466_,
		_w7539_,
		_w7540_,
		_w7541_
	);
	LUT3 #(
		.INIT('h2a)
	) name6192 (
		_w3243_,
		_w4474_,
		_w4475_,
		_w7542_
	);
	LUT4 #(
		.INIT('h5554)
	) name6193 (
		_w1916_,
		_w3101_,
		_w5455_,
		_w7542_,
		_w7543_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name6194 (
		_w4023_,
		_w4025_,
		_w4026_,
		_w4027_,
		_w7544_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6195 (
		_w1924_,
		_w4023_,
		_w4025_,
		_w4028_,
		_w7545_
	);
	LUT2 #(
		.INIT('h4)
	) name6196 (
		_w7544_,
		_w7545_,
		_w7546_
	);
	LUT4 #(
		.INIT('h20e4)
	) name6197 (
		_w1809_,
		_w1810_,
		_w1846_,
		_w1916_,
		_w7547_
	);
	LUT2 #(
		.INIT('h2)
	) name6198 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w7547_,
		_w7548_
	);
	LUT3 #(
		.INIT('h0b)
	) name6199 (
		_w7544_,
		_w7545_,
		_w7548_,
		_w7549_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6200 (
		_w1810_,
		_w7541_,
		_w7543_,
		_w7549_,
		_w7550_
	);
	LUT4 #(
		.INIT('h8000)
	) name6201 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w7530_,
		_w7551_
	);
	LUT3 #(
		.INIT('h6c)
	) name6202 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w7551_,
		_w7552_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6203 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w6378_,
		_w7551_,
		_w7553_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6204 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7554_
	);
	LUT4 #(
		.INIT('hb700)
	) name6205 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w2310_,
		_w6370_,
		_w7554_,
		_w7555_
	);
	LUT2 #(
		.INIT('h4)
	) name6206 (
		_w7553_,
		_w7555_,
		_w7556_
	);
	LUT3 #(
		.INIT('h2f)
	) name6207 (
		_w1933_,
		_w7550_,
		_w7556_,
		_w7557_
	);
	LUT3 #(
		.INIT('h08)
	) name6208 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7558_
	);
	LUT4 #(
		.INIT('h888a)
	) name6209 (
		_w3101_,
		_w4468_,
		_w4450_,
		_w5458_,
		_w7559_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6210 (
		_w3248_,
		_w3250_,
		_w4474_,
		_w4475_,
		_w7560_
	);
	LUT3 #(
		.INIT('h54)
	) name6211 (
		_w1916_,
		_w3101_,
		_w7560_,
		_w7561_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6212 (
		_w1810_,
		_w7558_,
		_w7559_,
		_w7561_,
		_w7562_
	);
	LUT3 #(
		.INIT('h13)
	) name6213 (
		_w3073_,
		_w3374_,
		_w5924_,
		_w7563_
	);
	LUT2 #(
		.INIT('h2)
	) name6214 (
		_w1924_,
		_w4030_,
		_w7564_
	);
	LUT4 #(
		.INIT('h028a)
	) name6215 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7565_
	);
	LUT3 #(
		.INIT('h0b)
	) name6216 (
		_w7563_,
		_w7564_,
		_w7565_,
		_w7566_
	);
	LUT4 #(
		.INIT('h070f)
	) name6217 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w6372_,
		_w7567_
	);
	LUT3 #(
		.INIT('h80)
	) name6218 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w6379_,
		_w7568_
	);
	LUT4 #(
		.INIT('h8000)
	) name6219 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w6379_,
		_w7569_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		_w7567_,
		_w7569_,
		_w7570_
	);
	LUT3 #(
		.INIT('h02)
	) name6221 (
		_w6378_,
		_w7567_,
		_w7569_,
		_w7571_
	);
	LUT4 #(
		.INIT('hb300)
	) name6222 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w2310_,
		_w6379_,
		_w6383_,
		_w7572_
	);
	LUT3 #(
		.INIT('h20)
	) name6223 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w1939_,
		_w7573_
	);
	LUT2 #(
		.INIT('h8)
	) name6224 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w3406_,
		_w7574_
	);
	LUT4 #(
		.INIT('h007f)
	) name6225 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w6379_,
		_w7573_,
		_w7574_,
		_w7575_
	);
	LUT3 #(
		.INIT('hd0)
	) name6226 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w7572_,
		_w7575_,
		_w7576_
	);
	LUT2 #(
		.INIT('h4)
	) name6227 (
		_w7571_,
		_w7576_,
		_w7577_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6228 (
		_w1933_,
		_w7562_,
		_w7566_,
		_w7577_,
		_w7578_
	);
	LUT3 #(
		.INIT('h08)
	) name6229 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7579_
	);
	LUT4 #(
		.INIT('haa20)
	) name6230 (
		_w1810_,
		_w4935_,
		_w4937_,
		_w7579_,
		_w7580_
	);
	LUT4 #(
		.INIT('h028a)
	) name6231 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7581_
	);
	LUT2 #(
		.INIT('h1)
	) name6232 (
		_w4939_,
		_w7581_,
		_w7582_
	);
	LUT4 #(
		.INIT('h8000)
	) name6233 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w6379_,
		_w7583_
	);
	LUT3 #(
		.INIT('h6c)
	) name6234 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w7568_,
		_w7584_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6235 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w6378_,
		_w7568_,
		_w7585_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6236 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7586_
	);
	LUT4 #(
		.INIT('hb700)
	) name6237 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		_w2310_,
		_w7568_,
		_w7586_,
		_w7587_
	);
	LUT2 #(
		.INIT('h4)
	) name6238 (
		_w7585_,
		_w7587_,
		_w7588_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6239 (
		_w1933_,
		_w7580_,
		_w7582_,
		_w7588_,
		_w7589_
	);
	LUT3 #(
		.INIT('h08)
	) name6240 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7590_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6241 (
		_w3237_,
		_w3247_,
		_w4476_,
		_w5455_,
		_w7591_
	);
	LUT4 #(
		.INIT('h1555)
	) name6242 (
		_w3101_,
		_w3247_,
		_w4477_,
		_w5455_,
		_w7592_
	);
	LUT4 #(
		.INIT('h1551)
	) name6243 (
		_w1916_,
		_w3101_,
		_w3313_,
		_w3312_,
		_w7593_
	);
	LUT4 #(
		.INIT('h1055)
	) name6244 (
		_w7590_,
		_w7591_,
		_w7592_,
		_w7593_,
		_w7594_
	);
	LUT4 #(
		.INIT('h028a)
	) name6245 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7595_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6246 (
		_w1924_,
		_w3377_,
		_w3382_,
		_w7595_,
		_w7596_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6247 (
		_w1810_,
		_w1933_,
		_w7594_,
		_w7596_,
		_w7597_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6248 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w6363_,
		_w6372_,
		_w7598_
	);
	LUT4 #(
		.INIT('h4888)
	) name6249 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		_w2310_,
		_w6379_,
		_w6363_,
		_w7599_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6250 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7600_
	);
	LUT4 #(
		.INIT('h0700)
	) name6251 (
		_w6378_,
		_w7598_,
		_w7599_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('hb)
	) name6252 (
		_w7597_,
		_w7601_,
		_w7602_
	);
	LUT3 #(
		.INIT('h08)
	) name6253 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7603_
	);
	LUT4 #(
		.INIT('haa20)
	) name6254 (
		_w1810_,
		_w4723_,
		_w4732_,
		_w7603_,
		_w7604_
	);
	LUT4 #(
		.INIT('h028a)
	) name6255 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7605_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6256 (
		_w1924_,
		_w4734_,
		_w4737_,
		_w7605_,
		_w7606_
	);
	LUT4 #(
		.INIT('h8000)
	) name6257 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		_w6379_,
		_w6363_,
		_w7607_
	);
	LUT4 #(
		.INIT('h74fc)
	) name6258 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w6997_,
		_w7607_,
		_w7608_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6259 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w3406_,
		_w6383_,
		_w7609_
	);
	LUT4 #(
		.INIT('hb700)
	) name6260 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w2310_,
		_w7607_,
		_w7609_,
		_w7610_
	);
	LUT3 #(
		.INIT('h70)
	) name6261 (
		_w6378_,
		_w7608_,
		_w7610_,
		_w7611_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6262 (
		_w1933_,
		_w7604_,
		_w7606_,
		_w7611_,
		_w7612_
	);
	LUT3 #(
		.INIT('h08)
	) name6263 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1842_,
		_w1915_,
		_w7613_
	);
	LUT4 #(
		.INIT('haa20)
	) name6264 (
		_w1810_,
		_w4704_,
		_w4705_,
		_w7613_,
		_w7614_
	);
	LUT4 #(
		.INIT('h028a)
	) name6265 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w7615_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6266 (
		_w1924_,
		_w3385_,
		_w3386_,
		_w7615_,
		_w7616_
	);
	LUT2 #(
		.INIT('h6)
	) name6267 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6374_,
		_w7617_
	);
	LUT3 #(
		.INIT('h60)
	) name6268 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6374_,
		_w6378_,
		_w7618_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6269 (
		_w2310_,
		_w6379_,
		_w6363_,
		_w6362_,
		_w7619_
	);
	LUT3 #(
		.INIT('ha2)
	) name6270 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6383_,
		_w7619_,
		_w7620_
	);
	LUT3 #(
		.INIT('h20)
	) name6271 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w1939_,
		_w7621_
	);
	LUT4 #(
		.INIT('h8000)
	) name6272 (
		_w6379_,
		_w6363_,
		_w6362_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h1)
	) name6273 (
		_w4717_,
		_w7622_,
		_w7623_
	);
	LUT3 #(
		.INIT('h10)
	) name6274 (
		_w7620_,
		_w7618_,
		_w7623_,
		_w7624_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6275 (
		_w1933_,
		_w7614_,
		_w7616_,
		_w7624_,
		_w7625_
	);
	LUT3 #(
		.INIT('h08)
	) name6276 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7626_
	);
	LUT4 #(
		.INIT('h028a)
	) name6277 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w5406_,
		_w7627_,
		_w7628_
	);
	LUT4 #(
		.INIT('h5700)
	) name6279 (
		_w1559_,
		_w5405_,
		_w7626_,
		_w7628_,
		_w7629_
	);
	LUT3 #(
		.INIT('h80)
	) name6280 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w7630_
	);
	LUT4 #(
		.INIT('h8000)
	) name6281 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w7631_
	);
	LUT3 #(
		.INIT('h6c)
	) name6282 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w7630_,
		_w7632_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6283 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w2283_,
		_w7630_,
		_w7633_
	);
	LUT3 #(
		.INIT('h80)
	) name6284 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w7634_
	);
	LUT4 #(
		.INIT('h0080)
	) name6285 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w6857_,
		_w7635_
	);
	LUT4 #(
		.INIT('h0080)
	) name6286 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w6857_,
		_w7636_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6287 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w1679_,
		_w7635_,
		_w7636_,
		_w7637_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6288 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7638_
	);
	LUT3 #(
		.INIT('h10)
	) name6289 (
		_w7637_,
		_w7633_,
		_w7638_,
		_w7639_
	);
	LUT3 #(
		.INIT('h2f)
	) name6290 (
		_w1678_,
		_w7629_,
		_w7639_,
		_w7640_
	);
	LUT4 #(
		.INIT('h2022)
	) name6291 (
		_w1559_,
		_w1661_,
		_w4812_,
		_w4829_,
		_w7641_
	);
	LUT4 #(
		.INIT('h20e4)
	) name6292 (
		_w1558_,
		_w1559_,
		_w1596_,
		_w1661_,
		_w7642_
	);
	LUT2 #(
		.INIT('h2)
	) name6293 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w7642_,
		_w7643_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6294 (
		_w1659_,
		_w4831_,
		_w4839_,
		_w7643_,
		_w7644_
	);
	LUT4 #(
		.INIT('h8848)
	) name6295 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w1679_,
		_w5730_,
		_w6857_,
		_w7645_
	);
	LUT3 #(
		.INIT('h6a)
	) name6296 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5730_,
		_w7646_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6297 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w2283_,
		_w5730_,
		_w7647_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6298 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7648_
	);
	LUT3 #(
		.INIT('h10)
	) name6299 (
		_w7647_,
		_w7645_,
		_w7648_,
		_w7649_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6300 (
		_w1678_,
		_w7641_,
		_w7644_,
		_w7649_,
		_w7650_
	);
	LUT3 #(
		.INIT('h08)
	) name6301 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7651_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6302 (
		_w4346_,
		_w4821_,
		_w4826_,
		_w5695_,
		_w7652_
	);
	LUT3 #(
		.INIT('h01)
	) name6303 (
		_w4214_,
		_w6845_,
		_w7652_,
		_w7653_
	);
	LUT3 #(
		.INIT('h07)
	) name6304 (
		_w4796_,
		_w4896_,
		_w4898_,
		_w7654_
	);
	LUT4 #(
		.INIT('h1115)
	) name6305 (
		_w1661_,
		_w4214_,
		_w4860_,
		_w7654_,
		_w7655_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6306 (
		_w1559_,
		_w7651_,
		_w7653_,
		_w7655_,
		_w7656_
	);
	LUT4 #(
		.INIT('h028a)
	) name6307 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7657_
	);
	LUT3 #(
		.INIT('h28)
	) name6308 (
		_w1659_,
		_w4873_,
		_w5715_,
		_w7658_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6309 (
		_w1659_,
		_w4873_,
		_w5715_,
		_w7657_,
		_w7659_
	);
	LUT4 #(
		.INIT('h8000)
	) name6310 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5730_,
		_w5731_,
		_w7660_
	);
	LUT3 #(
		.INIT('h6a)
	) name6311 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5732_,
		_w7661_
	);
	LUT4 #(
		.INIT('h6a00)
	) name6312 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5732_,
		_w5746_,
		_w7662_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6313 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7663_
	);
	LUT4 #(
		.INIT('hb700)
	) name6314 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w2242_,
		_w5732_,
		_w7663_,
		_w7664_
	);
	LUT2 #(
		.INIT('h4)
	) name6315 (
		_w7662_,
		_w7664_,
		_w7665_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6316 (
		_w1678_,
		_w7656_,
		_w7659_,
		_w7665_,
		_w7666_
	);
	LUT3 #(
		.INIT('h02)
	) name6317 (
		_w3335_,
		_w3339_,
		_w4018_,
		_w7667_
	);
	LUT3 #(
		.INIT('h87)
	) name6318 (
		_w3175_,
		_w3180_,
		_w3332_,
		_w7668_
	);
	LUT3 #(
		.INIT('h0e)
	) name6319 (
		_w3334_,
		_w4018_,
		_w7668_,
		_w7669_
	);
	LUT3 #(
		.INIT('h02)
	) name6320 (
		_w1924_,
		_w7669_,
		_w7667_,
		_w7670_
	);
	LUT3 #(
		.INIT('h87)
	) name6321 (
		_w3175_,
		_w3180_,
		_w3279_,
		_w7671_
	);
	LUT4 #(
		.INIT('ha802)
	) name6322 (
		_w3101_,
		_w3273_,
		_w3276_,
		_w7671_,
		_w7672_
	);
	LUT3 #(
		.INIT('h87)
	) name6323 (
		_w3175_,
		_w3180_,
		_w3181_,
		_w7673_
	);
	LUT4 #(
		.INIT('h0154)
	) name6324 (
		_w3101_,
		_w3197_,
		_w4000_,
		_w7673_,
		_w7674_
	);
	LUT3 #(
		.INIT('h02)
	) name6325 (
		_w1923_,
		_w7674_,
		_w7672_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name6326 (
		_w7670_,
		_w7675_,
		_w7676_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6327 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		_w1914_,
		_w1917_,
		_w1868_,
		_w7677_
	);
	LUT2 #(
		.INIT('h4)
	) name6328 (
		_w1862_,
		_w3279_,
		_w7678_
	);
	LUT3 #(
		.INIT('h40)
	) name6329 (
		_w1833_,
		_w1846_,
		_w3332_,
		_w7679_
	);
	LUT4 #(
		.INIT('h004f)
	) name6330 (
		_w1816_,
		_w1831_,
		_w3181_,
		_w7679_,
		_w7680_
	);
	LUT4 #(
		.INIT('h0400)
	) name6331 (
		_w7677_,
		_w7676_,
		_w7678_,
		_w7680_,
		_w7681_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6332 (
		\P1_InstAddrPointer_reg[3]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w3406_,
		_w3408_,
		_w7682_
	);
	LUT3 #(
		.INIT('h2f)
	) name6333 (
		_w1933_,
		_w7681_,
		_w7682_,
		_w7683_
	);
	LUT3 #(
		.INIT('h95)
	) name6334 (
		_w3288_,
		_w3108_,
		_w3113_,
		_w7684_
	);
	LUT4 #(
		.INIT('h4774)
	) name6335 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1916_,
		_w3285_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('h2)
	) name6336 (
		_w1810_,
		_w7685_,
		_w7686_
	);
	LUT3 #(
		.INIT('ha2)
	) name6337 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		_w1914_,
		_w1868_,
		_w7687_
	);
	LUT3 #(
		.INIT('h40)
	) name6338 (
		_w1833_,
		_w1846_,
		_w3327_,
		_w7688_
	);
	LUT4 #(
		.INIT('h004f)
	) name6339 (
		_w1816_,
		_w1831_,
		_w3115_,
		_w7688_,
		_w7689_
	);
	LUT2 #(
		.INIT('h4)
	) name6340 (
		_w3344_,
		_w4020_,
		_w7690_
	);
	LUT3 #(
		.INIT('h87)
	) name6341 (
		_w3108_,
		_w3113_,
		_w3327_,
		_w7691_
	);
	LUT4 #(
		.INIT('h0455)
	) name6342 (
		_w3330_,
		_w3335_,
		_w4018_,
		_w4019_,
		_w7692_
	);
	LUT3 #(
		.INIT('ha8)
	) name6343 (
		_w1924_,
		_w7691_,
		_w7692_,
		_w7693_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name6344 (
		_w1862_,
		_w3288_,
		_w7690_,
		_w7693_,
		_w7694_
	);
	LUT4 #(
		.INIT('h1000)
	) name6345 (
		_w7687_,
		_w7686_,
		_w7689_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h8)
	) name6346 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w3406_,
		_w7696_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6347 (
		\P1_InstAddrPointer_reg[5]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w3406_,
		_w3408_,
		_w7697_
	);
	LUT3 #(
		.INIT('h2f)
	) name6348 (
		_w1933_,
		_w7695_,
		_w7697_,
		_w7698_
	);
	LUT3 #(
		.INIT('h87)
	) name6349 (
		_w2803_,
		_w2808_,
		_w2811_,
		_w7699_
	);
	LUT4 #(
		.INIT('hb24d)
	) name6350 (
		_w2769_,
		_w2771_,
		_w2797_,
		_w7699_,
		_w7700_
	);
	LUT3 #(
		.INIT('h87)
	) name6351 (
		_w2803_,
		_w2808_,
		_w2922_,
		_w7701_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6352 (
		_w2755_,
		_w2919_,
		_w2924_,
		_w7701_,
		_w7702_
	);
	LUT4 #(
		.INIT('h5501)
	) name6353 (
		_w2173_,
		_w2755_,
		_w7700_,
		_w7702_,
		_w7703_
	);
	LUT3 #(
		.INIT('h01)
	) name6354 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7704_
	);
	LUT3 #(
		.INIT('h04)
	) name6355 (
		_w2060_,
		_w2041_,
		_w7704_,
		_w7705_
	);
	LUT2 #(
		.INIT('h4)
	) name6356 (
		_w7703_,
		_w7705_,
		_w7706_
	);
	LUT2 #(
		.INIT('h4)
	) name6357 (
		_w2117_,
		_w2922_,
		_w7707_
	);
	LUT3 #(
		.INIT('hb0)
	) name6358 (
		_w2073_,
		_w2086_,
		_w2811_,
		_w7708_
	);
	LUT4 #(
		.INIT('haaa2)
	) name6359 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2122_,
		_w2125_,
		_w2175_,
		_w7709_
	);
	LUT3 #(
		.INIT('ha6)
	) name6360 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		_w2098_,
		_w2770_,
		_w7710_
	);
	LUT3 #(
		.INIT('he0)
	) name6361 (
		_w2071_,
		_w2087_,
		_w7710_,
		_w7711_
	);
	LUT3 #(
		.INIT('h04)
	) name6362 (
		_w3006_,
		_w3010_,
		_w3011_,
		_w7712_
	);
	LUT3 #(
		.INIT('h87)
	) name6363 (
		_w2803_,
		_w2808_,
		_w3008_,
		_w7713_
	);
	LUT3 #(
		.INIT('h0e)
	) name6364 (
		_w3006_,
		_w3007_,
		_w7713_,
		_w7714_
	);
	LUT3 #(
		.INIT('h02)
	) name6365 (
		_w2181_,
		_w7714_,
		_w7712_,
		_w7715_
	);
	LUT3 #(
		.INIT('h01)
	) name6366 (
		_w7711_,
		_w7709_,
		_w7715_,
		_w7716_
	);
	LUT4 #(
		.INIT('h0100)
	) name6367 (
		_w7708_,
		_w7707_,
		_w7706_,
		_w7716_,
		_w7717_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6368 (
		\P3_InstAddrPointer_reg[3]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w3054_,
		_w3056_,
		_w7718_
	);
	LUT3 #(
		.INIT('h2f)
	) name6369 (
		_w1945_,
		_w7717_,
		_w7718_,
		_w7719_
	);
	LUT2 #(
		.INIT('h2)
	) name6370 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		_w7103_,
		_w7720_
	);
	LUT3 #(
		.INIT('h95)
	) name6371 (
		_w2930_,
		_w2849_,
		_w2854_,
		_w7721_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name6372 (
		_w2919_,
		_w2926_,
		_w2929_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h2)
	) name6373 (
		_w2180_,
		_w7722_,
		_w7723_
	);
	LUT4 #(
		.INIT('he000)
	) name6374 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2998_,
		_w7724_
	);
	LUT4 #(
		.INIT('h000b)
	) name6375 (
		_w2117_,
		_w2930_,
		_w7723_,
		_w7724_,
		_w7725_
	);
	LUT3 #(
		.INIT('hb0)
	) name6376 (
		_w2073_,
		_w2086_,
		_w2856_,
		_w7726_
	);
	LUT2 #(
		.INIT('h2)
	) name6377 (
		_w3014_,
		_w3016_,
		_w7727_
	);
	LUT3 #(
		.INIT('h87)
	) name6378 (
		_w2849_,
		_w2854_,
		_w2998_,
		_w7728_
	);
	LUT4 #(
		.INIT('h1055)
	) name6379 (
		_w2997_,
		_w3006_,
		_w3010_,
		_w3013_,
		_w7729_
	);
	LUT3 #(
		.INIT('ha8)
	) name6380 (
		_w2181_,
		_w7728_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h4)
	) name6381 (
		_w7727_,
		_w7730_,
		_w7731_
	);
	LUT3 #(
		.INIT('h10)
	) name6382 (
		_w7726_,
		_w7731_,
		_w7725_,
		_w7732_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6383 (
		\P3_InstAddrPointer_reg[5]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w3054_,
		_w3056_,
		_w7733_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6384 (
		_w1945_,
		_w7720_,
		_w7732_,
		_w7733_,
		_w7734_
	);
	LUT3 #(
		.INIT('hb0)
	) name6385 (
		_w1571_,
		_w1583_,
		_w4300_,
		_w7735_
	);
	LUT2 #(
		.INIT('h8)
	) name6386 (
		_w1640_,
		_w4384_,
		_w7736_
	);
	LUT3 #(
		.INIT('h87)
	) name6387 (
		_w4160_,
		_w4165_,
		_w4384_,
		_w7737_
	);
	LUT3 #(
		.INIT('h0e)
	) name6388 (
		_w4387_,
		_w4391_,
		_w7737_,
		_w7738_
	);
	LUT3 #(
		.INIT('h10)
	) name6389 (
		_w4387_,
		_w4391_,
		_w7737_,
		_w7739_
	);
	LUT3 #(
		.INIT('h02)
	) name6390 (
		_w1659_,
		_w7739_,
		_w7738_,
		_w7740_
	);
	LUT4 #(
		.INIT('h000b)
	) name6391 (
		_w1617_,
		_w4166_,
		_w7736_,
		_w7740_,
		_w7741_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name6392 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		_w1614_,
		_w1666_,
		_w1668_,
		_w7742_
	);
	LUT3 #(
		.INIT('h87)
	) name6393 (
		_w4160_,
		_w4165_,
		_w4166_,
		_w7743_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6394 (
		_w4214_,
		_w4142_,
		_w4168_,
		_w7743_,
		_w7744_
	);
	LUT3 #(
		.INIT('h87)
	) name6395 (
		_w4160_,
		_w4165_,
		_w4300_,
		_w7745_
	);
	LUT4 #(
		.INIT('h0154)
	) name6396 (
		_w4214_,
		_w4297_,
		_w4302_,
		_w7745_,
		_w7746_
	);
	LUT4 #(
		.INIT('h0002)
	) name6397 (
		_w1559_,
		_w1661_,
		_w7746_,
		_w7744_,
		_w7747_
	);
	LUT4 #(
		.INIT('h0100)
	) name6398 (
		_w7742_,
		_w7747_,
		_w7735_,
		_w7741_,
		_w7748_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6399 (
		\P2_InstAddrPointer_reg[3]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w2286_,
		_w4441_,
		_w7749_
	);
	LUT3 #(
		.INIT('h2f)
	) name6400 (
		_w1678_,
		_w7748_,
		_w7749_,
		_w7750_
	);
	LUT3 #(
		.INIT('h87)
	) name6401 (
		_w4192_,
		_w4197_,
		_w4379_,
		_w7751_
	);
	LUT3 #(
		.INIT('h82)
	) name6402 (
		_w1659_,
		_w4395_,
		_w7751_,
		_w7752_
	);
	LUT2 #(
		.INIT('h4)
	) name6403 (
		_w1617_,
		_w4198_,
		_w7753_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6404 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w1657_,
		_w6446_,
		_w6447_,
		_w7754_
	);
	LUT3 #(
		.INIT('h01)
	) name6405 (
		_w7753_,
		_w7754_,
		_w7752_,
		_w7755_
	);
	LUT3 #(
		.INIT('h87)
	) name6406 (
		_w4192_,
		_w4197_,
		_w4198_,
		_w7756_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name6407 (
		_w4142_,
		_w4170_,
		_w4173_,
		_w7756_,
		_w7757_
	);
	LUT4 #(
		.INIT('h808c)
	) name6408 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w1559_,
		_w1661_,
		_w7757_,
		_w7758_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name6409 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		_w1592_,
		_w1595_,
		_w4373_,
		_w7759_
	);
	LUT4 #(
		.INIT('hc800)
	) name6410 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w7759_,
		_w7760_
	);
	LUT4 #(
		.INIT('h004f)
	) name6411 (
		_w1571_,
		_w1583_,
		_w4287_,
		_w7760_,
		_w7761_
	);
	LUT2 #(
		.INIT('h4)
	) name6412 (
		_w7758_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w2286_,
		_w7763_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6414 (
		\P2_InstAddrPointer_reg[5]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w2286_,
		_w4441_,
		_w7764_
	);
	LUT4 #(
		.INIT('h2aff)
	) name6415 (
		_w1678_,
		_w7755_,
		_w7762_,
		_w7764_,
		_w7765_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name6416 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w7766_
	);
	LUT4 #(
		.INIT('hfc20)
	) name6417 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w7767_
	);
	LUT2 #(
		.INIT('h2)
	) name6418 (
		\P2_EAX_reg[31]/NET0131 ,
		_w7767_,
		_w7768_
	);
	LUT4 #(
		.INIT('h8000)
	) name6419 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		_w7769_
	);
	LUT4 #(
		.INIT('h8000)
	) name6420 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		\P2_EAX_reg[6]/NET0131 ,
		_w7769_,
		_w7770_
	);
	LUT4 #(
		.INIT('h8000)
	) name6421 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w7770_,
		_w7771_
	);
	LUT2 #(
		.INIT('h8)
	) name6422 (
		\P2_EAX_reg[10]/NET0131 ,
		_w7771_,
		_w7772_
	);
	LUT3 #(
		.INIT('h80)
	) name6423 (
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		_w7771_,
		_w7773_
	);
	LUT4 #(
		.INIT('h8000)
	) name6424 (
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		\P2_EAX_reg[12]/NET0131 ,
		_w7771_,
		_w7774_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		\P2_EAX_reg[13]/NET0131 ,
		_w7774_,
		_w7775_
	);
	LUT3 #(
		.INIT('h80)
	) name6426 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		_w7774_,
		_w7776_
	);
	LUT4 #(
		.INIT('h8000)
	) name6427 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		\P2_EAX_reg[15]/NET0131 ,
		_w7774_,
		_w7777_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[18]/NET0131 ,
		_w7778_
	);
	LUT3 #(
		.INIT('h80)
	) name6429 (
		\P2_EAX_reg[16]/NET0131 ,
		_w7777_,
		_w7778_,
		_w7779_
	);
	LUT4 #(
		.INIT('h8000)
	) name6430 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		_w7777_,
		_w7778_,
		_w7780_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		\P2_EAX_reg[21]/NET0131 ,
		\P2_EAX_reg[22]/NET0131 ,
		_w7781_
	);
	LUT3 #(
		.INIT('h80)
	) name6432 (
		\P2_EAX_reg[20]/NET0131 ,
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT3 #(
		.INIT('h80)
	) name6433 (
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		\P2_EAX_reg[25]/NET0131 ,
		_w7783_
	);
	LUT4 #(
		.INIT('h8000)
	) name6434 (
		\P2_EAX_reg[20]/NET0131 ,
		_w7780_,
		_w7781_,
		_w7783_,
		_w7784_
	);
	LUT2 #(
		.INIT('h8)
	) name6435 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		_w7785_
	);
	LUT3 #(
		.INIT('h80)
	) name6436 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		\P2_EAX_reg[28]/NET0131 ,
		_w7786_
	);
	LUT3 #(
		.INIT('h80)
	) name6437 (
		\P2_EAX_reg[29]/NET0131 ,
		_w7784_,
		_w7786_,
		_w7787_
	);
	LUT4 #(
		.INIT('h8000)
	) name6438 (
		\P2_EAX_reg[29]/NET0131 ,
		\P2_EAX_reg[30]/NET0131 ,
		_w7784_,
		_w7786_,
		_w7788_
	);
	LUT4 #(
		.INIT('h8000)
	) name6439 (
		_w1552_,
		_w1561_,
		_w1564_,
		_w1572_,
		_w7789_
	);
	LUT3 #(
		.INIT('h07)
	) name6440 (
		_w1549_,
		_w1553_,
		_w7789_,
		_w7790_
	);
	LUT3 #(
		.INIT('h13)
	) name6441 (
		_w1604_,
		_w1642_,
		_w7790_,
		_w7791_
	);
	LUT4 #(
		.INIT('h0103)
	) name6442 (
		_w1604_,
		_w1607_,
		_w1642_,
		_w7790_,
		_w7792_
	);
	LUT4 #(
		.INIT('h20aa)
	) name6443 (
		\P2_EAX_reg[31]/NET0131 ,
		_w7788_,
		_w7789_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h4)
	) name6444 (
		\P2_EAX_reg[31]/NET0131 ,
		_w7789_,
		_w7794_
	);
	LUT4 #(
		.INIT('h153f)
	) name6445 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1446_,
		_w1460_,
		_w7795_
	);
	LUT4 #(
		.INIT('h135f)
	) name6446 (
		\P2_InstQueue_reg[4][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1462_,
		_w1466_,
		_w7796_
	);
	LUT4 #(
		.INIT('h135f)
	) name6447 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1443_,
		_w1456_,
		_w7797_
	);
	LUT4 #(
		.INIT('h153f)
	) name6448 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[2][7]/NET0131 ,
		_w1453_,
		_w1447_,
		_w7798_
	);
	LUT4 #(
		.INIT('h8000)
	) name6449 (
		_w7797_,
		_w7798_,
		_w7795_,
		_w7796_,
		_w7799_
	);
	LUT4 #(
		.INIT('h153f)
	) name6450 (
		\P2_InstQueue_reg[6][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1449_,
		_w1450_,
		_w7800_
	);
	LUT4 #(
		.INIT('h135f)
	) name6451 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1452_,
		_w1459_,
		_w7801_
	);
	LUT4 #(
		.INIT('h135f)
	) name6452 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w1465_,
		_w1457_,
		_w7802_
	);
	LUT4 #(
		.INIT('h135f)
	) name6453 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1444_,
		_w1463_,
		_w7803_
	);
	LUT4 #(
		.INIT('h8000)
	) name6454 (
		_w7802_,
		_w7803_,
		_w7800_,
		_w7801_,
		_w7804_
	);
	LUT4 #(
		.INIT('h135f)
	) name6455 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7805_
	);
	LUT4 #(
		.INIT('h135f)
	) name6456 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7806_
	);
	LUT4 #(
		.INIT('h153f)
	) name6457 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7807_
	);
	LUT4 #(
		.INIT('h135f)
	) name6458 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7808_
	);
	LUT4 #(
		.INIT('h8000)
	) name6459 (
		_w7807_,
		_w7808_,
		_w7805_,
		_w7806_,
		_w7809_
	);
	LUT4 #(
		.INIT('h153f)
	) name6460 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7810_
	);
	LUT4 #(
		.INIT('h135f)
	) name6461 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7811_
	);
	LUT4 #(
		.INIT('h153f)
	) name6462 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7812_
	);
	LUT4 #(
		.INIT('h135f)
	) name6463 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7813_
	);
	LUT4 #(
		.INIT('h8000)
	) name6464 (
		_w7812_,
		_w7813_,
		_w7810_,
		_w7811_,
		_w7814_
	);
	LUT4 #(
		.INIT('h0777)
	) name6465 (
		_w7799_,
		_w7804_,
		_w7809_,
		_w7814_,
		_w7815_
	);
	LUT4 #(
		.INIT('h135f)
	) name6466 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[2][1]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7816_
	);
	LUT4 #(
		.INIT('h135f)
	) name6467 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		\P2_InstQueue_reg[15][1]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7817_
	);
	LUT4 #(
		.INIT('h153f)
	) name6468 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7818_
	);
	LUT4 #(
		.INIT('h135f)
	) name6469 (
		\P2_InstQueue_reg[3][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7819_
	);
	LUT4 #(
		.INIT('h8000)
	) name6470 (
		_w7818_,
		_w7819_,
		_w7816_,
		_w7817_,
		_w7820_
	);
	LUT4 #(
		.INIT('h153f)
	) name6471 (
		\P2_InstQueue_reg[1][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7821_
	);
	LUT4 #(
		.INIT('h135f)
	) name6472 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7822_
	);
	LUT4 #(
		.INIT('h153f)
	) name6473 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7823_
	);
	LUT4 #(
		.INIT('h135f)
	) name6474 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7824_
	);
	LUT4 #(
		.INIT('h8000)
	) name6475 (
		_w7823_,
		_w7824_,
		_w7821_,
		_w7822_,
		_w7825_
	);
	LUT2 #(
		.INIT('h8)
	) name6476 (
		_w7820_,
		_w7825_,
		_w7826_
	);
	LUT4 #(
		.INIT('h135f)
	) name6477 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7827_
	);
	LUT4 #(
		.INIT('h135f)
	) name6478 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[15][2]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7828_
	);
	LUT4 #(
		.INIT('h153f)
	) name6479 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7829_
	);
	LUT4 #(
		.INIT('h135f)
	) name6480 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7830_
	);
	LUT4 #(
		.INIT('h8000)
	) name6481 (
		_w7829_,
		_w7830_,
		_w7827_,
		_w7828_,
		_w7831_
	);
	LUT4 #(
		.INIT('h153f)
	) name6482 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7832_
	);
	LUT4 #(
		.INIT('h135f)
	) name6483 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7833_
	);
	LUT4 #(
		.INIT('h153f)
	) name6484 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7834_
	);
	LUT4 #(
		.INIT('h135f)
	) name6485 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7835_
	);
	LUT4 #(
		.INIT('h8000)
	) name6486 (
		_w7834_,
		_w7835_,
		_w7832_,
		_w7833_,
		_w7836_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		_w7831_,
		_w7836_,
		_w7837_
	);
	LUT3 #(
		.INIT('h02)
	) name6488 (
		_w7815_,
		_w7826_,
		_w7837_,
		_w7838_
	);
	LUT4 #(
		.INIT('h135f)
	) name6489 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7839_
	);
	LUT4 #(
		.INIT('h135f)
	) name6490 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[15][3]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7840_
	);
	LUT4 #(
		.INIT('h153f)
	) name6491 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7841_
	);
	LUT4 #(
		.INIT('h135f)
	) name6492 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7842_
	);
	LUT4 #(
		.INIT('h8000)
	) name6493 (
		_w7841_,
		_w7842_,
		_w7839_,
		_w7840_,
		_w7843_
	);
	LUT4 #(
		.INIT('h153f)
	) name6494 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7844_
	);
	LUT4 #(
		.INIT('h135f)
	) name6495 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7845_
	);
	LUT4 #(
		.INIT('h153f)
	) name6496 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7846_
	);
	LUT4 #(
		.INIT('h135f)
	) name6497 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7847_
	);
	LUT4 #(
		.INIT('h8000)
	) name6498 (
		_w7846_,
		_w7847_,
		_w7844_,
		_w7845_,
		_w7848_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		_w7843_,
		_w7848_,
		_w7849_
	);
	LUT4 #(
		.INIT('h0002)
	) name6500 (
		_w7815_,
		_w7826_,
		_w7837_,
		_w7849_,
		_w7850_
	);
	LUT4 #(
		.INIT('h135f)
	) name6501 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[2][4]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7851_
	);
	LUT4 #(
		.INIT('h135f)
	) name6502 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7852_
	);
	LUT4 #(
		.INIT('h153f)
	) name6503 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7853_
	);
	LUT4 #(
		.INIT('h135f)
	) name6504 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7854_
	);
	LUT4 #(
		.INIT('h8000)
	) name6505 (
		_w7853_,
		_w7854_,
		_w7851_,
		_w7852_,
		_w7855_
	);
	LUT4 #(
		.INIT('h153f)
	) name6506 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7856_
	);
	LUT4 #(
		.INIT('h135f)
	) name6507 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7857_
	);
	LUT4 #(
		.INIT('h153f)
	) name6508 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7858_
	);
	LUT4 #(
		.INIT('h135f)
	) name6509 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7859_
	);
	LUT4 #(
		.INIT('h8000)
	) name6510 (
		_w7858_,
		_w7859_,
		_w7856_,
		_w7857_,
		_w7860_
	);
	LUT2 #(
		.INIT('h8)
	) name6511 (
		_w7855_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h135f)
	) name6512 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7862_
	);
	LUT4 #(
		.INIT('h135f)
	) name6513 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[15][5]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7863_
	);
	LUT4 #(
		.INIT('h153f)
	) name6514 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7864_
	);
	LUT4 #(
		.INIT('h135f)
	) name6515 (
		\P2_InstQueue_reg[3][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7865_
	);
	LUT4 #(
		.INIT('h8000)
	) name6516 (
		_w7864_,
		_w7865_,
		_w7862_,
		_w7863_,
		_w7866_
	);
	LUT4 #(
		.INIT('h153f)
	) name6517 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7867_
	);
	LUT4 #(
		.INIT('h135f)
	) name6518 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7868_
	);
	LUT4 #(
		.INIT('h153f)
	) name6519 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7869_
	);
	LUT4 #(
		.INIT('h135f)
	) name6520 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7870_
	);
	LUT4 #(
		.INIT('h8000)
	) name6521 (
		_w7869_,
		_w7870_,
		_w7867_,
		_w7868_,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		_w7866_,
		_w7871_,
		_w7872_
	);
	LUT3 #(
		.INIT('h02)
	) name6523 (
		_w7850_,
		_w7861_,
		_w7872_,
		_w7873_
	);
	LUT4 #(
		.INIT('h135f)
	) name6524 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1447_,
		_w1457_,
		_w7874_
	);
	LUT4 #(
		.INIT('h135f)
	) name6525 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1443_,
		_w1459_,
		_w7875_
	);
	LUT4 #(
		.INIT('h153f)
	) name6526 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1446_,
		_w1456_,
		_w7876_
	);
	LUT4 #(
		.INIT('h135f)
	) name6527 (
		\P2_InstQueue_reg[3][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7877_
	);
	LUT4 #(
		.INIT('h8000)
	) name6528 (
		_w7876_,
		_w7877_,
		_w7874_,
		_w7875_,
		_w7878_
	);
	LUT4 #(
		.INIT('h153f)
	) name6529 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7879_
	);
	LUT4 #(
		.INIT('h135f)
	) name6530 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7880_
	);
	LUT4 #(
		.INIT('h153f)
	) name6531 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7881_
	);
	LUT4 #(
		.INIT('h135f)
	) name6532 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7882_
	);
	LUT4 #(
		.INIT('h8000)
	) name6533 (
		_w7881_,
		_w7882_,
		_w7879_,
		_w7880_,
		_w7883_
	);
	LUT2 #(
		.INIT('h8)
	) name6534 (
		_w7878_,
		_w7883_,
		_w7884_
	);
	LUT4 #(
		.INIT('h0002)
	) name6535 (
		_w7850_,
		_w7861_,
		_w7872_,
		_w7884_,
		_w7885_
	);
	LUT4 #(
		.INIT('h153f)
	) name6536 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1446_,
		_w1457_,
		_w7886_
	);
	LUT4 #(
		.INIT('h153f)
	) name6537 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[14][7]/NET0131 ,
		_w1443_,
		_w1447_,
		_w7887_
	);
	LUT4 #(
		.INIT('h135f)
	) name6538 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[15][7]/NET0131 ,
		_w1456_,
		_w1459_,
		_w7888_
	);
	LUT4 #(
		.INIT('h135f)
	) name6539 (
		\P2_InstQueue_reg[3][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1453_,
		_w1463_,
		_w7889_
	);
	LUT4 #(
		.INIT('h8000)
	) name6540 (
		_w7888_,
		_w7889_,
		_w7886_,
		_w7887_,
		_w7890_
	);
	LUT4 #(
		.INIT('h153f)
	) name6541 (
		\P2_InstQueue_reg[1][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1450_,
		_w1460_,
		_w7891_
	);
	LUT4 #(
		.INIT('h135f)
	) name6542 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1465_,
		_w1466_,
		_w7892_
	);
	LUT4 #(
		.INIT('h153f)
	) name6543 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1449_,
		_w1452_,
		_w7893_
	);
	LUT4 #(
		.INIT('h135f)
	) name6544 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1444_,
		_w1462_,
		_w7894_
	);
	LUT4 #(
		.INIT('h8000)
	) name6545 (
		_w7893_,
		_w7894_,
		_w7891_,
		_w7892_,
		_w7895_
	);
	LUT2 #(
		.INIT('h8)
	) name6546 (
		_w7890_,
		_w7895_,
		_w7896_
	);
	LUT4 #(
		.INIT('h0111)
	) name6547 (
		_w1592_,
		_w1595_,
		_w7890_,
		_w7895_,
		_w7897_
	);
	LUT3 #(
		.INIT('h80)
	) name6548 (
		_w1549_,
		_w1553_,
		_w7897_,
		_w7898_
	);
	LUT2 #(
		.INIT('h8)
	) name6549 (
		_w7885_,
		_w7898_,
		_w7899_
	);
	LUT3 #(
		.INIT('h07)
	) name6550 (
		_w7788_,
		_w7794_,
		_w7899_,
		_w7900_
	);
	LUT4 #(
		.INIT('hecee)
	) name6551 (
		_w1678_,
		_w7768_,
		_w7793_,
		_w7900_,
		_w7901_
	);
	LUT3 #(
		.INIT('h08)
	) name6552 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7902_
	);
	LUT4 #(
		.INIT('h1555)
	) name6553 (
		_w4261_,
		_w4231_,
		_w4244_,
		_w4258_,
		_w7903_
	);
	LUT3 #(
		.INIT('ha8)
	) name6554 (
		_w4214_,
		_w4862_,
		_w7903_,
		_w7904_
	);
	LUT4 #(
		.INIT('h4015)
	) name6555 (
		_w4214_,
		_w4339_,
		_w4348_,
		_w4349_,
		_w7905_
	);
	LUT2 #(
		.INIT('h1)
	) name6556 (
		_w1661_,
		_w7905_,
		_w7906_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6557 (
		_w1559_,
		_w7902_,
		_w7904_,
		_w7906_,
		_w7907_
	);
	LUT4 #(
		.INIT('h028a)
	) name6558 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7908_
	);
	LUT3 #(
		.INIT('h28)
	) name6559 (
		_w1659_,
		_w4417_,
		_w4418_,
		_w7909_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6560 (
		_w1659_,
		_w4417_,
		_w4418_,
		_w7908_,
		_w7910_
	);
	LUT3 #(
		.INIT('h08)
	) name6561 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w6857_,
		_w7911_
	);
	LUT3 #(
		.INIT('h48)
	) name6562 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w1679_,
		_w7911_,
		_w7912_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6563 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w5733_,
		_w7913_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6564 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7914_
	);
	LUT3 #(
		.INIT('h70)
	) name6565 (
		_w2283_,
		_w7913_,
		_w7914_,
		_w7915_
	);
	LUT2 #(
		.INIT('h4)
	) name6566 (
		_w7912_,
		_w7915_,
		_w7916_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6567 (
		_w1678_,
		_w7907_,
		_w7910_,
		_w7916_,
		_w7917_
	);
	LUT3 #(
		.INIT('h08)
	) name6568 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w1592_,
		_w1660_,
		_w7918_
	);
	LUT4 #(
		.INIT('haa20)
	) name6569 (
		_w1559_,
		_w5436_,
		_w5437_,
		_w7918_,
		_w7919_
	);
	LUT4 #(
		.INIT('h028a)
	) name6570 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7920_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6571 (
		_w1659_,
		_w4422_,
		_w4428_,
		_w7920_,
		_w7921_
	);
	LUT3 #(
		.INIT('h6a)
	) name6572 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5736_,
		_w5742_,
		_w7922_
	);
	LUT4 #(
		.INIT('h6a00)
	) name6573 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5736_,
		_w5742_,
		_w5746_,
		_w7923_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6574 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w2242_,
		_w5736_,
		_w7924_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6575 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7925_
	);
	LUT3 #(
		.INIT('h10)
	) name6576 (
		_w7924_,
		_w7923_,
		_w7925_,
		_w7926_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6577 (
		_w1678_,
		_w7919_,
		_w7921_,
		_w7926_,
		_w7927_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name6578 (
		_w4283_,
		_w4311_,
		_w4315_,
		_w4824_,
		_w7928_
	);
	LUT4 #(
		.INIT('h0015)
	) name6579 (
		_w4214_,
		_w4315_,
		_w4818_,
		_w7928_,
		_w7929_
	);
	LUT3 #(
		.INIT('h82)
	) name6580 (
		_w4214_,
		_w4223_,
		_w4807_,
		_w7930_
	);
	LUT4 #(
		.INIT('h4447)
	) name6581 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w1661_,
		_w7929_,
		_w7930_,
		_w7931_
	);
	LUT4 #(
		.INIT('h028a)
	) name6582 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w7932_
	);
	LUT4 #(
		.INIT('ha082)
	) name6583 (
		_w1659_,
		_w4401_,
		_w4403_,
		_w4869_,
		_w7933_
	);
	LUT2 #(
		.INIT('h1)
	) name6584 (
		_w7932_,
		_w7933_,
		_w7934_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6585 (
		_w1559_,
		_w1678_,
		_w7931_,
		_w7934_,
		_w7935_
	);
	LUT3 #(
		.INIT('h80)
	) name6586 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5723_,
		_w7936_
	);
	LUT4 #(
		.INIT('h8000)
	) name6587 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5723_,
		_w7937_
	);
	LUT2 #(
		.INIT('h6)
	) name6588 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w7937_,
		_w7938_
	);
	LUT3 #(
		.INIT('h48)
	) name6589 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w5746_,
		_w7937_,
		_w7939_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6590 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w2286_,
		_w5747_,
		_w7940_
	);
	LUT4 #(
		.INIT('hb700)
	) name6591 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w2242_,
		_w5724_,
		_w7940_,
		_w7941_
	);
	LUT2 #(
		.INIT('h4)
	) name6592 (
		_w7939_,
		_w7941_,
		_w7942_
	);
	LUT2 #(
		.INIT('hb)
	) name6593 (
		_w7935_,
		_w7942_,
		_w7943_
	);
	LUT3 #(
		.INIT('h02)
	) name6594 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7944_
	);
	LUT3 #(
		.INIT('ha8)
	) name6595 (
		_w2171_,
		_w5799_,
		_w7944_,
		_w7945_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6596 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7946_
	);
	LUT3 #(
		.INIT('h0b)
	) name6597 (
		_w5790_,
		_w5792_,
		_w7946_,
		_w7947_
	);
	LUT3 #(
		.INIT('h6a)
	) name6598 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5762_,
		_w7948_
	);
	LUT4 #(
		.INIT('h4111)
	) name6599 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5762_,
		_w7949_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6600 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2194_,
		_w5762_,
		_w7950_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6601 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w3055_,
		_w5762_,
		_w7951_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6602 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7952_
	);
	LUT4 #(
		.INIT('h4500)
	) name6603 (
		_w7951_,
		_w7949_,
		_w7950_,
		_w7952_,
		_w7953_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6604 (
		_w1945_,
		_w7945_,
		_w7947_,
		_w7953_,
		_w7954_
	);
	LUT3 #(
		.INIT('h02)
	) name6605 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2103_,
		_w2172_,
		_w7955_
	);
	LUT4 #(
		.INIT('h4105)
	) name6606 (
		_w2755_,
		_w2879_,
		_w2883_,
		_w2874_,
		_w7956_
	);
	LUT2 #(
		.INIT('h1)
	) name6607 (
		_w5357_,
		_w5358_,
		_w7957_
	);
	LUT3 #(
		.INIT('h20)
	) name6608 (
		_w2943_,
		_w4051_,
		_w4054_,
		_w7958_
	);
	LUT4 #(
		.INIT('h1115)
	) name6609 (
		_w2173_,
		_w2755_,
		_w7957_,
		_w7958_,
		_w7959_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6610 (
		_w2171_,
		_w7955_,
		_w7956_,
		_w7959_,
		_w7960_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6611 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w7961_
	);
	LUT3 #(
		.INIT('h6a)
	) name6612 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2733_,
		_w2986_,
		_w7962_
	);
	LUT4 #(
		.INIT('h0057)
	) name6613 (
		_w2990_,
		_w2993_,
		_w3020_,
		_w7962_,
		_w7963_
	);
	LUT4 #(
		.INIT('h222a)
	) name6614 (
		_w2181_,
		_w2991_,
		_w2993_,
		_w3020_,
		_w7964_
	);
	LUT2 #(
		.INIT('h4)
	) name6615 (
		_w7963_,
		_w7964_,
		_w7965_
	);
	LUT3 #(
		.INIT('h45)
	) name6616 (
		_w7961_,
		_w7963_,
		_w7964_,
		_w7966_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6617 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5762_,
		_w7967_
	);
	LUT2 #(
		.INIT('h8)
	) name6618 (
		_w3055_,
		_w7967_,
		_w7968_
	);
	LUT4 #(
		.INIT('h3313)
	) name6619 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w5762_,
		_w6938_,
		_w7969_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6620 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7970_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6621 (
		_w2194_,
		_w7447_,
		_w7969_,
		_w7970_,
		_w7971_
	);
	LUT2 #(
		.INIT('h4)
	) name6622 (
		_w7968_,
		_w7971_,
		_w7972_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6623 (
		_w1945_,
		_w7960_,
		_w7966_,
		_w7972_,
		_w7973_
	);
	LUT4 #(
		.INIT('h3133)
	) name6624 (
		_w2943_,
		_w2949_,
		_w4051_,
		_w4054_,
		_w7974_
	);
	LUT3 #(
		.INIT('ha8)
	) name6625 (
		_w2755_,
		_w2953_,
		_w7974_,
		_w7975_
	);
	LUT3 #(
		.INIT('h2a)
	) name6626 (
		_w2881_,
		_w4074_,
		_w4777_,
		_w7976_
	);
	LUT3 #(
		.INIT('h15)
	) name6627 (
		_w2755_,
		_w2874_,
		_w2884_,
		_w7977_
	);
	LUT3 #(
		.INIT('h45)
	) name6628 (
		_w2173_,
		_w7976_,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h2)
	) name6629 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w7422_,
		_w7979_
	);
	LUT4 #(
		.INIT('ha028)
	) name6630 (
		_w2181_,
		_w2991_,
		_w3023_,
		_w4088_,
		_w7980_
	);
	LUT2 #(
		.INIT('h1)
	) name6631 (
		_w7979_,
		_w7980_,
		_w7981_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6632 (
		_w2171_,
		_w7975_,
		_w7978_,
		_w7981_,
		_w7982_
	);
	LUT3 #(
		.INIT('h48)
	) name6633 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2194_,
		_w7447_,
		_w7983_
	);
	LUT2 #(
		.INIT('h6)
	) name6634 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w7441_,
		_w7984_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6635 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w3054_,
		_w5783_,
		_w7985_
	);
	LUT4 #(
		.INIT('hb700)
	) name6636 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w3055_,
		_w7441_,
		_w7985_,
		_w7986_
	);
	LUT2 #(
		.INIT('h4)
	) name6637 (
		_w7983_,
		_w7986_,
		_w7987_
	);
	LUT3 #(
		.INIT('h2f)
	) name6638 (
		_w1945_,
		_w7982_,
		_w7987_,
		_w7988_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6639 (
		_w2886_,
		_w4065_,
		_w4068_,
		_w4074_,
		_w7989_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name6640 (
		_w2955_,
		_w4051_,
		_w4054_,
		_w4056_,
		_w7990_
	);
	LUT4 #(
		.INIT('h5410)
	) name6641 (
		_w2173_,
		_w2755_,
		_w7989_,
		_w7990_,
		_w7991_
	);
	LUT2 #(
		.INIT('h2)
	) name6642 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w7422_,
		_w7992_
	);
	LUT3 #(
		.INIT('h6c)
	) name6643 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w3022_,
		_w7993_
	);
	LUT4 #(
		.INIT('h0080)
	) name6644 (
		\P3_InstAddrPointer_reg[15]/NET0131 ,
		_w2991_,
		_w3023_,
		_w4088_,
		_w7994_
	);
	LUT4 #(
		.INIT('haa2a)
	) name6645 (
		_w2181_,
		_w2991_,
		_w3024_,
		_w4088_,
		_w7995_
	);
	LUT3 #(
		.INIT('he0)
	) name6646 (
		_w7993_,
		_w7994_,
		_w7995_,
		_w7996_
	);
	LUT4 #(
		.INIT('h0155)
	) name6647 (
		_w7992_,
		_w7993_,
		_w7994_,
		_w7995_,
		_w7997_
	);
	LUT4 #(
		.INIT('h80aa)
	) name6648 (
		_w1945_,
		_w2171_,
		_w7991_,
		_w7997_,
		_w7998_
	);
	LUT3 #(
		.INIT('h15)
	) name6649 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w7443_,
		_w7999_
	);
	LUT2 #(
		.INIT('h8)
	) name6650 (
		_w5765_,
		_w7441_,
		_w8000_
	);
	LUT2 #(
		.INIT('h1)
	) name6651 (
		_w7999_,
		_w8000_,
		_w8001_
	);
	LUT3 #(
		.INIT('h02)
	) name6652 (
		_w6350_,
		_w7999_,
		_w8000_,
		_w8002_
	);
	LUT4 #(
		.INIT('h4888)
	) name6653 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2199_,
		_w5763_,
		_w5764_,
		_w8003_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6654 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8004_
	);
	LUT2 #(
		.INIT('h4)
	) name6655 (
		_w8003_,
		_w8004_,
		_w8005_
	);
	LUT2 #(
		.INIT('h4)
	) name6656 (
		_w8002_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('hb)
	) name6657 (
		_w7998_,
		_w8006_,
		_w8007_
	);
	LUT3 #(
		.INIT('h6a)
	) name6658 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2707_,
		_w2893_,
		_w8008_
	);
	LUT4 #(
		.INIT('h888a)
	) name6659 (
		_w2755_,
		_w2960_,
		_w4772_,
		_w8008_,
		_w8009_
	);
	LUT4 #(
		.INIT('h4000)
	) name6660 (
		_w2896_,
		_w4074_,
		_w4776_,
		_w4777_,
		_w8010_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6661 (
		_w2896_,
		_w4074_,
		_w4776_,
		_w4777_,
		_w8011_
	);
	LUT3 #(
		.INIT('h01)
	) name6662 (
		_w2755_,
		_w8011_,
		_w8010_,
		_w8012_
	);
	LUT3 #(
		.INIT('h02)
	) name6663 (
		_w2180_,
		_w8009_,
		_w8012_,
		_w8013_
	);
	LUT2 #(
		.INIT('h2)
	) name6664 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w7422_,
		_w8014_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6665 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2706_,
		_w3022_,
		_w8015_
	);
	LUT4 #(
		.INIT('h4448)
	) name6666 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2181_,
		_w3026_,
		_w7463_,
		_w8016_
	);
	LUT2 #(
		.INIT('h1)
	) name6667 (
		_w8014_,
		_w8016_,
		_w8017_
	);
	LUT3 #(
		.INIT('h80)
	) name6668 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5766_,
		_w8018_
	);
	LUT4 #(
		.INIT('h8000)
	) name6669 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5766_,
		_w8019_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6670 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5766_,
		_w8020_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6671 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2199_,
		_w5766_,
		_w8021_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6672 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8022_
	);
	LUT4 #(
		.INIT('h1300)
	) name6673 (
		_w6350_,
		_w8021_,
		_w8020_,
		_w8022_,
		_w8023_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6674 (
		_w1945_,
		_w8013_,
		_w8017_,
		_w8023_,
		_w8024_
	);
	LUT4 #(
		.INIT('h4447)
	) name6675 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w2173_,
		_w5352_,
		_w5364_,
		_w8025_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6676 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w8026_
	);
	LUT2 #(
		.INIT('h1)
	) name6677 (
		_w5366_,
		_w8026_,
		_w8027_
	);
	LUT4 #(
		.INIT('h08aa)
	) name6678 (
		_w1945_,
		_w2171_,
		_w8025_,
		_w8027_,
		_w8028_
	);
	LUT4 #(
		.INIT('h0080)
	) name6679 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5766_,
		_w5769_,
		_w6938_,
		_w8029_
	);
	LUT2 #(
		.INIT('h1)
	) name6680 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w8029_,
		_w8030_
	);
	LUT3 #(
		.INIT('ha2)
	) name6681 (
		_w2194_,
		_w5771_,
		_w6938_,
		_w8031_
	);
	LUT3 #(
		.INIT('h6c)
	) name6682 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w5770_,
		_w8032_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6683 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		_w3055_,
		_w5770_,
		_w8033_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6684 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8034_
	);
	LUT4 #(
		.INIT('h4500)
	) name6685 (
		_w8033_,
		_w8030_,
		_w8031_,
		_w8034_,
		_w8035_
	);
	LUT2 #(
		.INIT('hb)
	) name6686 (
		_w8028_,
		_w8035_,
		_w8036_
	);
	LUT3 #(
		.INIT('h02)
	) name6687 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w2103_,
		_w2172_,
		_w8037_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6688 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w8038_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6689 (
		_w2181_,
		_w3037_,
		_w3039_,
		_w8038_,
		_w8039_
	);
	LUT4 #(
		.INIT('h5700)
	) name6690 (
		_w2171_,
		_w5388_,
		_w8037_,
		_w8039_,
		_w8040_
	);
	LUT3 #(
		.INIT('h0e)
	) name6691 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w7495_,
		_w7512_,
		_w8041_
	);
	LUT4 #(
		.INIT('h60a0)
	) name6692 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w5772_,
		_w6350_,
		_w6941_,
		_w8042_
	);
	LUT4 #(
		.INIT('h1333)
	) name6693 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		_w5771_,
		_w5772_,
		_w8043_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6694 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		_w2199_,
		_w5771_,
		_w5773_,
		_w8044_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6695 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8045_
	);
	LUT3 #(
		.INIT('hb0)
	) name6696 (
		_w8043_,
		_w8044_,
		_w8045_,
		_w8046_
	);
	LUT2 #(
		.INIT('h4)
	) name6697 (
		_w8042_,
		_w8046_,
		_w8047_
	);
	LUT3 #(
		.INIT('h2f)
	) name6698 (
		_w1945_,
		_w8040_,
		_w8047_,
		_w8048_
	);
	LUT4 #(
		.INIT('h2022)
	) name6699 (
		_w2171_,
		_w2173_,
		_w5815_,
		_w5819_,
		_w8049_
	);
	LUT2 #(
		.INIT('h2)
	) name6700 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w7422_,
		_w8050_
	);
	LUT4 #(
		.INIT('h007d)
	) name6701 (
		_w2181_,
		_w2988_,
		_w4088_,
		_w8050_,
		_w8051_
	);
	LUT4 #(
		.INIT('h8000)
	) name6702 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5758_,
		_w8052_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name6703 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w5759_,
		_w8052_,
		_w8053_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6704 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w5758_,
		_w8054_
	);
	LUT3 #(
		.INIT('hc4)
	) name6705 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w8054_,
		_w8055_
	);
	LUT3 #(
		.INIT('he0)
	) name6706 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8053_,
		_w8055_,
		_w8056_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6707 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8057_
	);
	LUT3 #(
		.INIT('h70)
	) name6708 (
		_w3055_,
		_w8053_,
		_w8057_,
		_w8058_
	);
	LUT2 #(
		.INIT('h4)
	) name6709 (
		_w8056_,
		_w8058_,
		_w8059_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6710 (
		_w1945_,
		_w8049_,
		_w8051_,
		_w8059_,
		_w8060_
	);
	LUT4 #(
		.INIT('h7774)
	) name6711 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1916_,
		_w5906_,
		_w5905_,
		_w8061_
	);
	LUT4 #(
		.INIT('h028a)
	) name6712 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8062_
	);
	LUT4 #(
		.INIT('h0031)
	) name6713 (
		_w1810_,
		_w5909_,
		_w8061_,
		_w8062_,
		_w8063_
	);
	LUT3 #(
		.INIT('h6c)
	) name6714 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w7530_,
		_w8064_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6715 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w3407_,
		_w7530_,
		_w8065_
	);
	LUT4 #(
		.INIT('h8848)
	) name6716 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w1939_,
		_w6368_,
		_w7041_,
		_w8066_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6717 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8067_
	);
	LUT3 #(
		.INIT('h10)
	) name6718 (
		_w8066_,
		_w8065_,
		_w8067_,
		_w8068_
	);
	LUT3 #(
		.INIT('h2f)
	) name6719 (
		_w1933_,
		_w8063_,
		_w8068_,
		_w8069_
	);
	LUT3 #(
		.INIT('h08)
	) name6720 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8070_
	);
	LUT4 #(
		.INIT('h820a)
	) name6721 (
		_w3101_,
		_w3296_,
		_w3302_,
		_w3993_,
		_w8071_
	);
	LUT4 #(
		.INIT('h4554)
	) name6722 (
		_w1916_,
		_w3101_,
		_w3219_,
		_w4010_,
		_w8072_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6723 (
		_w1810_,
		_w8070_,
		_w8071_,
		_w8072_,
		_w8073_
	);
	LUT3 #(
		.INIT('h6c)
	) name6724 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w3361_,
		_w8074_
	);
	LUT4 #(
		.INIT('h0800)
	) name6725 (
		\P1_InstAddrPointer_reg[12]/NET0131 ,
		_w3362_,
		_w4023_,
		_w4025_,
		_w8075_
	);
	LUT3 #(
		.INIT('h28)
	) name6726 (
		_w1924_,
		_w8074_,
		_w8075_,
		_w8076_
	);
	LUT4 #(
		.INIT('h028a)
	) name6727 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8077_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6728 (
		_w1924_,
		_w8074_,
		_w8075_,
		_w8077_,
		_w8078_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6729 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w7530_,
		_w8079_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6730 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w2310_,
		_w6368_,
		_w8080_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6731 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8081_
	);
	LUT4 #(
		.INIT('h1300)
	) name6732 (
		_w6378_,
		_w8080_,
		_w8079_,
		_w8081_,
		_w8082_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6733 (
		_w1933_,
		_w8073_,
		_w8078_,
		_w8082_,
		_w8083_
	);
	LUT3 #(
		.INIT('h08)
	) name6734 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8084_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6735 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w3060_,
		_w3063_,
		_w3067_,
		_w8085_
	);
	LUT4 #(
		.INIT('h007f)
	) name6736 (
		_w3296_,
		_w3302_,
		_w3993_,
		_w8085_,
		_w8086_
	);
	LUT3 #(
		.INIT('ha8)
	) name6737 (
		_w3101_,
		_w7540_,
		_w8086_,
		_w8087_
	);
	LUT4 #(
		.INIT('h4554)
	) name6738 (
		_w1916_,
		_w3101_,
		_w3224_,
		_w3254_,
		_w8088_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6739 (
		_w1810_,
		_w8084_,
		_w8087_,
		_w8088_,
		_w8089_
	);
	LUT3 #(
		.INIT('h28)
	) name6740 (
		_w1924_,
		_w3364_,
		_w3369_,
		_w8090_
	);
	LUT4 #(
		.INIT('h028a)
	) name6741 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8091_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6742 (
		_w1924_,
		_w3364_,
		_w3369_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h6)
	) name6743 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w7551_,
		_w8093_
	);
	LUT3 #(
		.INIT('h48)
	) name6744 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w6378_,
		_w7551_,
		_w8094_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6745 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8095_
	);
	LUT4 #(
		.INIT('hb700)
	) name6746 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w2310_,
		_w6369_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h4)
	) name6747 (
		_w8094_,
		_w8096_,
		_w8097_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6748 (
		_w1933_,
		_w8089_,
		_w8092_,
		_w8097_,
		_w8098_
	);
	LUT3 #(
		.INIT('h08)
	) name6749 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8099_
	);
	LUT4 #(
		.INIT('h8222)
	) name6750 (
		_w3101_,
		_w3297_,
		_w4463_,
		_w4465_,
		_w8100_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6751 (
		_w3246_,
		_w4724_,
		_w4725_,
		_w4727_,
		_w8101_
	);
	LUT4 #(
		.INIT('h0054)
	) name6752 (
		_w1916_,
		_w3101_,
		_w8101_,
		_w8100_,
		_w8102_
	);
	LUT3 #(
		.INIT('h28)
	) name6753 (
		_w1924_,
		_w3368_,
		_w4735_,
		_w8103_
	);
	LUT4 #(
		.INIT('h028a)
	) name6754 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8104_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6755 (
		_w1924_,
		_w3368_,
		_w4735_,
		_w8104_,
		_w8105_
	);
	LUT4 #(
		.INIT('h5700)
	) name6756 (
		_w1810_,
		_w8099_,
		_w8102_,
		_w8105_,
		_w8106_
	);
	LUT4 #(
		.INIT('h0080)
	) name6757 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w6370_,
		_w7041_,
		_w8107_
	);
	LUT4 #(
		.INIT('h3313)
	) name6758 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w6370_,
		_w7041_,
		_w8108_
	);
	LUT3 #(
		.INIT('h02)
	) name6759 (
		_w1939_,
		_w8108_,
		_w8107_,
		_w8109_
	);
	LUT4 #(
		.INIT('h070f)
	) name6760 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w7551_,
		_w8110_
	);
	LUT2 #(
		.INIT('h1)
	) name6761 (
		_w6372_,
		_w8110_,
		_w8111_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6762 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8112_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6763 (
		_w3407_,
		_w6372_,
		_w8110_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h4)
	) name6764 (
		_w8109_,
		_w8113_,
		_w8114_
	);
	LUT3 #(
		.INIT('h2f)
	) name6765 (
		_w1933_,
		_w8106_,
		_w8114_,
		_w8115_
	);
	LUT4 #(
		.INIT('h4447)
	) name6766 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w1916_,
		_w5920_,
		_w5921_,
		_w8116_
	);
	LUT4 #(
		.INIT('h028a)
	) name6767 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8117_
	);
	LUT4 #(
		.INIT('h0031)
	) name6768 (
		_w1810_,
		_w5925_,
		_w8116_,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h6)
	) name6769 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6372_,
		_w8119_
	);
	LUT3 #(
		.INIT('h60)
	) name6770 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6372_,
		_w6378_,
		_w8120_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6771 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8121_
	);
	LUT4 #(
		.INIT('hb700)
	) name6772 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w2310_,
		_w6371_,
		_w8121_,
		_w8122_
	);
	LUT2 #(
		.INIT('h4)
	) name6773 (
		_w8120_,
		_w8122_,
		_w8123_
	);
	LUT3 #(
		.INIT('h2f)
	) name6774 (
		_w1933_,
		_w8118_,
		_w8123_,
		_w8124_
	);
	LUT3 #(
		.INIT('h08)
	) name6775 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8125_
	);
	LUT4 #(
		.INIT('h004f)
	) name6776 (
		_w5454_,
		_w5456_,
		_w5459_,
		_w8125_,
		_w8126_
	);
	LUT4 #(
		.INIT('h028a)
	) name6777 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8127_
	);
	LUT2 #(
		.INIT('h1)
	) name6778 (
		_w5461_,
		_w8127_,
		_w8128_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6779 (
		_w1810_,
		_w1933_,
		_w8126_,
		_w8128_,
		_w8129_
	);
	LUT3 #(
		.INIT('h6c)
	) name6780 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w6372_,
		_w8130_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6781 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w6372_,
		_w6378_,
		_w8131_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6782 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8132_
	);
	LUT4 #(
		.INIT('hb700)
	) name6783 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w2310_,
		_w6379_,
		_w8132_,
		_w8133_
	);
	LUT2 #(
		.INIT('h4)
	) name6784 (
		_w8131_,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('hb)
	) name6785 (
		_w8129_,
		_w8134_,
		_w8135_
	);
	LUT3 #(
		.INIT('h08)
	) name6786 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8136_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name6787 (
		_w3101_,
		_w3308_,
		_w3312_,
		_w3996_,
		_w8137_
	);
	LUT4 #(
		.INIT('h4111)
	) name6788 (
		_w3101_,
		_w3235_,
		_w3255_,
		_w4011_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name6789 (
		_w1916_,
		_w8138_,
		_w8139_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6790 (
		_w1810_,
		_w8136_,
		_w8137_,
		_w8139_,
		_w8140_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6791 (
		\P1_InstAddrPointer_reg[20]/NET0131 ,
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w3074_,
		_w3366_,
		_w8141_
	);
	LUT3 #(
		.INIT('h07)
	) name6792 (
		_w4016_,
		_w4030_,
		_w8141_,
		_w8142_
	);
	LUT3 #(
		.INIT('h2a)
	) name6793 (
		_w1924_,
		_w4017_,
		_w4030_,
		_w8143_
	);
	LUT4 #(
		.INIT('h028a)
	) name6794 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8144_
	);
	LUT3 #(
		.INIT('h0b)
	) name6795 (
		_w8142_,
		_w8143_,
		_w8144_,
		_w8145_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name6796 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w6373_,
		_w7583_,
		_w8146_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6797 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w2310_,
		_w6383_,
		_w7583_,
		_w8147_
	);
	LUT3 #(
		.INIT('h20)
	) name6798 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		_w1939_,
		_w8148_
	);
	LUT2 #(
		.INIT('h8)
	) name6799 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w3406_,
		_w8149_
	);
	LUT3 #(
		.INIT('h07)
	) name6800 (
		_w7583_,
		_w8148_,
		_w8149_,
		_w8150_
	);
	LUT4 #(
		.INIT('h1300)
	) name6801 (
		_w6378_,
		_w8147_,
		_w8146_,
		_w8150_,
		_w8151_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6802 (
		_w1933_,
		_w8140_,
		_w8145_,
		_w8151_,
		_w8152_
	);
	LUT3 #(
		.INIT('h08)
	) name6803 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8153_
	);
	LUT4 #(
		.INIT('h8222)
	) name6804 (
		_w3101_,
		_w3317_,
		_w3996_,
		_w4702_,
		_w8154_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name6805 (
		_w3239_,
		_w3240_,
		_w3255_,
		_w4011_,
		_w8155_
	);
	LUT3 #(
		.INIT('h15)
	) name6806 (
		_w3101_,
		_w3256_,
		_w4011_,
		_w8156_
	);
	LUT3 #(
		.INIT('h45)
	) name6807 (
		_w1916_,
		_w8155_,
		_w8156_,
		_w8157_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6808 (
		_w1810_,
		_w8153_,
		_w8154_,
		_w8157_,
		_w8158_
	);
	LUT4 #(
		.INIT('h028a)
	) name6809 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8159_
	);
	LUT4 #(
		.INIT('h1555)
	) name6810 (
		_w3380_,
		_w3383_,
		_w4017_,
		_w4030_,
		_w8160_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6811 (
		_w1924_,
		_w3384_,
		_w4017_,
		_w4030_,
		_w8161_
	);
	LUT3 #(
		.INIT('h45)
	) name6812 (
		_w8159_,
		_w8160_,
		_w8161_,
		_w8162_
	);
	LUT4 #(
		.INIT('h070f)
	) name6813 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w7607_,
		_w8163_
	);
	LUT2 #(
		.INIT('h1)
	) name6814 (
		_w6374_,
		_w8163_,
		_w8164_
	);
	LUT3 #(
		.INIT('h04)
	) name6815 (
		_w6374_,
		_w6378_,
		_w8163_,
		_w8165_
	);
	LUT3 #(
		.INIT('ha2)
	) name6816 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		_w6383_,
		_w7619_,
		_w8166_
	);
	LUT2 #(
		.INIT('h8)
	) name6817 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w3406_,
		_w8167_
	);
	LUT4 #(
		.INIT('h007f)
	) name6818 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w7607_,
		_w7619_,
		_w8167_,
		_w8168_
	);
	LUT2 #(
		.INIT('h4)
	) name6819 (
		_w8166_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h4)
	) name6820 (
		_w8165_,
		_w8169_,
		_w8170_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6821 (
		_w1933_,
		_w8158_,
		_w8162_,
		_w8170_,
		_w8171_
	);
	LUT4 #(
		.INIT('h1500)
	) name6822 (
		_w3268_,
		_w4455_,
		_w4458_,
		_w4461_,
		_w8172_
	);
	LUT4 #(
		.INIT('h80aa)
	) name6823 (
		_w3268_,
		_w4455_,
		_w4458_,
		_w4461_,
		_w8173_
	);
	LUT3 #(
		.INIT('h02)
	) name6824 (
		_w3101_,
		_w8173_,
		_w8172_,
		_w8174_
	);
	LUT4 #(
		.INIT('h3323)
	) name6825 (
		_w3102_,
		_w3210_,
		_w4005_,
		_w4472_,
		_w8175_
	);
	LUT4 #(
		.INIT('h0015)
	) name6826 (
		_w3101_,
		_w3210_,
		_w4724_,
		_w8175_,
		_w8176_
	);
	LUT4 #(
		.INIT('h4447)
	) name6827 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w1916_,
		_w8174_,
		_w8176_,
		_w8177_
	);
	LUT3 #(
		.INIT('h82)
	) name6828 (
		_w1924_,
		_w3358_,
		_w3356_,
		_w8178_
	);
	LUT4 #(
		.INIT('h028a)
	) name6829 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8179_
	);
	LUT4 #(
		.INIT('h007d)
	) name6830 (
		_w1924_,
		_w3358_,
		_w3356_,
		_w8179_,
		_w8180_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6831 (
		_w1810_,
		_w1933_,
		_w8177_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h6)
	) name6832 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w7529_,
		_w8182_
	);
	LUT3 #(
		.INIT('h41)
	) name6833 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w7529_,
		_w8183_
	);
	LUT4 #(
		.INIT('h78f0)
	) name6834 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w6365_,
		_w8184_
	);
	LUT3 #(
		.INIT('hc4)
	) name6835 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w8184_,
		_w8185_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6836 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8186_
	);
	LUT4 #(
		.INIT('hb700)
	) name6837 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w3407_,
		_w7529_,
		_w8186_,
		_w8187_
	);
	LUT3 #(
		.INIT('hb0)
	) name6838 (
		_w8183_,
		_w8185_,
		_w8187_,
		_w8188_
	);
	LUT2 #(
		.INIT('hb)
	) name6839 (
		_w8181_,
		_w8188_,
		_w8189_
	);
	LUT3 #(
		.INIT('h08)
	) name6840 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8190_
	);
	LUT4 #(
		.INIT('haa20)
	) name6841 (
		_w1559_,
		_w5869_,
		_w5872_,
		_w8190_,
		_w8191_
	);
	LUT4 #(
		.INIT('h028a)
	) name6842 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8192_
	);
	LUT2 #(
		.INIT('h1)
	) name6843 (
		_w5876_,
		_w8192_,
		_w8193_
	);
	LUT2 #(
		.INIT('h6)
	) name6844 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w7631_,
		_w8194_
	);
	LUT3 #(
		.INIT('h48)
	) name6845 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w5746_,
		_w7631_,
		_w8195_
	);
	LUT4 #(
		.INIT('h8000)
	) name6846 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w8196_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6847 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8197_
	);
	LUT4 #(
		.INIT('hb700)
	) name6848 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w2242_,
		_w5727_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h4)
	) name6849 (
		_w8195_,
		_w8198_,
		_w8199_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6850 (
		_w1678_,
		_w8191_,
		_w8193_,
		_w8199_,
		_w8200_
	);
	LUT3 #(
		.INIT('h08)
	) name6851 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8201_
	);
	LUT4 #(
		.INIT('haa20)
	) name6852 (
		_w1559_,
		_w5887_,
		_w5890_,
		_w8201_,
		_w8202_
	);
	LUT4 #(
		.INIT('h028a)
	) name6853 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8203_
	);
	LUT3 #(
		.INIT('h0b)
	) name6854 (
		_w5892_,
		_w5893_,
		_w8203_,
		_w8204_
	);
	LUT3 #(
		.INIT('h13)
	) name6855 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w7631_,
		_w8205_
	);
	LUT4 #(
		.INIT('h8000)
	) name6856 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w5728_,
		_w8206_
	);
	LUT2 #(
		.INIT('h8)
	) name6857 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w8206_,
		_w8207_
	);
	LUT2 #(
		.INIT('h1)
	) name6858 (
		_w8205_,
		_w8207_,
		_w8208_
	);
	LUT3 #(
		.INIT('h02)
	) name6859 (
		_w2283_,
		_w8205_,
		_w8207_,
		_w8209_
	);
	LUT3 #(
		.INIT('h13)
	) name6860 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w7636_,
		_w8210_
	);
	LUT3 #(
		.INIT('h8a)
	) name6861 (
		_w1679_,
		_w6857_,
		_w8206_,
		_w8211_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6862 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8212_
	);
	LUT3 #(
		.INIT('hb0)
	) name6863 (
		_w8210_,
		_w8211_,
		_w8212_,
		_w8213_
	);
	LUT2 #(
		.INIT('h4)
	) name6864 (
		_w8209_,
		_w8213_,
		_w8214_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6865 (
		_w1678_,
		_w8202_,
		_w8204_,
		_w8214_,
		_w8215_
	);
	LUT3 #(
		.INIT('h45)
	) name6866 (
		_w4240_,
		_w4807_,
		_w4810_,
		_w8216_
	);
	LUT3 #(
		.INIT('h2a)
	) name6867 (
		_w4214_,
		_w4796_,
		_w4799_,
		_w8217_
	);
	LUT2 #(
		.INIT('h4)
	) name6868 (
		_w8216_,
		_w8217_,
		_w8218_
	);
	LUT3 #(
		.INIT('h13)
	) name6869 (
		_w4328_,
		_w4823_,
		_w5889_,
		_w8219_
	);
	LUT4 #(
		.INIT('h4744)
	) name6870 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w1661_,
		_w8218_,
		_w8219_,
		_w8220_
	);
	LUT4 #(
		.INIT('h028a)
	) name6871 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8221_
	);
	LUT4 #(
		.INIT('h0080)
	) name6872 (
		_w4405_,
		_w4409_,
		_w4411_,
		_w4869_,
		_w8222_
	);
	LUT4 #(
		.INIT('h0f07)
	) name6873 (
		_w4405_,
		_w4409_,
		_w4411_,
		_w4869_,
		_w8223_
	);
	LUT3 #(
		.INIT('h02)
	) name6874 (
		_w1659_,
		_w8223_,
		_w8222_,
		_w8224_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6875 (
		_w1659_,
		_w4411_,
		_w4870_,
		_w8221_,
		_w8225_
	);
	LUT4 #(
		.INIT('h08cc)
	) name6876 (
		_w1559_,
		_w1678_,
		_w8220_,
		_w8225_,
		_w8226_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6877 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5727_,
		_w5728_,
		_w8227_
	);
	LUT4 #(
		.INIT('h4888)
	) name6878 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w2242_,
		_w5727_,
		_w5728_,
		_w8228_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6879 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8229_
	);
	LUT4 #(
		.INIT('h1300)
	) name6880 (
		_w5746_,
		_w8228_,
		_w8227_,
		_w8229_,
		_w8230_
	);
	LUT2 #(
		.INIT('hb)
	) name6881 (
		_w8226_,
		_w8230_,
		_w8231_
	);
	LUT3 #(
		.INIT('h08)
	) name6882 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8232_
	);
	LUT3 #(
		.INIT('h32)
	) name6883 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w4247_,
		_w4794_,
		_w8233_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6884 (
		_w4241_,
		_w4807_,
		_w4810_,
		_w8233_,
		_w8234_
	);
	LUT4 #(
		.INIT('h0020)
	) name6885 (
		_w4241_,
		_w4807_,
		_w4810_,
		_w8233_,
		_w8235_
	);
	LUT3 #(
		.INIT('h02)
	) name6886 (
		_w4214_,
		_w8235_,
		_w8234_,
		_w8236_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6887 (
		_w4336_,
		_w4818_,
		_w4903_,
		_w6883_,
		_w8237_
	);
	LUT4 #(
		.INIT('h5554)
	) name6888 (
		_w1661_,
		_w4214_,
		_w4855_,
		_w8237_,
		_w8238_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6889 (
		_w1559_,
		_w8232_,
		_w8236_,
		_w8238_,
		_w8239_
	);
	LUT4 #(
		.INIT('h028a)
	) name6890 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8240_
	);
	LUT3 #(
		.INIT('h28)
	) name6891 (
		_w1659_,
		_w6897_,
		_w6898_,
		_w8241_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6892 (
		_w1659_,
		_w6897_,
		_w6898_,
		_w8240_,
		_w8242_
	);
	LUT3 #(
		.INIT('h80)
	) name6893 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w5730_,
		_w8243_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name6894 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5730_,
		_w8244_
	);
	LUT4 #(
		.INIT('h60c0)
	) name6895 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w2242_,
		_w5730_,
		_w8245_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6896 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8246_
	);
	LUT4 #(
		.INIT('h0700)
	) name6897 (
		_w5746_,
		_w8244_,
		_w8245_,
		_w8246_,
		_w8247_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6898 (
		_w1678_,
		_w8239_,
		_w8242_,
		_w8247_,
		_w8248_
	);
	LUT3 #(
		.INIT('h08)
	) name6899 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8249_
	);
	LUT4 #(
		.INIT('h802a)
	) name6900 (
		_w4214_,
		_w4231_,
		_w4244_,
		_w4251_,
		_w8250_
	);
	LUT4 #(
		.INIT('h4554)
	) name6901 (
		_w1661_,
		_w4214_,
		_w4339_,
		_w4340_,
		_w8251_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6902 (
		_w1559_,
		_w8249_,
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT4 #(
		.INIT('h028a)
	) name6903 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8253_
	);
	LUT4 #(
		.INIT('h4000)
	) name6904 (
		_w4400_,
		_w4405_,
		_w4409_,
		_w4412_,
		_w8254_
	);
	LUT3 #(
		.INIT('h28)
	) name6905 (
		_w1659_,
		_w4413_,
		_w8254_,
		_w8255_
	);
	LUT4 #(
		.INIT('h0d07)
	) name6906 (
		_w1659_,
		_w4413_,
		_w8253_,
		_w8254_,
		_w8256_
	);
	LUT4 #(
		.INIT('h8000)
	) name6907 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w5730_,
		_w8257_
	);
	LUT2 #(
		.INIT('h6)
	) name6908 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w8257_,
		_w8258_
	);
	LUT3 #(
		.INIT('h48)
	) name6909 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w5746_,
		_w8257_,
		_w8259_
	);
	LUT4 #(
		.INIT('h8000)
	) name6910 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w5730_,
		_w8260_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6911 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8261_
	);
	LUT4 #(
		.INIT('hb700)
	) name6912 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w2242_,
		_w8243_,
		_w8261_,
		_w8262_
	);
	LUT2 #(
		.INIT('h4)
	) name6913 (
		_w8259_,
		_w8262_,
		_w8263_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6914 (
		_w1678_,
		_w8252_,
		_w8256_,
		_w8263_,
		_w8264_
	);
	LUT3 #(
		.INIT('h08)
	) name6915 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8265_
	);
	LUT4 #(
		.INIT('haa20)
	) name6916 (
		_w1559_,
		_w5417_,
		_w5419_,
		_w8265_,
		_w8266_
	);
	LUT4 #(
		.INIT('h028a)
	) name6917 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8267_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6918 (
		_w1659_,
		_w4865_,
		_w4872_,
		_w8267_,
		_w8268_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name6919 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w7660_,
		_w8257_,
		_w8269_
	);
	LUT3 #(
		.INIT('h32)
	) name6920 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w5732_,
		_w8260_,
		_w8270_
	);
	LUT4 #(
		.INIT('hc840)
	) name6921 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w8269_,
		_w8270_,
		_w8271_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6922 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8272_
	);
	LUT3 #(
		.INIT('h70)
	) name6923 (
		_w2283_,
		_w8269_,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h4)
	) name6924 (
		_w8271_,
		_w8273_,
		_w8274_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6925 (
		_w1678_,
		_w8266_,
		_w8268_,
		_w8274_,
		_w8275_
	);
	LUT3 #(
		.INIT('h54)
	) name6926 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1855_,
		_w1860_,
		_w8276_
	);
	LUT4 #(
		.INIT('haa2a)
	) name6927 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w1922_,
		_w5911_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h4)
	) name6928 (
		_w1862_,
		_w3272_,
		_w8278_
	);
	LUT3 #(
		.INIT('hb0)
	) name6929 (
		_w1816_,
		_w1831_,
		_w3196_,
		_w8279_
	);
	LUT4 #(
		.INIT('h40bf)
	) name6930 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3196_,
		_w8280_
	);
	LUT4 #(
		.INIT('h4114)
	) name6931 (
		_w3101_,
		_w3195_,
		_w3170_,
		_w3196_,
		_w8281_
	);
	LUT4 #(
		.INIT('h40bf)
	) name6932 (
		_w3189_,
		_w3187_,
		_w3194_,
		_w3272_,
		_w8282_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6933 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3154_,
		_w3275_,
		_w8282_,
		_w8283_
	);
	LUT4 #(
		.INIT('h0071)
	) name6934 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3154_,
		_w3275_,
		_w8282_,
		_w8284_
	);
	LUT3 #(
		.INIT('h02)
	) name6935 (
		_w3101_,
		_w8284_,
		_w8283_,
		_w8285_
	);
	LUT3 #(
		.INIT('h04)
	) name6936 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8286_
	);
	LUT2 #(
		.INIT('h2)
	) name6937 (
		_w1810_,
		_w8286_,
		_w8287_
	);
	LUT4 #(
		.INIT('hab00)
	) name6938 (
		_w1916_,
		_w8281_,
		_w8285_,
		_w8287_,
		_w8288_
	);
	LUT4 #(
		.INIT('haaa9)
	) name6939 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		_w1842_,
		_w1845_,
		_w3083_,
		_w8289_
	);
	LUT4 #(
		.INIT('h2b00)
	) name6940 (
		_w3154_,
		_w3155_,
		_w3337_,
		_w8280_,
		_w8290_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6941 (
		_w3154_,
		_w3155_,
		_w3337_,
		_w8280_,
		_w8291_
	);
	LUT4 #(
		.INIT('h0008)
	) name6942 (
		_w1809_,
		_w1846_,
		_w8291_,
		_w8290_,
		_w8292_
	);
	LUT3 #(
		.INIT('h0b)
	) name6943 (
		_w1833_,
		_w8289_,
		_w8292_,
		_w8293_
	);
	LUT2 #(
		.INIT('h4)
	) name6944 (
		_w8288_,
		_w8293_,
		_w8294_
	);
	LUT4 #(
		.INIT('h0100)
	) name6945 (
		_w8279_,
		_w8277_,
		_w8278_,
		_w8294_,
		_w8295_
	);
	LUT2 #(
		.INIT('h8)
	) name6946 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w3406_,
		_w8296_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6947 (
		\P1_InstAddrPointer_reg[2]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w3406_,
		_w3408_,
		_w8297_
	);
	LUT3 #(
		.INIT('h2f)
	) name6948 (
		_w1933_,
		_w8295_,
		_w8297_,
		_w8298_
	);
	LUT2 #(
		.INIT('h2)
	) name6949 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		_w7103_,
		_w8299_
	);
	LUT3 #(
		.INIT('hb0)
	) name6950 (
		_w2073_,
		_w2086_,
		_w2771_,
		_w8300_
	);
	LUT2 #(
		.INIT('h4)
	) name6951 (
		_w2117_,
		_w2917_,
		_w8301_
	);
	LUT3 #(
		.INIT('h87)
	) name6952 (
		_w2763_,
		_w2768_,
		_w2771_,
		_w8302_
	);
	LUT4 #(
		.INIT('hba45)
	) name6953 (
		_w3003_,
		_w3004_,
		_w3005_,
		_w8302_,
		_w8303_
	);
	LUT3 #(
		.INIT('h80)
	) name6954 (
		_w2060_,
		_w2041_,
		_w8303_,
		_w8304_
	);
	LUT4 #(
		.INIT('h00f1)
	) name6955 (
		_w2071_,
		_w2087_,
		_w2771_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h14)
	) name6956 (
		_w2755_,
		_w2797_,
		_w8302_,
		_w8306_
	);
	LUT3 #(
		.INIT('h87)
	) name6957 (
		_w2763_,
		_w2768_,
		_w2917_,
		_w8307_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6958 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2783_,
		_w2795_,
		_w8307_,
		_w8308_
	);
	LUT4 #(
		.INIT('h0071)
	) name6959 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2783_,
		_w2795_,
		_w8307_,
		_w8309_
	);
	LUT3 #(
		.INIT('h02)
	) name6960 (
		_w2755_,
		_w8309_,
		_w8308_,
		_w8310_
	);
	LUT3 #(
		.INIT('h02)
	) name6961 (
		_w2180_,
		_w8310_,
		_w8306_,
		_w8311_
	);
	LUT3 #(
		.INIT('h0d)
	) name6962 (
		_w2098_,
		_w8305_,
		_w8311_,
		_w8312_
	);
	LUT3 #(
		.INIT('h10)
	) name6963 (
		_w8301_,
		_w8300_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w3054_,
		_w8314_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6965 (
		\P3_InstAddrPointer_reg[2]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w3054_,
		_w3056_,
		_w8315_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6966 (
		_w1945_,
		_w8299_,
		_w8313_,
		_w8315_,
		_w8316_
	);
	LUT4 #(
		.INIT('haa8a)
	) name6967 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w1626_,
		_w1643_,
		_w1667_,
		_w8317_
	);
	LUT3 #(
		.INIT('h87)
	) name6968 (
		_w4109_,
		_w4114_,
		_w4291_,
		_w8318_
	);
	LUT4 #(
		.INIT('h54ab)
	) name6969 (
		_w4294_,
		_w4389_,
		_w4390_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		_w1558_,
		_w8319_,
		_w8320_
	);
	LUT4 #(
		.INIT('h00c8)
	) name6971 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w4291_,
		_w8321_
	);
	LUT3 #(
		.INIT('ha8)
	) name6972 (
		_w1596_,
		_w8320_,
		_w8321_,
		_w8322_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		_w1563_,
		_w4115_,
		_w8323_
	);
	LUT4 #(
		.INIT('hc666)
	) name6974 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w8324_
	);
	LUT4 #(
		.INIT('hec00)
	) name6975 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w8324_,
		_w8325_
	);
	LUT4 #(
		.INIT('hccc6)
	) name6976 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w1605_,
		_w1611_,
		_w8326_
	);
	LUT4 #(
		.INIT('hdc00)
	) name6977 (
		_w1501_,
		_w1566_,
		_w1568_,
		_w8326_,
		_w8327_
	);
	LUT4 #(
		.INIT('h2223)
	) name6978 (
		_w1602_,
		_w8323_,
		_w8325_,
		_w8327_,
		_w8328_
	);
	LUT3 #(
		.INIT('h10)
	) name6979 (
		_w8317_,
		_w8322_,
		_w8328_,
		_w8329_
	);
	LUT3 #(
		.INIT('h08)
	) name6980 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8330_
	);
	LUT3 #(
		.INIT('h87)
	) name6981 (
		_w4109_,
		_w4114_,
		_w4115_,
		_w8331_
	);
	LUT4 #(
		.INIT('h8e71)
	) name6982 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4127_,
		_w4140_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h2)
	) name6983 (
		_w4214_,
		_w8332_,
		_w8333_
	);
	LUT4 #(
		.INIT('h4554)
	) name6984 (
		_w1661_,
		_w4214_,
		_w4296_,
		_w8318_,
		_w8334_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6985 (
		_w1559_,
		_w8330_,
		_w8333_,
		_w8334_,
		_w8335_
	);
	LUT4 #(
		.INIT('h004f)
	) name6986 (
		_w1571_,
		_w1583_,
		_w4291_,
		_w8335_,
		_w8336_
	);
	LUT2 #(
		.INIT('h8)
	) name6987 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w2286_,
		_w8337_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6988 (
		\P2_InstAddrPointer_reg[2]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w2286_,
		_w4441_,
		_w8338_
	);
	LUT4 #(
		.INIT('h2aff)
	) name6989 (
		_w1678_,
		_w8329_,
		_w8336_,
		_w8338_,
		_w8339_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name6990 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w8340_
	);
	LUT4 #(
		.INIT('hfc20)
	) name6991 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w8341_
	);
	LUT2 #(
		.INIT('h2)
	) name6992 (
		\P3_EAX_reg[27]/NET0131 ,
		_w8341_,
		_w8342_
	);
	LUT4 #(
		.INIT('h8000)
	) name6993 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		_w8343_
	);
	LUT4 #(
		.INIT('h8000)
	) name6994 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		\P3_EAX_reg[6]/NET0131 ,
		_w8343_,
		_w8344_
	);
	LUT4 #(
		.INIT('h8000)
	) name6995 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		\P3_EAX_reg[9]/NET0131 ,
		_w8344_,
		_w8345_
	);
	LUT2 #(
		.INIT('h8)
	) name6996 (
		\P3_EAX_reg[10]/NET0131 ,
		_w8345_,
		_w8346_
	);
	LUT3 #(
		.INIT('h80)
	) name6997 (
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		_w8345_,
		_w8347_
	);
	LUT4 #(
		.INIT('h8000)
	) name6998 (
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		\P3_EAX_reg[12]/NET0131 ,
		_w8345_,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		\P3_EAX_reg[13]/NET0131 ,
		_w8348_,
		_w8349_
	);
	LUT3 #(
		.INIT('h80)
	) name7000 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		_w8348_,
		_w8350_
	);
	LUT4 #(
		.INIT('h8000)
	) name7001 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		\P3_EAX_reg[15]/NET0131 ,
		_w8348_,
		_w8351_
	);
	LUT2 #(
		.INIT('h8)
	) name7002 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		_w8352_
	);
	LUT3 #(
		.INIT('h80)
	) name7003 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[18]/NET0131 ,
		_w8353_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		_w8351_,
		_w8353_,
		_w8354_
	);
	LUT3 #(
		.INIT('h80)
	) name7005 (
		\P3_EAX_reg[19]/NET0131 ,
		_w8351_,
		_w8353_,
		_w8355_
	);
	LUT4 #(
		.INIT('h8000)
	) name7006 (
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		_w8351_,
		_w8353_,
		_w8356_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		_w8357_
	);
	LUT3 #(
		.INIT('h80)
	) name7008 (
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		_w8358_
	);
	LUT4 #(
		.INIT('h8000)
	) name7009 (
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		\P3_EAX_reg[24]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		_w8359_
	);
	LUT3 #(
		.INIT('h80)
	) name7010 (
		\P3_EAX_reg[21]/NET0131 ,
		_w8356_,
		_w8359_,
		_w8360_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		_w2063_,
		_w2075_,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name7012 (
		\P3_EAX_reg[26]/NET0131 ,
		\P3_EAX_reg[27]/NET0131 ,
		_w8362_
	);
	LUT4 #(
		.INIT('h8000)
	) name7013 (
		\P3_EAX_reg[21]/NET0131 ,
		_w8356_,
		_w8359_,
		_w8362_,
		_w8363_
	);
	LUT2 #(
		.INIT('h2)
	) name7014 (
		_w8361_,
		_w8363_,
		_w8364_
	);
	LUT4 #(
		.INIT('h60c0)
	) name7015 (
		\P3_EAX_reg[26]/NET0131 ,
		\P3_EAX_reg[27]/NET0131 ,
		_w8361_,
		_w8360_,
		_w8365_
	);
	LUT4 #(
		.INIT('h0800)
	) name7016 (
		_w2068_,
		_w2061_,
		_w2039_,
		_w2098_,
		_w8366_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name7017 (
		_w2107_,
		_w2087_,
		_w8366_,
		_w8361_,
		_w8367_
	);
	LUT3 #(
		.INIT('h01)
	) name7018 (
		\buf2_reg[27]/NET0131 ,
		_w2105_,
		_w2116_,
		_w8368_
	);
	LUT3 #(
		.INIT('h54)
	) name7019 (
		\P3_EAX_reg[27]/NET0131 ,
		_w2105_,
		_w2116_,
		_w8369_
	);
	LUT4 #(
		.INIT('h0008)
	) name7020 (
		_w2060_,
		_w2044_,
		_w8369_,
		_w8368_,
		_w8370_
	);
	LUT4 #(
		.INIT('h153f)
	) name7021 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8371_
	);
	LUT4 #(
		.INIT('h135f)
	) name7022 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8372_
	);
	LUT4 #(
		.INIT('h135f)
	) name7023 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8373_
	);
	LUT4 #(
		.INIT('h153f)
	) name7024 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8374_
	);
	LUT4 #(
		.INIT('h8000)
	) name7025 (
		_w8373_,
		_w8374_,
		_w8371_,
		_w8372_,
		_w8375_
	);
	LUT4 #(
		.INIT('h135f)
	) name7026 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8376_
	);
	LUT4 #(
		.INIT('h135f)
	) name7027 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8377_
	);
	LUT4 #(
		.INIT('h153f)
	) name7028 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8378_
	);
	LUT4 #(
		.INIT('h153f)
	) name7029 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8379_
	);
	LUT4 #(
		.INIT('h8000)
	) name7030 (
		_w8378_,
		_w8379_,
		_w8376_,
		_w8377_,
		_w8380_
	);
	LUT4 #(
		.INIT('h153f)
	) name7031 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1957_,
		_w1966_,
		_w8381_
	);
	LUT4 #(
		.INIT('h135f)
	) name7032 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1954_,
		_w1946_,
		_w8382_
	);
	LUT4 #(
		.INIT('h135f)
	) name7033 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1947_,
		_w1949_,
		_w8383_
	);
	LUT4 #(
		.INIT('h153f)
	) name7034 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w1956_,
		_w1950_,
		_w8384_
	);
	LUT4 #(
		.INIT('h8000)
	) name7035 (
		_w8383_,
		_w8384_,
		_w8381_,
		_w8382_,
		_w8385_
	);
	LUT4 #(
		.INIT('h135f)
	) name7036 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1952_,
		_w1967_,
		_w8386_
	);
	LUT4 #(
		.INIT('h153f)
	) name7037 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w1969_,
		_w1970_,
		_w8387_
	);
	LUT4 #(
		.INIT('h135f)
	) name7038 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1963_,
		_w1964_,
		_w8388_
	);
	LUT4 #(
		.INIT('h135f)
	) name7039 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w1960_,
		_w1961_,
		_w8389_
	);
	LUT4 #(
		.INIT('h8000)
	) name7040 (
		_w8388_,
		_w8389_,
		_w8386_,
		_w8387_,
		_w8390_
	);
	LUT4 #(
		.INIT('h0777)
	) name7041 (
		_w8375_,
		_w8380_,
		_w8385_,
		_w8390_,
		_w8391_
	);
	LUT4 #(
		.INIT('h153f)
	) name7042 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[14][1]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8392_
	);
	LUT4 #(
		.INIT('h135f)
	) name7043 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8393_
	);
	LUT4 #(
		.INIT('h135f)
	) name7044 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8394_
	);
	LUT4 #(
		.INIT('h153f)
	) name7045 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8395_
	);
	LUT4 #(
		.INIT('h8000)
	) name7046 (
		_w8394_,
		_w8395_,
		_w8392_,
		_w8393_,
		_w8396_
	);
	LUT4 #(
		.INIT('h135f)
	) name7047 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8397_
	);
	LUT4 #(
		.INIT('h135f)
	) name7048 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8398_
	);
	LUT4 #(
		.INIT('h153f)
	) name7049 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8399_
	);
	LUT4 #(
		.INIT('h153f)
	) name7050 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8400_
	);
	LUT4 #(
		.INIT('h8000)
	) name7051 (
		_w8399_,
		_w8400_,
		_w8397_,
		_w8398_,
		_w8401_
	);
	LUT2 #(
		.INIT('h8)
	) name7052 (
		_w8396_,
		_w8401_,
		_w8402_
	);
	LUT4 #(
		.INIT('h153f)
	) name7053 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8403_
	);
	LUT4 #(
		.INIT('h135f)
	) name7054 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8404_
	);
	LUT4 #(
		.INIT('h135f)
	) name7055 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8405_
	);
	LUT4 #(
		.INIT('h153f)
	) name7056 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8406_
	);
	LUT4 #(
		.INIT('h8000)
	) name7057 (
		_w8405_,
		_w8406_,
		_w8403_,
		_w8404_,
		_w8407_
	);
	LUT4 #(
		.INIT('h135f)
	) name7058 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8408_
	);
	LUT4 #(
		.INIT('h135f)
	) name7059 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8409_
	);
	LUT4 #(
		.INIT('h153f)
	) name7060 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8410_
	);
	LUT4 #(
		.INIT('h153f)
	) name7061 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8411_
	);
	LUT4 #(
		.INIT('h8000)
	) name7062 (
		_w8410_,
		_w8411_,
		_w8408_,
		_w8409_,
		_w8412_
	);
	LUT2 #(
		.INIT('h8)
	) name7063 (
		_w8407_,
		_w8412_,
		_w8413_
	);
	LUT3 #(
		.INIT('h02)
	) name7064 (
		_w8391_,
		_w8402_,
		_w8413_,
		_w8414_
	);
	LUT4 #(
		.INIT('h153f)
	) name7065 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8415_
	);
	LUT4 #(
		.INIT('h135f)
	) name7066 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8416_
	);
	LUT4 #(
		.INIT('h135f)
	) name7067 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8417_
	);
	LUT4 #(
		.INIT('h153f)
	) name7068 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8418_
	);
	LUT4 #(
		.INIT('h8000)
	) name7069 (
		_w8417_,
		_w8418_,
		_w8415_,
		_w8416_,
		_w8419_
	);
	LUT4 #(
		.INIT('h135f)
	) name7070 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8420_
	);
	LUT4 #(
		.INIT('h135f)
	) name7071 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[12][3]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8421_
	);
	LUT4 #(
		.INIT('h153f)
	) name7072 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8422_
	);
	LUT4 #(
		.INIT('h153f)
	) name7073 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8423_
	);
	LUT4 #(
		.INIT('h8000)
	) name7074 (
		_w8422_,
		_w8423_,
		_w8420_,
		_w8421_,
		_w8424_
	);
	LUT2 #(
		.INIT('h8)
	) name7075 (
		_w8419_,
		_w8424_,
		_w8425_
	);
	LUT4 #(
		.INIT('h0002)
	) name7076 (
		_w8391_,
		_w8402_,
		_w8413_,
		_w8425_,
		_w8426_
	);
	LUT4 #(
		.INIT('h153f)
	) name7077 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8427_
	);
	LUT4 #(
		.INIT('h135f)
	) name7078 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8428_
	);
	LUT4 #(
		.INIT('h135f)
	) name7079 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8429_
	);
	LUT4 #(
		.INIT('h153f)
	) name7080 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8430_
	);
	LUT4 #(
		.INIT('h8000)
	) name7081 (
		_w8429_,
		_w8430_,
		_w8427_,
		_w8428_,
		_w8431_
	);
	LUT4 #(
		.INIT('h135f)
	) name7082 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8432_
	);
	LUT4 #(
		.INIT('h135f)
	) name7083 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8433_
	);
	LUT4 #(
		.INIT('h153f)
	) name7084 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8434_
	);
	LUT4 #(
		.INIT('h153f)
	) name7085 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8435_
	);
	LUT4 #(
		.INIT('h8000)
	) name7086 (
		_w8434_,
		_w8435_,
		_w8432_,
		_w8433_,
		_w8436_
	);
	LUT2 #(
		.INIT('h8)
	) name7087 (
		_w8431_,
		_w8436_,
		_w8437_
	);
	LUT2 #(
		.INIT('h9)
	) name7088 (
		_w8426_,
		_w8437_,
		_w8438_
	);
	LUT3 #(
		.INIT('h02)
	) name7089 (
		\buf2_reg[11]/NET0131 ,
		_w2105_,
		_w2116_,
		_w8439_
	);
	LUT3 #(
		.INIT('h40)
	) name7090 (
		_w2060_,
		_w2047_,
		_w8439_,
		_w8440_
	);
	LUT4 #(
		.INIT('h0007)
	) name7091 (
		_w8366_,
		_w8438_,
		_w8370_,
		_w8440_,
		_w8441_
	);
	LUT4 #(
		.INIT('h5700)
	) name7092 (
		\P3_EAX_reg[27]/NET0131 ,
		_w2120_,
		_w8367_,
		_w8441_,
		_w8442_
	);
	LUT4 #(
		.INIT('hecee)
	) name7093 (
		_w1945_,
		_w8342_,
		_w8365_,
		_w8442_,
		_w8443_
	);
	LUT2 #(
		.INIT('h2)
	) name7094 (
		\P2_EAX_reg[27]/NET0131 ,
		_w7767_,
		_w8444_
	);
	LUT4 #(
		.INIT('h8f00)
	) name7095 (
		\P2_EAX_reg[26]/NET0131 ,
		_w7784_,
		_w7789_,
		_w7792_,
		_w8445_
	);
	LUT2 #(
		.INIT('h4)
	) name7096 (
		\P2_EAX_reg[27]/NET0131 ,
		_w7789_,
		_w8446_
	);
	LUT3 #(
		.INIT('h80)
	) name7097 (
		\P2_EAX_reg[26]/NET0131 ,
		_w7784_,
		_w8446_,
		_w8447_
	);
	LUT3 #(
		.INIT('h82)
	) name7098 (
		_w1596_,
		_w7850_,
		_w7861_,
		_w8448_
	);
	LUT2 #(
		.INIT('h8)
	) name7099 (
		_w1554_,
		_w8448_,
		_w8449_
	);
	LUT4 #(
		.INIT('hc444)
	) name7100 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[11]/NET0131 ,
		_w2255_,
		_w2260_,
		_w8450_
	);
	LUT4 #(
		.INIT('h0888)
	) name7101 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[11]/NET0131 ,
		_w2255_,
		_w2260_,
		_w8451_
	);
	LUT2 #(
		.INIT('h1)
	) name7102 (
		_w8450_,
		_w8451_,
		_w8452_
	);
	LUT2 #(
		.INIT('h2)
	) name7103 (
		_w1565_,
		_w8452_,
		_w8453_
	);
	LUT3 #(
		.INIT('h08)
	) name7104 (
		_w1501_,
		_w1568_,
		_w3552_,
		_w8454_
	);
	LUT3 #(
		.INIT('ha8)
	) name7105 (
		_w1606_,
		_w8453_,
		_w8454_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name7106 (
		_w8449_,
		_w8455_,
		_w8456_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7107 (
		\P2_EAX_reg[27]/NET0131 ,
		_w8445_,
		_w8447_,
		_w8456_,
		_w8457_
	);
	LUT3 #(
		.INIT('hce)
	) name7108 (
		_w1678_,
		_w8444_,
		_w8457_,
		_w8458_
	);
	LUT4 #(
		.INIT('hfffc)
	) name7109 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w8459_
	);
	LUT4 #(
		.INIT('hfda0)
	) name7110 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w8460_
	);
	LUT2 #(
		.INIT('h2)
	) name7111 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8460_,
		_w8461_
	);
	LUT3 #(
		.INIT('h72)
	) name7112 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8462_
	);
	LUT4 #(
		.INIT('h23af)
	) name7113 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2230_,
		_w2248_,
		_w8462_,
		_w8463_
	);
	LUT2 #(
		.INIT('h4)
	) name7114 (
		_w8461_,
		_w8463_,
		_w8464_
	);
	LUT4 #(
		.INIT('h10ff)
	) name7115 (
		_w1871_,
		_w1873_,
		_w1933_,
		_w8464_,
		_w8465_
	);
	LUT3 #(
		.INIT('h02)
	) name7116 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w3534_,
		_w3536_,
		_w8466_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7117 (
		_w3537_,
		_w3476_,
		_w3477_,
		_w8466_,
		_w8467_
	);
	LUT3 #(
		.INIT('h32)
	) name7118 (
		_w4953_,
		_w4956_,
		_w8467_,
		_w8468_
	);
	LUT4 #(
		.INIT('h08a2)
	) name7119 (
		_w3411_,
		_w3513_,
		_w3516_,
		_w3519_,
		_w8469_
	);
	LUT3 #(
		.INIT('hc4)
	) name7120 (
		_w3407_,
		_w3414_,
		_w8467_,
		_w8470_
	);
	LUT4 #(
		.INIT('hbe00)
	) name7121 (
		_w3411_,
		_w3493_,
		_w3531_,
		_w8470_,
		_w8471_
	);
	LUT2 #(
		.INIT('h2)
	) name7122 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w3545_,
		_w8472_
	);
	LUT4 #(
		.INIT('hc055)
	) name7123 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3534_,
		_w8473_
	);
	LUT3 #(
		.INIT('h31)
	) name7124 (
		_w2248_,
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7125 (
		_w8468_,
		_w8469_,
		_w8471_,
		_w8474_,
		_w8475_
	);
	LUT4 #(
		.INIT('hfda0)
	) name7126 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w8476_
	);
	LUT2 #(
		.INIT('h2)
	) name7127 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8476_,
		_w8477_
	);
	LUT3 #(
		.INIT('h72)
	) name7128 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8478_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name7129 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2215_,
		_w2216_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h4)
	) name7130 (
		_w8477_,
		_w8479_,
		_w8480_
	);
	LUT4 #(
		.INIT('h02ff)
	) name7131 (
		_w1945_,
		_w2131_,
		_w2133_,
		_w8480_,
		_w8481_
	);
	LUT4 #(
		.INIT('hfda0)
	) name7132 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w8482_
	);
	LUT2 #(
		.INIT('h2)
	) name7133 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8482_,
		_w8483_
	);
	LUT3 #(
		.INIT('h72)
	) name7134 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w8484_
	);
	LUT4 #(
		.INIT('h23af)
	) name7135 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2205_,
		_w2246_,
		_w8484_,
		_w8485_
	);
	LUT2 #(
		.INIT('h4)
	) name7136 (
		_w8483_,
		_w8485_,
		_w8486_
	);
	LUT4 #(
		.INIT('h10ff)
	) name7137 (
		_w1641_,
		_w1644_,
		_w1678_,
		_w8486_,
		_w8487_
	);
	LUT3 #(
		.INIT('h02)
	) name7138 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w3578_,
		_w3580_,
		_w8488_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7139 (
		_w3476_,
		_w3477_,
		_w3581_,
		_w8488_,
		_w8489_
	);
	LUT3 #(
		.INIT('h32)
	) name7140 (
		_w4953_,
		_w4990_,
		_w8489_,
		_w8490_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7141 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3572_,
		_w8491_
	);
	LUT3 #(
		.INIT('hc4)
	) name7142 (
		_w3407_,
		_w3575_,
		_w8489_,
		_w8492_
	);
	LUT4 #(
		.INIT('hf600)
	) name7143 (
		_w3493_,
		_w3531_,
		_w3572_,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h2)
	) name7144 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w3545_,
		_w8494_
	);
	LUT4 #(
		.INIT('hc055)
	) name7145 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3578_,
		_w8495_
	);
	LUT3 #(
		.INIT('h31)
	) name7146 (
		_w2248_,
		_w8494_,
		_w8495_,
		_w8496_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7147 (
		_w8490_,
		_w8491_,
		_w8493_,
		_w8496_,
		_w8497_
	);
	LUT3 #(
		.INIT('h02)
	) name7148 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w3536_,
		_w3412_,
		_w8498_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7149 (
		_w3476_,
		_w3477_,
		_w3597_,
		_w8498_,
		_w8499_
	);
	LUT3 #(
		.INIT('h32)
	) name7150 (
		_w4953_,
		_w5001_,
		_w8499_,
		_w8500_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7151 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3592_,
		_w8501_
	);
	LUT3 #(
		.INIT('hc4)
	) name7152 (
		_w3407_,
		_w3594_,
		_w8499_,
		_w8502_
	);
	LUT4 #(
		.INIT('hf600)
	) name7153 (
		_w3493_,
		_w3531_,
		_w3592_,
		_w8502_,
		_w8503_
	);
	LUT2 #(
		.INIT('h2)
	) name7154 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w3545_,
		_w8504_
	);
	LUT4 #(
		.INIT('hc055)
	) name7155 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3536_,
		_w8505_
	);
	LUT3 #(
		.INIT('h31)
	) name7156 (
		_w2248_,
		_w8504_,
		_w8505_,
		_w8506_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7157 (
		_w8500_,
		_w8501_,
		_w8503_,
		_w8506_,
		_w8507_
	);
	LUT3 #(
		.INIT('h02)
	) name7158 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w3534_,
		_w3611_,
		_w8508_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7159 (
		_w3476_,
		_w3477_,
		_w3612_,
		_w8508_,
		_w8509_
	);
	LUT3 #(
		.INIT('h32)
	) name7160 (
		_w4953_,
		_w5012_,
		_w8509_,
		_w8510_
	);
	LUT4 #(
		.INIT('h08a2)
	) name7161 (
		_w3412_,
		_w3513_,
		_w3516_,
		_w3519_,
		_w8511_
	);
	LUT3 #(
		.INIT('hc4)
	) name7162 (
		_w3407_,
		_w3608_,
		_w8509_,
		_w8512_
	);
	LUT4 #(
		.INIT('hbe00)
	) name7163 (
		_w3412_,
		_w3493_,
		_w3531_,
		_w8512_,
		_w8513_
	);
	LUT2 #(
		.INIT('h2)
	) name7164 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w3545_,
		_w8514_
	);
	LUT4 #(
		.INIT('hc055)
	) name7165 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3611_,
		_w8515_
	);
	LUT3 #(
		.INIT('h31)
	) name7166 (
		_w2248_,
		_w8514_,
		_w8515_,
		_w8516_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7167 (
		_w8510_,
		_w8511_,
		_w8513_,
		_w8516_,
		_w8517_
	);
	LUT3 #(
		.INIT('h02)
	) name7168 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w3572_,
		_w3611_,
		_w8518_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7169 (
		_w3476_,
		_w3477_,
		_w3626_,
		_w8518_,
		_w8519_
	);
	LUT3 #(
		.INIT('h32)
	) name7170 (
		_w4953_,
		_w5023_,
		_w8519_,
		_w8520_
	);
	LUT4 #(
		.INIT('h08a2)
	) name7171 (
		_w3536_,
		_w3513_,
		_w3516_,
		_w3519_,
		_w8521_
	);
	LUT3 #(
		.INIT('hc4)
	) name7172 (
		_w3407_,
		_w3623_,
		_w8519_,
		_w8522_
	);
	LUT4 #(
		.INIT('hbe00)
	) name7173 (
		_w3536_,
		_w3493_,
		_w3531_,
		_w8522_,
		_w8523_
	);
	LUT2 #(
		.INIT('h2)
	) name7174 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w3545_,
		_w8524_
	);
	LUT4 #(
		.INIT('hc055)
	) name7175 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3572_,
		_w8525_
	);
	LUT3 #(
		.INIT('h31)
	) name7176 (
		_w2248_,
		_w8524_,
		_w8525_,
		_w8526_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7177 (
		_w8520_,
		_w8521_,
		_w8523_,
		_w8526_,
		_w8527_
	);
	LUT3 #(
		.INIT('h02)
	) name7178 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w3572_,
		_w3573_,
		_w8528_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7179 (
		_w3476_,
		_w3477_,
		_w3574_,
		_w8528_,
		_w8529_
	);
	LUT3 #(
		.INIT('h32)
	) name7180 (
		_w4953_,
		_w5034_,
		_w8529_,
		_w8530_
	);
	LUT4 #(
		.INIT('h08a2)
	) name7181 (
		_w3534_,
		_w3513_,
		_w3516_,
		_w3519_,
		_w8531_
	);
	LUT3 #(
		.INIT('hc4)
	) name7182 (
		_w3407_,
		_w3637_,
		_w8529_,
		_w8532_
	);
	LUT4 #(
		.INIT('hbe00)
	) name7183 (
		_w3534_,
		_w3493_,
		_w3531_,
		_w8532_,
		_w8533_
	);
	LUT2 #(
		.INIT('h2)
	) name7184 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w3545_,
		_w8534_
	);
	LUT4 #(
		.INIT('hc055)
	) name7185 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3573_,
		_w8535_
	);
	LUT3 #(
		.INIT('h31)
	) name7186 (
		_w2248_,
		_w8534_,
		_w8535_,
		_w8536_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7187 (
		_w8530_,
		_w8531_,
		_w8533_,
		_w8536_,
		_w8537_
	);
	LUT3 #(
		.INIT('h02)
	) name7188 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w3580_,
		_w3573_,
		_w8538_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7189 (
		_w3476_,
		_w3477_,
		_w3653_,
		_w8538_,
		_w8539_
	);
	LUT3 #(
		.INIT('h32)
	) name7190 (
		_w4953_,
		_w5045_,
		_w8539_,
		_w8540_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7191 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3611_,
		_w8541_
	);
	LUT3 #(
		.INIT('hc4)
	) name7192 (
		_w3407_,
		_w3650_,
		_w8539_,
		_w8542_
	);
	LUT4 #(
		.INIT('hf600)
	) name7193 (
		_w3493_,
		_w3531_,
		_w3611_,
		_w8542_,
		_w8543_
	);
	LUT2 #(
		.INIT('h2)
	) name7194 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w3545_,
		_w8544_
	);
	LUT4 #(
		.INIT('hc055)
	) name7195 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3580_,
		_w8545_
	);
	LUT3 #(
		.INIT('h31)
	) name7196 (
		_w2248_,
		_w8544_,
		_w8545_,
		_w8546_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7197 (
		_w8540_,
		_w8541_,
		_w8543_,
		_w8546_,
		_w8547_
	);
	LUT3 #(
		.INIT('h02)
	) name7198 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w3578_,
		_w3667_,
		_w8548_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7199 (
		_w3476_,
		_w3477_,
		_w3668_,
		_w8548_,
		_w8549_
	);
	LUT3 #(
		.INIT('h32)
	) name7200 (
		_w4953_,
		_w5056_,
		_w8549_,
		_w8550_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7201 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3573_,
		_w8551_
	);
	LUT3 #(
		.INIT('hc4)
	) name7202 (
		_w3407_,
		_w3664_,
		_w8549_,
		_w8552_
	);
	LUT4 #(
		.INIT('hf600)
	) name7203 (
		_w3493_,
		_w3531_,
		_w3573_,
		_w8552_,
		_w8553_
	);
	LUT2 #(
		.INIT('h2)
	) name7204 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w3545_,
		_w8554_
	);
	LUT4 #(
		.INIT('hc055)
	) name7205 (
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3667_,
		_w8555_
	);
	LUT3 #(
		.INIT('h31)
	) name7206 (
		_w2248_,
		_w8554_,
		_w8555_,
		_w8556_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7207 (
		_w8550_,
		_w8551_,
		_w8553_,
		_w8556_,
		_w8557_
	);
	LUT3 #(
		.INIT('h02)
	) name7208 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w3667_,
		_w3683_,
		_w8558_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7209 (
		_w3476_,
		_w3477_,
		_w3698_,
		_w8558_,
		_w8559_
	);
	LUT3 #(
		.INIT('h32)
	) name7210 (
		_w4953_,
		_w5067_,
		_w8559_,
		_w8560_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7211 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3580_,
		_w8561_
	);
	LUT3 #(
		.INIT('hc4)
	) name7212 (
		_w3407_,
		_w3695_,
		_w8559_,
		_w8562_
	);
	LUT4 #(
		.INIT('hf600)
	) name7213 (
		_w3493_,
		_w3531_,
		_w3580_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h2)
	) name7214 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w3545_,
		_w8564_
	);
	LUT4 #(
		.INIT('hc055)
	) name7215 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3683_,
		_w8565_
	);
	LUT3 #(
		.INIT('h31)
	) name7216 (
		_w2248_,
		_w8564_,
		_w8565_,
		_w8566_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7217 (
		_w8560_,
		_w8561_,
		_w8563_,
		_w8566_,
		_w8567_
	);
	LUT3 #(
		.INIT('h02)
	) name7218 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w3682_,
		_w3683_,
		_w8568_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7219 (
		_w3476_,
		_w3477_,
		_w3684_,
		_w8568_,
		_w8569_
	);
	LUT3 #(
		.INIT('h32)
	) name7220 (
		_w4953_,
		_w5078_,
		_w8569_,
		_w8570_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7221 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3578_,
		_w8571_
	);
	LUT3 #(
		.INIT('hc4)
	) name7222 (
		_w3407_,
		_w3679_,
		_w8569_,
		_w8572_
	);
	LUT4 #(
		.INIT('hf600)
	) name7223 (
		_w3493_,
		_w3531_,
		_w3578_,
		_w8572_,
		_w8573_
	);
	LUT2 #(
		.INIT('h2)
	) name7224 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w3545_,
		_w8574_
	);
	LUT4 #(
		.INIT('hc055)
	) name7225 (
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3682_,
		_w8575_
	);
	LUT3 #(
		.INIT('h31)
	) name7226 (
		_w2248_,
		_w8574_,
		_w8575_,
		_w8576_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7227 (
		_w8570_,
		_w8571_,
		_w8573_,
		_w8576_,
		_w8577_
	);
	LUT3 #(
		.INIT('h02)
	) name7228 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w3682_,
		_w3712_,
		_w8578_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7229 (
		_w3476_,
		_w3477_,
		_w3713_,
		_w8578_,
		_w8579_
	);
	LUT3 #(
		.INIT('h32)
	) name7230 (
		_w4953_,
		_w5089_,
		_w8579_,
		_w8580_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7231 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3667_,
		_w8581_
	);
	LUT3 #(
		.INIT('hc4)
	) name7232 (
		_w3407_,
		_w3709_,
		_w8579_,
		_w8582_
	);
	LUT4 #(
		.INIT('hf600)
	) name7233 (
		_w3493_,
		_w3531_,
		_w3667_,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h2)
	) name7234 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w3545_,
		_w8584_
	);
	LUT4 #(
		.INIT('hc055)
	) name7235 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3712_,
		_w8585_
	);
	LUT3 #(
		.INIT('h31)
	) name7236 (
		_w2248_,
		_w8584_,
		_w8585_,
		_w8586_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7237 (
		_w8580_,
		_w8581_,
		_w8583_,
		_w8586_,
		_w8587_
	);
	LUT3 #(
		.INIT('h02)
	) name7238 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w3712_,
		_w3727_,
		_w8588_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7239 (
		_w3476_,
		_w3477_,
		_w3728_,
		_w8588_,
		_w8589_
	);
	LUT3 #(
		.INIT('h32)
	) name7240 (
		_w4953_,
		_w5100_,
		_w8589_,
		_w8590_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7241 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3683_,
		_w8591_
	);
	LUT3 #(
		.INIT('hc4)
	) name7242 (
		_w3407_,
		_w3724_,
		_w8589_,
		_w8592_
	);
	LUT4 #(
		.INIT('hf600)
	) name7243 (
		_w3493_,
		_w3531_,
		_w3683_,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h2)
	) name7244 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w3545_,
		_w8594_
	);
	LUT4 #(
		.INIT('hc055)
	) name7245 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3727_,
		_w8595_
	);
	LUT3 #(
		.INIT('h31)
	) name7246 (
		_w2248_,
		_w8594_,
		_w8595_,
		_w8596_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7247 (
		_w8590_,
		_w8591_,
		_w8593_,
		_w8596_,
		_w8597_
	);
	LUT3 #(
		.INIT('h02)
	) name7248 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w3727_,
		_w3742_,
		_w8598_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7249 (
		_w3476_,
		_w3477_,
		_w3743_,
		_w8598_,
		_w8599_
	);
	LUT3 #(
		.INIT('h32)
	) name7250 (
		_w4953_,
		_w5111_,
		_w8599_,
		_w8600_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7251 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3682_,
		_w8601_
	);
	LUT3 #(
		.INIT('hc4)
	) name7252 (
		_w3407_,
		_w3739_,
		_w8599_,
		_w8602_
	);
	LUT4 #(
		.INIT('hf600)
	) name7253 (
		_w3493_,
		_w3531_,
		_w3682_,
		_w8602_,
		_w8603_
	);
	LUT2 #(
		.INIT('h2)
	) name7254 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w3545_,
		_w8604_
	);
	LUT4 #(
		.INIT('hc055)
	) name7255 (
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3742_,
		_w8605_
	);
	LUT3 #(
		.INIT('h31)
	) name7256 (
		_w2248_,
		_w8604_,
		_w8605_,
		_w8606_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7257 (
		_w8600_,
		_w8601_,
		_w8603_,
		_w8606_,
		_w8607_
	);
	LUT3 #(
		.INIT('h02)
	) name7258 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w3592_,
		_w3742_,
		_w8608_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7259 (
		_w3476_,
		_w3477_,
		_w3757_,
		_w8608_,
		_w8609_
	);
	LUT3 #(
		.INIT('h32)
	) name7260 (
		_w4953_,
		_w5122_,
		_w8609_,
		_w8610_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7261 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3712_,
		_w8611_
	);
	LUT3 #(
		.INIT('hc4)
	) name7262 (
		_w3407_,
		_w3754_,
		_w8609_,
		_w8612_
	);
	LUT4 #(
		.INIT('hf600)
	) name7263 (
		_w3493_,
		_w3531_,
		_w3712_,
		_w8612_,
		_w8613_
	);
	LUT2 #(
		.INIT('h2)
	) name7264 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w3545_,
		_w8614_
	);
	LUT4 #(
		.INIT('hc055)
	) name7265 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3592_,
		_w8615_
	);
	LUT3 #(
		.INIT('h31)
	) name7266 (
		_w2248_,
		_w8614_,
		_w8615_,
		_w8616_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7267 (
		_w8610_,
		_w8611_,
		_w8613_,
		_w8616_,
		_w8617_
	);
	LUT3 #(
		.INIT('h02)
	) name7268 (
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w3411_,
		_w3592_,
		_w8618_
	);
	LUT4 #(
		.INIT('h00f1)
	) name7269 (
		_w3476_,
		_w3477_,
		_w3593_,
		_w8618_,
		_w8619_
	);
	LUT3 #(
		.INIT('h32)
	) name7270 (
		_w4953_,
		_w5133_,
		_w8619_,
		_w8620_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7271 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3727_,
		_w8621_
	);
	LUT3 #(
		.INIT('hc4)
	) name7272 (
		_w3407_,
		_w3768_,
		_w8619_,
		_w8622_
	);
	LUT4 #(
		.INIT('hf600)
	) name7273 (
		_w3493_,
		_w3531_,
		_w3727_,
		_w8622_,
		_w8623_
	);
	LUT2 #(
		.INIT('h2)
	) name7274 (
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w3545_,
		_w8624_
	);
	LUT4 #(
		.INIT('hc055)
	) name7275 (
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3411_,
		_w8625_
	);
	LUT3 #(
		.INIT('h31)
	) name7276 (
		_w2248_,
		_w8624_,
		_w8625_,
		_w8626_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7277 (
		_w8620_,
		_w8621_,
		_w8623_,
		_w8626_,
		_w8627_
	);
	LUT3 #(
		.INIT('h02)
	) name7278 (
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w3411_,
		_w3412_,
		_w8628_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7279 (
		_w3413_,
		_w3476_,
		_w3477_,
		_w8628_,
		_w8629_
	);
	LUT3 #(
		.INIT('h32)
	) name7280 (
		_w4953_,
		_w5144_,
		_w8629_,
		_w8630_
	);
	LUT4 #(
		.INIT('h2d00)
	) name7281 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3742_,
		_w8631_
	);
	LUT3 #(
		.INIT('hc4)
	) name7282 (
		_w3407_,
		_w3781_,
		_w8629_,
		_w8632_
	);
	LUT4 #(
		.INIT('hf600)
	) name7283 (
		_w3493_,
		_w3531_,
		_w3742_,
		_w8632_,
		_w8633_
	);
	LUT2 #(
		.INIT('h2)
	) name7284 (
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w3545_,
		_w8634_
	);
	LUT4 #(
		.INIT('hc055)
	) name7285 (
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1719_,
		_w1724_,
		_w3412_,
		_w8635_
	);
	LUT3 #(
		.INIT('h31)
	) name7286 (
		_w2248_,
		_w8634_,
		_w8635_,
		_w8636_
	);
	LUT4 #(
		.INIT('h45ff)
	) name7287 (
		_w8630_,
		_w8631_,
		_w8633_,
		_w8636_,
		_w8637_
	);
	LUT4 #(
		.INIT('h4447)
	) name7288 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w1661_,
		_w6431_,
		_w6432_,
		_w8638_
	);
	LUT4 #(
		.INIT('h028a)
	) name7289 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8639_
	);
	LUT4 #(
		.INIT('h007d)
	) name7290 (
		_w1659_,
		_w4399_,
		_w6435_,
		_w8639_,
		_w8640_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7291 (
		_w1559_,
		_w1678_,
		_w8638_,
		_w8640_,
		_w8641_
	);
	LUT4 #(
		.INIT('h0080)
	) name7292 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5723_,
		_w6857_,
		_w8642_
	);
	LUT4 #(
		.INIT('h3313)
	) name7293 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5723_,
		_w6857_,
		_w8643_
	);
	LUT3 #(
		.INIT('h02)
	) name7294 (
		_w1679_,
		_w8643_,
		_w8642_,
		_w8644_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7295 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w5723_,
		_w8645_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7296 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8646_
	);
	LUT3 #(
		.INIT('h70)
	) name7297 (
		_w2283_,
		_w8645_,
		_w8646_,
		_w8647_
	);
	LUT2 #(
		.INIT('h4)
	) name7298 (
		_w8644_,
		_w8647_,
		_w8648_
	);
	LUT2 #(
		.INIT('hb)
	) name7299 (
		_w8641_,
		_w8648_,
		_w8649_
	);
	LUT4 #(
		.INIT('h7774)
	) name7300 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w1661_,
		_w6459_,
		_w6457_,
		_w8650_
	);
	LUT4 #(
		.INIT('h028a)
	) name7301 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8651_
	);
	LUT3 #(
		.INIT('h0b)
	) name7302 (
		_w6462_,
		_w6463_,
		_w8651_,
		_w8652_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7303 (
		_w1559_,
		_w1678_,
		_w8650_,
		_w8652_,
		_w8653_
	);
	LUT3 #(
		.INIT('h13)
	) name7304 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w7937_,
		_w8654_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w7630_,
		_w8654_,
		_w8655_
	);
	LUT4 #(
		.INIT('h70d0)
	) name7306 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w1679_,
		_w5725_,
		_w8656_
	);
	LUT4 #(
		.INIT('hab00)
	) name7307 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7630_,
		_w8654_,
		_w8656_,
		_w8657_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7308 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8658_
	);
	LUT4 #(
		.INIT('hfd00)
	) name7309 (
		_w2283_,
		_w7630_,
		_w8654_,
		_w8658_,
		_w8659_
	);
	LUT2 #(
		.INIT('h4)
	) name7310 (
		_w8657_,
		_w8659_,
		_w8660_
	);
	LUT2 #(
		.INIT('hb)
	) name7311 (
		_w8653_,
		_w8660_,
		_w8661_
	);
	LUT4 #(
		.INIT('h0f07)
	) name7312 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2944_,
		_w4052_,
		_w4051_,
		_w8662_
	);
	LUT3 #(
		.INIT('ha8)
	) name7313 (
		_w2755_,
		_w7424_,
		_w8662_,
		_w8663_
	);
	LUT3 #(
		.INIT('h2a)
	) name7314 (
		_w2869_,
		_w4066_,
		_w4074_,
		_w8664_
	);
	LUT2 #(
		.INIT('h1)
	) name7315 (
		_w2755_,
		_w2874_,
		_w8665_
	);
	LUT3 #(
		.INIT('h45)
	) name7316 (
		_w2173_,
		_w8664_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h2)
	) name7317 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		_w7422_,
		_w8667_
	);
	LUT4 #(
		.INIT('h3313)
	) name7318 (
		\P3_InstAddrPointer_reg[9]/NET0131 ,
		_w2987_,
		_w2988_,
		_w4088_,
		_w8668_
	);
	LUT3 #(
		.INIT('h02)
	) name7319 (
		_w2181_,
		_w5789_,
		_w8668_,
		_w8669_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7320 (
		_w2181_,
		_w2987_,
		_w5788_,
		_w8667_,
		_w8670_
	);
	LUT4 #(
		.INIT('hdf00)
	) name7321 (
		_w2171_,
		_w8663_,
		_w8666_,
		_w8670_,
		_w8671_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name7322 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w8672_
	);
	LUT3 #(
		.INIT('h6a)
	) name7323 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w8673_
	);
	LUT4 #(
		.INIT('hc840)
	) name7324 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w8672_,
		_w8673_,
		_w8674_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7325 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8675_
	);
	LUT3 #(
		.INIT('h70)
	) name7326 (
		_w3055_,
		_w8672_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h4)
	) name7327 (
		_w8674_,
		_w8676_,
		_w8677_
	);
	LUT3 #(
		.INIT('h2f)
	) name7328 (
		_w1945_,
		_w8671_,
		_w8677_,
		_w8678_
	);
	LUT3 #(
		.INIT('h02)
	) name7329 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2103_,
		_w2172_,
		_w8679_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7330 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w8680_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7331 (
		_w2181_,
		_w3018_,
		_w6392_,
		_w8680_,
		_w8681_
	);
	LUT4 #(
		.INIT('h5700)
	) name7332 (
		_w2171_,
		_w6390_,
		_w8679_,
		_w8681_,
		_w8682_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7333 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5758_,
		_w8683_
	);
	LUT3 #(
		.INIT('h6c)
	) name7334 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5758_,
		_w8684_
	);
	LUT4 #(
		.INIT('hc840)
	) name7335 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w8683_,
		_w8684_,
		_w8685_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7336 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8686_
	);
	LUT3 #(
		.INIT('h70)
	) name7337 (
		_w3055_,
		_w8683_,
		_w8686_,
		_w8687_
	);
	LUT2 #(
		.INIT('h4)
	) name7338 (
		_w8685_,
		_w8687_,
		_w8688_
	);
	LUT3 #(
		.INIT('h2f)
	) name7339 (
		_w1945_,
		_w8682_,
		_w8688_,
		_w8689_
	);
	LUT3 #(
		.INIT('h02)
	) name7340 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2103_,
		_w2172_,
		_w8690_
	);
	LUT4 #(
		.INIT('haa20)
	) name7341 (
		_w2171_,
		_w6407_,
		_w6410_,
		_w8690_,
		_w8691_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name7342 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w8692_
	);
	LUT4 #(
		.INIT('h00fd)
	) name7343 (
		_w2181_,
		_w6414_,
		_w6412_,
		_w8692_,
		_w8693_
	);
	LUT3 #(
		.INIT('h6c)
	) name7344 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w8694_
	);
	LUT4 #(
		.INIT('h4105)
	) name7345 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w8695_
	);
	LUT4 #(
		.INIT('h70d0)
	) name7346 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2194_,
		_w5760_,
		_w8696_
	);
	LUT4 #(
		.INIT('h60c0)
	) name7347 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w3055_,
		_w5760_,
		_w8697_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7348 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w3054_,
		_w5783_,
		_w8698_
	);
	LUT4 #(
		.INIT('h4500)
	) name7349 (
		_w8697_,
		_w8695_,
		_w8696_,
		_w8698_,
		_w8699_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7350 (
		_w1945_,
		_w8691_,
		_w8693_,
		_w8699_,
		_w8700_
	);
	LUT3 #(
		.INIT('h08)
	) name7351 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8701_
	);
	LUT4 #(
		.INIT('h002f)
	) name7352 (
		_w3101_,
		_w5852_,
		_w5853_,
		_w8701_,
		_w8702_
	);
	LUT4 #(
		.INIT('h028a)
	) name7353 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8703_
	);
	LUT2 #(
		.INIT('h1)
	) name7354 (
		_w5855_,
		_w8703_,
		_w8704_
	);
	LUT4 #(
		.INIT('h08cc)
	) name7355 (
		_w1810_,
		_w1933_,
		_w8702_,
		_w8704_,
		_w8705_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name7356 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w7529_,
		_w8706_
	);
	LUT3 #(
		.INIT('h6a)
	) name7357 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w6367_,
		_w8707_
	);
	LUT4 #(
		.INIT('hc840)
	) name7358 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w8706_,
		_w8707_,
		_w8708_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7359 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8709_
	);
	LUT3 #(
		.INIT('h70)
	) name7360 (
		_w3407_,
		_w8706_,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h4)
	) name7361 (
		_w8708_,
		_w8710_,
		_w8711_
	);
	LUT2 #(
		.INIT('hb)
	) name7362 (
		_w8705_,
		_w8711_,
		_w8712_
	);
	LUT3 #(
		.INIT('h08)
	) name7363 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8713_
	);
	LUT4 #(
		.INIT('h9a55)
	) name7364 (
		_w3269_,
		_w3285_,
		_w3290_,
		_w3294_,
		_w8714_
	);
	LUT4 #(
		.INIT('h1141)
	) name7365 (
		_w3101_,
		_w3102_,
		_w4005_,
		_w4472_,
		_w8715_
	);
	LUT4 #(
		.INIT('h0051)
	) name7366 (
		_w1916_,
		_w3101_,
		_w8714_,
		_w8715_,
		_w8716_
	);
	LUT3 #(
		.INIT('h87)
	) name7367 (
		_w3095_,
		_w3100_,
		_w3348_,
		_w8717_
	);
	LUT4 #(
		.INIT('h4500)
	) name7368 (
		_w3351_,
		_w4020_,
		_w4021_,
		_w8717_,
		_w8718_
	);
	LUT4 #(
		.INIT('h00ba)
	) name7369 (
		_w3351_,
		_w4020_,
		_w4021_,
		_w8717_,
		_w8719_
	);
	LUT3 #(
		.INIT('h02)
	) name7370 (
		_w1924_,
		_w8719_,
		_w8718_,
		_w8720_
	);
	LUT4 #(
		.INIT('h028a)
	) name7371 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8721_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7372 (
		_w1924_,
		_w4022_,
		_w8717_,
		_w8721_,
		_w8722_
	);
	LUT4 #(
		.INIT('h5700)
	) name7373 (
		_w1810_,
		_w8713_,
		_w8716_,
		_w8722_,
		_w8723_
	);
	LUT4 #(
		.INIT('h78f0)
	) name7374 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w6365_,
		_w8724_
	);
	LUT2 #(
		.INIT('h8)
	) name7375 (
		_w6378_,
		_w8724_,
		_w8725_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7376 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8726_
	);
	LUT4 #(
		.INIT('hb700)
	) name7377 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w2310_,
		_w6366_,
		_w8726_,
		_w8727_
	);
	LUT2 #(
		.INIT('h4)
	) name7378 (
		_w8725_,
		_w8727_,
		_w8728_
	);
	LUT3 #(
		.INIT('h2f)
	) name7379 (
		_w1933_,
		_w8723_,
		_w8728_,
		_w8729_
	);
	LUT3 #(
		.INIT('h08)
	) name7380 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1842_,
		_w1915_,
		_w8730_
	);
	LUT3 #(
		.INIT('h82)
	) name7381 (
		_w3101_,
		_w3267_,
		_w3296_,
		_w8731_
	);
	LUT3 #(
		.INIT('h8a)
	) name7382 (
		_w3211_,
		_w4003_,
		_w4007_,
		_w8732_
	);
	LUT4 #(
		.INIT('h5554)
	) name7383 (
		_w1916_,
		_w3101_,
		_w3214_,
		_w8732_,
		_w8733_
	);
	LUT4 #(
		.INIT('h8a88)
	) name7384 (
		_w1810_,
		_w8730_,
		_w8731_,
		_w8733_,
		_w8734_
	);
	LUT3 #(
		.INIT('h6a)
	) name7385 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w3064_,
		_w3347_,
		_w8735_
	);
	LUT4 #(
		.INIT('h8a20)
	) name7386 (
		_w1924_,
		_w4023_,
		_w4024_,
		_w8735_,
		_w8736_
	);
	LUT4 #(
		.INIT('h028a)
	) name7387 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w8737_
	);
	LUT2 #(
		.INIT('h1)
	) name7388 (
		_w8736_,
		_w8737_,
		_w8738_
	);
	LUT3 #(
		.INIT('h6c)
	) name7389 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w7529_,
		_w8739_
	);
	LUT4 #(
		.INIT('h4105)
	) name7390 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w7529_,
		_w8740_
	);
	LUT4 #(
		.INIT('h70d0)
	) name7391 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w1939_,
		_w6367_,
		_w8741_
	);
	LUT4 #(
		.INIT('h60c0)
	) name7392 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w3407_,
		_w7529_,
		_w8742_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7393 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w3406_,
		_w6383_,
		_w8743_
	);
	LUT4 #(
		.INIT('h4500)
	) name7394 (
		_w8742_,
		_w8740_,
		_w8741_,
		_w8743_,
		_w8744_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7395 (
		_w1933_,
		_w8734_,
		_w8738_,
		_w8744_,
		_w8745_
	);
	LUT3 #(
		.INIT('h08)
	) name7396 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w1592_,
		_w1660_,
		_w8746_
	);
	LUT4 #(
		.INIT('haa20)
	) name7397 (
		_w1559_,
		_w5838_,
		_w5841_,
		_w8746_,
		_w8747_
	);
	LUT4 #(
		.INIT('h028a)
	) name7398 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w8748_
	);
	LUT2 #(
		.INIT('h1)
	) name7399 (
		_w5843_,
		_w8748_,
		_w8749_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name7400 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w8750_
	);
	LUT3 #(
		.INIT('h6a)
	) name7401 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w8751_
	);
	LUT4 #(
		.INIT('hc840)
	) name7402 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w8750_,
		_w8751_,
		_w8752_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7403 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w2286_,
		_w5747_,
		_w8753_
	);
	LUT3 #(
		.INIT('h70)
	) name7404 (
		_w2283_,
		_w8750_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h4)
	) name7405 (
		_w8752_,
		_w8754_,
		_w8755_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7406 (
		_w1678_,
		_w8747_,
		_w8749_,
		_w8755_,
		_w8756_
	);
	LUT3 #(
		.INIT('h80)
	) name7407 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2788_,
		_w2793_,
		_w8757_
	);
	LUT3 #(
		.INIT('h6a)
	) name7408 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2788_,
		_w2793_,
		_w8758_
	);
	LUT4 #(
		.INIT('h0004)
	) name7409 (
		_w2060_,
		_w2041_,
		_w2173_,
		_w8758_,
		_w8759_
	);
	LUT4 #(
		.INIT('h8000)
	) name7410 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w8758_,
		_w8760_
	);
	LUT2 #(
		.INIT('h1)
	) name7411 (
		_w8759_,
		_w8760_,
		_w8761_
	);
	LUT4 #(
		.INIT('h0010)
	) name7412 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2073_,
		_w2086_,
		_w2099_,
		_w8762_
	);
	LUT4 #(
		.INIT('h0002)
	) name7413 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2064_,
		_w8763_
	);
	LUT3 #(
		.INIT('h40)
	) name7414 (
		_w2174_,
		_w2176_,
		_w8763_,
		_w8764_
	);
	LUT4 #(
		.INIT('h222a)
	) name7415 (
		_w1945_,
		_w8761_,
		_w8762_,
		_w8764_,
		_w8765_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7416 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w3054_,
		_w3056_,
		_w8766_
	);
	LUT2 #(
		.INIT('hb)
	) name7417 (
		_w8765_,
		_w8766_,
		_w8767_
	);
	LUT3 #(
		.INIT('h8a)
	) name7418 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w4784_,
		_w4785_,
		_w8768_
	);
	LUT2 #(
		.INIT('h1)
	) name7419 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2117_,
		_w8769_
	);
	LUT3 #(
		.INIT('h0b)
	) name7420 (
		_w2073_,
		_w2086_,
		_w3002_,
		_w8770_
	);
	LUT3 #(
		.INIT('h6a)
	) name7421 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2777_,
		_w2782_,
		_w8771_
	);
	LUT3 #(
		.INIT('h78)
	) name7422 (
		_w2777_,
		_w2782_,
		_w3002_,
		_w8772_
	);
	LUT4 #(
		.INIT('h4501)
	) name7423 (
		_w2755_,
		_w8757_,
		_w8772_,
		_w8771_,
		_w8773_
	);
	LUT3 #(
		.INIT('h28)
	) name7424 (
		_w2755_,
		_w2795_,
		_w8771_,
		_w8774_
	);
	LUT3 #(
		.INIT('h54)
	) name7425 (
		_w2173_,
		_w8773_,
		_w8774_,
		_w8775_
	);
	LUT4 #(
		.INIT('h4447)
	) name7426 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2173_,
		_w8773_,
		_w8774_,
		_w8776_
	);
	LUT2 #(
		.INIT('h2)
	) name7427 (
		_w2171_,
		_w8776_,
		_w8777_
	);
	LUT3 #(
		.INIT('h6c)
	) name7428 (
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		_w2098_,
		_w8778_
	);
	LUT3 #(
		.INIT('he4)
	) name7429 (
		_w3005_,
		_w8772_,
		_w8771_,
		_w8779_
	);
	LUT4 #(
		.INIT('h8000)
	) name7430 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w8779_,
		_w8780_
	);
	LUT4 #(
		.INIT('h001f)
	) name7431 (
		_w2071_,
		_w2087_,
		_w8778_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h4)
	) name7432 (
		_w8777_,
		_w8781_,
		_w8782_
	);
	LUT4 #(
		.INIT('h0100)
	) name7433 (
		_w8768_,
		_w8770_,
		_w8769_,
		_w8782_,
		_w8783_
	);
	LUT2 #(
		.INIT('h8)
	) name7434 (
		\P3_rEIP_reg[1]/NET0131 ,
		_w3054_,
		_w8784_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7435 (
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w3054_,
		_w3056_,
		_w8785_
	);
	LUT3 #(
		.INIT('h2f)
	) name7436 (
		_w1945_,
		_w8783_,
		_w8785_,
		_w8786_
	);
	LUT4 #(
		.INIT('h0010)
	) name7437 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1571_,
		_w1583_,
		_w1640_,
		_w8787_
	);
	LUT4 #(
		.INIT('h0080)
	) name7438 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1570_,
		_w1643_,
		_w1667_,
		_w8788_
	);
	LUT3 #(
		.INIT('h6a)
	) name7439 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w4133_,
		_w4138_,
		_w8789_
	);
	LUT2 #(
		.INIT('h1)
	) name7440 (
		_w1661_,
		_w8789_,
		_w8790_
	);
	LUT3 #(
		.INIT('h56)
	) name7441 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		_w1661_,
		_w4139_,
		_w8791_
	);
	LUT2 #(
		.INIT('h2)
	) name7442 (
		_w1559_,
		_w8791_,
		_w8792_
	);
	LUT3 #(
		.INIT('h80)
	) name7443 (
		_w1558_,
		_w1596_,
		_w8789_,
		_w8793_
	);
	LUT2 #(
		.INIT('h1)
	) name7444 (
		_w8792_,
		_w8793_,
		_w8794_
	);
	LUT4 #(
		.INIT('h02aa)
	) name7445 (
		_w1678_,
		_w8787_,
		_w8788_,
		_w8794_,
		_w8795_
	);
	LUT2 #(
		.INIT('h8)
	) name7446 (
		\P2_rEIP_reg[0]/NET0131 ,
		_w2286_,
		_w8796_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7447 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w2286_,
		_w4441_,
		_w8797_
	);
	LUT2 #(
		.INIT('hb)
	) name7448 (
		_w8795_,
		_w8797_,
		_w8798_
	);
	LUT3 #(
		.INIT('h2a)
	) name7449 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1808_,
		_w1914_,
		_w8799_
	);
	LUT4 #(
		.INIT('h5545)
	) name7450 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1816_,
		_w1831_,
		_w1847_,
		_w8800_
	);
	LUT3 #(
		.INIT('h6a)
	) name7451 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w3162_,
		_w3167_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name7452 (
		_w1916_,
		_w8801_,
		_w8802_
	);
	LUT3 #(
		.INIT('h56)
	) name7453 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		_w1916_,
		_w3168_,
		_w8803_
	);
	LUT2 #(
		.INIT('h2)
	) name7454 (
		_w1810_,
		_w8803_,
		_w8804_
	);
	LUT3 #(
		.INIT('h80)
	) name7455 (
		_w1809_,
		_w1846_,
		_w8801_,
		_w8805_
	);
	LUT2 #(
		.INIT('h1)
	) name7456 (
		_w8804_,
		_w8805_,
		_w8806_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7457 (
		_w1933_,
		_w8800_,
		_w8799_,
		_w8806_,
		_w8807_
	);
	LUT2 #(
		.INIT('h8)
	) name7458 (
		\P1_rEIP_reg[0]/NET0131 ,
		_w3406_,
		_w8808_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7459 (
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w3406_,
		_w3408_,
		_w8809_
	);
	LUT2 #(
		.INIT('hb)
	) name7460 (
		_w8807_,
		_w8809_,
		_w8810_
	);
	LUT3 #(
		.INIT('hb0)
	) name7461 (
		_w1571_,
		_w1583_,
		_w4293_,
		_w8811_
	);
	LUT4 #(
		.INIT('hec00)
	) name7462 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1606_,
		_w8812_
	);
	LUT2 #(
		.INIT('h1)
	) name7463 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1563_,
		_w8813_
	);
	LUT2 #(
		.INIT('h4)
	) name7464 (
		_w8812_,
		_w8813_,
		_w8814_
	);
	LUT4 #(
		.INIT('hec00)
	) name7465 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w1605_,
		_w8815_
	);
	LUT4 #(
		.INIT('h0002)
	) name7466 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1626_,
		_w1667_,
		_w8815_,
		_w8816_
	);
	LUT3 #(
		.INIT('h87)
	) name7467 (
		_w4121_,
		_w4126_,
		_w4293_,
		_w8817_
	);
	LUT3 #(
		.INIT('h6a)
	) name7468 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w4121_,
		_w4126_,
		_w8818_
	);
	LUT4 #(
		.INIT('h4051)
	) name7469 (
		_w4214_,
		_w4295_,
		_w8818_,
		_w8817_,
		_w8819_
	);
	LUT3 #(
		.INIT('h28)
	) name7470 (
		_w4214_,
		_w4140_,
		_w8818_,
		_w8820_
	);
	LUT4 #(
		.INIT('h4447)
	) name7471 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1661_,
		_w8819_,
		_w8820_,
		_w8821_
	);
	LUT2 #(
		.INIT('h2)
	) name7472 (
		_w1559_,
		_w8821_,
		_w8822_
	);
	LUT3 #(
		.INIT('ha9)
	) name7473 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1605_,
		_w1611_,
		_w8823_
	);
	LUT3 #(
		.INIT('hd8)
	) name7474 (
		_w4390_,
		_w8818_,
		_w8817_,
		_w8824_
	);
	LUT3 #(
		.INIT('h80)
	) name7475 (
		_w1558_,
		_w1596_,
		_w8824_,
		_w8825_
	);
	LUT4 #(
		.INIT('hccc6)
	) name7476 (
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		_w1592_,
		_w1595_,
		_w8826_
	);
	LUT4 #(
		.INIT('hc800)
	) name7477 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w8826_,
		_w8827_
	);
	LUT4 #(
		.INIT('h0007)
	) name7478 (
		_w4927_,
		_w8823_,
		_w8825_,
		_w8827_,
		_w8828_
	);
	LUT4 #(
		.INIT('h5400)
	) name7479 (
		_w8822_,
		_w8814_,
		_w8816_,
		_w8828_,
		_w8829_
	);
	LUT2 #(
		.INIT('h8)
	) name7480 (
		\P2_rEIP_reg[1]/NET0131 ,
		_w2286_,
		_w8830_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7481 (
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w2286_,
		_w4441_,
		_w8831_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7482 (
		_w1678_,
		_w8811_,
		_w8829_,
		_w8831_,
		_w8832_
	);
	LUT3 #(
		.INIT('h31)
	) name7483 (
		_w1852_,
		_w1921_,
		_w3399_,
		_w8833_
	);
	LUT3 #(
		.INIT('h2a)
	) name7484 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1810_,
		_w1916_,
		_w8834_
	);
	LUT3 #(
		.INIT('h15)
	) name7485 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1805_,
		_w1806_,
		_w8835_
	);
	LUT3 #(
		.INIT('h70)
	) name7486 (
		_w1920_,
		_w4739_,
		_w8835_,
		_w8836_
	);
	LUT4 #(
		.INIT('h007f)
	) name7487 (
		_w1914_,
		_w8833_,
		_w8834_,
		_w8836_,
		_w8837_
	);
	LUT4 #(
		.INIT('hfb00)
	) name7488 (
		_w1816_,
		_w1831_,
		_w1847_,
		_w3155_,
		_w8838_
	);
	LUT3 #(
		.INIT('h87)
	) name7489 (
		_w3148_,
		_w3153_,
		_w3155_,
		_w8839_
	);
	LUT3 #(
		.INIT('h6a)
	) name7490 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w3148_,
		_w3153_,
		_w8840_
	);
	LUT4 #(
		.INIT('h4051)
	) name7491 (
		_w3101_,
		_w3169_,
		_w8840_,
		_w8839_,
		_w8841_
	);
	LUT3 #(
		.INIT('h28)
	) name7492 (
		_w3101_,
		_w3275_,
		_w8840_,
		_w8842_
	);
	LUT4 #(
		.INIT('h2220)
	) name7493 (
		_w1810_,
		_w1916_,
		_w8841_,
		_w8842_,
		_w8843_
	);
	LUT3 #(
		.INIT('hd8)
	) name7494 (
		_w3337_,
		_w8840_,
		_w8839_,
		_w8844_
	);
	LUT3 #(
		.INIT('h80)
	) name7495 (
		_w1809_,
		_w1846_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h1)
	) name7496 (
		_w8843_,
		_w8845_,
		_w8846_
	);
	LUT3 #(
		.INIT('h06)
	) name7497 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		_w1867_,
		_w4710_,
		_w8847_
	);
	LUT2 #(
		.INIT('h2)
	) name7498 (
		_w8846_,
		_w8847_,
		_w8848_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7499 (
		_w1933_,
		_w8838_,
		_w8837_,
		_w8848_,
		_w8849_
	);
	LUT2 #(
		.INIT('h8)
	) name7500 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w3406_,
		_w8850_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7501 (
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w3406_,
		_w3408_,
		_w8851_
	);
	LUT2 #(
		.INIT('hb)
	) name7502 (
		_w8849_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h2)
	) name7503 (
		\P3_EAX_reg[31]/NET0131 ,
		_w8341_,
		_w8853_
	);
	LUT3 #(
		.INIT('h80)
	) name7504 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w8363_,
		_w8854_
	);
	LUT4 #(
		.INIT('h8000)
	) name7505 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		\P3_EAX_reg[30]/NET0131 ,
		_w8363_,
		_w8855_
	);
	LUT3 #(
		.INIT('h48)
	) name7506 (
		\P3_EAX_reg[31]/NET0131 ,
		_w8361_,
		_w8855_,
		_w8856_
	);
	LUT4 #(
		.INIT('h153f)
	) name7507 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8857_
	);
	LUT4 #(
		.INIT('h135f)
	) name7508 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8858_
	);
	LUT4 #(
		.INIT('h135f)
	) name7509 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8859_
	);
	LUT4 #(
		.INIT('h153f)
	) name7510 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8860_
	);
	LUT4 #(
		.INIT('h8000)
	) name7511 (
		_w8859_,
		_w8860_,
		_w8857_,
		_w8858_,
		_w8861_
	);
	LUT4 #(
		.INIT('h135f)
	) name7512 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8862_
	);
	LUT4 #(
		.INIT('h135f)
	) name7513 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8863_
	);
	LUT4 #(
		.INIT('h153f)
	) name7514 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8864_
	);
	LUT4 #(
		.INIT('h153f)
	) name7515 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8865_
	);
	LUT4 #(
		.INIT('h8000)
	) name7516 (
		_w8864_,
		_w8865_,
		_w8862_,
		_w8863_,
		_w8866_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		_w8861_,
		_w8866_,
		_w8867_
	);
	LUT4 #(
		.INIT('h153f)
	) name7518 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8868_
	);
	LUT4 #(
		.INIT('h135f)
	) name7519 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8869_
	);
	LUT4 #(
		.INIT('h135f)
	) name7520 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8870_
	);
	LUT4 #(
		.INIT('h153f)
	) name7521 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8871_
	);
	LUT4 #(
		.INIT('h8000)
	) name7522 (
		_w8870_,
		_w8871_,
		_w8868_,
		_w8869_,
		_w8872_
	);
	LUT4 #(
		.INIT('h135f)
	) name7523 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8873_
	);
	LUT4 #(
		.INIT('h135f)
	) name7524 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8874_
	);
	LUT4 #(
		.INIT('h153f)
	) name7525 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8875_
	);
	LUT4 #(
		.INIT('h153f)
	) name7526 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8876_
	);
	LUT4 #(
		.INIT('h8000)
	) name7527 (
		_w8875_,
		_w8876_,
		_w8873_,
		_w8874_,
		_w8877_
	);
	LUT2 #(
		.INIT('h8)
	) name7528 (
		_w8872_,
		_w8877_,
		_w8878_
	);
	LUT4 #(
		.INIT('h0002)
	) name7529 (
		_w8426_,
		_w8437_,
		_w8867_,
		_w8878_,
		_w8879_
	);
	LUT4 #(
		.INIT('h153f)
	) name7530 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1956_,
		_w1947_,
		_w8880_
	);
	LUT4 #(
		.INIT('h135f)
	) name7531 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w1949_,
		_w1963_,
		_w8881_
	);
	LUT4 #(
		.INIT('h135f)
	) name7532 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1969_,
		_w1964_,
		_w8882_
	);
	LUT4 #(
		.INIT('h153f)
	) name7533 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1957_,
		_w1970_,
		_w8883_
	);
	LUT4 #(
		.INIT('h8000)
	) name7534 (
		_w8882_,
		_w8883_,
		_w8880_,
		_w8881_,
		_w8884_
	);
	LUT4 #(
		.INIT('h135f)
	) name7535 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w1966_,
		_w1967_,
		_w8885_
	);
	LUT4 #(
		.INIT('h135f)
	) name7536 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w1954_,
		_w1950_,
		_w8886_
	);
	LUT4 #(
		.INIT('h153f)
	) name7537 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1946_,
		_w1960_,
		_w8887_
	);
	LUT4 #(
		.INIT('h153f)
	) name7538 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1952_,
		_w1961_,
		_w8888_
	);
	LUT4 #(
		.INIT('h8000)
	) name7539 (
		_w8887_,
		_w8888_,
		_w8885_,
		_w8886_,
		_w8889_
	);
	LUT2 #(
		.INIT('h8)
	) name7540 (
		_w8884_,
		_w8889_,
		_w8890_
	);
	LUT3 #(
		.INIT('h08)
	) name7541 (
		_w8366_,
		_w8879_,
		_w8890_,
		_w8891_
	);
	LUT3 #(
		.INIT('h01)
	) name7542 (
		_w2120_,
		_w2121_,
		_w8367_,
		_w8892_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7543 (
		\P3_EAX_reg[31]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w8893_
	);
	LUT2 #(
		.INIT('h1)
	) name7544 (
		_w8891_,
		_w8893_,
		_w8894_
	);
	LUT4 #(
		.INIT('hecee)
	) name7545 (
		_w1945_,
		_w8853_,
		_w8856_,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h2)
	) name7546 (
		\P3_EAX_reg[30]/NET0131 ,
		_w8341_,
		_w8896_
	);
	LUT3 #(
		.INIT('h48)
	) name7547 (
		\P3_EAX_reg[30]/NET0131 ,
		_w8361_,
		_w8854_,
		_w8897_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7548 (
		\P3_EAX_reg[30]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w8898_
	);
	LUT3 #(
		.INIT('h82)
	) name7549 (
		_w8366_,
		_w8879_,
		_w8890_,
		_w8899_
	);
	LUT3 #(
		.INIT('h80)
	) name7550 (
		\buf2_reg[30]/NET0131 ,
		_w2060_,
		_w2044_,
		_w8900_
	);
	LUT3 #(
		.INIT('h20)
	) name7551 (
		\buf2_reg[14]/NET0131 ,
		_w2060_,
		_w2047_,
		_w8901_
	);
	LUT3 #(
		.INIT('ha8)
	) name7552 (
		_w2119_,
		_w8900_,
		_w8901_,
		_w8902_
	);
	LUT2 #(
		.INIT('h1)
	) name7553 (
		_w8899_,
		_w8902_,
		_w8903_
	);
	LUT2 #(
		.INIT('h4)
	) name7554 (
		_w8898_,
		_w8903_,
		_w8904_
	);
	LUT4 #(
		.INIT('hecee)
	) name7555 (
		_w1945_,
		_w8896_,
		_w8897_,
		_w8904_,
		_w8905_
	);
	LUT4 #(
		.INIT('h8000)
	) name7556 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w8906_
	);
	LUT4 #(
		.INIT('h8000)
	) name7557 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w8906_,
		_w8907_
	);
	LUT4 #(
		.INIT('h8000)
	) name7558 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w8907_,
		_w8908_
	);
	LUT2 #(
		.INIT('h8)
	) name7559 (
		\P3_EBX_reg[10]/NET0131 ,
		_w8908_,
		_w8909_
	);
	LUT3 #(
		.INIT('h80)
	) name7560 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		_w8908_,
		_w8910_
	);
	LUT4 #(
		.INIT('h8000)
	) name7561 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[12]/NET0131 ,
		_w8908_,
		_w8911_
	);
	LUT2 #(
		.INIT('h8)
	) name7562 (
		\P3_EBX_reg[13]/NET0131 ,
		_w8911_,
		_w8912_
	);
	LUT3 #(
		.INIT('h80)
	) name7563 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		_w8911_,
		_w8913_
	);
	LUT4 #(
		.INIT('h8000)
	) name7564 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[15]/NET0131 ,
		_w8911_,
		_w8914_
	);
	LUT2 #(
		.INIT('h8)
	) name7565 (
		\P3_EBX_reg[16]/NET0131 ,
		_w8914_,
		_w8915_
	);
	LUT3 #(
		.INIT('h80)
	) name7566 (
		\P3_EBX_reg[16]/NET0131 ,
		\P3_EBX_reg[17]/NET0131 ,
		_w8914_,
		_w8916_
	);
	LUT4 #(
		.INIT('h8000)
	) name7567 (
		\P3_EBX_reg[16]/NET0131 ,
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		_w8914_,
		_w8917_
	);
	LUT4 #(
		.INIT('h8000)
	) name7568 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[23]/NET0131 ,
		_w8918_
	);
	LUT3 #(
		.INIT('h80)
	) name7569 (
		\P3_EBX_reg[19]/NET0131 ,
		_w8917_,
		_w8918_,
		_w8919_
	);
	LUT4 #(
		.INIT('h8000)
	) name7570 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[24]/NET0131 ,
		_w8917_,
		_w8918_,
		_w8920_
	);
	LUT4 #(
		.INIT('h8000)
	) name7571 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		\P3_EBX_reg[29]/NET0131 ,
		_w8921_
	);
	LUT4 #(
		.INIT('h8000)
	) name7572 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[30]/NET0131 ,
		_w8920_,
		_w8921_,
		_w8922_
	);
	LUT3 #(
		.INIT('h80)
	) name7573 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w8923_
	);
	LUT3 #(
		.INIT('h08)
	) name7574 (
		_w2075_,
		_w2083_,
		_w2070_,
		_w8924_
	);
	LUT2 #(
		.INIT('h1)
	) name7575 (
		_w8923_,
		_w8924_,
		_w8925_
	);
	LUT3 #(
		.INIT('h02)
	) name7576 (
		\P3_EBX_reg[31]/NET0131 ,
		_w8923_,
		_w8924_,
		_w8926_
	);
	LUT3 #(
		.INIT('h20)
	) name7577 (
		_w8879_,
		_w8890_,
		_w8923_,
		_w8927_
	);
	LUT2 #(
		.INIT('h1)
	) name7578 (
		_w8926_,
		_w8927_,
		_w8928_
	);
	LUT4 #(
		.INIT('hb700)
	) name7579 (
		\P3_EBX_reg[31]/NET0131 ,
		_w2084_,
		_w8922_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h2)
	) name7580 (
		\P3_EBX_reg[31]/NET0131 ,
		_w8341_,
		_w8930_
	);
	LUT3 #(
		.INIT('hf2)
	) name7581 (
		_w1945_,
		_w8929_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h2)
	) name7582 (
		\P2_EAX_reg[30]/NET0131 ,
		_w7767_,
		_w8932_
	);
	LUT4 #(
		.INIT('h8008)
	) name7583 (
		_w1554_,
		_w1596_,
		_w7885_,
		_w7896_,
		_w8933_
	);
	LUT4 #(
		.INIT('h0080)
	) name7584 (
		_w1501_,
		_w1568_,
		_w1606_,
		_w4968_,
		_w8934_
	);
	LUT4 #(
		.INIT('h3111)
	) name7585 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[14]/NET0131 ,
		_w2255_,
		_w2260_,
		_w8935_
	);
	LUT4 #(
		.INIT('h0222)
	) name7586 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[14]/NET0131 ,
		_w2255_,
		_w2260_,
		_w8936_
	);
	LUT2 #(
		.INIT('h1)
	) name7587 (
		_w8935_,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h8)
	) name7588 (
		_w1606_,
		_w8937_,
		_w8938_
	);
	LUT2 #(
		.INIT('h8)
	) name7589 (
		_w1565_,
		_w8938_,
		_w8939_
	);
	LUT2 #(
		.INIT('h1)
	) name7590 (
		_w8934_,
		_w8939_,
		_w8940_
	);
	LUT4 #(
		.INIT('h0d00)
	) name7591 (
		\P2_EAX_reg[30]/NET0131 ,
		_w7792_,
		_w8933_,
		_w8940_,
		_w8941_
	);
	LUT4 #(
		.INIT('h9f00)
	) name7592 (
		\P2_EAX_reg[30]/NET0131 ,
		_w7787_,
		_w7789_,
		_w8941_,
		_w8942_
	);
	LUT3 #(
		.INIT('hce)
	) name7593 (
		_w1678_,
		_w8932_,
		_w8942_,
		_w8943_
	);
	LUT4 #(
		.INIT('h8000)
	) name7594 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w8944_
	);
	LUT4 #(
		.INIT('h8000)
	) name7595 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w8944_,
		_w8945_
	);
	LUT4 #(
		.INIT('h8000)
	) name7596 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w8945_,
		_w8946_
	);
	LUT2 #(
		.INIT('h8)
	) name7597 (
		\P2_EBX_reg[10]/NET0131 ,
		_w8946_,
		_w8947_
	);
	LUT3 #(
		.INIT('h80)
	) name7598 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		_w8946_,
		_w8948_
	);
	LUT4 #(
		.INIT('h8000)
	) name7599 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[12]/NET0131 ,
		_w8946_,
		_w8949_
	);
	LUT2 #(
		.INIT('h8)
	) name7600 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		_w8950_
	);
	LUT2 #(
		.INIT('h8)
	) name7601 (
		_w8949_,
		_w8950_,
		_w8951_
	);
	LUT3 #(
		.INIT('h80)
	) name7602 (
		\P2_EBX_reg[15]/NET0131 ,
		_w8949_,
		_w8950_,
		_w8952_
	);
	LUT4 #(
		.INIT('h8000)
	) name7603 (
		\P2_EBX_reg[15]/NET0131 ,
		\P2_EBX_reg[16]/NET0131 ,
		_w8949_,
		_w8950_,
		_w8953_
	);
	LUT2 #(
		.INIT('h8)
	) name7604 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w8954_
	);
	LUT3 #(
		.INIT('h80)
	) name7605 (
		\P2_EBX_reg[19]/NET0131 ,
		_w8953_,
		_w8954_,
		_w8955_
	);
	LUT4 #(
		.INIT('h8000)
	) name7606 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w8956_
	);
	LUT4 #(
		.INIT('h8000)
	) name7607 (
		\P2_EBX_reg[19]/NET0131 ,
		_w8953_,
		_w8954_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h8)
	) name7608 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		_w8958_
	);
	LUT3 #(
		.INIT('h80)
	) name7609 (
		\P2_EBX_reg[26]/NET0131 ,
		_w8957_,
		_w8958_,
		_w8959_
	);
	LUT4 #(
		.INIT('h8000)
	) name7610 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[27]/NET0131 ,
		_w8957_,
		_w8958_,
		_w8960_
	);
	LUT4 #(
		.INIT('hf870)
	) name7611 (
		_w1503_,
		_w1549_,
		_w1578_,
		_w1596_,
		_w8961_
	);
	LUT4 #(
		.INIT('h3f15)
	) name7612 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1550_,
		_w8448_,
		_w8961_,
		_w8962_
	);
	LUT4 #(
		.INIT('hb700)
	) name7613 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1578_,
		_w8959_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h2)
	) name7614 (
		\P2_EBX_reg[27]/NET0131 ,
		_w7767_,
		_w8964_
	);
	LUT3 #(
		.INIT('hf2)
	) name7615 (
		_w1678_,
		_w8963_,
		_w8964_,
		_w8965_
	);
	LUT3 #(
		.INIT('h80)
	) name7616 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w8960_,
		_w8966_
	);
	LUT4 #(
		.INIT('h8000)
	) name7617 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		\P2_EBX_reg[30]/NET0131 ,
		_w8960_,
		_w8967_
	);
	LUT3 #(
		.INIT('h80)
	) name7618 (
		_w1503_,
		_w1549_,
		_w7897_,
		_w8968_
	);
	LUT4 #(
		.INIT('h31f5)
	) name7619 (
		\P2_EBX_reg[31]/NET0131 ,
		_w7885_,
		_w8961_,
		_w8968_,
		_w8969_
	);
	LUT4 #(
		.INIT('hb700)
	) name7620 (
		\P2_EBX_reg[31]/NET0131 ,
		_w1578_,
		_w8967_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h2)
	) name7621 (
		\P2_EBX_reg[31]/NET0131 ,
		_w7767_,
		_w8971_
	);
	LUT3 #(
		.INIT('hf2)
	) name7622 (
		_w1678_,
		_w8970_,
		_w8971_,
		_w8972_
	);
	LUT4 #(
		.INIT('h8000)
	) name7623 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w8973_
	);
	LUT4 #(
		.INIT('h8000)
	) name7624 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w8973_,
		_w8974_
	);
	LUT4 #(
		.INIT('h8000)
	) name7625 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h8)
	) name7626 (
		\P1_EBX_reg[10]/NET0131 ,
		_w8975_,
		_w8976_
	);
	LUT3 #(
		.INIT('h80)
	) name7627 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		_w8975_,
		_w8977_
	);
	LUT4 #(
		.INIT('h8000)
	) name7628 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w8975_,
		_w8978_
	);
	LUT2 #(
		.INIT('h8)
	) name7629 (
		\P1_EBX_reg[13]/NET0131 ,
		_w8978_,
		_w8979_
	);
	LUT3 #(
		.INIT('h80)
	) name7630 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		_w8978_,
		_w8980_
	);
	LUT4 #(
		.INIT('h8000)
	) name7631 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w8978_,
		_w8981_
	);
	LUT2 #(
		.INIT('h8)
	) name7632 (
		\P1_EBX_reg[16]/NET0131 ,
		_w8981_,
		_w8982_
	);
	LUT3 #(
		.INIT('h80)
	) name7633 (
		\P1_EBX_reg[16]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		_w8981_,
		_w8983_
	);
	LUT4 #(
		.INIT('h8000)
	) name7634 (
		\P1_EBX_reg[16]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w8981_,
		_w8984_
	);
	LUT4 #(
		.INIT('h8000)
	) name7635 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		_w8985_
	);
	LUT3 #(
		.INIT('h80)
	) name7636 (
		\P1_EBX_reg[19]/NET0131 ,
		_w8984_,
		_w8985_,
		_w8986_
	);
	LUT4 #(
		.INIT('h8000)
	) name7637 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[24]/NET0131 ,
		_w8984_,
		_w8985_,
		_w8987_
	);
	LUT3 #(
		.INIT('h80)
	) name7638 (
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h8)
	) name7639 (
		\P1_EBX_reg[27]/NET0131 ,
		\P1_EBX_reg[28]/NET0131 ,
		_w8989_
	);
	LUT4 #(
		.INIT('h8000)
	) name7640 (
		\P1_EBX_reg[27]/NET0131 ,
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w8990_
	);
	LUT4 #(
		.INIT('h8000)
	) name7641 (
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w8987_,
		_w8990_,
		_w8991_
	);
	LUT4 #(
		.INIT('h0777)
	) name7642 (
		_w1750_,
		_w1813_,
		_w1826_,
		_w1828_,
		_w8992_
	);
	LUT2 #(
		.INIT('h1)
	) name7643 (
		_w1863_,
		_w8992_,
		_w8993_
	);
	LUT3 #(
		.INIT('ha8)
	) name7644 (
		\P1_EBX_reg[31]/NET0131 ,
		_w1863_,
		_w8992_,
		_w8994_
	);
	LUT4 #(
		.INIT('h153f)
	) name7645 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1689_,
		_w1702_,
		_w8995_
	);
	LUT4 #(
		.INIT('h135f)
	) name7646 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1692_,
		_w1709_,
		_w8996_
	);
	LUT4 #(
		.INIT('h153f)
	) name7647 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1691_,
		_w1705_,
		_w8997_
	);
	LUT4 #(
		.INIT('h153f)
	) name7648 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[13][7]/NET0131 ,
		_w1694_,
		_w1703_,
		_w8998_
	);
	LUT4 #(
		.INIT('h8000)
	) name7649 (
		_w8997_,
		_w8998_,
		_w8995_,
		_w8996_,
		_w8999_
	);
	LUT4 #(
		.INIT('h135f)
	) name7650 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1699_,
		_w1711_,
		_w9000_
	);
	LUT4 #(
		.INIT('h153f)
	) name7651 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[15][7]/NET0131 ,
		_w1698_,
		_w1712_,
		_w9001_
	);
	LUT4 #(
		.INIT('h135f)
	) name7652 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1696_,
		_w1688_,
		_w9002_
	);
	LUT4 #(
		.INIT('h135f)
	) name7653 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1708_,
		_w1706_,
		_w9003_
	);
	LUT4 #(
		.INIT('h8000)
	) name7654 (
		_w9002_,
		_w9003_,
		_w9000_,
		_w9001_,
		_w9004_
	);
	LUT4 #(
		.INIT('h153f)
	) name7655 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1709_,
		_w1711_,
		_w9005_
	);
	LUT4 #(
		.INIT('h135f)
	) name7656 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1694_,
		_w1692_,
		_w9006_
	);
	LUT4 #(
		.INIT('h135f)
	) name7657 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1712_,
		_w1703_,
		_w9007_
	);
	LUT4 #(
		.INIT('h135f)
	) name7658 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1696_,
		_w1691_,
		_w9008_
	);
	LUT4 #(
		.INIT('h8000)
	) name7659 (
		_w9007_,
		_w9008_,
		_w9005_,
		_w9006_,
		_w9009_
	);
	LUT4 #(
		.INIT('h135f)
	) name7660 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1699_,
		_w1688_,
		_w9010_
	);
	LUT4 #(
		.INIT('h153f)
	) name7661 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1702_,
		_w1705_,
		_w9011_
	);
	LUT4 #(
		.INIT('h135f)
	) name7662 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w1698_,
		_w1708_,
		_w9012_
	);
	LUT4 #(
		.INIT('h153f)
	) name7663 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1689_,
		_w1706_,
		_w9013_
	);
	LUT4 #(
		.INIT('h8000)
	) name7664 (
		_w9012_,
		_w9013_,
		_w9010_,
		_w9011_,
		_w9014_
	);
	LUT4 #(
		.INIT('h0777)
	) name7665 (
		_w8999_,
		_w9004_,
		_w9009_,
		_w9014_,
		_w9015_
	);
	LUT4 #(
		.INIT('h153f)
	) name7666 (
		\P1_InstQueue_reg[7][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1691_,
		_w1702_,
		_w9016_
	);
	LUT4 #(
		.INIT('h135f)
	) name7667 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9017_
	);
	LUT4 #(
		.INIT('h153f)
	) name7668 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1709_,
		_w1703_,
		_w9018_
	);
	LUT4 #(
		.INIT('h153f)
	) name7669 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9019_
	);
	LUT4 #(
		.INIT('h8000)
	) name7670 (
		_w9018_,
		_w9019_,
		_w9016_,
		_w9017_,
		_w9020_
	);
	LUT4 #(
		.INIT('h135f)
	) name7671 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1708_,
		_w1706_,
		_w9021_
	);
	LUT4 #(
		.INIT('h135f)
	) name7672 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1711_,
		_w1705_,
		_w9022_
	);
	LUT4 #(
		.INIT('h153f)
	) name7673 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9023_
	);
	LUT4 #(
		.INIT('h135f)
	) name7674 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1696_,
		_w1699_,
		_w9024_
	);
	LUT4 #(
		.INIT('h8000)
	) name7675 (
		_w9023_,
		_w9024_,
		_w9021_,
		_w9022_,
		_w9025_
	);
	LUT2 #(
		.INIT('h8)
	) name7676 (
		_w9020_,
		_w9025_,
		_w9026_
	);
	LUT4 #(
		.INIT('h135f)
	) name7677 (
		\P1_InstQueue_reg[15][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1696_,
		_w1709_,
		_w9027_
	);
	LUT4 #(
		.INIT('h135f)
	) name7678 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1694_,
		_w1692_,
		_w9028_
	);
	LUT4 #(
		.INIT('h153f)
	) name7679 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1691_,
		_w1712_,
		_w9029_
	);
	LUT4 #(
		.INIT('h135f)
	) name7680 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[13][2]/NET0131 ,
		_w1711_,
		_w1703_,
		_w9030_
	);
	LUT4 #(
		.INIT('h8000)
	) name7681 (
		_w9029_,
		_w9030_,
		_w9027_,
		_w9028_,
		_w9031_
	);
	LUT4 #(
		.INIT('h153f)
	) name7682 (
		\P1_InstQueue_reg[3][2]/NET0131 ,
		\P1_InstQueue_reg[4][2]/NET0131 ,
		_w1688_,
		_w1706_,
		_w9032_
	);
	LUT4 #(
		.INIT('h153f)
	) name7683 (
		\P1_InstQueue_reg[1][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1702_,
		_w1705_,
		_w9033_
	);
	LUT4 #(
		.INIT('h135f)
	) name7684 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[11][2]/NET0131 ,
		_w1698_,
		_w1708_,
		_w9034_
	);
	LUT4 #(
		.INIT('h135f)
	) name7685 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1699_,
		_w1689_,
		_w9035_
	);
	LUT4 #(
		.INIT('h8000)
	) name7686 (
		_w9034_,
		_w9035_,
		_w9032_,
		_w9033_,
		_w9036_
	);
	LUT2 #(
		.INIT('h8)
	) name7687 (
		_w9031_,
		_w9036_,
		_w9037_
	);
	LUT3 #(
		.INIT('h02)
	) name7688 (
		_w9015_,
		_w9026_,
		_w9037_,
		_w9038_
	);
	LUT4 #(
		.INIT('h153f)
	) name7689 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1691_,
		_w1702_,
		_w9039_
	);
	LUT4 #(
		.INIT('h135f)
	) name7690 (
		\P1_InstQueue_reg[4][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9040_
	);
	LUT4 #(
		.INIT('h153f)
	) name7691 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1709_,
		_w1703_,
		_w9041_
	);
	LUT4 #(
		.INIT('h153f)
	) name7692 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9042_
	);
	LUT4 #(
		.INIT('h8000)
	) name7693 (
		_w9041_,
		_w9042_,
		_w9039_,
		_w9040_,
		_w9043_
	);
	LUT4 #(
		.INIT('h153f)
	) name7694 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[2][3]/NET0131 ,
		_w1699_,
		_w1708_,
		_w9044_
	);
	LUT4 #(
		.INIT('h135f)
	) name7695 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w1711_,
		_w1705_,
		_w9045_
	);
	LUT4 #(
		.INIT('h153f)
	) name7696 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[14][3]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9046_
	);
	LUT4 #(
		.INIT('h135f)
	) name7697 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1696_,
		_w1706_,
		_w9047_
	);
	LUT4 #(
		.INIT('h8000)
	) name7698 (
		_w9046_,
		_w9047_,
		_w9044_,
		_w9045_,
		_w9048_
	);
	LUT2 #(
		.INIT('h8)
	) name7699 (
		_w9043_,
		_w9048_,
		_w9049_
	);
	LUT4 #(
		.INIT('h0002)
	) name7700 (
		_w9015_,
		_w9026_,
		_w9037_,
		_w9049_,
		_w9050_
	);
	LUT4 #(
		.INIT('h153f)
	) name7701 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1702_,
		_w1703_,
		_w9051_
	);
	LUT4 #(
		.INIT('h135f)
	) name7702 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9052_
	);
	LUT4 #(
		.INIT('h153f)
	) name7703 (
		\P1_InstQueue_reg[6][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1691_,
		_w1709_,
		_w9053_
	);
	LUT4 #(
		.INIT('h153f)
	) name7704 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9054_
	);
	LUT4 #(
		.INIT('h8000)
	) name7705 (
		_w9053_,
		_w9054_,
		_w9051_,
		_w9052_,
		_w9055_
	);
	LUT4 #(
		.INIT('h153f)
	) name7706 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w1699_,
		_w1708_,
		_w9056_
	);
	LUT4 #(
		.INIT('h135f)
	) name7707 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1696_,
		_w1705_,
		_w9057_
	);
	LUT4 #(
		.INIT('h153f)
	) name7708 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[14][4]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9058_
	);
	LUT4 #(
		.INIT('h135f)
	) name7709 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1711_,
		_w1706_,
		_w9059_
	);
	LUT4 #(
		.INIT('h8000)
	) name7710 (
		_w9058_,
		_w9059_,
		_w9056_,
		_w9057_,
		_w9060_
	);
	LUT2 #(
		.INIT('h8)
	) name7711 (
		_w9055_,
		_w9060_,
		_w9061_
	);
	LUT4 #(
		.INIT('h153f)
	) name7712 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1702_,
		_w1703_,
		_w9062_
	);
	LUT4 #(
		.INIT('h135f)
	) name7713 (
		\P1_InstQueue_reg[4][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9063_
	);
	LUT4 #(
		.INIT('h153f)
	) name7714 (
		\P1_InstQueue_reg[6][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1691_,
		_w1709_,
		_w9064_
	);
	LUT4 #(
		.INIT('h153f)
	) name7715 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9065_
	);
	LUT4 #(
		.INIT('h8000)
	) name7716 (
		_w9064_,
		_w9065_,
		_w9062_,
		_w9063_,
		_w9066_
	);
	LUT4 #(
		.INIT('h153f)
	) name7717 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1699_,
		_w1708_,
		_w9067_
	);
	LUT4 #(
		.INIT('h135f)
	) name7718 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1696_,
		_w1705_,
		_w9068_
	);
	LUT4 #(
		.INIT('h153f)
	) name7719 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[14][5]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9069_
	);
	LUT4 #(
		.INIT('h135f)
	) name7720 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1711_,
		_w1706_,
		_w9070_
	);
	LUT4 #(
		.INIT('h8000)
	) name7721 (
		_w9069_,
		_w9070_,
		_w9067_,
		_w9068_,
		_w9071_
	);
	LUT2 #(
		.INIT('h8)
	) name7722 (
		_w9066_,
		_w9071_,
		_w9072_
	);
	LUT3 #(
		.INIT('h02)
	) name7723 (
		_w9050_,
		_w9061_,
		_w9072_,
		_w9073_
	);
	LUT4 #(
		.INIT('h153f)
	) name7724 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1702_,
		_w1703_,
		_w9074_
	);
	LUT4 #(
		.INIT('h135f)
	) name7725 (
		\P1_InstQueue_reg[4][6]/NET0131 ,
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9075_
	);
	LUT4 #(
		.INIT('h153f)
	) name7726 (
		\P1_InstQueue_reg[6][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1691_,
		_w1709_,
		_w9076_
	);
	LUT4 #(
		.INIT('h153f)
	) name7727 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9077_
	);
	LUT4 #(
		.INIT('h8000)
	) name7728 (
		_w9076_,
		_w9077_,
		_w9074_,
		_w9075_,
		_w9078_
	);
	LUT4 #(
		.INIT('h153f)
	) name7729 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[2][6]/NET0131 ,
		_w1699_,
		_w1708_,
		_w9079_
	);
	LUT4 #(
		.INIT('h135f)
	) name7730 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1696_,
		_w1705_,
		_w9080_
	);
	LUT4 #(
		.INIT('h153f)
	) name7731 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[14][6]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9081_
	);
	LUT4 #(
		.INIT('h135f)
	) name7732 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1711_,
		_w1706_,
		_w9082_
	);
	LUT4 #(
		.INIT('h8000)
	) name7733 (
		_w9081_,
		_w9082_,
		_w9079_,
		_w9080_,
		_w9083_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		_w9078_,
		_w9083_,
		_w9084_
	);
	LUT4 #(
		.INIT('h0002)
	) name7735 (
		_w9050_,
		_w9061_,
		_w9072_,
		_w9084_,
		_w9085_
	);
	LUT4 #(
		.INIT('h153f)
	) name7736 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1702_,
		_w1703_,
		_w9086_
	);
	LUT4 #(
		.INIT('h135f)
	) name7737 (
		\P1_InstQueue_reg[4][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1688_,
		_w1692_,
		_w9087_
	);
	LUT4 #(
		.INIT('h153f)
	) name7738 (
		\P1_InstQueue_reg[6][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1691_,
		_w1709_,
		_w9088_
	);
	LUT4 #(
		.INIT('h153f)
	) name7739 (
		\P1_InstQueue_reg[12][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1689_,
		_w1712_,
		_w9089_
	);
	LUT4 #(
		.INIT('h8000)
	) name7740 (
		_w9088_,
		_w9089_,
		_w9086_,
		_w9087_,
		_w9090_
	);
	LUT4 #(
		.INIT('h153f)
	) name7741 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[2][7]/NET0131 ,
		_w1699_,
		_w1708_,
		_w9091_
	);
	LUT4 #(
		.INIT('h135f)
	) name7742 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[1][7]/NET0131 ,
		_w1696_,
		_w1705_,
		_w9092_
	);
	LUT4 #(
		.INIT('h153f)
	) name7743 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[14][7]/NET0131 ,
		_w1694_,
		_w1698_,
		_w9093_
	);
	LUT4 #(
		.INIT('h135f)
	) name7744 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1711_,
		_w1706_,
		_w9094_
	);
	LUT4 #(
		.INIT('h8000)
	) name7745 (
		_w9093_,
		_w9094_,
		_w9091_,
		_w9092_,
		_w9095_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		_w9090_,
		_w9095_,
		_w9096_
	);
	LUT4 #(
		.INIT('h0111)
	) name7747 (
		_w1842_,
		_w1845_,
		_w9090_,
		_w9095_,
		_w9097_
	);
	LUT3 #(
		.INIT('h80)
	) name7748 (
		_w1814_,
		_w9085_,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h1)
	) name7749 (
		_w8994_,
		_w9098_,
		_w9099_
	);
	LUT4 #(
		.INIT('hb700)
	) name7750 (
		\P1_EBX_reg[31]/NET0131 ,
		_w1829_,
		_w8991_,
		_w9099_,
		_w9100_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name7751 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9101_
	);
	LUT4 #(
		.INIT('hfc20)
	) name7752 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9102_
	);
	LUT2 #(
		.INIT('h2)
	) name7753 (
		\P1_EBX_reg[31]/NET0131 ,
		_w9102_,
		_w9103_
	);
	LUT3 #(
		.INIT('hf2)
	) name7754 (
		_w1933_,
		_w9100_,
		_w9103_,
		_w9104_
	);
	LUT4 #(
		.INIT('hc444)
	) name7755 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9105_
	);
	LUT4 #(
		.INIT('h0888)
	) name7756 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[24]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9106_
	);
	LUT3 #(
		.INIT('ha8)
	) name7757 (
		_w2250_,
		_w9105_,
		_w9106_,
		_w9107_
	);
	LUT4 #(
		.INIT('hc444)
	) name7758 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[16]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9108_
	);
	LUT4 #(
		.INIT('h0888)
	) name7759 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[16]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9109_
	);
	LUT2 #(
		.INIT('h1)
	) name7760 (
		_w9108_,
		_w9109_,
		_w9110_
	);
	LUT3 #(
		.INIT('ha8)
	) name7761 (
		_w2264_,
		_w9108_,
		_w9109_,
		_w9111_
	);
	LUT3 #(
		.INIT('ha8)
	) name7762 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9107_,
		_w9111_,
		_w9112_
	);
	LUT4 #(
		.INIT('hc444)
	) name7763 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9113_
	);
	LUT4 #(
		.INIT('h0888)
	) name7764 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[0]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9114_
	);
	LUT2 #(
		.INIT('h1)
	) name7765 (
		_w9113_,
		_w9114_,
		_w9115_
	);
	LUT3 #(
		.INIT('h02)
	) name7766 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w2271_,
		_w2272_,
		_w9116_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7767 (
		_w2273_,
		_w9113_,
		_w9114_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h1)
	) name7768 (
		_w2280_,
		_w9117_,
		_w9118_
	);
	LUT3 #(
		.INIT('ha8)
	) name7769 (
		_w1679_,
		_w9112_,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h2)
	) name7770 (
		_w2283_,
		_w9117_,
		_w9120_
	);
	LUT4 #(
		.INIT('hc055)
	) name7771 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2272_,
		_w9121_
	);
	LUT2 #(
		.INIT('h2)
	) name7772 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w2288_,
		_w9122_
	);
	LUT3 #(
		.INIT('h0d)
	) name7773 (
		_w2246_,
		_w9121_,
		_w9122_,
		_w9123_
	);
	LUT2 #(
		.INIT('h4)
	) name7774 (
		_w9120_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('hb)
	) name7775 (
		_w9119_,
		_w9124_,
		_w9125_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name7776 (
		_w1945_,
		_w2141_,
		_w2138_,
		_w2149_,
		_w9126_
	);
	LUT4 #(
		.INIT('h0880)
	) name7777 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w9127_
	);
	LUT3 #(
		.INIT('ha8)
	) name7778 (
		_w2216_,
		_w2220_,
		_w9127_,
		_w9128_
	);
	LUT4 #(
		.INIT('hfffc)
	) name7779 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9129_
	);
	LUT4 #(
		.INIT('h9f15)
	) name7780 (
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1953_,
		_w2215_,
		_w8476_,
		_w9130_
	);
	LUT2 #(
		.INIT('h4)
	) name7781 (
		_w9128_,
		_w9130_,
		_w9131_
	);
	LUT2 #(
		.INIT('hb)
	) name7782 (
		_w9126_,
		_w9131_,
		_w9132_
	);
	LUT4 #(
		.INIT('h0880)
	) name7783 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w9133_
	);
	LUT3 #(
		.INIT('ha8)
	) name7784 (
		_w2205_,
		_w2206_,
		_w9133_,
		_w9134_
	);
	LUT4 #(
		.INIT('h9f15)
	) name7785 (
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1440_,
		_w2246_,
		_w8482_,
		_w9135_
	);
	LUT2 #(
		.INIT('h4)
	) name7786 (
		_w9134_,
		_w9135_,
		_w9136_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7787 (
		_w1599_,
		_w1619_,
		_w1678_,
		_w9136_,
		_w9137_
	);
	LUT3 #(
		.INIT('ha8)
	) name7788 (
		_w2315_,
		_w9105_,
		_w9106_,
		_w9138_
	);
	LUT3 #(
		.INIT('ha8)
	) name7789 (
		_w2317_,
		_w9108_,
		_w9109_,
		_w9139_
	);
	LUT3 #(
		.INIT('ha8)
	) name7790 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9138_,
		_w9139_,
		_w9140_
	);
	LUT3 #(
		.INIT('h02)
	) name7791 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w2320_,
		_w2322_,
		_w9141_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7792 (
		_w2323_,
		_w9113_,
		_w9114_,
		_w9141_,
		_w9142_
	);
	LUT2 #(
		.INIT('h1)
	) name7793 (
		_w2327_,
		_w9142_,
		_w9143_
	);
	LUT3 #(
		.INIT('ha8)
	) name7794 (
		_w1679_,
		_w9140_,
		_w9143_,
		_w9144_
	);
	LUT2 #(
		.INIT('h2)
	) name7795 (
		_w2283_,
		_w9142_,
		_w9145_
	);
	LUT4 #(
		.INIT('hc055)
	) name7796 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2320_,
		_w9146_
	);
	LUT2 #(
		.INIT('h2)
	) name7797 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		_w2288_,
		_w9147_
	);
	LUT3 #(
		.INIT('h0d)
	) name7798 (
		_w2246_,
		_w9146_,
		_w9147_,
		_w9148_
	);
	LUT2 #(
		.INIT('h4)
	) name7799 (
		_w9145_,
		_w9148_,
		_w9149_
	);
	LUT2 #(
		.INIT('hb)
	) name7800 (
		_w9144_,
		_w9149_,
		_w9150_
	);
	LUT3 #(
		.INIT('ha8)
	) name7801 (
		_w2250_,
		_w9108_,
		_w9109_,
		_w9151_
	);
	LUT3 #(
		.INIT('ha8)
	) name7802 (
		_w2349_,
		_w9105_,
		_w9106_,
		_w9152_
	);
	LUT3 #(
		.INIT('ha8)
	) name7803 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9151_,
		_w9152_,
		_w9153_
	);
	LUT3 #(
		.INIT('h02)
	) name7804 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w2271_,
		_w2264_,
		_w9154_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7805 (
		_w2346_,
		_w9113_,
		_w9114_,
		_w9154_,
		_w9155_
	);
	LUT2 #(
		.INIT('h1)
	) name7806 (
		_w2351_,
		_w9155_,
		_w9156_
	);
	LUT3 #(
		.INIT('ha8)
	) name7807 (
		_w1679_,
		_w9153_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h2)
	) name7808 (
		_w2283_,
		_w9155_,
		_w9158_
	);
	LUT4 #(
		.INIT('hc055)
	) name7809 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2271_,
		_w9159_
	);
	LUT2 #(
		.INIT('h2)
	) name7810 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		_w2288_,
		_w9160_
	);
	LUT3 #(
		.INIT('h0d)
	) name7811 (
		_w2246_,
		_w9159_,
		_w9160_,
		_w9161_
	);
	LUT2 #(
		.INIT('h4)
	) name7812 (
		_w9158_,
		_w9161_,
		_w9162_
	);
	LUT2 #(
		.INIT('hb)
	) name7813 (
		_w9157_,
		_w9162_,
		_w9163_
	);
	LUT3 #(
		.INIT('ha8)
	) name7814 (
		_w2264_,
		_w9105_,
		_w9106_,
		_w9164_
	);
	LUT3 #(
		.INIT('ha8)
	) name7815 (
		_w2271_,
		_w9108_,
		_w9109_,
		_w9165_
	);
	LUT3 #(
		.INIT('ha8)
	) name7816 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9164_,
		_w9165_,
		_w9166_
	);
	LUT3 #(
		.INIT('h02)
	) name7817 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w2272_,
		_w2376_,
		_w9167_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7818 (
		_w2377_,
		_w9113_,
		_w9114_,
		_w9167_,
		_w9168_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		_w2380_,
		_w9168_,
		_w9169_
	);
	LUT3 #(
		.INIT('ha8)
	) name7820 (
		_w1679_,
		_w9166_,
		_w9169_,
		_w9170_
	);
	LUT2 #(
		.INIT('h2)
	) name7821 (
		_w2283_,
		_w9168_,
		_w9171_
	);
	LUT4 #(
		.INIT('hc055)
	) name7822 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2376_,
		_w9172_
	);
	LUT2 #(
		.INIT('h2)
	) name7823 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		_w2288_,
		_w9173_
	);
	LUT3 #(
		.INIT('h0d)
	) name7824 (
		_w2246_,
		_w9172_,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('h4)
	) name7825 (
		_w9171_,
		_w9174_,
		_w9175_
	);
	LUT2 #(
		.INIT('hb)
	) name7826 (
		_w9170_,
		_w9175_,
		_w9176_
	);
	LUT3 #(
		.INIT('ha8)
	) name7827 (
		_w2271_,
		_w9105_,
		_w9106_,
		_w9177_
	);
	LUT3 #(
		.INIT('ha8)
	) name7828 (
		_w2272_,
		_w9108_,
		_w9109_,
		_w9178_
	);
	LUT3 #(
		.INIT('ha8)
	) name7829 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9177_,
		_w9178_,
		_w9179_
	);
	LUT3 #(
		.INIT('h02)
	) name7830 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w2315_,
		_w2376_,
		_w9180_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7831 (
		_w2402_,
		_w9113_,
		_w9114_,
		_w9180_,
		_w9181_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		_w2405_,
		_w9181_,
		_w9182_
	);
	LUT3 #(
		.INIT('ha8)
	) name7833 (
		_w1679_,
		_w9179_,
		_w9182_,
		_w9183_
	);
	LUT2 #(
		.INIT('h2)
	) name7834 (
		_w2283_,
		_w9181_,
		_w9184_
	);
	LUT4 #(
		.INIT('hc055)
	) name7835 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2315_,
		_w9185_
	);
	LUT2 #(
		.INIT('h2)
	) name7836 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		_w2288_,
		_w9186_
	);
	LUT3 #(
		.INIT('h0d)
	) name7837 (
		_w2246_,
		_w9185_,
		_w9186_,
		_w9187_
	);
	LUT2 #(
		.INIT('h4)
	) name7838 (
		_w9184_,
		_w9187_,
		_w9188_
	);
	LUT2 #(
		.INIT('hb)
	) name7839 (
		_w9183_,
		_w9188_,
		_w9189_
	);
	LUT3 #(
		.INIT('ha8)
	) name7840 (
		_w2272_,
		_w9105_,
		_w9106_,
		_w9190_
	);
	LUT3 #(
		.INIT('ha8)
	) name7841 (
		_w2376_,
		_w9108_,
		_w9109_,
		_w9191_
	);
	LUT3 #(
		.INIT('ha8)
	) name7842 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9190_,
		_w9191_,
		_w9192_
	);
	LUT3 #(
		.INIT('h02)
	) name7843 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w2315_,
		_w2317_,
		_w9193_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7844 (
		_w2326_,
		_w9113_,
		_w9114_,
		_w9193_,
		_w9194_
	);
	LUT2 #(
		.INIT('h1)
	) name7845 (
		_w2429_,
		_w9194_,
		_w9195_
	);
	LUT3 #(
		.INIT('ha8)
	) name7846 (
		_w1679_,
		_w9192_,
		_w9195_,
		_w9196_
	);
	LUT2 #(
		.INIT('h2)
	) name7847 (
		_w2283_,
		_w9194_,
		_w9197_
	);
	LUT4 #(
		.INIT('hc055)
	) name7848 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2317_,
		_w9198_
	);
	LUT2 #(
		.INIT('h2)
	) name7849 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		_w2288_,
		_w9199_
	);
	LUT3 #(
		.INIT('h0d)
	) name7850 (
		_w2246_,
		_w9198_,
		_w9199_,
		_w9200_
	);
	LUT2 #(
		.INIT('h4)
	) name7851 (
		_w9197_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('hb)
	) name7852 (
		_w9196_,
		_w9201_,
		_w9202_
	);
	LUT3 #(
		.INIT('ha8)
	) name7853 (
		_w2376_,
		_w9105_,
		_w9106_,
		_w9203_
	);
	LUT3 #(
		.INIT('ha8)
	) name7854 (
		_w2315_,
		_w9108_,
		_w9109_,
		_w9204_
	);
	LUT3 #(
		.INIT('ha8)
	) name7855 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9203_,
		_w9204_,
		_w9205_
	);
	LUT3 #(
		.INIT('h02)
	) name7856 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w2322_,
		_w2317_,
		_w9206_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7857 (
		_w2451_,
		_w9113_,
		_w9114_,
		_w9206_,
		_w9207_
	);
	LUT2 #(
		.INIT('h1)
	) name7858 (
		_w2454_,
		_w9207_,
		_w9208_
	);
	LUT3 #(
		.INIT('ha8)
	) name7859 (
		_w1679_,
		_w9205_,
		_w9208_,
		_w9209_
	);
	LUT2 #(
		.INIT('h2)
	) name7860 (
		_w2283_,
		_w9207_,
		_w9210_
	);
	LUT4 #(
		.INIT('hc055)
	) name7861 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2322_,
		_w9211_
	);
	LUT2 #(
		.INIT('h2)
	) name7862 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w2288_,
		_w9212_
	);
	LUT3 #(
		.INIT('h0d)
	) name7863 (
		_w2246_,
		_w9211_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h4)
	) name7864 (
		_w9210_,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('hb)
	) name7865 (
		_w9209_,
		_w9214_,
		_w9215_
	);
	LUT3 #(
		.INIT('ha8)
	) name7866 (
		_w2317_,
		_w9105_,
		_w9106_,
		_w9216_
	);
	LUT3 #(
		.INIT('ha8)
	) name7867 (
		_w2322_,
		_w9108_,
		_w9109_,
		_w9217_
	);
	LUT3 #(
		.INIT('ha8)
	) name7868 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9216_,
		_w9217_,
		_w9218_
	);
	LUT3 #(
		.INIT('h02)
	) name7869 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w2320_,
		_w2473_,
		_w9219_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7870 (
		_w2474_,
		_w9113_,
		_w9114_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w2477_,
		_w9220_,
		_w9221_
	);
	LUT3 #(
		.INIT('ha8)
	) name7872 (
		_w1679_,
		_w9218_,
		_w9221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h2)
	) name7873 (
		_w2283_,
		_w9220_,
		_w9223_
	);
	LUT4 #(
		.INIT('hc055)
	) name7874 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2473_,
		_w9224_
	);
	LUT2 #(
		.INIT('h2)
	) name7875 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w2288_,
		_w9225_
	);
	LUT3 #(
		.INIT('h0d)
	) name7876 (
		_w2246_,
		_w9224_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h4)
	) name7877 (
		_w9223_,
		_w9226_,
		_w9227_
	);
	LUT2 #(
		.INIT('hb)
	) name7878 (
		_w9222_,
		_w9227_,
		_w9228_
	);
	LUT3 #(
		.INIT('ha8)
	) name7879 (
		_w2320_,
		_w9108_,
		_w9109_,
		_w9229_
	);
	LUT3 #(
		.INIT('ha8)
	) name7880 (
		_w2322_,
		_w9105_,
		_w9106_,
		_w9230_
	);
	LUT3 #(
		.INIT('ha8)
	) name7881 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9229_,
		_w9230_,
		_w9231_
	);
	LUT3 #(
		.INIT('h02)
	) name7882 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w2473_,
		_w2502_,
		_w9232_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7883 (
		_w2503_,
		_w9113_,
		_w9114_,
		_w9232_,
		_w9233_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w2506_,
		_w9233_,
		_w9234_
	);
	LUT3 #(
		.INIT('ha8)
	) name7885 (
		_w1679_,
		_w9231_,
		_w9234_,
		_w9235_
	);
	LUT2 #(
		.INIT('h2)
	) name7886 (
		_w2283_,
		_w9233_,
		_w9236_
	);
	LUT4 #(
		.INIT('hc055)
	) name7887 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2502_,
		_w9237_
	);
	LUT2 #(
		.INIT('h2)
	) name7888 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w2288_,
		_w9238_
	);
	LUT3 #(
		.INIT('h0d)
	) name7889 (
		_w2246_,
		_w9237_,
		_w9238_,
		_w9239_
	);
	LUT2 #(
		.INIT('h4)
	) name7890 (
		_w9236_,
		_w9239_,
		_w9240_
	);
	LUT2 #(
		.INIT('hb)
	) name7891 (
		_w9235_,
		_w9240_,
		_w9241_
	);
	LUT3 #(
		.INIT('ha8)
	) name7892 (
		_w2320_,
		_w9105_,
		_w9106_,
		_w9242_
	);
	LUT3 #(
		.INIT('ha8)
	) name7893 (
		_w2473_,
		_w9108_,
		_w9109_,
		_w9243_
	);
	LUT3 #(
		.INIT('ha8)
	) name7894 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9242_,
		_w9243_,
		_w9244_
	);
	LUT3 #(
		.INIT('h02)
	) name7895 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w2502_,
		_w2528_,
		_w9245_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7896 (
		_w2529_,
		_w9113_,
		_w9114_,
		_w9245_,
		_w9246_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		_w2532_,
		_w9246_,
		_w9247_
	);
	LUT3 #(
		.INIT('ha8)
	) name7898 (
		_w1679_,
		_w9244_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h2)
	) name7899 (
		_w2283_,
		_w9246_,
		_w9249_
	);
	LUT4 #(
		.INIT('hc055)
	) name7900 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2528_,
		_w9250_
	);
	LUT2 #(
		.INIT('h2)
	) name7901 (
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w2288_,
		_w9251_
	);
	LUT3 #(
		.INIT('h0d)
	) name7902 (
		_w2246_,
		_w9250_,
		_w9251_,
		_w9252_
	);
	LUT2 #(
		.INIT('h4)
	) name7903 (
		_w9249_,
		_w9252_,
		_w9253_
	);
	LUT2 #(
		.INIT('hb)
	) name7904 (
		_w9248_,
		_w9253_,
		_w9254_
	);
	LUT3 #(
		.INIT('ha8)
	) name7905 (
		_w2473_,
		_w9105_,
		_w9106_,
		_w9255_
	);
	LUT3 #(
		.INIT('ha8)
	) name7906 (
		_w2502_,
		_w9108_,
		_w9109_,
		_w9256_
	);
	LUT3 #(
		.INIT('ha8)
	) name7907 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9255_,
		_w9256_,
		_w9257_
	);
	LUT3 #(
		.INIT('h02)
	) name7908 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w2528_,
		_w2554_,
		_w9258_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7909 (
		_w2555_,
		_w9113_,
		_w9114_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h1)
	) name7910 (
		_w2558_,
		_w9259_,
		_w9260_
	);
	LUT3 #(
		.INIT('ha8)
	) name7911 (
		_w1679_,
		_w9257_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h2)
	) name7912 (
		_w2283_,
		_w9259_,
		_w9262_
	);
	LUT4 #(
		.INIT('hc055)
	) name7913 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2554_,
		_w9263_
	);
	LUT2 #(
		.INIT('h2)
	) name7914 (
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w2288_,
		_w9264_
	);
	LUT3 #(
		.INIT('h0d)
	) name7915 (
		_w2246_,
		_w9263_,
		_w9264_,
		_w9265_
	);
	LUT2 #(
		.INIT('h4)
	) name7916 (
		_w9262_,
		_w9265_,
		_w9266_
	);
	LUT2 #(
		.INIT('hb)
	) name7917 (
		_w9261_,
		_w9266_,
		_w9267_
	);
	LUT3 #(
		.INIT('ha8)
	) name7918 (
		_w2502_,
		_w9105_,
		_w9106_,
		_w9268_
	);
	LUT3 #(
		.INIT('ha8)
	) name7919 (
		_w2528_,
		_w9108_,
		_w9109_,
		_w9269_
	);
	LUT3 #(
		.INIT('ha8)
	) name7920 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9268_,
		_w9269_,
		_w9270_
	);
	LUT3 #(
		.INIT('h02)
	) name7921 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w2554_,
		_w2580_,
		_w9271_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7922 (
		_w2581_,
		_w9113_,
		_w9114_,
		_w9271_,
		_w9272_
	);
	LUT2 #(
		.INIT('h1)
	) name7923 (
		_w2584_,
		_w9272_,
		_w9273_
	);
	LUT3 #(
		.INIT('ha8)
	) name7924 (
		_w1679_,
		_w9270_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h2)
	) name7925 (
		_w2283_,
		_w9272_,
		_w9275_
	);
	LUT4 #(
		.INIT('hc055)
	) name7926 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2580_,
		_w9276_
	);
	LUT2 #(
		.INIT('h2)
	) name7927 (
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w2288_,
		_w9277_
	);
	LUT3 #(
		.INIT('h0d)
	) name7928 (
		_w2246_,
		_w9276_,
		_w9277_,
		_w9278_
	);
	LUT2 #(
		.INIT('h4)
	) name7929 (
		_w9275_,
		_w9278_,
		_w9279_
	);
	LUT2 #(
		.INIT('hb)
	) name7930 (
		_w9274_,
		_w9279_,
		_w9280_
	);
	LUT3 #(
		.INIT('ha8)
	) name7931 (
		_w2528_,
		_w9105_,
		_w9106_,
		_w9281_
	);
	LUT3 #(
		.INIT('ha8)
	) name7932 (
		_w2554_,
		_w9108_,
		_w9109_,
		_w9282_
	);
	LUT3 #(
		.INIT('ha8)
	) name7933 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9281_,
		_w9282_,
		_w9283_
	);
	LUT3 #(
		.INIT('h02)
	) name7934 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w2580_,
		_w2606_,
		_w9284_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7935 (
		_w2607_,
		_w9113_,
		_w9114_,
		_w9284_,
		_w9285_
	);
	LUT2 #(
		.INIT('h1)
	) name7936 (
		_w2610_,
		_w9285_,
		_w9286_
	);
	LUT3 #(
		.INIT('ha8)
	) name7937 (
		_w1679_,
		_w9283_,
		_w9286_,
		_w9287_
	);
	LUT2 #(
		.INIT('h2)
	) name7938 (
		_w2283_,
		_w9285_,
		_w9288_
	);
	LUT4 #(
		.INIT('hc055)
	) name7939 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2606_,
		_w9289_
	);
	LUT2 #(
		.INIT('h2)
	) name7940 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w2288_,
		_w9290_
	);
	LUT3 #(
		.INIT('h0d)
	) name7941 (
		_w2246_,
		_w9289_,
		_w9290_,
		_w9291_
	);
	LUT2 #(
		.INIT('h4)
	) name7942 (
		_w9288_,
		_w9291_,
		_w9292_
	);
	LUT2 #(
		.INIT('hb)
	) name7943 (
		_w9287_,
		_w9292_,
		_w9293_
	);
	LUT3 #(
		.INIT('ha8)
	) name7944 (
		_w2554_,
		_w9105_,
		_w9106_,
		_w9294_
	);
	LUT3 #(
		.INIT('ha8)
	) name7945 (
		_w2580_,
		_w9108_,
		_w9109_,
		_w9295_
	);
	LUT3 #(
		.INIT('ha8)
	) name7946 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9294_,
		_w9295_,
		_w9296_
	);
	LUT3 #(
		.INIT('h02)
	) name7947 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w2349_,
		_w2606_,
		_w9297_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7948 (
		_w2632_,
		_w9113_,
		_w9114_,
		_w9297_,
		_w9298_
	);
	LUT2 #(
		.INIT('h1)
	) name7949 (
		_w2635_,
		_w9298_,
		_w9299_
	);
	LUT3 #(
		.INIT('ha8)
	) name7950 (
		_w1679_,
		_w9296_,
		_w9299_,
		_w9300_
	);
	LUT2 #(
		.INIT('h2)
	) name7951 (
		_w2283_,
		_w9298_,
		_w9301_
	);
	LUT4 #(
		.INIT('hc055)
	) name7952 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2349_,
		_w9302_
	);
	LUT2 #(
		.INIT('h2)
	) name7953 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w2288_,
		_w9303_
	);
	LUT3 #(
		.INIT('h0d)
	) name7954 (
		_w2246_,
		_w9302_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('h4)
	) name7955 (
		_w9301_,
		_w9304_,
		_w9305_
	);
	LUT2 #(
		.INIT('hb)
	) name7956 (
		_w9300_,
		_w9305_,
		_w9306_
	);
	LUT3 #(
		.INIT('ha8)
	) name7957 (
		_w2580_,
		_w9105_,
		_w9106_,
		_w9307_
	);
	LUT3 #(
		.INIT('ha8)
	) name7958 (
		_w2606_,
		_w9108_,
		_w9109_,
		_w9308_
	);
	LUT3 #(
		.INIT('ha8)
	) name7959 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9307_,
		_w9308_,
		_w9309_
	);
	LUT3 #(
		.INIT('h02)
	) name7960 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w2250_,
		_w2349_,
		_w9310_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7961 (
		_w2350_,
		_w9113_,
		_w9114_,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h1)
	) name7962 (
		_w2659_,
		_w9311_,
		_w9312_
	);
	LUT3 #(
		.INIT('ha8)
	) name7963 (
		_w1679_,
		_w9309_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h2)
	) name7964 (
		_w2283_,
		_w9311_,
		_w9314_
	);
	LUT4 #(
		.INIT('hc055)
	) name7965 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2250_,
		_w9315_
	);
	LUT2 #(
		.INIT('h2)
	) name7966 (
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w2288_,
		_w9316_
	);
	LUT3 #(
		.INIT('h0d)
	) name7967 (
		_w2246_,
		_w9315_,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h4)
	) name7968 (
		_w9314_,
		_w9317_,
		_w9318_
	);
	LUT2 #(
		.INIT('hb)
	) name7969 (
		_w9313_,
		_w9318_,
		_w9319_
	);
	LUT3 #(
		.INIT('ha8)
	) name7970 (
		_w2606_,
		_w9105_,
		_w9106_,
		_w9320_
	);
	LUT3 #(
		.INIT('ha8)
	) name7971 (
		_w2349_,
		_w9108_,
		_w9109_,
		_w9321_
	);
	LUT3 #(
		.INIT('ha8)
	) name7972 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9320_,
		_w9321_,
		_w9322_
	);
	LUT3 #(
		.INIT('h02)
	) name7973 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w2250_,
		_w2264_,
		_w9323_
	);
	LUT4 #(
		.INIT('h00ab)
	) name7974 (
		_w2279_,
		_w9113_,
		_w9114_,
		_w9323_,
		_w9324_
	);
	LUT2 #(
		.INIT('h1)
	) name7975 (
		_w2683_,
		_w9324_,
		_w9325_
	);
	LUT3 #(
		.INIT('ha8)
	) name7976 (
		_w1679_,
		_w9322_,
		_w9325_,
		_w9326_
	);
	LUT2 #(
		.INIT('h2)
	) name7977 (
		_w2283_,
		_w9324_,
		_w9327_
	);
	LUT4 #(
		.INIT('hc055)
	) name7978 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1455_,
		_w1468_,
		_w2264_,
		_w9328_
	);
	LUT2 #(
		.INIT('h2)
	) name7979 (
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w2288_,
		_w9329_
	);
	LUT3 #(
		.INIT('h0d)
	) name7980 (
		_w2246_,
		_w9328_,
		_w9329_,
		_w9330_
	);
	LUT2 #(
		.INIT('h4)
	) name7981 (
		_w9327_,
		_w9330_,
		_w9331_
	);
	LUT2 #(
		.INIT('hb)
	) name7982 (
		_w9326_,
		_w9331_,
		_w9332_
	);
	LUT3 #(
		.INIT('h08)
	) name7983 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w1592_,
		_w1660_,
		_w9333_
	);
	LUT4 #(
		.INIT('haa20)
	) name7984 (
		_w1559_,
		_w7112_,
		_w7114_,
		_w9333_,
		_w9334_
	);
	LUT4 #(
		.INIT('h028a)
	) name7985 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w9335_
	);
	LUT4 #(
		.INIT('h00d7)
	) name7986 (
		_w1659_,
		_w7119_,
		_w7120_,
		_w9335_,
		_w9336_
	);
	LUT4 #(
		.INIT('h8000)
	) name7987 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9337_
	);
	LUT4 #(
		.INIT('h7f80)
	) name7988 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9338_
	);
	LUT3 #(
		.INIT('h78)
	) name7989 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w9339_
	);
	LUT4 #(
		.INIT('hc840)
	) name7990 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w9338_,
		_w9339_,
		_w9340_
	);
	LUT2 #(
		.INIT('h2)
	) name7991 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w5747_,
		_w9341_
	);
	LUT4 #(
		.INIT('h135f)
	) name7992 (
		\P2_rEIP_reg[4]/NET0131 ,
		_w2283_,
		_w2286_,
		_w9338_,
		_w9342_
	);
	LUT3 #(
		.INIT('h10)
	) name7993 (
		_w9340_,
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT4 #(
		.INIT('h8aff)
	) name7994 (
		_w1678_,
		_w9334_,
		_w9336_,
		_w9343_,
		_w9344_
	);
	LUT4 #(
		.INIT('h0880)
	) name7995 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w9345_
	);
	LUT3 #(
		.INIT('ha8)
	) name7996 (
		_w2230_,
		_w2231_,
		_w9345_,
		_w9346_
	);
	LUT4 #(
		.INIT('h9f15)
	) name7997 (
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w1695_,
		_w2248_,
		_w8460_,
		_w9347_
	);
	LUT2 #(
		.INIT('h4)
	) name7998 (
		_w9346_,
		_w9347_,
		_w9348_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7999 (
		_w1900_,
		_w1905_,
		_w1933_,
		_w9348_,
		_w9349_
	);
	LUT2 #(
		.INIT('h2)
	) name8000 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w7422_,
		_w9350_
	);
	LUT3 #(
		.INIT('h87)
	) name8001 (
		_w2818_,
		_w2823_,
		_w2996_,
		_w9351_
	);
	LUT4 #(
		.INIT('hf400)
	) name8002 (
		_w3006_,
		_w3010_,
		_w3011_,
		_w9351_,
		_w9352_
	);
	LUT4 #(
		.INIT('h000b)
	) name8003 (
		_w3006_,
		_w3010_,
		_w3011_,
		_w9351_,
		_w9353_
	);
	LUT3 #(
		.INIT('h02)
	) name8004 (
		_w2181_,
		_w9353_,
		_w9352_,
		_w9354_
	);
	LUT3 #(
		.INIT('h95)
	) name8005 (
		_w2920_,
		_w2818_,
		_w2823_,
		_w9355_
	);
	LUT4 #(
		.INIT('h000b)
	) name8006 (
		_w2796_,
		_w2925_,
		_w4045_,
		_w9355_,
		_w9356_
	);
	LUT4 #(
		.INIT('hf400)
	) name8007 (
		_w2796_,
		_w2925_,
		_w4045_,
		_w9355_,
		_w9357_
	);
	LUT3 #(
		.INIT('h02)
	) name8008 (
		_w2180_,
		_w9357_,
		_w9356_,
		_w9358_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8009 (
		_w1945_,
		_w9350_,
		_w9354_,
		_w9358_,
		_w9359_
	);
	LUT3 #(
		.INIT('h80)
	) name8010 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9360_
	);
	LUT4 #(
		.INIT('h8000)
	) name8011 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9361_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8012 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9362_
	);
	LUT4 #(
		.INIT('hf400)
	) name8013 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w9362_,
		_w9363_
	);
	LUT2 #(
		.INIT('h2)
	) name8014 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w5783_,
		_w9364_
	);
	LUT3 #(
		.INIT('h78)
	) name8015 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w9365_
	);
	LUT3 #(
		.INIT('h80)
	) name8016 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w9365_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name8017 (
		\P3_rEIP_reg[4]/NET0131 ,
		_w3054_,
		_w9367_
	);
	LUT4 #(
		.INIT('h0001)
	) name8018 (
		_w9366_,
		_w9364_,
		_w9363_,
		_w9367_,
		_w9368_
	);
	LUT2 #(
		.INIT('hb)
	) name8019 (
		_w9359_,
		_w9368_,
		_w9369_
	);
	LUT3 #(
		.INIT('h08)
	) name8020 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w1842_,
		_w1915_,
		_w9370_
	);
	LUT4 #(
		.INIT('haa20)
	) name8021 (
		_w1810_,
		_w7061_,
		_w7063_,
		_w9370_,
		_w9371_
	);
	LUT4 #(
		.INIT('h028a)
	) name8022 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w9372_
	);
	LUT4 #(
		.INIT('h007d)
	) name8023 (
		_w1924_,
		_w3342_,
		_w7072_,
		_w9372_,
		_w9373_
	);
	LUT4 #(
		.INIT('h8000)
	) name8024 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9374_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8025 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9375_
	);
	LUT4 #(
		.INIT('hf400)
	) name8026 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3407_,
		_w9375_,
		_w9376_
	);
	LUT2 #(
		.INIT('h2)
	) name8027 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w6383_,
		_w9377_
	);
	LUT3 #(
		.INIT('h78)
	) name8028 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w9378_
	);
	LUT3 #(
		.INIT('h80)
	) name8029 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w9378_,
		_w9379_
	);
	LUT4 #(
		.INIT('h0001)
	) name8030 (
		_w7078_,
		_w9379_,
		_w9377_,
		_w9376_,
		_w9380_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8031 (
		_w1933_,
		_w9371_,
		_w9373_,
		_w9380_,
		_w9381_
	);
	LUT2 #(
		.INIT('h4)
	) name8032 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w9382_
	);
	LUT4 #(
		.INIT('h8008)
	) name8033 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstAddrPointer_reg[0]/NET0131 ,
		\P1_InstAddrPointer_reg[1]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w9383_
	);
	LUT3 #(
		.INIT('ha8)
	) name8034 (
		_w2230_,
		_w9382_,
		_w9383_,
		_w9384_
	);
	LUT4 #(
		.INIT('h9f13)
	) name8035 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P1_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2248_,
		_w8460_,
		_w9385_
	);
	LUT2 #(
		.INIT('h4)
	) name8036 (
		_w9384_,
		_w9385_,
		_w9386_
	);
	LUT4 #(
		.INIT('he0ff)
	) name8037 (
		_w1849_,
		_w1869_,
		_w1933_,
		_w9386_,
		_w9387_
	);
	LUT4 #(
		.INIT('hef00)
	) name8038 (
		_w1884_,
		_w1882_,
		_w1892_,
		_w1933_,
		_w9388_
	);
	LUT2 #(
		.INIT('h4)
	) name8039 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w9389_
	);
	LUT3 #(
		.INIT('ha8)
	) name8040 (
		_w2230_,
		_w9345_,
		_w9389_,
		_w9390_
	);
	LUT4 #(
		.INIT('hcf45)
	) name8041 (
		\P1_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1883_,
		_w2248_,
		_w8460_,
		_w9391_
	);
	LUT2 #(
		.INIT('h4)
	) name8042 (
		_w9390_,
		_w9391_,
		_w9392_
	);
	LUT2 #(
		.INIT('hb)
	) name8043 (
		_w9388_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h4)
	) name8044 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w9394_
	);
	LUT3 #(
		.INIT('ha8)
	) name8045 (
		_w2216_,
		_w9127_,
		_w9394_,
		_w9395_
	);
	LUT4 #(
		.INIT('hcf45)
	) name8046 (
		\P3_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2156_,
		_w2215_,
		_w8476_,
		_w9396_
	);
	LUT2 #(
		.INIT('h4)
	) name8047 (
		_w9395_,
		_w9396_,
		_w9397_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8048 (
		_w1945_,
		_w2155_,
		_w2161_,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h4)
	) name8049 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w9399_
	);
	LUT3 #(
		.INIT('ha8)
	) name8050 (
		_w2205_,
		_w9133_,
		_w9399_,
		_w9400_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8051 (
		\P2_InstQueueRd_Addr_reg[3]/NET0131 ,
		_w1623_,
		_w2246_,
		_w8482_,
		_w9401_
	);
	LUT2 #(
		.INIT('h4)
	) name8052 (
		_w9400_,
		_w9401_,
		_w9402_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name8053 (
		_w1624_,
		_w1637_,
		_w1678_,
		_w9402_,
		_w9403_
	);
	LUT4 #(
		.INIT('h888a)
	) name8054 (
		_w1945_,
		_w2101_,
		_w2118_,
		_w2129_,
		_w9404_
	);
	LUT2 #(
		.INIT('h4)
	) name8055 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w9405_
	);
	LUT4 #(
		.INIT('h8008)
	) name8056 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstAddrPointer_reg[0]/NET0131 ,
		\P3_InstAddrPointer_reg[1]/NET0131 ,
		\P3_InstAddrPointer_reg[31]/NET0131 ,
		_w9406_
	);
	LUT3 #(
		.INIT('ha8)
	) name8057 (
		_w2216_,
		_w9405_,
		_w9406_,
		_w9407_
	);
	LUT4 #(
		.INIT('h9f13)
	) name8058 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P3_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2215_,
		_w8476_,
		_w9408_
	);
	LUT2 #(
		.INIT('h4)
	) name8059 (
		_w9407_,
		_w9408_,
		_w9409_
	);
	LUT2 #(
		.INIT('hb)
	) name8060 (
		_w9404_,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h4)
	) name8061 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w9411_
	);
	LUT4 #(
		.INIT('h8008)
	) name8062 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstAddrPointer_reg[0]/NET0131 ,
		\P2_InstAddrPointer_reg[1]/NET0131 ,
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w9412_
	);
	LUT3 #(
		.INIT('ha8)
	) name8063 (
		_w2205_,
		_w9411_,
		_w9412_,
		_w9413_
	);
	LUT4 #(
		.INIT('h9f13)
	) name8064 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		\P2_InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2246_,
		_w8482_,
		_w9414_
	);
	LUT2 #(
		.INIT('h4)
	) name8065 (
		_w9413_,
		_w9414_,
		_w9415_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name8066 (
		_w1647_,
		_w1650_,
		_w1678_,
		_w9415_,
		_w9416_
	);
	LUT2 #(
		.INIT('h2)
	) name8067 (
		\P1_EAX_reg[26]/NET0131 ,
		_w9102_,
		_w9417_
	);
	LUT4 #(
		.INIT('h8000)
	) name8068 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w9418_
	);
	LUT4 #(
		.INIT('h8000)
	) name8069 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w9418_,
		_w9419_
	);
	LUT4 #(
		.INIT('h8000)
	) name8070 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		\P1_EAX_reg[10]/NET0131 ,
		_w9420_,
		_w9421_
	);
	LUT3 #(
		.INIT('h80)
	) name8072 (
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		_w9420_,
		_w9422_
	);
	LUT4 #(
		.INIT('h8000)
	) name8073 (
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w9420_,
		_w9423_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		\P1_EAX_reg[13]/NET0131 ,
		_w9423_,
		_w9424_
	);
	LUT3 #(
		.INIT('h80)
	) name8075 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		_w9423_,
		_w9425_
	);
	LUT4 #(
		.INIT('h8000)
	) name8076 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		_w9423_,
		_w9426_
	);
	LUT2 #(
		.INIT('h8)
	) name8077 (
		\P1_EAX_reg[16]/NET0131 ,
		_w9426_,
		_w9427_
	);
	LUT2 #(
		.INIT('h8)
	) name8078 (
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[18]/NET0131 ,
		_w9428_
	);
	LUT3 #(
		.INIT('h80)
	) name8079 (
		\P1_EAX_reg[16]/NET0131 ,
		_w9426_,
		_w9428_,
		_w9429_
	);
	LUT4 #(
		.INIT('h8000)
	) name8080 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		_w9426_,
		_w9428_,
		_w9430_
	);
	LUT2 #(
		.INIT('h8)
	) name8081 (
		\P1_EAX_reg[20]/NET0131 ,
		\P1_EAX_reg[21]/NET0131 ,
		_w9431_
	);
	LUT3 #(
		.INIT('h80)
	) name8082 (
		\P1_EAX_reg[20]/NET0131 ,
		\P1_EAX_reg[21]/NET0131 ,
		\P1_EAX_reg[22]/NET0131 ,
		_w9432_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		\P1_EAX_reg[23]/NET0131 ,
		\P1_EAX_reg[24]/NET0131 ,
		_w9433_
	);
	LUT3 #(
		.INIT('h80)
	) name8084 (
		_w9430_,
		_w9432_,
		_w9433_,
		_w9434_
	);
	LUT4 #(
		.INIT('h8000)
	) name8085 (
		\P1_EAX_reg[25]/NET0131 ,
		_w9430_,
		_w9432_,
		_w9433_,
		_w9435_
	);
	LUT4 #(
		.INIT('h00ec)
	) name8086 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w1867_,
		_w9436_
	);
	LUT4 #(
		.INIT('h00fb)
	) name8087 (
		_w1827_,
		_w1854_,
		_w1832_,
		_w1864_,
		_w9437_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8088 (
		_w1827_,
		_w9435_,
		_w9436_,
		_w9437_,
		_w9438_
	);
	LUT3 #(
		.INIT('h40)
	) name8089 (
		\P1_EAX_reg[26]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9439_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8090 (
		_w9015_,
		_w9026_,
		_w9037_,
		_w9049_,
		_w9440_
	);
	LUT3 #(
		.INIT('h02)
	) name8091 (
		_w1846_,
		_w9050_,
		_w9440_,
		_w9441_
	);
	LUT4 #(
		.INIT('h0080)
	) name8092 (
		_w1725_,
		_w1802_,
		_w1867_,
		_w3522_,
		_w9442_
	);
	LUT3 #(
		.INIT('h08)
	) name8093 (
		_w1795_,
		_w1867_,
		_w3449_,
		_w9443_
	);
	LUT4 #(
		.INIT('h0013)
	) name8094 (
		_w1832_,
		_w9442_,
		_w9441_,
		_w9443_,
		_w9444_
	);
	LUT3 #(
		.INIT('h70)
	) name8095 (
		_w9435_,
		_w9439_,
		_w9444_,
		_w9445_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8096 (
		\P1_EAX_reg[26]/NET0131 ,
		_w1933_,
		_w9438_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('he)
	) name8097 (
		_w9417_,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h2)
	) name8098 (
		\P2_uWord_reg[12]/NET0131 ,
		_w7767_,
		_w9448_
	);
	LUT4 #(
		.INIT('h0222)
	) name8099 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[12]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9449_
	);
	LUT4 #(
		.INIT('h3111)
	) name8100 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[12]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9450_
	);
	LUT3 #(
		.INIT('h01)
	) name8101 (
		_w1605_,
		_w9450_,
		_w9449_,
		_w9451_
	);
	LUT2 #(
		.INIT('h8)
	) name8102 (
		_w1565_,
		_w9451_,
		_w9452_
	);
	LUT4 #(
		.INIT('h0001)
	) name8103 (
		\P2_EAX_reg[13]/NET0131 ,
		\P2_EAX_reg[14]/NET0131 ,
		\P2_EAX_reg[15]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		_w9453_
	);
	LUT4 #(
		.INIT('h0001)
	) name8104 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		\P2_EAX_reg[12]/NET0131 ,
		_w9454_
	);
	LUT4 #(
		.INIT('h0001)
	) name8105 (
		\P2_EAX_reg[6]/NET0131 ,
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w9455_
	);
	LUT4 #(
		.INIT('h0001)
	) name8106 (
		\P2_EAX_reg[2]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w9456_
	);
	LUT4 #(
		.INIT('h8000)
	) name8107 (
		_w9455_,
		_w9456_,
		_w9453_,
		_w9454_,
		_w9457_
	);
	LUT4 #(
		.INIT('h0080)
	) name8108 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9457_,
		_w9458_
	);
	LUT4 #(
		.INIT('h8000)
	) name8109 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w9458_,
		_w9459_
	);
	LUT3 #(
		.INIT('h80)
	) name8110 (
		_w7781_,
		_w7783_,
		_w9459_,
		_w9460_
	);
	LUT4 #(
		.INIT('h8000)
	) name8111 (
		_w7781_,
		_w7783_,
		_w7785_,
		_w9459_,
		_w9461_
	);
	LUT2 #(
		.INIT('h8)
	) name8112 (
		\P2_EAX_reg[28]/NET0131 ,
		_w9461_,
		_w9462_
	);
	LUT3 #(
		.INIT('h48)
	) name8113 (
		\P2_EAX_reg[28]/NET0131 ,
		_w1566_,
		_w9461_,
		_w9463_
	);
	LUT3 #(
		.INIT('h54)
	) name8114 (
		_w1602_,
		_w9452_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h2)
	) name8115 (
		_w1566_,
		_w1602_,
		_w9465_
	);
	LUT3 #(
		.INIT('hf1)
	) name8116 (
		_w1565_,
		_w1566_,
		_w1602_,
		_w9466_
	);
	LUT4 #(
		.INIT('h004e)
	) name8117 (
		_w1565_,
		_w1566_,
		_w1605_,
		_w1602_,
		_w9467_
	);
	LUT2 #(
		.INIT('h2)
	) name8118 (
		\P2_uWord_reg[12]/NET0131 ,
		_w9467_,
		_w9468_
	);
	LUT4 #(
		.INIT('heeec)
	) name8119 (
		_w1678_,
		_w9448_,
		_w9464_,
		_w9468_,
		_w9469_
	);
	LUT4 #(
		.INIT('hfc23)
	) name8120 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9470_
	);
	LUT2 #(
		.INIT('h2)
	) name8121 (
		_w1797_,
		_w1852_,
		_w9471_
	);
	LUT3 #(
		.INIT('hf1)
	) name8122 (
		_w1795_,
		_w1797_,
		_w1852_,
		_w9472_
	);
	LUT4 #(
		.INIT('h040e)
	) name8123 (
		_w1795_,
		_w1797_,
		_w1852_,
		_w1861_,
		_w9473_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8124 (
		\P1_uWord_reg[12]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w9474_
	);
	LUT3 #(
		.INIT('h02)
	) name8125 (
		_w1795_,
		_w1861_,
		_w3464_,
		_w9475_
	);
	LUT2 #(
		.INIT('h8)
	) name8126 (
		\P1_EAX_reg[25]/NET0131 ,
		\P1_EAX_reg[26]/NET0131 ,
		_w9476_
	);
	LUT3 #(
		.INIT('h80)
	) name8127 (
		\P1_EAX_reg[25]/NET0131 ,
		\P1_EAX_reg[26]/NET0131 ,
		\P1_EAX_reg[27]/NET0131 ,
		_w9477_
	);
	LUT4 #(
		.INIT('h0001)
	) name8128 (
		\P1_EAX_reg[13]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w9478_
	);
	LUT4 #(
		.INIT('h0001)
	) name8129 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[10]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w9479_
	);
	LUT4 #(
		.INIT('h0001)
	) name8130 (
		\P1_EAX_reg[6]/NET0131 ,
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w9480_
	);
	LUT4 #(
		.INIT('h0001)
	) name8131 (
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w9481_
	);
	LUT4 #(
		.INIT('h8000)
	) name8132 (
		_w9480_,
		_w9481_,
		_w9478_,
		_w9479_,
		_w9482_
	);
	LUT4 #(
		.INIT('h0080)
	) name8133 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9482_,
		_w9483_
	);
	LUT4 #(
		.INIT('h8000)
	) name8134 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		_w9431_,
		_w9483_,
		_w9484_
	);
	LUT2 #(
		.INIT('h8)
	) name8135 (
		\P1_EAX_reg[22]/NET0131 ,
		_w9484_,
		_w9485_
	);
	LUT3 #(
		.INIT('h80)
	) name8136 (
		\P1_EAX_reg[22]/NET0131 ,
		_w9433_,
		_w9484_,
		_w9486_
	);
	LUT4 #(
		.INIT('h8000)
	) name8137 (
		\P1_EAX_reg[22]/NET0131 ,
		_w9433_,
		_w9477_,
		_w9484_,
		_w9487_
	);
	LUT3 #(
		.INIT('h48)
	) name8138 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1797_,
		_w9487_,
		_w9488_
	);
	LUT3 #(
		.INIT('hd0)
	) name8139 (
		_w1842_,
		_w1851_,
		_w1933_,
		_w9489_
	);
	LUT3 #(
		.INIT('he0)
	) name8140 (
		_w9475_,
		_w9488_,
		_w9489_,
		_w9490_
	);
	LUT2 #(
		.INIT('he)
	) name8141 (
		_w9474_,
		_w9490_,
		_w9491_
	);
	LUT2 #(
		.INIT('h2)
	) name8142 (
		\P3_EAX_reg[26]/NET0131 ,
		_w8341_,
		_w9492_
	);
	LUT3 #(
		.INIT('h48)
	) name8143 (
		\P3_EAX_reg[26]/NET0131 ,
		_w8361_,
		_w8360_,
		_w9493_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8144 (
		\P3_EAX_reg[26]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w9494_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8145 (
		_w8391_,
		_w8402_,
		_w8413_,
		_w8425_,
		_w9495_
	);
	LUT3 #(
		.INIT('h02)
	) name8146 (
		_w2098_,
		_w8426_,
		_w9495_,
		_w9496_
	);
	LUT2 #(
		.INIT('h8)
	) name8147 (
		_w2087_,
		_w9496_,
		_w9497_
	);
	LUT3 #(
		.INIT('h80)
	) name8148 (
		\buf2_reg[26]/NET0131 ,
		_w2060_,
		_w2044_,
		_w9498_
	);
	LUT3 #(
		.INIT('h20)
	) name8149 (
		\buf2_reg[10]/NET0131 ,
		_w2060_,
		_w2047_,
		_w9499_
	);
	LUT3 #(
		.INIT('ha8)
	) name8150 (
		_w2119_,
		_w9498_,
		_w9499_,
		_w9500_
	);
	LUT2 #(
		.INIT('h1)
	) name8151 (
		_w9497_,
		_w9500_,
		_w9501_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8152 (
		_w1945_,
		_w9493_,
		_w9494_,
		_w9501_,
		_w9502_
	);
	LUT2 #(
		.INIT('he)
	) name8153 (
		_w9492_,
		_w9502_,
		_w9503_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name8154 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2084_,
		_w8920_,
		_w8921_,
		_w9504_
	);
	LUT3 #(
		.INIT('ha8)
	) name8155 (
		\P3_EBX_reg[30]/NET0131 ,
		_w8925_,
		_w9504_,
		_w9505_
	);
	LUT3 #(
		.INIT('h90)
	) name8156 (
		_w8879_,
		_w8890_,
		_w8923_,
		_w9506_
	);
	LUT3 #(
		.INIT('h40)
	) name8157 (
		\P3_EBX_reg[30]/NET0131 ,
		_w2075_,
		_w2083_,
		_w9507_
	);
	LUT4 #(
		.INIT('h8000)
	) name8158 (
		\P3_EBX_reg[25]/NET0131 ,
		_w8920_,
		_w8921_,
		_w9507_,
		_w9508_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		_w9506_,
		_w9508_,
		_w9509_
	);
	LUT2 #(
		.INIT('h2)
	) name8160 (
		\P3_EBX_reg[30]/NET0131 ,
		_w8341_,
		_w9510_
	);
	LUT4 #(
		.INIT('hff8a)
	) name8161 (
		_w1945_,
		_w9505_,
		_w9509_,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h2)
	) name8162 (
		\P2_EAX_reg[26]/NET0131 ,
		_w7767_,
		_w9512_
	);
	LUT3 #(
		.INIT('h60)
	) name8163 (
		\P2_EAX_reg[26]/NET0131 ,
		_w7784_,
		_w7789_,
		_w9513_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8164 (
		\P2_EAX_reg[26]/NET0131 ,
		_w1604_,
		_w1642_,
		_w7790_,
		_w9514_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name8165 (
		\P2_EAX_reg[26]/NET0131 ,
		_w1592_,
		_w1605_,
		_w1601_,
		_w9515_
	);
	LUT3 #(
		.INIT('hd1)
	) name8166 (
		\P2_EAX_reg[26]/NET0131 ,
		_w1606_,
		_w5478_,
		_w9516_
	);
	LUT3 #(
		.INIT('h08)
	) name8167 (
		_w1501_,
		_w1568_,
		_w9516_,
		_w9517_
	);
	LUT4 #(
		.INIT('hfd00)
	) name8168 (
		_w7815_,
		_w7826_,
		_w7837_,
		_w7849_,
		_w9518_
	);
	LUT3 #(
		.INIT('h02)
	) name8169 (
		_w1596_,
		_w7850_,
		_w9518_,
		_w9519_
	);
	LUT4 #(
		.INIT('h0222)
	) name8170 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[10]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9520_
	);
	LUT4 #(
		.INIT('h3111)
	) name8171 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[10]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9521_
	);
	LUT3 #(
		.INIT('h01)
	) name8172 (
		_w1605_,
		_w9521_,
		_w9520_,
		_w9522_
	);
	LUT3 #(
		.INIT('h23)
	) name8173 (
		_w1602_,
		_w9515_,
		_w9522_,
		_w9523_
	);
	LUT2 #(
		.INIT('h2)
	) name8174 (
		_w1565_,
		_w9523_,
		_w9524_
	);
	LUT4 #(
		.INIT('h0007)
	) name8175 (
		_w1554_,
		_w9519_,
		_w9524_,
		_w9517_,
		_w9525_
	);
	LUT2 #(
		.INIT('h4)
	) name8176 (
		_w9514_,
		_w9525_,
		_w9526_
	);
	LUT4 #(
		.INIT('hecee)
	) name8177 (
		_w1678_,
		_w9512_,
		_w9513_,
		_w9526_,
		_w9527_
	);
	LUT3 #(
		.INIT('h70)
	) name8178 (
		_w2054_,
		_w2059_,
		_w2116_,
		_w9528_
	);
	LUT4 #(
		.INIT('haaa2)
	) name8179 (
		_w1945_,
		_w2047_,
		_w2105_,
		_w9528_,
		_w9529_
	);
	LUT3 #(
		.INIT('ha2)
	) name8180 (
		\P3_uWord_reg[12]/NET0131 ,
		_w8341_,
		_w9529_,
		_w9530_
	);
	LUT3 #(
		.INIT('h02)
	) name8181 (
		\buf2_reg[12]/NET0131 ,
		_w2105_,
		_w2116_,
		_w9531_
	);
	LUT3 #(
		.INIT('h40)
	) name8182 (
		_w2060_,
		_w2047_,
		_w9531_,
		_w9532_
	);
	LUT4 #(
		.INIT('h0001)
	) name8183 (
		\P3_EAX_reg[13]/NET0131 ,
		\P3_EAX_reg[14]/NET0131 ,
		\P3_EAX_reg[15]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		_w9533_
	);
	LUT4 #(
		.INIT('h0001)
	) name8184 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[10]/NET0131 ,
		\P3_EAX_reg[11]/NET0131 ,
		\P3_EAX_reg[12]/NET0131 ,
		_w9534_
	);
	LUT4 #(
		.INIT('h0001)
	) name8185 (
		\P3_EAX_reg[6]/NET0131 ,
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		\P3_EAX_reg[9]/NET0131 ,
		_w9535_
	);
	LUT4 #(
		.INIT('h0001)
	) name8186 (
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		_w9536_
	);
	LUT4 #(
		.INIT('h8000)
	) name8187 (
		_w9535_,
		_w9536_,
		_w9533_,
		_w9534_,
		_w9537_
	);
	LUT4 #(
		.INIT('h0080)
	) name8188 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w8352_,
		_w9537_,
		_w9538_
	);
	LUT4 #(
		.INIT('h8000)
	) name8189 (
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		\P3_EAX_reg[21]/NET0131 ,
		_w9538_,
		_w9539_
	);
	LUT2 #(
		.INIT('h8)
	) name8190 (
		_w8357_,
		_w9539_,
		_w9540_
	);
	LUT4 #(
		.INIT('h8000)
	) name8191 (
		\P3_EAX_reg[24]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		_w8357_,
		_w9539_,
		_w9541_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		_w8362_,
		_w9541_,
		_w9542_
	);
	LUT3 #(
		.INIT('h08)
	) name8193 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w9543_
	);
	LUT3 #(
		.INIT('h80)
	) name8194 (
		\P3_EAX_reg[28]/NET0131 ,
		_w8362_,
		_w9541_,
		_w9544_
	);
	LUT4 #(
		.INIT('h2313)
	) name8195 (
		\P3_EAX_reg[28]/NET0131 ,
		_w9532_,
		_w9543_,
		_w9542_,
		_w9545_
	);
	LUT3 #(
		.INIT('hce)
	) name8196 (
		_w1945_,
		_w9530_,
		_w9545_,
		_w9546_
	);
	LUT4 #(
		.INIT('h7774)
	) name8197 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w1661_,
		_w7746_,
		_w7744_,
		_w9547_
	);
	LUT4 #(
		.INIT('h028a)
	) name8198 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w9548_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8199 (
		_w1659_,
		_w7739_,
		_w7738_,
		_w9548_,
		_w9549_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8200 (
		_w1559_,
		_w1678_,
		_w9547_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h8)
	) name8201 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w2211_,
		_w9551_
	);
	LUT3 #(
		.INIT('h78)
	) name8202 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9552_
	);
	LUT4 #(
		.INIT('h135f)
	) name8203 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w2283_,
		_w2286_,
		_w9552_,
		_w9553_
	);
	LUT4 #(
		.INIT('h001f)
	) name8204 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9554_
	);
	LUT4 #(
		.INIT('he000)
	) name8205 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9555_
	);
	LUT3 #(
		.INIT('h02)
	) name8206 (
		_w1679_,
		_w9554_,
		_w9555_,
		_w9556_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8207 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9557_
	);
	LUT2 #(
		.INIT('h2)
	) name8208 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		_w9557_,
		_w9558_
	);
	LUT4 #(
		.INIT('h0100)
	) name8209 (
		_w9556_,
		_w9558_,
		_w9551_,
		_w9553_,
		_w9559_
	);
	LUT2 #(
		.INIT('hb)
	) name8210 (
		_w9550_,
		_w9559_,
		_w9560_
	);
	LUT4 #(
		.INIT('h808c)
	) name8211 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w1559_,
		_w1661_,
		_w7757_,
		_w9561_
	);
	LUT4 #(
		.INIT('h028a)
	) name8212 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w9562_
	);
	LUT4 #(
		.INIT('h007d)
	) name8213 (
		_w1659_,
		_w4395_,
		_w7751_,
		_w9562_,
		_w9563_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8214 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5722_,
		_w9337_,
		_w9564_
	);
	LUT2 #(
		.INIT('h8)
	) name8215 (
		_w5746_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h2)
	) name8216 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w5747_,
		_w9566_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8217 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w9567_
	);
	LUT3 #(
		.INIT('h80)
	) name8218 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w9567_,
		_w9568_
	);
	LUT3 #(
		.INIT('h01)
	) name8219 (
		_w7763_,
		_w9568_,
		_w9566_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name8220 (
		_w9565_,
		_w9569_,
		_w9570_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8221 (
		_w1678_,
		_w9561_,
		_w9563_,
		_w9570_,
		_w9571_
	);
	LUT3 #(
		.INIT('h08)
	) name8222 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1592_,
		_w1660_,
		_w9572_
	);
	LUT4 #(
		.INIT('h028a)
	) name8223 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1558_,
		_w1559_,
		_w1596_,
		_w9573_
	);
	LUT4 #(
		.INIT('h00d7)
	) name8224 (
		_w1659_,
		_w7133_,
		_w7134_,
		_w9573_,
		_w9574_
	);
	LUT4 #(
		.INIT('h5700)
	) name8225 (
		_w1559_,
		_w7131_,
		_w9572_,
		_w9574_,
		_w9575_
	);
	LUT3 #(
		.INIT('h6c)
	) name8226 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w5723_,
		_w9576_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8227 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w2283_,
		_w5723_,
		_w9577_
	);
	LUT4 #(
		.INIT('h8848)
	) name8228 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w1679_,
		_w5723_,
		_w6857_,
		_w9578_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8229 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w2286_,
		_w5747_,
		_w9579_
	);
	LUT3 #(
		.INIT('h10)
	) name8230 (
		_w9578_,
		_w9577_,
		_w9579_,
		_w9580_
	);
	LUT3 #(
		.INIT('h2f)
	) name8231 (
		_w1678_,
		_w9575_,
		_w9580_,
		_w9581_
	);
	LUT4 #(
		.INIT('h00a8)
	) name8232 (
		_w2180_,
		_w2755_,
		_w7700_,
		_w7702_,
		_w9582_
	);
	LUT2 #(
		.INIT('h2)
	) name8233 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w7422_,
		_w9583_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8234 (
		_w1945_,
		_w7715_,
		_w9582_,
		_w9583_,
		_w9584_
	);
	LUT2 #(
		.INIT('h8)
	) name8235 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w2225_,
		_w9585_
	);
	LUT3 #(
		.INIT('h78)
	) name8236 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9586_
	);
	LUT4 #(
		.INIT('h0777)
	) name8237 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w3054_,
		_w3055_,
		_w9586_,
		_w9587_
	);
	LUT4 #(
		.INIT('h001f)
	) name8238 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9588_
	);
	LUT4 #(
		.INIT('he000)
	) name8239 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9589_
	);
	LUT3 #(
		.INIT('h02)
	) name8240 (
		_w2194_,
		_w9588_,
		_w9589_,
		_w9590_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8241 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9591_
	);
	LUT2 #(
		.INIT('h2)
	) name8242 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		_w9591_,
		_w9592_
	);
	LUT4 #(
		.INIT('h0100)
	) name8243 (
		_w9590_,
		_w9592_,
		_w9585_,
		_w9587_,
		_w9593_
	);
	LUT2 #(
		.INIT('hb)
	) name8244 (
		_w9584_,
		_w9593_,
		_w9594_
	);
	LUT3 #(
		.INIT('h01)
	) name8245 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2103_,
		_w2172_,
		_w9595_
	);
	LUT3 #(
		.INIT('h04)
	) name8246 (
		_w2060_,
		_w2041_,
		_w9595_,
		_w9596_
	);
	LUT3 #(
		.INIT('hb0)
	) name8247 (
		_w2173_,
		_w7722_,
		_w9596_,
		_w9597_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8248 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w9598_
	);
	LUT4 #(
		.INIT('h000b)
	) name8249 (
		_w7727_,
		_w7730_,
		_w9598_,
		_w9597_,
		_w9599_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8250 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w5757_,
		_w9361_,
		_w9600_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8251 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w9601_
	);
	LUT3 #(
		.INIT('hc4)
	) name8252 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w9601_,
		_w9602_
	);
	LUT3 #(
		.INIT('he0)
	) name8253 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9600_,
		_w9602_,
		_w9603_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8254 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w3054_,
		_w5783_,
		_w9604_
	);
	LUT3 #(
		.INIT('h70)
	) name8255 (
		_w3055_,
		_w9600_,
		_w9604_,
		_w9605_
	);
	LUT2 #(
		.INIT('h4)
	) name8256 (
		_w9603_,
		_w9605_,
		_w9606_
	);
	LUT3 #(
		.INIT('h2f)
	) name8257 (
		_w1945_,
		_w9599_,
		_w9606_,
		_w9607_
	);
	LUT4 #(
		.INIT('h4510)
	) name8258 (
		_w2173_,
		_w4047_,
		_w4048_,
		_w7096_,
		_w9608_
	);
	LUT3 #(
		.INIT('h01)
	) name8259 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2103_,
		_w2172_,
		_w9609_
	);
	LUT3 #(
		.INIT('h04)
	) name8260 (
		_w2060_,
		_w2041_,
		_w9609_,
		_w9610_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8261 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w9611_
	);
	LUT4 #(
		.INIT('h1011)
	) name8262 (
		_w7105_,
		_w9611_,
		_w9608_,
		_w9610_,
		_w9612_
	);
	LUT3 #(
		.INIT('h6c)
	) name8263 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5758_,
		_w9613_
	);
	LUT4 #(
		.INIT('h4105)
	) name8264 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5758_,
		_w9614_
	);
	LUT4 #(
		.INIT('h70d0)
	) name8265 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2194_,
		_w5758_,
		_w9615_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8266 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w3055_,
		_w5758_,
		_w9616_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8267 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w3054_,
		_w5783_,
		_w9617_
	);
	LUT4 #(
		.INIT('h4500)
	) name8268 (
		_w9616_,
		_w9614_,
		_w9615_,
		_w9617_,
		_w9618_
	);
	LUT3 #(
		.INIT('h2f)
	) name8269 (
		_w1945_,
		_w9612_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h2)
	) name8270 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w7547_,
		_w9620_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8271 (
		_w1933_,
		_w7670_,
		_w7675_,
		_w9620_,
		_w9621_
	);
	LUT2 #(
		.INIT('h8)
	) name8272 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w2234_,
		_w9622_
	);
	LUT3 #(
		.INIT('h78)
	) name8273 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9623_
	);
	LUT4 #(
		.INIT('h0777)
	) name8274 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w3406_,
		_w3407_,
		_w9623_,
		_w9624_
	);
	LUT4 #(
		.INIT('h001f)
	) name8275 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9625_
	);
	LUT4 #(
		.INIT('he000)
	) name8276 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9626_
	);
	LUT3 #(
		.INIT('h02)
	) name8277 (
		_w1939_,
		_w9625_,
		_w9626_,
		_w9627_
	);
	LUT4 #(
		.INIT('hfe35)
	) name8278 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9628_
	);
	LUT2 #(
		.INIT('h2)
	) name8279 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w9628_,
		_w9629_
	);
	LUT4 #(
		.INIT('h0100)
	) name8280 (
		_w9627_,
		_w9629_,
		_w9622_,
		_w9624_,
		_w9630_
	);
	LUT2 #(
		.INIT('hb)
	) name8281 (
		_w9621_,
		_w9630_,
		_w9631_
	);
	LUT4 #(
		.INIT('h4774)
	) name8282 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1916_,
		_w3285_,
		_w7684_,
		_w9632_
	);
	LUT2 #(
		.INIT('h2)
	) name8283 (
		_w1810_,
		_w9632_,
		_w9633_
	);
	LUT4 #(
		.INIT('h028a)
	) name8284 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w9634_
	);
	LUT3 #(
		.INIT('h0b)
	) name8285 (
		_w7690_,
		_w7693_,
		_w9634_,
		_w9635_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name8286 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w6364_,
		_w9374_,
		_w9636_
	);
	LUT2 #(
		.INIT('h8)
	) name8287 (
		_w6378_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h2)
	) name8288 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w6383_,
		_w9638_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8289 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w9639_
	);
	LUT3 #(
		.INIT('h80)
	) name8290 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w9639_,
		_w9640_
	);
	LUT3 #(
		.INIT('h01)
	) name8291 (
		_w7696_,
		_w9640_,
		_w9638_,
		_w9641_
	);
	LUT2 #(
		.INIT('h4)
	) name8292 (
		_w9637_,
		_w9641_,
		_w9642_
	);
	LUT4 #(
		.INIT('h8aff)
	) name8293 (
		_w1933_,
		_w9633_,
		_w9635_,
		_w9642_,
		_w9643_
	);
	LUT4 #(
		.INIT('h5070)
	) name8294 (
		_w1810_,
		_w1916_,
		_w6357_,
		_w7085_,
		_w9644_
	);
	LUT4 #(
		.INIT('h00df)
	) name8295 (
		_w1810_,
		_w1916_,
		_w7085_,
		_w7089_,
		_w9645_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8296 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1933_,
		_w9644_,
		_w9645_,
		_w9646_
	);
	LUT3 #(
		.INIT('h6c)
	) name8297 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w6365_,
		_w9647_
	);
	LUT4 #(
		.INIT('h4105)
	) name8298 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w6365_,
		_w9648_
	);
	LUT4 #(
		.INIT('h70d0)
	) name8299 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w1939_,
		_w6365_,
		_w9649_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8300 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w3407_,
		_w6365_,
		_w9650_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8301 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w3406_,
		_w6383_,
		_w9651_
	);
	LUT4 #(
		.INIT('h4500)
	) name8302 (
		_w9650_,
		_w9648_,
		_w9649_,
		_w9651_,
		_w9652_
	);
	LUT2 #(
		.INIT('hb)
	) name8303 (
		_w9646_,
		_w9652_,
		_w9653_
	);
	LUT2 #(
		.INIT('h2)
	) name8304 (
		\P1_EAX_reg[29]/NET0131 ,
		_w9102_,
		_w9654_
	);
	LUT4 #(
		.INIT('h8000)
	) name8305 (
		_w9430_,
		_w9432_,
		_w9433_,
		_w9477_,
		_w9655_
	);
	LUT3 #(
		.INIT('h80)
	) name8306 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w9655_,
		_w9656_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8307 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w1827_,
		_w9655_,
		_w9657_
	);
	LUT4 #(
		.INIT('h8008)
	) name8308 (
		_w1832_,
		_w1846_,
		_w9073_,
		_w9084_,
		_w9658_
	);
	LUT4 #(
		.INIT('h0080)
	) name8309 (
		_w1725_,
		_w1802_,
		_w1867_,
		_w4502_,
		_w9659_
	);
	LUT3 #(
		.INIT('h08)
	) name8310 (
		_w1795_,
		_w1867_,
		_w3467_,
		_w9660_
	);
	LUT2 #(
		.INIT('h1)
	) name8311 (
		_w9659_,
		_w9660_,
		_w9661_
	);
	LUT4 #(
		.INIT('h7500)
	) name8312 (
		\P1_EAX_reg[29]/NET0131 ,
		_w9436_,
		_w9437_,
		_w9661_,
		_w9662_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8313 (
		_w1933_,
		_w9658_,
		_w9657_,
		_w9662_,
		_w9663_
	);
	LUT2 #(
		.INIT('he)
	) name8314 (
		_w9654_,
		_w9663_,
		_w9664_
	);
	LUT2 #(
		.INIT('h2)
	) name8315 (
		\P3_EAX_reg[29]/NET0131 ,
		_w8341_,
		_w9665_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8316 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w8361_,
		_w8363_,
		_w9666_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8317 (
		\P3_EAX_reg[29]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w9667_
	);
	LUT4 #(
		.INIT('h02fd)
	) name8318 (
		_w8426_,
		_w8437_,
		_w8867_,
		_w8878_,
		_w9668_
	);
	LUT2 #(
		.INIT('h8)
	) name8319 (
		_w8366_,
		_w9668_,
		_w9669_
	);
	LUT3 #(
		.INIT('h80)
	) name8320 (
		\buf2_reg[29]/NET0131 ,
		_w2060_,
		_w2044_,
		_w9670_
	);
	LUT3 #(
		.INIT('h20)
	) name8321 (
		\buf2_reg[13]/NET0131 ,
		_w2060_,
		_w2047_,
		_w9671_
	);
	LUT3 #(
		.INIT('ha8)
	) name8322 (
		_w2119_,
		_w9670_,
		_w9671_,
		_w9672_
	);
	LUT2 #(
		.INIT('h1)
	) name8323 (
		_w9669_,
		_w9672_,
		_w9673_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name8324 (
		_w1945_,
		_w9666_,
		_w9667_,
		_w9673_,
		_w9674_
	);
	LUT2 #(
		.INIT('he)
	) name8325 (
		_w9665_,
		_w9674_,
		_w9675_
	);
	LUT2 #(
		.INIT('h4)
	) name8326 (
		_w7777_,
		_w7789_,
		_w9676_
	);
	LUT3 #(
		.INIT('h60)
	) name8327 (
		\P2_EAX_reg[15]/NET0131 ,
		_w7776_,
		_w7789_,
		_w9677_
	);
	LUT4 #(
		.INIT('h153f)
	) name8328 (
		\P2_InstQueue_reg[10][7]/NET0131 ,
		\P2_InstQueue_reg[3][7]/NET0131 ,
		_w1462_,
		_w1465_,
		_w9678_
	);
	LUT4 #(
		.INIT('h153f)
	) name8329 (
		\P2_InstQueue_reg[14][7]/NET0131 ,
		\P2_InstQueue_reg[1][7]/NET0131 ,
		_w1453_,
		_w1447_,
		_w9679_
	);
	LUT4 #(
		.INIT('h153f)
	) name8330 (
		\P2_InstQueue_reg[2][7]/NET0131 ,
		\P2_InstQueue_reg[5][7]/NET0131 ,
		_w1450_,
		_w1446_,
		_w9680_
	);
	LUT4 #(
		.INIT('h135f)
	) name8331 (
		\P2_InstQueue_reg[12][7]/NET0131 ,
		\P2_InstQueue_reg[6][7]/NET0131 ,
		_w1443_,
		_w1466_,
		_w9681_
	);
	LUT4 #(
		.INIT('h8000)
	) name8332 (
		_w9680_,
		_w9681_,
		_w9678_,
		_w9679_,
		_w9682_
	);
	LUT4 #(
		.INIT('h153f)
	) name8333 (
		\P2_InstQueue_reg[15][7]/NET0131 ,
		\P2_InstQueue_reg[4][7]/NET0131 ,
		_w1463_,
		_w1460_,
		_w9683_
	);
	LUT4 #(
		.INIT('h135f)
	) name8334 (
		\P2_InstQueue_reg[11][7]/NET0131 ,
		\P2_InstQueue_reg[8][7]/NET0131 ,
		_w1452_,
		_w1456_,
		_w9684_
	);
	LUT4 #(
		.INIT('h153f)
	) name8335 (
		\P2_InstQueue_reg[0][7]/NET0131 ,
		\P2_InstQueue_reg[7][7]/NET0131 ,
		_w1449_,
		_w1457_,
		_w9685_
	);
	LUT4 #(
		.INIT('h153f)
	) name8336 (
		\P2_InstQueue_reg[13][7]/NET0131 ,
		\P2_InstQueue_reg[9][7]/NET0131 ,
		_w1444_,
		_w1459_,
		_w9686_
	);
	LUT4 #(
		.INIT('h8000)
	) name8337 (
		_w9685_,
		_w9686_,
		_w9683_,
		_w9684_,
		_w9687_
	);
	LUT4 #(
		.INIT('h0111)
	) name8338 (
		_w1592_,
		_w1595_,
		_w9682_,
		_w9687_,
		_w9688_
	);
	LUT3 #(
		.INIT('h80)
	) name8339 (
		_w1549_,
		_w1553_,
		_w9688_,
		_w9689_
	);
	LUT4 #(
		.INIT('h0222)
	) name8340 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[15]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9690_
	);
	LUT4 #(
		.INIT('h3111)
	) name8341 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[15]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9691_
	);
	LUT3 #(
		.INIT('h01)
	) name8342 (
		_w1605_,
		_w9691_,
		_w9690_,
		_w9692_
	);
	LUT3 #(
		.INIT('h13)
	) name8343 (
		_w1656_,
		_w9689_,
		_w9692_,
		_w9693_
	);
	LUT4 #(
		.INIT('h0d00)
	) name8344 (
		\P2_EAX_reg[15]/NET0131 ,
		_w7792_,
		_w9677_,
		_w9693_,
		_w9694_
	);
	LUT2 #(
		.INIT('h2)
	) name8345 (
		\P2_EAX_reg[15]/NET0131 ,
		_w7767_,
		_w9695_
	);
	LUT3 #(
		.INIT('hf2)
	) name8346 (
		_w1678_,
		_w9694_,
		_w9695_,
		_w9696_
	);
	LUT2 #(
		.INIT('h2)
	) name8347 (
		\P2_EAX_reg[29]/NET0131 ,
		_w7767_,
		_w9697_
	);
	LUT4 #(
		.INIT('h6a00)
	) name8348 (
		\P2_EAX_reg[29]/NET0131 ,
		_w7784_,
		_w7786_,
		_w7789_,
		_w9698_
	);
	LUT4 #(
		.INIT('h8008)
	) name8349 (
		_w1554_,
		_w1596_,
		_w7873_,
		_w7884_,
		_w9699_
	);
	LUT4 #(
		.INIT('hc444)
	) name8350 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[13]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9700_
	);
	LUT4 #(
		.INIT('h0888)
	) name8351 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[13]/NET0131 ,
		_w2255_,
		_w2260_,
		_w9701_
	);
	LUT2 #(
		.INIT('h1)
	) name8352 (
		_w9700_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h2)
	) name8353 (
		_w1565_,
		_w9702_,
		_w9703_
	);
	LUT3 #(
		.INIT('h08)
	) name8354 (
		_w1501_,
		_w1568_,
		_w6493_,
		_w9704_
	);
	LUT3 #(
		.INIT('ha8)
	) name8355 (
		_w1606_,
		_w9703_,
		_w9704_,
		_w9705_
	);
	LUT4 #(
		.INIT('h000d)
	) name8356 (
		\P2_EAX_reg[29]/NET0131 ,
		_w7792_,
		_w9699_,
		_w9705_,
		_w9706_
	);
	LUT4 #(
		.INIT('hecee)
	) name8357 (
		_w1678_,
		_w9697_,
		_w9698_,
		_w9706_,
		_w9707_
	);
	LUT4 #(
		.INIT('h60c0)
	) name8358 (
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w1829_,
		_w8987_,
		_w9708_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name8359 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1846_,
		_w9038_,
		_w9049_,
		_w9709_
	);
	LUT4 #(
		.INIT('hfd31)
	) name8360 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1814_,
		_w1829_,
		_w9709_,
		_w9710_
	);
	LUT2 #(
		.INIT('h2)
	) name8361 (
		\P1_EBX_reg[26]/NET0131 ,
		_w9102_,
		_w9711_
	);
	LUT4 #(
		.INIT('hff8a)
	) name8362 (
		_w1933_,
		_w9708_,
		_w9710_,
		_w9711_,
		_w9712_
	);
	LUT4 #(
		.INIT('h4888)
	) name8363 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1578_,
		_w8957_,
		_w8958_,
		_w9713_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name8364 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1596_,
		_w7838_,
		_w7849_,
		_w9714_
	);
	LUT4 #(
		.INIT('h002a)
	) name8365 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1503_,
		_w1549_,
		_w1578_,
		_w9715_
	);
	LUT3 #(
		.INIT('h0d)
	) name8366 (
		_w1550_,
		_w9714_,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h2)
	) name8367 (
		\P2_EBX_reg[26]/NET0131 ,
		_w7767_,
		_w9717_
	);
	LUT4 #(
		.INIT('hff8a)
	) name8368 (
		_w1678_,
		_w9713_,
		_w9716_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h2)
	) name8369 (
		\P1_EAX_reg[15]/NET0131 ,
		_w9102_,
		_w9719_
	);
	LUT3 #(
		.INIT('h08)
	) name8370 (
		_w1804_,
		_w1826_,
		_w9425_,
		_w9720_
	);
	LUT4 #(
		.INIT('haa8a)
	) name8371 (
		\P1_EAX_reg[15]/NET0131 ,
		_w9436_,
		_w9437_,
		_w9720_,
		_w9721_
	);
	LUT2 #(
		.INIT('h2)
	) name8372 (
		\P1_EAX_reg[14]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		_w9722_
	);
	LUT4 #(
		.INIT('h8000)
	) name8373 (
		_w1804_,
		_w1826_,
		_w9424_,
		_w9722_,
		_w9723_
	);
	LUT4 #(
		.INIT('h135f)
	) name8374 (
		\P1_InstQueue_reg[2][7]/NET0131 ,
		\P1_InstQueue_reg[6][7]/NET0131 ,
		_w1688_,
		_w1689_,
		_w9724_
	);
	LUT4 #(
		.INIT('h153f)
	) name8375 (
		\P1_InstQueue_reg[15][7]/NET0131 ,
		\P1_InstQueue_reg[9][7]/NET0131 ,
		_w1708_,
		_w1705_,
		_w9725_
	);
	LUT4 #(
		.INIT('h153f)
	) name8376 (
		\P1_InstQueue_reg[1][7]/NET0131 ,
		\P1_InstQueue_reg[3][7]/NET0131 ,
		_w1692_,
		_w1706_,
		_w9726_
	);
	LUT4 #(
		.INIT('h135f)
	) name8377 (
		\P1_InstQueue_reg[13][7]/NET0131 ,
		\P1_InstQueue_reg[4][7]/NET0131 ,
		_w1696_,
		_w1709_,
		_w9727_
	);
	LUT4 #(
		.INIT('h8000)
	) name8378 (
		_w9726_,
		_w9727_,
		_w9724_,
		_w9725_,
		_w9728_
	);
	LUT4 #(
		.INIT('h153f)
	) name8379 (
		\P1_InstQueue_reg[11][7]/NET0131 ,
		\P1_InstQueue_reg[7][7]/NET0131 ,
		_w1691_,
		_w1703_,
		_w9729_
	);
	LUT4 #(
		.INIT('h135f)
	) name8380 (
		\P1_InstQueue_reg[10][7]/NET0131 ,
		\P1_InstQueue_reg[5][7]/NET0131 ,
		_w1712_,
		_w1702_,
		_w9730_
	);
	LUT4 #(
		.INIT('h135f)
	) name8381 (
		\P1_InstQueue_reg[14][7]/NET0131 ,
		\P1_InstQueue_reg[8][7]/NET0131 ,
		_w1698_,
		_w1711_,
		_w9731_
	);
	LUT4 #(
		.INIT('h153f)
	) name8382 (
		\P1_InstQueue_reg[0][7]/NET0131 ,
		\P1_InstQueue_reg[12][7]/NET0131 ,
		_w1694_,
		_w1699_,
		_w9732_
	);
	LUT4 #(
		.INIT('h8000)
	) name8383 (
		_w9731_,
		_w9732_,
		_w9729_,
		_w9730_,
		_w9733_
	);
	LUT4 #(
		.INIT('h0111)
	) name8384 (
		_w1842_,
		_w1845_,
		_w9728_,
		_w9733_,
		_w9734_
	);
	LUT4 #(
		.INIT('h4000)
	) name8385 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w9734_,
		_w9735_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8386 (
		_w1855_,
		_w1861_,
		_w3460_,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h4)
	) name8387 (
		_w9723_,
		_w9736_,
		_w9737_
	);
	LUT4 #(
		.INIT('hecee)
	) name8388 (
		_w1933_,
		_w9719_,
		_w9721_,
		_w9737_,
		_w9738_
	);
	LUT3 #(
		.INIT('h28)
	) name8389 (
		_w3411_,
		_w3513_,
		_w3516_,
		_w9739_
	);
	LUT4 #(
		.INIT('h2ad5)
	) name8390 (
		_w3425_,
		_w3454_,
		_w3483_,
		_w3500_,
		_w9740_
	);
	LUT3 #(
		.INIT('hc8)
	) name8391 (
		_w3411_,
		_w4956_,
		_w9740_,
		_w9741_
	);
	LUT3 #(
		.INIT('h02)
	) name8392 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w3534_,
		_w3536_,
		_w9742_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8393 (
		_w3537_,
		_w3469_,
		_w3470_,
		_w9742_,
		_w9743_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8394 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3413_,
		_w4953_,
		_w9744_
	);
	LUT2 #(
		.INIT('h4)
	) name8395 (
		_w9743_,
		_w9744_,
		_w9745_
	);
	LUT2 #(
		.INIT('h2)
	) name8396 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w3545_,
		_w9746_
	);
	LUT4 #(
		.INIT('hc055)
	) name8397 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3534_,
		_w9747_
	);
	LUT3 #(
		.INIT('h31)
	) name8398 (
		_w2248_,
		_w9746_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h4)
	) name8399 (
		_w9745_,
		_w9748_,
		_w9749_
	);
	LUT3 #(
		.INIT('h4f)
	) name8400 (
		_w9739_,
		_w9741_,
		_w9749_,
		_w9750_
	);
	LUT3 #(
		.INIT('h01)
	) name8401 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1605_,
		_w1611_,
		_w9751_
	);
	LUT3 #(
		.INIT('h02)
	) name8402 (
		_w1566_,
		_w1602_,
		_w9751_,
		_w9752_
	);
	LUT4 #(
		.INIT('h0001)
	) name8403 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w9753_
	);
	LUT4 #(
		.INIT('h0100)
	) name8404 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w9753_,
		_w9754_
	);
	LUT4 #(
		.INIT('h0100)
	) name8405 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w9754_,
		_w9755_
	);
	LUT4 #(
		.INIT('h0100)
	) name8406 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[12]/NET0131 ,
		_w9755_,
		_w9756_
	);
	LUT4 #(
		.INIT('h0001)
	) name8407 (
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[15]/NET0131 ,
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[17]/NET0131 ,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name8408 (
		\P2_EBX_reg[18]/NET0131 ,
		\P2_EBX_reg[19]/NET0131 ,
		_w9758_
	);
	LUT4 #(
		.INIT('h4000)
	) name8409 (
		\P2_EBX_reg[13]/NET0131 ,
		_w9756_,
		_w9757_,
		_w9758_,
		_w9759_
	);
	LUT2 #(
		.INIT('h1)
	) name8410 (
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w9760_
	);
	LUT4 #(
		.INIT('h1000)
	) name8411 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		_w9759_,
		_w9760_,
		_w9761_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		_w9762_
	);
	LUT2 #(
		.INIT('h1)
	) name8413 (
		\P2_EBX_reg[27]/NET0131 ,
		\P2_EBX_reg[28]/NET0131 ,
		_w9763_
	);
	LUT4 #(
		.INIT('h4000)
	) name8414 (
		\P2_EBX_reg[26]/NET0131 ,
		_w9761_,
		_w9762_,
		_w9763_,
		_w9764_
	);
	LUT3 #(
		.INIT('h02)
	) name8415 (
		_w1565_,
		_w1602_,
		_w1673_,
		_w9765_
	);
	LUT4 #(
		.INIT('h0004)
	) name8416 (
		\P2_EBX_reg[30]/NET0131 ,
		_w1565_,
		_w1602_,
		_w1673_,
		_w9766_
	);
	LUT4 #(
		.INIT('h2333)
	) name8417 (
		\P2_EBX_reg[29]/NET0131 ,
		_w9752_,
		_w9764_,
		_w9766_,
		_w9767_
	);
	LUT4 #(
		.INIT('h8000)
	) name8418 (
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w9768_
	);
	LUT3 #(
		.INIT('h80)
	) name8419 (
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w9769_
	);
	LUT4 #(
		.INIT('h8000)
	) name8420 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9768_,
		_w9769_,
		_w9770_
	);
	LUT2 #(
		.INIT('h8)
	) name8421 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w9771_
	);
	LUT3 #(
		.INIT('h80)
	) name8422 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9772_
	);
	LUT2 #(
		.INIT('h8)
	) name8423 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w9773_
	);
	LUT3 #(
		.INIT('h80)
	) name8424 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w9774_
	);
	LUT4 #(
		.INIT('h8000)
	) name8425 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w9775_
	);
	LUT2 #(
		.INIT('h8)
	) name8426 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9775_,
		_w9776_
	);
	LUT3 #(
		.INIT('h80)
	) name8427 (
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w9775_,
		_w9777_
	);
	LUT4 #(
		.INIT('h8000)
	) name8428 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9777_,
		_w9778_
	);
	LUT3 #(
		.INIT('h80)
	) name8429 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w9778_,
		_w9779_
	);
	LUT4 #(
		.INIT('h8000)
	) name8430 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w9778_,
		_w9780_
	);
	LUT3 #(
		.INIT('h80)
	) name8431 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w9780_,
		_w9781_
	);
	LUT4 #(
		.INIT('h8000)
	) name8432 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9780_,
		_w9782_
	);
	LUT3 #(
		.INIT('h80)
	) name8433 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9782_,
		_w9783_
	);
	LUT4 #(
		.INIT('h8000)
	) name8434 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w9782_,
		_w9784_
	);
	LUT3 #(
		.INIT('h80)
	) name8435 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9784_,
		_w9785_
	);
	LUT4 #(
		.INIT('hf5f1)
	) name8436 (
		_w1565_,
		_w1566_,
		_w1602_,
		_w1611_,
		_w9786_
	);
	LUT2 #(
		.INIT('h2)
	) name8437 (
		_w1673_,
		_w9786_,
		_w9787_
	);
	LUT4 #(
		.INIT('h00fe)
	) name8438 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1602_,
		_w9788_
	);
	LUT4 #(
		.INIT('h9f15)
	) name8439 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w9785_,
		_w9787_,
		_w9788_,
		_w9789_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8440 (
		\P2_EBX_reg[31]/NET0131 ,
		_w1678_,
		_w9767_,
		_w9789_,
		_w9790_
	);
	LUT2 #(
		.INIT('h8)
	) name8441 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w9791_
	);
	LUT2 #(
		.INIT('h4)
	) name8442 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w9792_
	);
	LUT2 #(
		.INIT('h8)
	) name8443 (
		_w8260_,
		_w9792_,
		_w9793_
	);
	LUT3 #(
		.INIT('h80)
	) name8444 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		_w5736_,
		_w9793_,
		_w9794_
	);
	LUT4 #(
		.INIT('h8000)
	) name8445 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		_w5736_,
		_w9793_,
		_w9795_
	);
	LUT2 #(
		.INIT('h8)
	) name8446 (
		_w5741_,
		_w9795_,
		_w9796_
	);
	LUT3 #(
		.INIT('h40)
	) name8447 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w5741_,
		_w9795_,
		_w9797_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name8448 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9791_,
		_w9797_,
		_w9798_
	);
	LUT4 #(
		.INIT('hfe25)
	) name8449 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9799_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8450 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2211_,
		_w9799_,
		_w9800_
	);
	LUT3 #(
		.INIT('hd0)
	) name8451 (
		_w1679_,
		_w9798_,
		_w9800_,
		_w9801_
	);
	LUT2 #(
		.INIT('hb)
	) name8452 (
		_w9790_,
		_w9801_,
		_w9802_
	);
	LUT3 #(
		.INIT('h60)
	) name8453 (
		_w3513_,
		_w3516_,
		_w3572_,
		_w9803_
	);
	LUT3 #(
		.INIT('hc8)
	) name8454 (
		_w3572_,
		_w4990_,
		_w9740_,
		_w9804_
	);
	LUT3 #(
		.INIT('h02)
	) name8455 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w3578_,
		_w3580_,
		_w9805_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8456 (
		_w3469_,
		_w3470_,
		_w3581_,
		_w9805_,
		_w9806_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8457 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3574_,
		_w4953_,
		_w9807_
	);
	LUT2 #(
		.INIT('h4)
	) name8458 (
		_w9806_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h2)
	) name8459 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w3545_,
		_w9809_
	);
	LUT4 #(
		.INIT('hc055)
	) name8460 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3578_,
		_w9810_
	);
	LUT3 #(
		.INIT('h31)
	) name8461 (
		_w2248_,
		_w9809_,
		_w9810_,
		_w9811_
	);
	LUT2 #(
		.INIT('h4)
	) name8462 (
		_w9808_,
		_w9811_,
		_w9812_
	);
	LUT3 #(
		.INIT('h4f)
	) name8463 (
		_w9803_,
		_w9804_,
		_w9812_,
		_w9813_
	);
	LUT3 #(
		.INIT('h60)
	) name8464 (
		_w3513_,
		_w3516_,
		_w3592_,
		_w9814_
	);
	LUT3 #(
		.INIT('hc8)
	) name8465 (
		_w3592_,
		_w5001_,
		_w9740_,
		_w9815_
	);
	LUT3 #(
		.INIT('h02)
	) name8466 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		_w3536_,
		_w3412_,
		_w9816_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8467 (
		_w3469_,
		_w3470_,
		_w3597_,
		_w9816_,
		_w9817_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8468 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3593_,
		_w4953_,
		_w9818_
	);
	LUT2 #(
		.INIT('h4)
	) name8469 (
		_w9817_,
		_w9818_,
		_w9819_
	);
	LUT2 #(
		.INIT('h2)
	) name8470 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		_w3545_,
		_w9820_
	);
	LUT4 #(
		.INIT('hc055)
	) name8471 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3536_,
		_w9821_
	);
	LUT3 #(
		.INIT('h31)
	) name8472 (
		_w2248_,
		_w9820_,
		_w9821_,
		_w9822_
	);
	LUT2 #(
		.INIT('h4)
	) name8473 (
		_w9819_,
		_w9822_,
		_w9823_
	);
	LUT3 #(
		.INIT('h4f)
	) name8474 (
		_w9814_,
		_w9815_,
		_w9823_,
		_w9824_
	);
	LUT3 #(
		.INIT('h28)
	) name8475 (
		_w3412_,
		_w3513_,
		_w3516_,
		_w9825_
	);
	LUT3 #(
		.INIT('hc8)
	) name8476 (
		_w3412_,
		_w5012_,
		_w9740_,
		_w9826_
	);
	LUT3 #(
		.INIT('h02)
	) name8477 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w3534_,
		_w3611_,
		_w9827_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8478 (
		_w3469_,
		_w3470_,
		_w3612_,
		_w9827_,
		_w9828_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8479 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3597_,
		_w4953_,
		_w9829_
	);
	LUT2 #(
		.INIT('h4)
	) name8480 (
		_w9828_,
		_w9829_,
		_w9830_
	);
	LUT2 #(
		.INIT('h2)
	) name8481 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w3545_,
		_w9831_
	);
	LUT4 #(
		.INIT('hc055)
	) name8482 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3611_,
		_w9832_
	);
	LUT3 #(
		.INIT('h31)
	) name8483 (
		_w2248_,
		_w9831_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h4)
	) name8484 (
		_w9830_,
		_w9833_,
		_w9834_
	);
	LUT3 #(
		.INIT('h4f)
	) name8485 (
		_w9825_,
		_w9826_,
		_w9834_,
		_w9835_
	);
	LUT3 #(
		.INIT('h28)
	) name8486 (
		_w3536_,
		_w3513_,
		_w3516_,
		_w9836_
	);
	LUT3 #(
		.INIT('hc8)
	) name8487 (
		_w3536_,
		_w5023_,
		_w9740_,
		_w9837_
	);
	LUT3 #(
		.INIT('h02)
	) name8488 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w3572_,
		_w3611_,
		_w9838_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8489 (
		_w3469_,
		_w3470_,
		_w3626_,
		_w9838_,
		_w9839_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8490 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3537_,
		_w4953_,
		_w9840_
	);
	LUT2 #(
		.INIT('h4)
	) name8491 (
		_w9839_,
		_w9840_,
		_w9841_
	);
	LUT2 #(
		.INIT('h2)
	) name8492 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w3545_,
		_w9842_
	);
	LUT4 #(
		.INIT('hc055)
	) name8493 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3572_,
		_w9843_
	);
	LUT3 #(
		.INIT('h31)
	) name8494 (
		_w2248_,
		_w9842_,
		_w9843_,
		_w9844_
	);
	LUT2 #(
		.INIT('h4)
	) name8495 (
		_w9841_,
		_w9844_,
		_w9845_
	);
	LUT3 #(
		.INIT('h4f)
	) name8496 (
		_w9836_,
		_w9837_,
		_w9845_,
		_w9846_
	);
	LUT3 #(
		.INIT('h28)
	) name8497 (
		_w3534_,
		_w3513_,
		_w3516_,
		_w9847_
	);
	LUT3 #(
		.INIT('hc8)
	) name8498 (
		_w3534_,
		_w5034_,
		_w9740_,
		_w9848_
	);
	LUT3 #(
		.INIT('h02)
	) name8499 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w3572_,
		_w3573_,
		_w9849_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8500 (
		_w3469_,
		_w3470_,
		_w3574_,
		_w9849_,
		_w9850_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8501 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3612_,
		_w4953_,
		_w9851_
	);
	LUT2 #(
		.INIT('h4)
	) name8502 (
		_w9850_,
		_w9851_,
		_w9852_
	);
	LUT2 #(
		.INIT('h2)
	) name8503 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w3545_,
		_w9853_
	);
	LUT4 #(
		.INIT('hc055)
	) name8504 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3573_,
		_w9854_
	);
	LUT3 #(
		.INIT('h31)
	) name8505 (
		_w2248_,
		_w9853_,
		_w9854_,
		_w9855_
	);
	LUT2 #(
		.INIT('h4)
	) name8506 (
		_w9852_,
		_w9855_,
		_w9856_
	);
	LUT3 #(
		.INIT('h4f)
	) name8507 (
		_w9847_,
		_w9848_,
		_w9856_,
		_w9857_
	);
	LUT3 #(
		.INIT('h60)
	) name8508 (
		_w3513_,
		_w3516_,
		_w3611_,
		_w9858_
	);
	LUT3 #(
		.INIT('hc8)
	) name8509 (
		_w3611_,
		_w5045_,
		_w9740_,
		_w9859_
	);
	LUT3 #(
		.INIT('h02)
	) name8510 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w3580_,
		_w3573_,
		_w9860_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8511 (
		_w3469_,
		_w3470_,
		_w3653_,
		_w9860_,
		_w9861_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8512 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3626_,
		_w4953_,
		_w9862_
	);
	LUT2 #(
		.INIT('h4)
	) name8513 (
		_w9861_,
		_w9862_,
		_w9863_
	);
	LUT2 #(
		.INIT('h2)
	) name8514 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w3545_,
		_w9864_
	);
	LUT4 #(
		.INIT('hc055)
	) name8515 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3580_,
		_w9865_
	);
	LUT3 #(
		.INIT('h31)
	) name8516 (
		_w2248_,
		_w9864_,
		_w9865_,
		_w9866_
	);
	LUT2 #(
		.INIT('h4)
	) name8517 (
		_w9863_,
		_w9866_,
		_w9867_
	);
	LUT3 #(
		.INIT('h4f)
	) name8518 (
		_w9858_,
		_w9859_,
		_w9867_,
		_w9868_
	);
	LUT3 #(
		.INIT('h60)
	) name8519 (
		_w3513_,
		_w3516_,
		_w3573_,
		_w9869_
	);
	LUT3 #(
		.INIT('hc8)
	) name8520 (
		_w3573_,
		_w5056_,
		_w9740_,
		_w9870_
	);
	LUT3 #(
		.INIT('h02)
	) name8521 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w3578_,
		_w3667_,
		_w9871_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8522 (
		_w3469_,
		_w3470_,
		_w3668_,
		_w9871_,
		_w9872_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8523 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3653_,
		_w4953_,
		_w9873_
	);
	LUT2 #(
		.INIT('h4)
	) name8524 (
		_w9872_,
		_w9873_,
		_w9874_
	);
	LUT2 #(
		.INIT('h2)
	) name8525 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w3545_,
		_w9875_
	);
	LUT4 #(
		.INIT('hc055)
	) name8526 (
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3667_,
		_w9876_
	);
	LUT3 #(
		.INIT('h31)
	) name8527 (
		_w2248_,
		_w9875_,
		_w9876_,
		_w9877_
	);
	LUT2 #(
		.INIT('h4)
	) name8528 (
		_w9874_,
		_w9877_,
		_w9878_
	);
	LUT3 #(
		.INIT('h4f)
	) name8529 (
		_w9869_,
		_w9870_,
		_w9878_,
		_w9879_
	);
	LUT3 #(
		.INIT('h60)
	) name8530 (
		_w3513_,
		_w3516_,
		_w3580_,
		_w9880_
	);
	LUT3 #(
		.INIT('hc8)
	) name8531 (
		_w3580_,
		_w5067_,
		_w9740_,
		_w9881_
	);
	LUT3 #(
		.INIT('h02)
	) name8532 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w3667_,
		_w3683_,
		_w9882_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8533 (
		_w3469_,
		_w3470_,
		_w3698_,
		_w9882_,
		_w9883_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8534 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3581_,
		_w4953_,
		_w9884_
	);
	LUT2 #(
		.INIT('h4)
	) name8535 (
		_w9883_,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h2)
	) name8536 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w3545_,
		_w9886_
	);
	LUT4 #(
		.INIT('hc055)
	) name8537 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3683_,
		_w9887_
	);
	LUT3 #(
		.INIT('h31)
	) name8538 (
		_w2248_,
		_w9886_,
		_w9887_,
		_w9888_
	);
	LUT2 #(
		.INIT('h4)
	) name8539 (
		_w9885_,
		_w9888_,
		_w9889_
	);
	LUT3 #(
		.INIT('h4f)
	) name8540 (
		_w9880_,
		_w9881_,
		_w9889_,
		_w9890_
	);
	LUT3 #(
		.INIT('h60)
	) name8541 (
		_w3513_,
		_w3516_,
		_w3578_,
		_w9891_
	);
	LUT3 #(
		.INIT('hc8)
	) name8542 (
		_w3578_,
		_w5078_,
		_w9740_,
		_w9892_
	);
	LUT3 #(
		.INIT('h02)
	) name8543 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w3682_,
		_w3683_,
		_w9893_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8544 (
		_w3469_,
		_w3470_,
		_w3684_,
		_w9893_,
		_w9894_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8545 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3668_,
		_w4953_,
		_w9895_
	);
	LUT2 #(
		.INIT('h4)
	) name8546 (
		_w9894_,
		_w9895_,
		_w9896_
	);
	LUT2 #(
		.INIT('h2)
	) name8547 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w3545_,
		_w9897_
	);
	LUT4 #(
		.INIT('hc055)
	) name8548 (
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3682_,
		_w9898_
	);
	LUT3 #(
		.INIT('h31)
	) name8549 (
		_w2248_,
		_w9897_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h4)
	) name8550 (
		_w9896_,
		_w9899_,
		_w9900_
	);
	LUT3 #(
		.INIT('h4f)
	) name8551 (
		_w9891_,
		_w9892_,
		_w9900_,
		_w9901_
	);
	LUT3 #(
		.INIT('h60)
	) name8552 (
		_w3513_,
		_w3516_,
		_w3667_,
		_w9902_
	);
	LUT3 #(
		.INIT('hc8)
	) name8553 (
		_w3667_,
		_w5089_,
		_w9740_,
		_w9903_
	);
	LUT3 #(
		.INIT('h02)
	) name8554 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w3682_,
		_w3712_,
		_w9904_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8555 (
		_w3469_,
		_w3470_,
		_w3713_,
		_w9904_,
		_w9905_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8556 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3698_,
		_w4953_,
		_w9906_
	);
	LUT2 #(
		.INIT('h4)
	) name8557 (
		_w9905_,
		_w9906_,
		_w9907_
	);
	LUT2 #(
		.INIT('h2)
	) name8558 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w3545_,
		_w9908_
	);
	LUT4 #(
		.INIT('hc055)
	) name8559 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3712_,
		_w9909_
	);
	LUT3 #(
		.INIT('h31)
	) name8560 (
		_w2248_,
		_w9908_,
		_w9909_,
		_w9910_
	);
	LUT2 #(
		.INIT('h4)
	) name8561 (
		_w9907_,
		_w9910_,
		_w9911_
	);
	LUT3 #(
		.INIT('h4f)
	) name8562 (
		_w9902_,
		_w9903_,
		_w9911_,
		_w9912_
	);
	LUT3 #(
		.INIT('h60)
	) name8563 (
		_w3513_,
		_w3516_,
		_w3683_,
		_w9913_
	);
	LUT3 #(
		.INIT('hc8)
	) name8564 (
		_w3683_,
		_w5100_,
		_w9740_,
		_w9914_
	);
	LUT3 #(
		.INIT('h02)
	) name8565 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w3712_,
		_w3727_,
		_w9915_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8566 (
		_w3469_,
		_w3470_,
		_w3728_,
		_w9915_,
		_w9916_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8567 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3684_,
		_w4953_,
		_w9917_
	);
	LUT2 #(
		.INIT('h4)
	) name8568 (
		_w9916_,
		_w9917_,
		_w9918_
	);
	LUT2 #(
		.INIT('h2)
	) name8569 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w3545_,
		_w9919_
	);
	LUT4 #(
		.INIT('hc055)
	) name8570 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3727_,
		_w9920_
	);
	LUT3 #(
		.INIT('h31)
	) name8571 (
		_w2248_,
		_w9919_,
		_w9920_,
		_w9921_
	);
	LUT2 #(
		.INIT('h4)
	) name8572 (
		_w9918_,
		_w9921_,
		_w9922_
	);
	LUT3 #(
		.INIT('h4f)
	) name8573 (
		_w9913_,
		_w9914_,
		_w9922_,
		_w9923_
	);
	LUT3 #(
		.INIT('h60)
	) name8574 (
		_w3513_,
		_w3516_,
		_w3682_,
		_w9924_
	);
	LUT3 #(
		.INIT('hc8)
	) name8575 (
		_w3682_,
		_w5111_,
		_w9740_,
		_w9925_
	);
	LUT3 #(
		.INIT('h02)
	) name8576 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w3727_,
		_w3742_,
		_w9926_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8577 (
		_w3469_,
		_w3470_,
		_w3743_,
		_w9926_,
		_w9927_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8578 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3713_,
		_w4953_,
		_w9928_
	);
	LUT2 #(
		.INIT('h4)
	) name8579 (
		_w9927_,
		_w9928_,
		_w9929_
	);
	LUT2 #(
		.INIT('h2)
	) name8580 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w3545_,
		_w9930_
	);
	LUT4 #(
		.INIT('hc055)
	) name8581 (
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3742_,
		_w9931_
	);
	LUT3 #(
		.INIT('h31)
	) name8582 (
		_w2248_,
		_w9930_,
		_w9931_,
		_w9932_
	);
	LUT2 #(
		.INIT('h4)
	) name8583 (
		_w9929_,
		_w9932_,
		_w9933_
	);
	LUT3 #(
		.INIT('h4f)
	) name8584 (
		_w9924_,
		_w9925_,
		_w9933_,
		_w9934_
	);
	LUT3 #(
		.INIT('h60)
	) name8585 (
		_w3513_,
		_w3516_,
		_w3712_,
		_w9935_
	);
	LUT3 #(
		.INIT('hc8)
	) name8586 (
		_w3712_,
		_w5122_,
		_w9740_,
		_w9936_
	);
	LUT3 #(
		.INIT('h02)
	) name8587 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w3592_,
		_w3742_,
		_w9937_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8588 (
		_w3469_,
		_w3470_,
		_w3757_,
		_w9937_,
		_w9938_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8589 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3728_,
		_w4953_,
		_w9939_
	);
	LUT2 #(
		.INIT('h4)
	) name8590 (
		_w9938_,
		_w9939_,
		_w9940_
	);
	LUT2 #(
		.INIT('h2)
	) name8591 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w3545_,
		_w9941_
	);
	LUT4 #(
		.INIT('hc055)
	) name8592 (
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3592_,
		_w9942_
	);
	LUT3 #(
		.INIT('h31)
	) name8593 (
		_w2248_,
		_w9941_,
		_w9942_,
		_w9943_
	);
	LUT2 #(
		.INIT('h4)
	) name8594 (
		_w9940_,
		_w9943_,
		_w9944_
	);
	LUT3 #(
		.INIT('h4f)
	) name8595 (
		_w9935_,
		_w9936_,
		_w9944_,
		_w9945_
	);
	LUT3 #(
		.INIT('h60)
	) name8596 (
		_w3513_,
		_w3516_,
		_w3727_,
		_w9946_
	);
	LUT3 #(
		.INIT('hc8)
	) name8597 (
		_w3727_,
		_w5133_,
		_w9740_,
		_w9947_
	);
	LUT3 #(
		.INIT('h02)
	) name8598 (
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w3411_,
		_w3592_,
		_w9948_
	);
	LUT4 #(
		.INIT('h00f1)
	) name8599 (
		_w3469_,
		_w3470_,
		_w3593_,
		_w9948_,
		_w9949_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8600 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3743_,
		_w4953_,
		_w9950_
	);
	LUT2 #(
		.INIT('h4)
	) name8601 (
		_w9949_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h2)
	) name8602 (
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w3545_,
		_w9952_
	);
	LUT4 #(
		.INIT('hc055)
	) name8603 (
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3411_,
		_w9953_
	);
	LUT3 #(
		.INIT('h31)
	) name8604 (
		_w2248_,
		_w9952_,
		_w9953_,
		_w9954_
	);
	LUT2 #(
		.INIT('h4)
	) name8605 (
		_w9951_,
		_w9954_,
		_w9955_
	);
	LUT3 #(
		.INIT('h4f)
	) name8606 (
		_w9946_,
		_w9947_,
		_w9955_,
		_w9956_
	);
	LUT3 #(
		.INIT('h60)
	) name8607 (
		_w3513_,
		_w3516_,
		_w3742_,
		_w9957_
	);
	LUT3 #(
		.INIT('hc8)
	) name8608 (
		_w3742_,
		_w5144_,
		_w9740_,
		_w9958_
	);
	LUT3 #(
		.INIT('h02)
	) name8609 (
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w3411_,
		_w3412_,
		_w9959_
	);
	LUT4 #(
		.INIT('h00ab)
	) name8610 (
		_w3413_,
		_w3469_,
		_w3470_,
		_w9959_,
		_w9960_
	);
	LUT4 #(
		.INIT('h00fd)
	) name8611 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w3407_,
		_w3757_,
		_w4953_,
		_w9961_
	);
	LUT2 #(
		.INIT('h4)
	) name8612 (
		_w9960_,
		_w9961_,
		_w9962_
	);
	LUT2 #(
		.INIT('h2)
	) name8613 (
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w3545_,
		_w9963_
	);
	LUT4 #(
		.INIT('hc055)
	) name8614 (
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1742_,
		_w1747_,
		_w3412_,
		_w9964_
	);
	LUT3 #(
		.INIT('h31)
	) name8615 (
		_w2248_,
		_w9963_,
		_w9964_,
		_w9965_
	);
	LUT2 #(
		.INIT('h4)
	) name8616 (
		_w9962_,
		_w9965_,
		_w9966_
	);
	LUT3 #(
		.INIT('h4f)
	) name8617 (
		_w9957_,
		_w9958_,
		_w9966_,
		_w9967_
	);
	LUT4 #(
		.INIT('h070f)
	) name8618 (
		\P1_EAX_reg[22]/NET0131 ,
		\P1_EAX_reg[23]/NET0131 ,
		\P1_EAX_reg[24]/NET0131 ,
		_w9484_,
		_w9968_
	);
	LUT3 #(
		.INIT('h02)
	) name8619 (
		_w1797_,
		_w9486_,
		_w9968_,
		_w9969_
	);
	LUT4 #(
		.INIT('h0008)
	) name8620 (
		_w1797_,
		_w1859_,
		_w9486_,
		_w9968_,
		_w9970_
	);
	LUT4 #(
		.INIT('hf020)
	) name8621 (
		\P1_Datao_reg[24]/NET0131 ,
		_w1860_,
		_w1933_,
		_w9970_,
		_w9971_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8622 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w9972_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8623 (
		\P1_Datao_reg[24]/NET0131 ,
		\P1_uWord_reg[8]/NET0131 ,
		_w1935_,
		_w9972_,
		_w9973_
	);
	LUT2 #(
		.INIT('hb)
	) name8624 (
		_w9971_,
		_w9973_,
		_w9974_
	);
	LUT4 #(
		.INIT('h4080)
	) name8625 (
		\P3_EAX_reg[24]/NET0131 ,
		_w2060_,
		_w2047_,
		_w9540_,
		_w9975_
	);
	LUT4 #(
		.INIT('h115d)
	) name8626 (
		\datao[24]_pad ,
		_w2112_,
		_w2114_,
		_w9975_,
		_w9976_
	);
	LUT4 #(
		.INIT('h0040)
	) name8627 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9977_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8628 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w9978_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8629 (
		\P3_uWord_reg[8]/NET0131 ,
		\datao[24]_pad ,
		_w9977_,
		_w9978_,
		_w9979_
	);
	LUT3 #(
		.INIT('h2f)
	) name8630 (
		_w1945_,
		_w9976_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h2)
	) name8631 (
		\datao[28]_pad ,
		_w2115_,
		_w9981_
	);
	LUT4 #(
		.INIT('h1020)
	) name8632 (
		\P3_EAX_reg[28]/NET0131 ,
		_w2111_,
		_w9543_,
		_w9542_,
		_w9982_
	);
	LUT4 #(
		.INIT('h5f13)
	) name8633 (
		\P3_uWord_reg[12]/NET0131 ,
		\datao[28]_pad ,
		_w9977_,
		_w9978_,
		_w9983_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name8634 (
		_w1945_,
		_w9981_,
		_w9982_,
		_w9983_,
		_w9984_
	);
	LUT4 #(
		.INIT('h4080)
	) name8635 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1797_,
		_w1859_,
		_w9487_,
		_w9985_
	);
	LUT4 #(
		.INIT('hf020)
	) name8636 (
		\P1_Datao_reg[28]/NET0131 ,
		_w1860_,
		_w1933_,
		_w9985_,
		_w9986_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8637 (
		\P1_Datao_reg[28]/NET0131 ,
		\P1_uWord_reg[12]/NET0131 ,
		_w1935_,
		_w9972_,
		_w9987_
	);
	LUT2 #(
		.INIT('hb)
	) name8638 (
		_w9986_,
		_w9987_,
		_w9988_
	);
	LUT3 #(
		.INIT('h40)
	) name8639 (
		_w1501_,
		_w1568_,
		_w1611_,
		_w9989_
	);
	LUT4 #(
		.INIT('h8000)
	) name8640 (
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		_w7781_,
		_w9459_,
		_w9990_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name8641 (
		\P2_EAX_reg[23]/NET0131 ,
		\P2_EAX_reg[24]/NET0131 ,
		_w7781_,
		_w9459_,
		_w9991_
	);
	LUT4 #(
		.INIT('h2220)
	) name8642 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w9991_,
		_w9992_
	);
	LUT4 #(
		.INIT('haaa2)
	) name8643 (
		\P2_Datao_reg[24]/NET0131 ,
		_w4927_,
		_w9989_,
		_w9992_,
		_w9993_
	);
	LUT4 #(
		.INIT('h0200)
	) name8644 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w9991_,
		_w9994_
	);
	LUT4 #(
		.INIT('h0040)
	) name8645 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9995_
	);
	LUT4 #(
		.INIT('hfc60)
	) name8646 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w9996_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8647 (
		\P2_Datao_reg[24]/NET0131 ,
		\P2_uWord_reg[8]/NET0131 ,
		_w9995_,
		_w9996_,
		_w9997_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name8648 (
		_w1678_,
		_w9993_,
		_w9994_,
		_w9997_,
		_w9998_
	);
	LUT4 #(
		.INIT('h4080)
	) name8649 (
		\P2_EAX_reg[28]/NET0131 ,
		_w1566_,
		_w1674_,
		_w9461_,
		_w9999_
	);
	LUT4 #(
		.INIT('h0075)
	) name8650 (
		\P2_Datao_reg[28]/NET0131 ,
		_w1602_,
		_w1616_,
		_w9999_,
		_w10000_
	);
	LUT4 #(
		.INIT('h3f15)
	) name8651 (
		\P2_Datao_reg[28]/NET0131 ,
		\P2_uWord_reg[12]/NET0131 ,
		_w9995_,
		_w9996_,
		_w10001_
	);
	LUT3 #(
		.INIT('h2f)
	) name8652 (
		_w1678_,
		_w10000_,
		_w10001_,
		_w10002_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8653 (
		\P2_uWord_reg[8]/NET0131 ,
		_w1678_,
		_w7767_,
		_w9467_,
		_w10003_
	);
	LUT4 #(
		.INIT('h0222)
	) name8654 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[8]/NET0131 ,
		_w2255_,
		_w2260_,
		_w10004_
	);
	LUT4 #(
		.INIT('h3111)
	) name8655 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[8]/NET0131 ,
		_w2255_,
		_w2260_,
		_w10005_
	);
	LUT3 #(
		.INIT('h01)
	) name8656 (
		_w1605_,
		_w10005_,
		_w10004_,
		_w10006_
	);
	LUT2 #(
		.INIT('h8)
	) name8657 (
		_w1565_,
		_w10006_,
		_w10007_
	);
	LUT4 #(
		.INIT('h153f)
	) name8658 (
		_w1565_,
		_w1566_,
		_w9991_,
		_w10006_,
		_w10008_
	);
	LUT3 #(
		.INIT('hd0)
	) name8659 (
		_w1592_,
		_w1601_,
		_w1678_,
		_w10009_
	);
	LUT2 #(
		.INIT('h4)
	) name8660 (
		_w10008_,
		_w10009_,
		_w10010_
	);
	LUT2 #(
		.INIT('he)
	) name8661 (
		_w10003_,
		_w10010_,
		_w10011_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8662 (
		\P1_uWord_reg[8]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w10012_
	);
	LUT3 #(
		.INIT('h02)
	) name8663 (
		_w1795_,
		_w1861_,
		_w3435_,
		_w10013_
	);
	LUT3 #(
		.INIT('ha8)
	) name8664 (
		_w9489_,
		_w9969_,
		_w10013_,
		_w10014_
	);
	LUT2 #(
		.INIT('he)
	) name8665 (
		_w10012_,
		_w10014_,
		_w10015_
	);
	LUT4 #(
		.INIT('h4c44)
	) name8666 (
		_w1933_,
		_w9102_,
		_w9436_,
		_w9437_,
		_w10016_
	);
	LUT2 #(
		.INIT('h2)
	) name8667 (
		_w1846_,
		_w3195_,
		_w10017_
	);
	LUT4 #(
		.INIT('h4000)
	) name8668 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10017_,
		_w10018_
	);
	LUT2 #(
		.INIT('h2)
	) name8669 (
		_w1867_,
		_w3481_,
		_w10019_
	);
	LUT4 #(
		.INIT('hec00)
	) name8670 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10019_,
		_w10020_
	);
	LUT3 #(
		.INIT('h78)
	) name8671 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		_w10021_
	);
	LUT3 #(
		.INIT('h80)
	) name8672 (
		_w1804_,
		_w1826_,
		_w10021_,
		_w10022_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8673 (
		_w1933_,
		_w10020_,
		_w10018_,
		_w10022_,
		_w10023_
	);
	LUT3 #(
		.INIT('hf2)
	) name8674 (
		\P1_EAX_reg[2]/NET0131 ,
		_w10016_,
		_w10023_,
		_w10024_
	);
	LUT2 #(
		.INIT('h2)
	) name8675 (
		\P3_EAX_reg[10]/NET0131 ,
		_w8341_,
		_w10025_
	);
	LUT3 #(
		.INIT('h08)
	) name8676 (
		_w2063_,
		_w2075_,
		_w8346_,
		_w10026_
	);
	LUT4 #(
		.INIT('h0001)
	) name8677 (
		_w2120_,
		_w2121_,
		_w8367_,
		_w10026_,
		_w10027_
	);
	LUT3 #(
		.INIT('h08)
	) name8678 (
		\buf2_reg[10]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10028_
	);
	LUT4 #(
		.INIT('h153f)
	) name8679 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1954_,
		_w1961_,
		_w10029_
	);
	LUT4 #(
		.INIT('h153f)
	) name8680 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10030_
	);
	LUT4 #(
		.INIT('h153f)
	) name8681 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1946_,
		_w1967_,
		_w10031_
	);
	LUT4 #(
		.INIT('h135f)
	) name8682 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1966_,
		_w1969_,
		_w10032_
	);
	LUT4 #(
		.INIT('h8000)
	) name8683 (
		_w10031_,
		_w10032_,
		_w10029_,
		_w10030_,
		_w10033_
	);
	LUT4 #(
		.INIT('h135f)
	) name8684 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w1956_,
		_w1957_,
		_w10034_
	);
	LUT4 #(
		.INIT('h153f)
	) name8685 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10035_
	);
	LUT4 #(
		.INIT('h135f)
	) name8686 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1960_,
		_w1964_,
		_w10036_
	);
	LUT4 #(
		.INIT('h153f)
	) name8687 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1949_,
		_w1963_,
		_w10037_
	);
	LUT4 #(
		.INIT('h8000)
	) name8688 (
		_w10036_,
		_w10037_,
		_w10034_,
		_w10035_,
		_w10038_
	);
	LUT2 #(
		.INIT('h8)
	) name8689 (
		_w10033_,
		_w10038_,
		_w10039_
	);
	LUT4 #(
		.INIT('h4000)
	) name8690 (
		\P3_EAX_reg[10]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8345_,
		_w10040_
	);
	LUT3 #(
		.INIT('h0d)
	) name8691 (
		_w8366_,
		_w10039_,
		_w10040_,
		_w10041_
	);
	LUT2 #(
		.INIT('h4)
	) name8692 (
		_w10028_,
		_w10041_,
		_w10042_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8693 (
		\P3_EAX_reg[10]/NET0131 ,
		_w1945_,
		_w10027_,
		_w10042_,
		_w10043_
	);
	LUT2 #(
		.INIT('he)
	) name8694 (
		_w10025_,
		_w10043_,
		_w10044_
	);
	LUT4 #(
		.INIT('h0111)
	) name8695 (
		_w1842_,
		_w1845_,
		_w3175_,
		_w3180_,
		_w10045_
	);
	LUT4 #(
		.INIT('h4000)
	) name8696 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h2)
	) name8697 (
		_w1867_,
		_w3428_,
		_w10047_
	);
	LUT4 #(
		.INIT('hec00)
	) name8698 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10047_,
		_w10048_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8699 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w10049_
	);
	LUT3 #(
		.INIT('h80)
	) name8700 (
		_w1804_,
		_w1826_,
		_w10049_,
		_w10050_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8701 (
		_w1933_,
		_w10048_,
		_w10046_,
		_w10050_,
		_w10051_
	);
	LUT3 #(
		.INIT('hf2)
	) name8702 (
		\P1_EAX_reg[3]/NET0131 ,
		_w10016_,
		_w10051_,
		_w10052_
	);
	LUT2 #(
		.INIT('h2)
	) name8703 (
		\P3_EAX_reg[11]/NET0131 ,
		_w8341_,
		_w10053_
	);
	LUT4 #(
		.INIT('h135f)
	) name8704 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[11][3]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10054_
	);
	LUT4 #(
		.INIT('h135f)
	) name8705 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10055_
	);
	LUT4 #(
		.INIT('h135f)
	) name8706 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10056_
	);
	LUT4 #(
		.INIT('h153f)
	) name8707 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10057_
	);
	LUT4 #(
		.INIT('h8000)
	) name8708 (
		_w10056_,
		_w10057_,
		_w10054_,
		_w10055_,
		_w10058_
	);
	LUT4 #(
		.INIT('h135f)
	) name8709 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10059_
	);
	LUT4 #(
		.INIT('h153f)
	) name8710 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10060_
	);
	LUT4 #(
		.INIT('h153f)
	) name8711 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10061_
	);
	LUT4 #(
		.INIT('h153f)
	) name8712 (
		\P3_InstQueue_reg[7][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10062_
	);
	LUT4 #(
		.INIT('h8000)
	) name8713 (
		_w10061_,
		_w10062_,
		_w10059_,
		_w10060_,
		_w10063_
	);
	LUT2 #(
		.INIT('h8)
	) name8714 (
		_w10058_,
		_w10063_,
		_w10064_
	);
	LUT3 #(
		.INIT('h08)
	) name8715 (
		_w2063_,
		_w2075_,
		_w8347_,
		_w10065_
	);
	LUT4 #(
		.INIT('h4000)
	) name8716 (
		\P3_EAX_reg[11]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8346_,
		_w10066_
	);
	LUT4 #(
		.INIT('hd800)
	) name8717 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w8439_,
		_w10067_
	);
	LUT4 #(
		.INIT('h0031)
	) name8718 (
		_w8366_,
		_w10066_,
		_w10064_,
		_w10067_,
		_w10068_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8719 (
		\P3_EAX_reg[11]/NET0131 ,
		_w1945_,
		_w10027_,
		_w10068_,
		_w10069_
	);
	LUT2 #(
		.INIT('he)
	) name8720 (
		_w10053_,
		_w10069_,
		_w10070_
	);
	LUT2 #(
		.INIT('h2)
	) name8721 (
		\P3_EAX_reg[12]/NET0131 ,
		_w8341_,
		_w10071_
	);
	LUT4 #(
		.INIT('h5553)
	) name8722 (
		\P3_EAX_reg[12]/NET0131 ,
		\buf2_reg[12]/NET0131 ,
		_w2105_,
		_w2116_,
		_w10072_
	);
	LUT4 #(
		.INIT('h00d8)
	) name8723 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w10072_,
		_w10073_
	);
	LUT4 #(
		.INIT('h135f)
	) name8724 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10074_
	);
	LUT4 #(
		.INIT('h135f)
	) name8725 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10075_
	);
	LUT4 #(
		.INIT('h135f)
	) name8726 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10076_
	);
	LUT4 #(
		.INIT('h153f)
	) name8727 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10077_
	);
	LUT4 #(
		.INIT('h8000)
	) name8728 (
		_w10076_,
		_w10077_,
		_w10074_,
		_w10075_,
		_w10078_
	);
	LUT4 #(
		.INIT('h135f)
	) name8729 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10079_
	);
	LUT4 #(
		.INIT('h153f)
	) name8730 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10080_
	);
	LUT4 #(
		.INIT('h153f)
	) name8731 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10081_
	);
	LUT4 #(
		.INIT('h153f)
	) name8732 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10082_
	);
	LUT4 #(
		.INIT('h8000)
	) name8733 (
		_w10081_,
		_w10082_,
		_w10079_,
		_w10080_,
		_w10083_
	);
	LUT2 #(
		.INIT('h8)
	) name8734 (
		_w10078_,
		_w10083_,
		_w10084_
	);
	LUT4 #(
		.INIT('h4000)
	) name8735 (
		\P3_EAX_reg[12]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8347_,
		_w10085_
	);
	LUT4 #(
		.INIT('h000d)
	) name8736 (
		_w8366_,
		_w10084_,
		_w10073_,
		_w10085_,
		_w10086_
	);
	LUT4 #(
		.INIT('h5700)
	) name8737 (
		\P3_EAX_reg[12]/NET0131 ,
		_w8367_,
		_w10065_,
		_w10086_,
		_w10087_
	);
	LUT3 #(
		.INIT('hce)
	) name8738 (
		_w1945_,
		_w10071_,
		_w10087_,
		_w10088_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8739 (
		_w1945_,
		_w2120_,
		_w2121_,
		_w8367_,
		_w10089_
	);
	LUT4 #(
		.INIT('h4080)
	) name8740 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8348_,
		_w10090_
	);
	LUT4 #(
		.INIT('h135f)
	) name8741 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10091_
	);
	LUT4 #(
		.INIT('h135f)
	) name8742 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10092_
	);
	LUT4 #(
		.INIT('h135f)
	) name8743 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10093_
	);
	LUT4 #(
		.INIT('h153f)
	) name8744 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10094_
	);
	LUT4 #(
		.INIT('h8000)
	) name8745 (
		_w10093_,
		_w10094_,
		_w10091_,
		_w10092_,
		_w10095_
	);
	LUT4 #(
		.INIT('h135f)
	) name8746 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10096_
	);
	LUT4 #(
		.INIT('h153f)
	) name8747 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10097_
	);
	LUT4 #(
		.INIT('h153f)
	) name8748 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10098_
	);
	LUT4 #(
		.INIT('h153f)
	) name8749 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10099_
	);
	LUT4 #(
		.INIT('h8000)
	) name8750 (
		_w10098_,
		_w10099_,
		_w10096_,
		_w10097_,
		_w10100_
	);
	LUT2 #(
		.INIT('h8)
	) name8751 (
		_w10095_,
		_w10100_,
		_w10101_
	);
	LUT2 #(
		.INIT('h2)
	) name8752 (
		_w8366_,
		_w10101_,
		_w10102_
	);
	LUT3 #(
		.INIT('h08)
	) name8753 (
		\buf2_reg[13]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10103_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8754 (
		_w1945_,
		_w10102_,
		_w10103_,
		_w10090_,
		_w10104_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8755 (
		\P3_EAX_reg[13]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10104_,
		_w10105_
	);
	LUT4 #(
		.INIT('h4080)
	) name8756 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8349_,
		_w10106_
	);
	LUT3 #(
		.INIT('h08)
	) name8757 (
		\buf2_reg[14]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10107_
	);
	LUT4 #(
		.INIT('h135f)
	) name8758 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10108_
	);
	LUT4 #(
		.INIT('h135f)
	) name8759 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10109_
	);
	LUT4 #(
		.INIT('h135f)
	) name8760 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10110_
	);
	LUT4 #(
		.INIT('h153f)
	) name8761 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10111_
	);
	LUT4 #(
		.INIT('h8000)
	) name8762 (
		_w10110_,
		_w10111_,
		_w10108_,
		_w10109_,
		_w10112_
	);
	LUT4 #(
		.INIT('h135f)
	) name8763 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10113_
	);
	LUT4 #(
		.INIT('h153f)
	) name8764 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10114_
	);
	LUT4 #(
		.INIT('h153f)
	) name8765 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10115_
	);
	LUT4 #(
		.INIT('h153f)
	) name8766 (
		\P3_InstQueue_reg[7][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10116_
	);
	LUT4 #(
		.INIT('h8000)
	) name8767 (
		_w10115_,
		_w10116_,
		_w10113_,
		_w10114_,
		_w10117_
	);
	LUT2 #(
		.INIT('h8)
	) name8768 (
		_w10112_,
		_w10117_,
		_w10118_
	);
	LUT2 #(
		.INIT('h2)
	) name8769 (
		_w8366_,
		_w10118_,
		_w10119_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8770 (
		_w1945_,
		_w10107_,
		_w10119_,
		_w10106_,
		_w10120_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8771 (
		\P3_EAX_reg[14]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10120_,
		_w10121_
	);
	LUT3 #(
		.INIT('h08)
	) name8772 (
		_w2063_,
		_w2075_,
		_w8351_,
		_w10122_
	);
	LUT4 #(
		.INIT('h4080)
	) name8773 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8350_,
		_w10123_
	);
	LUT3 #(
		.INIT('h02)
	) name8774 (
		\buf2_reg[15]/NET0131 ,
		_w2105_,
		_w2116_,
		_w10124_
	);
	LUT4 #(
		.INIT('hd800)
	) name8775 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w10124_,
		_w10125_
	);
	LUT4 #(
		.INIT('h135f)
	) name8776 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		\P3_InstQueue_reg[11][7]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10126_
	);
	LUT4 #(
		.INIT('h135f)
	) name8777 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10127_
	);
	LUT4 #(
		.INIT('h135f)
	) name8778 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10128_
	);
	LUT4 #(
		.INIT('h153f)
	) name8779 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10129_
	);
	LUT4 #(
		.INIT('h8000)
	) name8780 (
		_w10128_,
		_w10129_,
		_w10126_,
		_w10127_,
		_w10130_
	);
	LUT4 #(
		.INIT('h135f)
	) name8781 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10131_
	);
	LUT4 #(
		.INIT('h153f)
	) name8782 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10132_
	);
	LUT4 #(
		.INIT('h153f)
	) name8783 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10133_
	);
	LUT4 #(
		.INIT('h153f)
	) name8784 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10134_
	);
	LUT4 #(
		.INIT('h8000)
	) name8785 (
		_w10133_,
		_w10134_,
		_w10131_,
		_w10132_,
		_w10135_
	);
	LUT2 #(
		.INIT('h8)
	) name8786 (
		_w10130_,
		_w10135_,
		_w10136_
	);
	LUT4 #(
		.INIT('h0301)
	) name8787 (
		_w8366_,
		_w10125_,
		_w10123_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h2)
	) name8788 (
		_w1945_,
		_w10137_,
		_w10138_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8789 (
		\P3_EAX_reg[15]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10138_,
		_w10139_
	);
	LUT3 #(
		.INIT('h02)
	) name8790 (
		_w1855_,
		_w1861_,
		_w3442_,
		_w10140_
	);
	LUT4 #(
		.INIT('h0111)
	) name8791 (
		_w1842_,
		_w1845_,
		_w3136_,
		_w3141_,
		_w10141_
	);
	LUT4 #(
		.INIT('h4000)
	) name8792 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('h6)
	) name8793 (
		\P1_EAX_reg[4]/NET0131 ,
		_w9418_,
		_w10143_
	);
	LUT3 #(
		.INIT('h80)
	) name8794 (
		_w1804_,
		_w1826_,
		_w10143_,
		_w10144_
	);
	LUT2 #(
		.INIT('h1)
	) name8795 (
		_w10142_,
		_w10144_,
		_w10145_
	);
	LUT3 #(
		.INIT('h8a)
	) name8796 (
		_w1933_,
		_w10140_,
		_w10145_,
		_w10146_
	);
	LUT3 #(
		.INIT('hf2)
	) name8797 (
		\P1_EAX_reg[4]/NET0131 ,
		_w10016_,
		_w10146_,
		_w10147_
	);
	LUT2 #(
		.INIT('h2)
	) name8798 (
		\P3_EAX_reg[1]/NET0131 ,
		_w8341_,
		_w10148_
	);
	LUT3 #(
		.INIT('h40)
	) name8799 (
		\P3_EAX_reg[0]/NET0131 ,
		_w2063_,
		_w2075_,
		_w10149_
	);
	LUT4 #(
		.INIT('h0001)
	) name8800 (
		_w2120_,
		_w2121_,
		_w8367_,
		_w10149_,
		_w10150_
	);
	LUT3 #(
		.INIT('h02)
	) name8801 (
		\buf2_reg[1]/NET0131 ,
		_w2105_,
		_w2116_,
		_w10151_
	);
	LUT4 #(
		.INIT('hd800)
	) name8802 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w10151_,
		_w10152_
	);
	LUT2 #(
		.INIT('h2)
	) name8803 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		_w10153_
	);
	LUT3 #(
		.INIT('h80)
	) name8804 (
		_w2063_,
		_w2075_,
		_w10153_,
		_w10154_
	);
	LUT4 #(
		.INIT('h000b)
	) name8805 (
		_w2783_,
		_w8366_,
		_w10152_,
		_w10154_,
		_w10155_
	);
	LUT4 #(
		.INIT('h08cc)
	) name8806 (
		\P3_EAX_reg[1]/NET0131 ,
		_w1945_,
		_w10150_,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('he)
	) name8807 (
		_w10148_,
		_w10156_,
		_w10157_
	);
	LUT3 #(
		.INIT('h02)
	) name8808 (
		_w1855_,
		_w1861_,
		_w3452_,
		_w10158_
	);
	LUT4 #(
		.INIT('h0111)
	) name8809 (
		_w1842_,
		_w1845_,
		_w3108_,
		_w3113_,
		_w10159_
	);
	LUT4 #(
		.INIT('h4000)
	) name8810 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10159_,
		_w10160_
	);
	LUT3 #(
		.INIT('h6c)
	) name8811 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w9418_,
		_w10161_
	);
	LUT3 #(
		.INIT('h80)
	) name8812 (
		_w1804_,
		_w1826_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('h1)
	) name8813 (
		_w10160_,
		_w10162_,
		_w10163_
	);
	LUT3 #(
		.INIT('h8a)
	) name8814 (
		_w1933_,
		_w10158_,
		_w10163_,
		_w10164_
	);
	LUT3 #(
		.INIT('hf2)
	) name8815 (
		\P1_EAX_reg[5]/NET0131 ,
		_w10016_,
		_w10164_,
		_w10165_
	);
	LUT3 #(
		.INIT('h08)
	) name8816 (
		\buf2_reg[2]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10166_
	);
	LUT3 #(
		.INIT('h78)
	) name8817 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		_w10167_
	);
	LUT3 #(
		.INIT('h80)
	) name8818 (
		_w2063_,
		_w2075_,
		_w10167_,
		_w10168_
	);
	LUT3 #(
		.INIT('h0b)
	) name8819 (
		_w2769_,
		_w8366_,
		_w10168_,
		_w10169_
	);
	LUT3 #(
		.INIT('h8a)
	) name8820 (
		_w1945_,
		_w10166_,
		_w10169_,
		_w10170_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8821 (
		\P3_EAX_reg[2]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10170_,
		_w10171_
	);
	LUT3 #(
		.INIT('h08)
	) name8822 (
		\buf2_reg[3]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10172_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8823 (
		\P3_EAX_reg[0]/NET0131 ,
		\P3_EAX_reg[1]/NET0131 ,
		\P3_EAX_reg[2]/NET0131 ,
		\P3_EAX_reg[3]/NET0131 ,
		_w10173_
	);
	LUT3 #(
		.INIT('h80)
	) name8824 (
		_w2063_,
		_w2075_,
		_w10173_,
		_w10174_
	);
	LUT3 #(
		.INIT('h0b)
	) name8825 (
		_w2809_,
		_w8366_,
		_w10174_,
		_w10175_
	);
	LUT3 #(
		.INIT('h8a)
	) name8826 (
		_w1945_,
		_w10172_,
		_w10175_,
		_w10176_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8827 (
		\P3_EAX_reg[3]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10176_,
		_w10177_
	);
	LUT3 #(
		.INIT('h02)
	) name8828 (
		_w1855_,
		_w1861_,
		_w3438_,
		_w10178_
	);
	LUT4 #(
		.INIT('h0111)
	) name8829 (
		_w1842_,
		_w1845_,
		_w3095_,
		_w3100_,
		_w10179_
	);
	LUT4 #(
		.INIT('h4000)
	) name8830 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('h6)
	) name8831 (
		\P1_EAX_reg[7]/NET0131 ,
		_w9419_,
		_w10181_
	);
	LUT3 #(
		.INIT('h80)
	) name8832 (
		_w1804_,
		_w1826_,
		_w10181_,
		_w10182_
	);
	LUT2 #(
		.INIT('h1)
	) name8833 (
		_w10180_,
		_w10182_,
		_w10183_
	);
	LUT3 #(
		.INIT('h8a)
	) name8834 (
		_w1933_,
		_w10178_,
		_w10183_,
		_w10184_
	);
	LUT3 #(
		.INIT('hf2)
	) name8835 (
		\P1_EAX_reg[7]/NET0131 ,
		_w10016_,
		_w10184_,
		_w10185_
	);
	LUT3 #(
		.INIT('h08)
	) name8836 (
		\buf2_reg[4]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10186_
	);
	LUT2 #(
		.INIT('h6)
	) name8837 (
		\P3_EAX_reg[4]/NET0131 ,
		_w8343_,
		_w10187_
	);
	LUT3 #(
		.INIT('h80)
	) name8838 (
		_w2063_,
		_w2075_,
		_w10187_,
		_w10188_
	);
	LUT3 #(
		.INIT('h0b)
	) name8839 (
		_w2824_,
		_w8366_,
		_w10188_,
		_w10189_
	);
	LUT3 #(
		.INIT('h8a)
	) name8840 (
		_w1945_,
		_w10186_,
		_w10189_,
		_w10190_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8841 (
		\P3_EAX_reg[4]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10190_,
		_w10191_
	);
	LUT3 #(
		.INIT('h08)
	) name8842 (
		\buf2_reg[5]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10192_
	);
	LUT3 #(
		.INIT('h6c)
	) name8843 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		_w8343_,
		_w10193_
	);
	LUT3 #(
		.INIT('h80)
	) name8844 (
		_w2063_,
		_w2075_,
		_w10193_,
		_w10194_
	);
	LUT3 #(
		.INIT('h0b)
	) name8845 (
		_w2855_,
		_w8366_,
		_w10194_,
		_w10195_
	);
	LUT3 #(
		.INIT('h8a)
	) name8846 (
		_w1945_,
		_w10192_,
		_w10195_,
		_w10196_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8847 (
		\P3_EAX_reg[5]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10196_,
		_w10197_
	);
	LUT3 #(
		.INIT('h08)
	) name8848 (
		\buf2_reg[6]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10198_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8849 (
		\P3_EAX_reg[4]/NET0131 ,
		\P3_EAX_reg[5]/NET0131 ,
		\P3_EAX_reg[6]/NET0131 ,
		_w8343_,
		_w10199_
	);
	LUT3 #(
		.INIT('h80)
	) name8850 (
		_w2063_,
		_w2075_,
		_w10199_,
		_w10200_
	);
	LUT3 #(
		.INIT('h0b)
	) name8851 (
		_w2842_,
		_w8366_,
		_w10200_,
		_w10201_
	);
	LUT3 #(
		.INIT('h8a)
	) name8852 (
		_w1945_,
		_w10198_,
		_w10201_,
		_w10202_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8853 (
		\P3_EAX_reg[6]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10202_,
		_w10203_
	);
	LUT3 #(
		.INIT('h08)
	) name8854 (
		\buf2_reg[7]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10204_
	);
	LUT2 #(
		.INIT('h6)
	) name8855 (
		\P3_EAX_reg[7]/NET0131 ,
		_w8344_,
		_w10205_
	);
	LUT3 #(
		.INIT('h80)
	) name8856 (
		_w2063_,
		_w2075_,
		_w10205_,
		_w10206_
	);
	LUT3 #(
		.INIT('h0b)
	) name8857 (
		_w2755_,
		_w8366_,
		_w10206_,
		_w10207_
	);
	LUT3 #(
		.INIT('h8a)
	) name8858 (
		_w1945_,
		_w10204_,
		_w10207_,
		_w10208_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8859 (
		\P3_EAX_reg[7]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10208_,
		_w10209_
	);
	LUT3 #(
		.INIT('h08)
	) name8860 (
		\buf2_reg[8]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10210_
	);
	LUT4 #(
		.INIT('h135f)
	) name8861 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w1961_,
		_w1963_,
		_w10211_
	);
	LUT4 #(
		.INIT('h135f)
	) name8862 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w1956_,
		_w1969_,
		_w10212_
	);
	LUT4 #(
		.INIT('h135f)
	) name8863 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w1966_,
		_w1967_,
		_w10213_
	);
	LUT4 #(
		.INIT('h153f)
	) name8864 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w1947_,
		_w1950_,
		_w10214_
	);
	LUT4 #(
		.INIT('h8000)
	) name8865 (
		_w10213_,
		_w10214_,
		_w10211_,
		_w10212_,
		_w10215_
	);
	LUT4 #(
		.INIT('h135f)
	) name8866 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1957_,
		_w1946_,
		_w10216_
	);
	LUT4 #(
		.INIT('h153f)
	) name8867 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10217_
	);
	LUT4 #(
		.INIT('h153f)
	) name8868 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1949_,
		_w1960_,
		_w10218_
	);
	LUT4 #(
		.INIT('h153f)
	) name8869 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1954_,
		_w1964_,
		_w10219_
	);
	LUT4 #(
		.INIT('h8000)
	) name8870 (
		_w10218_,
		_w10219_,
		_w10216_,
		_w10217_,
		_w10220_
	);
	LUT2 #(
		.INIT('h8)
	) name8871 (
		_w10215_,
		_w10220_,
		_w10221_
	);
	LUT3 #(
		.INIT('h6c)
	) name8872 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		_w8344_,
		_w10222_
	);
	LUT3 #(
		.INIT('h80)
	) name8873 (
		_w2063_,
		_w2075_,
		_w10222_,
		_w10223_
	);
	LUT3 #(
		.INIT('h0d)
	) name8874 (
		_w8366_,
		_w10221_,
		_w10223_,
		_w10224_
	);
	LUT3 #(
		.INIT('h8a)
	) name8875 (
		_w1945_,
		_w10210_,
		_w10224_,
		_w10225_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8876 (
		\P3_EAX_reg[8]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10225_,
		_w10226_
	);
	LUT3 #(
		.INIT('h08)
	) name8877 (
		\buf2_reg[9]/NET0131 ,
		_w2108_,
		_w2116_,
		_w10227_
	);
	LUT4 #(
		.INIT('h153f)
	) name8878 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1954_,
		_w1961_,
		_w10228_
	);
	LUT4 #(
		.INIT('h135f)
	) name8879 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w1950_,
		_w1969_,
		_w10229_
	);
	LUT4 #(
		.INIT('h153f)
	) name8880 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1946_,
		_w1967_,
		_w10230_
	);
	LUT4 #(
		.INIT('h153f)
	) name8881 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1966_,
		_w1963_,
		_w10231_
	);
	LUT4 #(
		.INIT('h8000)
	) name8882 (
		_w10230_,
		_w10231_,
		_w10228_,
		_w10229_,
		_w10232_
	);
	LUT4 #(
		.INIT('h153f)
	) name8883 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1957_,
		_w1947_,
		_w10233_
	);
	LUT4 #(
		.INIT('h153f)
	) name8884 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1952_,
		_w1970_,
		_w10234_
	);
	LUT4 #(
		.INIT('h135f)
	) name8885 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1960_,
		_w1964_,
		_w10235_
	);
	LUT4 #(
		.INIT('h135f)
	) name8886 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1956_,
		_w1949_,
		_w10236_
	);
	LUT4 #(
		.INIT('h8000)
	) name8887 (
		_w10235_,
		_w10236_,
		_w10233_,
		_w10234_,
		_w10237_
	);
	LUT2 #(
		.INIT('h8)
	) name8888 (
		_w10232_,
		_w10237_,
		_w10238_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8889 (
		\P3_EAX_reg[7]/NET0131 ,
		\P3_EAX_reg[8]/NET0131 ,
		\P3_EAX_reg[9]/NET0131 ,
		_w8344_,
		_w10239_
	);
	LUT3 #(
		.INIT('h80)
	) name8890 (
		_w2063_,
		_w2075_,
		_w10239_,
		_w10240_
	);
	LUT3 #(
		.INIT('h0d)
	) name8891 (
		_w8366_,
		_w10238_,
		_w10240_,
		_w10241_
	);
	LUT3 #(
		.INIT('h8a)
	) name8892 (
		_w1945_,
		_w10227_,
		_w10241_,
		_w10242_
	);
	LUT4 #(
		.INIT('hffa2)
	) name8893 (
		\P3_EAX_reg[9]/NET0131 ,
		_w8341_,
		_w10089_,
		_w10242_,
		_w10243_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name8894 (
		\P2_EAX_reg[0]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10244_
	);
	LUT2 #(
		.INIT('h2)
	) name8895 (
		_w1606_,
		_w9115_,
		_w10245_
	);
	LUT4 #(
		.INIT('hec00)
	) name8896 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w10245_,
		_w10246_
	);
	LUT2 #(
		.INIT('h4)
	) name8897 (
		\P2_EAX_reg[0]/NET0131 ,
		_w7789_,
		_w10247_
	);
	LUT4 #(
		.INIT('h0111)
	) name8898 (
		_w1592_,
		_w1595_,
		_w4133_,
		_w4138_,
		_w10248_
	);
	LUT3 #(
		.INIT('h80)
	) name8899 (
		_w1549_,
		_w1553_,
		_w10248_,
		_w10249_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8900 (
		_w1678_,
		_w10247_,
		_w10249_,
		_w10246_,
		_w10250_
	);
	LUT2 #(
		.INIT('he)
	) name8901 (
		_w10244_,
		_w10250_,
		_w10251_
	);
	LUT2 #(
		.INIT('h2)
	) name8902 (
		\P3_EBX_reg[29]/NET0131 ,
		_w8341_,
		_w10252_
	);
	LUT3 #(
		.INIT('h80)
	) name8903 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		_w8920_,
		_w10253_
	);
	LUT4 #(
		.INIT('h8000)
	) name8904 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		_w8920_,
		_w10254_
	);
	LUT3 #(
		.INIT('h80)
	) name8905 (
		\P3_EBX_reg[28]/NET0131 ,
		_w9504_,
		_w10254_,
		_w10255_
	);
	LUT2 #(
		.INIT('h8)
	) name8906 (
		_w8923_,
		_w9668_,
		_w10256_
	);
	LUT4 #(
		.INIT('h0057)
	) name8907 (
		\P3_EBX_reg[29]/NET0131 ,
		_w8925_,
		_w9504_,
		_w10256_,
		_w10257_
	);
	LUT4 #(
		.INIT('hecee)
	) name8908 (
		_w1945_,
		_w10252_,
		_w10255_,
		_w10257_,
		_w10258_
	);
	LUT4 #(
		.INIT('h135f)
	) name8909 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[5][0]/NET0131 ,
		_w1712_,
		_w1702_,
		_w10259_
	);
	LUT4 #(
		.INIT('h153f)
	) name8910 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1711_,
		_w1705_,
		_w10260_
	);
	LUT4 #(
		.INIT('h135f)
	) name8911 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1696_,
		_w1706_,
		_w10261_
	);
	LUT4 #(
		.INIT('h135f)
	) name8912 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1694_,
		_w1692_,
		_w10262_
	);
	LUT4 #(
		.INIT('h8000)
	) name8913 (
		_w10261_,
		_w10262_,
		_w10259_,
		_w10260_,
		_w10263_
	);
	LUT4 #(
		.INIT('h135f)
	) name8914 (
		\P1_InstQueue_reg[14][0]/NET0131 ,
		\P1_InstQueue_reg[4][0]/NET0131 ,
		_w1698_,
		_w1709_,
		_w10264_
	);
	LUT4 #(
		.INIT('h153f)
	) name8915 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1708_,
		_w1703_,
		_w10265_
	);
	LUT4 #(
		.INIT('h135f)
	) name8916 (
		\P1_InstQueue_reg[2][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1688_,
		_w1689_,
		_w10266_
	);
	LUT4 #(
		.INIT('h135f)
	) name8917 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1699_,
		_w1691_,
		_w10267_
	);
	LUT4 #(
		.INIT('h8000)
	) name8918 (
		_w10266_,
		_w10267_,
		_w10264_,
		_w10265_,
		_w10268_
	);
	LUT4 #(
		.INIT('h0111)
	) name8919 (
		_w1842_,
		_w1845_,
		_w10263_,
		_w10268_,
		_w10269_
	);
	LUT4 #(
		.INIT('h4000)
	) name8920 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10269_,
		_w10270_
	);
	LUT2 #(
		.INIT('h2)
	) name8921 (
		_w1867_,
		_w3435_,
		_w10271_
	);
	LUT4 #(
		.INIT('hec00)
	) name8922 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10271_,
		_w10272_
	);
	LUT3 #(
		.INIT('h6c)
	) name8923 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		_w9419_,
		_w10273_
	);
	LUT3 #(
		.INIT('h80)
	) name8924 (
		_w1804_,
		_w1826_,
		_w10273_,
		_w10274_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8925 (
		_w1933_,
		_w10272_,
		_w10270_,
		_w10274_,
		_w10275_
	);
	LUT3 #(
		.INIT('hf2)
	) name8926 (
		\P1_EAX_reg[8]/NET0131 ,
		_w10016_,
		_w10275_,
		_w10276_
	);
	LUT2 #(
		.INIT('h2)
	) name8927 (
		\P2_EAX_reg[10]/NET0131 ,
		_w7767_,
		_w10277_
	);
	LUT2 #(
		.INIT('h4)
	) name8928 (
		_w7772_,
		_w7789_,
		_w10278_
	);
	LUT4 #(
		.INIT('h153f)
	) name8929 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[3][2]/NET0131 ,
		_w1462_,
		_w1465_,
		_w10279_
	);
	LUT4 #(
		.INIT('h153f)
	) name8930 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[1][2]/NET0131 ,
		_w1453_,
		_w1447_,
		_w10280_
	);
	LUT4 #(
		.INIT('h153f)
	) name8931 (
		\P2_InstQueue_reg[2][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1450_,
		_w1446_,
		_w10281_
	);
	LUT4 #(
		.INIT('h135f)
	) name8932 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1443_,
		_w1466_,
		_w10282_
	);
	LUT4 #(
		.INIT('h8000)
	) name8933 (
		_w10281_,
		_w10282_,
		_w10279_,
		_w10280_,
		_w10283_
	);
	LUT4 #(
		.INIT('h153f)
	) name8934 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10284_
	);
	LUT4 #(
		.INIT('h135f)
	) name8935 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1452_,
		_w1456_,
		_w10285_
	);
	LUT4 #(
		.INIT('h153f)
	) name8936 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1449_,
		_w1457_,
		_w10286_
	);
	LUT4 #(
		.INIT('h153f)
	) name8937 (
		\P2_InstQueue_reg[13][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1444_,
		_w1459_,
		_w10287_
	);
	LUT4 #(
		.INIT('h8000)
	) name8938 (
		_w10286_,
		_w10287_,
		_w10284_,
		_w10285_,
		_w10288_
	);
	LUT4 #(
		.INIT('h0111)
	) name8939 (
		_w1592_,
		_w1595_,
		_w10283_,
		_w10288_,
		_w10289_
	);
	LUT3 #(
		.INIT('h80)
	) name8940 (
		_w1549_,
		_w1553_,
		_w10289_,
		_w10290_
	);
	LUT3 #(
		.INIT('h40)
	) name8941 (
		\P2_EAX_reg[10]/NET0131 ,
		_w7771_,
		_w7789_,
		_w10291_
	);
	LUT4 #(
		.INIT('h0007)
	) name8942 (
		_w1656_,
		_w9522_,
		_w10290_,
		_w10291_,
		_w10292_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8943 (
		\P2_EAX_reg[10]/NET0131 ,
		_w7792_,
		_w10278_,
		_w10292_,
		_w10293_
	);
	LUT3 #(
		.INIT('hce)
	) name8944 (
		_w1678_,
		_w10277_,
		_w10293_,
		_w10294_
	);
	LUT2 #(
		.INIT('h2)
	) name8945 (
		\P2_EAX_reg[11]/NET0131 ,
		_w7767_,
		_w10295_
	);
	LUT4 #(
		.INIT('h153f)
	) name8946 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[3][3]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10296_
	);
	LUT4 #(
		.INIT('h153f)
	) name8947 (
		\P2_InstQueue_reg[13][3]/NET0131 ,
		\P2_InstQueue_reg[1][3]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10297_
	);
	LUT4 #(
		.INIT('h153f)
	) name8948 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1450_,
		_w1465_,
		_w10298_
	);
	LUT4 #(
		.INIT('h153f)
	) name8949 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10299_
	);
	LUT4 #(
		.INIT('h8000)
	) name8950 (
		_w10298_,
		_w10299_,
		_w10296_,
		_w10297_,
		_w10300_
	);
	LUT4 #(
		.INIT('h135f)
	) name8951 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1443_,
		_w1446_,
		_w10301_
	);
	LUT4 #(
		.INIT('h153f)
	) name8952 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10302_
	);
	LUT4 #(
		.INIT('h135f)
	) name8953 (
		\P2_InstQueue_reg[6][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1466_,
		_w1456_,
		_w10303_
	);
	LUT4 #(
		.INIT('h153f)
	) name8954 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1444_,
		_w1447_,
		_w10304_
	);
	LUT4 #(
		.INIT('h8000)
	) name8955 (
		_w10303_,
		_w10304_,
		_w10301_,
		_w10302_,
		_w10305_
	);
	LUT4 #(
		.INIT('h0111)
	) name8956 (
		_w1592_,
		_w1595_,
		_w10300_,
		_w10305_,
		_w10306_
	);
	LUT3 #(
		.INIT('h80)
	) name8957 (
		_w1549_,
		_w1553_,
		_w10306_,
		_w10307_
	);
	LUT3 #(
		.INIT('h20)
	) name8958 (
		\P2_EAX_reg[10]/NET0131 ,
		\P2_EAX_reg[11]/NET0131 ,
		_w7771_,
		_w10308_
	);
	LUT2 #(
		.INIT('h8)
	) name8959 (
		_w7789_,
		_w10308_,
		_w10309_
	);
	LUT4 #(
		.INIT('h000b)
	) name8960 (
		_w8452_,
		_w8812_,
		_w10307_,
		_w10309_,
		_w10310_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8961 (
		\P2_EAX_reg[11]/NET0131 ,
		_w7792_,
		_w10278_,
		_w10310_,
		_w10311_
	);
	LUT3 #(
		.INIT('hce)
	) name8962 (
		_w1678_,
		_w10295_,
		_w10311_,
		_w10312_
	);
	LUT2 #(
		.INIT('h2)
	) name8963 (
		\P2_EAX_reg[12]/NET0131 ,
		_w7767_,
		_w10313_
	);
	LUT2 #(
		.INIT('h4)
	) name8964 (
		_w7774_,
		_w7789_,
		_w10314_
	);
	LUT3 #(
		.INIT('h40)
	) name8965 (
		\P2_EAX_reg[12]/NET0131 ,
		_w7773_,
		_w7789_,
		_w10315_
	);
	LUT4 #(
		.INIT('h153f)
	) name8966 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[3][4]/NET0131 ,
		_w1462_,
		_w1465_,
		_w10316_
	);
	LUT4 #(
		.INIT('h153f)
	) name8967 (
		\P2_InstQueue_reg[14][4]/NET0131 ,
		\P2_InstQueue_reg[1][4]/NET0131 ,
		_w1453_,
		_w1447_,
		_w10317_
	);
	LUT4 #(
		.INIT('h153f)
	) name8968 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1450_,
		_w1446_,
		_w10318_
	);
	LUT4 #(
		.INIT('h135f)
	) name8969 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1443_,
		_w1466_,
		_w10319_
	);
	LUT4 #(
		.INIT('h8000)
	) name8970 (
		_w10318_,
		_w10319_,
		_w10316_,
		_w10317_,
		_w10320_
	);
	LUT4 #(
		.INIT('h153f)
	) name8971 (
		\P2_InstQueue_reg[15][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10321_
	);
	LUT4 #(
		.INIT('h135f)
	) name8972 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1452_,
		_w1456_,
		_w10322_
	);
	LUT4 #(
		.INIT('h153f)
	) name8973 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1449_,
		_w1457_,
		_w10323_
	);
	LUT4 #(
		.INIT('h153f)
	) name8974 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1444_,
		_w1459_,
		_w10324_
	);
	LUT4 #(
		.INIT('h8000)
	) name8975 (
		_w10323_,
		_w10324_,
		_w10321_,
		_w10322_,
		_w10325_
	);
	LUT4 #(
		.INIT('h0111)
	) name8976 (
		_w1592_,
		_w1595_,
		_w10320_,
		_w10325_,
		_w10326_
	);
	LUT3 #(
		.INIT('h80)
	) name8977 (
		_w1549_,
		_w1553_,
		_w10326_,
		_w10327_
	);
	LUT4 #(
		.INIT('h0007)
	) name8978 (
		_w1656_,
		_w9451_,
		_w10315_,
		_w10327_,
		_w10328_
	);
	LUT4 #(
		.INIT('h5d00)
	) name8979 (
		\P2_EAX_reg[12]/NET0131 ,
		_w7792_,
		_w10314_,
		_w10328_,
		_w10329_
	);
	LUT3 #(
		.INIT('hce)
	) name8980 (
		_w1678_,
		_w10313_,
		_w10329_,
		_w10330_
	);
	LUT3 #(
		.INIT('h02)
	) name8981 (
		_w1855_,
		_w1861_,
		_w3474_,
		_w10331_
	);
	LUT4 #(
		.INIT('h0111)
	) name8982 (
		_w1842_,
		_w1845_,
		_w3121_,
		_w3126_,
		_w10332_
	);
	LUT4 #(
		.INIT('h4000)
	) name8983 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10332_,
		_w10333_
	);
	LUT4 #(
		.INIT('h78f0)
	) name8984 (
		\P1_EAX_reg[4]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w9418_,
		_w10334_
	);
	LUT3 #(
		.INIT('h80)
	) name8985 (
		_w1804_,
		_w1826_,
		_w10334_,
		_w10335_
	);
	LUT2 #(
		.INIT('h1)
	) name8986 (
		_w10333_,
		_w10335_,
		_w10336_
	);
	LUT3 #(
		.INIT('h8a)
	) name8987 (
		_w1933_,
		_w10331_,
		_w10336_,
		_w10337_
	);
	LUT3 #(
		.INIT('hf2)
	) name8988 (
		\P1_EAX_reg[6]/NET0131 ,
		_w10016_,
		_w10337_,
		_w10338_
	);
	LUT3 #(
		.INIT('h02)
	) name8989 (
		_w1855_,
		_w1861_,
		_w3445_,
		_w10339_
	);
	LUT4 #(
		.INIT('h153f)
	) name8990 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1691_,
		_w1703_,
		_w10340_
	);
	LUT4 #(
		.INIT('h153f)
	) name8991 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[5][1]/NET0131 ,
		_w1702_,
		_w1705_,
		_w10341_
	);
	LUT4 #(
		.INIT('h135f)
	) name8992 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1696_,
		_w1706_,
		_w10342_
	);
	LUT4 #(
		.INIT('h135f)
	) name8993 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1694_,
		_w1692_,
		_w10343_
	);
	LUT4 #(
		.INIT('h8000)
	) name8994 (
		_w10342_,
		_w10343_,
		_w10340_,
		_w10341_,
		_w10344_
	);
	LUT4 #(
		.INIT('h135f)
	) name8995 (
		\P1_InstQueue_reg[14][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1698_,
		_w1689_,
		_w10345_
	);
	LUT4 #(
		.INIT('h153f)
	) name8996 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1711_,
		_w1712_,
		_w10346_
	);
	LUT4 #(
		.INIT('h135f)
	) name8997 (
		\P1_InstQueue_reg[2][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1688_,
		_w1708_,
		_w10347_
	);
	LUT4 #(
		.INIT('h135f)
	) name8998 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[4][1]/NET0131 ,
		_w1699_,
		_w1709_,
		_w10348_
	);
	LUT4 #(
		.INIT('h8000)
	) name8999 (
		_w10347_,
		_w10348_,
		_w10345_,
		_w10346_,
		_w10349_
	);
	LUT4 #(
		.INIT('h0111)
	) name9000 (
		_w1842_,
		_w1845_,
		_w10344_,
		_w10349_,
		_w10350_
	);
	LUT4 #(
		.INIT('h4000)
	) name9001 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10350_,
		_w10351_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9002 (
		\P1_EAX_reg[7]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w9419_,
		_w10352_
	);
	LUT3 #(
		.INIT('h80)
	) name9003 (
		_w1804_,
		_w1826_,
		_w10352_,
		_w10353_
	);
	LUT2 #(
		.INIT('h1)
	) name9004 (
		_w10351_,
		_w10353_,
		_w10354_
	);
	LUT3 #(
		.INIT('h8a)
	) name9005 (
		_w1933_,
		_w10339_,
		_w10354_,
		_w10355_
	);
	LUT3 #(
		.INIT('hf2)
	) name9006 (
		\P1_EAX_reg[9]/NET0131 ,
		_w10016_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h2)
	) name9007 (
		\P2_EAX_reg[13]/NET0131 ,
		_w7767_,
		_w10357_
	);
	LUT3 #(
		.INIT('h40)
	) name9008 (
		\P2_EAX_reg[13]/NET0131 ,
		_w7774_,
		_w7789_,
		_w10358_
	);
	LUT2 #(
		.INIT('h2)
	) name9009 (
		_w1606_,
		_w9702_,
		_w10359_
	);
	LUT4 #(
		.INIT('hec00)
	) name9010 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w10359_,
		_w10360_
	);
	LUT4 #(
		.INIT('h153f)
	) name9011 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10361_
	);
	LUT4 #(
		.INIT('h153f)
	) name9012 (
		\P2_InstQueue_reg[13][5]/NET0131 ,
		\P2_InstQueue_reg[1][5]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10362_
	);
	LUT4 #(
		.INIT('h153f)
	) name9013 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[5][5]/NET0131 ,
		_w1450_,
		_w1465_,
		_w10363_
	);
	LUT4 #(
		.INIT('h153f)
	) name9014 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10364_
	);
	LUT4 #(
		.INIT('h8000)
	) name9015 (
		_w10363_,
		_w10364_,
		_w10361_,
		_w10362_,
		_w10365_
	);
	LUT4 #(
		.INIT('h135f)
	) name9016 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1443_,
		_w1446_,
		_w10366_
	);
	LUT4 #(
		.INIT('h153f)
	) name9017 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10367_
	);
	LUT4 #(
		.INIT('h135f)
	) name9018 (
		\P2_InstQueue_reg[6][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1466_,
		_w1456_,
		_w10368_
	);
	LUT4 #(
		.INIT('h153f)
	) name9019 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1444_,
		_w1447_,
		_w10369_
	);
	LUT4 #(
		.INIT('h8000)
	) name9020 (
		_w10368_,
		_w10369_,
		_w10366_,
		_w10367_,
		_w10370_
	);
	LUT4 #(
		.INIT('h0111)
	) name9021 (
		_w1592_,
		_w1595_,
		_w10365_,
		_w10370_,
		_w10371_
	);
	LUT3 #(
		.INIT('h80)
	) name9022 (
		_w1549_,
		_w1553_,
		_w10371_,
		_w10372_
	);
	LUT3 #(
		.INIT('h01)
	) name9023 (
		_w10360_,
		_w10372_,
		_w10358_,
		_w10373_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9024 (
		\P2_EAX_reg[13]/NET0131 ,
		_w7792_,
		_w10314_,
		_w10373_,
		_w10374_
	);
	LUT3 #(
		.INIT('hce)
	) name9025 (
		_w1678_,
		_w10357_,
		_w10374_,
		_w10375_
	);
	LUT2 #(
		.INIT('h2)
	) name9026 (
		\P2_EAX_reg[14]/NET0131 ,
		_w7767_,
		_w10376_
	);
	LUT2 #(
		.INIT('h4)
	) name9027 (
		_w7775_,
		_w7789_,
		_w10377_
	);
	LUT3 #(
		.INIT('h40)
	) name9028 (
		\P2_EAX_reg[14]/NET0131 ,
		_w7775_,
		_w7789_,
		_w10378_
	);
	LUT4 #(
		.INIT('hec00)
	) name9029 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w8938_,
		_w10379_
	);
	LUT4 #(
		.INIT('h153f)
	) name9030 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10380_
	);
	LUT4 #(
		.INIT('h153f)
	) name9031 (
		\P2_InstQueue_reg[13][6]/NET0131 ,
		\P2_InstQueue_reg[1][6]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10381_
	);
	LUT4 #(
		.INIT('h153f)
	) name9032 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1450_,
		_w1465_,
		_w10382_
	);
	LUT4 #(
		.INIT('h153f)
	) name9033 (
		\P2_InstQueue_reg[15][6]/NET0131 ,
		\P2_InstQueue_reg[4][6]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10383_
	);
	LUT4 #(
		.INIT('h8000)
	) name9034 (
		_w10382_,
		_w10383_,
		_w10380_,
		_w10381_,
		_w10384_
	);
	LUT4 #(
		.INIT('h135f)
	) name9035 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[2][6]/NET0131 ,
		_w1443_,
		_w1446_,
		_w10385_
	);
	LUT4 #(
		.INIT('h153f)
	) name9036 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10386_
	);
	LUT4 #(
		.INIT('h135f)
	) name9037 (
		\P2_InstQueue_reg[6][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1466_,
		_w1456_,
		_w10387_
	);
	LUT4 #(
		.INIT('h153f)
	) name9038 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1444_,
		_w1447_,
		_w10388_
	);
	LUT4 #(
		.INIT('h8000)
	) name9039 (
		_w10387_,
		_w10388_,
		_w10385_,
		_w10386_,
		_w10389_
	);
	LUT4 #(
		.INIT('h0111)
	) name9040 (
		_w1592_,
		_w1595_,
		_w10384_,
		_w10389_,
		_w10390_
	);
	LUT3 #(
		.INIT('h80)
	) name9041 (
		_w1549_,
		_w1553_,
		_w10390_,
		_w10391_
	);
	LUT3 #(
		.INIT('h01)
	) name9042 (
		_w10379_,
		_w10391_,
		_w10378_,
		_w10392_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9043 (
		\P2_EAX_reg[14]/NET0131 ,
		_w7792_,
		_w10377_,
		_w10392_,
		_w10393_
	);
	LUT3 #(
		.INIT('hce)
	) name9044 (
		_w1678_,
		_w10376_,
		_w10393_,
		_w10394_
	);
	LUT2 #(
		.INIT('h2)
	) name9045 (
		\P2_EAX_reg[1]/NET0131 ,
		_w7767_,
		_w10395_
	);
	LUT2 #(
		.INIT('h2)
	) name9046 (
		_w1606_,
		_w7156_,
		_w10396_
	);
	LUT4 #(
		.INIT('hec00)
	) name9047 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w10396_,
		_w10397_
	);
	LUT4 #(
		.INIT('h0111)
	) name9048 (
		_w1592_,
		_w1595_,
		_w4121_,
		_w4126_,
		_w10398_
	);
	LUT3 #(
		.INIT('h80)
	) name9049 (
		_w1549_,
		_w1553_,
		_w10398_,
		_w10399_
	);
	LUT2 #(
		.INIT('h2)
	) name9050 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		_w10400_
	);
	LUT2 #(
		.INIT('h8)
	) name9051 (
		_w7789_,
		_w10400_,
		_w10401_
	);
	LUT3 #(
		.INIT('h01)
	) name9052 (
		_w10397_,
		_w10399_,
		_w10401_,
		_w10402_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9053 (
		\P2_EAX_reg[1]/NET0131 ,
		_w7792_,
		_w10247_,
		_w10402_,
		_w10403_
	);
	LUT3 #(
		.INIT('hce)
	) name9054 (
		_w1678_,
		_w10395_,
		_w10403_,
		_w10404_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9055 (
		\P2_EAX_reg[2]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10405_
	);
	LUT4 #(
		.INIT('h0111)
	) name9056 (
		_w1592_,
		_w1595_,
		_w4109_,
		_w4114_,
		_w10406_
	);
	LUT3 #(
		.INIT('h80)
	) name9057 (
		_w1549_,
		_w1553_,
		_w10406_,
		_w10407_
	);
	LUT3 #(
		.INIT('h78)
	) name9058 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		_w10408_
	);
	LUT2 #(
		.INIT('h8)
	) name9059 (
		_w7789_,
		_w10408_,
		_w10409_
	);
	LUT4 #(
		.INIT('h000b)
	) name9060 (
		_w5487_,
		_w8812_,
		_w10407_,
		_w10409_,
		_w10410_
	);
	LUT2 #(
		.INIT('h2)
	) name9061 (
		_w1678_,
		_w10410_,
		_w10411_
	);
	LUT2 #(
		.INIT('he)
	) name9062 (
		_w10405_,
		_w10411_,
		_w10412_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9063 (
		\P2_EAX_reg[3]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10413_
	);
	LUT4 #(
		.INIT('h0111)
	) name9064 (
		_w1592_,
		_w1595_,
		_w4160_,
		_w4165_,
		_w10414_
	);
	LUT3 #(
		.INIT('h80)
	) name9065 (
		_w1549_,
		_w1553_,
		_w10414_,
		_w10415_
	);
	LUT4 #(
		.INIT('h7f80)
	) name9066 (
		\P2_EAX_reg[0]/NET0131 ,
		\P2_EAX_reg[1]/NET0131 ,
		\P2_EAX_reg[2]/NET0131 ,
		\P2_EAX_reg[3]/NET0131 ,
		_w10416_
	);
	LUT2 #(
		.INIT('h8)
	) name9067 (
		_w7789_,
		_w10416_,
		_w10417_
	);
	LUT4 #(
		.INIT('h000b)
	) name9068 (
		_w3561_,
		_w8812_,
		_w10415_,
		_w10417_,
		_w10418_
	);
	LUT2 #(
		.INIT('h2)
	) name9069 (
		_w1678_,
		_w10418_,
		_w10419_
	);
	LUT2 #(
		.INIT('he)
	) name9070 (
		_w10413_,
		_w10419_,
		_w10420_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9071 (
		\P2_EAX_reg[4]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10421_
	);
	LUT4 #(
		.INIT('h0111)
	) name9072 (
		_w1592_,
		_w1595_,
		_w4147_,
		_w4152_,
		_w10422_
	);
	LUT3 #(
		.INIT('h80)
	) name9073 (
		_w1549_,
		_w1553_,
		_w10422_,
		_w10423_
	);
	LUT2 #(
		.INIT('h6)
	) name9074 (
		\P2_EAX_reg[4]/NET0131 ,
		_w7769_,
		_w10424_
	);
	LUT2 #(
		.INIT('h8)
	) name9075 (
		_w7789_,
		_w10424_,
		_w10425_
	);
	LUT4 #(
		.INIT('h000b)
	) name9076 (
		_w2276_,
		_w8812_,
		_w10423_,
		_w10425_,
		_w10426_
	);
	LUT2 #(
		.INIT('h2)
	) name9077 (
		_w1678_,
		_w10426_,
		_w10427_
	);
	LUT2 #(
		.INIT('he)
	) name9078 (
		_w10421_,
		_w10427_,
		_w10428_
	);
	LUT4 #(
		.INIT('h135f)
	) name9079 (
		\P1_InstQueue_reg[2][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1688_,
		_w1691_,
		_w10429_
	);
	LUT4 #(
		.INIT('h135f)
	) name9080 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w1712_,
		_w1705_,
		_w10430_
	);
	LUT4 #(
		.INIT('h135f)
	) name9081 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w1696_,
		_w1706_,
		_w10431_
	);
	LUT4 #(
		.INIT('h135f)
	) name9082 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1698_,
		_w1692_,
		_w10432_
	);
	LUT4 #(
		.INIT('h8000)
	) name9083 (
		_w10431_,
		_w10432_,
		_w10429_,
		_w10430_,
		_w10433_
	);
	LUT4 #(
		.INIT('h135f)
	) name9084 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1709_,
		_w1711_,
		_w10434_
	);
	LUT4 #(
		.INIT('h153f)
	) name9085 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1689_,
		_w1703_,
		_w10435_
	);
	LUT4 #(
		.INIT('h135f)
	) name9086 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[5][2]/NET0131 ,
		_w1694_,
		_w1702_,
		_w10436_
	);
	LUT4 #(
		.INIT('h135f)
	) name9087 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1699_,
		_w1708_,
		_w10437_
	);
	LUT4 #(
		.INIT('h8000)
	) name9088 (
		_w10436_,
		_w10437_,
		_w10434_,
		_w10435_,
		_w10438_
	);
	LUT4 #(
		.INIT('h0111)
	) name9089 (
		_w1842_,
		_w1845_,
		_w10433_,
		_w10438_,
		_w10439_
	);
	LUT4 #(
		.INIT('h4000)
	) name9090 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10439_,
		_w10440_
	);
	LUT2 #(
		.INIT('h2)
	) name9091 (
		_w1867_,
		_w3449_,
		_w10441_
	);
	LUT4 #(
		.INIT('hec00)
	) name9092 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10441_,
		_w10442_
	);
	LUT2 #(
		.INIT('h6)
	) name9093 (
		\P1_EAX_reg[10]/NET0131 ,
		_w9420_,
		_w10443_
	);
	LUT3 #(
		.INIT('h80)
	) name9094 (
		_w1804_,
		_w1826_,
		_w10443_,
		_w10444_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9095 (
		_w1933_,
		_w10442_,
		_w10440_,
		_w10444_,
		_w10445_
	);
	LUT3 #(
		.INIT('hf2)
	) name9096 (
		\P1_EAX_reg[10]/NET0131 ,
		_w10016_,
		_w10445_,
		_w10446_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9097 (
		\P2_EAX_reg[5]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10447_
	);
	LUT4 #(
		.INIT('h0111)
	) name9098 (
		_w1592_,
		_w1595_,
		_w4192_,
		_w4197_,
		_w10448_
	);
	LUT3 #(
		.INIT('h80)
	) name9099 (
		_w1549_,
		_w1553_,
		_w10448_,
		_w10449_
	);
	LUT3 #(
		.INIT('h6c)
	) name9100 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		_w7769_,
		_w10450_
	);
	LUT2 #(
		.INIT('h8)
	) name9101 (
		_w7789_,
		_w10450_,
		_w10451_
	);
	LUT4 #(
		.INIT('h000b)
	) name9102 (
		_w6502_,
		_w8812_,
		_w10449_,
		_w10451_,
		_w10452_
	);
	LUT2 #(
		.INIT('h2)
	) name9103 (
		_w1678_,
		_w10452_,
		_w10453_
	);
	LUT2 #(
		.INIT('he)
	) name9104 (
		_w10447_,
		_w10453_,
		_w10454_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9105 (
		\P2_EAX_reg[6]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10455_
	);
	LUT4 #(
		.INIT('h0111)
	) name9106 (
		_w1592_,
		_w1595_,
		_w4178_,
		_w4183_,
		_w10456_
	);
	LUT3 #(
		.INIT('h80)
	) name9107 (
		_w1549_,
		_w1553_,
		_w10456_,
		_w10457_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9108 (
		\P2_EAX_reg[4]/NET0131 ,
		\P2_EAX_reg[5]/NET0131 ,
		\P2_EAX_reg[6]/NET0131 ,
		_w7769_,
		_w10458_
	);
	LUT2 #(
		.INIT('h8)
	) name9109 (
		_w7789_,
		_w10458_,
		_w10459_
	);
	LUT4 #(
		.INIT('h000b)
	) name9110 (
		_w4977_,
		_w8812_,
		_w10457_,
		_w10459_,
		_w10460_
	);
	LUT2 #(
		.INIT('h2)
	) name9111 (
		_w1678_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('he)
	) name9112 (
		_w10455_,
		_w10461_,
		_w10462_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9113 (
		\P2_EAX_reg[8]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10463_
	);
	LUT4 #(
		.INIT('h153f)
	) name9114 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1462_,
		_w1457_,
		_w10464_
	);
	LUT4 #(
		.INIT('h153f)
	) name9115 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[1][0]/NET0131 ,
		_w1453_,
		_w1459_,
		_w10465_
	);
	LUT4 #(
		.INIT('h153f)
	) name9116 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1450_,
		_w1465_,
		_w10466_
	);
	LUT4 #(
		.INIT('h153f)
	) name9117 (
		\P2_InstQueue_reg[15][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10467_
	);
	LUT4 #(
		.INIT('h8000)
	) name9118 (
		_w10466_,
		_w10467_,
		_w10464_,
		_w10465_,
		_w10468_
	);
	LUT4 #(
		.INIT('h135f)
	) name9119 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[2][0]/NET0131 ,
		_w1443_,
		_w1446_,
		_w10469_
	);
	LUT4 #(
		.INIT('h153f)
	) name9120 (
		\P2_InstQueue_reg[11][0]/NET0131 ,
		\P2_InstQueue_reg[7][0]/NET0131 ,
		_w1449_,
		_w1452_,
		_w10470_
	);
	LUT4 #(
		.INIT('h135f)
	) name9121 (
		\P2_InstQueue_reg[6][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1466_,
		_w1456_,
		_w10471_
	);
	LUT4 #(
		.INIT('h153f)
	) name9122 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1444_,
		_w1447_,
		_w10472_
	);
	LUT4 #(
		.INIT('h8000)
	) name9123 (
		_w10471_,
		_w10472_,
		_w10469_,
		_w10470_,
		_w10473_
	);
	LUT4 #(
		.INIT('h0111)
	) name9124 (
		_w1592_,
		_w1595_,
		_w10468_,
		_w10473_,
		_w10474_
	);
	LUT3 #(
		.INIT('h80)
	) name9125 (
		_w1549_,
		_w1553_,
		_w10474_,
		_w10475_
	);
	LUT3 #(
		.INIT('h6c)
	) name9126 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		_w7770_,
		_w10476_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		_w7789_,
		_w10476_,
		_w10477_
	);
	LUT4 #(
		.INIT('h0007)
	) name9128 (
		_w1656_,
		_w10006_,
		_w10475_,
		_w10477_,
		_w10478_
	);
	LUT2 #(
		.INIT('h2)
	) name9129 (
		_w1678_,
		_w10478_,
		_w10479_
	);
	LUT2 #(
		.INIT('he)
	) name9130 (
		_w10463_,
		_w10479_,
		_w10480_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9131 (
		\P2_EAX_reg[9]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w10481_
	);
	LUT4 #(
		.INIT('h3111)
	) name9132 (
		\P2_Address_reg[29]/NET0131 ,
		\buf2_reg[9]/NET0131 ,
		_w2255_,
		_w2260_,
		_w10482_
	);
	LUT4 #(
		.INIT('h0222)
	) name9133 (
		\P2_Address_reg[29]/NET0131 ,
		\buf1_reg[9]/NET0131 ,
		_w2255_,
		_w2260_,
		_w10483_
	);
	LUT2 #(
		.INIT('h1)
	) name9134 (
		_w10482_,
		_w10483_,
		_w10484_
	);
	LUT2 #(
		.INIT('h8)
	) name9135 (
		_w1606_,
		_w10484_,
		_w10485_
	);
	LUT4 #(
		.INIT('hec00)
	) name9136 (
		_w1501_,
		_w1565_,
		_w1568_,
		_w10485_,
		_w10486_
	);
	LUT4 #(
		.INIT('h153f)
	) name9137 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1462_,
		_w1465_,
		_w10487_
	);
	LUT4 #(
		.INIT('h153f)
	) name9138 (
		\P2_InstQueue_reg[14][1]/NET0131 ,
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1453_,
		_w1447_,
		_w10488_
	);
	LUT4 #(
		.INIT('h153f)
	) name9139 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1450_,
		_w1446_,
		_w10489_
	);
	LUT4 #(
		.INIT('h135f)
	) name9140 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1443_,
		_w1466_,
		_w10490_
	);
	LUT4 #(
		.INIT('h8000)
	) name9141 (
		_w10489_,
		_w10490_,
		_w10487_,
		_w10488_,
		_w10491_
	);
	LUT4 #(
		.INIT('h153f)
	) name9142 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1463_,
		_w1460_,
		_w10492_
	);
	LUT4 #(
		.INIT('h135f)
	) name9143 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1452_,
		_w1456_,
		_w10493_
	);
	LUT4 #(
		.INIT('h153f)
	) name9144 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[7][1]/NET0131 ,
		_w1449_,
		_w1457_,
		_w10494_
	);
	LUT4 #(
		.INIT('h153f)
	) name9145 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1444_,
		_w1459_,
		_w10495_
	);
	LUT4 #(
		.INIT('h8000)
	) name9146 (
		_w10494_,
		_w10495_,
		_w10492_,
		_w10493_,
		_w10496_
	);
	LUT4 #(
		.INIT('h0111)
	) name9147 (
		_w1592_,
		_w1595_,
		_w10491_,
		_w10496_,
		_w10497_
	);
	LUT3 #(
		.INIT('h80)
	) name9148 (
		_w1549_,
		_w1553_,
		_w10497_,
		_w10498_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9149 (
		\P2_EAX_reg[7]/NET0131 ,
		\P2_EAX_reg[8]/NET0131 ,
		\P2_EAX_reg[9]/NET0131 ,
		_w7770_,
		_w10499_
	);
	LUT2 #(
		.INIT('h8)
	) name9150 (
		_w7789_,
		_w10499_,
		_w10500_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9151 (
		_w1678_,
		_w10486_,
		_w10498_,
		_w10500_,
		_w10501_
	);
	LUT2 #(
		.INIT('he)
	) name9152 (
		_w10481_,
		_w10501_,
		_w10502_
	);
	LUT2 #(
		.INIT('h2)
	) name9153 (
		\P1_EAX_reg[11]/NET0131 ,
		_w9102_,
		_w10503_
	);
	LUT3 #(
		.INIT('h08)
	) name9154 (
		_w1804_,
		_w1826_,
		_w9422_,
		_w10504_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9155 (
		\P1_EAX_reg[11]/NET0131 ,
		_w9436_,
		_w9437_,
		_w10504_,
		_w10505_
	);
	LUT4 #(
		.INIT('h4000)
	) name9156 (
		\P1_EAX_reg[11]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9421_,
		_w10506_
	);
	LUT2 #(
		.INIT('h2)
	) name9157 (
		_w1867_,
		_w3431_,
		_w10507_
	);
	LUT4 #(
		.INIT('hec00)
	) name9158 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10507_,
		_w10508_
	);
	LUT4 #(
		.INIT('h135f)
	) name9159 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1688_,
		_w1689_,
		_w10509_
	);
	LUT4 #(
		.INIT('h153f)
	) name9160 (
		\P1_InstQueue_reg[15][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1708_,
		_w1705_,
		_w10510_
	);
	LUT4 #(
		.INIT('h153f)
	) name9161 (
		\P1_InstQueue_reg[1][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1692_,
		_w1706_,
		_w10511_
	);
	LUT4 #(
		.INIT('h135f)
	) name9162 (
		\P1_InstQueue_reg[13][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1696_,
		_w1709_,
		_w10512_
	);
	LUT4 #(
		.INIT('h8000)
	) name9163 (
		_w10511_,
		_w10512_,
		_w10509_,
		_w10510_,
		_w10513_
	);
	LUT4 #(
		.INIT('h135f)
	) name9164 (
		\P1_InstQueue_reg[7][3]/NET0131 ,
		\P1_InstQueue_reg[8][3]/NET0131 ,
		_w1691_,
		_w1711_,
		_w10514_
	);
	LUT4 #(
		.INIT('h135f)
	) name9165 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[11][3]/NET0131 ,
		_w1712_,
		_w1703_,
		_w10515_
	);
	LUT4 #(
		.INIT('h135f)
	) name9166 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[5][3]/NET0131 ,
		_w1698_,
		_w1702_,
		_w10516_
	);
	LUT4 #(
		.INIT('h153f)
	) name9167 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[12][3]/NET0131 ,
		_w1694_,
		_w1699_,
		_w10517_
	);
	LUT4 #(
		.INIT('h8000)
	) name9168 (
		_w10516_,
		_w10517_,
		_w10514_,
		_w10515_,
		_w10518_
	);
	LUT4 #(
		.INIT('h0111)
	) name9169 (
		_w1842_,
		_w1845_,
		_w10513_,
		_w10518_,
		_w10519_
	);
	LUT4 #(
		.INIT('h4000)
	) name9170 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10519_,
		_w10520_
	);
	LUT3 #(
		.INIT('h01)
	) name9171 (
		_w10508_,
		_w10520_,
		_w10506_,
		_w10521_
	);
	LUT4 #(
		.INIT('hecee)
	) name9172 (
		_w1933_,
		_w10503_,
		_w10505_,
		_w10521_,
		_w10522_
	);
	LUT4 #(
		.INIT('h8000)
	) name9173 (
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w8987_,
		_w8989_,
		_w10523_
	);
	LUT3 #(
		.INIT('ha8)
	) name9174 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1863_,
		_w8992_,
		_w10524_
	);
	LUT4 #(
		.INIT('h8008)
	) name9175 (
		_w1814_,
		_w1846_,
		_w9073_,
		_w9084_,
		_w10525_
	);
	LUT2 #(
		.INIT('h1)
	) name9176 (
		_w10524_,
		_w10525_,
		_w10526_
	);
	LUT4 #(
		.INIT('hb700)
	) name9177 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1829_,
		_w10523_,
		_w10526_,
		_w10527_
	);
	LUT2 #(
		.INIT('h2)
	) name9178 (
		\P1_EBX_reg[29]/NET0131 ,
		_w9102_,
		_w10528_
	);
	LUT3 #(
		.INIT('hf2)
	) name9179 (
		_w1933_,
		_w10527_,
		_w10528_,
		_w10529_
	);
	LUT4 #(
		.INIT('h60c0)
	) name9180 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w1578_,
		_w8960_,
		_w10530_
	);
	LUT4 #(
		.INIT('h8008)
	) name9181 (
		_w1550_,
		_w1596_,
		_w7873_,
		_w7884_,
		_w10531_
	);
	LUT2 #(
		.INIT('h2)
	) name9182 (
		\P2_EBX_reg[29]/NET0131 ,
		_w8961_,
		_w10532_
	);
	LUT2 #(
		.INIT('h1)
	) name9183 (
		_w10531_,
		_w10532_,
		_w10533_
	);
	LUT2 #(
		.INIT('h2)
	) name9184 (
		\P2_EBX_reg[29]/NET0131 ,
		_w7767_,
		_w10534_
	);
	LUT4 #(
		.INIT('hff8a)
	) name9185 (
		_w1678_,
		_w10530_,
		_w10533_,
		_w10534_,
		_w10535_
	);
	LUT2 #(
		.INIT('h2)
	) name9186 (
		\P1_EAX_reg[14]/NET0131 ,
		_w9102_,
		_w10536_
	);
	LUT3 #(
		.INIT('h08)
	) name9187 (
		_w1804_,
		_w1826_,
		_w9424_,
		_w10537_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9188 (
		\P1_EAX_reg[14]/NET0131 ,
		_w9436_,
		_w9437_,
		_w10537_,
		_w10538_
	);
	LUT3 #(
		.INIT('h02)
	) name9189 (
		_w1855_,
		_w1861_,
		_w3457_,
		_w10539_
	);
	LUT4 #(
		.INIT('h4000)
	) name9190 (
		\P1_EAX_reg[14]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9424_,
		_w10540_
	);
	LUT4 #(
		.INIT('h135f)
	) name9191 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1688_,
		_w1691_,
		_w10541_
	);
	LUT4 #(
		.INIT('h153f)
	) name9192 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1711_,
		_w1705_,
		_w10542_
	);
	LUT4 #(
		.INIT('h153f)
	) name9193 (
		\P1_InstQueue_reg[1][6]/NET0131 ,
		\P1_InstQueue_reg[3][6]/NET0131 ,
		_w1692_,
		_w1706_,
		_w10543_
	);
	LUT4 #(
		.INIT('h135f)
	) name9194 (
		\P1_InstQueue_reg[12][6]/NET0131 ,
		\P1_InstQueue_reg[13][6]/NET0131 ,
		_w1694_,
		_w1696_,
		_w10544_
	);
	LUT4 #(
		.INIT('h8000)
	) name9195 (
		_w10543_,
		_w10544_,
		_w10541_,
		_w10542_,
		_w10545_
	);
	LUT4 #(
		.INIT('h135f)
	) name9196 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1698_,
		_w1689_,
		_w10546_
	);
	LUT4 #(
		.INIT('h135f)
	) name9197 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[11][6]/NET0131 ,
		_w1712_,
		_w1703_,
		_w10547_
	);
	LUT4 #(
		.INIT('h153f)
	) name9198 (
		\P1_InstQueue_reg[5][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1708_,
		_w1702_,
		_w10548_
	);
	LUT4 #(
		.INIT('h135f)
	) name9199 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1699_,
		_w1709_,
		_w10549_
	);
	LUT4 #(
		.INIT('h8000)
	) name9200 (
		_w10548_,
		_w10549_,
		_w10546_,
		_w10547_,
		_w10550_
	);
	LUT4 #(
		.INIT('h0111)
	) name9201 (
		_w1842_,
		_w1845_,
		_w10545_,
		_w10550_,
		_w10551_
	);
	LUT4 #(
		.INIT('h4000)
	) name9202 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('h1)
	) name9203 (
		_w10540_,
		_w10552_,
		_w10553_
	);
	LUT2 #(
		.INIT('h4)
	) name9204 (
		_w10539_,
		_w10553_,
		_w10554_
	);
	LUT4 #(
		.INIT('hecee)
	) name9205 (
		_w1933_,
		_w10536_,
		_w10538_,
		_w10554_,
		_w10555_
	);
	LUT2 #(
		.INIT('h2)
	) name9206 (
		\P1_EAX_reg[13]/NET0131 ,
		_w9102_,
		_w10556_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9207 (
		\P1_EAX_reg[13]/NET0131 ,
		_w9436_,
		_w9437_,
		_w10537_,
		_w10557_
	);
	LUT4 #(
		.INIT('h4000)
	) name9208 (
		\P1_EAX_reg[13]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9423_,
		_w10558_
	);
	LUT4 #(
		.INIT('h153f)
	) name9209 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[2][5]/NET0131 ,
		_w1688_,
		_w1712_,
		_w10559_
	);
	LUT4 #(
		.INIT('h153f)
	) name9210 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1691_,
		_w1705_,
		_w10560_
	);
	LUT4 #(
		.INIT('h135f)
	) name9211 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1696_,
		_w1706_,
		_w10561_
	);
	LUT4 #(
		.INIT('h135f)
	) name9212 (
		\P1_InstQueue_reg[3][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1692_,
		_w1711_,
		_w10562_
	);
	LUT4 #(
		.INIT('h8000)
	) name9213 (
		_w10561_,
		_w10562_,
		_w10559_,
		_w10560_,
		_w10563_
	);
	LUT4 #(
		.INIT('h135f)
	) name9214 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1698_,
		_w1709_,
		_w10564_
	);
	LUT4 #(
		.INIT('h135f)
	) name9215 (
		\P1_InstQueue_reg[12][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1694_,
		_w1708_,
		_w10565_
	);
	LUT4 #(
		.INIT('h153f)
	) name9216 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[5][5]/NET0131 ,
		_w1702_,
		_w1703_,
		_w10566_
	);
	LUT4 #(
		.INIT('h135f)
	) name9217 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1699_,
		_w1689_,
		_w10567_
	);
	LUT4 #(
		.INIT('h8000)
	) name9218 (
		_w10566_,
		_w10567_,
		_w10564_,
		_w10565_,
		_w10568_
	);
	LUT4 #(
		.INIT('h0111)
	) name9219 (
		_w1842_,
		_w1845_,
		_w10563_,
		_w10568_,
		_w10569_
	);
	LUT4 #(
		.INIT('h4000)
	) name9220 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10569_,
		_w10570_
	);
	LUT4 #(
		.INIT('h00fd)
	) name9221 (
		_w1855_,
		_w1861_,
		_w3467_,
		_w10570_,
		_w10571_
	);
	LUT2 #(
		.INIT('h4)
	) name9222 (
		_w10558_,
		_w10571_,
		_w10572_
	);
	LUT4 #(
		.INIT('hecee)
	) name9223 (
		_w1933_,
		_w10556_,
		_w10557_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h2)
	) name9224 (
		\P1_EAX_reg[12]/NET0131 ,
		_w9102_,
		_w10574_
	);
	LUT2 #(
		.INIT('h2)
	) name9225 (
		_w1867_,
		_w3464_,
		_w10575_
	);
	LUT3 #(
		.INIT('hd1)
	) name9226 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1867_,
		_w3464_,
		_w10576_
	);
	LUT4 #(
		.INIT('h00ec)
	) name9227 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w10576_,
		_w10577_
	);
	LUT4 #(
		.INIT('h4000)
	) name9228 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9422_,
		_w10578_
	);
	LUT4 #(
		.INIT('h153f)
	) name9229 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[12][4]/NET0131 ,
		_w1694_,
		_w1699_,
		_w10579_
	);
	LUT4 #(
		.INIT('h135f)
	) name9230 (
		\P1_InstQueue_reg[3][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1692_,
		_w1708_,
		_w10580_
	);
	LUT4 #(
		.INIT('h135f)
	) name9231 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[15][4]/NET0131 ,
		_w1696_,
		_w1705_,
		_w10581_
	);
	LUT4 #(
		.INIT('h135f)
	) name9232 (
		\P1_InstQueue_reg[7][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1691_,
		_w1711_,
		_w10582_
	);
	LUT4 #(
		.INIT('h8000)
	) name9233 (
		_w10581_,
		_w10582_,
		_w10579_,
		_w10580_,
		_w10583_
	);
	LUT4 #(
		.INIT('h135f)
	) name9234 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1698_,
		_w1689_,
		_w10584_
	);
	LUT4 #(
		.INIT('h153f)
	) name9235 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[2][4]/NET0131 ,
		_w1688_,
		_w1712_,
		_w10585_
	);
	LUT4 #(
		.INIT('h135f)
	) name9236 (
		\P1_InstQueue_reg[4][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1709_,
		_w1702_,
		_w10586_
	);
	LUT4 #(
		.INIT('h135f)
	) name9237 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1703_,
		_w1706_,
		_w10587_
	);
	LUT4 #(
		.INIT('h8000)
	) name9238 (
		_w10586_,
		_w10587_,
		_w10584_,
		_w10585_,
		_w10588_
	);
	LUT4 #(
		.INIT('h0111)
	) name9239 (
		_w1842_,
		_w1845_,
		_w10583_,
		_w10588_,
		_w10589_
	);
	LUT4 #(
		.INIT('h4000)
	) name9240 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10589_,
		_w10590_
	);
	LUT3 #(
		.INIT('h01)
	) name9241 (
		_w10578_,
		_w10590_,
		_w10577_,
		_w10591_
	);
	LUT4 #(
		.INIT('h5d00)
	) name9242 (
		\P1_EAX_reg[12]/NET0131 ,
		_w9437_,
		_w10504_,
		_w10591_,
		_w10592_
	);
	LUT3 #(
		.INIT('hce)
	) name9243 (
		_w1933_,
		_w10574_,
		_w10592_,
		_w10593_
	);
	LUT3 #(
		.INIT('ha2)
	) name9244 (
		\P3_uWord_reg[8]/NET0131 ,
		_w8341_,
		_w9529_,
		_w10594_
	);
	LUT2 #(
		.INIT('h2)
	) name9245 (
		_w1945_,
		_w2105_,
		_w10595_
	);
	LUT3 #(
		.INIT('h2a)
	) name9246 (
		\buf2_reg[8]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w10596_
	);
	LUT3 #(
		.INIT('h40)
	) name9247 (
		_w2060_,
		_w2047_,
		_w10596_,
		_w10597_
	);
	LUT3 #(
		.INIT('hc8)
	) name9248 (
		_w9975_,
		_w10595_,
		_w10597_,
		_w10598_
	);
	LUT2 #(
		.INIT('he)
	) name9249 (
		_w10594_,
		_w10598_,
		_w10599_
	);
	LUT2 #(
		.INIT('h2)
	) name9250 (
		\P1_EAX_reg[1]/NET0131 ,
		_w9102_,
		_w10600_
	);
	LUT3 #(
		.INIT('h40)
	) name9251 (
		\P1_EAX_reg[0]/NET0131 ,
		_w1804_,
		_w1826_,
		_w10601_
	);
	LUT4 #(
		.INIT('haa8a)
	) name9252 (
		\P1_EAX_reg[1]/NET0131 ,
		_w9436_,
		_w9437_,
		_w10601_,
		_w10602_
	);
	LUT3 #(
		.INIT('h02)
	) name9253 (
		_w1855_,
		_w1861_,
		_w3478_,
		_w10603_
	);
	LUT4 #(
		.INIT('h0111)
	) name9254 (
		_w1842_,
		_w1845_,
		_w3148_,
		_w3153_,
		_w10604_
	);
	LUT4 #(
		.INIT('h4000)
	) name9255 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w10604_,
		_w10605_
	);
	LUT2 #(
		.INIT('h2)
	) name9256 (
		\P1_EAX_reg[0]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w10606_
	);
	LUT3 #(
		.INIT('h80)
	) name9257 (
		_w1804_,
		_w1826_,
		_w10606_,
		_w10607_
	);
	LUT2 #(
		.INIT('h1)
	) name9258 (
		_w10605_,
		_w10607_,
		_w10608_
	);
	LUT2 #(
		.INIT('h4)
	) name9259 (
		_w10603_,
		_w10608_,
		_w10609_
	);
	LUT4 #(
		.INIT('hecee)
	) name9260 (
		_w1933_,
		_w10600_,
		_w10602_,
		_w10609_,
		_w10610_
	);
	LUT4 #(
		.INIT('h0001)
	) name9261 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10611_
	);
	LUT3 #(
		.INIT('hc8)
	) name9262 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		_w2215_,
		_w10611_,
		_w10612_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9263 (
		_w1988_,
		_w1993_,
		_w10611_,
		_w10612_,
		_w10613_
	);
	LUT4 #(
		.INIT('h2000)
	) name9264 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10614_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w10615_
	);
	LUT4 #(
		.INIT('h4000)
	) name9266 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10616_
	);
	LUT4 #(
		.INIT('h9fff)
	) name9267 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10617_
	);
	LUT4 #(
		.INIT('h030b)
	) name9268 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10617_,
		_w10618_
	);
	LUT3 #(
		.INIT('h80)
	) name9269 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w10619_
	);
	LUT4 #(
		.INIT('h8000)
	) name9270 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10620_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name9271 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10621_
	);
	LUT4 #(
		.INIT('hfd14)
	) name9272 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w10622_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9273 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w10623_
	);
	LUT4 #(
		.INIT('h153f)
	) name9274 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10614_,
		_w10616_,
		_w10624_
	);
	LUT2 #(
		.INIT('h2)
	) name9275 (
		_w2199_,
		_w10624_,
		_w10625_
	);
	LUT3 #(
		.INIT('h02)
	) name9276 (
		\buf2_reg[4]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10626_
	);
	LUT3 #(
		.INIT('h01)
	) name9277 (
		_w10623_,
		_w10625_,
		_w10626_,
		_w10627_
	);
	LUT2 #(
		.INIT('hb)
	) name9278 (
		_w10613_,
		_w10627_,
		_w10628_
	);
	LUT3 #(
		.INIT('h20)
	) name9279 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10629_
	);
	LUT4 #(
		.INIT('h0400)
	) name9280 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10630_
	);
	LUT3 #(
		.INIT('hc8)
	) name9281 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		_w2215_,
		_w10630_,
		_w10631_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9282 (
		_w1988_,
		_w1993_,
		_w10630_,
		_w10631_,
		_w10632_
	);
	LUT4 #(
		.INIT('h0080)
	) name9283 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10633_
	);
	LUT3 #(
		.INIT('h10)
	) name9284 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10634_
	);
	LUT4 #(
		.INIT('h0100)
	) name9285 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10635_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name9286 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10636_
	);
	LUT4 #(
		.INIT('h030b)
	) name9287 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10636_,
		_w10637_
	);
	LUT2 #(
		.INIT('h9)
	) name9288 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w10638_
	);
	LUT4 #(
		.INIT('h0600)
	) name9289 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10639_
	);
	LUT4 #(
		.INIT('h222a)
	) name9290 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w10640_
	);
	LUT4 #(
		.INIT('h153f)
	) name9291 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10633_,
		_w10635_,
		_w10641_
	);
	LUT2 #(
		.INIT('h2)
	) name9292 (
		_w2199_,
		_w10641_,
		_w10642_
	);
	LUT3 #(
		.INIT('h20)
	) name9293 (
		\buf2_reg[4]/NET0131 ,
		_w10637_,
		_w10639_,
		_w10643_
	);
	LUT3 #(
		.INIT('h01)
	) name9294 (
		_w10640_,
		_w10642_,
		_w10643_,
		_w10644_
	);
	LUT2 #(
		.INIT('hb)
	) name9295 (
		_w10632_,
		_w10644_,
		_w10645_
	);
	LUT4 #(
		.INIT('h0800)
	) name9296 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10646_
	);
	LUT3 #(
		.INIT('hc8)
	) name9297 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w2215_,
		_w10646_,
		_w10647_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9298 (
		_w1988_,
		_w1993_,
		_w10646_,
		_w10647_,
		_w10648_
	);
	LUT4 #(
		.INIT('h0200)
	) name9299 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10649_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name9300 (
		_w2194_,
		_w3055_,
		_w10629_,
		_w10649_,
		_w10650_
	);
	LUT3 #(
		.INIT('ha2)
	) name9301 (
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w10622_,
		_w10650_,
		_w10651_
	);
	LUT4 #(
		.INIT('h0200)
	) name9302 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10652_
	);
	LUT4 #(
		.INIT('h27ff)
	) name9303 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10634_,
		_w10653_
	);
	LUT4 #(
		.INIT('h2000)
	) name9304 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w10654_
	);
	LUT4 #(
		.INIT('hce00)
	) name9305 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w10654_,
		_w10655_
	);
	LUT3 #(
		.INIT('h0d)
	) name9306 (
		_w2199_,
		_w10653_,
		_w10655_,
		_w10656_
	);
	LUT2 #(
		.INIT('h4)
	) name9307 (
		_w10651_,
		_w10656_,
		_w10657_
	);
	LUT2 #(
		.INIT('hb)
	) name9308 (
		_w10648_,
		_w10657_,
		_w10658_
	);
	LUT4 #(
		.INIT('h1000)
	) name9309 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10659_
	);
	LUT3 #(
		.INIT('hc8)
	) name9310 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w2215_,
		_w10659_,
		_w10660_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9311 (
		_w1988_,
		_w1993_,
		_w10659_,
		_w10660_,
		_w10661_
	);
	LUT4 #(
		.INIT('h0b03)
	) name9312 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10639_,
		_w10662_
	);
	LUT4 #(
		.INIT('he7ff)
	) name9313 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10663_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9314 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w10664_
	);
	LUT4 #(
		.INIT('h135f)
	) name9315 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10630_,
		_w10652_,
		_w10665_
	);
	LUT2 #(
		.INIT('h2)
	) name9316 (
		_w2199_,
		_w10665_,
		_w10666_
	);
	LUT3 #(
		.INIT('h02)
	) name9317 (
		\buf2_reg[4]/NET0131 ,
		_w10662_,
		_w10663_,
		_w10667_
	);
	LUT3 #(
		.INIT('h01)
	) name9318 (
		_w10664_,
		_w10666_,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('hb)
	) name9319 (
		_w10661_,
		_w10668_,
		_w10669_
	);
	LUT3 #(
		.INIT('hc8)
	) name9320 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w2215_,
		_w10614_,
		_w10670_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9321 (
		_w1988_,
		_w1993_,
		_w10614_,
		_w10670_,
		_w10671_
	);
	LUT4 #(
		.INIT('hcfff)
	) name9322 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10672_
	);
	LUT4 #(
		.INIT('h0800)
	) name9323 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10673_
	);
	LUT3 #(
		.INIT('h23)
	) name9324 (
		_w3055_,
		_w6349_,
		_w10673_,
		_w10674_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name9325 (
		_w2194_,
		_w3055_,
		_w10672_,
		_w10673_,
		_w10675_
	);
	LUT3 #(
		.INIT('ha2)
	) name9326 (
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w10622_,
		_w10675_,
		_w10676_
	);
	LUT4 #(
		.INIT('h27ff)
	) name9327 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10629_,
		_w10677_
	);
	LUT2 #(
		.INIT('h2)
	) name9328 (
		\buf2_reg[4]/NET0131 ,
		_w10672_,
		_w10678_
	);
	LUT4 #(
		.INIT('h31f5)
	) name9329 (
		_w2199_,
		_w10674_,
		_w10677_,
		_w10678_,
		_w10679_
	);
	LUT2 #(
		.INIT('h4)
	) name9330 (
		_w10676_,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('hb)
	) name9331 (
		_w10671_,
		_w10680_,
		_w10681_
	);
	LUT3 #(
		.INIT('hc8)
	) name9332 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w2215_,
		_w10616_,
		_w10682_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9333 (
		_w1988_,
		_w1993_,
		_w10616_,
		_w10682_,
		_w10683_
	);
	LUT4 #(
		.INIT('h030b)
	) name9334 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10663_,
		_w10684_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name9335 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w10685_
	);
	LUT4 #(
		.INIT('h153f)
	) name9336 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10646_,
		_w10659_,
		_w10686_
	);
	LUT2 #(
		.INIT('h2)
	) name9337 (
		_w2199_,
		_w10686_,
		_w10687_
	);
	LUT3 #(
		.INIT('h02)
	) name9338 (
		\buf2_reg[4]/NET0131 ,
		_w10617_,
		_w10684_,
		_w10688_
	);
	LUT3 #(
		.INIT('h01)
	) name9339 (
		_w10685_,
		_w10687_,
		_w10688_,
		_w10689_
	);
	LUT2 #(
		.INIT('hb)
	) name9340 (
		_w10683_,
		_w10689_,
		_w10690_
	);
	LUT3 #(
		.INIT('hc8)
	) name9341 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w2215_,
		_w10620_,
		_w10691_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9342 (
		_w1988_,
		_w1993_,
		_w10620_,
		_w10691_,
		_w10692_
	);
	LUT4 #(
		.INIT('h030b)
	) name9343 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10672_,
		_w10693_
	);
	LUT4 #(
		.INIT('h3fff)
	) name9344 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10694_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9345 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w10695_
	);
	LUT4 #(
		.INIT('h135f)
	) name9346 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10614_,
		_w10659_,
		_w10696_
	);
	LUT2 #(
		.INIT('h2)
	) name9347 (
		_w2199_,
		_w10696_,
		_w10697_
	);
	LUT3 #(
		.INIT('h02)
	) name9348 (
		\buf2_reg[4]/NET0131 ,
		_w10693_,
		_w10694_,
		_w10698_
	);
	LUT3 #(
		.INIT('h01)
	) name9349 (
		_w10695_,
		_w10697_,
		_w10698_,
		_w10699_
	);
	LUT2 #(
		.INIT('hb)
	) name9350 (
		_w10692_,
		_w10699_,
		_w10700_
	);
	LUT4 #(
		.INIT('h0002)
	) name9351 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10701_
	);
	LUT3 #(
		.INIT('hc8)
	) name9352 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w2215_,
		_w10701_,
		_w10702_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9353 (
		_w1988_,
		_w1993_,
		_w10701_,
		_w10702_,
		_w10703_
	);
	LUT4 #(
		.INIT('h030b)
	) name9354 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10694_,
		_w10704_
	);
	LUT4 #(
		.INIT('hfffc)
	) name9355 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10705_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9356 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w10706_
	);
	LUT4 #(
		.INIT('h153f)
	) name9357 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10616_,
		_w10620_,
		_w10707_
	);
	LUT2 #(
		.INIT('h2)
	) name9358 (
		_w2199_,
		_w10707_,
		_w10708_
	);
	LUT3 #(
		.INIT('h02)
	) name9359 (
		\buf2_reg[4]/NET0131 ,
		_w10704_,
		_w10705_,
		_w10709_
	);
	LUT3 #(
		.INIT('h01)
	) name9360 (
		_w10706_,
		_w10708_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('hb)
	) name9361 (
		_w10703_,
		_w10710_,
		_w10711_
	);
	LUT3 #(
		.INIT('h02)
	) name9362 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10712_
	);
	LUT4 #(
		.INIT('h0004)
	) name9363 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10713_
	);
	LUT3 #(
		.INIT('hc8)
	) name9364 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w2215_,
		_w10713_,
		_w10714_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9365 (
		_w1988_,
		_w1993_,
		_w10713_,
		_w10714_,
		_w10715_
	);
	LUT4 #(
		.INIT('h030b)
	) name9366 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10621_,
		_w10716_
	);
	LUT4 #(
		.INIT('h0006)
	) name9367 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10717_
	);
	LUT4 #(
		.INIT('h222a)
	) name9368 (
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w10718_
	);
	LUT4 #(
		.INIT('h135f)
	) name9369 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10611_,
		_w10620_,
		_w10719_
	);
	LUT2 #(
		.INIT('h2)
	) name9370 (
		_w2199_,
		_w10719_,
		_w10720_
	);
	LUT3 #(
		.INIT('h20)
	) name9371 (
		\buf2_reg[4]/NET0131 ,
		_w10716_,
		_w10717_,
		_w10721_
	);
	LUT3 #(
		.INIT('h01)
	) name9372 (
		_w10718_,
		_w10720_,
		_w10721_,
		_w10722_
	);
	LUT2 #(
		.INIT('hb)
	) name9373 (
		_w10715_,
		_w10722_,
		_w10723_
	);
	LUT4 #(
		.INIT('h0008)
	) name9374 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10724_
	);
	LUT3 #(
		.INIT('hc8)
	) name9375 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w2215_,
		_w10724_,
		_w10725_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9376 (
		_w1988_,
		_w1993_,
		_w10724_,
		_w10725_,
		_w10726_
	);
	LUT4 #(
		.INIT('h030b)
	) name9377 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10705_,
		_w10727_
	);
	LUT4 #(
		.INIT('h222a)
	) name9378 (
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w10728_
	);
	LUT4 #(
		.INIT('h153f)
	) name9379 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10611_,
		_w10701_,
		_w10729_
	);
	LUT2 #(
		.INIT('h2)
	) name9380 (
		_w2199_,
		_w10729_,
		_w10730_
	);
	LUT3 #(
		.INIT('h08)
	) name9381 (
		\buf2_reg[4]/NET0131 ,
		_w10712_,
		_w10727_,
		_w10731_
	);
	LUT3 #(
		.INIT('h01)
	) name9382 (
		_w10728_,
		_w10730_,
		_w10731_,
		_w10732_
	);
	LUT2 #(
		.INIT('hb)
	) name9383 (
		_w10726_,
		_w10732_,
		_w10733_
	);
	LUT4 #(
		.INIT('h0010)
	) name9384 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10734_
	);
	LUT3 #(
		.INIT('hc8)
	) name9385 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w2215_,
		_w10734_,
		_w10735_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9386 (
		_w1988_,
		_w1993_,
		_w10734_,
		_w10735_,
		_w10736_
	);
	LUT4 #(
		.INIT('h0b03)
	) name9387 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10717_,
		_w10737_
	);
	LUT4 #(
		.INIT('hffe7)
	) name9388 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10738_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9389 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w10739_
	);
	LUT4 #(
		.INIT('h153f)
	) name9390 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10701_,
		_w10713_,
		_w10740_
	);
	LUT2 #(
		.INIT('h2)
	) name9391 (
		_w2199_,
		_w10740_,
		_w10741_
	);
	LUT3 #(
		.INIT('h02)
	) name9392 (
		\buf2_reg[4]/NET0131 ,
		_w10737_,
		_w10738_,
		_w10742_
	);
	LUT3 #(
		.INIT('h01)
	) name9393 (
		_w10739_,
		_w10741_,
		_w10742_,
		_w10743_
	);
	LUT2 #(
		.INIT('hb)
	) name9394 (
		_w10736_,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('h0020)
	) name9395 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10745_
	);
	LUT3 #(
		.INIT('hc8)
	) name9396 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w2215_,
		_w10745_,
		_w10746_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9397 (
		_w1988_,
		_w1993_,
		_w10745_,
		_w10746_,
		_w10747_
	);
	LUT4 #(
		.INIT('hffcf)
	) name9398 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10748_
	);
	LUT4 #(
		.INIT('h0008)
	) name9399 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10749_
	);
	LUT3 #(
		.INIT('h23)
	) name9400 (
		_w3055_,
		_w6349_,
		_w10749_,
		_w10750_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name9401 (
		_w2194_,
		_w3055_,
		_w10748_,
		_w10749_,
		_w10751_
	);
	LUT3 #(
		.INIT('ha2)
	) name9402 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		_w10622_,
		_w10751_,
		_w10752_
	);
	LUT4 #(
		.INIT('h27ff)
	) name9403 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10712_,
		_w10753_
	);
	LUT2 #(
		.INIT('h2)
	) name9404 (
		\buf2_reg[4]/NET0131 ,
		_w10748_,
		_w10754_
	);
	LUT4 #(
		.INIT('h31f5)
	) name9405 (
		_w2199_,
		_w10750_,
		_w10753_,
		_w10754_,
		_w10755_
	);
	LUT2 #(
		.INIT('h4)
	) name9406 (
		_w10752_,
		_w10755_,
		_w10756_
	);
	LUT2 #(
		.INIT('hb)
	) name9407 (
		_w10747_,
		_w10756_,
		_w10757_
	);
	LUT4 #(
		.INIT('h0040)
	) name9408 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10758_
	);
	LUT3 #(
		.INIT('hc8)
	) name9409 (
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w2215_,
		_w10758_,
		_w10759_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9410 (
		_w1988_,
		_w1993_,
		_w10758_,
		_w10759_,
		_w10760_
	);
	LUT4 #(
		.INIT('h030b)
	) name9411 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10738_,
		_w10761_
	);
	LUT4 #(
		.INIT('hff9f)
	) name9412 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10762_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9413 (
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w10763_
	);
	LUT4 #(
		.INIT('h153f)
	) name9414 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10724_,
		_w10734_,
		_w10764_
	);
	LUT2 #(
		.INIT('h2)
	) name9415 (
		_w2199_,
		_w10764_,
		_w10765_
	);
	LUT3 #(
		.INIT('h02)
	) name9416 (
		\buf2_reg[4]/NET0131 ,
		_w10761_,
		_w10762_,
		_w10766_
	);
	LUT3 #(
		.INIT('h01)
	) name9417 (
		_w10763_,
		_w10765_,
		_w10766_,
		_w10767_
	);
	LUT2 #(
		.INIT('hb)
	) name9418 (
		_w10760_,
		_w10767_,
		_w10768_
	);
	LUT3 #(
		.INIT('hc8)
	) name9419 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w2215_,
		_w10633_,
		_w10769_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9420 (
		_w1988_,
		_w1993_,
		_w10633_,
		_w10769_,
		_w10770_
	);
	LUT4 #(
		.INIT('h030b)
	) name9421 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10748_,
		_w10771_
	);
	LUT4 #(
		.INIT('hff3f)
	) name9422 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w10772_
	);
	LUT4 #(
		.INIT('h2a22)
	) name9423 (
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w10773_
	);
	LUT4 #(
		.INIT('h153f)
	) name9424 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10734_,
		_w10745_,
		_w10774_
	);
	LUT2 #(
		.INIT('h2)
	) name9425 (
		_w2199_,
		_w10774_,
		_w10775_
	);
	LUT3 #(
		.INIT('h02)
	) name9426 (
		\buf2_reg[4]/NET0131 ,
		_w10771_,
		_w10772_,
		_w10776_
	);
	LUT3 #(
		.INIT('h01)
	) name9427 (
		_w10773_,
		_w10775_,
		_w10776_,
		_w10777_
	);
	LUT2 #(
		.INIT('hb)
	) name9428 (
		_w10770_,
		_w10777_,
		_w10778_
	);
	LUT3 #(
		.INIT('hc8)
	) name9429 (
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w2215_,
		_w10635_,
		_w10779_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9430 (
		_w1988_,
		_w1993_,
		_w10635_,
		_w10779_,
		_w10780_
	);
	LUT4 #(
		.INIT('h030b)
	) name9431 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w10762_,
		_w10781_
	);
	LUT4 #(
		.INIT('h22a2)
	) name9432 (
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w10782_
	);
	LUT4 #(
		.INIT('h153f)
	) name9433 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10745_,
		_w10758_,
		_w10783_
	);
	LUT2 #(
		.INIT('h2)
	) name9434 (
		_w2199_,
		_w10783_,
		_w10784_
	);
	LUT3 #(
		.INIT('h02)
	) name9435 (
		\buf2_reg[4]/NET0131 ,
		_w10636_,
		_w10781_,
		_w10785_
	);
	LUT3 #(
		.INIT('h01)
	) name9436 (
		_w10782_,
		_w10784_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('hb)
	) name9437 (
		_w10780_,
		_w10786_,
		_w10787_
	);
	LUT3 #(
		.INIT('hc8)
	) name9438 (
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w2215_,
		_w10652_,
		_w10788_
	);
	LUT4 #(
		.INIT('h7f00)
	) name9439 (
		_w1988_,
		_w1993_,
		_w10652_,
		_w10788_,
		_w10789_
	);
	LUT4 #(
		.INIT('h135f)
	) name9440 (
		\buf2_reg[20]/NET0131 ,
		\buf2_reg[28]/NET0131 ,
		_w10633_,
		_w10758_,
		_w10790_
	);
	LUT4 #(
		.INIT('hef00)
	) name9441 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w10791_
	);
	LUT4 #(
		.INIT('h1000)
	) name9442 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w10792_
	);
	LUT4 #(
		.INIT('hddd0)
	) name9443 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w10791_,
		_w10792_,
		_w10793_
	);
	LUT4 #(
		.INIT('hcc08)
	) name9444 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w10790_,
		_w10793_,
		_w10794_
	);
	LUT3 #(
		.INIT('ha8)
	) name9445 (
		_w3055_,
		_w10791_,
		_w10792_,
		_w10795_
	);
	LUT2 #(
		.INIT('h2)
	) name9446 (
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w10622_,
		_w10796_
	);
	LUT2 #(
		.INIT('h1)
	) name9447 (
		_w10795_,
		_w10796_,
		_w10797_
	);
	LUT2 #(
		.INIT('h4)
	) name9448 (
		_w10794_,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('hb)
	) name9449 (
		_w10789_,
		_w10798_,
		_w10799_
	);
	LUT2 #(
		.INIT('h6)
	) name9450 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10800_
	);
	LUT2 #(
		.INIT('h4)
	) name9451 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w10801_
	);
	LUT2 #(
		.INIT('h8)
	) name9452 (
		_w6367_,
		_w10801_,
		_w10802_
	);
	LUT4 #(
		.INIT('h8000)
	) name9453 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w6368_,
		_w10802_,
		_w10803_
	);
	LUT3 #(
		.INIT('h06)
	) name9454 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10803_,
		_w10804_
	);
	LUT2 #(
		.INIT('h2)
	) name9455 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w10805_
	);
	LUT2 #(
		.INIT('h2)
	) name9456 (
		_w1939_,
		_w10805_,
		_w10806_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9457 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8093_,
		_w10804_,
		_w10806_,
		_w10807_
	);
	LUT4 #(
		.INIT('h00fe)
	) name9458 (
		_w1795_,
		_w1797_,
		_w1802_,
		_w1852_,
		_w10808_
	);
	LUT2 #(
		.INIT('h2)
	) name9459 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10808_,
		_w10809_
	);
	LUT4 #(
		.INIT('h8000)
	) name9460 (
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w10810_
	);
	LUT4 #(
		.INIT('h8000)
	) name9461 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w10810_,
		_w10811_
	);
	LUT4 #(
		.INIT('h8000)
	) name9462 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10811_,
		_w10812_
	);
	LUT3 #(
		.INIT('h80)
	) name9463 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w10812_,
		_w10813_
	);
	LUT4 #(
		.INIT('h8000)
	) name9464 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w10812_,
		_w10814_
	);
	LUT3 #(
		.INIT('h84)
	) name9465 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w1930_,
		_w10814_,
		_w10815_
	);
	LUT4 #(
		.INIT('h2010)
	) name9466 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w1858_,
		_w1930_,
		_w10814_,
		_w10816_
	);
	LUT3 #(
		.INIT('h01)
	) name9467 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10817_
	);
	LUT4 #(
		.INIT('h3332)
	) name9468 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10818_
	);
	LUT3 #(
		.INIT('h02)
	) name9469 (
		_w1797_,
		_w10818_,
		_w10816_,
		_w10819_
	);
	LUT4 #(
		.INIT('h0001)
	) name9470 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w10820_
	);
	LUT4 #(
		.INIT('h0100)
	) name9471 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w10820_,
		_w10821_
	);
	LUT4 #(
		.INIT('h0100)
	) name9472 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w10821_,
		_w10822_
	);
	LUT4 #(
		.INIT('h0100)
	) name9473 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w10822_,
		_w10823_
	);
	LUT3 #(
		.INIT('h8c)
	) name9474 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10823_,
		_w10824_
	);
	LUT3 #(
		.INIT('h21)
	) name9475 (
		\P1_EBX_reg[14]/NET0131 ,
		_w1930_,
		_w10824_,
		_w10825_
	);
	LUT2 #(
		.INIT('h2)
	) name9476 (
		_w1795_,
		_w10815_,
		_w10826_
	);
	LUT4 #(
		.INIT('h4544)
	) name9477 (
		_w1852_,
		_w10819_,
		_w10825_,
		_w10826_,
		_w10827_
	);
	LUT4 #(
		.INIT('hfe25)
	) name9478 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w10828_
	);
	LUT2 #(
		.INIT('h2)
	) name9479 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10828_,
		_w10829_
	);
	LUT3 #(
		.INIT('h07)
	) name9480 (
		\P1_PhyAddrPointer_reg[14]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10830_
	);
	LUT2 #(
		.INIT('h4)
	) name9481 (
		_w10829_,
		_w10830_,
		_w10831_
	);
	LUT4 #(
		.INIT('h5700)
	) name9482 (
		_w1933_,
		_w10809_,
		_w10827_,
		_w10831_,
		_w10832_
	);
	LUT2 #(
		.INIT('hb)
	) name9483 (
		_w10807_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h8)
	) name9484 (
		_w6370_,
		_w10802_,
		_w10834_
	);
	LUT3 #(
		.INIT('h06)
	) name9485 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10834_,
		_w10835_
	);
	LUT2 #(
		.INIT('h2)
	) name9486 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w10836_
	);
	LUT2 #(
		.INIT('h2)
	) name9487 (
		_w1939_,
		_w10836_,
		_w10837_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9488 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7552_,
		_w10835_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h2)
	) name9489 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w10808_,
		_w10839_
	);
	LUT4 #(
		.INIT('h9030)
	) name9490 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w1930_,
		_w10814_,
		_w10840_
	);
	LUT4 #(
		.INIT('h3332)
	) name9491 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10841_
	);
	LUT4 #(
		.INIT('h080a)
	) name9492 (
		_w1797_,
		_w1858_,
		_w10841_,
		_w10840_,
		_w10842_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9493 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10823_,
		_w10843_
	);
	LUT3 #(
		.INIT('h21)
	) name9494 (
		\P1_EBX_reg[15]/NET0131 ,
		_w1930_,
		_w10843_,
		_w10844_
	);
	LUT2 #(
		.INIT('h2)
	) name9495 (
		_w1795_,
		_w10840_,
		_w10845_
	);
	LUT4 #(
		.INIT('h4544)
	) name9496 (
		_w1852_,
		_w10842_,
		_w10844_,
		_w10845_,
		_w10846_
	);
	LUT2 #(
		.INIT('h2)
	) name9497 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w10828_,
		_w10847_
	);
	LUT3 #(
		.INIT('h07)
	) name9498 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10848_
	);
	LUT2 #(
		.INIT('h4)
	) name9499 (
		_w10847_,
		_w10848_,
		_w10849_
	);
	LUT4 #(
		.INIT('h5700)
	) name9500 (
		_w1933_,
		_w10839_,
		_w10846_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('hb)
	) name9501 (
		_w10838_,
		_w10850_,
		_w10851_
	);
	LUT3 #(
		.INIT('h80)
	) name9502 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		_w6370_,
		_w10802_,
		_w10852_
	);
	LUT4 #(
		.INIT('hf096)
	) name9503 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w8111_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h2)
	) name9504 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10854_
	);
	LUT2 #(
		.INIT('h2)
	) name9505 (
		_w1939_,
		_w10854_,
		_w10855_
	);
	LUT3 #(
		.INIT('he0)
	) name9506 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w10853_,
		_w10855_,
		_w10856_
	);
	LUT2 #(
		.INIT('h2)
	) name9507 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w10808_,
		_w10857_
	);
	LUT4 #(
		.INIT('h8000)
	) name9508 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10814_,
		_w10858_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9509 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w10814_,
		_w10859_
	);
	LUT3 #(
		.INIT('h04)
	) name9510 (
		_w1858_,
		_w1930_,
		_w10859_,
		_w10860_
	);
	LUT4 #(
		.INIT('h3332)
	) name9511 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[16]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10861_
	);
	LUT2 #(
		.INIT('h2)
	) name9512 (
		_w1797_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h1)
	) name9513 (
		\P1_EBX_reg[14]/NET0131 ,
		\P1_EBX_reg[15]/NET0131 ,
		_w10863_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9514 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10823_,
		_w10863_,
		_w10864_
	);
	LUT3 #(
		.INIT('h21)
	) name9515 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1930_,
		_w10864_,
		_w10865_
	);
	LUT3 #(
		.INIT('ha2)
	) name9516 (
		_w1795_,
		_w1930_,
		_w10859_,
		_w10866_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name9517 (
		_w10860_,
		_w10862_,
		_w10865_,
		_w10866_,
		_w10867_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name9518 (
		_w1852_,
		_w1933_,
		_w10857_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h2)
	) name9519 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w10828_,
		_w10869_
	);
	LUT3 #(
		.INIT('h07)
	) name9520 (
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10870_
	);
	LUT2 #(
		.INIT('h4)
	) name9521 (
		_w10869_,
		_w10870_,
		_w10871_
	);
	LUT2 #(
		.INIT('h4)
	) name9522 (
		_w10868_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('hb)
	) name9523 (
		_w10856_,
		_w10872_,
		_w10873_
	);
	LUT4 #(
		.INIT('h8000)
	) name9524 (
		\P1_PhyAddrPointer_reg[15]/NET0131 ,
		\P1_PhyAddrPointer_reg[16]/NET0131 ,
		_w6370_,
		_w10802_,
		_w10874_
	);
	LUT3 #(
		.INIT('h06)
	) name9525 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10874_,
		_w10875_
	);
	LUT2 #(
		.INIT('h2)
	) name9526 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w10876_
	);
	LUT2 #(
		.INIT('h2)
	) name9527 (
		_w1939_,
		_w10876_,
		_w10877_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9528 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8119_,
		_w10875_,
		_w10877_,
		_w10878_
	);
	LUT3 #(
		.INIT('h84)
	) name9529 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1930_,
		_w10858_,
		_w10879_
	);
	LUT4 #(
		.INIT('h3222)
	) name9530 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[17]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10880_
	);
	LUT4 #(
		.INIT('h000d)
	) name9531 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w10880_,
		_w10881_
	);
	LUT4 #(
		.INIT('h7b00)
	) name9532 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1930_,
		_w10858_,
		_w10881_,
		_w10882_
	);
	LUT4 #(
		.INIT('ha200)
	) name9533 (
		\P1_EBX_reg[17]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w10883_
	);
	LUT3 #(
		.INIT('h08)
	) name9534 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1842_,
		_w1851_,
		_w10884_
	);
	LUT2 #(
		.INIT('h1)
	) name9535 (
		_w10883_,
		_w10884_,
		_w10885_
	);
	LUT3 #(
		.INIT('h8a)
	) name9536 (
		_w1797_,
		_w10882_,
		_w10885_,
		_w10886_
	);
	LUT4 #(
		.INIT('hf301)
	) name9537 (
		_w1795_,
		_w1797_,
		_w1802_,
		_w1852_,
		_w10887_
	);
	LUT2 #(
		.INIT('h8)
	) name9538 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w10887_,
		_w10888_
	);
	LUT4 #(
		.INIT('h1000)
	) name9539 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[16]/NET0131 ,
		_w10823_,
		_w10863_,
		_w10889_
	);
	LUT4 #(
		.INIT('h0509)
	) name9540 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w10889_,
		_w10890_
	);
	LUT3 #(
		.INIT('h02)
	) name9541 (
		_w4709_,
		_w10879_,
		_w10890_,
		_w10891_
	);
	LUT4 #(
		.INIT('haaa8)
	) name9542 (
		_w1933_,
		_w10888_,
		_w10886_,
		_w10891_,
		_w10892_
	);
	LUT2 #(
		.INIT('h2)
	) name9543 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w10828_,
		_w10893_
	);
	LUT3 #(
		.INIT('h07)
	) name9544 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10894_
	);
	LUT2 #(
		.INIT('h4)
	) name9545 (
		_w10893_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h4)
	) name9546 (
		_w10892_,
		_w10895_,
		_w10896_
	);
	LUT2 #(
		.INIT('hb)
	) name9547 (
		_w10878_,
		_w10896_,
		_w10897_
	);
	LUT3 #(
		.INIT('h80)
	) name9548 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6372_,
		_w10852_,
		_w10898_
	);
	LUT4 #(
		.INIT('hf096)
	) name9549 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w8130_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h2)
	) name9550 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10900_
	);
	LUT2 #(
		.INIT('h2)
	) name9551 (
		_w1939_,
		_w10900_,
		_w10901_
	);
	LUT3 #(
		.INIT('he0)
	) name9552 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w10899_,
		_w10901_,
		_w10902_
	);
	LUT2 #(
		.INIT('h2)
	) name9553 (
		\P1_rEIP_reg[18]/NET0131 ,
		_w10808_,
		_w10903_
	);
	LUT4 #(
		.INIT('h3332)
	) name9554 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10904_
	);
	LUT3 #(
		.INIT('h02)
	) name9555 (
		_w1797_,
		_w1852_,
		_w10904_,
		_w10905_
	);
	LUT3 #(
		.INIT('h8c)
	) name9556 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10889_,
		_w10906_
	);
	LUT4 #(
		.INIT('hd0e0)
	) name9557 (
		\P1_EBX_reg[18]/NET0131 ,
		_w1930_,
		_w4709_,
		_w10906_,
		_w10907_
	);
	LUT3 #(
		.INIT('h80)
	) name9558 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10858_,
		_w10908_
	);
	LUT3 #(
		.INIT('h6c)
	) name9559 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10858_,
		_w10909_
	);
	LUT4 #(
		.INIT('h0020)
	) name9560 (
		_w1797_,
		_w1852_,
		_w1858_,
		_w10904_,
		_w10910_
	);
	LUT3 #(
		.INIT('h02)
	) name9561 (
		_w1930_,
		_w10909_,
		_w10910_,
		_w10911_
	);
	LUT4 #(
		.INIT('h5501)
	) name9562 (
		_w10903_,
		_w10905_,
		_w10907_,
		_w10911_,
		_w10912_
	);
	LUT2 #(
		.INIT('h2)
	) name9563 (
		\P1_rEIP_reg[18]/NET0131 ,
		_w10828_,
		_w10913_
	);
	LUT3 #(
		.INIT('h07)
	) name9564 (
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10914_
	);
	LUT2 #(
		.INIT('h4)
	) name9565 (
		_w10913_,
		_w10914_,
		_w10915_
	);
	LUT3 #(
		.INIT('hd0)
	) name9566 (
		_w1933_,
		_w10912_,
		_w10915_,
		_w10916_
	);
	LUT2 #(
		.INIT('hb)
	) name9567 (
		_w10902_,
		_w10916_,
		_w10917_
	);
	LUT4 #(
		.INIT('h8000)
	) name9568 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		\P1_PhyAddrPointer_reg[18]/NET0131 ,
		_w6372_,
		_w10852_,
		_w10918_
	);
	LUT3 #(
		.INIT('h06)
	) name9569 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10918_,
		_w10919_
	);
	LUT2 #(
		.INIT('h2)
	) name9570 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w10920_
	);
	LUT2 #(
		.INIT('h2)
	) name9571 (
		_w1939_,
		_w10920_,
		_w10921_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9572 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7570_,
		_w10919_,
		_w10921_,
		_w10922_
	);
	LUT4 #(
		.INIT('h8000)
	) name9573 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w10858_,
		_w10923_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9574 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w10858_,
		_w10924_
	);
	LUT4 #(
		.INIT('h3222)
	) name9575 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[19]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10925_
	);
	LUT4 #(
		.INIT('h000d)
	) name9576 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w10925_,
		_w10926_
	);
	LUT3 #(
		.INIT('h08)
	) name9577 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w1842_,
		_w1851_,
		_w10927_
	);
	LUT4 #(
		.INIT('ha200)
	) name9578 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w10928_
	);
	LUT2 #(
		.INIT('h1)
	) name9579 (
		_w10927_,
		_w10928_,
		_w10929_
	);
	LUT4 #(
		.INIT('h2f00)
	) name9580 (
		_w1930_,
		_w10924_,
		_w10926_,
		_w10929_,
		_w10930_
	);
	LUT2 #(
		.INIT('h2)
	) name9581 (
		_w1797_,
		_w10930_,
		_w10931_
	);
	LUT2 #(
		.INIT('h8)
	) name9582 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10887_,
		_w10932_
	);
	LUT2 #(
		.INIT('h1)
	) name9583 (
		\P1_EBX_reg[17]/NET0131 ,
		\P1_EBX_reg[18]/NET0131 ,
		_w10933_
	);
	LUT3 #(
		.INIT('h2a)
	) name9584 (
		\P1_EBX_reg[31]/NET0131 ,
		_w10889_,
		_w10933_,
		_w10934_
	);
	LUT3 #(
		.INIT('h21)
	) name9585 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1930_,
		_w10934_,
		_w10935_
	);
	LUT3 #(
		.INIT('hc4)
	) name9586 (
		_w1930_,
		_w4709_,
		_w10924_,
		_w10936_
	);
	LUT3 #(
		.INIT('h45)
	) name9587 (
		_w10932_,
		_w10935_,
		_w10936_,
		_w10937_
	);
	LUT2 #(
		.INIT('h2)
	) name9588 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10828_,
		_w10938_
	);
	LUT3 #(
		.INIT('h07)
	) name9589 (
		\P1_PhyAddrPointer_reg[19]/NET0131 ,
		_w2234_,
		_w3406_,
		_w10939_
	);
	LUT2 #(
		.INIT('h4)
	) name9590 (
		_w10938_,
		_w10939_,
		_w10940_
	);
	LUT4 #(
		.INIT('h7500)
	) name9591 (
		_w1933_,
		_w10931_,
		_w10937_,
		_w10940_,
		_w10941_
	);
	LUT2 #(
		.INIT('hb)
	) name9592 (
		_w10922_,
		_w10941_,
		_w10942_
	);
	LUT4 #(
		.INIT('h3993)
	) name9593 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10943_
	);
	LUT2 #(
		.INIT('h2)
	) name9594 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w10944_
	);
	LUT2 #(
		.INIT('h2)
	) name9595 (
		_w1939_,
		_w10944_,
		_w10945_
	);
	LUT2 #(
		.INIT('h2)
	) name9596 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w10808_,
		_w10946_
	);
	LUT2 #(
		.INIT('h6)
	) name9597 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		_w10947_
	);
	LUT3 #(
		.INIT('h90)
	) name9598 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10948_
	);
	LUT2 #(
		.INIT('h1)
	) name9599 (
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10949_
	);
	LUT2 #(
		.INIT('h1)
	) name9600 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w10950_
	);
	LUT4 #(
		.INIT('h0111)
	) name9601 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10951_
	);
	LUT4 #(
		.INIT('h00fe)
	) name9602 (
		_w1930_,
		_w10949_,
		_w10948_,
		_w10951_,
		_w10952_
	);
	LUT3 #(
		.INIT('h02)
	) name9603 (
		_w1795_,
		_w1852_,
		_w10952_,
		_w10953_
	);
	LUT3 #(
		.INIT('h02)
	) name9604 (
		_w1802_,
		_w1852_,
		_w1848_,
		_w10954_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9605 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10955_
	);
	LUT3 #(
		.INIT('h10)
	) name9606 (
		_w1858_,
		_w1861_,
		_w10950_,
		_w10956_
	);
	LUT2 #(
		.INIT('h1)
	) name9607 (
		_w10955_,
		_w10956_,
		_w10957_
	);
	LUT3 #(
		.INIT('h02)
	) name9608 (
		_w1797_,
		_w1852_,
		_w10957_,
		_w10958_
	);
	LUT3 #(
		.INIT('h01)
	) name9609 (
		_w10954_,
		_w10958_,
		_w10953_,
		_w10959_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9610 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w2234_,
		_w10828_,
		_w10960_
	);
	LUT4 #(
		.INIT('h7500)
	) name9611 (
		_w1933_,
		_w10946_,
		_w10959_,
		_w10960_,
		_w10961_
	);
	LUT4 #(
		.INIT('he0ff)
	) name9612 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w10943_,
		_w10945_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h8)
	) name9613 (
		_w7569_,
		_w10852_,
		_w10963_
	);
	LUT3 #(
		.INIT('h06)
	) name9614 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10963_,
		_w10964_
	);
	LUT2 #(
		.INIT('h2)
	) name9615 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10965_
	);
	LUT2 #(
		.INIT('h2)
	) name9616 (
		_w1939_,
		_w10965_,
		_w10966_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9617 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7584_,
		_w10964_,
		_w10966_,
		_w10967_
	);
	LUT2 #(
		.INIT('h2)
	) name9618 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w10808_,
		_w10968_
	);
	LUT4 #(
		.INIT('h3332)
	) name9619 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w1858_,
		_w1861_,
		_w10969_
	);
	LUT2 #(
		.INIT('h2)
	) name9620 (
		_w1797_,
		_w10969_,
		_w10970_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9621 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10889_,
		_w10933_,
		_w10971_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9622 (
		\P1_EBX_reg[20]/NET0131 ,
		_w1795_,
		_w1930_,
		_w10971_,
		_w10972_
	);
	LUT2 #(
		.INIT('h8)
	) name9623 (
		\P1_rEIP_reg[19]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10973_
	);
	LUT4 #(
		.INIT('h8000)
	) name9624 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10858_,
		_w10973_,
		_w10974_
	);
	LUT4 #(
		.INIT('hf070)
	) name9625 (
		_w1797_,
		_w1858_,
		_w1930_,
		_w10969_,
		_w10975_
	);
	LUT4 #(
		.INIT('h9300)
	) name9626 (
		\P1_rEIP_reg[19]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w10908_,
		_w10975_,
		_w10976_
	);
	LUT4 #(
		.INIT('h0054)
	) name9627 (
		_w1852_,
		_w10970_,
		_w10972_,
		_w10976_,
		_w10977_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9628 (
		\P1_PhyAddrPointer_reg[20]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w2234_,
		_w10828_,
		_w10978_
	);
	LUT4 #(
		.INIT('h5700)
	) name9629 (
		_w1933_,
		_w10968_,
		_w10977_,
		_w10978_,
		_w10979_
	);
	LUT2 #(
		.INIT('hb)
	) name9630 (
		_w10967_,
		_w10979_,
		_w10980_
	);
	LUT3 #(
		.INIT('h80)
	) name9631 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w7583_,
		_w10852_,
		_w10981_
	);
	LUT3 #(
		.INIT('h06)
	) name9632 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10981_,
		_w10982_
	);
	LUT2 #(
		.INIT('h2)
	) name9633 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w10983_
	);
	LUT2 #(
		.INIT('h2)
	) name9634 (
		_w1939_,
		_w10983_,
		_w10984_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9635 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8146_,
		_w10982_,
		_w10984_,
		_w10985_
	);
	LUT4 #(
		.INIT('h3222)
	) name9636 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w10986_
	);
	LUT4 #(
		.INIT('h000d)
	) name9637 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w10986_,
		_w10987_
	);
	LUT4 #(
		.INIT('h7b00)
	) name9638 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w1930_,
		_w10974_,
		_w10987_,
		_w10988_
	);
	LUT4 #(
		.INIT('ha200)
	) name9639 (
		\P1_EBX_reg[21]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w10989_
	);
	LUT3 #(
		.INIT('h08)
	) name9640 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w1842_,
		_w1851_,
		_w10990_
	);
	LUT2 #(
		.INIT('h1)
	) name9641 (
		_w10989_,
		_w10990_,
		_w10991_
	);
	LUT3 #(
		.INIT('h8a)
	) name9642 (
		_w1797_,
		_w10988_,
		_w10991_,
		_w10992_
	);
	LUT2 #(
		.INIT('h8)
	) name9643 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w10887_,
		_w10993_
	);
	LUT4 #(
		.INIT('h1000)
	) name9644 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w10889_,
		_w10933_,
		_w10994_
	);
	LUT4 #(
		.INIT('h0509)
	) name9645 (
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w10994_,
		_w10995_
	);
	LUT4 #(
		.INIT('h70b0)
	) name9646 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w1930_,
		_w4709_,
		_w10974_,
		_w10996_
	);
	LUT3 #(
		.INIT('h45)
	) name9647 (
		_w10993_,
		_w10995_,
		_w10996_,
		_w10997_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9648 (
		\P1_PhyAddrPointer_reg[21]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w2234_,
		_w10828_,
		_w10998_
	);
	LUT4 #(
		.INIT('h7500)
	) name9649 (
		_w1933_,
		_w10992_,
		_w10997_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('hb)
	) name9650 (
		_w10985_,
		_w10999_,
		_w11000_
	);
	LUT4 #(
		.INIT('h8000)
	) name9651 (
		\P1_PhyAddrPointer_reg[17]/NET0131 ,
		_w6363_,
		_w6372_,
		_w10852_,
		_w11001_
	);
	LUT3 #(
		.INIT('h06)
	) name9652 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11001_,
		_w11002_
	);
	LUT2 #(
		.INIT('h2)
	) name9653 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w11003_
	);
	LUT2 #(
		.INIT('h2)
	) name9654 (
		_w1939_,
		_w11003_,
		_w11004_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9655 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7598_,
		_w11002_,
		_w11004_,
		_w11005_
	);
	LUT2 #(
		.INIT('h2)
	) name9656 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w10808_,
		_w11006_
	);
	LUT4 #(
		.INIT('h3332)
	) name9657 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11007_
	);
	LUT2 #(
		.INIT('h2)
	) name9658 (
		_w1797_,
		_w11007_,
		_w11008_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		_w11009_
	);
	LUT4 #(
		.INIT('h4000)
	) name9660 (
		\P1_EBX_reg[19]/NET0131 ,
		_w10889_,
		_w10933_,
		_w11009_,
		_w11010_
	);
	LUT4 #(
		.INIT('h0509)
	) name9661 (
		\P1_EBX_reg[22]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w11010_,
		_w11011_
	);
	LUT3 #(
		.INIT('h31)
	) name9662 (
		_w1795_,
		_w11008_,
		_w11011_,
		_w11012_
	);
	LUT4 #(
		.INIT('hf070)
	) name9663 (
		_w1797_,
		_w1858_,
		_w1930_,
		_w11007_,
		_w11013_
	);
	LUT4 #(
		.INIT('h9300)
	) name9664 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w10974_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h1)
	) name9665 (
		_w1852_,
		_w11014_,
		_w11015_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9666 (
		_w1933_,
		_w11006_,
		_w11012_,
		_w11015_,
		_w11016_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9667 (
		\P1_PhyAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11017_
	);
	LUT3 #(
		.INIT('hef)
	) name9668 (
		_w11016_,
		_w11005_,
		_w11017_,
		_w11018_
	);
	LUT2 #(
		.INIT('h8)
	) name9669 (
		_w6996_,
		_w10852_,
		_w11019_
	);
	LUT3 #(
		.INIT('h06)
	) name9670 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('h2)
	) name9671 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w11021_
	);
	LUT2 #(
		.INIT('h2)
	) name9672 (
		_w1939_,
		_w11021_,
		_w11022_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9673 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6998_,
		_w11020_,
		_w11022_,
		_w11023_
	);
	LUT3 #(
		.INIT('h80)
	) name9674 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w11024_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9675 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w10974_,
		_w11025_
	);
	LUT2 #(
		.INIT('h2)
	) name9676 (
		_w1930_,
		_w11025_,
		_w11026_
	);
	LUT4 #(
		.INIT('h3222)
	) name9677 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w11027_
	);
	LUT3 #(
		.INIT('h08)
	) name9678 (
		_w1797_,
		_w1859_,
		_w11027_,
		_w11028_
	);
	LUT3 #(
		.INIT('h01)
	) name9679 (
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		\P1_EBX_reg[22]/NET0131 ,
		_w11029_
	);
	LUT4 #(
		.INIT('h4000)
	) name9680 (
		\P1_EBX_reg[19]/NET0131 ,
		_w10889_,
		_w10933_,
		_w11029_,
		_w11030_
	);
	LUT4 #(
		.INIT('h0509)
	) name9681 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w11030_,
		_w11031_
	);
	LUT3 #(
		.INIT('h31)
	) name9682 (
		_w4709_,
		_w11028_,
		_w11031_,
		_w11032_
	);
	LUT4 #(
		.INIT('ha200)
	) name9683 (
		\P1_EBX_reg[23]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w11033_
	);
	LUT3 #(
		.INIT('h08)
	) name9684 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w1842_,
		_w1851_,
		_w11034_
	);
	LUT2 #(
		.INIT('h1)
	) name9685 (
		_w11033_,
		_w11034_,
		_w11035_
	);
	LUT2 #(
		.INIT('h2)
	) name9686 (
		_w1797_,
		_w11035_,
		_w11036_
	);
	LUT3 #(
		.INIT('h07)
	) name9687 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w10887_,
		_w11036_,
		_w11037_
	);
	LUT4 #(
		.INIT('h02aa)
	) name9688 (
		_w1933_,
		_w11026_,
		_w11032_,
		_w11037_,
		_w11038_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9689 (
		\P1_PhyAddrPointer_reg[23]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11039_
	);
	LUT3 #(
		.INIT('hef)
	) name9690 (
		_w11038_,
		_w11023_,
		_w11039_,
		_w11040_
	);
	LUT4 #(
		.INIT('h4000)
	) name9691 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w11041_
	);
	LUT3 #(
		.INIT('h06)
	) name9692 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11041_,
		_w11042_
	);
	LUT2 #(
		.INIT('h2)
	) name9693 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w11043_
	);
	LUT2 #(
		.INIT('h2)
	) name9694 (
		_w1679_,
		_w11043_,
		_w11044_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9695 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8750_,
		_w11042_,
		_w11044_,
		_w11045_
	);
	LUT4 #(
		.INIT('h0a06)
	) name9696 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w9755_,
		_w11046_
	);
	LUT4 #(
		.INIT('h0104)
	) name9697 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w1605_,
		_w9770_,
		_w11047_
	);
	LUT2 #(
		.INIT('h1)
	) name9698 (
		_w11046_,
		_w11047_,
		_w11048_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9699 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[10]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11049_
	);
	LUT4 #(
		.INIT('h1040)
	) name9700 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		_w1612_,
		_w9770_,
		_w11050_
	);
	LUT2 #(
		.INIT('h1)
	) name9701 (
		_w11049_,
		_w11050_,
		_w11051_
	);
	LUT4 #(
		.INIT('hf531)
	) name9702 (
		_w1565_,
		_w1566_,
		_w11048_,
		_w11051_,
		_w11052_
	);
	LUT4 #(
		.INIT('h5750)
	) name9703 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w1569_,
		_w1602_,
		_w11052_,
		_w11053_
	);
	LUT2 #(
		.INIT('h2)
	) name9704 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w9799_,
		_w11054_
	);
	LUT3 #(
		.INIT('h07)
	) name9705 (
		\P2_PhyAddrPointer_reg[10]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11055_
	);
	LUT2 #(
		.INIT('h4)
	) name9706 (
		_w11054_,
		_w11055_,
		_w11056_
	);
	LUT3 #(
		.INIT('hd0)
	) name9707 (
		_w1678_,
		_w11053_,
		_w11056_,
		_w11057_
	);
	LUT2 #(
		.INIT('hb)
	) name9708 (
		_w11045_,
		_w11057_,
		_w11058_
	);
	LUT2 #(
		.INIT('h8)
	) name9709 (
		_w6361_,
		_w11001_,
		_w11059_
	);
	LUT4 #(
		.INIT('hf096)
	) name9710 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w7608_,
		_w11059_,
		_w11060_
	);
	LUT2 #(
		.INIT('h2)
	) name9711 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w11061_
	);
	LUT2 #(
		.INIT('h2)
	) name9712 (
		_w1939_,
		_w11061_,
		_w11062_
	);
	LUT3 #(
		.INIT('he0)
	) name9713 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w11060_,
		_w11062_,
		_w11063_
	);
	LUT4 #(
		.INIT('h8444)
	) name9714 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w1930_,
		_w10974_,
		_w11024_,
		_w11064_
	);
	LUT4 #(
		.INIT('h3222)
	) name9715 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[24]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w11065_
	);
	LUT4 #(
		.INIT('h000d)
	) name9716 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w11065_,
		_w11066_
	);
	LUT4 #(
		.INIT('ha200)
	) name9717 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w11067_
	);
	LUT3 #(
		.INIT('h08)
	) name9718 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w1842_,
		_w1851_,
		_w11068_
	);
	LUT2 #(
		.INIT('h1)
	) name9719 (
		_w11067_,
		_w11068_,
		_w11069_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9720 (
		_w1797_,
		_w11064_,
		_w11066_,
		_w11069_,
		_w11070_
	);
	LUT3 #(
		.INIT('h8c)
	) name9721 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11030_,
		_w11071_
	);
	LUT3 #(
		.INIT('h21)
	) name9722 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1930_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h2)
	) name9723 (
		_w4709_,
		_w11064_,
		_w11073_
	);
	LUT2 #(
		.INIT('h8)
	) name9724 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w10887_,
		_w11074_
	);
	LUT4 #(
		.INIT('h000b)
	) name9725 (
		_w11072_,
		_w11073_,
		_w11074_,
		_w11070_,
		_w11075_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9726 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11076_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name9727 (
		_w1933_,
		_w11075_,
		_w11063_,
		_w11076_,
		_w11077_
	);
	LUT3 #(
		.INIT('h06)
	) name9728 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9792_,
		_w11078_
	);
	LUT4 #(
		.INIT('hf999)
	) name9729 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w7634_,
		_w9792_,
		_w11079_
	);
	LUT2 #(
		.INIT('h2)
	) name9730 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w11080_
	);
	LUT2 #(
		.INIT('h2)
	) name9731 (
		_w1679_,
		_w11080_,
		_w11081_
	);
	LUT4 #(
		.INIT('heb00)
	) name9732 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7632_,
		_w11079_,
		_w11081_,
		_w11082_
	);
	LUT3 #(
		.INIT('h8c)
	) name9733 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w11083_
	);
	LUT4 #(
		.INIT('hfd00)
	) name9734 (
		_w1566_,
		_w1602_,
		_w9751_,
		_w11083_,
		_w11084_
	);
	LUT4 #(
		.INIT('h00a8)
	) name9735 (
		\P2_EBX_reg[11]/NET0131 ,
		_w9752_,
		_w9765_,
		_w11084_,
		_w11085_
	);
	LUT3 #(
		.INIT('h6c)
	) name9736 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w9770_,
		_w11086_
	);
	LUT3 #(
		.INIT('h20)
	) name9737 (
		_w1673_,
		_w9786_,
		_w11086_,
		_w11087_
	);
	LUT4 #(
		.INIT('h2030)
	) name9738 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w11088_
	);
	LUT4 #(
		.INIT('h0200)
	) name9739 (
		_w1565_,
		_w1602_,
		_w1673_,
		_w11088_,
		_w11089_
	);
	LUT3 #(
		.INIT('h0d)
	) name9740 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w9788_,
		_w11089_,
		_w11090_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name9741 (
		_w1678_,
		_w11087_,
		_w11085_,
		_w11090_,
		_w11091_
	);
	LUT2 #(
		.INIT('h2)
	) name9742 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w9799_,
		_w11092_
	);
	LUT3 #(
		.INIT('h07)
	) name9743 (
		\P2_PhyAddrPointer_reg[11]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11093_
	);
	LUT2 #(
		.INIT('h4)
	) name9744 (
		_w11092_,
		_w11093_,
		_w11094_
	);
	LUT2 #(
		.INIT('h4)
	) name9745 (
		_w11091_,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('hb)
	) name9746 (
		_w11082_,
		_w11095_,
		_w11096_
	);
	LUT3 #(
		.INIT('h80)
	) name9747 (
		\P1_PhyAddrPointer_reg[24]/NET0131 ,
		_w6361_,
		_w11001_,
		_w11097_
	);
	LUT3 #(
		.INIT('h06)
	) name9748 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('h2)
	) name9749 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w11099_
	);
	LUT2 #(
		.INIT('h2)
	) name9750 (
		_w1939_,
		_w11099_,
		_w11100_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9751 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8164_,
		_w11098_,
		_w11100_,
		_w11101_
	);
	LUT4 #(
		.INIT('h1f0f)
	) name9752 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11030_,
		_w11102_
	);
	LUT3 #(
		.INIT('h12)
	) name9753 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1930_,
		_w11102_,
		_w11103_
	);
	LUT4 #(
		.INIT('h1333)
	) name9754 (
		\P1_rEIP_reg[24]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w10974_,
		_w11024_,
		_w11104_
	);
	LUT4 #(
		.INIT('h8000)
	) name9755 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		\P1_rEIP_reg[24]/NET0131 ,
		_w11105_
	);
	LUT4 #(
		.INIT('h8000)
	) name9756 (
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w11106_
	);
	LUT2 #(
		.INIT('h8)
	) name9757 (
		_w11105_,
		_w11106_,
		_w11107_
	);
	LUT3 #(
		.INIT('h80)
	) name9758 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w10858_,
		_w11107_,
		_w11108_
	);
	LUT4 #(
		.INIT('h444c)
	) name9759 (
		_w1930_,
		_w4709_,
		_w11104_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h2)
	) name9760 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w10808_,
		_w11110_
	);
	LUT4 #(
		.INIT('h3332)
	) name9761 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11111_
	);
	LUT3 #(
		.INIT('h02)
	) name9762 (
		_w1797_,
		_w1852_,
		_w11111_,
		_w11112_
	);
	LUT4 #(
		.INIT('h5700)
	) name9763 (
		_w10817_,
		_w11104_,
		_w11108_,
		_w11112_,
		_w11113_
	);
	LUT4 #(
		.INIT('h1011)
	) name9764 (
		_w11110_,
		_w11113_,
		_w11103_,
		_w11109_,
		_w11114_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9765 (
		\P1_PhyAddrPointer_reg[25]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11115_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name9766 (
		_w1933_,
		_w11114_,
		_w11101_,
		_w11115_,
		_w11116_
	);
	LUT4 #(
		.INIT('h8000)
	) name9767 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w5725_,
		_w5726_,
		_w9792_,
		_w11117_
	);
	LUT3 #(
		.INIT('h06)
	) name9768 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11117_,
		_w11118_
	);
	LUT2 #(
		.INIT('h2)
	) name9769 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w11119_
	);
	LUT2 #(
		.INIT('h2)
	) name9770 (
		_w1679_,
		_w11119_,
		_w11120_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9771 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8194_,
		_w11118_,
		_w11120_,
		_w11121_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9772 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[12]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11122_
	);
	LUT4 #(
		.INIT('h4888)
	) name9773 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w1673_,
		_w9771_,
		_w9770_,
		_w11123_
	);
	LUT3 #(
		.INIT('h23)
	) name9774 (
		_w1611_,
		_w11122_,
		_w11123_,
		_w11124_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9775 (
		\P2_EBX_reg[10]/NET0131 ,
		\P2_EBX_reg[11]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9755_,
		_w11125_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name9776 (
		\P2_EBX_reg[12]/NET0131 ,
		_w1673_,
		_w11123_,
		_w11125_,
		_w11126_
	);
	LUT4 #(
		.INIT('hf351)
	) name9777 (
		_w1565_,
		_w1566_,
		_w11124_,
		_w11126_,
		_w11127_
	);
	LUT4 #(
		.INIT('h5750)
	) name9778 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w1569_,
		_w1602_,
		_w11127_,
		_w11128_
	);
	LUT2 #(
		.INIT('h2)
	) name9779 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w9799_,
		_w11129_
	);
	LUT3 #(
		.INIT('h07)
	) name9780 (
		\P2_PhyAddrPointer_reg[12]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11130_
	);
	LUT2 #(
		.INIT('h4)
	) name9781 (
		_w11129_,
		_w11130_,
		_w11131_
	);
	LUT3 #(
		.INIT('hd0)
	) name9782 (
		_w1678_,
		_w11128_,
		_w11131_,
		_w11132_
	);
	LUT2 #(
		.INIT('hb)
	) name9783 (
		_w11121_,
		_w11132_,
		_w11133_
	);
	LUT2 #(
		.INIT('h8)
	) name9784 (
		_w8196_,
		_w9792_,
		_w11134_
	);
	LUT3 #(
		.INIT('h06)
	) name9785 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11134_,
		_w11135_
	);
	LUT2 #(
		.INIT('h2)
	) name9786 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w11136_
	);
	LUT2 #(
		.INIT('h2)
	) name9787 (
		_w1679_,
		_w11136_,
		_w11137_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9788 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8208_,
		_w11135_,
		_w11137_,
		_w11138_
	);
	LUT2 #(
		.INIT('h2)
	) name9789 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w9788_,
		_w11139_
	);
	LUT4 #(
		.INIT('h9500)
	) name9790 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9751_,
		_w11140_
	);
	LUT4 #(
		.INIT('h3332)
	) name9791 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[13]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11141_
	);
	LUT3 #(
		.INIT('h02)
	) name9792 (
		_w1566_,
		_w11141_,
		_w11140_,
		_w11142_
	);
	LUT4 #(
		.INIT('h0509)
	) name9793 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w9756_,
		_w11143_
	);
	LUT4 #(
		.INIT('h8444)
	) name9794 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w1673_,
		_w9770_,
		_w9772_,
		_w11144_
	);
	LUT3 #(
		.INIT('h02)
	) name9795 (
		_w1565_,
		_w11144_,
		_w11143_,
		_w11145_
	);
	LUT3 #(
		.INIT('h54)
	) name9796 (
		_w1602_,
		_w11142_,
		_w11145_,
		_w11146_
	);
	LUT2 #(
		.INIT('h2)
	) name9797 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w9799_,
		_w11147_
	);
	LUT3 #(
		.INIT('h07)
	) name9798 (
		\P2_PhyAddrPointer_reg[13]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11148_
	);
	LUT2 #(
		.INIT('h4)
	) name9799 (
		_w11147_,
		_w11148_,
		_w11149_
	);
	LUT4 #(
		.INIT('h5700)
	) name9800 (
		_w1678_,
		_w11139_,
		_w11146_,
		_w11149_,
		_w11150_
	);
	LUT2 #(
		.INIT('hb)
	) name9801 (
		_w11138_,
		_w11150_,
		_w11151_
	);
	LUT2 #(
		.INIT('h8)
	) name9802 (
		_w6362_,
		_w11001_,
		_w11152_
	);
	LUT4 #(
		.INIT('hf096)
	) name9803 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w7617_,
		_w11152_,
		_w11153_
	);
	LUT2 #(
		.INIT('h2)
	) name9804 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w11154_
	);
	LUT2 #(
		.INIT('h2)
	) name9805 (
		_w1939_,
		_w11154_,
		_w11155_
	);
	LUT3 #(
		.INIT('he0)
	) name9806 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w11153_,
		_w11155_,
		_w11156_
	);
	LUT2 #(
		.INIT('h1)
	) name9807 (
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		_w11157_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9808 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11030_,
		_w11157_,
		_w11158_
	);
	LUT4 #(
		.INIT('h8000)
	) name9809 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w10858_,
		_w11107_,
		_w11159_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name9810 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w10858_,
		_w11107_,
		_w11160_
	);
	LUT3 #(
		.INIT('hc4)
	) name9811 (
		_w1930_,
		_w4709_,
		_w11160_,
		_w11161_
	);
	LUT4 #(
		.INIT('hde00)
	) name9812 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1930_,
		_w11158_,
		_w11161_,
		_w11162_
	);
	LUT2 #(
		.INIT('h8)
	) name9813 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w10887_,
		_w11163_
	);
	LUT4 #(
		.INIT('h3222)
	) name9814 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w11164_
	);
	LUT4 #(
		.INIT('h000d)
	) name9815 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w11164_,
		_w11165_
	);
	LUT4 #(
		.INIT('ha200)
	) name9816 (
		\P1_EBX_reg[26]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w11166_
	);
	LUT3 #(
		.INIT('h08)
	) name9817 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w1842_,
		_w1851_,
		_w11167_
	);
	LUT2 #(
		.INIT('h1)
	) name9818 (
		_w11166_,
		_w11167_,
		_w11168_
	);
	LUT4 #(
		.INIT('h2f00)
	) name9819 (
		_w1930_,
		_w11160_,
		_w11165_,
		_w11168_,
		_w11169_
	);
	LUT3 #(
		.INIT('h31)
	) name9820 (
		_w1797_,
		_w11163_,
		_w11169_,
		_w11170_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9821 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		\P1_rEIP_reg[26]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11171_
	);
	LUT4 #(
		.INIT('h7500)
	) name9822 (
		_w1933_,
		_w11162_,
		_w11170_,
		_w11171_,
		_w11172_
	);
	LUT2 #(
		.INIT('hb)
	) name9823 (
		_w11156_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h8)
	) name9824 (
		_w5728_,
		_w11117_,
		_w11174_
	);
	LUT3 #(
		.INIT('h06)
	) name9825 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11174_,
		_w11175_
	);
	LUT2 #(
		.INIT('h2)
	) name9826 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w11176_
	);
	LUT2 #(
		.INIT('h2)
	) name9827 (
		_w1679_,
		_w11176_,
		_w11177_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9828 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8227_,
		_w11175_,
		_w11177_,
		_w11178_
	);
	LUT2 #(
		.INIT('h2)
	) name9829 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9788_,
		_w11179_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name9830 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w9770_,
		_w9772_,
		_w11180_
	);
	LUT2 #(
		.INIT('h2)
	) name9831 (
		_w9751_,
		_w11180_,
		_w11181_
	);
	LUT4 #(
		.INIT('h3332)
	) name9832 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11182_
	);
	LUT3 #(
		.INIT('h02)
	) name9833 (
		_w1566_,
		_w11182_,
		_w11181_,
		_w11183_
	);
	LUT3 #(
		.INIT('h8c)
	) name9834 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9756_,
		_w11184_
	);
	LUT3 #(
		.INIT('h21)
	) name9835 (
		\P2_EBX_reg[14]/NET0131 ,
		_w1673_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h2)
	) name9836 (
		_w1673_,
		_w11180_,
		_w11186_
	);
	LUT2 #(
		.INIT('h2)
	) name9837 (
		_w1565_,
		_w11186_,
		_w11187_
	);
	LUT4 #(
		.INIT('h4544)
	) name9838 (
		_w1602_,
		_w11183_,
		_w11185_,
		_w11187_,
		_w11188_
	);
	LUT2 #(
		.INIT('h2)
	) name9839 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w9799_,
		_w11189_
	);
	LUT3 #(
		.INIT('h07)
	) name9840 (
		\P2_PhyAddrPointer_reg[14]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11190_
	);
	LUT2 #(
		.INIT('h4)
	) name9841 (
		_w11189_,
		_w11190_,
		_w11191_
	);
	LUT4 #(
		.INIT('h5700)
	) name9842 (
		_w1678_,
		_w11179_,
		_w11188_,
		_w11191_,
		_w11192_
	);
	LUT2 #(
		.INIT('hb)
	) name9843 (
		_w11178_,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h8)
	) name9844 (
		_w5730_,
		_w9792_,
		_w11194_
	);
	LUT3 #(
		.INIT('h06)
	) name9845 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11194_,
		_w11195_
	);
	LUT2 #(
		.INIT('h2)
	) name9846 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w11196_
	);
	LUT2 #(
		.INIT('h2)
	) name9847 (
		_w1679_,
		_w11196_,
		_w11197_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9848 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7646_,
		_w11195_,
		_w11197_,
		_w11198_
	);
	LUT2 #(
		.INIT('h2)
	) name9849 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9788_,
		_w11199_
	);
	LUT4 #(
		.INIT('h3332)
	) name9850 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[15]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11200_
	);
	LUT2 #(
		.INIT('h2)
	) name9851 (
		_w1566_,
		_w11200_,
		_w11201_
	);
	LUT4 #(
		.INIT('he0f0)
	) name9852 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9756_,
		_w11202_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9853 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1565_,
		_w1673_,
		_w11202_,
		_w11203_
	);
	LUT4 #(
		.INIT('h8000)
	) name9854 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9773_,
		_w11204_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name9855 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9773_,
		_w11205_
	);
	LUT2 #(
		.INIT('h2)
	) name9856 (
		_w1673_,
		_w11205_,
		_w11206_
	);
	LUT4 #(
		.INIT('hf700)
	) name9857 (
		_w1566_,
		_w1611_,
		_w11200_,
		_w11206_,
		_w11207_
	);
	LUT4 #(
		.INIT('h0504)
	) name9858 (
		_w1602_,
		_w11201_,
		_w11207_,
		_w11203_,
		_w11208_
	);
	LUT2 #(
		.INIT('h2)
	) name9859 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9799_,
		_w11209_
	);
	LUT3 #(
		.INIT('h07)
	) name9860 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11210_
	);
	LUT2 #(
		.INIT('h4)
	) name9861 (
		_w11209_,
		_w11210_,
		_w11211_
	);
	LUT4 #(
		.INIT('h5700)
	) name9862 (
		_w1678_,
		_w11199_,
		_w11208_,
		_w11211_,
		_w11212_
	);
	LUT2 #(
		.INIT('hb)
	) name9863 (
		_w11198_,
		_w11212_,
		_w11213_
	);
	LUT3 #(
		.INIT('h80)
	) name9864 (
		\P1_PhyAddrPointer_reg[26]/NET0131 ,
		_w6362_,
		_w11001_,
		_w11214_
	);
	LUT3 #(
		.INIT('h06)
	) name9865 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11214_,
		_w11215_
	);
	LUT2 #(
		.INIT('h2)
	) name9866 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w11216_
	);
	LUT2 #(
		.INIT('h2)
	) name9867 (
		_w1939_,
		_w11216_,
		_w11217_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9868 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7025_,
		_w11215_,
		_w11217_,
		_w11218_
	);
	LUT3 #(
		.INIT('h01)
	) name9869 (
		\P1_EBX_reg[24]/NET0131 ,
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		_w11219_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9870 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11030_,
		_w11219_,
		_w11220_
	);
	LUT4 #(
		.INIT('h70b0)
	) name9871 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w1930_,
		_w4709_,
		_w11159_,
		_w11221_
	);
	LUT4 #(
		.INIT('hde00)
	) name9872 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1930_,
		_w11220_,
		_w11221_,
		_w11222_
	);
	LUT2 #(
		.INIT('h8)
	) name9873 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w10887_,
		_w11223_
	);
	LUT4 #(
		.INIT('h3222)
	) name9874 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w11224_
	);
	LUT4 #(
		.INIT('h000d)
	) name9875 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w11224_,
		_w11225_
	);
	LUT4 #(
		.INIT('h7b00)
	) name9876 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w1930_,
		_w11159_,
		_w11225_,
		_w11226_
	);
	LUT4 #(
		.INIT('ha200)
	) name9877 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w11227_
	);
	LUT3 #(
		.INIT('h08)
	) name9878 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w1842_,
		_w1851_,
		_w11228_
	);
	LUT2 #(
		.INIT('h1)
	) name9879 (
		_w11227_,
		_w11228_,
		_w11229_
	);
	LUT4 #(
		.INIT('h1311)
	) name9880 (
		_w1797_,
		_w11223_,
		_w11226_,
		_w11229_,
		_w11230_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9881 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11231_
	);
	LUT4 #(
		.INIT('h7500)
	) name9882 (
		_w1933_,
		_w11222_,
		_w11230_,
		_w11231_,
		_w11232_
	);
	LUT2 #(
		.INIT('hb)
	) name9883 (
		_w11218_,
		_w11232_,
		_w11233_
	);
	LUT3 #(
		.INIT('h80)
	) name9884 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		_w5730_,
		_w9792_,
		_w11234_
	);
	LUT3 #(
		.INIT('h06)
	) name9885 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11234_,
		_w11235_
	);
	LUT2 #(
		.INIT('h2)
	) name9886 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w11236_
	);
	LUT2 #(
		.INIT('h2)
	) name9887 (
		_w1679_,
		_w11236_,
		_w11237_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9888 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8244_,
		_w11235_,
		_w11237_,
		_w11238_
	);
	LUT2 #(
		.INIT('h2)
	) name9889 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9788_,
		_w11239_
	);
	LUT4 #(
		.INIT('h3332)
	) name9890 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[16]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11240_
	);
	LUT2 #(
		.INIT('h2)
	) name9891 (
		_w1566_,
		_w11240_,
		_w11241_
	);
	LUT4 #(
		.INIT('h0100)
	) name9892 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		\P2_EBX_reg[15]/NET0131 ,
		_w9756_,
		_w11242_
	);
	LUT4 #(
		.INIT('h0509)
	) name9893 (
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w11242_,
		_w11243_
	);
	LUT3 #(
		.INIT('h31)
	) name9894 (
		_w1565_,
		_w11241_,
		_w11243_,
		_w11244_
	);
	LUT3 #(
		.INIT('h80)
	) name9895 (
		_w9770_,
		_w9772_,
		_w9775_,
		_w11245_
	);
	LUT4 #(
		.INIT('hcc04)
	) name9896 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w1673_,
		_w11204_,
		_w11245_,
		_w11246_
	);
	LUT4 #(
		.INIT('hf700)
	) name9897 (
		_w1566_,
		_w1611_,
		_w11240_,
		_w11246_,
		_w11247_
	);
	LUT2 #(
		.INIT('h1)
	) name9898 (
		_w1602_,
		_w11247_,
		_w11248_
	);
	LUT4 #(
		.INIT('h8a88)
	) name9899 (
		_w1678_,
		_w11239_,
		_w11244_,
		_w11248_,
		_w11249_
	);
	LUT2 #(
		.INIT('h2)
	) name9900 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9799_,
		_w11250_
	);
	LUT3 #(
		.INIT('h07)
	) name9901 (
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11251_
	);
	LUT2 #(
		.INIT('h4)
	) name9902 (
		_w11250_,
		_w11251_,
		_w11252_
	);
	LUT2 #(
		.INIT('h4)
	) name9903 (
		_w11249_,
		_w11252_,
		_w11253_
	);
	LUT2 #(
		.INIT('hb)
	) name9904 (
		_w11238_,
		_w11253_,
		_w11254_
	);
	LUT4 #(
		.INIT('h8000)
	) name9905 (
		\P2_PhyAddrPointer_reg[15]/NET0131 ,
		\P2_PhyAddrPointer_reg[16]/NET0131 ,
		_w5730_,
		_w9792_,
		_w11255_
	);
	LUT3 #(
		.INIT('h06)
	) name9906 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h2)
	) name9907 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w11257_
	);
	LUT2 #(
		.INIT('h2)
	) name9908 (
		_w1679_,
		_w11257_,
		_w11258_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9909 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8258_,
		_w11256_,
		_w11258_,
		_w11259_
	);
	LUT4 #(
		.INIT('hfb01)
	) name9910 (
		_w1565_,
		_w1566_,
		_w1568_,
		_w1602_,
		_w11260_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name9911 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9775_,
		_w11261_
	);
	LUT3 #(
		.INIT('h40)
	) name9912 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1612_,
		_w11261_,
		_w11262_
	);
	LUT4 #(
		.INIT('hccc8)
	) name9913 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[17]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11263_
	);
	LUT3 #(
		.INIT('h0d)
	) name9914 (
		_w1592_,
		_w1601_,
		_w11263_,
		_w11264_
	);
	LUT2 #(
		.INIT('h4)
	) name9915 (
		_w11262_,
		_w11264_,
		_w11265_
	);
	LUT2 #(
		.INIT('h2)
	) name9916 (
		_w1566_,
		_w11265_,
		_w11266_
	);
	LUT3 #(
		.INIT('ha8)
	) name9917 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w11260_,
		_w11266_,
		_w11267_
	);
	LUT3 #(
		.INIT('h8c)
	) name9918 (
		\P2_EBX_reg[16]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11242_,
		_w11268_
	);
	LUT3 #(
		.INIT('h10)
	) name9919 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1605_,
		_w11261_,
		_w11269_
	);
	LUT4 #(
		.INIT('h00ed)
	) name9920 (
		\P2_EBX_reg[17]/NET0131 ,
		_w1673_,
		_w11268_,
		_w11269_,
		_w11270_
	);
	LUT4 #(
		.INIT('h3032)
	) name9921 (
		_w1565_,
		_w1602_,
		_w11266_,
		_w11270_,
		_w11271_
	);
	LUT2 #(
		.INIT('h2)
	) name9922 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w9799_,
		_w11272_
	);
	LUT3 #(
		.INIT('h07)
	) name9923 (
		\P2_PhyAddrPointer_reg[17]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11273_
	);
	LUT2 #(
		.INIT('h4)
	) name9924 (
		_w11272_,
		_w11273_,
		_w11274_
	);
	LUT4 #(
		.INIT('h5700)
	) name9925 (
		_w1678_,
		_w11267_,
		_w11271_,
		_w11274_,
		_w11275_
	);
	LUT2 #(
		.INIT('hb)
	) name9926 (
		_w11259_,
		_w11275_,
		_w11276_
	);
	LUT4 #(
		.INIT('h8000)
	) name9927 (
		\P1_PhyAddrPointer_reg[27]/NET0131 ,
		_w6362_,
		_w6380_,
		_w11001_,
		_w11277_
	);
	LUT3 #(
		.INIT('h06)
	) name9928 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11277_,
		_w11278_
	);
	LUT2 #(
		.INIT('h2)
	) name9929 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w11279_
	);
	LUT2 #(
		.INIT('h2)
	) name9930 (
		_w1939_,
		_w11279_,
		_w11280_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9931 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7039_,
		_w11278_,
		_w11280_,
		_w11281_
	);
	LUT4 #(
		.INIT('h1000)
	) name9932 (
		\P1_EBX_reg[23]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w11030_,
		_w11219_,
		_w11282_
	);
	LUT4 #(
		.INIT('h0509)
	) name9933 (
		\P1_EBX_reg[28]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w11282_,
		_w11283_
	);
	LUT4 #(
		.INIT('h9030)
	) name9934 (
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w1930_,
		_w11159_,
		_w11284_
	);
	LUT2 #(
		.INIT('h2)
	) name9935 (
		_w4709_,
		_w11284_,
		_w11285_
	);
	LUT2 #(
		.INIT('h2)
	) name9936 (
		\P1_rEIP_reg[28]/NET0131 ,
		_w10808_,
		_w11286_
	);
	LUT4 #(
		.INIT('h3332)
	) name9937 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[28]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11287_
	);
	LUT3 #(
		.INIT('h02)
	) name9938 (
		_w1797_,
		_w1852_,
		_w11287_,
		_w11288_
	);
	LUT4 #(
		.INIT('h1033)
	) name9939 (
		_w1858_,
		_w11286_,
		_w11284_,
		_w11288_,
		_w11289_
	);
	LUT4 #(
		.INIT('h20aa)
	) name9940 (
		_w1933_,
		_w11283_,
		_w11285_,
		_w11289_,
		_w11290_
	);
	LUT4 #(
		.INIT('h5f13)
	) name9941 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11291_
	);
	LUT3 #(
		.INIT('hef)
	) name9942 (
		_w11290_,
		_w11281_,
		_w11291_,
		_w11292_
	);
	LUT3 #(
		.INIT('h06)
	) name9943 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9793_,
		_w11293_
	);
	LUT2 #(
		.INIT('h2)
	) name9944 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		_w11294_
	);
	LUT2 #(
		.INIT('h2)
	) name9945 (
		_w1679_,
		_w11294_,
		_w11295_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9946 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8269_,
		_w11293_,
		_w11295_,
		_w11296_
	);
	LUT2 #(
		.INIT('h2)
	) name9947 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w9788_,
		_w11297_
	);
	LUT4 #(
		.INIT('h3332)
	) name9948 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11298_
	);
	LUT2 #(
		.INIT('h2)
	) name9949 (
		_w1566_,
		_w11298_,
		_w11299_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name9950 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9756_,
		_w9757_,
		_w11300_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name9951 (
		\P2_EBX_reg[18]/NET0131 ,
		_w1565_,
		_w1673_,
		_w11300_,
		_w11301_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name9952 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9776_,
		_w11302_
	);
	LUT2 #(
		.INIT('h2)
	) name9953 (
		_w1673_,
		_w11302_,
		_w11303_
	);
	LUT4 #(
		.INIT('hf700)
	) name9954 (
		_w1566_,
		_w1611_,
		_w11298_,
		_w11303_,
		_w11304_
	);
	LUT4 #(
		.INIT('h0504)
	) name9955 (
		_w1602_,
		_w11299_,
		_w11304_,
		_w11301_,
		_w11305_
	);
	LUT2 #(
		.INIT('h2)
	) name9956 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w9799_,
		_w11306_
	);
	LUT3 #(
		.INIT('h07)
	) name9957 (
		\P2_PhyAddrPointer_reg[18]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11307_
	);
	LUT2 #(
		.INIT('h4)
	) name9958 (
		_w11306_,
		_w11307_,
		_w11308_
	);
	LUT4 #(
		.INIT('h5700)
	) name9959 (
		_w1678_,
		_w11297_,
		_w11305_,
		_w11308_,
		_w11309_
	);
	LUT2 #(
		.INIT('hb)
	) name9960 (
		_w11296_,
		_w11309_,
		_w11310_
	);
	LUT4 #(
		.INIT('heda5)
	) name9961 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5732_,
		_w5745_,
		_w9793_,
		_w11311_
	);
	LUT2 #(
		.INIT('h2)
	) name9962 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w11312_
	);
	LUT2 #(
		.INIT('h2)
	) name9963 (
		_w1679_,
		_w11312_,
		_w11313_
	);
	LUT4 #(
		.INIT('heb00)
	) name9964 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7661_,
		_w11311_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h2)
	) name9965 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9788_,
		_w11315_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name9966 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9770_,
		_w9772_,
		_w9777_,
		_w11316_
	);
	LUT2 #(
		.INIT('h2)
	) name9967 (
		_w9751_,
		_w11316_,
		_w11317_
	);
	LUT4 #(
		.INIT('h3332)
	) name9968 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[19]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11318_
	);
	LUT3 #(
		.INIT('h02)
	) name9969 (
		_w1566_,
		_w11318_,
		_w11317_,
		_w11319_
	);
	LUT4 #(
		.INIT('h1000)
	) name9970 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w9756_,
		_w9757_,
		_w11320_
	);
	LUT4 #(
		.INIT('h0509)
	) name9971 (
		\P2_EBX_reg[19]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w11320_,
		_w11321_
	);
	LUT2 #(
		.INIT('h2)
	) name9972 (
		_w1673_,
		_w11316_,
		_w11322_
	);
	LUT2 #(
		.INIT('h2)
	) name9973 (
		_w1565_,
		_w11322_,
		_w11323_
	);
	LUT4 #(
		.INIT('h4544)
	) name9974 (
		_w1602_,
		_w11319_,
		_w11321_,
		_w11323_,
		_w11324_
	);
	LUT2 #(
		.INIT('h2)
	) name9975 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w9799_,
		_w11325_
	);
	LUT3 #(
		.INIT('h07)
	) name9976 (
		\P2_PhyAddrPointer_reg[19]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11326_
	);
	LUT2 #(
		.INIT('h4)
	) name9977 (
		_w11325_,
		_w11326_,
		_w11327_
	);
	LUT4 #(
		.INIT('h5700)
	) name9978 (
		_w1678_,
		_w11315_,
		_w11324_,
		_w11327_,
		_w11328_
	);
	LUT2 #(
		.INIT('hb)
	) name9979 (
		_w11314_,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h1)
	) name9980 (
		\P1_EBX_reg[27]/NET0131 ,
		\P1_EBX_reg[28]/NET0131 ,
		_w11330_
	);
	LUT4 #(
		.INIT('h4000)
	) name9981 (
		\P1_EBX_reg[23]/NET0131 ,
		_w11030_,
		_w11219_,
		_w11330_,
		_w11331_
	);
	LUT4 #(
		.INIT('h0509)
	) name9982 (
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w11331_,
		_w11332_
	);
	LUT4 #(
		.INIT('h8000)
	) name9983 (
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w11159_,
		_w11333_
	);
	LUT4 #(
		.INIT('h78f0)
	) name9984 (
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w11159_,
		_w11334_
	);
	LUT3 #(
		.INIT('hc4)
	) name9985 (
		_w1930_,
		_w4709_,
		_w11334_,
		_w11335_
	);
	LUT2 #(
		.INIT('h4)
	) name9986 (
		_w11332_,
		_w11335_,
		_w11336_
	);
	LUT4 #(
		.INIT('h3222)
	) name9987 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[29]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w11337_
	);
	LUT4 #(
		.INIT('h000d)
	) name9988 (
		_w1842_,
		_w1851_,
		_w1858_,
		_w11337_,
		_w11338_
	);
	LUT4 #(
		.INIT('ha200)
	) name9989 (
		\P1_EBX_reg[29]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1858_,
		_w11339_
	);
	LUT3 #(
		.INIT('h08)
	) name9990 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w1842_,
		_w1851_,
		_w11340_
	);
	LUT2 #(
		.INIT('h1)
	) name9991 (
		_w11339_,
		_w11340_,
		_w11341_
	);
	LUT4 #(
		.INIT('h2f00)
	) name9992 (
		_w1930_,
		_w11334_,
		_w11338_,
		_w11341_,
		_w11342_
	);
	LUT2 #(
		.INIT('h8)
	) name9993 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w10887_,
		_w11343_
	);
	LUT3 #(
		.INIT('h0d)
	) name9994 (
		_w1797_,
		_w11342_,
		_w11343_,
		_w11344_
	);
	LUT3 #(
		.INIT('h8a)
	) name9995 (
		_w1933_,
		_w11336_,
		_w11344_,
		_w11345_
	);
	LUT4 #(
		.INIT('h143c)
	) name9996 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11277_,
		_w11346_
	);
	LUT2 #(
		.INIT('h2)
	) name9997 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w11347_
	);
	LUT2 #(
		.INIT('h2)
	) name9998 (
		_w1939_,
		_w11347_,
		_w11348_
	);
	LUT4 #(
		.INIT('hbe00)
	) name9999 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7051_,
		_w11346_,
		_w11348_,
		_w11349_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10000 (
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11350_
	);
	LUT2 #(
		.INIT('h4)
	) name10001 (
		_w11349_,
		_w11350_,
		_w11351_
	);
	LUT2 #(
		.INIT('hb)
	) name10002 (
		_w11345_,
		_w11351_,
		_w11352_
	);
	LUT3 #(
		.INIT('h28)
	) name10003 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11353_
	);
	LUT2 #(
		.INIT('h2)
	) name10004 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w11354_
	);
	LUT2 #(
		.INIT('h2)
	) name10005 (
		_w1679_,
		_w11354_,
		_w11355_
	);
	LUT4 #(
		.INIT('heb00)
	) name10006 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w11353_,
		_w11355_,
		_w11356_
	);
	LUT2 #(
		.INIT('h2)
	) name10007 (
		\P2_rEIP_reg[1]/NET0131 ,
		_w9788_,
		_w11357_
	);
	LUT2 #(
		.INIT('h6)
	) name10008 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		_w11358_
	);
	LUT3 #(
		.INIT('h90)
	) name10009 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11359_
	);
	LUT2 #(
		.INIT('h1)
	) name10010 (
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11360_
	);
	LUT2 #(
		.INIT('h1)
	) name10011 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w11361_
	);
	LUT4 #(
		.INIT('h0111)
	) name10012 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w11362_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10013 (
		_w1673_,
		_w11360_,
		_w11359_,
		_w11362_,
		_w11363_
	);
	LUT2 #(
		.INIT('h2)
	) name10014 (
		_w1565_,
		_w11363_,
		_w11364_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10015 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11365_
	);
	LUT3 #(
		.INIT('h10)
	) name10016 (
		_w1605_,
		_w1611_,
		_w11361_,
		_w11366_
	);
	LUT2 #(
		.INIT('h1)
	) name10017 (
		_w11365_,
		_w11366_,
		_w11367_
	);
	LUT4 #(
		.INIT('hf351)
	) name10018 (
		_w1566_,
		_w1568_,
		_w1646_,
		_w11367_,
		_w11368_
	);
	LUT3 #(
		.INIT('h45)
	) name10019 (
		_w1602_,
		_w11364_,
		_w11368_,
		_w11369_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10020 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11370_
	);
	LUT4 #(
		.INIT('h5700)
	) name10021 (
		_w1678_,
		_w11357_,
		_w11369_,
		_w11370_,
		_w11371_
	);
	LUT2 #(
		.INIT('hb)
	) name10022 (
		_w11356_,
		_w11371_,
		_w11372_
	);
	LUT3 #(
		.INIT('h80)
	) name10023 (
		_w5733_,
		_w8260_,
		_w9792_,
		_w11373_
	);
	LUT3 #(
		.INIT('h06)
	) name10024 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11373_,
		_w11374_
	);
	LUT2 #(
		.INIT('h2)
	) name10025 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w11375_
	);
	LUT2 #(
		.INIT('h2)
	) name10026 (
		_w1679_,
		_w11375_,
		_w11376_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10027 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7373_,
		_w11374_,
		_w11376_,
		_w11377_
	);
	LUT4 #(
		.INIT('h1040)
	) name10028 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w1612_,
		_w9778_,
		_w11378_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10029 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[20]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11379_
	);
	LUT3 #(
		.INIT('h0d)
	) name10030 (
		_w1592_,
		_w1601_,
		_w11379_,
		_w11380_
	);
	LUT2 #(
		.INIT('h4)
	) name10031 (
		_w11378_,
		_w11380_,
		_w11381_
	);
	LUT2 #(
		.INIT('h2)
	) name10032 (
		_w1566_,
		_w11381_,
		_w11382_
	);
	LUT3 #(
		.INIT('ha8)
	) name10033 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w11260_,
		_w11382_,
		_w11383_
	);
	LUT4 #(
		.INIT('h0a06)
	) name10034 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w9759_,
		_w11384_
	);
	LUT4 #(
		.INIT('h0104)
	) name10035 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w1605_,
		_w9778_,
		_w11385_
	);
	LUT4 #(
		.INIT('h1113)
	) name10036 (
		_w1565_,
		_w11382_,
		_w11384_,
		_w11385_,
		_w11386_
	);
	LUT4 #(
		.INIT('hc0c4)
	) name10037 (
		_w1602_,
		_w1678_,
		_w11383_,
		_w11386_,
		_w11387_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10038 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11388_
	);
	LUT2 #(
		.INIT('h4)
	) name10039 (
		_w11387_,
		_w11388_,
		_w11389_
	);
	LUT2 #(
		.INIT('hb)
	) name10040 (
		_w11377_,
		_w11389_,
		_w11390_
	);
	LUT4 #(
		.INIT('h8000)
	) name10041 (
		\P2_PhyAddrPointer_reg[20]/NET0131 ,
		_w5733_,
		_w8260_,
		_w9792_,
		_w11391_
	);
	LUT3 #(
		.INIT('h06)
	) name10042 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11391_,
		_w11392_
	);
	LUT2 #(
		.INIT('h2)
	) name10043 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w11393_
	);
	LUT2 #(
		.INIT('h2)
	) name10044 (
		_w1679_,
		_w11393_,
		_w11394_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10045 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7913_,
		_w11392_,
		_w11394_,
		_w11395_
	);
	LUT2 #(
		.INIT('h2)
	) name10046 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w9788_,
		_w11396_
	);
	LUT4 #(
		.INIT('h3332)
	) name10047 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11397_
	);
	LUT3 #(
		.INIT('h02)
	) name10048 (
		_w1566_,
		_w1602_,
		_w11397_,
		_w11398_
	);
	LUT3 #(
		.INIT('h8c)
	) name10049 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9759_,
		_w11399_
	);
	LUT4 #(
		.INIT('hd0e0)
	) name10050 (
		\P2_EBX_reg[21]/NET0131 ,
		_w1673_,
		_w6439_,
		_w11399_,
		_w11400_
	);
	LUT4 #(
		.INIT('h0020)
	) name10051 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w11397_,
		_w11401_
	);
	LUT4 #(
		.INIT('h9030)
	) name10052 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w1673_,
		_w9778_,
		_w11402_
	);
	LUT2 #(
		.INIT('h4)
	) name10053 (
		_w11401_,
		_w11402_,
		_w11403_
	);
	LUT4 #(
		.INIT('h5501)
	) name10054 (
		_w11396_,
		_w11398_,
		_w11400_,
		_w11403_,
		_w11404_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10055 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11405_
	);
	LUT3 #(
		.INIT('hd0)
	) name10056 (
		_w1678_,
		_w11404_,
		_w11405_,
		_w11406_
	);
	LUT2 #(
		.INIT('hb)
	) name10057 (
		_w11395_,
		_w11406_,
		_w11407_
	);
	LUT2 #(
		.INIT('h6)
	) name10058 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w11408_
	);
	LUT4 #(
		.INIT('hf906)
	) name10059 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10801_,
		_w11408_,
		_w11409_
	);
	LUT2 #(
		.INIT('h2)
	) name10060 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w11410_
	);
	LUT2 #(
		.INIT('h2)
	) name10061 (
		_w1939_,
		_w11410_,
		_w11411_
	);
	LUT2 #(
		.INIT('h2)
	) name10062 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w10808_,
		_w11412_
	);
	LUT3 #(
		.INIT('h14)
	) name10063 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w11413_
	);
	LUT2 #(
		.INIT('h4)
	) name10064 (
		_w1861_,
		_w11413_,
		_w11414_
	);
	LUT3 #(
		.INIT('he0)
	) name10065 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11415_
	);
	LUT3 #(
		.INIT('h12)
	) name10066 (
		\P1_EBX_reg[2]/NET0131 ,
		_w1930_,
		_w11415_,
		_w11416_
	);
	LUT2 #(
		.INIT('h1)
	) name10067 (
		_w11414_,
		_w11416_,
		_w11417_
	);
	LUT3 #(
		.INIT('h02)
	) name10068 (
		_w1795_,
		_w1852_,
		_w11417_,
		_w11418_
	);
	LUT3 #(
		.INIT('h08)
	) name10069 (
		_w1802_,
		_w1895_,
		_w1852_,
		_w11419_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10070 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11420_
	);
	LUT3 #(
		.INIT('h10)
	) name10071 (
		_w1858_,
		_w1861_,
		_w11413_,
		_w11421_
	);
	LUT2 #(
		.INIT('h1)
	) name10072 (
		_w11420_,
		_w11421_,
		_w11422_
	);
	LUT3 #(
		.INIT('h02)
	) name10073 (
		_w1797_,
		_w1852_,
		_w11422_,
		_w11423_
	);
	LUT3 #(
		.INIT('h01)
	) name10074 (
		_w11419_,
		_w11423_,
		_w11418_,
		_w11424_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10075 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11425_
	);
	LUT4 #(
		.INIT('h7500)
	) name10076 (
		_w1933_,
		_w11412_,
		_w11424_,
		_w11425_,
		_w11426_
	);
	LUT4 #(
		.INIT('he0ff)
	) name10077 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w11409_,
		_w11411_,
		_w11426_,
		_w11427_
	);
	LUT2 #(
		.INIT('h8)
	) name10078 (
		\P2_PhyAddrPointer_reg[21]/NET0131 ,
		_w11391_,
		_w11428_
	);
	LUT3 #(
		.INIT('h06)
	) name10079 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h2)
	) name10080 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w11430_
	);
	LUT2 #(
		.INIT('h2)
	) name10081 (
		_w1679_,
		_w11430_,
		_w11431_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10082 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7385_,
		_w11429_,
		_w11431_,
		_w11432_
	);
	LUT2 #(
		.INIT('h2)
	) name10083 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w9788_,
		_w11433_
	);
	LUT4 #(
		.INIT('h3332)
	) name10084 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11434_
	);
	LUT2 #(
		.INIT('h2)
	) name10085 (
		_w1566_,
		_w11434_,
		_w11435_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10086 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9759_,
		_w11436_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name10087 (
		\P2_EBX_reg[22]/NET0131 ,
		_w1565_,
		_w1673_,
		_w11436_,
		_w11437_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10088 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w9778_,
		_w11438_
	);
	LUT4 #(
		.INIT('hf070)
	) name10089 (
		_w1566_,
		_w1611_,
		_w1673_,
		_w11434_,
		_w11439_
	);
	LUT3 #(
		.INIT('h45)
	) name10090 (
		_w1602_,
		_w11438_,
		_w11439_,
		_w11440_
	);
	LUT4 #(
		.INIT('h0155)
	) name10091 (
		_w11433_,
		_w11435_,
		_w11437_,
		_w11440_,
		_w11441_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10092 (
		\P2_PhyAddrPointer_reg[22]/NET0131 ,
		\P2_rEIP_reg[22]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11442_
	);
	LUT3 #(
		.INIT('hd0)
	) name10093 (
		_w1678_,
		_w11441_,
		_w11442_,
		_w11443_
	);
	LUT2 #(
		.INIT('hb)
	) name10094 (
		_w11432_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h8)
	) name10095 (
		_w5734_,
		_w11391_,
		_w11445_
	);
	LUT3 #(
		.INIT('h06)
	) name10096 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11445_,
		_w11446_
	);
	LUT2 #(
		.INIT('h2)
	) name10097 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w11447_
	);
	LUT2 #(
		.INIT('h2)
	) name10098 (
		_w1679_,
		_w11447_,
		_w11448_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10099 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6861_,
		_w11446_,
		_w11448_,
		_w11449_
	);
	LUT2 #(
		.INIT('h2)
	) name10100 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9788_,
		_w11450_
	);
	LUT4 #(
		.INIT('h3332)
	) name10101 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11451_
	);
	LUT3 #(
		.INIT('h02)
	) name10102 (
		_w1566_,
		_w1602_,
		_w11451_,
		_w11452_
	);
	LUT4 #(
		.INIT('h0100)
	) name10103 (
		\P2_EBX_reg[20]/NET0131 ,
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		_w9759_,
		_w11453_
	);
	LUT4 #(
		.INIT('h0509)
	) name10104 (
		\P2_EBX_reg[23]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w11453_,
		_w11454_
	);
	LUT2 #(
		.INIT('h6)
	) name10105 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9780_,
		_w11455_
	);
	LUT4 #(
		.INIT('h0800)
	) name10106 (
		\P2_EBX_reg[23]/NET0131 ,
		_w1566_,
		_w1602_,
		_w1611_,
		_w11456_
	);
	LUT3 #(
		.INIT('h02)
	) name10107 (
		_w1673_,
		_w11456_,
		_w11455_,
		_w11457_
	);
	LUT4 #(
		.INIT('h00ce)
	) name10108 (
		_w6439_,
		_w11452_,
		_w11454_,
		_w11457_,
		_w11458_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10109 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11459_
	);
	LUT4 #(
		.INIT('h5700)
	) name10110 (
		_w1678_,
		_w11450_,
		_w11458_,
		_w11459_,
		_w11460_
	);
	LUT2 #(
		.INIT('hb)
	) name10111 (
		_w11449_,
		_w11460_,
		_w11461_
	);
	LUT4 #(
		.INIT('hebc3)
	) name10112 (
		\P2_PhyAddrPointer_reg[23]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11445_,
		_w11462_
	);
	LUT2 #(
		.INIT('h2)
	) name10113 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w11463_
	);
	LUT2 #(
		.INIT('h2)
	) name10114 (
		_w1679_,
		_w11463_,
		_w11464_
	);
	LUT4 #(
		.INIT('heb00)
	) name10115 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7403_,
		_w11462_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h2)
	) name10116 (
		\P2_rEIP_reg[24]/NET0131 ,
		_w9788_,
		_w11466_
	);
	LUT4 #(
		.INIT('h00a8)
	) name10117 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w11467_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10118 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9465_,
		_w9761_,
		_w11467_,
		_w11468_
	);
	LUT3 #(
		.INIT('h04)
	) name10119 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1565_,
		_w1602_,
		_w11469_
	);
	LUT3 #(
		.INIT('h20)
	) name10120 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9761_,
		_w11469_,
		_w11470_
	);
	LUT3 #(
		.INIT('h6c)
	) name10121 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w9780_,
		_w11471_
	);
	LUT4 #(
		.INIT('h0800)
	) name10122 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1566_,
		_w1602_,
		_w1611_,
		_w11472_
	);
	LUT3 #(
		.INIT('h02)
	) name10123 (
		_w1673_,
		_w11472_,
		_w11471_,
		_w11473_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10124 (
		_w9787_,
		_w11470_,
		_w11468_,
		_w11473_,
		_w11474_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10125 (
		\P2_PhyAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11475_
	);
	LUT4 #(
		.INIT('h5700)
	) name10126 (
		_w1678_,
		_w11466_,
		_w11474_,
		_w11475_,
		_w11476_
	);
	LUT2 #(
		.INIT('hb)
	) name10127 (
		_w11465_,
		_w11476_,
		_w11477_
	);
	LUT3 #(
		.INIT('h06)
	) name10128 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9794_,
		_w11478_
	);
	LUT2 #(
		.INIT('h2)
	) name10129 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w11479_
	);
	LUT2 #(
		.INIT('h2)
	) name10130 (
		_w1679_,
		_w11479_,
		_w11480_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10131 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7922_,
		_w11478_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h2)
	) name10132 (
		\P2_rEIP_reg[25]/NET0131 ,
		_w9788_,
		_w11482_
	);
	LUT4 #(
		.INIT('h3332)
	) name10133 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[25]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11483_
	);
	LUT3 #(
		.INIT('h02)
	) name10134 (
		_w1566_,
		_w1602_,
		_w11483_,
		_w11484_
	);
	LUT3 #(
		.INIT('h8c)
	) name10135 (
		\P2_EBX_reg[24]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9761_,
		_w11485_
	);
	LUT4 #(
		.INIT('hd0e0)
	) name10136 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1673_,
		_w6439_,
		_w11485_,
		_w11486_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10137 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w9780_,
		_w11487_
	);
	LUT4 #(
		.INIT('h0800)
	) name10138 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1566_,
		_w1602_,
		_w1611_,
		_w11488_
	);
	LUT3 #(
		.INIT('h02)
	) name10139 (
		_w1673_,
		_w11488_,
		_w11487_,
		_w11489_
	);
	LUT4 #(
		.INIT('h5501)
	) name10140 (
		_w11482_,
		_w11484_,
		_w11486_,
		_w11489_,
		_w11490_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10141 (
		\P2_PhyAddrPointer_reg[25]/NET0131 ,
		\P2_rEIP_reg[25]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11491_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name10142 (
		_w1678_,
		_w11490_,
		_w11481_,
		_w11491_,
		_w11492_
	);
	LUT3 #(
		.INIT('h40)
	) name10143 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w11493_
	);
	LUT3 #(
		.INIT('h06)
	) name10144 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11493_,
		_w11494_
	);
	LUT2 #(
		.INIT('h2)
	) name10145 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w11495_
	);
	LUT2 #(
		.INIT('h2)
	) name10146 (
		_w1939_,
		_w11495_,
		_w11496_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10147 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w9623_,
		_w11494_,
		_w11496_,
		_w11497_
	);
	LUT2 #(
		.INIT('h2)
	) name10148 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w10808_,
		_w11498_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10149 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11499_
	);
	LUT4 #(
		.INIT('h1540)
	) name10150 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w11500_
	);
	LUT3 #(
		.INIT('h10)
	) name10151 (
		_w1858_,
		_w1861_,
		_w11500_,
		_w11501_
	);
	LUT2 #(
		.INIT('h1)
	) name10152 (
		_w11499_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h2)
	) name10153 (
		_w1797_,
		_w11502_,
		_w11503_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10154 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11504_
	);
	LUT3 #(
		.INIT('h12)
	) name10155 (
		\P1_EBX_reg[3]/NET0131 ,
		_w1930_,
		_w11504_,
		_w11505_
	);
	LUT2 #(
		.INIT('h4)
	) name10156 (
		_w1861_,
		_w11500_,
		_w11506_
	);
	LUT2 #(
		.INIT('h1)
	) name10157 (
		_w11505_,
		_w11506_,
		_w11507_
	);
	LUT4 #(
		.INIT('hf351)
	) name10158 (
		_w1795_,
		_w1802_,
		_w1883_,
		_w11507_,
		_w11508_
	);
	LUT3 #(
		.INIT('h45)
	) name10159 (
		_w1852_,
		_w11503_,
		_w11508_,
		_w11509_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10160 (
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		_w2234_,
		_w10828_,
		_w11510_
	);
	LUT4 #(
		.INIT('h5700)
	) name10161 (
		_w1933_,
		_w11498_,
		_w11509_,
		_w11510_,
		_w11511_
	);
	LUT2 #(
		.INIT('hb)
	) name10162 (
		_w11497_,
		_w11511_,
		_w11512_
	);
	LUT4 #(
		.INIT('hf096)
	) name10163 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w7413_,
		_w9795_,
		_w11513_
	);
	LUT2 #(
		.INIT('h2)
	) name10164 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w11514_
	);
	LUT2 #(
		.INIT('h2)
	) name10165 (
		_w1679_,
		_w11514_,
		_w11515_
	);
	LUT3 #(
		.INIT('he0)
	) name10166 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w11513_,
		_w11515_,
		_w11516_
	);
	LUT2 #(
		.INIT('h2)
	) name10167 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9788_,
		_w11517_
	);
	LUT4 #(
		.INIT('h3332)
	) name10168 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[26]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11518_
	);
	LUT3 #(
		.INIT('h02)
	) name10169 (
		_w1566_,
		_w1602_,
		_w11518_,
		_w11519_
	);
	LUT3 #(
		.INIT('h2a)
	) name10170 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9761_,
		_w9762_,
		_w11520_
	);
	LUT4 #(
		.INIT('hd0e0)
	) name10171 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1673_,
		_w6439_,
		_w11520_,
		_w11521_
	);
	LUT2 #(
		.INIT('h6)
	) name10172 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9782_,
		_w11522_
	);
	LUT4 #(
		.INIT('h0800)
	) name10173 (
		\P2_EBX_reg[26]/NET0131 ,
		_w1566_,
		_w1602_,
		_w1611_,
		_w11523_
	);
	LUT3 #(
		.INIT('h02)
	) name10174 (
		_w1673_,
		_w11523_,
		_w11522_,
		_w11524_
	);
	LUT4 #(
		.INIT('h5501)
	) name10175 (
		_w11517_,
		_w11519_,
		_w11521_,
		_w11524_,
		_w11525_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10176 (
		\P2_PhyAddrPointer_reg[26]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11526_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name10177 (
		_w1678_,
		_w11525_,
		_w11516_,
		_w11526_,
		_w11527_
	);
	LUT4 #(
		.INIT('heda5)
	) name10178 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5738_,
		_w5745_,
		_w9793_,
		_w11528_
	);
	LUT2 #(
		.INIT('h2)
	) name10179 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w11529_
	);
	LUT2 #(
		.INIT('h2)
	) name10180 (
		_w1679_,
		_w11529_,
		_w11530_
	);
	LUT4 #(
		.INIT('heb00)
	) name10181 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6877_,
		_w11528_,
		_w11530_,
		_w11531_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10182 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9761_,
		_w9762_,
		_w11532_
	);
	LUT4 #(
		.INIT('h9030)
	) name10183 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w1673_,
		_w9782_,
		_w11533_
	);
	LUT2 #(
		.INIT('h2)
	) name10184 (
		_w6439_,
		_w11533_,
		_w11534_
	);
	LUT4 #(
		.INIT('hde00)
	) name10185 (
		\P2_EBX_reg[27]/NET0131 ,
		_w1673_,
		_w11532_,
		_w11534_,
		_w11535_
	);
	LUT2 #(
		.INIT('h2)
	) name10186 (
		\P2_rEIP_reg[27]/NET0131 ,
		_w9788_,
		_w11536_
	);
	LUT4 #(
		.INIT('h3332)
	) name10187 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[27]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11537_
	);
	LUT3 #(
		.INIT('h02)
	) name10188 (
		_w1566_,
		_w1602_,
		_w11537_,
		_w11538_
	);
	LUT3 #(
		.INIT('hb0)
	) name10189 (
		_w1611_,
		_w11533_,
		_w11538_,
		_w11539_
	);
	LUT2 #(
		.INIT('h1)
	) name10190 (
		_w11536_,
		_w11539_,
		_w11540_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10191 (
		\P2_PhyAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11541_
	);
	LUT4 #(
		.INIT('h7500)
	) name10192 (
		_w1678_,
		_w11535_,
		_w11540_,
		_w11541_,
		_w11542_
	);
	LUT2 #(
		.INIT('hb)
	) name10193 (
		_w11531_,
		_w11542_,
		_w11543_
	);
	LUT3 #(
		.INIT('h48)
	) name10194 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w1673_,
		_w9783_,
		_w11544_
	);
	LUT4 #(
		.INIT('h1000)
	) name10195 (
		\P2_EBX_reg[26]/NET0131 ,
		\P2_EBX_reg[27]/NET0131 ,
		_w9761_,
		_w9762_,
		_w11545_
	);
	LUT4 #(
		.INIT('h0a06)
	) name10196 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w11545_,
		_w11546_
	);
	LUT3 #(
		.INIT('ha8)
	) name10197 (
		_w6439_,
		_w11544_,
		_w11546_,
		_w11547_
	);
	LUT2 #(
		.INIT('h8)
	) name10198 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w11260_,
		_w11548_
	);
	LUT4 #(
		.INIT('hc535)
	) name10199 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w1673_,
		_w9783_,
		_w11549_
	);
	LUT4 #(
		.INIT('ha88a)
	) name10200 (
		\P2_EBX_reg[28]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w11550_
	);
	LUT4 #(
		.INIT('h04f7)
	) name10201 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w1592_,
		_w1601_,
		_w11550_,
		_w11551_
	);
	LUT4 #(
		.INIT('h08aa)
	) name10202 (
		_w1566_,
		_w1674_,
		_w11549_,
		_w11551_,
		_w11552_
	);
	LUT2 #(
		.INIT('h1)
	) name10203 (
		_w11548_,
		_w11552_,
		_w11553_
	);
	LUT3 #(
		.INIT('h8a)
	) name10204 (
		_w1678_,
		_w11547_,
		_w11553_,
		_w11554_
	);
	LUT3 #(
		.INIT('h06)
	) name10205 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9796_,
		_w11555_
	);
	LUT2 #(
		.INIT('h2)
	) name10206 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w11556_
	);
	LUT2 #(
		.INIT('h2)
	) name10207 (
		_w1679_,
		_w11556_,
		_w11557_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10208 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6908_,
		_w11555_,
		_w11557_,
		_w11558_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10209 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11559_
	);
	LUT2 #(
		.INIT('h4)
	) name10210 (
		_w11558_,
		_w11559_,
		_w11560_
	);
	LUT2 #(
		.INIT('hb)
	) name10211 (
		_w11554_,
		_w11560_,
		_w11561_
	);
	LUT4 #(
		.INIT('h4000)
	) name10212 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		\P1_PhyAddrPointer_reg[3]/NET0131 ,
		_w11562_
	);
	LUT3 #(
		.INIT('h06)
	) name10213 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11562_,
		_w11563_
	);
	LUT2 #(
		.INIT('h2)
	) name10214 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w11564_
	);
	LUT2 #(
		.INIT('h2)
	) name10215 (
		_w1939_,
		_w11564_,
		_w11565_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10216 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w9375_,
		_w11563_,
		_w11565_,
		_w11566_
	);
	LUT4 #(
		.INIT('h0309)
	) name10217 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w1930_,
		_w10820_,
		_w11567_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10218 (
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w11568_
	);
	LUT2 #(
		.INIT('h2)
	) name10219 (
		_w1930_,
		_w11568_,
		_w11569_
	);
	LUT2 #(
		.INIT('h1)
	) name10220 (
		_w11567_,
		_w11569_,
		_w11570_
	);
	LUT3 #(
		.INIT('h20)
	) name10221 (
		_w1795_,
		_w1852_,
		_w11570_,
		_w11571_
	);
	LUT4 #(
		.INIT('h3332)
	) name10222 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11572_
	);
	LUT4 #(
		.INIT('h0001)
	) name10223 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11568_,
		_w11573_
	);
	LUT2 #(
		.INIT('h1)
	) name10224 (
		_w11572_,
		_w11573_,
		_w11574_
	);
	LUT3 #(
		.INIT('h20)
	) name10225 (
		_w1797_,
		_w1852_,
		_w11574_,
		_w11575_
	);
	LUT4 #(
		.INIT('h000d)
	) name10226 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w10808_,
		_w11571_,
		_w11575_,
		_w11576_
	);
	LUT2 #(
		.INIT('h2)
	) name10227 (
		\P1_rEIP_reg[4]/NET0131 ,
		_w10828_,
		_w11577_
	);
	LUT3 #(
		.INIT('h07)
	) name10228 (
		\P1_PhyAddrPointer_reg[4]/NET0131 ,
		_w2234_,
		_w3406_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name10229 (
		_w11577_,
		_w11578_,
		_w11579_
	);
	LUT3 #(
		.INIT('hd0)
	) name10230 (
		_w1933_,
		_w11576_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('hb)
	) name10231 (
		_w11566_,
		_w11580_,
		_w11581_
	);
	LUT3 #(
		.INIT('h4c)
	) name10232 (
		\P2_PhyAddrPointer_reg[28]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5743_,
		_w11582_
	);
	LUT4 #(
		.INIT('h00f9)
	) name10233 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w9795_,
		_w11582_,
		_w11583_
	);
	LUT2 #(
		.INIT('h2)
	) name10234 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w11584_
	);
	LUT2 #(
		.INIT('h2)
	) name10235 (
		_w1679_,
		_w11584_,
		_w11585_
	);
	LUT4 #(
		.INIT('heb00)
	) name10236 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6919_,
		_w11583_,
		_w11585_,
		_w11586_
	);
	LUT4 #(
		.INIT('h0509)
	) name10237 (
		\P2_EBX_reg[29]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w1673_,
		_w9764_,
		_w11587_
	);
	LUT4 #(
		.INIT('h70b0)
	) name10238 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w1673_,
		_w6439_,
		_w9784_,
		_w11588_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10239 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[29]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11589_
	);
	LUT3 #(
		.INIT('h0d)
	) name10240 (
		_w1592_,
		_w1601_,
		_w11589_,
		_w11590_
	);
	LUT4 #(
		.INIT('h9f00)
	) name10241 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w9784_,
		_w9751_,
		_w11590_,
		_w11591_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name10242 (
		\P2_rEIP_reg[29]/NET0131 ,
		_w1566_,
		_w11260_,
		_w11591_,
		_w11592_
	);
	LUT3 #(
		.INIT('h02)
	) name10243 (
		_w1566_,
		_w1602_,
		_w11591_,
		_w11593_
	);
	LUT4 #(
		.INIT('h000b)
	) name10244 (
		_w11587_,
		_w11588_,
		_w11592_,
		_w11593_,
		_w11594_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10245 (
		\P2_PhyAddrPointer_reg[29]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11595_
	);
	LUT4 #(
		.INIT('hceff)
	) name10246 (
		_w1678_,
		_w11586_,
		_w11594_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h6)
	) name10247 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w11597_
	);
	LUT2 #(
		.INIT('h2)
	) name10248 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w11598_
	);
	LUT2 #(
		.INIT('h2)
	) name10249 (
		_w1679_,
		_w11598_,
		_w11599_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10250 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w11078_,
		_w11597_,
		_w11599_,
		_w11600_
	);
	LUT2 #(
		.INIT('h2)
	) name10251 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w9788_,
		_w11601_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10252 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11602_
	);
	LUT3 #(
		.INIT('h14)
	) name10253 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w11603_
	);
	LUT3 #(
		.INIT('h10)
	) name10254 (
		_w1605_,
		_w1611_,
		_w11603_,
		_w11604_
	);
	LUT2 #(
		.INIT('h1)
	) name10255 (
		_w11602_,
		_w11604_,
		_w11605_
	);
	LUT2 #(
		.INIT('h2)
	) name10256 (
		_w1566_,
		_w11605_,
		_w11606_
	);
	LUT2 #(
		.INIT('h4)
	) name10257 (
		_w1605_,
		_w11603_,
		_w11607_
	);
	LUT3 #(
		.INIT('he0)
	) name10258 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11608_
	);
	LUT3 #(
		.INIT('h12)
	) name10259 (
		\P2_EBX_reg[2]/NET0131 ,
		_w1673_,
		_w11608_,
		_w11609_
	);
	LUT2 #(
		.INIT('h1)
	) name10260 (
		_w11607_,
		_w11609_,
		_w11610_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10261 (
		_w1442_,
		_w1565_,
		_w1568_,
		_w11610_,
		_w11611_
	);
	LUT3 #(
		.INIT('h45)
	) name10262 (
		_w1602_,
		_w11606_,
		_w11611_,
		_w11612_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10263 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11613_
	);
	LUT4 #(
		.INIT('h5700)
	) name10264 (
		_w1678_,
		_w11601_,
		_w11612_,
		_w11613_,
		_w11614_
	);
	LUT2 #(
		.INIT('hb)
	) name10265 (
		_w11600_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h8)
	) name10266 (
		_w6365_,
		_w10801_,
		_w11616_
	);
	LUT3 #(
		.INIT('h06)
	) name10267 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11616_,
		_w11617_
	);
	LUT2 #(
		.INIT('h2)
	) name10268 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w11618_
	);
	LUT2 #(
		.INIT('h2)
	) name10269 (
		_w1939_,
		_w11618_,
		_w11619_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10270 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w9647_,
		_w11617_,
		_w11619_,
		_w11620_
	);
	LUT4 #(
		.INIT('h9030)
	) name10271 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w1930_,
		_w10810_,
		_w11621_
	);
	LUT4 #(
		.INIT('h3332)
	) name10272 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11622_
	);
	LUT3 #(
		.INIT('h0b)
	) name10273 (
		_w1858_,
		_w11621_,
		_w11622_,
		_w11623_
	);
	LUT3 #(
		.INIT('h20)
	) name10274 (
		_w1797_,
		_w1852_,
		_w11623_,
		_w11624_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10275 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w10820_,
		_w11625_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name10276 (
		\P1_EBX_reg[6]/NET0131 ,
		_w1930_,
		_w11621_,
		_w11625_,
		_w11626_
	);
	LUT3 #(
		.INIT('h20)
	) name10277 (
		_w1795_,
		_w1852_,
		_w11626_,
		_w11627_
	);
	LUT4 #(
		.INIT('h000d)
	) name10278 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w10808_,
		_w11624_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h2)
	) name10279 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w10828_,
		_w11629_
	);
	LUT3 #(
		.INIT('h07)
	) name10280 (
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w2234_,
		_w3406_,
		_w11630_
	);
	LUT2 #(
		.INIT('h4)
	) name10281 (
		_w11629_,
		_w11630_,
		_w11631_
	);
	LUT3 #(
		.INIT('hd0)
	) name10282 (
		_w1933_,
		_w11628_,
		_w11631_,
		_w11632_
	);
	LUT2 #(
		.INIT('hb)
	) name10283 (
		_w11620_,
		_w11632_,
		_w11633_
	);
	LUT3 #(
		.INIT('h40)
	) name10284 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w11634_
	);
	LUT3 #(
		.INIT('h06)
	) name10285 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11634_,
		_w11635_
	);
	LUT2 #(
		.INIT('h2)
	) name10286 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w11636_
	);
	LUT2 #(
		.INIT('h2)
	) name10287 (
		_w1679_,
		_w11636_,
		_w11637_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10288 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9552_,
		_w11635_,
		_w11637_,
		_w11638_
	);
	LUT2 #(
		.INIT('h2)
	) name10289 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w9788_,
		_w11639_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10290 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11640_
	);
	LUT4 #(
		.INIT('h1540)
	) name10291 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w11641_
	);
	LUT3 #(
		.INIT('h10)
	) name10292 (
		_w1605_,
		_w1611_,
		_w11641_,
		_w11642_
	);
	LUT2 #(
		.INIT('h1)
	) name10293 (
		_w11640_,
		_w11642_,
		_w11643_
	);
	LUT2 #(
		.INIT('h2)
	) name10294 (
		_w1566_,
		_w11643_,
		_w11644_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10295 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w11645_
	);
	LUT3 #(
		.INIT('h12)
	) name10296 (
		\P2_EBX_reg[3]/NET0131 ,
		_w1673_,
		_w11645_,
		_w11646_
	);
	LUT2 #(
		.INIT('h4)
	) name10297 (
		_w1605_,
		_w11641_,
		_w11647_
	);
	LUT2 #(
		.INIT('h1)
	) name10298 (
		_w11646_,
		_w11647_,
		_w11648_
	);
	LUT4 #(
		.INIT('h3f15)
	) name10299 (
		_w1565_,
		_w1568_,
		_w1623_,
		_w11648_,
		_w11649_
	);
	LUT3 #(
		.INIT('h45)
	) name10300 (
		_w1602_,
		_w11644_,
		_w11649_,
		_w11650_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10301 (
		\P2_PhyAddrPointer_reg[3]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		_w2211_,
		_w9799_,
		_w11651_
	);
	LUT4 #(
		.INIT('h5700)
	) name10302 (
		_w1678_,
		_w11639_,
		_w11650_,
		_w11651_,
		_w11652_
	);
	LUT2 #(
		.INIT('hb)
	) name10303 (
		_w11638_,
		_w11652_,
		_w11653_
	);
	LUT4 #(
		.INIT('heda5)
	) name10304 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5721_,
		_w5745_,
		_w9792_,
		_w11654_
	);
	LUT2 #(
		.INIT('h2)
	) name10305 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w11655_
	);
	LUT2 #(
		.INIT('h2)
	) name10306 (
		_w1679_,
		_w11655_,
		_w11656_
	);
	LUT4 #(
		.INIT('heb00)
	) name10307 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9338_,
		_w11654_,
		_w11656_,
		_w11657_
	);
	LUT2 #(
		.INIT('h2)
	) name10308 (
		\P2_EBX_reg[31]/NET0131 ,
		_w9753_,
		_w11658_
	);
	LUT4 #(
		.INIT('hfd00)
	) name10309 (
		_w1566_,
		_w1602_,
		_w9751_,
		_w11658_,
		_w11659_
	);
	LUT4 #(
		.INIT('h00a8)
	) name10310 (
		\P2_EBX_reg[4]/NET0131 ,
		_w9752_,
		_w9765_,
		_w11659_,
		_w11660_
	);
	LUT3 #(
		.INIT('h02)
	) name10311 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		_w9753_,
		_w11661_
	);
	LUT4 #(
		.INIT('h0200)
	) name10312 (
		_w1565_,
		_w1602_,
		_w1673_,
		_w11661_,
		_w11662_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10313 (
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w11663_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name10314 (
		_w1673_,
		_w9786_,
		_w11662_,
		_w11663_,
		_w11664_
	);
	LUT3 #(
		.INIT('h8a)
	) name10315 (
		_w1678_,
		_w11660_,
		_w11664_,
		_w11665_
	);
	LUT4 #(
		.INIT('h08aa)
	) name10316 (
		\P2_rEIP_reg[4]/NET0131 ,
		_w1678_,
		_w9788_,
		_w9799_,
		_w11666_
	);
	LUT3 #(
		.INIT('h07)
	) name10317 (
		\P2_PhyAddrPointer_reg[4]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11667_
	);
	LUT2 #(
		.INIT('h4)
	) name10318 (
		_w11666_,
		_w11667_,
		_w11668_
	);
	LUT2 #(
		.INIT('h4)
	) name10319 (
		_w11665_,
		_w11668_,
		_w11669_
	);
	LUT2 #(
		.INIT('hb)
	) name10320 (
		_w11657_,
		_w11669_,
		_w11670_
	);
	LUT4 #(
		.INIT('h4000)
	) name10321 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[6]/NET0131 ,
		_w6365_,
		_w11671_
	);
	LUT3 #(
		.INIT('h06)
	) name10322 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11671_,
		_w11672_
	);
	LUT2 #(
		.INIT('h2)
	) name10323 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w11673_
	);
	LUT2 #(
		.INIT('h2)
	) name10324 (
		_w1939_,
		_w11673_,
		_w11674_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10325 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8724_,
		_w11672_,
		_w11674_,
		_w11675_
	);
	LUT2 #(
		.INIT('h2)
	) name10326 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w10808_,
		_w11676_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10327 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w10810_,
		_w11677_
	);
	LUT3 #(
		.INIT('he2)
	) name10328 (
		\P1_EBX_reg[7]/NET0131 ,
		_w10817_,
		_w11677_,
		_w11678_
	);
	LUT2 #(
		.INIT('h8)
	) name10329 (
		_w1797_,
		_w11678_,
		_w11679_
	);
	LUT4 #(
		.INIT('h0309)
	) name10330 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		_w1930_,
		_w10821_,
		_w11680_
	);
	LUT2 #(
		.INIT('h2)
	) name10331 (
		_w1930_,
		_w11677_,
		_w11681_
	);
	LUT3 #(
		.INIT('h02)
	) name10332 (
		_w1795_,
		_w11681_,
		_w11680_,
		_w11682_
	);
	LUT3 #(
		.INIT('h54)
	) name10333 (
		_w1852_,
		_w11679_,
		_w11682_,
		_w11683_
	);
	LUT2 #(
		.INIT('h2)
	) name10334 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w10828_,
		_w11684_
	);
	LUT3 #(
		.INIT('h07)
	) name10335 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w2234_,
		_w3406_,
		_w11685_
	);
	LUT2 #(
		.INIT('h4)
	) name10336 (
		_w11684_,
		_w11685_,
		_w11686_
	);
	LUT4 #(
		.INIT('h5700)
	) name10337 (
		_w1933_,
		_w11676_,
		_w11683_,
		_w11686_,
		_w11687_
	);
	LUT2 #(
		.INIT('hb)
	) name10338 (
		_w11675_,
		_w11687_,
		_w11688_
	);
	LUT2 #(
		.INIT('h8)
	) name10339 (
		\P1_PhyAddrPointer_reg[7]/NET0131 ,
		_w11671_,
		_w11689_
	);
	LUT3 #(
		.INIT('h06)
	) name10340 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w11689_,
		_w11690_
	);
	LUT2 #(
		.INIT('h2)
	) name10341 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w11691_
	);
	LUT2 #(
		.INIT('h2)
	) name10342 (
		_w1939_,
		_w11691_,
		_w11692_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10343 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8182_,
		_w11690_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h2)
	) name10344 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w10808_,
		_w11694_
	);
	LUT4 #(
		.INIT('h3aca)
	) name10345 (
		\P1_EBX_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w10817_,
		_w10811_,
		_w11695_
	);
	LUT2 #(
		.INIT('h8)
	) name10346 (
		_w1797_,
		_w11695_,
		_w11696_
	);
	LUT3 #(
		.INIT('h8a)
	) name10347 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		_w10821_,
		_w11697_
	);
	LUT3 #(
		.INIT('h21)
	) name10348 (
		\P1_EBX_reg[8]/NET0131 ,
		_w1930_,
		_w11697_,
		_w11698_
	);
	LUT3 #(
		.INIT('h84)
	) name10349 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w1930_,
		_w10811_,
		_w11699_
	);
	LUT3 #(
		.INIT('h02)
	) name10350 (
		_w1795_,
		_w11699_,
		_w11698_,
		_w11700_
	);
	LUT3 #(
		.INIT('h54)
	) name10351 (
		_w1852_,
		_w11696_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h2)
	) name10352 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w10828_,
		_w11702_
	);
	LUT3 #(
		.INIT('h07)
	) name10353 (
		\P1_PhyAddrPointer_reg[8]/NET0131 ,
		_w2234_,
		_w3406_,
		_w11703_
	);
	LUT2 #(
		.INIT('h4)
	) name10354 (
		_w11702_,
		_w11703_,
		_w11704_
	);
	LUT4 #(
		.INIT('h5700)
	) name10355 (
		_w1933_,
		_w11694_,
		_w11701_,
		_w11704_,
		_w11705_
	);
	LUT2 #(
		.INIT('hb)
	) name10356 (
		_w11693_,
		_w11705_,
		_w11706_
	);
	LUT2 #(
		.INIT('h8)
	) name10357 (
		_w5723_,
		_w9792_,
		_w11707_
	);
	LUT3 #(
		.INIT('h06)
	) name10358 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w11707_,
		_w11708_
	);
	LUT2 #(
		.INIT('h2)
	) name10359 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w11709_
	);
	LUT2 #(
		.INIT('h2)
	) name10360 (
		_w1679_,
		_w11709_,
		_w11710_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10361 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9576_,
		_w11708_,
		_w11710_,
		_w11711_
	);
	LUT3 #(
		.INIT('h6c)
	) name10362 (
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		_w9768_,
		_w11712_
	);
	LUT3 #(
		.INIT('h20)
	) name10363 (
		_w1673_,
		_w9786_,
		_w11712_,
		_w11713_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10364 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		_w9753_,
		_w11714_
	);
	LUT4 #(
		.INIT('h08aa)
	) name10365 (
		\P2_EBX_reg[6]/NET0131 ,
		_w1566_,
		_w1602_,
		_w11714_,
		_w11715_
	);
	LUT3 #(
		.INIT('he0)
	) name10366 (
		_w9752_,
		_w9765_,
		_w11715_,
		_w11716_
	);
	LUT2 #(
		.INIT('h4)
	) name10367 (
		\P2_EBX_reg[6]/NET0131 ,
		_w11714_,
		_w11717_
	);
	LUT4 #(
		.INIT('h0200)
	) name10368 (
		_w1565_,
		_w1602_,
		_w1673_,
		_w11717_,
		_w11718_
	);
	LUT3 #(
		.INIT('h0d)
	) name10369 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w9788_,
		_w11718_,
		_w11719_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10370 (
		_w1678_,
		_w11716_,
		_w11713_,
		_w11719_,
		_w11720_
	);
	LUT2 #(
		.INIT('h2)
	) name10371 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w9799_,
		_w11721_
	);
	LUT3 #(
		.INIT('h07)
	) name10372 (
		\P2_PhyAddrPointer_reg[6]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11722_
	);
	LUT2 #(
		.INIT('h4)
	) name10373 (
		_w11721_,
		_w11722_,
		_w11723_
	);
	LUT2 #(
		.INIT('h4)
	) name10374 (
		_w11720_,
		_w11723_,
		_w11724_
	);
	LUT2 #(
		.INIT('hb)
	) name10375 (
		_w11711_,
		_w11724_,
		_w11725_
	);
	LUT4 #(
		.INIT('hd7c3)
	) name10376 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5745_,
		_w7936_,
		_w11726_
	);
	LUT2 #(
		.INIT('h2)
	) name10377 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w11727_
	);
	LUT2 #(
		.INIT('h2)
	) name10378 (
		_w1679_,
		_w11727_,
		_w11728_
	);
	LUT4 #(
		.INIT('heb00)
	) name10379 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8645_,
		_w11726_,
		_w11728_,
		_w11729_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10380 (
		\P2_rEIP_reg[5]/NET0131 ,
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w9768_,
		_w11730_
	);
	LUT3 #(
		.INIT('he2)
	) name10381 (
		\P2_EBX_reg[7]/NET0131 ,
		_w9751_,
		_w11730_,
		_w11731_
	);
	LUT3 #(
		.INIT('h20)
	) name10382 (
		_w1566_,
		_w1602_,
		_w11731_,
		_w11732_
	);
	LUT2 #(
		.INIT('h2)
	) name10383 (
		_w1673_,
		_w11730_,
		_w11733_
	);
	LUT4 #(
		.INIT('h0309)
	) name10384 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		_w1673_,
		_w9754_,
		_w11734_
	);
	LUT2 #(
		.INIT('h1)
	) name10385 (
		_w11733_,
		_w11734_,
		_w11735_
	);
	LUT3 #(
		.INIT('h20)
	) name10386 (
		_w1565_,
		_w1602_,
		_w11735_,
		_w11736_
	);
	LUT4 #(
		.INIT('h000d)
	) name10387 (
		\P2_rEIP_reg[7]/NET0131 ,
		_w9788_,
		_w11732_,
		_w11736_,
		_w11737_
	);
	LUT2 #(
		.INIT('h2)
	) name10388 (
		\P2_rEIP_reg[7]/NET0131 ,
		_w9799_,
		_w11738_
	);
	LUT3 #(
		.INIT('h07)
	) name10389 (
		\P2_PhyAddrPointer_reg[7]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11739_
	);
	LUT2 #(
		.INIT('h4)
	) name10390 (
		_w11738_,
		_w11739_,
		_w11740_
	);
	LUT3 #(
		.INIT('hd0)
	) name10391 (
		_w1678_,
		_w11737_,
		_w11740_,
		_w11741_
	);
	LUT2 #(
		.INIT('hb)
	) name10392 (
		_w11729_,
		_w11741_,
		_w11742_
	);
	LUT3 #(
		.INIT('h06)
	) name10393 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w10802_,
		_w11743_
	);
	LUT2 #(
		.INIT('h2)
	) name10394 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w11744_
	);
	LUT2 #(
		.INIT('h2)
	) name10395 (
		_w1939_,
		_w11744_,
		_w11745_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10396 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8739_,
		_w11743_,
		_w11745_,
		_w11746_
	);
	LUT2 #(
		.INIT('h2)
	) name10397 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w10808_,
		_w11747_
	);
	LUT4 #(
		.INIT('h9030)
	) name10398 (
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10817_,
		_w10811_,
		_w11748_
	);
	LUT4 #(
		.INIT('h3332)
	) name10399 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w1858_,
		_w1861_,
		_w11749_
	);
	LUT3 #(
		.INIT('h02)
	) name10400 (
		_w1797_,
		_w11749_,
		_w11748_,
		_w11750_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10401 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		_w10821_,
		_w11751_
	);
	LUT3 #(
		.INIT('h21)
	) name10402 (
		\P1_EBX_reg[9]/NET0131 ,
		_w1930_,
		_w11751_,
		_w11752_
	);
	LUT4 #(
		.INIT('h9030)
	) name10403 (
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w1930_,
		_w10811_,
		_w11753_
	);
	LUT3 #(
		.INIT('h02)
	) name10404 (
		_w1795_,
		_w11753_,
		_w11752_,
		_w11754_
	);
	LUT3 #(
		.INIT('h54)
	) name10405 (
		_w1852_,
		_w11750_,
		_w11754_,
		_w11755_
	);
	LUT2 #(
		.INIT('h2)
	) name10406 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w10828_,
		_w11756_
	);
	LUT3 #(
		.INIT('h07)
	) name10407 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w2234_,
		_w3406_,
		_w11757_
	);
	LUT2 #(
		.INIT('h4)
	) name10408 (
		_w11756_,
		_w11757_,
		_w11758_
	);
	LUT4 #(
		.INIT('h5700)
	) name10409 (
		_w1933_,
		_w11747_,
		_w11755_,
		_w11758_,
		_w11759_
	);
	LUT2 #(
		.INIT('hb)
	) name10410 (
		_w11746_,
		_w11759_,
		_w11760_
	);
	LUT4 #(
		.INIT('heda5)
	) name10411 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5724_,
		_w5745_,
		_w9792_,
		_w11761_
	);
	LUT2 #(
		.INIT('h2)
	) name10412 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w11762_
	);
	LUT2 #(
		.INIT('h2)
	) name10413 (
		_w1679_,
		_w11762_,
		_w11763_
	);
	LUT4 #(
		.INIT('heb00)
	) name10414 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w7938_,
		_w11761_,
		_w11763_,
		_w11764_
	);
	LUT3 #(
		.INIT('h8a)
	) name10415 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		_w9754_,
		_w11765_
	);
	LUT4 #(
		.INIT('h1444)
	) name10416 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w9768_,
		_w9769_,
		_w11766_
	);
	LUT2 #(
		.INIT('h4)
	) name10417 (
		_w1605_,
		_w11766_,
		_w11767_
	);
	LUT4 #(
		.INIT('h00ed)
	) name10418 (
		\P2_EBX_reg[8]/NET0131 ,
		_w1673_,
		_w11765_,
		_w11767_,
		_w11768_
	);
	LUT4 #(
		.INIT('hccc8)
	) name10419 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		_w1605_,
		_w1611_,
		_w11769_
	);
	LUT3 #(
		.INIT('h07)
	) name10420 (
		_w1612_,
		_w11766_,
		_w11769_,
		_w11770_
	);
	LUT4 #(
		.INIT('hf531)
	) name10421 (
		_w1565_,
		_w1566_,
		_w11768_,
		_w11770_,
		_w11771_
	);
	LUT4 #(
		.INIT('h5750)
	) name10422 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w1569_,
		_w1602_,
		_w11771_,
		_w11772_
	);
	LUT2 #(
		.INIT('h2)
	) name10423 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9799_,
		_w11773_
	);
	LUT3 #(
		.INIT('h07)
	) name10424 (
		\P2_PhyAddrPointer_reg[8]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11774_
	);
	LUT2 #(
		.INIT('h4)
	) name10425 (
		_w11773_,
		_w11774_,
		_w11775_
	);
	LUT3 #(
		.INIT('hd0)
	) name10426 (
		_w1678_,
		_w11772_,
		_w11775_,
		_w11776_
	);
	LUT2 #(
		.INIT('hb)
	) name10427 (
		_w11764_,
		_w11776_,
		_w11777_
	);
	LUT4 #(
		.INIT('heda5)
	) name10428 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5725_,
		_w5745_,
		_w9792_,
		_w11778_
	);
	LUT2 #(
		.INIT('h2)
	) name10429 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w11779_
	);
	LUT2 #(
		.INIT('h2)
	) name10430 (
		_w1679_,
		_w11779_,
		_w11780_
	);
	LUT4 #(
		.INIT('heb00)
	) name10431 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w8655_,
		_w11778_,
		_w11780_,
		_w11781_
	);
	LUT2 #(
		.INIT('h2)
	) name10432 (
		\P2_rEIP_reg[9]/NET0131 ,
		_w9788_,
		_w11782_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10433 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w9768_,
		_w9769_,
		_w11783_
	);
	LUT3 #(
		.INIT('he2)
	) name10434 (
		\P2_EBX_reg[9]/NET0131 ,
		_w9751_,
		_w11783_,
		_w11784_
	);
	LUT2 #(
		.INIT('h8)
	) name10435 (
		_w1566_,
		_w11784_,
		_w11785_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10436 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		_w9754_,
		_w11786_
	);
	LUT3 #(
		.INIT('h21)
	) name10437 (
		\P2_EBX_reg[9]/NET0131 ,
		_w1673_,
		_w11786_,
		_w11787_
	);
	LUT2 #(
		.INIT('h2)
	) name10438 (
		_w1673_,
		_w11783_,
		_w11788_
	);
	LUT3 #(
		.INIT('h02)
	) name10439 (
		_w1565_,
		_w11788_,
		_w11787_,
		_w11789_
	);
	LUT3 #(
		.INIT('h54)
	) name10440 (
		_w1602_,
		_w11785_,
		_w11789_,
		_w11790_
	);
	LUT2 #(
		.INIT('h2)
	) name10441 (
		\P2_rEIP_reg[9]/NET0131 ,
		_w9799_,
		_w11791_
	);
	LUT3 #(
		.INIT('h07)
	) name10442 (
		\P2_PhyAddrPointer_reg[9]/NET0131 ,
		_w2211_,
		_w2286_,
		_w11792_
	);
	LUT2 #(
		.INIT('h4)
	) name10443 (
		_w11791_,
		_w11792_,
		_w11793_
	);
	LUT4 #(
		.INIT('h5700)
	) name10444 (
		_w1678_,
		_w11782_,
		_w11790_,
		_w11793_,
		_w11794_
	);
	LUT2 #(
		.INIT('hb)
	) name10445 (
		_w11781_,
		_w11794_,
		_w11795_
	);
	LUT4 #(
		.INIT('h4000)
	) name10446 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w5758_,
		_w11796_
	);
	LUT3 #(
		.INIT('h80)
	) name10447 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w5760_,
		_w11796_,
		_w11797_
	);
	LUT4 #(
		.INIT('h0514)
	) name10448 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8672_,
		_w11797_,
		_w11798_
	);
	LUT2 #(
		.INIT('h2)
	) name10449 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w11799_
	);
	LUT2 #(
		.INIT('h2)
	) name10450 (
		_w2194_,
		_w11799_,
		_w11800_
	);
	LUT4 #(
		.INIT('haa02)
	) name10451 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11801_
	);
	LUT2 #(
		.INIT('h4)
	) name10452 (
		_w2111_,
		_w2187_,
		_w11802_
	);
	LUT4 #(
		.INIT('h8000)
	) name10453 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w11803_
	);
	LUT4 #(
		.INIT('h8000)
	) name10454 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w11803_,
		_w11804_
	);
	LUT3 #(
		.INIT('h80)
	) name10455 (
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w11804_,
		_w11805_
	);
	LUT4 #(
		.INIT('h8000)
	) name10456 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w11804_,
		_w11806_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10457 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w11804_,
		_w11807_
	);
	LUT2 #(
		.INIT('h2)
	) name10458 (
		_w11802_,
		_w11807_,
		_w11808_
	);
	LUT3 #(
		.INIT('h45)
	) name10459 (
		\P3_EBX_reg[10]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11809_
	);
	LUT4 #(
		.INIT('h0008)
	) name10460 (
		_w2060_,
		_w2047_,
		_w11809_,
		_w11808_,
		_w11810_
	);
	LUT4 #(
		.INIT('h0001)
	) name10461 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w11811_
	);
	LUT4 #(
		.INIT('h0100)
	) name10462 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w11811_,
		_w11812_
	);
	LUT4 #(
		.INIT('h0100)
	) name10463 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w11812_,
		_w11813_
	);
	LUT4 #(
		.INIT('h0509)
	) name10464 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w11813_,
		_w11814_
	);
	LUT2 #(
		.INIT('h2)
	) name10465 (
		_w2187_,
		_w11807_,
		_w11815_
	);
	LUT4 #(
		.INIT('h0004)
	) name10466 (
		_w2060_,
		_w2047_,
		_w11815_,
		_w11814_,
		_w11816_
	);
	LUT4 #(
		.INIT('h2223)
	) name10467 (
		_w2105_,
		_w11801_,
		_w11810_,
		_w11816_,
		_w11817_
	);
	LUT4 #(
		.INIT('hfe25)
	) name10468 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w11818_
	);
	LUT2 #(
		.INIT('h2)
	) name10469 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w11818_,
		_w11819_
	);
	LUT3 #(
		.INIT('h07)
	) name10470 (
		\P3_PhyAddrPointer_reg[10]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11820_
	);
	LUT2 #(
		.INIT('h4)
	) name10471 (
		_w11819_,
		_w11820_,
		_w11821_
	);
	LUT3 #(
		.INIT('hd0)
	) name10472 (
		_w1945_,
		_w11817_,
		_w11821_,
		_w11822_
	);
	LUT3 #(
		.INIT('h4f)
	) name10473 (
		_w11798_,
		_w11800_,
		_w11822_,
		_w11823_
	);
	LUT2 #(
		.INIT('h4)
	) name10474 (
		_w8672_,
		_w11797_,
		_w11824_
	);
	LUT4 #(
		.INIT('h0514)
	) name10475 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7429_,
		_w11824_,
		_w11825_
	);
	LUT2 #(
		.INIT('h2)
	) name10476 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w11826_
	);
	LUT2 #(
		.INIT('h2)
	) name10477 (
		_w2194_,
		_w11826_,
		_w11827_
	);
	LUT3 #(
		.INIT('h8c)
	) name10478 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11813_,
		_w11828_
	);
	LUT3 #(
		.INIT('h21)
	) name10479 (
		\P3_EBX_reg[11]/NET0131 ,
		_w2187_,
		_w11828_,
		_w11829_
	);
	LUT3 #(
		.INIT('h84)
	) name10480 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w2187_,
		_w11806_,
		_w11830_
	);
	LUT3 #(
		.INIT('h04)
	) name10481 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w11831_
	);
	LUT4 #(
		.INIT('h0004)
	) name10482 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w11830_,
		_w11832_
	);
	LUT2 #(
		.INIT('h4)
	) name10483 (
		_w11829_,
		_w11832_,
		_w11833_
	);
	LUT4 #(
		.INIT('haa02)
	) name10484 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11834_
	);
	LUT4 #(
		.INIT('h2010)
	) name10485 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11806_,
		_w11835_
	);
	LUT3 #(
		.INIT('h45)
	) name10486 (
		\P3_EBX_reg[11]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11836_
	);
	LUT4 #(
		.INIT('h0008)
	) name10487 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w11836_,
		_w11837_
	);
	LUT3 #(
		.INIT('h45)
	) name10488 (
		_w11834_,
		_w11835_,
		_w11837_,
		_w11838_
	);
	LUT2 #(
		.INIT('h2)
	) name10489 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w11818_,
		_w11839_
	);
	LUT3 #(
		.INIT('h07)
	) name10490 (
		\P3_PhyAddrPointer_reg[11]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11840_
	);
	LUT2 #(
		.INIT('h4)
	) name10491 (
		_w11839_,
		_w11840_,
		_w11841_
	);
	LUT4 #(
		.INIT('h7500)
	) name10492 (
		_w1945_,
		_w11833_,
		_w11838_,
		_w11841_,
		_w11842_
	);
	LUT3 #(
		.INIT('h4f)
	) name10493 (
		_w11825_,
		_w11827_,
		_w11842_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name10494 (
		_w7429_,
		_w11824_,
		_w11844_
	);
	LUT4 #(
		.INIT('h0514)
	) name10495 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7948_,
		_w11844_,
		_w11845_
	);
	LUT2 #(
		.INIT('h2)
	) name10496 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w11846_
	);
	LUT2 #(
		.INIT('h2)
	) name10497 (
		_w2194_,
		_w11846_,
		_w11847_
	);
	LUT4 #(
		.INIT('haa02)
	) name10498 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11848_
	);
	LUT4 #(
		.INIT('h9030)
	) name10499 (
		\P3_rEIP_reg[11]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w2187_,
		_w11806_,
		_w11849_
	);
	LUT3 #(
		.INIT('h45)
	) name10500 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11850_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10501 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11813_,
		_w11851_
	);
	LUT3 #(
		.INIT('h21)
	) name10502 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2187_,
		_w11851_,
		_w11852_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name10503 (
		_w2060_,
		_w2047_,
		_w11850_,
		_w11852_,
		_w11853_
	);
	LUT4 #(
		.INIT('h0080)
	) name10504 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w11850_,
		_w11854_
	);
	LUT4 #(
		.INIT('h5501)
	) name10505 (
		_w2105_,
		_w11849_,
		_w11853_,
		_w11854_,
		_w11855_
	);
	LUT2 #(
		.INIT('h2)
	) name10506 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w11818_,
		_w11856_
	);
	LUT3 #(
		.INIT('h07)
	) name10507 (
		\P3_PhyAddrPointer_reg[12]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11857_
	);
	LUT2 #(
		.INIT('h4)
	) name10508 (
		_w11856_,
		_w11857_,
		_w11858_
	);
	LUT4 #(
		.INIT('h5700)
	) name10509 (
		_w1945_,
		_w11848_,
		_w11855_,
		_w11858_,
		_w11859_
	);
	LUT3 #(
		.INIT('h4f)
	) name10510 (
		_w11845_,
		_w11847_,
		_w11859_,
		_w11860_
	);
	LUT3 #(
		.INIT('h10)
	) name10511 (
		_w7429_,
		_w7948_,
		_w11824_,
		_w11861_
	);
	LUT4 #(
		.INIT('h0514)
	) name10512 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7967_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h2)
	) name10513 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w11863_
	);
	LUT2 #(
		.INIT('h2)
	) name10514 (
		_w2194_,
		_w11863_,
		_w11864_
	);
	LUT4 #(
		.INIT('haa02)
	) name10515 (
		\P3_rEIP_reg[13]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11865_
	);
	LUT3 #(
		.INIT('h45)
	) name10516 (
		\P3_EBX_reg[13]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11866_
	);
	LUT4 #(
		.INIT('h0100)
	) name10517 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		\P3_EBX_reg[12]/NET0131 ,
		_w11813_,
		_w11867_
	);
	LUT4 #(
		.INIT('h0509)
	) name10518 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w11867_,
		_w11868_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name10519 (
		_w2060_,
		_w2047_,
		_w11866_,
		_w11868_,
		_w11869_
	);
	LUT4 #(
		.INIT('h0080)
	) name10520 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w11866_,
		_w11870_
	);
	LUT4 #(
		.INIT('h8000)
	) name10521 (
		\P3_rEIP_reg[11]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w11806_,
		_w11871_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10522 (
		\P3_rEIP_reg[11]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w11806_,
		_w11872_
	);
	LUT2 #(
		.INIT('h2)
	) name10523 (
		_w2187_,
		_w11872_,
		_w11873_
	);
	LUT4 #(
		.INIT('h0045)
	) name10524 (
		_w2105_,
		_w11870_,
		_w11873_,
		_w11869_,
		_w11874_
	);
	LUT2 #(
		.INIT('h2)
	) name10525 (
		\P3_rEIP_reg[13]/NET0131 ,
		_w11818_,
		_w11875_
	);
	LUT3 #(
		.INIT('h07)
	) name10526 (
		\P3_PhyAddrPointer_reg[13]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11876_
	);
	LUT2 #(
		.INIT('h4)
	) name10527 (
		_w11875_,
		_w11876_,
		_w11877_
	);
	LUT4 #(
		.INIT('h5700)
	) name10528 (
		_w1945_,
		_w11865_,
		_w11874_,
		_w11877_,
		_w11878_
	);
	LUT3 #(
		.INIT('h4f)
	) name10529 (
		_w11862_,
		_w11864_,
		_w11878_,
		_w11879_
	);
	LUT4 #(
		.INIT('h0100)
	) name10530 (
		_w7429_,
		_w7948_,
		_w7967_,
		_w11824_,
		_w11880_
	);
	LUT4 #(
		.INIT('h0514)
	) name10531 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7984_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h2)
	) name10532 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w11882_
	);
	LUT2 #(
		.INIT('h2)
	) name10533 (
		_w2194_,
		_w11882_,
		_w11883_
	);
	LUT4 #(
		.INIT('haa02)
	) name10534 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11884_
	);
	LUT3 #(
		.INIT('h84)
	) name10535 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w11802_,
		_w11871_,
		_w11885_
	);
	LUT3 #(
		.INIT('h45)
	) name10536 (
		\P3_EBX_reg[14]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11886_
	);
	LUT4 #(
		.INIT('h0008)
	) name10537 (
		_w2060_,
		_w2047_,
		_w11886_,
		_w11885_,
		_w11887_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name10538 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11867_,
		_w11888_
	);
	LUT2 #(
		.INIT('h1)
	) name10539 (
		_w2187_,
		_w11888_,
		_w11889_
	);
	LUT3 #(
		.INIT('h84)
	) name10540 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w2187_,
		_w11871_,
		_w11890_
	);
	LUT3 #(
		.INIT('h04)
	) name10541 (
		_w2060_,
		_w2047_,
		_w11890_,
		_w11891_
	);
	LUT4 #(
		.INIT('h4544)
	) name10542 (
		_w2105_,
		_w11887_,
		_w11889_,
		_w11891_,
		_w11892_
	);
	LUT2 #(
		.INIT('h2)
	) name10543 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w11818_,
		_w11893_
	);
	LUT3 #(
		.INIT('h07)
	) name10544 (
		\P3_PhyAddrPointer_reg[14]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11894_
	);
	LUT2 #(
		.INIT('h4)
	) name10545 (
		_w11893_,
		_w11894_,
		_w11895_
	);
	LUT4 #(
		.INIT('h5700)
	) name10546 (
		_w1945_,
		_w11884_,
		_w11892_,
		_w11895_,
		_w11896_
	);
	LUT3 #(
		.INIT('h4f)
	) name10547 (
		_w11881_,
		_w11883_,
		_w11896_,
		_w11897_
	);
	LUT2 #(
		.INIT('h4)
	) name10548 (
		_w7984_,
		_w11880_,
		_w11898_
	);
	LUT4 #(
		.INIT('h0514)
	) name10549 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7445_,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('h2)
	) name10550 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w11900_
	);
	LUT2 #(
		.INIT('h2)
	) name10551 (
		_w2194_,
		_w11900_,
		_w11901_
	);
	LUT4 #(
		.INIT('haa02)
	) name10552 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11902_
	);
	LUT3 #(
		.INIT('h45)
	) name10553 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11903_
	);
	LUT3 #(
		.INIT('h08)
	) name10554 (
		_w2060_,
		_w2047_,
		_w11903_,
		_w11904_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10555 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11867_,
		_w11905_
	);
	LUT3 #(
		.INIT('h21)
	) name10556 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2187_,
		_w11905_,
		_w11906_
	);
	LUT3 #(
		.INIT('h31)
	) name10557 (
		_w2106_,
		_w11904_,
		_w11906_,
		_w11907_
	);
	LUT3 #(
		.INIT('h6c)
	) name10558 (
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w11871_,
		_w11908_
	);
	LUT4 #(
		.INIT('h0080)
	) name10559 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w11903_,
		_w11909_
	);
	LUT4 #(
		.INIT('h5551)
	) name10560 (
		_w2105_,
		_w2187_,
		_w11908_,
		_w11909_,
		_w11910_
	);
	LUT4 #(
		.INIT('h8a88)
	) name10561 (
		_w1945_,
		_w11902_,
		_w11907_,
		_w11910_,
		_w11911_
	);
	LUT2 #(
		.INIT('h2)
	) name10562 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w11818_,
		_w11912_
	);
	LUT3 #(
		.INIT('h07)
	) name10563 (
		\P3_PhyAddrPointer_reg[15]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11913_
	);
	LUT2 #(
		.INIT('h4)
	) name10564 (
		_w11912_,
		_w11913_,
		_w11914_
	);
	LUT2 #(
		.INIT('h4)
	) name10565 (
		_w11911_,
		_w11914_,
		_w11915_
	);
	LUT3 #(
		.INIT('h4f)
	) name10566 (
		_w11899_,
		_w11901_,
		_w11915_,
		_w11916_
	);
	LUT4 #(
		.INIT('h0e00)
	) name10567 (
		_w7442_,
		_w7444_,
		_w7984_,
		_w11880_,
		_w11917_
	);
	LUT4 #(
		.INIT('h0514)
	) name10568 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8001_,
		_w11917_,
		_w11918_
	);
	LUT2 #(
		.INIT('h2)
	) name10569 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w11919_
	);
	LUT2 #(
		.INIT('h2)
	) name10570 (
		_w2194_,
		_w11919_,
		_w11920_
	);
	LUT2 #(
		.INIT('h8)
	) name10571 (
		\P3_EBX_reg[15]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11921_
	);
	LUT4 #(
		.INIT('h2221)
	) name10572 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2187_,
		_w11905_,
		_w11921_,
		_w11922_
	);
	LUT4 #(
		.INIT('h8000)
	) name10573 (
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w11871_,
		_w11923_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10574 (
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w11871_,
		_w11924_
	);
	LUT2 #(
		.INIT('h2)
	) name10575 (
		_w2187_,
		_w11924_,
		_w11925_
	);
	LUT3 #(
		.INIT('h02)
	) name10576 (
		_w11831_,
		_w11922_,
		_w11925_,
		_w11926_
	);
	LUT4 #(
		.INIT('haa02)
	) name10577 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11927_
	);
	LUT2 #(
		.INIT('h2)
	) name10578 (
		_w11802_,
		_w11924_,
		_w11928_
	);
	LUT3 #(
		.INIT('h45)
	) name10579 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11929_
	);
	LUT4 #(
		.INIT('h0008)
	) name10580 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w11929_,
		_w11930_
	);
	LUT3 #(
		.INIT('h45)
	) name10581 (
		_w11927_,
		_w11928_,
		_w11930_,
		_w11931_
	);
	LUT2 #(
		.INIT('h2)
	) name10582 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w11818_,
		_w11932_
	);
	LUT3 #(
		.INIT('h07)
	) name10583 (
		\P3_PhyAddrPointer_reg[16]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11933_
	);
	LUT2 #(
		.INIT('h4)
	) name10584 (
		_w11932_,
		_w11933_,
		_w11934_
	);
	LUT4 #(
		.INIT('h7500)
	) name10585 (
		_w1945_,
		_w11926_,
		_w11931_,
		_w11934_,
		_w11935_
	);
	LUT3 #(
		.INIT('h4f)
	) name10586 (
		_w11918_,
		_w11920_,
		_w11935_,
		_w11936_
	);
	LUT2 #(
		.INIT('h4)
	) name10587 (
		_w8001_,
		_w11917_,
		_w11937_
	);
	LUT3 #(
		.INIT('h15)
	) name10588 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5765_,
		_w7441_,
		_w11938_
	);
	LUT2 #(
		.INIT('h1)
	) name10589 (
		_w8018_,
		_w11938_,
		_w11939_
	);
	LUT4 #(
		.INIT('h0154)
	) name10590 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w11937_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h2)
	) name10591 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w11941_
	);
	LUT2 #(
		.INIT('h2)
	) name10592 (
		_w2194_,
		_w11941_,
		_w11942_
	);
	LUT3 #(
		.INIT('h84)
	) name10593 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2187_,
		_w11923_,
		_w11943_
	);
	LUT4 #(
		.INIT('h3222)
	) name10594 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[17]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w11944_
	);
	LUT3 #(
		.INIT('h01)
	) name10595 (
		_w2111_,
		_w2105_,
		_w11944_,
		_w11945_
	);
	LUT4 #(
		.INIT('h7b00)
	) name10596 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2187_,
		_w11923_,
		_w11945_,
		_w11946_
	);
	LUT4 #(
		.INIT('h335f)
	) name10597 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w2111_,
		_w2105_,
		_w11947_
	);
	LUT3 #(
		.INIT('h8a)
	) name10598 (
		_w2113_,
		_w11946_,
		_w11947_,
		_w11948_
	);
	LUT4 #(
		.INIT('hdf03)
	) name10599 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11949_
	);
	LUT2 #(
		.INIT('h8)
	) name10600 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w11949_,
		_w11950_
	);
	LUT2 #(
		.INIT('h1)
	) name10601 (
		\P3_EBX_reg[15]/NET0131 ,
		\P3_EBX_reg[16]/NET0131 ,
		_w11951_
	);
	LUT4 #(
		.INIT('h1000)
	) name10602 (
		\P3_EBX_reg[13]/NET0131 ,
		\P3_EBX_reg[14]/NET0131 ,
		_w11867_,
		_w11951_,
		_w11952_
	);
	LUT4 #(
		.INIT('h0509)
	) name10603 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w11952_,
		_w11953_
	);
	LUT3 #(
		.INIT('h02)
	) name10604 (
		_w11831_,
		_w11943_,
		_w11953_,
		_w11954_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10605 (
		_w1945_,
		_w11950_,
		_w11948_,
		_w11954_,
		_w11955_
	);
	LUT2 #(
		.INIT('h2)
	) name10606 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w11818_,
		_w11956_
	);
	LUT3 #(
		.INIT('h07)
	) name10607 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11957_
	);
	LUT2 #(
		.INIT('h4)
	) name10608 (
		_w11956_,
		_w11957_,
		_w11958_
	);
	LUT2 #(
		.INIT('h4)
	) name10609 (
		_w11955_,
		_w11958_,
		_w11959_
	);
	LUT3 #(
		.INIT('h4f)
	) name10610 (
		_w11940_,
		_w11942_,
		_w11959_,
		_w11960_
	);
	LUT3 #(
		.INIT('h04)
	) name10611 (
		_w8001_,
		_w11917_,
		_w11939_,
		_w11961_
	);
	LUT4 #(
		.INIT('h0514)
	) name10612 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8020_,
		_w11961_,
		_w11962_
	);
	LUT2 #(
		.INIT('h2)
	) name10613 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w11963_
	);
	LUT2 #(
		.INIT('h2)
	) name10614 (
		_w2194_,
		_w11963_,
		_w11964_
	);
	LUT4 #(
		.INIT('haa02)
	) name10615 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11965_
	);
	LUT3 #(
		.INIT('h45)
	) name10616 (
		\P3_EBX_reg[18]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11966_
	);
	LUT3 #(
		.INIT('h08)
	) name10617 (
		_w2060_,
		_w2047_,
		_w11966_,
		_w11967_
	);
	LUT3 #(
		.INIT('h73)
	) name10618 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11952_,
		_w11968_
	);
	LUT4 #(
		.INIT('hc8c4)
	) name10619 (
		\P3_EBX_reg[18]/NET0131 ,
		_w2106_,
		_w2187_,
		_w11968_,
		_w11969_
	);
	LUT2 #(
		.INIT('h8)
	) name10620 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w11970_
	);
	LUT3 #(
		.INIT('h6c)
	) name10621 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w11923_,
		_w11971_
	);
	LUT4 #(
		.INIT('h0080)
	) name10622 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w11966_,
		_w11972_
	);
	LUT4 #(
		.INIT('h5551)
	) name10623 (
		_w2105_,
		_w2187_,
		_w11971_,
		_w11972_,
		_w11973_
	);
	LUT4 #(
		.INIT('h0155)
	) name10624 (
		_w11965_,
		_w11967_,
		_w11969_,
		_w11973_,
		_w11974_
	);
	LUT2 #(
		.INIT('h2)
	) name10625 (
		\P3_rEIP_reg[18]/NET0131 ,
		_w11818_,
		_w11975_
	);
	LUT3 #(
		.INIT('h07)
	) name10626 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11976_
	);
	LUT2 #(
		.INIT('h4)
	) name10627 (
		_w11975_,
		_w11976_,
		_w11977_
	);
	LUT3 #(
		.INIT('hd0)
	) name10628 (
		_w1945_,
		_w11974_,
		_w11977_,
		_w11978_
	);
	LUT3 #(
		.INIT('h4f)
	) name10629 (
		_w11962_,
		_w11964_,
		_w11978_,
		_w11979_
	);
	LUT3 #(
		.INIT('h32)
	) name10630 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w7467_,
		_w8019_,
		_w11980_
	);
	LUT3 #(
		.INIT('hba)
	) name10631 (
		_w5779_,
		_w8020_,
		_w11961_,
		_w11981_
	);
	LUT2 #(
		.INIT('h2)
	) name10632 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w11982_
	);
	LUT2 #(
		.INIT('h2)
	) name10633 (
		_w2194_,
		_w11982_,
		_w11983_
	);
	LUT4 #(
		.INIT('heb00)
	) name10634 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w11980_,
		_w11981_,
		_w11983_,
		_w11984_
	);
	LUT4 #(
		.INIT('haa02)
	) name10635 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w11985_
	);
	LUT3 #(
		.INIT('h45)
	) name10636 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11986_
	);
	LUT3 #(
		.INIT('h08)
	) name10637 (
		_w2060_,
		_w2047_,
		_w11986_,
		_w11987_
	);
	LUT2 #(
		.INIT('h1)
	) name10638 (
		\P3_EBX_reg[17]/NET0131 ,
		\P3_EBX_reg[18]/NET0131 ,
		_w11988_
	);
	LUT3 #(
		.INIT('h2a)
	) name10639 (
		\P3_EBX_reg[31]/NET0131 ,
		_w11952_,
		_w11988_,
		_w11989_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name10640 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2106_,
		_w2187_,
		_w11989_,
		_w11990_
	);
	LUT3 #(
		.INIT('h6a)
	) name10641 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11923_,
		_w11970_,
		_w11991_
	);
	LUT4 #(
		.INIT('h0080)
	) name10642 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w11986_,
		_w11992_
	);
	LUT4 #(
		.INIT('h5551)
	) name10643 (
		_w2105_,
		_w2187_,
		_w11991_,
		_w11992_,
		_w11993_
	);
	LUT4 #(
		.INIT('h0155)
	) name10644 (
		_w11985_,
		_w11987_,
		_w11990_,
		_w11993_,
		_w11994_
	);
	LUT2 #(
		.INIT('h2)
	) name10645 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11818_,
		_w11995_
	);
	LUT3 #(
		.INIT('h07)
	) name10646 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2225_,
		_w3054_,
		_w11996_
	);
	LUT2 #(
		.INIT('h4)
	) name10647 (
		_w11995_,
		_w11996_,
		_w11997_
	);
	LUT3 #(
		.INIT('hd0)
	) name10648 (
		_w1945_,
		_w11994_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('hb)
	) name10649 (
		_w11984_,
		_w11998_,
		_w11999_
	);
	LUT4 #(
		.INIT('h5014)
	) name10650 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5779_,
		_w12000_
	);
	LUT2 #(
		.INIT('h2)
	) name10651 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w12001_
	);
	LUT2 #(
		.INIT('h2)
	) name10652 (
		_w2194_,
		_w12001_,
		_w12002_
	);
	LUT4 #(
		.INIT('haa02)
	) name10653 (
		\P3_rEIP_reg[1]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12003_
	);
	LUT2 #(
		.INIT('h6)
	) name10654 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		_w12004_
	);
	LUT3 #(
		.INIT('h90)
	) name10655 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12005_
	);
	LUT2 #(
		.INIT('h1)
	) name10656 (
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12006_
	);
	LUT2 #(
		.INIT('h1)
	) name10657 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w12007_
	);
	LUT4 #(
		.INIT('h0111)
	) name10658 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12008_
	);
	LUT4 #(
		.INIT('h00fe)
	) name10659 (
		_w2187_,
		_w12006_,
		_w12005_,
		_w12008_,
		_w12009_
	);
	LUT3 #(
		.INIT('h04)
	) name10660 (
		_w2060_,
		_w2047_,
		_w12009_,
		_w12010_
	);
	LUT2 #(
		.INIT('h8)
	) name10661 (
		_w2044_,
		_w2100_,
		_w12011_
	);
	LUT3 #(
		.INIT('h8a)
	) name10662 (
		\P3_EBX_reg[1]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12012_
	);
	LUT3 #(
		.INIT('h10)
	) name10663 (
		_w2111_,
		_w2116_,
		_w12007_,
		_w12013_
	);
	LUT2 #(
		.INIT('h1)
	) name10664 (
		_w12012_,
		_w12013_,
		_w12014_
	);
	LUT3 #(
		.INIT('h08)
	) name10665 (
		_w2060_,
		_w2047_,
		_w12014_,
		_w12015_
	);
	LUT4 #(
		.INIT('h5554)
	) name10666 (
		_w2105_,
		_w12011_,
		_w12015_,
		_w12010_,
		_w12016_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10667 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12017_
	);
	LUT4 #(
		.INIT('h5700)
	) name10668 (
		_w1945_,
		_w12003_,
		_w12016_,
		_w12017_,
		_w12018_
	);
	LUT3 #(
		.INIT('h4f)
	) name10669 (
		_w12000_,
		_w12002_,
		_w12018_,
		_w12019_
	);
	LUT4 #(
		.INIT('h8111)
	) name10670 (
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5767_,
		_w12020_
	);
	LUT4 #(
		.INIT('h0400)
	) name10671 (
		_w8001_,
		_w11917_,
		_w11939_,
		_w12020_,
		_w12021_
	);
	LUT4 #(
		.INIT('h0514)
	) name10672 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7469_,
		_w12021_,
		_w12022_
	);
	LUT2 #(
		.INIT('h2)
	) name10673 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w12023_
	);
	LUT2 #(
		.INIT('h2)
	) name10674 (
		_w2194_,
		_w12023_,
		_w12024_
	);
	LUT3 #(
		.INIT('h80)
	) name10675 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w12025_
	);
	LUT4 #(
		.INIT('h8000)
	) name10676 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w12026_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10677 (
		\P3_rEIP_reg[19]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w11923_,
		_w11970_,
		_w12027_
	);
	LUT4 #(
		.INIT('h3222)
	) name10678 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12028_
	);
	LUT3 #(
		.INIT('h01)
	) name10679 (
		_w2111_,
		_w2105_,
		_w12028_,
		_w12029_
	);
	LUT4 #(
		.INIT('h335f)
	) name10680 (
		\P3_EBX_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w2111_,
		_w2105_,
		_w12030_
	);
	LUT4 #(
		.INIT('h2f00)
	) name10681 (
		_w2187_,
		_w12027_,
		_w12029_,
		_w12030_,
		_w12031_
	);
	LUT2 #(
		.INIT('h2)
	) name10682 (
		_w2113_,
		_w12031_,
		_w12032_
	);
	LUT2 #(
		.INIT('h8)
	) name10683 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w11949_,
		_w12033_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10684 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w11952_,
		_w11988_,
		_w12034_
	);
	LUT3 #(
		.INIT('h21)
	) name10685 (
		\P3_EBX_reg[20]/NET0131 ,
		_w2187_,
		_w12034_,
		_w12035_
	);
	LUT3 #(
		.INIT('hc4)
	) name10686 (
		_w2187_,
		_w11831_,
		_w12027_,
		_w12036_
	);
	LUT3 #(
		.INIT('h45)
	) name10687 (
		_w12033_,
		_w12035_,
		_w12036_,
		_w12037_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10688 (
		\P3_PhyAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12038_
	);
	LUT4 #(
		.INIT('h7500)
	) name10689 (
		_w1945_,
		_w12032_,
		_w12037_,
		_w12038_,
		_w12039_
	);
	LUT3 #(
		.INIT('h4f)
	) name10690 (
		_w12022_,
		_w12024_,
		_w12039_,
		_w12040_
	);
	LUT3 #(
		.INIT('hba)
	) name10691 (
		_w5779_,
		_w7469_,
		_w12021_,
		_w12041_
	);
	LUT2 #(
		.INIT('h2)
	) name10692 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w12042_
	);
	LUT2 #(
		.INIT('h2)
	) name10693 (
		_w2194_,
		_w12042_,
		_w12043_
	);
	LUT4 #(
		.INIT('heb00)
	) name10694 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8032_,
		_w12041_,
		_w12043_,
		_w12044_
	);
	LUT2 #(
		.INIT('h1)
	) name10695 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		_w12045_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name10696 (
		\P3_EBX_reg[31]/NET0131 ,
		_w11952_,
		_w11988_,
		_w12045_,
		_w12046_
	);
	LUT3 #(
		.INIT('h21)
	) name10697 (
		\P3_EBX_reg[21]/NET0131 ,
		_w2187_,
		_w12046_,
		_w12047_
	);
	LUT4 #(
		.INIT('h8444)
	) name10698 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w2187_,
		_w11923_,
		_w12026_,
		_w12048_
	);
	LUT2 #(
		.INIT('h2)
	) name10699 (
		_w11831_,
		_w12048_,
		_w12049_
	);
	LUT4 #(
		.INIT('haa02)
	) name10700 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12050_
	);
	LUT4 #(
		.INIT('h8444)
	) name10701 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w11802_,
		_w11923_,
		_w12026_,
		_w12051_
	);
	LUT3 #(
		.INIT('h45)
	) name10702 (
		\P3_EBX_reg[21]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12052_
	);
	LUT4 #(
		.INIT('h0008)
	) name10703 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12052_,
		_w12053_
	);
	LUT3 #(
		.INIT('h45)
	) name10704 (
		_w12050_,
		_w12051_,
		_w12053_,
		_w12054_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10705 (
		_w1945_,
		_w12047_,
		_w12049_,
		_w12054_,
		_w12055_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10706 (
		\P3_PhyAddrPointer_reg[21]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12056_
	);
	LUT2 #(
		.INIT('h4)
	) name10707 (
		_w12055_,
		_w12056_,
		_w12057_
	);
	LUT2 #(
		.INIT('hb)
	) name10708 (
		_w12044_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h1)
	) name10709 (
		_w7469_,
		_w8032_,
		_w12059_
	);
	LUT2 #(
		.INIT('h8)
	) name10710 (
		_w12021_,
		_w12059_,
		_w12060_
	);
	LUT4 #(
		.INIT('h0514)
	) name10711 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7481_,
		_w12060_,
		_w12061_
	);
	LUT2 #(
		.INIT('h2)
	) name10712 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w12062_
	);
	LUT2 #(
		.INIT('h2)
	) name10713 (
		_w2194_,
		_w12062_,
		_w12063_
	);
	LUT4 #(
		.INIT('haa02)
	) name10714 (
		\P3_rEIP_reg[22]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12064_
	);
	LUT3 #(
		.INIT('h45)
	) name10715 (
		\P3_EBX_reg[22]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12065_
	);
	LUT3 #(
		.INIT('h08)
	) name10716 (
		_w2060_,
		_w2047_,
		_w12065_,
		_w12066_
	);
	LUT4 #(
		.INIT('h4000)
	) name10717 (
		\P3_EBX_reg[21]/NET0131 ,
		_w11952_,
		_w11988_,
		_w12045_,
		_w12067_
	);
	LUT4 #(
		.INIT('h0509)
	) name10718 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w12067_,
		_w12068_
	);
	LUT2 #(
		.INIT('h8)
	) name10719 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w12069_
	);
	LUT3 #(
		.INIT('h80)
	) name10720 (
		_w11923_,
		_w12026_,
		_w12069_,
		_w12070_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10721 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w11923_,
		_w12026_,
		_w12071_
	);
	LUT4 #(
		.INIT('h0080)
	) name10722 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w12065_,
		_w12072_
	);
	LUT4 #(
		.INIT('h5551)
	) name10723 (
		_w2105_,
		_w2187_,
		_w12071_,
		_w12072_,
		_w12073_
	);
	LUT4 #(
		.INIT('hce00)
	) name10724 (
		_w2106_,
		_w12066_,
		_w12068_,
		_w12073_,
		_w12074_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10725 (
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12075_
	);
	LUT4 #(
		.INIT('h5700)
	) name10726 (
		_w1945_,
		_w12064_,
		_w12074_,
		_w12075_,
		_w12076_
	);
	LUT3 #(
		.INIT('h4f)
	) name10727 (
		_w12061_,
		_w12063_,
		_w12076_,
		_w12077_
	);
	LUT3 #(
		.INIT('h40)
	) name10728 (
		_w7481_,
		_w12021_,
		_w12059_,
		_w12078_
	);
	LUT4 #(
		.INIT('h0514)
	) name10729 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w6943_,
		_w12078_,
		_w12079_
	);
	LUT2 #(
		.INIT('h2)
	) name10730 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w12080_
	);
	LUT2 #(
		.INIT('h2)
	) name10731 (
		_w2194_,
		_w12080_,
		_w12081_
	);
	LUT2 #(
		.INIT('h4)
	) name10732 (
		_w12079_,
		_w12081_,
		_w12082_
	);
	LUT4 #(
		.INIT('haa02)
	) name10733 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12083_
	);
	LUT4 #(
		.INIT('h8000)
	) name10734 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w11923_,
		_w12026_,
		_w12069_,
		_w12084_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name10735 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w11923_,
		_w12026_,
		_w12069_,
		_w12085_
	);
	LUT3 #(
		.INIT('h45)
	) name10736 (
		\P3_EBX_reg[23]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12086_
	);
	LUT3 #(
		.INIT('h08)
	) name10737 (
		_w2060_,
		_w2047_,
		_w12086_,
		_w12087_
	);
	LUT3 #(
		.INIT('hd0)
	) name10738 (
		_w11802_,
		_w12085_,
		_w12087_,
		_w12088_
	);
	LUT3 #(
		.INIT('h8c)
	) name10739 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12067_,
		_w12089_
	);
	LUT3 #(
		.INIT('ha2)
	) name10740 (
		_w2106_,
		_w2187_,
		_w12085_,
		_w12090_
	);
	LUT4 #(
		.INIT('hde00)
	) name10741 (
		\P3_EBX_reg[23]/NET0131 ,
		_w2187_,
		_w12089_,
		_w12090_,
		_w12091_
	);
	LUT4 #(
		.INIT('h2223)
	) name10742 (
		_w2105_,
		_w12083_,
		_w12088_,
		_w12091_,
		_w12092_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10743 (
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12093_
	);
	LUT3 #(
		.INIT('hd0)
	) name10744 (
		_w1945_,
		_w12092_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('hb)
	) name10745 (
		_w12082_,
		_w12094_,
		_w12095_
	);
	LUT4 #(
		.INIT('h8103)
	) name10746 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[22]/NET0131 ,
		\P3_PhyAddrPointer_reg[23]/NET0131 ,
		_w5771_,
		_w12096_
	);
	LUT3 #(
		.INIT('h80)
	) name10747 (
		_w12021_,
		_w12059_,
		_w12096_,
		_w12097_
	);
	LUT4 #(
		.INIT('h0514)
	) name10748 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w7496_,
		_w12097_,
		_w12098_
	);
	LUT2 #(
		.INIT('h2)
	) name10749 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w12099_
	);
	LUT2 #(
		.INIT('h2)
	) name10750 (
		_w2194_,
		_w12099_,
		_w12100_
	);
	LUT2 #(
		.INIT('h1)
	) name10751 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[23]/NET0131 ,
		_w12101_
	);
	LUT3 #(
		.INIT('h2a)
	) name10752 (
		\P3_EBX_reg[31]/NET0131 ,
		_w12067_,
		_w12101_,
		_w12102_
	);
	LUT4 #(
		.INIT('h70b0)
	) name10753 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2187_,
		_w11831_,
		_w12084_,
		_w12103_
	);
	LUT4 #(
		.INIT('hde00)
	) name10754 (
		\P3_EBX_reg[24]/NET0131 ,
		_w2187_,
		_w12102_,
		_w12103_,
		_w12104_
	);
	LUT4 #(
		.INIT('h3222)
	) name10755 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[24]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12105_
	);
	LUT3 #(
		.INIT('h01)
	) name10756 (
		_w2111_,
		_w2105_,
		_w12105_,
		_w12106_
	);
	LUT4 #(
		.INIT('h7b00)
	) name10757 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2187_,
		_w12084_,
		_w12106_,
		_w12107_
	);
	LUT4 #(
		.INIT('h335f)
	) name10758 (
		\P3_EBX_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w2111_,
		_w2105_,
		_w12108_
	);
	LUT2 #(
		.INIT('h8)
	) name10759 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w11949_,
		_w12109_
	);
	LUT4 #(
		.INIT('h0075)
	) name10760 (
		_w2113_,
		_w12107_,
		_w12108_,
		_w12109_,
		_w12110_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10761 (
		\P3_PhyAddrPointer_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12111_
	);
	LUT4 #(
		.INIT('h7500)
	) name10762 (
		_w1945_,
		_w12104_,
		_w12110_,
		_w12111_,
		_w12112_
	);
	LUT3 #(
		.INIT('h4f)
	) name10763 (
		_w12098_,
		_w12100_,
		_w12112_,
		_w12113_
	);
	LUT3 #(
		.INIT('hba)
	) name10764 (
		_w5779_,
		_w7496_,
		_w12097_,
		_w12114_
	);
	LUT2 #(
		.INIT('h2)
	) name10765 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w12115_
	);
	LUT2 #(
		.INIT('h2)
	) name10766 (
		_w2194_,
		_w12115_,
		_w12116_
	);
	LUT4 #(
		.INIT('heb00)
	) name10767 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w8041_,
		_w12114_,
		_w12116_,
		_w12117_
	);
	LUT2 #(
		.INIT('h8)
	) name10768 (
		\P3_rEIP_reg[23]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w12118_
	);
	LUT3 #(
		.INIT('h80)
	) name10769 (
		\P3_rEIP_reg[23]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w12119_
	);
	LUT4 #(
		.INIT('h8000)
	) name10770 (
		_w11923_,
		_w12026_,
		_w12069_,
		_w12119_,
		_w12120_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10771 (
		\P3_rEIP_reg[23]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w12070_,
		_w12121_
	);
	LUT4 #(
		.INIT('h3222)
	) name10772 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[25]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12122_
	);
	LUT3 #(
		.INIT('h01)
	) name10773 (
		_w2111_,
		_w2105_,
		_w12122_,
		_w12123_
	);
	LUT4 #(
		.INIT('h335f)
	) name10774 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w2111_,
		_w2105_,
		_w12124_
	);
	LUT4 #(
		.INIT('h2f00)
	) name10775 (
		_w2187_,
		_w12121_,
		_w12123_,
		_w12124_,
		_w12125_
	);
	LUT2 #(
		.INIT('h2)
	) name10776 (
		_w2113_,
		_w12125_,
		_w12126_
	);
	LUT2 #(
		.INIT('h8)
	) name10777 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w11949_,
		_w12127_
	);
	LUT3 #(
		.INIT('h01)
	) name10778 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[23]/NET0131 ,
		\P3_EBX_reg[24]/NET0131 ,
		_w12128_
	);
	LUT3 #(
		.INIT('h2a)
	) name10779 (
		\P3_EBX_reg[31]/NET0131 ,
		_w12067_,
		_w12128_,
		_w12129_
	);
	LUT3 #(
		.INIT('h21)
	) name10780 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2187_,
		_w12129_,
		_w12130_
	);
	LUT3 #(
		.INIT('hc4)
	) name10781 (
		_w2187_,
		_w11831_,
		_w12121_,
		_w12131_
	);
	LUT3 #(
		.INIT('h45)
	) name10782 (
		_w12127_,
		_w12130_,
		_w12131_,
		_w12132_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10783 (
		\P3_PhyAddrPointer_reg[25]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12133_
	);
	LUT4 #(
		.INIT('h7500)
	) name10784 (
		_w1945_,
		_w12126_,
		_w12132_,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('hb)
	) name10785 (
		_w12117_,
		_w12134_,
		_w12135_
	);
	LUT2 #(
		.INIT('h1)
	) name10786 (
		_w7496_,
		_w8041_,
		_w12136_
	);
	LUT3 #(
		.INIT('h15)
	) name10787 (
		_w5779_,
		_w12097_,
		_w12136_,
		_w12137_
	);
	LUT2 #(
		.INIT('h2)
	) name10788 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w12138_
	);
	LUT2 #(
		.INIT('h2)
	) name10789 (
		_w2194_,
		_w12138_,
		_w12139_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10790 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w7513_,
		_w12137_,
		_w12139_,
		_w12140_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name10791 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12067_,
		_w12128_,
		_w12141_
	);
	LUT4 #(
		.INIT('h70b0)
	) name10792 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2187_,
		_w11831_,
		_w12120_,
		_w12142_
	);
	LUT4 #(
		.INIT('hde00)
	) name10793 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2187_,
		_w12141_,
		_w12142_,
		_w12143_
	);
	LUT4 #(
		.INIT('haa02)
	) name10794 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12144_
	);
	LUT3 #(
		.INIT('h45)
	) name10795 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12145_
	);
	LUT4 #(
		.INIT('h0008)
	) name10796 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12145_,
		_w12146_
	);
	LUT4 #(
		.INIT('h7b00)
	) name10797 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w11802_,
		_w12120_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h1)
	) name10798 (
		_w12144_,
		_w12147_,
		_w12148_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10799 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12149_
	);
	LUT4 #(
		.INIT('h7500)
	) name10800 (
		_w1945_,
		_w12143_,
		_w12148_,
		_w12149_,
		_w12150_
	);
	LUT2 #(
		.INIT('hb)
	) name10801 (
		_w12140_,
		_w12150_,
		_w12151_
	);
	LUT4 #(
		.INIT('h4555)
	) name10802 (
		_w5779_,
		_w7513_,
		_w12097_,
		_w12136_,
		_w12152_
	);
	LUT2 #(
		.INIT('h2)
	) name10803 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w12153_
	);
	LUT2 #(
		.INIT('h2)
	) name10804 (
		_w2194_,
		_w12153_,
		_w12154_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10805 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6956_,
		_w12152_,
		_w12154_,
		_w12155_
	);
	LUT4 #(
		.INIT('h1000)
	) name10806 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		_w12067_,
		_w12128_,
		_w12156_
	);
	LUT4 #(
		.INIT('h0509)
	) name10807 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h8)
	) name10808 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w12158_
	);
	LUT4 #(
		.INIT('h9030)
	) name10809 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w2187_,
		_w12120_,
		_w12159_
	);
	LUT2 #(
		.INIT('h2)
	) name10810 (
		_w11831_,
		_w12159_,
		_w12160_
	);
	LUT2 #(
		.INIT('h8)
	) name10811 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w11949_,
		_w12161_
	);
	LUT4 #(
		.INIT('h60c0)
	) name10812 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w11802_,
		_w12120_,
		_w12162_
	);
	LUT3 #(
		.INIT('h8a)
	) name10813 (
		\P3_EBX_reg[27]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12163_
	);
	LUT2 #(
		.INIT('h1)
	) name10814 (
		_w2105_,
		_w12163_,
		_w12164_
	);
	LUT2 #(
		.INIT('h4)
	) name10815 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w2105_,
		_w12165_
	);
	LUT3 #(
		.INIT('h08)
	) name10816 (
		_w2060_,
		_w2047_,
		_w12165_,
		_w12166_
	);
	LUT4 #(
		.INIT('h1055)
	) name10817 (
		_w12161_,
		_w12162_,
		_w12164_,
		_w12166_,
		_w12167_
	);
	LUT4 #(
		.INIT('h20aa)
	) name10818 (
		_w1945_,
		_w12157_,
		_w12160_,
		_w12167_,
		_w12168_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10819 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12169_
	);
	LUT2 #(
		.INIT('h4)
	) name10820 (
		_w12168_,
		_w12169_,
		_w12170_
	);
	LUT2 #(
		.INIT('hb)
	) name10821 (
		_w12155_,
		_w12170_,
		_w12171_
	);
	LUT3 #(
		.INIT('h8c)
	) name10822 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12156_,
		_w12172_
	);
	LUT4 #(
		.INIT('h8444)
	) name10823 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w2187_,
		_w12120_,
		_w12158_,
		_w12173_
	);
	LUT2 #(
		.INIT('h2)
	) name10824 (
		_w11831_,
		_w12173_,
		_w12174_
	);
	LUT4 #(
		.INIT('hde00)
	) name10825 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2187_,
		_w12172_,
		_w12174_,
		_w12175_
	);
	LUT4 #(
		.INIT('h4888)
	) name10826 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w11802_,
		_w12120_,
		_w12158_,
		_w12176_
	);
	LUT3 #(
		.INIT('h8a)
	) name10827 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12177_
	);
	LUT2 #(
		.INIT('h1)
	) name10828 (
		_w2105_,
		_w12177_,
		_w12178_
	);
	LUT4 #(
		.INIT('h1311)
	) name10829 (
		_w2113_,
		_w11949_,
		_w12176_,
		_w12178_,
		_w12179_
	);
	LUT4 #(
		.INIT('h4440)
	) name10830 (
		_w2105_,
		_w2113_,
		_w12177_,
		_w12176_,
		_w12180_
	);
	LUT3 #(
		.INIT('h0d)
	) name10831 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w12179_,
		_w12180_,
		_w12181_
	);
	LUT3 #(
		.INIT('h8a)
	) name10832 (
		_w1945_,
		_w12175_,
		_w12181_,
		_w12182_
	);
	LUT4 #(
		.INIT('hc0c1)
	) name10833 (
		\P3_PhyAddrPointer_reg[26]/NET0131 ,
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		_w5775_,
		_w7512_,
		_w12183_
	);
	LUT4 #(
		.INIT('h1555)
	) name10834 (
		_w5779_,
		_w12097_,
		_w12136_,
		_w12183_,
		_w12184_
	);
	LUT2 #(
		.INIT('h2)
	) name10835 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w12185_
	);
	LUT2 #(
		.INIT('h2)
	) name10836 (
		_w2194_,
		_w12185_,
		_w12186_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10837 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6967_,
		_w12184_,
		_w12186_,
		_w12187_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10838 (
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12188_
	);
	LUT3 #(
		.INIT('hef)
	) name10839 (
		_w12182_,
		_w12187_,
		_w12188_,
		_w12189_
	);
	LUT2 #(
		.INIT('h1)
	) name10840 (
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		_w12190_
	);
	LUT3 #(
		.INIT('h2a)
	) name10841 (
		\P3_EBX_reg[31]/NET0131 ,
		_w12156_,
		_w12190_,
		_w12191_
	);
	LUT3 #(
		.INIT('h80)
	) name10842 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w12192_
	);
	LUT4 #(
		.INIT('h8000)
	) name10843 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w12193_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name10844 (
		\P3_rEIP_reg[28]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w12120_,
		_w12158_,
		_w12194_
	);
	LUT3 #(
		.INIT('hc4)
	) name10845 (
		_w2187_,
		_w11831_,
		_w12194_,
		_w12195_
	);
	LUT4 #(
		.INIT('hde00)
	) name10846 (
		\P3_EBX_reg[29]/NET0131 ,
		_w2187_,
		_w12191_,
		_w12195_,
		_w12196_
	);
	LUT2 #(
		.INIT('h8)
	) name10847 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w11949_,
		_w12197_
	);
	LUT3 #(
		.INIT('h8a)
	) name10848 (
		\P3_EBX_reg[29]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12198_
	);
	LUT2 #(
		.INIT('h1)
	) name10849 (
		_w2105_,
		_w12198_,
		_w12199_
	);
	LUT2 #(
		.INIT('h4)
	) name10850 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w2105_,
		_w12200_
	);
	LUT3 #(
		.INIT('h08)
	) name10851 (
		_w2060_,
		_w2047_,
		_w12200_,
		_w12201_
	);
	LUT4 #(
		.INIT('h8f00)
	) name10852 (
		_w11802_,
		_w12194_,
		_w12199_,
		_w12201_,
		_w12202_
	);
	LUT2 #(
		.INIT('h1)
	) name10853 (
		_w12197_,
		_w12202_,
		_w12203_
	);
	LUT3 #(
		.INIT('h8a)
	) name10854 (
		_w1945_,
		_w12196_,
		_w12203_,
		_w12204_
	);
	LUT2 #(
		.INIT('h4)
	) name10855 (
		_w6967_,
		_w12183_,
		_w12205_
	);
	LUT4 #(
		.INIT('h1555)
	) name10856 (
		_w5779_,
		_w12097_,
		_w12136_,
		_w12205_,
		_w12206_
	);
	LUT2 #(
		.INIT('h2)
	) name10857 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w12207_
	);
	LUT2 #(
		.INIT('h2)
	) name10858 (
		_w2194_,
		_w12207_,
		_w12208_
	);
	LUT4 #(
		.INIT('hbe00)
	) name10859 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6985_,
		_w12206_,
		_w12208_,
		_w12209_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10860 (
		\P3_PhyAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12210_
	);
	LUT3 #(
		.INIT('hef)
	) name10861 (
		_w12204_,
		_w12209_,
		_w12210_,
		_w12211_
	);
	LUT2 #(
		.INIT('h4)
	) name10862 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w12212_
	);
	LUT2 #(
		.INIT('h6)
	) name10863 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w12213_
	);
	LUT4 #(
		.INIT('h0154)
	) name10864 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w12212_,
		_w12213_,
		_w12214_
	);
	LUT2 #(
		.INIT('h2)
	) name10865 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w12215_
	);
	LUT2 #(
		.INIT('h2)
	) name10866 (
		_w2194_,
		_w12215_,
		_w12216_
	);
	LUT4 #(
		.INIT('haa02)
	) name10867 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12217_
	);
	LUT3 #(
		.INIT('h14)
	) name10868 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w12218_
	);
	LUT2 #(
		.INIT('h4)
	) name10869 (
		_w2116_,
		_w12218_,
		_w12219_
	);
	LUT3 #(
		.INIT('he0)
	) name10870 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12220_
	);
	LUT3 #(
		.INIT('h12)
	) name10871 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2187_,
		_w12220_,
		_w12221_
	);
	LUT2 #(
		.INIT('h1)
	) name10872 (
		_w12219_,
		_w12221_,
		_w12222_
	);
	LUT3 #(
		.INIT('h04)
	) name10873 (
		_w2060_,
		_w2047_,
		_w12222_,
		_w12223_
	);
	LUT2 #(
		.INIT('h8)
	) name10874 (
		_w2044_,
		_w2140_,
		_w12224_
	);
	LUT3 #(
		.INIT('h8a)
	) name10875 (
		\P3_EBX_reg[2]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12225_
	);
	LUT3 #(
		.INIT('h10)
	) name10876 (
		_w2111_,
		_w2116_,
		_w12218_,
		_w12226_
	);
	LUT2 #(
		.INIT('h1)
	) name10877 (
		_w12225_,
		_w12226_,
		_w12227_
	);
	LUT3 #(
		.INIT('h08)
	) name10878 (
		_w2060_,
		_w2047_,
		_w12227_,
		_w12228_
	);
	LUT4 #(
		.INIT('h5554)
	) name10879 (
		_w2105_,
		_w12224_,
		_w12228_,
		_w12223_,
		_w12229_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10880 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12230_
	);
	LUT4 #(
		.INIT('h5700)
	) name10881 (
		_w1945_,
		_w12217_,
		_w12229_,
		_w12230_,
		_w12231_
	);
	LUT3 #(
		.INIT('h4f)
	) name10882 (
		_w12214_,
		_w12216_,
		_w12231_,
		_w12232_
	);
	LUT4 #(
		.INIT('hc888)
	) name10883 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w12233_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		\P3_EBX_reg[29]/NET0131 ,
		\P3_EBX_reg[30]/NET0131 ,
		_w12234_
	);
	LUT2 #(
		.INIT('h8)
	) name10885 (
		_w12233_,
		_w12234_,
		_w12235_
	);
	LUT3 #(
		.INIT('h80)
	) name10886 (
		_w12156_,
		_w12190_,
		_w12235_,
		_w12236_
	);
	LUT3 #(
		.INIT('h80)
	) name10887 (
		\P3_rEIP_reg[30]/NET0131 ,
		_w12120_,
		_w12193_,
		_w12237_
	);
	LUT3 #(
		.INIT('h48)
	) name10888 (
		\P3_rEIP_reg[31]/NET0131 ,
		_w2187_,
		_w12237_,
		_w12238_
	);
	LUT3 #(
		.INIT('ha8)
	) name10889 (
		_w2106_,
		_w12236_,
		_w12238_,
		_w12239_
	);
	LUT4 #(
		.INIT('hc535)
	) name10890 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w2187_,
		_w12237_,
		_w12240_
	);
	LUT3 #(
		.INIT('h08)
	) name10891 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w12241_
	);
	LUT2 #(
		.INIT('h4)
	) name10892 (
		_w12240_,
		_w12241_,
		_w12242_
	);
	LUT4 #(
		.INIT('haa02)
	) name10893 (
		\P3_rEIP_reg[31]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12243_
	);
	LUT4 #(
		.INIT('h0080)
	) name10894 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w2105_,
		_w12244_
	);
	LUT3 #(
		.INIT('h13)
	) name10895 (
		\P3_EBX_reg[31]/NET0131 ,
		_w12243_,
		_w12244_,
		_w12245_
	);
	LUT4 #(
		.INIT('hab00)
	) name10896 (
		_w2105_,
		_w12239_,
		_w12242_,
		_w12245_,
		_w12246_
	);
	LUT2 #(
		.INIT('h8)
	) name10897 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w12247_
	);
	LUT3 #(
		.INIT('h81)
	) name10898 (
		\P3_PhyAddrPointer_reg[27]/NET0131 ,
		\P3_PhyAddrPointer_reg[28]/NET0131 ,
		_w5775_,
		_w12248_
	);
	LUT3 #(
		.INIT('h10)
	) name10899 (
		_w6348_,
		_w6985_,
		_w12248_,
		_w12249_
	);
	LUT4 #(
		.INIT('h4000)
	) name10900 (
		_w7513_,
		_w12097_,
		_w12136_,
		_w12249_,
		_w12250_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name10901 (
		_w2194_,
		_w5780_,
		_w12247_,
		_w12250_,
		_w12251_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10902 (
		\P3_PhyAddrPointer_reg[31]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12252_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name10903 (
		_w1945_,
		_w12246_,
		_w12251_,
		_w12252_,
		_w12253_
	);
	LUT3 #(
		.INIT('h40)
	) name10904 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w12254_
	);
	LUT4 #(
		.INIT('h0514)
	) name10905 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w9586_,
		_w12254_,
		_w12255_
	);
	LUT2 #(
		.INIT('h2)
	) name10906 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w12256_
	);
	LUT2 #(
		.INIT('h2)
	) name10907 (
		_w2194_,
		_w12256_,
		_w12257_
	);
	LUT4 #(
		.INIT('haa02)
	) name10908 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12258_
	);
	LUT3 #(
		.INIT('h8a)
	) name10909 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12259_
	);
	LUT4 #(
		.INIT('h1540)
	) name10910 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w12260_
	);
	LUT3 #(
		.INIT('h10)
	) name10911 (
		_w2111_,
		_w2116_,
		_w12260_,
		_w12261_
	);
	LUT2 #(
		.INIT('h1)
	) name10912 (
		_w12259_,
		_w12261_,
		_w12262_
	);
	LUT3 #(
		.INIT('h08)
	) name10913 (
		_w2060_,
		_w2047_,
		_w12262_,
		_w12263_
	);
	LUT2 #(
		.INIT('h2)
	) name10914 (
		_w2044_,
		_w2156_,
		_w12264_
	);
	LUT4 #(
		.INIT('hfe00)
	) name10915 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w12265_
	);
	LUT3 #(
		.INIT('h12)
	) name10916 (
		\P3_EBX_reg[3]/NET0131 ,
		_w2187_,
		_w12265_,
		_w12266_
	);
	LUT2 #(
		.INIT('h4)
	) name10917 (
		_w2116_,
		_w12260_,
		_w12267_
	);
	LUT2 #(
		.INIT('h1)
	) name10918 (
		_w12266_,
		_w12267_,
		_w12268_
	);
	LUT3 #(
		.INIT('h04)
	) name10919 (
		_w2060_,
		_w2047_,
		_w12268_,
		_w12269_
	);
	LUT4 #(
		.INIT('h5554)
	) name10920 (
		_w2105_,
		_w12264_,
		_w12269_,
		_w12263_,
		_w12270_
	);
	LUT4 #(
		.INIT('h5f13)
	) name10921 (
		\P3_PhyAddrPointer_reg[3]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12271_
	);
	LUT4 #(
		.INIT('h5700)
	) name10922 (
		_w1945_,
		_w12258_,
		_w12270_,
		_w12271_,
		_w12272_
	);
	LUT3 #(
		.INIT('h4f)
	) name10923 (
		_w12255_,
		_w12257_,
		_w12272_,
		_w12273_
	);
	LUT3 #(
		.INIT('hdc)
	) name10924 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w5779_,
		_w9360_,
		_w12274_
	);
	LUT2 #(
		.INIT('h2)
	) name10925 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w12275_
	);
	LUT2 #(
		.INIT('h2)
	) name10926 (
		_w2194_,
		_w12275_,
		_w12276_
	);
	LUT4 #(
		.INIT('heb00)
	) name10927 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9362_,
		_w12274_,
		_w12276_,
		_w12277_
	);
	LUT2 #(
		.INIT('h2)
	) name10928 (
		\P3_EBX_reg[31]/NET0131 ,
		_w11811_,
		_w12278_
	);
	LUT4 #(
		.INIT('hf700)
	) name10929 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w12278_,
		_w12279_
	);
	LUT3 #(
		.INIT('h02)
	) name10930 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		_w11811_,
		_w12280_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name10931 (
		_w2060_,
		_w2047_,
		_w2187_,
		_w12280_,
		_w12281_
	);
	LUT4 #(
		.INIT('h7f80)
	) name10932 (
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w12282_
	);
	LUT2 #(
		.INIT('h2)
	) name10933 (
		_w2187_,
		_w12282_,
		_w12283_
	);
	LUT2 #(
		.INIT('h1)
	) name10934 (
		_w2105_,
		_w12283_,
		_w12284_
	);
	LUT4 #(
		.INIT('h4c00)
	) name10935 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w12284_,
		_w12285_
	);
	LUT4 #(
		.INIT('h2f00)
	) name10936 (
		\P3_EBX_reg[4]/NET0131 ,
		_w12279_,
		_w12281_,
		_w12285_,
		_w12286_
	);
	LUT4 #(
		.INIT('haa02)
	) name10937 (
		\P3_rEIP_reg[4]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12287_
	);
	LUT3 #(
		.INIT('h07)
	) name10938 (
		\P3_EBX_reg[4]/NET0131 ,
		_w12244_,
		_w12287_,
		_w12288_
	);
	LUT2 #(
		.INIT('h2)
	) name10939 (
		\P3_rEIP_reg[4]/NET0131 ,
		_w11818_,
		_w12289_
	);
	LUT3 #(
		.INIT('h07)
	) name10940 (
		\P3_PhyAddrPointer_reg[4]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12290_
	);
	LUT2 #(
		.INIT('h4)
	) name10941 (
		_w12289_,
		_w12290_,
		_w12291_
	);
	LUT4 #(
		.INIT('h7500)
	) name10942 (
		_w1945_,
		_w12286_,
		_w12288_,
		_w12291_,
		_w12292_
	);
	LUT2 #(
		.INIT('hb)
	) name10943 (
		_w12277_,
		_w12292_,
		_w12293_
	);
	LUT3 #(
		.INIT('h40)
	) name10944 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5758_,
		_w12294_
	);
	LUT4 #(
		.INIT('h0514)
	) name10945 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w9613_,
		_w12294_,
		_w12295_
	);
	LUT2 #(
		.INIT('h2)
	) name10946 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w12296_
	);
	LUT2 #(
		.INIT('h2)
	) name10947 (
		_w2194_,
		_w12296_,
		_w12297_
	);
	LUT3 #(
		.INIT('h6c)
	) name10948 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w11803_,
		_w12298_
	);
	LUT3 #(
		.INIT('he2)
	) name10949 (
		\P3_EBX_reg[6]/NET0131 ,
		_w11802_,
		_w12298_,
		_w12299_
	);
	LUT4 #(
		.INIT('h0800)
	) name10950 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12299_,
		_w12300_
	);
	LUT4 #(
		.INIT('haa02)
	) name10951 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12301_
	);
	LUT4 #(
		.INIT('h9030)
	) name10952 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w2187_,
		_w11803_,
		_w12302_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name10953 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		_w11811_,
		_w12303_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name10954 (
		\P3_EBX_reg[6]/NET0131 ,
		_w2187_,
		_w12302_,
		_w12303_,
		_w12304_
	);
	LUT4 #(
		.INIT('h0400)
	) name10955 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12304_,
		_w12305_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10956 (
		_w1945_,
		_w12301_,
		_w12305_,
		_w12300_,
		_w12306_
	);
	LUT2 #(
		.INIT('h2)
	) name10957 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w11818_,
		_w12307_
	);
	LUT3 #(
		.INIT('h07)
	) name10958 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12308_
	);
	LUT2 #(
		.INIT('h4)
	) name10959 (
		_w12307_,
		_w12308_,
		_w12309_
	);
	LUT2 #(
		.INIT('h4)
	) name10960 (
		_w12306_,
		_w12309_,
		_w12310_
	);
	LUT3 #(
		.INIT('h4f)
	) name10961 (
		_w12295_,
		_w12297_,
		_w12310_,
		_w12311_
	);
	LUT4 #(
		.INIT('h0514)
	) name10962 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8683_,
		_w11796_,
		_w12312_
	);
	LUT2 #(
		.INIT('h2)
	) name10963 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w12313_
	);
	LUT2 #(
		.INIT('h2)
	) name10964 (
		_w2194_,
		_w12313_,
		_w12314_
	);
	LUT4 #(
		.INIT('h78f0)
	) name10965 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w11803_,
		_w12315_
	);
	LUT3 #(
		.INIT('he2)
	) name10966 (
		\P3_EBX_reg[7]/NET0131 ,
		_w11802_,
		_w12315_,
		_w12316_
	);
	LUT4 #(
		.INIT('h0800)
	) name10967 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12316_,
		_w12317_
	);
	LUT4 #(
		.INIT('haa02)
	) name10968 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12318_
	);
	LUT2 #(
		.INIT('h2)
	) name10969 (
		_w2187_,
		_w12315_,
		_w12319_
	);
	LUT4 #(
		.INIT('h0309)
	) name10970 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		_w2187_,
		_w11812_,
		_w12320_
	);
	LUT2 #(
		.INIT('h1)
	) name10971 (
		_w12319_,
		_w12320_,
		_w12321_
	);
	LUT4 #(
		.INIT('h0400)
	) name10972 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12321_,
		_w12322_
	);
	LUT4 #(
		.INIT('haaa8)
	) name10973 (
		_w1945_,
		_w12318_,
		_w12322_,
		_w12317_,
		_w12323_
	);
	LUT2 #(
		.INIT('h2)
	) name10974 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w11818_,
		_w12324_
	);
	LUT3 #(
		.INIT('h07)
	) name10975 (
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12325_
	);
	LUT2 #(
		.INIT('h4)
	) name10976 (
		_w12324_,
		_w12325_,
		_w12326_
	);
	LUT2 #(
		.INIT('h4)
	) name10977 (
		_w12323_,
		_w12326_,
		_w12327_
	);
	LUT3 #(
		.INIT('h4f)
	) name10978 (
		_w12312_,
		_w12314_,
		_w12327_,
		_w12328_
	);
	LUT4 #(
		.INIT('h8000)
	) name10979 (
		\P3_PhyAddrPointer_reg[6]/NET0131 ,
		\P3_PhyAddrPointer_reg[7]/NET0131 ,
		_w5758_,
		_w12212_,
		_w12329_
	);
	LUT4 #(
		.INIT('h0514)
	) name10980 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8053_,
		_w12329_,
		_w12330_
	);
	LUT2 #(
		.INIT('h2)
	) name10981 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w12331_
	);
	LUT2 #(
		.INIT('h2)
	) name10982 (
		_w2194_,
		_w12331_,
		_w12332_
	);
	LUT4 #(
		.INIT('haa02)
	) name10983 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12333_
	);
	LUT3 #(
		.INIT('h84)
	) name10984 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w2187_,
		_w11804_,
		_w12334_
	);
	LUT3 #(
		.INIT('h45)
	) name10985 (
		\P3_EBX_reg[8]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12335_
	);
	LUT3 #(
		.INIT('h8a)
	) name10986 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		_w11812_,
		_w12336_
	);
	LUT3 #(
		.INIT('h21)
	) name10987 (
		\P3_EBX_reg[8]/NET0131 ,
		_w2187_,
		_w12336_,
		_w12337_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name10988 (
		_w2060_,
		_w2047_,
		_w12335_,
		_w12337_,
		_w12338_
	);
	LUT4 #(
		.INIT('h0080)
	) name10989 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w12335_,
		_w12339_
	);
	LUT4 #(
		.INIT('h5501)
	) name10990 (
		_w2105_,
		_w12334_,
		_w12338_,
		_w12339_,
		_w12340_
	);
	LUT2 #(
		.INIT('h2)
	) name10991 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w11818_,
		_w12341_
	);
	LUT3 #(
		.INIT('h07)
	) name10992 (
		\P3_PhyAddrPointer_reg[8]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12342_
	);
	LUT2 #(
		.INIT('h4)
	) name10993 (
		_w12341_,
		_w12342_,
		_w12343_
	);
	LUT4 #(
		.INIT('h5700)
	) name10994 (
		_w1945_,
		_w12333_,
		_w12340_,
		_w12343_,
		_w12344_
	);
	LUT3 #(
		.INIT('h4f)
	) name10995 (
		_w12330_,
		_w12332_,
		_w12344_,
		_w12345_
	);
	LUT3 #(
		.INIT('h40)
	) name10996 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w5760_,
		_w12346_
	);
	LUT4 #(
		.INIT('h0514)
	) name10997 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w5779_,
		_w8694_,
		_w12346_,
		_w12347_
	);
	LUT2 #(
		.INIT('h2)
	) name10998 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w12348_
	);
	LUT2 #(
		.INIT('h2)
	) name10999 (
		_w2194_,
		_w12348_,
		_w12349_
	);
	LUT4 #(
		.INIT('haa02)
	) name11000 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12350_
	);
	LUT4 #(
		.INIT('h9030)
	) name11001 (
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w2187_,
		_w11804_,
		_w12351_
	);
	LUT2 #(
		.INIT('h4)
	) name11002 (
		_w2111_,
		_w12351_,
		_w12352_
	);
	LUT3 #(
		.INIT('h45)
	) name11003 (
		\P3_EBX_reg[9]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12353_
	);
	LUT4 #(
		.INIT('h0008)
	) name11004 (
		_w2060_,
		_w2047_,
		_w12352_,
		_w12353_,
		_w12354_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11005 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		_w11812_,
		_w12355_
	);
	LUT3 #(
		.INIT('h21)
	) name11006 (
		\P3_EBX_reg[9]/NET0131 ,
		_w2187_,
		_w12355_,
		_w12356_
	);
	LUT4 #(
		.INIT('h0004)
	) name11007 (
		_w2060_,
		_w2047_,
		_w12351_,
		_w12356_,
		_w12357_
	);
	LUT4 #(
		.INIT('h2223)
	) name11008 (
		_w2105_,
		_w12350_,
		_w12354_,
		_w12357_,
		_w12358_
	);
	LUT2 #(
		.INIT('h2)
	) name11009 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w11818_,
		_w12359_
	);
	LUT3 #(
		.INIT('h07)
	) name11010 (
		\P3_PhyAddrPointer_reg[9]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12360_
	);
	LUT2 #(
		.INIT('h4)
	) name11011 (
		_w12359_,
		_w12360_,
		_w12361_
	);
	LUT3 #(
		.INIT('hd0)
	) name11012 (
		_w1945_,
		_w12358_,
		_w12361_,
		_w12362_
	);
	LUT3 #(
		.INIT('h4f)
	) name11013 (
		_w12347_,
		_w12349_,
		_w12362_,
		_w12363_
	);
	LUT3 #(
		.INIT('h80)
	) name11014 (
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w6367_,
		_w10801_,
		_w12364_
	);
	LUT3 #(
		.INIT('h06)
	) name11015 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w12364_,
		_w12365_
	);
	LUT2 #(
		.INIT('h2)
	) name11016 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		_w12366_
	);
	LUT2 #(
		.INIT('h2)
	) name11017 (
		_w1939_,
		_w12366_,
		_w12367_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11018 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8706_,
		_w12365_,
		_w12367_,
		_w12368_
	);
	LUT2 #(
		.INIT('h2)
	) name11019 (
		\P1_rEIP_reg[10]/NET0131 ,
		_w10808_,
		_w12369_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name11020 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w10811_,
		_w12370_
	);
	LUT2 #(
		.INIT('h2)
	) name11021 (
		_w10817_,
		_w12370_,
		_w12371_
	);
	LUT4 #(
		.INIT('h3332)
	) name11022 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[10]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12372_
	);
	LUT3 #(
		.INIT('h02)
	) name11023 (
		_w1797_,
		_w12372_,
		_w12371_,
		_w12373_
	);
	LUT4 #(
		.INIT('h0509)
	) name11024 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w10822_,
		_w12374_
	);
	LUT2 #(
		.INIT('h2)
	) name11025 (
		_w1930_,
		_w12370_,
		_w12375_
	);
	LUT3 #(
		.INIT('h02)
	) name11026 (
		_w1795_,
		_w12375_,
		_w12374_,
		_w12376_
	);
	LUT3 #(
		.INIT('h54)
	) name11027 (
		_w1852_,
		_w12373_,
		_w12376_,
		_w12377_
	);
	LUT2 #(
		.INIT('h2)
	) name11028 (
		\P1_rEIP_reg[10]/NET0131 ,
		_w10828_,
		_w12378_
	);
	LUT3 #(
		.INIT('h07)
	) name11029 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		_w2234_,
		_w3406_,
		_w12379_
	);
	LUT2 #(
		.INIT('h4)
	) name11030 (
		_w12378_,
		_w12379_,
		_w12380_
	);
	LUT4 #(
		.INIT('h5700)
	) name11031 (
		_w1933_,
		_w12369_,
		_w12377_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('hb)
	) name11032 (
		_w12368_,
		_w12381_,
		_w12382_
	);
	LUT4 #(
		.INIT('h8000)
	) name11033 (
		\P1_PhyAddrPointer_reg[10]/NET0131 ,
		\P1_PhyAddrPointer_reg[9]/NET0131 ,
		_w6367_,
		_w10801_,
		_w12383_
	);
	LUT3 #(
		.INIT('h06)
	) name11034 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w12383_,
		_w12384_
	);
	LUT2 #(
		.INIT('h2)
	) name11035 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w12385_
	);
	LUT2 #(
		.INIT('h2)
	) name11036 (
		_w1939_,
		_w12385_,
		_w12386_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11037 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w7531_,
		_w12384_,
		_w12386_,
		_w12387_
	);
	LUT2 #(
		.INIT('h2)
	) name11038 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10808_,
		_w12388_
	);
	LUT3 #(
		.INIT('h84)
	) name11039 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10817_,
		_w10812_,
		_w12389_
	);
	LUT4 #(
		.INIT('h3332)
	) name11040 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12390_
	);
	LUT3 #(
		.INIT('h02)
	) name11041 (
		_w1797_,
		_w12390_,
		_w12389_,
		_w12391_
	);
	LUT3 #(
		.INIT('h8c)
	) name11042 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10822_,
		_w12392_
	);
	LUT3 #(
		.INIT('h21)
	) name11043 (
		\P1_EBX_reg[11]/NET0131 ,
		_w1930_,
		_w12392_,
		_w12393_
	);
	LUT3 #(
		.INIT('h84)
	) name11044 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w1930_,
		_w10812_,
		_w12394_
	);
	LUT3 #(
		.INIT('h02)
	) name11045 (
		_w1795_,
		_w12394_,
		_w12393_,
		_w12395_
	);
	LUT3 #(
		.INIT('h54)
	) name11046 (
		_w1852_,
		_w12391_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h2)
	) name11047 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10828_,
		_w12397_
	);
	LUT3 #(
		.INIT('h07)
	) name11048 (
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w2234_,
		_w3406_,
		_w12398_
	);
	LUT2 #(
		.INIT('h4)
	) name11049 (
		_w12397_,
		_w12398_,
		_w12399_
	);
	LUT4 #(
		.INIT('h5700)
	) name11050 (
		_w1933_,
		_w12388_,
		_w12396_,
		_w12399_,
		_w12400_
	);
	LUT2 #(
		.INIT('hb)
	) name11051 (
		_w12387_,
		_w12400_,
		_w12401_
	);
	LUT3 #(
		.INIT('h40)
	) name11052 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		\P1_PhyAddrPointer_reg[11]/NET0131 ,
		_w7530_,
		_w12402_
	);
	LUT3 #(
		.INIT('h06)
	) name11053 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w12402_,
		_w12403_
	);
	LUT2 #(
		.INIT('h2)
	) name11054 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w12404_
	);
	LUT2 #(
		.INIT('h2)
	) name11055 (
		_w1939_,
		_w12404_,
		_w12405_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11056 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8064_,
		_w12403_,
		_w12405_,
		_w12406_
	);
	LUT2 #(
		.INIT('h2)
	) name11057 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w10808_,
		_w12407_
	);
	LUT4 #(
		.INIT('h9030)
	) name11058 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w1930_,
		_w10812_,
		_w12408_
	);
	LUT2 #(
		.INIT('h4)
	) name11059 (
		_w1858_,
		_w12408_,
		_w12409_
	);
	LUT4 #(
		.INIT('h3332)
	) name11060 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[12]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12410_
	);
	LUT3 #(
		.INIT('h02)
	) name11061 (
		_w1797_,
		_w12410_,
		_w12409_,
		_w12411_
	);
	LUT4 #(
		.INIT('he0f0)
	) name11062 (
		\P1_EBX_reg[10]/NET0131 ,
		\P1_EBX_reg[11]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w10822_,
		_w12412_
	);
	LUT3 #(
		.INIT('h21)
	) name11063 (
		\P1_EBX_reg[12]/NET0131 ,
		_w1930_,
		_w12412_,
		_w12413_
	);
	LUT3 #(
		.INIT('h02)
	) name11064 (
		_w1795_,
		_w12408_,
		_w12413_,
		_w12414_
	);
	LUT3 #(
		.INIT('h54)
	) name11065 (
		_w1852_,
		_w12411_,
		_w12414_,
		_w12415_
	);
	LUT2 #(
		.INIT('h2)
	) name11066 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w10828_,
		_w12416_
	);
	LUT3 #(
		.INIT('h07)
	) name11067 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w2234_,
		_w3406_,
		_w12417_
	);
	LUT2 #(
		.INIT('h4)
	) name11068 (
		_w12416_,
		_w12417_,
		_w12418_
	);
	LUT4 #(
		.INIT('h5700)
	) name11069 (
		_w1933_,
		_w12407_,
		_w12415_,
		_w12418_,
		_w12419_
	);
	LUT2 #(
		.INIT('hb)
	) name11070 (
		_w12406_,
		_w12419_,
		_w12420_
	);
	LUT3 #(
		.INIT('h80)
	) name11071 (
		\P1_PhyAddrPointer_reg[12]/NET0131 ,
		_w6368_,
		_w10802_,
		_w12421_
	);
	LUT3 #(
		.INIT('h06)
	) name11072 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w12421_,
		_w12422_
	);
	LUT2 #(
		.INIT('h2)
	) name11073 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w12423_
	);
	LUT2 #(
		.INIT('h2)
	) name11074 (
		_w1939_,
		_w12423_,
		_w12424_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11075 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w8079_,
		_w12422_,
		_w12424_,
		_w12425_
	);
	LUT2 #(
		.INIT('h2)
	) name11076 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w10808_,
		_w12426_
	);
	LUT4 #(
		.INIT('h78f0)
	) name11077 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w10812_,
		_w12427_
	);
	LUT2 #(
		.INIT('h2)
	) name11078 (
		_w1930_,
		_w12427_,
		_w12428_
	);
	LUT3 #(
		.INIT('h04)
	) name11079 (
		_w1858_,
		_w1930_,
		_w12427_,
		_w12429_
	);
	LUT4 #(
		.INIT('h3332)
	) name11080 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[13]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12430_
	);
	LUT3 #(
		.INIT('h02)
	) name11081 (
		_w1797_,
		_w12430_,
		_w12429_,
		_w12431_
	);
	LUT4 #(
		.INIT('h0509)
	) name11082 (
		\P1_EBX_reg[13]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1930_,
		_w10823_,
		_w12432_
	);
	LUT3 #(
		.INIT('h02)
	) name11083 (
		_w1795_,
		_w12428_,
		_w12432_,
		_w12433_
	);
	LUT3 #(
		.INIT('h54)
	) name11084 (
		_w1852_,
		_w12431_,
		_w12433_,
		_w12434_
	);
	LUT2 #(
		.INIT('h2)
	) name11085 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w10828_,
		_w12435_
	);
	LUT3 #(
		.INIT('h07)
	) name11086 (
		\P1_PhyAddrPointer_reg[13]/NET0131 ,
		_w2234_,
		_w3406_,
		_w12436_
	);
	LUT2 #(
		.INIT('h4)
	) name11087 (
		_w12435_,
		_w12436_,
		_w12437_
	);
	LUT4 #(
		.INIT('h5700)
	) name11088 (
		_w1933_,
		_w12426_,
		_w12434_,
		_w12437_,
		_w12438_
	);
	LUT2 #(
		.INIT('hb)
	) name11089 (
		_w12425_,
		_w12438_,
		_w12439_
	);
	LUT3 #(
		.INIT('h20)
	) name11090 (
		_w1559_,
		_w8333_,
		_w8334_,
		_w12440_
	);
	LUT3 #(
		.INIT('h80)
	) name11091 (
		_w1558_,
		_w1596_,
		_w8319_,
		_w12441_
	);
	LUT3 #(
		.INIT('h0d)
	) name11092 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w7642_,
		_w12441_,
		_w12442_
	);
	LUT4 #(
		.INIT('hf400)
	) name11093 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2283_,
		_w11597_,
		_w12443_
	);
	LUT2 #(
		.INIT('h2)
	) name11094 (
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w5747_,
		_w12444_
	);
	LUT3 #(
		.INIT('h20)
	) name11095 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[2]/NET0131 ,
		_w1679_,
		_w12445_
	);
	LUT4 #(
		.INIT('h0001)
	) name11096 (
		_w8337_,
		_w12445_,
		_w12443_,
		_w12444_,
		_w12446_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11097 (
		_w1678_,
		_w12440_,
		_w12442_,
		_w12446_,
		_w12447_
	);
	LUT3 #(
		.INIT('h04)
	) name11098 (
		\P2_RequestPending_reg/NET0131 ,
		_w1592_,
		_w1601_,
		_w12448_
	);
	LUT4 #(
		.INIT('h00fe)
	) name11099 (
		_w1607_,
		_w1613_,
		_w1603_,
		_w12448_,
		_w12449_
	);
	LUT4 #(
		.INIT('h0002)
	) name11100 (
		\P2_RequestPending_reg/NET0131 ,
		_w1565_,
		_w1566_,
		_w1568_,
		_w12450_
	);
	LUT3 #(
		.INIT('h04)
	) name11101 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12451_
	);
	LUT2 #(
		.INIT('h1)
	) name11102 (
		_w12450_,
		_w12451_,
		_w12452_
	);
	LUT2 #(
		.INIT('h2)
	) name11103 (
		\P2_RequestPending_reg/NET0131 ,
		_w7766_,
		_w12453_
	);
	LUT3 #(
		.INIT('h02)
	) name11104 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w12454_
	);
	LUT4 #(
		.INIT('hfff4)
	) name11105 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w12455_
	);
	LUT3 #(
		.INIT('h70)
	) name11106 (
		_w2210_,
		_w12454_,
		_w12455_,
		_w12456_
	);
	LUT2 #(
		.INIT('h4)
	) name11107 (
		_w12453_,
		_w12456_,
		_w12457_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11108 (
		_w1678_,
		_w12449_,
		_w12452_,
		_w12457_,
		_w12458_
	);
	LUT2 #(
		.INIT('h2)
	) name11109 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w7422_,
		_w12459_
	);
	LUT4 #(
		.INIT('h8000)
	) name11110 (
		_w2060_,
		_w2041_,
		_w2098_,
		_w8303_,
		_w12460_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11111 (
		_w2180_,
		_w8310_,
		_w8306_,
		_w12460_,
		_w12461_
	);
	LUT2 #(
		.INIT('h2)
	) name11112 (
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w5783_,
		_w12462_
	);
	LUT4 #(
		.INIT('hf400)
	) name11113 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w12213_,
		_w12463_
	);
	LUT3 #(
		.INIT('h20)
	) name11114 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[2]/NET0131 ,
		_w2194_,
		_w12464_
	);
	LUT4 #(
		.INIT('h0001)
	) name11115 (
		_w8314_,
		_w12463_,
		_w12464_,
		_w12462_,
		_w12465_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11116 (
		_w1945_,
		_w12459_,
		_w12461_,
		_w12465_,
		_w12466_
	);
	LUT3 #(
		.INIT('h40)
	) name11117 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2060_,
		_w2047_,
		_w12467_
	);
	LUT4 #(
		.INIT('h0004)
	) name11118 (
		_w2048_,
		_w2122_,
		_w2125_,
		_w12467_,
		_w12468_
	);
	LUT4 #(
		.INIT('h5551)
	) name11119 (
		_w2105_,
		_w2122_,
		_w2125_,
		_w12467_,
		_w12469_
	);
	LUT4 #(
		.INIT('hcc08)
	) name11120 (
		\P3_RequestPending_reg/NET0131 ,
		_w1945_,
		_w12468_,
		_w12469_,
		_w12470_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name11121 (
		\P3_RequestPending_reg/NET0131 ,
		_w2116_,
		_w8340_,
		_w9977_,
		_w12471_
	);
	LUT4 #(
		.INIT('hfff4)
	) name11122 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w12472_
	);
	LUT2 #(
		.INIT('h4)
	) name11123 (
		_w12471_,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('hb)
	) name11124 (
		_w12470_,
		_w12473_,
		_w12474_
	);
	LUT3 #(
		.INIT('h02)
	) name11125 (
		_w1923_,
		_w8281_,
		_w8285_,
		_w12475_
	);
	LUT3 #(
		.INIT('h0d)
	) name11126 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w7547_,
		_w8292_,
		_w12476_
	);
	LUT4 #(
		.INIT('hf400)
	) name11127 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3407_,
		_w11408_,
		_w12477_
	);
	LUT2 #(
		.INIT('h2)
	) name11128 (
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w6383_,
		_w12478_
	);
	LUT3 #(
		.INIT('h20)
	) name11129 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[2]/NET0131 ,
		_w1939_,
		_w12479_
	);
	LUT4 #(
		.INIT('h0001)
	) name11130 (
		_w8296_,
		_w12479_,
		_w12477_,
		_w12478_,
		_w12480_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11131 (
		_w1933_,
		_w12475_,
		_w12476_,
		_w12480_,
		_w12481_
	);
	LUT3 #(
		.INIT('h04)
	) name11132 (
		\P1_RequestPending_reg/NET0131 ,
		_w1842_,
		_w1851_,
		_w12482_
	);
	LUT4 #(
		.INIT('h0045)
	) name11133 (
		_w1803_,
		_w1866_,
		_w1867_,
		_w12482_,
		_w12483_
	);
	LUT4 #(
		.INIT('h0002)
	) name11134 (
		\P1_RequestPending_reg/NET0131 ,
		_w1795_,
		_w1797_,
		_w1802_,
		_w12484_
	);
	LUT3 #(
		.INIT('h04)
	) name11135 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1797_,
		_w1852_,
		_w12485_
	);
	LUT2 #(
		.INIT('h1)
	) name11136 (
		_w12484_,
		_w12485_,
		_w12486_
	);
	LUT4 #(
		.INIT('h80aa)
	) name11137 (
		\P1_RequestPending_reg/NET0131 ,
		_w1861_,
		_w1935_,
		_w9101_,
		_w12487_
	);
	LUT2 #(
		.INIT('h2)
	) name11138 (
		_w3544_,
		_w12487_,
		_w12488_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11139 (
		_w1933_,
		_w12483_,
		_w12486_,
		_w12488_,
		_w12489_
	);
	LUT4 #(
		.INIT('h080a)
	) name11140 (
		\P1_Datao_reg[20]/NET0131 ,
		_w1725_,
		_w1797_,
		_w1802_,
		_w12490_
	);
	LUT4 #(
		.INIT('hccdc)
	) name11141 (
		_w1725_,
		_w1797_,
		_w1802_,
		_w1859_,
		_w12491_
	);
	LUT4 #(
		.INIT('h8000)
	) name11142 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		\P1_EAX_reg[20]/NET0131 ,
		_w9483_,
		_w12492_
	);
	LUT4 #(
		.INIT('h78f0)
	) name11143 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		\P1_EAX_reg[20]/NET0131 ,
		_w9483_,
		_w12493_
	);
	LUT3 #(
		.INIT('he2)
	) name11144 (
		\P1_Datao_reg[20]/NET0131 ,
		_w1859_,
		_w12493_,
		_w12494_
	);
	LUT4 #(
		.INIT('ha888)
	) name11145 (
		_w1933_,
		_w12490_,
		_w12491_,
		_w12494_,
		_w12495_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11146 (
		\P1_Datao_reg[20]/NET0131 ,
		\P1_uWord_reg[4]/NET0131 ,
		_w1935_,
		_w9972_,
		_w12496_
	);
	LUT2 #(
		.INIT('hb)
	) name11147 (
		_w12495_,
		_w12496_,
		_w12497_
	);
	LUT3 #(
		.INIT('h6c)
	) name11148 (
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		_w9538_,
		_w12498_
	);
	LUT4 #(
		.INIT('h0800)
	) name11149 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12498_,
		_w12499_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name11150 (
		\datao[20]_pad ,
		_w2111_,
		_w2115_,
		_w12499_,
		_w12500_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11151 (
		\P3_uWord_reg[4]/NET0131 ,
		\datao[20]_pad ,
		_w9977_,
		_w9978_,
		_w12501_
	);
	LUT3 #(
		.INIT('h2f)
	) name11152 (
		_w1945_,
		_w12500_,
		_w12501_,
		_w12502_
	);
	LUT4 #(
		.INIT('h78f0)
	) name11153 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		\P2_EAX_reg[20]/NET0131 ,
		_w9458_,
		_w12503_
	);
	LUT2 #(
		.INIT('h1)
	) name11154 (
		_w1611_,
		_w12503_,
		_w12504_
	);
	LUT3 #(
		.INIT('h02)
	) name11155 (
		_w1566_,
		_w1602_,
		_w12504_,
		_w12505_
	);
	LUT4 #(
		.INIT('haaa2)
	) name11156 (
		\P2_Datao_reg[20]/NET0131 ,
		_w4927_,
		_w9989_,
		_w12505_,
		_w12506_
	);
	LUT3 #(
		.INIT('h80)
	) name11157 (
		_w1566_,
		_w1674_,
		_w12503_,
		_w12507_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11158 (
		\P2_Datao_reg[20]/NET0131 ,
		\P2_uWord_reg[4]/NET0131 ,
		_w9995_,
		_w9996_,
		_w12508_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11159 (
		_w1678_,
		_w12506_,
		_w12507_,
		_w12508_,
		_w12509_
	);
	LUT2 #(
		.INIT('h2)
	) name11160 (
		\P1_EAX_reg[25]/NET0131 ,
		_w9102_,
		_w12510_
	);
	LUT3 #(
		.INIT('h48)
	) name11161 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1827_,
		_w9434_,
		_w12511_
	);
	LUT3 #(
		.INIT('h08)
	) name11162 (
		_w1725_,
		_w1802_,
		_w3519_,
		_w12512_
	);
	LUT2 #(
		.INIT('h2)
	) name11163 (
		_w1795_,
		_w3445_,
		_w12513_
	);
	LUT4 #(
		.INIT('h08a2)
	) name11164 (
		_w1846_,
		_w9015_,
		_w9026_,
		_w9037_,
		_w12514_
	);
	LUT4 #(
		.INIT('h4000)
	) name11165 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w12514_,
		_w12515_
	);
	LUT4 #(
		.INIT('h0057)
	) name11166 (
		_w1867_,
		_w12512_,
		_w12513_,
		_w12515_,
		_w12516_
	);
	LUT4 #(
		.INIT('h7500)
	) name11167 (
		\P1_EAX_reg[25]/NET0131 ,
		_w9436_,
		_w9437_,
		_w12516_,
		_w12517_
	);
	LUT4 #(
		.INIT('hecee)
	) name11168 (
		_w1933_,
		_w12510_,
		_w12511_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h2)
	) name11169 (
		\P2_uWord_reg[4]/NET0131 ,
		_w7767_,
		_w12519_
	);
	LUT3 #(
		.INIT('h80)
	) name11170 (
		\P2_uWord_reg[4]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12520_
	);
	LUT3 #(
		.INIT('h0d)
	) name11171 (
		_w1606_,
		_w2276_,
		_w12520_,
		_w12521_
	);
	LUT2 #(
		.INIT('h2)
	) name11172 (
		_w1565_,
		_w12521_,
		_w12522_
	);
	LUT4 #(
		.INIT('haa02)
	) name11173 (
		\P2_uWord_reg[4]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12523_
	);
	LUT3 #(
		.INIT('h20)
	) name11174 (
		_w1566_,
		_w1602_,
		_w12503_,
		_w12524_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11175 (
		_w1678_,
		_w12523_,
		_w12524_,
		_w12522_,
		_w12525_
	);
	LUT2 #(
		.INIT('he)
	) name11176 (
		_w12519_,
		_w12525_,
		_w12526_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11177 (
		\P1_uWord_reg[4]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w12527_
	);
	LUT3 #(
		.INIT('h20)
	) name11178 (
		_w1797_,
		_w1852_,
		_w12493_,
		_w12528_
	);
	LUT3 #(
		.INIT('h08)
	) name11179 (
		_w1795_,
		_w1867_,
		_w3442_,
		_w12529_
	);
	LUT3 #(
		.INIT('ha8)
	) name11180 (
		_w1933_,
		_w12528_,
		_w12529_,
		_w12530_
	);
	LUT2 #(
		.INIT('he)
	) name11181 (
		_w12527_,
		_w12530_,
		_w12531_
	);
	LUT2 #(
		.INIT('h2)
	) name11182 (
		\P3_EAX_reg[25]/NET0131 ,
		_w8341_,
		_w12532_
	);
	LUT4 #(
		.INIT('h1333)
	) name11183 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		_w8356_,
		_w8358_,
		_w12533_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11184 (
		\P3_EAX_reg[21]/NET0131 ,
		_w8361_,
		_w8356_,
		_w8359_,
		_w12534_
	);
	LUT2 #(
		.INIT('h4)
	) name11185 (
		_w12533_,
		_w12534_,
		_w12535_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11186 (
		\P3_EAX_reg[25]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w12536_
	);
	LUT3 #(
		.INIT('h2d)
	) name11187 (
		_w8391_,
		_w8402_,
		_w8413_,
		_w12537_
	);
	LUT2 #(
		.INIT('h8)
	) name11188 (
		_w8366_,
		_w12537_,
		_w12538_
	);
	LUT3 #(
		.INIT('h80)
	) name11189 (
		\buf2_reg[25]/NET0131 ,
		_w2060_,
		_w2044_,
		_w12539_
	);
	LUT3 #(
		.INIT('h20)
	) name11190 (
		\buf2_reg[9]/NET0131 ,
		_w2060_,
		_w2047_,
		_w12540_
	);
	LUT3 #(
		.INIT('ha8)
	) name11191 (
		_w2119_,
		_w12539_,
		_w12540_,
		_w12541_
	);
	LUT2 #(
		.INIT('h1)
	) name11192 (
		_w12538_,
		_w12541_,
		_w12542_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11193 (
		_w1945_,
		_w12535_,
		_w12536_,
		_w12542_,
		_w12543_
	);
	LUT2 #(
		.INIT('he)
	) name11194 (
		_w12532_,
		_w12543_,
		_w12544_
	);
	LUT2 #(
		.INIT('h2)
	) name11195 (
		\P2_EAX_reg[25]/NET0131 ,
		_w7767_,
		_w12545_
	);
	LUT4 #(
		.INIT('h8000)
	) name11196 (
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[23]/NET0131 ,
		_w7780_,
		_w7781_,
		_w12546_
	);
	LUT4 #(
		.INIT('hb030)
	) name11197 (
		\P2_EAX_reg[24]/NET0131 ,
		_w7789_,
		_w7791_,
		_w12546_,
		_w12547_
	);
	LUT2 #(
		.INIT('h4)
	) name11198 (
		\P2_EAX_reg[25]/NET0131 ,
		_w7789_,
		_w12548_
	);
	LUT3 #(
		.INIT('hd1)
	) name11199 (
		\P2_EAX_reg[25]/NET0131 ,
		_w1606_,
		_w7147_,
		_w12549_
	);
	LUT3 #(
		.INIT('h08)
	) name11200 (
		_w1501_,
		_w1568_,
		_w12549_,
		_w12550_
	);
	LUT4 #(
		.INIT('h08a2)
	) name11201 (
		_w1596_,
		_w7815_,
		_w7826_,
		_w7837_,
		_w12551_
	);
	LUT3 #(
		.INIT('h80)
	) name11202 (
		_w1549_,
		_w1553_,
		_w12551_,
		_w12552_
	);
	LUT3 #(
		.INIT('h1d)
	) name11203 (
		\P2_EAX_reg[25]/NET0131 ,
		_w1606_,
		_w10484_,
		_w12553_
	);
	LUT2 #(
		.INIT('h2)
	) name11204 (
		_w1565_,
		_w12553_,
		_w12554_
	);
	LUT3 #(
		.INIT('h01)
	) name11205 (
		_w12552_,
		_w12554_,
		_w12550_,
		_w12555_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11206 (
		\P2_EAX_reg[24]/NET0131 ,
		_w12546_,
		_w12548_,
		_w12555_,
		_w12556_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11207 (
		\P2_EAX_reg[25]/NET0131 ,
		_w1678_,
		_w12547_,
		_w12556_,
		_w12557_
	);
	LUT2 #(
		.INIT('he)
	) name11208 (
		_w12545_,
		_w12557_,
		_w12558_
	);
	LUT2 #(
		.INIT('h2)
	) name11209 (
		\P3_uWord_reg[4]/NET0131 ,
		_w8341_,
		_w12559_
	);
	LUT4 #(
		.INIT('h55f3)
	) name11210 (
		\P3_uWord_reg[4]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w2105_,
		_w2116_,
		_w12560_
	);
	LUT3 #(
		.INIT('h04)
	) name11211 (
		_w2060_,
		_w2047_,
		_w12560_,
		_w12561_
	);
	LUT3 #(
		.INIT('ha2)
	) name11212 (
		\P3_uWord_reg[4]/NET0131 ,
		_w2047_,
		_w2105_,
		_w12562_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11213 (
		_w1945_,
		_w12499_,
		_w12561_,
		_w12562_,
		_w12563_
	);
	LUT2 #(
		.INIT('he)
	) name11214 (
		_w12559_,
		_w12563_,
		_w12564_
	);
	LUT4 #(
		.INIT('h20aa)
	) name11215 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w12565_
	);
	LUT3 #(
		.INIT('hc8)
	) name11216 (
		\P3_InstQueue_reg[0][7]/NET0131 ,
		_w2215_,
		_w10611_,
		_w12566_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11217 (
		_w1977_,
		_w1982_,
		_w10611_,
		_w12566_,
		_w12567_
	);
	LUT4 #(
		.INIT('h8000)
	) name11218 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10616_,
		_w12568_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11219 (
		\buf2_reg[7]/NET0131 ,
		_w10618_,
		_w10621_,
		_w12568_,
		_w12569_
	);
	LUT3 #(
		.INIT('hef)
	) name11220 (
		_w12567_,
		_w12565_,
		_w12569_,
		_w12570_
	);
	LUT4 #(
		.INIT('h222a)
	) name11221 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w12571_
	);
	LUT3 #(
		.INIT('hc8)
	) name11222 (
		\P3_InstQueue_reg[10][7]/NET0131 ,
		_w2215_,
		_w10630_,
		_w12572_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11223 (
		_w1977_,
		_w1982_,
		_w10630_,
		_w12572_,
		_w12573_
	);
	LUT4 #(
		.INIT('h8000)
	) name11224 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10635_,
		_w12574_
	);
	LUT4 #(
		.INIT('h00df)
	) name11225 (
		\buf2_reg[7]/NET0131 ,
		_w10637_,
		_w10639_,
		_w12574_,
		_w12575_
	);
	LUT3 #(
		.INIT('hef)
	) name11226 (
		_w12573_,
		_w12571_,
		_w12575_,
		_w12576_
	);
	LUT3 #(
		.INIT('hc8)
	) name11227 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		_w2215_,
		_w10646_,
		_w12577_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11228 (
		_w1977_,
		_w1982_,
		_w10646_,
		_w12577_,
		_w12578_
	);
	LUT3 #(
		.INIT('ha2)
	) name11229 (
		\P3_InstQueue_reg[11][7]/NET0131 ,
		_w10622_,
		_w10650_,
		_w12579_
	);
	LUT4 #(
		.INIT('h8000)
	) name11230 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10652_,
		_w12580_
	);
	LUT4 #(
		.INIT('h2000)
	) name11231 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w12581_
	);
	LUT4 #(
		.INIT('hce00)
	) name11232 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w12581_,
		_w12582_
	);
	LUT2 #(
		.INIT('h1)
	) name11233 (
		_w12580_,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h4)
	) name11234 (
		_w12579_,
		_w12583_,
		_w12584_
	);
	LUT2 #(
		.INIT('hb)
	) name11235 (
		_w12578_,
		_w12584_,
		_w12585_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11236 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w12586_
	);
	LUT3 #(
		.INIT('hc8)
	) name11237 (
		\P3_InstQueue_reg[12][7]/NET0131 ,
		_w2215_,
		_w10659_,
		_w12587_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11238 (
		_w1977_,
		_w1982_,
		_w10659_,
		_w12587_,
		_w12588_
	);
	LUT4 #(
		.INIT('h8000)
	) name11239 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10630_,
		_w12589_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11240 (
		\buf2_reg[7]/NET0131 ,
		_w10662_,
		_w10663_,
		_w12589_,
		_w12590_
	);
	LUT3 #(
		.INIT('hef)
	) name11241 (
		_w12588_,
		_w12586_,
		_w12590_,
		_w12591_
	);
	LUT3 #(
		.INIT('hc8)
	) name11242 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w2215_,
		_w10614_,
		_w12592_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11243 (
		_w1977_,
		_w1982_,
		_w10614_,
		_w12592_,
		_w12593_
	);
	LUT2 #(
		.INIT('h4)
	) name11244 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w10672_,
		_w12594_
	);
	LUT2 #(
		.INIT('h1)
	) name11245 (
		\buf2_reg[7]/NET0131 ,
		_w10672_,
		_w12595_
	);
	LUT3 #(
		.INIT('h02)
	) name11246 (
		_w10674_,
		_w12595_,
		_w12594_,
		_w12596_
	);
	LUT4 #(
		.INIT('h8000)
	) name11247 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10646_,
		_w12597_
	);
	LUT2 #(
		.INIT('h2)
	) name11248 (
		\P3_InstQueue_reg[13][7]/NET0131 ,
		_w10622_,
		_w12598_
	);
	LUT2 #(
		.INIT('h1)
	) name11249 (
		_w12597_,
		_w12598_,
		_w12599_
	);
	LUT2 #(
		.INIT('h4)
	) name11250 (
		_w12596_,
		_w12599_,
		_w12600_
	);
	LUT2 #(
		.INIT('hb)
	) name11251 (
		_w12593_,
		_w12600_,
		_w12601_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11252 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w12602_
	);
	LUT3 #(
		.INIT('hc8)
	) name11253 (
		\P3_InstQueue_reg[14][7]/NET0131 ,
		_w2215_,
		_w10616_,
		_w12603_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11254 (
		_w1977_,
		_w1982_,
		_w10616_,
		_w12603_,
		_w12604_
	);
	LUT4 #(
		.INIT('h8000)
	) name11255 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10659_,
		_w12605_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11256 (
		\buf2_reg[7]/NET0131 ,
		_w10617_,
		_w10684_,
		_w12605_,
		_w12606_
	);
	LUT3 #(
		.INIT('hef)
	) name11257 (
		_w12604_,
		_w12602_,
		_w12606_,
		_w12607_
	);
	LUT3 #(
		.INIT('hc8)
	) name11258 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w2215_,
		_w10620_,
		_w12608_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11259 (
		_w1977_,
		_w1982_,
		_w10620_,
		_w12608_,
		_w12609_
	);
	LUT3 #(
		.INIT('hac)
	) name11260 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w10694_,
		_w12610_
	);
	LUT4 #(
		.INIT('h8000)
	) name11261 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10614_,
		_w12611_
	);
	LUT2 #(
		.INIT('h2)
	) name11262 (
		\P3_InstQueue_reg[15][7]/NET0131 ,
		_w10622_,
		_w12612_
	);
	LUT4 #(
		.INIT('h0203)
	) name11263 (
		_w10693_,
		_w12611_,
		_w12612_,
		_w12610_,
		_w12613_
	);
	LUT2 #(
		.INIT('hb)
	) name11264 (
		_w12609_,
		_w12613_,
		_w12614_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11265 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w12615_
	);
	LUT3 #(
		.INIT('hc8)
	) name11266 (
		\P3_InstQueue_reg[1][7]/NET0131 ,
		_w2215_,
		_w10701_,
		_w12616_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11267 (
		_w1977_,
		_w1982_,
		_w10701_,
		_w12616_,
		_w12617_
	);
	LUT4 #(
		.INIT('h8000)
	) name11268 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10620_,
		_w12618_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11269 (
		\buf2_reg[7]/NET0131 ,
		_w10704_,
		_w10705_,
		_w12618_,
		_w12619_
	);
	LUT3 #(
		.INIT('hef)
	) name11270 (
		_w12617_,
		_w12615_,
		_w12619_,
		_w12620_
	);
	LUT4 #(
		.INIT('h222a)
	) name11271 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w12621_
	);
	LUT3 #(
		.INIT('hc8)
	) name11272 (
		\P3_InstQueue_reg[2][7]/NET0131 ,
		_w2215_,
		_w10713_,
		_w12622_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11273 (
		_w1977_,
		_w1982_,
		_w10713_,
		_w12622_,
		_w12623_
	);
	LUT4 #(
		.INIT('h8000)
	) name11274 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10611_,
		_w12624_
	);
	LUT4 #(
		.INIT('h00df)
	) name11275 (
		\buf2_reg[7]/NET0131 ,
		_w10716_,
		_w10717_,
		_w12624_,
		_w12625_
	);
	LUT3 #(
		.INIT('hef)
	) name11276 (
		_w12623_,
		_w12621_,
		_w12625_,
		_w12626_
	);
	LUT4 #(
		.INIT('h222a)
	) name11277 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w12627_
	);
	LUT3 #(
		.INIT('hc8)
	) name11278 (
		\P3_InstQueue_reg[3][7]/NET0131 ,
		_w2215_,
		_w10724_,
		_w12628_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11279 (
		_w1977_,
		_w1982_,
		_w10724_,
		_w12628_,
		_w12629_
	);
	LUT4 #(
		.INIT('h8000)
	) name11280 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10701_,
		_w12630_
	);
	LUT4 #(
		.INIT('h00f7)
	) name11281 (
		\buf2_reg[7]/NET0131 ,
		_w10712_,
		_w10727_,
		_w12630_,
		_w12631_
	);
	LUT3 #(
		.INIT('hef)
	) name11282 (
		_w12629_,
		_w12627_,
		_w12631_,
		_w12632_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11283 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w12633_
	);
	LUT3 #(
		.INIT('hc8)
	) name11284 (
		\P3_InstQueue_reg[4][7]/NET0131 ,
		_w2215_,
		_w10734_,
		_w12634_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11285 (
		_w1977_,
		_w1982_,
		_w10734_,
		_w12634_,
		_w12635_
	);
	LUT4 #(
		.INIT('h8000)
	) name11286 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10713_,
		_w12636_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11287 (
		\buf2_reg[7]/NET0131 ,
		_w10737_,
		_w10738_,
		_w12636_,
		_w12637_
	);
	LUT3 #(
		.INIT('hef)
	) name11288 (
		_w12635_,
		_w12633_,
		_w12637_,
		_w12638_
	);
	LUT3 #(
		.INIT('hc8)
	) name11289 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w2215_,
		_w10745_,
		_w12639_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11290 (
		_w1977_,
		_w1982_,
		_w10745_,
		_w12639_,
		_w12640_
	);
	LUT2 #(
		.INIT('h4)
	) name11291 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w10748_,
		_w12641_
	);
	LUT2 #(
		.INIT('h1)
	) name11292 (
		\buf2_reg[7]/NET0131 ,
		_w10748_,
		_w12642_
	);
	LUT3 #(
		.INIT('h02)
	) name11293 (
		_w10750_,
		_w12642_,
		_w12641_,
		_w12643_
	);
	LUT4 #(
		.INIT('h8000)
	) name11294 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10724_,
		_w12644_
	);
	LUT2 #(
		.INIT('h2)
	) name11295 (
		\P3_InstQueue_reg[5][7]/NET0131 ,
		_w10622_,
		_w12645_
	);
	LUT2 #(
		.INIT('h1)
	) name11296 (
		_w12644_,
		_w12645_,
		_w12646_
	);
	LUT2 #(
		.INIT('h4)
	) name11297 (
		_w12643_,
		_w12646_,
		_w12647_
	);
	LUT2 #(
		.INIT('hb)
	) name11298 (
		_w12640_,
		_w12647_,
		_w12648_
	);
	LUT4 #(
		.INIT('h2a22)
	) name11299 (
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w12649_
	);
	LUT3 #(
		.INIT('hc8)
	) name11300 (
		\P3_InstQueue_reg[6][7]/NET0131 ,
		_w2215_,
		_w10758_,
		_w12650_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11301 (
		_w1977_,
		_w1982_,
		_w10758_,
		_w12650_,
		_w12651_
	);
	LUT4 #(
		.INIT('h8000)
	) name11302 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10734_,
		_w12652_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11303 (
		\buf2_reg[7]/NET0131 ,
		_w10761_,
		_w10762_,
		_w12652_,
		_w12653_
	);
	LUT3 #(
		.INIT('hef)
	) name11304 (
		_w12651_,
		_w12649_,
		_w12653_,
		_w12654_
	);
	LUT3 #(
		.INIT('hc8)
	) name11305 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w2215_,
		_w10633_,
		_w12655_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11306 (
		_w1977_,
		_w1982_,
		_w10633_,
		_w12655_,
		_w12656_
	);
	LUT3 #(
		.INIT('hac)
	) name11307 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w10772_,
		_w12657_
	);
	LUT4 #(
		.INIT('h8000)
	) name11308 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10745_,
		_w12658_
	);
	LUT2 #(
		.INIT('h2)
	) name11309 (
		\P3_InstQueue_reg[7][7]/NET0131 ,
		_w10622_,
		_w12659_
	);
	LUT4 #(
		.INIT('h0203)
	) name11310 (
		_w10771_,
		_w12658_,
		_w12659_,
		_w12657_,
		_w12660_
	);
	LUT2 #(
		.INIT('hb)
	) name11311 (
		_w12656_,
		_w12660_,
		_w12661_
	);
	LUT4 #(
		.INIT('h22a2)
	) name11312 (
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w12662_
	);
	LUT3 #(
		.INIT('hc8)
	) name11313 (
		\P3_InstQueue_reg[8][7]/NET0131 ,
		_w2215_,
		_w10635_,
		_w12663_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11314 (
		_w1977_,
		_w1982_,
		_w10635_,
		_w12663_,
		_w12664_
	);
	LUT4 #(
		.INIT('h8000)
	) name11315 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10758_,
		_w12665_
	);
	LUT4 #(
		.INIT('h00fd)
	) name11316 (
		\buf2_reg[7]/NET0131 ,
		_w10636_,
		_w10781_,
		_w12665_,
		_w12666_
	);
	LUT3 #(
		.INIT('hef)
	) name11317 (
		_w12664_,
		_w12662_,
		_w12666_,
		_w12667_
	);
	LUT3 #(
		.INIT('hc8)
	) name11318 (
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w2215_,
		_w10652_,
		_w12668_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11319 (
		_w1977_,
		_w1982_,
		_w10652_,
		_w12668_,
		_w12669_
	);
	LUT3 #(
		.INIT('h02)
	) name11320 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w3055_,
		_w10772_,
		_w12670_
	);
	LUT4 #(
		.INIT('h1000)
	) name11321 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w12671_
	);
	LUT4 #(
		.INIT('hef00)
	) name11322 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w12672_
	);
	LUT3 #(
		.INIT('h54)
	) name11323 (
		_w6349_,
		_w12671_,
		_w12672_,
		_w12673_
	);
	LUT4 #(
		.INIT('h8000)
	) name11324 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2194_,
		_w10633_,
		_w12674_
	);
	LUT2 #(
		.INIT('h2)
	) name11325 (
		\P3_InstQueue_reg[9][7]/NET0131 ,
		_w10622_,
		_w12675_
	);
	LUT4 #(
		.INIT('h1011)
	) name11326 (
		_w12674_,
		_w12675_,
		_w12670_,
		_w12673_,
		_w12676_
	);
	LUT2 #(
		.INIT('hb)
	) name11327 (
		_w12669_,
		_w12676_,
		_w12677_
	);
	LUT4 #(
		.INIT('h550d)
	) name11328 (
		\P3_MemoryFetch_reg/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12678_
	);
	LUT4 #(
		.INIT('hfc23)
	) name11329 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w12679_
	);
	LUT3 #(
		.INIT('hc4)
	) name11330 (
		\P3_MemoryFetch_reg/NET0131 ,
		_w9129_,
		_w12679_,
		_w12680_
	);
	LUT3 #(
		.INIT('h2f)
	) name11331 (
		_w1945_,
		_w12678_,
		_w12680_,
		_w12681_
	);
	LUT3 #(
		.INIT('ha2)
	) name11332 (
		\P1_MemoryFetch_reg/NET0131 ,
		_w1802_,
		_w1852_,
		_w12682_
	);
	LUT3 #(
		.INIT('hc4)
	) name11333 (
		\P1_MemoryFetch_reg/NET0131 ,
		_w8459_,
		_w9470_,
		_w12683_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name11334 (
		_w1933_,
		_w9472_,
		_w12682_,
		_w12683_,
		_w12684_
	);
	LUT3 #(
		.INIT('ha2)
	) name11335 (
		\P2_MemoryFetch_reg/NET0131 ,
		_w1568_,
		_w1602_,
		_w12685_
	);
	LUT4 #(
		.INIT('hfc23)
	) name11336 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w12686_
	);
	LUT3 #(
		.INIT('hc4)
	) name11337 (
		\P2_MemoryFetch_reg/NET0131 ,
		_w2287_,
		_w12686_,
		_w12687_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name11338 (
		_w1678_,
		_w9466_,
		_w12685_,
		_w12687_,
		_w12688_
	);
	LUT4 #(
		.INIT('h08aa)
	) name11339 (
		\P2_rEIP_reg[0]/NET0131 ,
		_w1673_,
		_w9786_,
		_w9788_,
		_w12689_
	);
	LUT3 #(
		.INIT('h04)
	) name11340 (
		\P2_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1568_,
		_w1602_,
		_w12690_
	);
	LUT4 #(
		.INIT('h0057)
	) name11341 (
		\P2_EBX_reg[0]/NET0131 ,
		_w9752_,
		_w9765_,
		_w12690_,
		_w12691_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11342 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		_w1679_,
		_w2211_,
		_w12692_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11343 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w1679_,
		_w9799_,
		_w12693_
	);
	LUT2 #(
		.INIT('h1)
	) name11344 (
		_w12692_,
		_w12693_,
		_w12694_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11345 (
		_w1678_,
		_w12689_,
		_w12691_,
		_w12694_,
		_w12695_
	);
	LUT3 #(
		.INIT('h8c)
	) name11346 (
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w11331_,
		_w12696_
	);
	LUT4 #(
		.INIT('h70b0)
	) name11347 (
		\P1_rEIP_reg[30]/NET0131 ,
		_w1930_,
		_w4709_,
		_w11333_,
		_w12697_
	);
	LUT4 #(
		.INIT('hde00)
	) name11348 (
		\P1_EBX_reg[30]/NET0131 ,
		_w1930_,
		_w12696_,
		_w12697_,
		_w12698_
	);
	LUT2 #(
		.INIT('h2)
	) name11349 (
		\P1_rEIP_reg[30]/NET0131 ,
		_w10808_,
		_w12699_
	);
	LUT4 #(
		.INIT('h3332)
	) name11350 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12700_
	);
	LUT3 #(
		.INIT('h02)
	) name11351 (
		_w1797_,
		_w1852_,
		_w12700_,
		_w12701_
	);
	LUT4 #(
		.INIT('h7b00)
	) name11352 (
		\P1_rEIP_reg[30]/NET0131 ,
		_w10817_,
		_w11333_,
		_w12701_,
		_w12702_
	);
	LUT2 #(
		.INIT('h1)
	) name11353 (
		_w12699_,
		_w12702_,
		_w12703_
	);
	LUT3 #(
		.INIT('h8a)
	) name11354 (
		_w1933_,
		_w12698_,
		_w12703_,
		_w12704_
	);
	LUT3 #(
		.INIT('h80)
	) name11355 (
		\P1_PhyAddrPointer_reg[28]/NET0131 ,
		\P1_PhyAddrPointer_reg[29]/NET0131 ,
		_w11277_,
		_w12705_
	);
	LUT4 #(
		.INIT('h1141)
	) name11356 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6377_,
		_w10800_,
		_w12705_,
		_w12706_
	);
	LUT2 #(
		.INIT('h2)
	) name11357 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w12707_
	);
	LUT2 #(
		.INIT('h2)
	) name11358 (
		_w1939_,
		_w12707_,
		_w12708_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11359 (
		\P1_PhyAddrPointer_reg[30]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w2234_,
		_w10828_,
		_w12709_
	);
	LUT3 #(
		.INIT('hb0)
	) name11360 (
		_w12706_,
		_w12708_,
		_w12709_,
		_w12710_
	);
	LUT2 #(
		.INIT('hb)
	) name11361 (
		_w12704_,
		_w12710_,
		_w12711_
	);
	LUT4 #(
		.INIT('h60c0)
	) name11362 (
		\P1_rEIP_reg[30]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w1930_,
		_w11333_,
		_w12712_
	);
	LUT2 #(
		.INIT('h4)
	) name11363 (
		\P1_EBX_reg[30]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w12713_
	);
	LUT2 #(
		.INIT('h8)
	) name11364 (
		_w11337_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h8)
	) name11365 (
		_w11331_,
		_w12714_,
		_w12715_
	);
	LUT3 #(
		.INIT('ha8)
	) name11366 (
		_w4709_,
		_w12712_,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h2)
	) name11367 (
		\P1_rEIP_reg[31]/NET0131 ,
		_w10808_,
		_w12717_
	);
	LUT4 #(
		.INIT('h9030)
	) name11368 (
		\P1_rEIP_reg[30]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w10817_,
		_w11333_,
		_w12718_
	);
	LUT4 #(
		.INIT('h3332)
	) name11369 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[31]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12719_
	);
	LUT3 #(
		.INIT('h02)
	) name11370 (
		_w1797_,
		_w1852_,
		_w12719_,
		_w12720_
	);
	LUT3 #(
		.INIT('h45)
	) name11371 (
		_w12717_,
		_w12718_,
		_w12720_,
		_w12721_
	);
	LUT3 #(
		.INIT('h8a)
	) name11372 (
		_w1933_,
		_w12716_,
		_w12721_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name11373 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w12723_
	);
	LUT2 #(
		.INIT('h1)
	) name11374 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w6377_,
		_w12724_
	);
	LUT4 #(
		.INIT('h070f)
	) name11375 (
		_w10800_,
		_w12705_,
		_w12723_,
		_w12724_,
		_w12725_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11376 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w2234_,
		_w10828_,
		_w12726_
	);
	LUT3 #(
		.INIT('hd0)
	) name11377 (
		_w1939_,
		_w12725_,
		_w12726_,
		_w12727_
	);
	LUT2 #(
		.INIT('hb)
	) name11378 (
		_w12722_,
		_w12727_,
		_w12728_
	);
	LUT2 #(
		.INIT('h8)
	) name11379 (
		_w6364_,
		_w10801_,
		_w12729_
	);
	LUT3 #(
		.INIT('h06)
	) name11380 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w12729_,
		_w12730_
	);
	LUT2 #(
		.INIT('h2)
	) name11381 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w12731_
	);
	LUT2 #(
		.INIT('h2)
	) name11382 (
		_w1939_,
		_w12731_,
		_w12732_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11383 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w9636_,
		_w12730_,
		_w12732_,
		_w12733_
	);
	LUT3 #(
		.INIT('h84)
	) name11384 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w1930_,
		_w10810_,
		_w12734_
	);
	LUT4 #(
		.INIT('h2010)
	) name11385 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w1858_,
		_w1930_,
		_w10810_,
		_w12735_
	);
	LUT4 #(
		.INIT('h3332)
	) name11386 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12736_
	);
	LUT2 #(
		.INIT('h1)
	) name11387 (
		_w12735_,
		_w12736_,
		_w12737_
	);
	LUT3 #(
		.INIT('h20)
	) name11388 (
		_w1797_,
		_w1852_,
		_w12737_,
		_w12738_
	);
	LUT3 #(
		.INIT('h8a)
	) name11389 (
		\P1_EBX_reg[31]/NET0131 ,
		\P1_EBX_reg[4]/NET0131 ,
		_w10820_,
		_w12739_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name11390 (
		\P1_EBX_reg[5]/NET0131 ,
		_w1930_,
		_w12734_,
		_w12739_,
		_w12740_
	);
	LUT3 #(
		.INIT('h20)
	) name11391 (
		_w1795_,
		_w1852_,
		_w12740_,
		_w12741_
	);
	LUT4 #(
		.INIT('h000d)
	) name11392 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w10808_,
		_w12738_,
		_w12741_,
		_w12742_
	);
	LUT2 #(
		.INIT('h2)
	) name11393 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w10828_,
		_w12743_
	);
	LUT3 #(
		.INIT('h07)
	) name11394 (
		\P1_PhyAddrPointer_reg[5]/NET0131 ,
		_w2234_,
		_w3406_,
		_w12744_
	);
	LUT2 #(
		.INIT('h4)
	) name11395 (
		_w12743_,
		_w12744_,
		_w12745_
	);
	LUT3 #(
		.INIT('hd0)
	) name11396 (
		_w1933_,
		_w12742_,
		_w12745_,
		_w12746_
	);
	LUT2 #(
		.INIT('hb)
	) name11397 (
		_w12733_,
		_w12746_,
		_w12747_
	);
	LUT3 #(
		.INIT('h8c)
	) name11398 (
		\P2_EBX_reg[29]/NET0131 ,
		\P2_EBX_reg[31]/NET0131 ,
		_w9764_,
		_w12748_
	);
	LUT4 #(
		.INIT('h9030)
	) name11399 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w1673_,
		_w9784_,
		_w12749_
	);
	LUT2 #(
		.INIT('h2)
	) name11400 (
		_w6439_,
		_w12749_,
		_w12750_
	);
	LUT4 #(
		.INIT('hde00)
	) name11401 (
		\P2_EBX_reg[30]/NET0131 ,
		_w1673_,
		_w12748_,
		_w12750_,
		_w12751_
	);
	LUT2 #(
		.INIT('h2)
	) name11402 (
		\P2_rEIP_reg[30]/NET0131 ,
		_w9788_,
		_w12752_
	);
	LUT4 #(
		.INIT('h9300)
	) name11403 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9784_,
		_w9751_,
		_w12753_
	);
	LUT4 #(
		.INIT('h3332)
	) name11404 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_EBX_reg[30]/NET0131 ,
		_w1605_,
		_w1611_,
		_w12754_
	);
	LUT3 #(
		.INIT('h02)
	) name11405 (
		_w1566_,
		_w1602_,
		_w12754_,
		_w12755_
	);
	LUT3 #(
		.INIT('h45)
	) name11406 (
		_w12752_,
		_w12753_,
		_w12755_,
		_w12756_
	);
	LUT3 #(
		.INIT('h8a)
	) name11407 (
		_w1678_,
		_w12751_,
		_w12756_,
		_w12757_
	);
	LUT4 #(
		.INIT('h0c6c)
	) name11408 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5744_,
		_w9796_,
		_w12758_
	);
	LUT2 #(
		.INIT('h2)
	) name11409 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w12759_
	);
	LUT2 #(
		.INIT('h2)
	) name11410 (
		_w1679_,
		_w12759_,
		_w12760_
	);
	LUT4 #(
		.INIT('hbe00)
	) name11411 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w6327_,
		_w12758_,
		_w12760_,
		_w12761_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11412 (
		\P2_PhyAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2211_,
		_w9799_,
		_w12762_
	);
	LUT2 #(
		.INIT('h4)
	) name11413 (
		_w12761_,
		_w12762_,
		_w12763_
	);
	LUT2 #(
		.INIT('hb)
	) name11414 (
		_w12757_,
		_w12763_,
		_w12764_
	);
	LUT4 #(
		.INIT('heda5)
	) name11415 (
		\P2_PhyAddrPointer_reg[31]/NET0131 ,
		_w5722_,
		_w5745_,
		_w9792_,
		_w12765_
	);
	LUT2 #(
		.INIT('h2)
	) name11416 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w12766_
	);
	LUT2 #(
		.INIT('h2)
	) name11417 (
		_w1679_,
		_w12766_,
		_w12767_
	);
	LUT4 #(
		.INIT('heb00)
	) name11418 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w9564_,
		_w12765_,
		_w12767_,
		_w12768_
	);
	LUT3 #(
		.INIT('h8a)
	) name11419 (
		\P2_EBX_reg[31]/NET0131 ,
		\P2_EBX_reg[4]/NET0131 ,
		_w9753_,
		_w12769_
	);
	LUT2 #(
		.INIT('h6)
	) name11420 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w9768_,
		_w12770_
	);
	LUT3 #(
		.INIT('h84)
	) name11421 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w1673_,
		_w9768_,
		_w12771_
	);
	LUT4 #(
		.INIT('h00de)
	) name11422 (
		\P2_EBX_reg[5]/NET0131 ,
		_w1673_,
		_w12769_,
		_w12771_,
		_w12772_
	);
	LUT3 #(
		.INIT('h20)
	) name11423 (
		_w1565_,
		_w1602_,
		_w12772_,
		_w12773_
	);
	LUT3 #(
		.INIT('he2)
	) name11424 (
		\P2_EBX_reg[5]/NET0131 ,
		_w9751_,
		_w12770_,
		_w12774_
	);
	LUT3 #(
		.INIT('h20)
	) name11425 (
		_w1566_,
		_w1602_,
		_w12774_,
		_w12775_
	);
	LUT4 #(
		.INIT('h000d)
	) name11426 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w9788_,
		_w12773_,
		_w12775_,
		_w12776_
	);
	LUT2 #(
		.INIT('h2)
	) name11427 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w9799_,
		_w12777_
	);
	LUT3 #(
		.INIT('h07)
	) name11428 (
		\P2_PhyAddrPointer_reg[5]/NET0131 ,
		_w2211_,
		_w2286_,
		_w12778_
	);
	LUT2 #(
		.INIT('h4)
	) name11429 (
		_w12777_,
		_w12778_,
		_w12779_
	);
	LUT3 #(
		.INIT('hd0)
	) name11430 (
		_w1678_,
		_w12776_,
		_w12779_,
		_w12780_
	);
	LUT2 #(
		.INIT('hb)
	) name11431 (
		_w12768_,
		_w12780_,
		_w12781_
	);
	LUT4 #(
		.INIT('h4c00)
	) name11432 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w2187_,
		_w12782_
	);
	LUT3 #(
		.INIT('ha8)
	) name11433 (
		\P3_rEIP_reg[0]/NET0131 ,
		_w2178_,
		_w12782_,
		_w12783_
	);
	LUT2 #(
		.INIT('h4)
	) name11434 (
		\P3_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2044_,
		_w12784_
	);
	LUT4 #(
		.INIT('h7f33)
	) name11435 (
		_w2060_,
		_w2047_,
		_w2111_,
		_w2187_,
		_w12785_
	);
	LUT4 #(
		.INIT('h3032)
	) name11436 (
		\P3_EBX_reg[0]/NET0131 ,
		_w2105_,
		_w12784_,
		_w12785_,
		_w12786_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11437 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w2194_,
		_w2225_,
		_w12787_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11438 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w2194_,
		_w11818_,
		_w12788_
	);
	LUT2 #(
		.INIT('h1)
	) name11439 (
		_w12787_,
		_w12788_,
		_w12789_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11440 (
		_w1945_,
		_w12783_,
		_w12786_,
		_w12789_,
		_w12790_
	);
	LUT2 #(
		.INIT('h4)
	) name11441 (
		_w5779_,
		_w6985_,
		_w12791_
	);
	LUT4 #(
		.INIT('h4441)
	) name11442 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w6348_,
		_w12206_,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h2)
	) name11443 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w12793_
	);
	LUT2 #(
		.INIT('h2)
	) name11444 (
		_w2194_,
		_w12793_,
		_w12794_
	);
	LUT4 #(
		.INIT('h0001)
	) name11445 (
		\P3_EBX_reg[26]/NET0131 ,
		\P3_EBX_reg[27]/NET0131 ,
		\P3_EBX_reg[28]/NET0131 ,
		\P3_EBX_reg[29]/NET0131 ,
		_w12795_
	);
	LUT4 #(
		.INIT('h4000)
	) name11446 (
		\P3_EBX_reg[25]/NET0131 ,
		_w12067_,
		_w12128_,
		_w12795_,
		_w12796_
	);
	LUT4 #(
		.INIT('h0509)
	) name11447 (
		\P3_EBX_reg[30]/NET0131 ,
		\P3_EBX_reg[31]/NET0131 ,
		_w2187_,
		_w12796_,
		_w12797_
	);
	LUT4 #(
		.INIT('h8444)
	) name11448 (
		\P3_rEIP_reg[30]/NET0131 ,
		_w2187_,
		_w12120_,
		_w12193_,
		_w12798_
	);
	LUT2 #(
		.INIT('h2)
	) name11449 (
		_w11831_,
		_w12798_,
		_w12799_
	);
	LUT4 #(
		.INIT('haa02)
	) name11450 (
		\P3_rEIP_reg[30]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12800_
	);
	LUT3 #(
		.INIT('h45)
	) name11451 (
		\P3_EBX_reg[30]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12801_
	);
	LUT4 #(
		.INIT('h0008)
	) name11452 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12801_,
		_w12802_
	);
	LUT4 #(
		.INIT('h040f)
	) name11453 (
		_w2111_,
		_w12798_,
		_w12800_,
		_w12802_,
		_w12803_
	);
	LUT4 #(
		.INIT('h20aa)
	) name11454 (
		_w1945_,
		_w12797_,
		_w12799_,
		_w12803_,
		_w12804_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11455 (
		\P3_PhyAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2225_,
		_w11818_,
		_w12805_
	);
	LUT2 #(
		.INIT('h4)
	) name11456 (
		_w12804_,
		_w12805_,
		_w12806_
	);
	LUT3 #(
		.INIT('h4f)
	) name11457 (
		_w12792_,
		_w12794_,
		_w12806_,
		_w12807_
	);
	LUT3 #(
		.INIT('hec)
	) name11458 (
		_w5757_,
		_w5779_,
		_w12212_,
		_w12808_
	);
	LUT2 #(
		.INIT('h2)
	) name11459 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w12809_
	);
	LUT2 #(
		.INIT('h2)
	) name11460 (
		_w2194_,
		_w12809_,
		_w12810_
	);
	LUT4 #(
		.INIT('heb00)
	) name11461 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w9600_,
		_w12808_,
		_w12810_,
		_w12811_
	);
	LUT4 #(
		.INIT('h2010)
	) name11462 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2111_,
		_w2187_,
		_w11803_,
		_w12812_
	);
	LUT3 #(
		.INIT('h45)
	) name11463 (
		\P3_EBX_reg[5]/NET0131 ,
		_w2111_,
		_w2187_,
		_w12813_
	);
	LUT2 #(
		.INIT('h1)
	) name11464 (
		_w12812_,
		_w12813_,
		_w12814_
	);
	LUT4 #(
		.INIT('h0800)
	) name11465 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12814_,
		_w12815_
	);
	LUT4 #(
		.INIT('haa02)
	) name11466 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2044_,
		_w2047_,
		_w2105_,
		_w12816_
	);
	LUT3 #(
		.INIT('h84)
	) name11467 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2187_,
		_w11803_,
		_w12817_
	);
	LUT3 #(
		.INIT('h8a)
	) name11468 (
		\P3_EBX_reg[31]/NET0131 ,
		\P3_EBX_reg[4]/NET0131 ,
		_w11811_,
		_w12818_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name11469 (
		\P3_EBX_reg[5]/NET0131 ,
		_w2187_,
		_w12817_,
		_w12818_,
		_w12819_
	);
	LUT4 #(
		.INIT('h0400)
	) name11470 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w12819_,
		_w12820_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11471 (
		_w1945_,
		_w12816_,
		_w12820_,
		_w12815_,
		_w12821_
	);
	LUT2 #(
		.INIT('h2)
	) name11472 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w11818_,
		_w12822_
	);
	LUT3 #(
		.INIT('h07)
	) name11473 (
		\P3_PhyAddrPointer_reg[5]/NET0131 ,
		_w2225_,
		_w3054_,
		_w12823_
	);
	LUT2 #(
		.INIT('h4)
	) name11474 (
		_w12822_,
		_w12823_,
		_w12824_
	);
	LUT2 #(
		.INIT('h4)
	) name11475 (
		_w12821_,
		_w12824_,
		_w12825_
	);
	LUT2 #(
		.INIT('hb)
	) name11476 (
		_w12811_,
		_w12825_,
		_w12826_
	);
	LUT2 #(
		.INIT('h8)
	) name11477 (
		_w1797_,
		_w10817_,
		_w12827_
	);
	LUT3 #(
		.INIT('ha2)
	) name11478 (
		\P1_rEIP_reg[0]/NET0131 ,
		_w10808_,
		_w12827_,
		_w12828_
	);
	LUT4 #(
		.INIT('h0444)
	) name11479 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w12829_
	);
	LUT4 #(
		.INIT('hc888)
	) name11480 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w12830_
	);
	LUT4 #(
		.INIT('h020f)
	) name11481 (
		_w1842_,
		_w1851_,
		_w12829_,
		_w12830_,
		_w12831_
	);
	LUT2 #(
		.INIT('h2)
	) name11482 (
		_w1795_,
		_w12831_,
		_w12832_
	);
	LUT4 #(
		.INIT('hccc8)
	) name11483 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_EBX_reg[0]/NET0131 ,
		_w1858_,
		_w1861_,
		_w12833_
	);
	LUT4 #(
		.INIT('h23af)
	) name11484 (
		\P1_InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1797_,
		_w1802_,
		_w12833_,
		_w12834_
	);
	LUT3 #(
		.INIT('h32)
	) name11485 (
		_w1852_,
		_w12832_,
		_w12834_,
		_w12835_
	);
	LUT4 #(
		.INIT('hcc40)
	) name11486 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		_w1939_,
		_w2234_,
		_w12836_
	);
	LUT4 #(
		.INIT('h80cc)
	) name11487 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w1939_,
		_w10828_,
		_w12837_
	);
	LUT2 #(
		.INIT('h1)
	) name11488 (
		_w12836_,
		_w12837_,
		_w12838_
	);
	LUT4 #(
		.INIT('h8aff)
	) name11489 (
		_w1933_,
		_w12828_,
		_w12835_,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h2)
	) name11490 (
		\datao[27]_pad ,
		_w2115_,
		_w12840_
	);
	LUT3 #(
		.INIT('h13)
	) name11491 (
		\P3_EAX_reg[26]/NET0131 ,
		\P3_EAX_reg[27]/NET0131 ,
		_w9541_,
		_w12841_
	);
	LUT4 #(
		.INIT('h0004)
	) name11492 (
		_w2111_,
		_w9543_,
		_w9542_,
		_w12841_,
		_w12842_
	);
	LUT4 #(
		.INIT('h5f13)
	) name11493 (
		\P3_uWord_reg[11]/NET0131 ,
		\datao[27]_pad ,
		_w9977_,
		_w9978_,
		_w12843_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11494 (
		_w1945_,
		_w12840_,
		_w12842_,
		_w12843_,
		_w12844_
	);
	LUT2 #(
		.INIT('h2)
	) name11495 (
		\P1_Datao_reg[27]/NET0131 ,
		_w1860_,
		_w12845_
	);
	LUT4 #(
		.INIT('h8000)
	) name11496 (
		\P1_EAX_reg[22]/NET0131 ,
		\P1_EAX_reg[25]/NET0131 ,
		_w9433_,
		_w9484_,
		_w12846_
	);
	LUT3 #(
		.INIT('h13)
	) name11497 (
		\P1_EAX_reg[26]/NET0131 ,
		\P1_EAX_reg[27]/NET0131 ,
		_w12846_,
		_w12847_
	);
	LUT2 #(
		.INIT('h2)
	) name11498 (
		_w1797_,
		_w9487_,
		_w12848_
	);
	LUT3 #(
		.INIT('h20)
	) name11499 (
		_w1859_,
		_w12847_,
		_w12848_,
		_w12849_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11500 (
		\P1_Datao_reg[27]/NET0131 ,
		\P1_uWord_reg[11]/NET0131 ,
		_w1935_,
		_w9972_,
		_w12850_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11501 (
		_w1933_,
		_w12845_,
		_w12849_,
		_w12850_,
		_w12851_
	);
	LUT4 #(
		.INIT('h0903)
	) name11502 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		_w1611_,
		_w9460_,
		_w12852_
	);
	LUT4 #(
		.INIT('h5445)
	) name11503 (
		\P2_Datao_reg[27]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w12853_
	);
	LUT3 #(
		.INIT('h02)
	) name11504 (
		_w1566_,
		_w1602_,
		_w12853_,
		_w12854_
	);
	LUT2 #(
		.INIT('h4)
	) name11505 (
		_w12852_,
		_w12854_,
		_w12855_
	);
	LUT3 #(
		.INIT('ha2)
	) name11506 (
		\P2_Datao_reg[27]/NET0131 ,
		_w4927_,
		_w9989_,
		_w12856_
	);
	LUT4 #(
		.INIT('h3f15)
	) name11507 (
		\P2_Datao_reg[27]/NET0131 ,
		\P2_uWord_reg[11]/NET0131 ,
		_w9995_,
		_w9996_,
		_w12857_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name11508 (
		_w1678_,
		_w12855_,
		_w12856_,
		_w12857_,
		_w12858_
	);
	LUT2 #(
		.INIT('h2)
	) name11509 (
		\P1_EAX_reg[23]/NET0131 ,
		_w9102_,
		_w12859_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name11510 (
		\P1_EAX_reg[23]/NET0131 ,
		_w1827_,
		_w9430_,
		_w9432_,
		_w12860_
	);
	LUT4 #(
		.INIT('h4888)
	) name11511 (
		\P1_EAX_reg[23]/NET0131 ,
		_w1827_,
		_w9430_,
		_w9432_,
		_w12861_
	);
	LUT4 #(
		.INIT('h0080)
	) name11512 (
		_w1725_,
		_w1802_,
		_w1867_,
		_w3507_,
		_w12862_
	);
	LUT4 #(
		.INIT('h7888)
	) name11513 (
		_w8999_,
		_w9004_,
		_w9009_,
		_w9014_,
		_w12863_
	);
	LUT2 #(
		.INIT('h8)
	) name11514 (
		_w1846_,
		_w12863_,
		_w12864_
	);
	LUT4 #(
		.INIT('h4000)
	) name11515 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w12864_,
		_w12865_
	);
	LUT3 #(
		.INIT('h08)
	) name11516 (
		_w1795_,
		_w1867_,
		_w3438_,
		_w12866_
	);
	LUT3 #(
		.INIT('h01)
	) name11517 (
		_w12865_,
		_w12866_,
		_w12862_,
		_w12867_
	);
	LUT4 #(
		.INIT('h7500)
	) name11518 (
		\P1_EAX_reg[23]/NET0131 ,
		_w9436_,
		_w9437_,
		_w12867_,
		_w12868_
	);
	LUT4 #(
		.INIT('hecee)
	) name11519 (
		_w1933_,
		_w12859_,
		_w12861_,
		_w12868_,
		_w12869_
	);
	LUT3 #(
		.INIT('h80)
	) name11520 (
		\P2_lWord_reg[0]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12870_
	);
	LUT3 #(
		.INIT('h0d)
	) name11521 (
		_w1606_,
		_w9115_,
		_w12870_,
		_w12871_
	);
	LUT2 #(
		.INIT('h2)
	) name11522 (
		_w1565_,
		_w12871_,
		_w12872_
	);
	LUT4 #(
		.INIT('haa02)
	) name11523 (
		\P2_lWord_reg[0]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12873_
	);
	LUT3 #(
		.INIT('h08)
	) name11524 (
		\P2_EAX_reg[0]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12874_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11525 (
		_w1678_,
		_w12873_,
		_w12872_,
		_w12874_,
		_w12875_
	);
	LUT2 #(
		.INIT('h2)
	) name11526 (
		\P2_lWord_reg[0]/NET0131 ,
		_w7767_,
		_w12876_
	);
	LUT2 #(
		.INIT('he)
	) name11527 (
		_w12875_,
		_w12876_,
		_w12877_
	);
	LUT2 #(
		.INIT('h2)
	) name11528 (
		\P2_lWord_reg[10]/NET0131 ,
		_w7767_,
		_w12878_
	);
	LUT3 #(
		.INIT('h80)
	) name11529 (
		\P2_lWord_reg[10]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12879_
	);
	LUT3 #(
		.INIT('h0b)
	) name11530 (
		_w1602_,
		_w9522_,
		_w12879_,
		_w12880_
	);
	LUT2 #(
		.INIT('h2)
	) name11531 (
		_w1565_,
		_w12880_,
		_w12881_
	);
	LUT3 #(
		.INIT('h08)
	) name11532 (
		\P2_EAX_reg[10]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12882_
	);
	LUT4 #(
		.INIT('haa02)
	) name11533 (
		\P2_lWord_reg[10]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12883_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11534 (
		_w1678_,
		_w12882_,
		_w12883_,
		_w12881_,
		_w12884_
	);
	LUT2 #(
		.INIT('he)
	) name11535 (
		_w12878_,
		_w12884_,
		_w12885_
	);
	LUT2 #(
		.INIT('h2)
	) name11536 (
		\P2_lWord_reg[11]/NET0131 ,
		_w7767_,
		_w12886_
	);
	LUT3 #(
		.INIT('h80)
	) name11537 (
		\P2_lWord_reg[11]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12887_
	);
	LUT3 #(
		.INIT('h54)
	) name11538 (
		_w1605_,
		_w8450_,
		_w8451_,
		_w12888_
	);
	LUT3 #(
		.INIT('h23)
	) name11539 (
		_w1602_,
		_w12887_,
		_w12888_,
		_w12889_
	);
	LUT2 #(
		.INIT('h2)
	) name11540 (
		_w1565_,
		_w12889_,
		_w12890_
	);
	LUT3 #(
		.INIT('h08)
	) name11541 (
		\P2_EAX_reg[11]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12891_
	);
	LUT4 #(
		.INIT('haa02)
	) name11542 (
		\P2_lWord_reg[11]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12892_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11543 (
		_w1678_,
		_w12891_,
		_w12892_,
		_w12890_,
		_w12893_
	);
	LUT2 #(
		.INIT('he)
	) name11544 (
		_w12886_,
		_w12893_,
		_w12894_
	);
	LUT2 #(
		.INIT('h2)
	) name11545 (
		\P1_EAX_reg[24]/NET0131 ,
		_w9102_,
		_w12895_
	);
	LUT3 #(
		.INIT('ha2)
	) name11546 (
		\P1_EAX_reg[24]/NET0131 ,
		_w9437_,
		_w12860_,
		_w12896_
	);
	LUT3 #(
		.INIT('h40)
	) name11547 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1804_,
		_w1826_,
		_w12897_
	);
	LUT4 #(
		.INIT('h8000)
	) name11548 (
		\P1_EAX_reg[23]/NET0131 ,
		_w9430_,
		_w9432_,
		_w12897_,
		_w12898_
	);
	LUT3 #(
		.INIT('hd1)
	) name11549 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1867_,
		_w3435_,
		_w12899_
	);
	LUT2 #(
		.INIT('h2)
	) name11550 (
		_w1795_,
		_w12899_,
		_w12900_
	);
	LUT3 #(
		.INIT('h82)
	) name11551 (
		_w1846_,
		_w9015_,
		_w9026_,
		_w12901_
	);
	LUT4 #(
		.INIT('h4000)
	) name11552 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w12901_,
		_w12902_
	);
	LUT3 #(
		.INIT('hd1)
	) name11553 (
		\P1_EAX_reg[24]/NET0131 ,
		_w1867_,
		_w3516_,
		_w12903_
	);
	LUT3 #(
		.INIT('h08)
	) name11554 (
		_w1725_,
		_w1802_,
		_w12903_,
		_w12904_
	);
	LUT3 #(
		.INIT('h01)
	) name11555 (
		_w12902_,
		_w12904_,
		_w12900_,
		_w12905_
	);
	LUT2 #(
		.INIT('h4)
	) name11556 (
		_w12898_,
		_w12905_,
		_w12906_
	);
	LUT4 #(
		.INIT('hecee)
	) name11557 (
		_w1933_,
		_w12895_,
		_w12896_,
		_w12906_,
		_w12907_
	);
	LUT2 #(
		.INIT('h2)
	) name11558 (
		\P2_lWord_reg[12]/NET0131 ,
		_w7767_,
		_w12908_
	);
	LUT3 #(
		.INIT('h80)
	) name11559 (
		\P2_lWord_reg[12]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12909_
	);
	LUT3 #(
		.INIT('h0b)
	) name11560 (
		_w1602_,
		_w9451_,
		_w12909_,
		_w12910_
	);
	LUT2 #(
		.INIT('h2)
	) name11561 (
		_w1565_,
		_w12910_,
		_w12911_
	);
	LUT3 #(
		.INIT('h08)
	) name11562 (
		\P2_EAX_reg[12]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12912_
	);
	LUT4 #(
		.INIT('haa02)
	) name11563 (
		\P2_lWord_reg[12]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12913_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11564 (
		_w1678_,
		_w12912_,
		_w12913_,
		_w12911_,
		_w12914_
	);
	LUT2 #(
		.INIT('he)
	) name11565 (
		_w12908_,
		_w12914_,
		_w12915_
	);
	LUT2 #(
		.INIT('h2)
	) name11566 (
		\P2_lWord_reg[13]/NET0131 ,
		_w7767_,
		_w12916_
	);
	LUT3 #(
		.INIT('h80)
	) name11567 (
		\P2_lWord_reg[13]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12917_
	);
	LUT3 #(
		.INIT('h0d)
	) name11568 (
		_w1606_,
		_w9702_,
		_w12917_,
		_w12918_
	);
	LUT2 #(
		.INIT('h2)
	) name11569 (
		_w1565_,
		_w12918_,
		_w12919_
	);
	LUT4 #(
		.INIT('haa02)
	) name11570 (
		\P2_lWord_reg[13]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12920_
	);
	LUT3 #(
		.INIT('h08)
	) name11571 (
		\P2_EAX_reg[13]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12921_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11572 (
		_w1678_,
		_w12920_,
		_w12919_,
		_w12921_,
		_w12922_
	);
	LUT2 #(
		.INIT('he)
	) name11573 (
		_w12916_,
		_w12922_,
		_w12923_
	);
	LUT2 #(
		.INIT('h2)
	) name11574 (
		\P2_lWord_reg[14]/NET0131 ,
		_w7767_,
		_w12924_
	);
	LUT3 #(
		.INIT('h80)
	) name11575 (
		\P2_lWord_reg[14]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12925_
	);
	LUT3 #(
		.INIT('h07)
	) name11576 (
		_w1606_,
		_w8937_,
		_w12925_,
		_w12926_
	);
	LUT2 #(
		.INIT('h2)
	) name11577 (
		_w1565_,
		_w12926_,
		_w12927_
	);
	LUT4 #(
		.INIT('haa02)
	) name11578 (
		\P2_lWord_reg[14]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12928_
	);
	LUT3 #(
		.INIT('h08)
	) name11579 (
		\P2_EAX_reg[14]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12929_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11580 (
		_w1678_,
		_w12928_,
		_w12927_,
		_w12929_,
		_w12930_
	);
	LUT2 #(
		.INIT('he)
	) name11581 (
		_w12924_,
		_w12930_,
		_w12931_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11582 (
		\P2_lWord_reg[15]/NET0131 ,
		_w1678_,
		_w7767_,
		_w9467_,
		_w12932_
	);
	LUT4 #(
		.INIT('h135f)
	) name11583 (
		\P2_EAX_reg[15]/NET0131 ,
		_w1565_,
		_w1566_,
		_w9692_,
		_w12933_
	);
	LUT2 #(
		.INIT('h2)
	) name11584 (
		_w10009_,
		_w12933_,
		_w12934_
	);
	LUT2 #(
		.INIT('he)
	) name11585 (
		_w12932_,
		_w12934_,
		_w12935_
	);
	LUT3 #(
		.INIT('h80)
	) name11586 (
		\P2_lWord_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12936_
	);
	LUT3 #(
		.INIT('h0d)
	) name11587 (
		_w1606_,
		_w7156_,
		_w12936_,
		_w12937_
	);
	LUT2 #(
		.INIT('h2)
	) name11588 (
		_w1565_,
		_w12937_,
		_w12938_
	);
	LUT4 #(
		.INIT('haa02)
	) name11589 (
		\P2_lWord_reg[1]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12939_
	);
	LUT3 #(
		.INIT('h08)
	) name11590 (
		\P2_EAX_reg[1]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12940_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11591 (
		_w1678_,
		_w12939_,
		_w12938_,
		_w12940_,
		_w12941_
	);
	LUT2 #(
		.INIT('h2)
	) name11592 (
		\P2_lWord_reg[1]/NET0131 ,
		_w7767_,
		_w12942_
	);
	LUT2 #(
		.INIT('he)
	) name11593 (
		_w12941_,
		_w12942_,
		_w12943_
	);
	LUT3 #(
		.INIT('h80)
	) name11594 (
		\P2_lWord_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12944_
	);
	LUT3 #(
		.INIT('h0d)
	) name11595 (
		_w1606_,
		_w5487_,
		_w12944_,
		_w12945_
	);
	LUT2 #(
		.INIT('h2)
	) name11596 (
		_w1565_,
		_w12945_,
		_w12946_
	);
	LUT4 #(
		.INIT('haa02)
	) name11597 (
		\P2_lWord_reg[2]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12947_
	);
	LUT3 #(
		.INIT('h08)
	) name11598 (
		\P2_EAX_reg[2]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12948_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11599 (
		_w1678_,
		_w12947_,
		_w12946_,
		_w12948_,
		_w12949_
	);
	LUT2 #(
		.INIT('h2)
	) name11600 (
		\P2_lWord_reg[2]/NET0131 ,
		_w7767_,
		_w12950_
	);
	LUT2 #(
		.INIT('he)
	) name11601 (
		_w12949_,
		_w12950_,
		_w12951_
	);
	LUT3 #(
		.INIT('h80)
	) name11602 (
		\P2_lWord_reg[3]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12952_
	);
	LUT3 #(
		.INIT('h0d)
	) name11603 (
		_w1606_,
		_w3561_,
		_w12952_,
		_w12953_
	);
	LUT2 #(
		.INIT('h2)
	) name11604 (
		_w1565_,
		_w12953_,
		_w12954_
	);
	LUT4 #(
		.INIT('haa02)
	) name11605 (
		\P2_lWord_reg[3]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12955_
	);
	LUT3 #(
		.INIT('h08)
	) name11606 (
		\P2_EAX_reg[3]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12956_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11607 (
		_w1678_,
		_w12955_,
		_w12954_,
		_w12956_,
		_w12957_
	);
	LUT2 #(
		.INIT('h2)
	) name11608 (
		\P2_lWord_reg[3]/NET0131 ,
		_w7767_,
		_w12958_
	);
	LUT2 #(
		.INIT('he)
	) name11609 (
		_w12957_,
		_w12958_,
		_w12959_
	);
	LUT3 #(
		.INIT('h80)
	) name11610 (
		\P2_lWord_reg[4]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12960_
	);
	LUT3 #(
		.INIT('h0d)
	) name11611 (
		_w1606_,
		_w2276_,
		_w12960_,
		_w12961_
	);
	LUT2 #(
		.INIT('h2)
	) name11612 (
		_w1565_,
		_w12961_,
		_w12962_
	);
	LUT4 #(
		.INIT('haa02)
	) name11613 (
		\P2_lWord_reg[4]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12963_
	);
	LUT3 #(
		.INIT('h08)
	) name11614 (
		\P2_EAX_reg[4]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12964_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11615 (
		_w1678_,
		_w12963_,
		_w12962_,
		_w12964_,
		_w12965_
	);
	LUT2 #(
		.INIT('h2)
	) name11616 (
		\P2_lWord_reg[4]/NET0131 ,
		_w7767_,
		_w12966_
	);
	LUT2 #(
		.INIT('he)
	) name11617 (
		_w12965_,
		_w12966_,
		_w12967_
	);
	LUT3 #(
		.INIT('h80)
	) name11618 (
		\P2_lWord_reg[5]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12968_
	);
	LUT3 #(
		.INIT('h0d)
	) name11619 (
		_w1606_,
		_w6502_,
		_w12968_,
		_w12969_
	);
	LUT2 #(
		.INIT('h2)
	) name11620 (
		_w1565_,
		_w12969_,
		_w12970_
	);
	LUT4 #(
		.INIT('haa02)
	) name11621 (
		\P2_lWord_reg[5]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12971_
	);
	LUT3 #(
		.INIT('h08)
	) name11622 (
		\P2_EAX_reg[5]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12972_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11623 (
		_w1678_,
		_w12971_,
		_w12970_,
		_w12972_,
		_w12973_
	);
	LUT2 #(
		.INIT('h2)
	) name11624 (
		\P2_lWord_reg[5]/NET0131 ,
		_w7767_,
		_w12974_
	);
	LUT2 #(
		.INIT('he)
	) name11625 (
		_w12973_,
		_w12974_,
		_w12975_
	);
	LUT3 #(
		.INIT('h80)
	) name11626 (
		\P2_lWord_reg[6]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12976_
	);
	LUT3 #(
		.INIT('h54)
	) name11627 (
		_w1605_,
		_w4975_,
		_w4976_,
		_w12977_
	);
	LUT3 #(
		.INIT('h23)
	) name11628 (
		_w1602_,
		_w12976_,
		_w12977_,
		_w12978_
	);
	LUT2 #(
		.INIT('h2)
	) name11629 (
		_w1565_,
		_w12978_,
		_w12979_
	);
	LUT3 #(
		.INIT('h08)
	) name11630 (
		\P2_EAX_reg[6]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12980_
	);
	LUT4 #(
		.INIT('haa02)
	) name11631 (
		\P2_lWord_reg[6]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12981_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11632 (
		_w1678_,
		_w12980_,
		_w12981_,
		_w12979_,
		_w12982_
	);
	LUT2 #(
		.INIT('h2)
	) name11633 (
		\P2_lWord_reg[6]/NET0131 ,
		_w7767_,
		_w12983_
	);
	LUT2 #(
		.INIT('he)
	) name11634 (
		_w12982_,
		_w12983_,
		_w12984_
	);
	LUT3 #(
		.INIT('h80)
	) name11635 (
		\P2_lWord_reg[7]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12985_
	);
	LUT3 #(
		.INIT('h0d)
	) name11636 (
		_w1606_,
		_w2295_,
		_w12985_,
		_w12986_
	);
	LUT2 #(
		.INIT('h2)
	) name11637 (
		_w1565_,
		_w12986_,
		_w12987_
	);
	LUT4 #(
		.INIT('haa02)
	) name11638 (
		\P2_lWord_reg[7]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12988_
	);
	LUT3 #(
		.INIT('h08)
	) name11639 (
		\P2_EAX_reg[7]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12989_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11640 (
		_w1678_,
		_w12988_,
		_w12987_,
		_w12989_,
		_w12990_
	);
	LUT2 #(
		.INIT('h2)
	) name11641 (
		\P2_lWord_reg[7]/NET0131 ,
		_w7767_,
		_w12991_
	);
	LUT2 #(
		.INIT('he)
	) name11642 (
		_w12990_,
		_w12991_,
		_w12992_
	);
	LUT2 #(
		.INIT('h2)
	) name11643 (
		\P2_lWord_reg[8]/NET0131 ,
		_w7767_,
		_w12993_
	);
	LUT3 #(
		.INIT('h80)
	) name11644 (
		\P2_lWord_reg[8]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w12994_
	);
	LUT3 #(
		.INIT('h0b)
	) name11645 (
		_w1602_,
		_w10006_,
		_w12994_,
		_w12995_
	);
	LUT2 #(
		.INIT('h2)
	) name11646 (
		_w1565_,
		_w12995_,
		_w12996_
	);
	LUT3 #(
		.INIT('h08)
	) name11647 (
		\P2_EAX_reg[8]/NET0131 ,
		_w1566_,
		_w1602_,
		_w12997_
	);
	LUT4 #(
		.INIT('haa02)
	) name11648 (
		\P2_lWord_reg[8]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w12998_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11649 (
		_w1678_,
		_w12997_,
		_w12998_,
		_w12996_,
		_w12999_
	);
	LUT2 #(
		.INIT('he)
	) name11650 (
		_w12993_,
		_w12999_,
		_w13000_
	);
	LUT2 #(
		.INIT('h2)
	) name11651 (
		\P2_lWord_reg[9]/NET0131 ,
		_w7767_,
		_w13001_
	);
	LUT3 #(
		.INIT('h80)
	) name11652 (
		\P2_lWord_reg[9]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13002_
	);
	LUT3 #(
		.INIT('h07)
	) name11653 (
		_w1606_,
		_w10484_,
		_w13002_,
		_w13003_
	);
	LUT2 #(
		.INIT('h2)
	) name11654 (
		_w1565_,
		_w13003_,
		_w13004_
	);
	LUT4 #(
		.INIT('haa02)
	) name11655 (
		\P2_lWord_reg[9]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w13005_
	);
	LUT3 #(
		.INIT('h08)
	) name11656 (
		\P2_EAX_reg[9]/NET0131 ,
		_w1566_,
		_w1602_,
		_w13006_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11657 (
		_w1678_,
		_w13005_,
		_w13004_,
		_w13006_,
		_w13007_
	);
	LUT2 #(
		.INIT('he)
	) name11658 (
		_w13001_,
		_w13007_,
		_w13008_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11659 (
		\P2_uWord_reg[11]/NET0131 ,
		_w1678_,
		_w7767_,
		_w9467_,
		_w13009_
	);
	LUT4 #(
		.INIT('h60c0)
	) name11660 (
		\P2_EAX_reg[26]/NET0131 ,
		\P2_EAX_reg[27]/NET0131 ,
		_w1566_,
		_w9460_,
		_w13010_
	);
	LUT2 #(
		.INIT('h8)
	) name11661 (
		_w1565_,
		_w12888_,
		_w13011_
	);
	LUT3 #(
		.INIT('ha8)
	) name11662 (
		_w10009_,
		_w13010_,
		_w13011_,
		_w13012_
	);
	LUT2 #(
		.INIT('he)
	) name11663 (
		_w13009_,
		_w13012_,
		_w13013_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name11664 (
		\P1_uWord_reg[11]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w13014_
	);
	LUT3 #(
		.INIT('h02)
	) name11665 (
		_w1795_,
		_w1861_,
		_w3431_,
		_w13015_
	);
	LUT4 #(
		.INIT('haa20)
	) name11666 (
		_w9489_,
		_w12847_,
		_w12848_,
		_w13015_,
		_w13016_
	);
	LUT2 #(
		.INIT('he)
	) name11667 (
		_w13014_,
		_w13016_,
		_w13017_
	);
	LUT2 #(
		.INIT('h2)
	) name11668 (
		\P1_EAX_reg[28]/NET0131 ,
		_w9102_,
		_w13018_
	);
	LUT3 #(
		.INIT('h48)
	) name11669 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1827_,
		_w9655_,
		_w13019_
	);
	LUT2 #(
		.INIT('h2)
	) name11670 (
		_w1795_,
		_w1867_,
		_w13020_
	);
	LUT4 #(
		.INIT('h08a2)
	) name11671 (
		_w1846_,
		_w9050_,
		_w9061_,
		_w9072_,
		_w13021_
	);
	LUT2 #(
		.INIT('h8)
	) name11672 (
		_w1795_,
		_w10575_,
		_w13022_
	);
	LUT2 #(
		.INIT('h8)
	) name11673 (
		_w1867_,
		_w3529_,
		_w13023_
	);
	LUT4 #(
		.INIT('h5504)
	) name11674 (
		\P1_EAX_reg[28]/NET0131 ,
		_w1842_,
		_w1851_,
		_w1861_,
		_w13024_
	);
	LUT4 #(
		.INIT('h0008)
	) name11675 (
		_w1725_,
		_w1802_,
		_w13024_,
		_w13023_,
		_w13025_
	);
	LUT4 #(
		.INIT('h0013)
	) name11676 (
		_w1832_,
		_w13022_,
		_w13021_,
		_w13025_,
		_w13026_
	);
	LUT4 #(
		.INIT('h5d00)
	) name11677 (
		\P1_EAX_reg[28]/NET0131 ,
		_w9437_,
		_w13020_,
		_w13026_,
		_w13027_
	);
	LUT4 #(
		.INIT('hecee)
	) name11678 (
		_w1933_,
		_w13018_,
		_w13019_,
		_w13027_,
		_w13028_
	);
	LUT3 #(
		.INIT('h08)
	) name11679 (
		\buf2_reg[0]/NET0131 ,
		_w2108_,
		_w2116_,
		_w13029_
	);
	LUT3 #(
		.INIT('h0b)
	) name11680 (
		_w2794_,
		_w8366_,
		_w10149_,
		_w13030_
	);
	LUT3 #(
		.INIT('h8a)
	) name11681 (
		_w1945_,
		_w13029_,
		_w13030_,
		_w13031_
	);
	LUT4 #(
		.INIT('hffa2)
	) name11682 (
		\P3_EAX_reg[0]/NET0131 ,
		_w8341_,
		_w10089_,
		_w13031_,
		_w13032_
	);
	LUT2 #(
		.INIT('h2)
	) name11683 (
		\P3_EAX_reg[16]/NET0131 ,
		_w8341_,
		_w13033_
	);
	LUT3 #(
		.INIT('ha8)
	) name11684 (
		\P3_EAX_reg[16]/NET0131 ,
		_w8367_,
		_w10122_,
		_w13034_
	);
	LUT2 #(
		.INIT('h8)
	) name11685 (
		\P3_EAX_reg[16]/NET0131 ,
		_w8351_,
		_w13035_
	);
	LUT4 #(
		.INIT('h40c0)
	) name11686 (
		\P3_EAX_reg[16]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8351_,
		_w13036_
	);
	LUT4 #(
		.INIT('h4000)
	) name11687 (
		\P3_EAX_reg[16]/NET0131 ,
		_w2063_,
		_w2075_,
		_w8351_,
		_w13037_
	);
	LUT4 #(
		.INIT('h5553)
	) name11688 (
		\P3_EAX_reg[16]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13038_
	);
	LUT3 #(
		.INIT('h04)
	) name11689 (
		_w2060_,
		_w2047_,
		_w13038_,
		_w13039_
	);
	LUT4 #(
		.INIT('h135f)
	) name11690 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w1956_,
		_w1947_,
		_w13040_
	);
	LUT4 #(
		.INIT('h153f)
	) name11691 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w1946_,
		_w1950_,
		_w13041_
	);
	LUT4 #(
		.INIT('h153f)
	) name11692 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w1969_,
		_w1963_,
		_w13042_
	);
	LUT4 #(
		.INIT('h135f)
	) name11693 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w1966_,
		_w1967_,
		_w13043_
	);
	LUT4 #(
		.INIT('h8000)
	) name11694 (
		_w13042_,
		_w13043_,
		_w13040_,
		_w13041_,
		_w13044_
	);
	LUT4 #(
		.INIT('h135f)
	) name11695 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w1954_,
		_w1960_,
		_w13045_
	);
	LUT4 #(
		.INIT('h135f)
	) name11696 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w1957_,
		_w1949_,
		_w13046_
	);
	LUT4 #(
		.INIT('h135f)
	) name11697 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w1970_,
		_w1964_,
		_w13047_
	);
	LUT4 #(
		.INIT('h153f)
	) name11698 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w1952_,
		_w1961_,
		_w13048_
	);
	LUT4 #(
		.INIT('h8000)
	) name11699 (
		_w13047_,
		_w13048_,
		_w13045_,
		_w13046_,
		_w13049_
	);
	LUT2 #(
		.INIT('h8)
	) name11700 (
		_w13044_,
		_w13049_,
		_w13050_
	);
	LUT4 #(
		.INIT('h5553)
	) name11701 (
		\P3_EAX_reg[16]/NET0131 ,
		\buf2_reg[16]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13051_
	);
	LUT3 #(
		.INIT('h08)
	) name11702 (
		_w2060_,
		_w2044_,
		_w13051_,
		_w13052_
	);
	LUT4 #(
		.INIT('h000d)
	) name11703 (
		_w8366_,
		_w13050_,
		_w13052_,
		_w13039_,
		_w13053_
	);
	LUT2 #(
		.INIT('h4)
	) name11704 (
		_w13037_,
		_w13053_,
		_w13054_
	);
	LUT4 #(
		.INIT('hecee)
	) name11705 (
		_w1945_,
		_w13033_,
		_w13034_,
		_w13054_,
		_w13055_
	);
	LUT2 #(
		.INIT('h2)
	) name11706 (
		\P3_EAX_reg[17]/NET0131 ,
		_w8341_,
		_w13056_
	);
	LUT4 #(
		.INIT('h0001)
	) name11707 (
		_w2120_,
		_w2121_,
		_w8367_,
		_w13036_,
		_w13057_
	);
	LUT3 #(
		.INIT('h40)
	) name11708 (
		\P3_EAX_reg[17]/NET0131 ,
		_w2063_,
		_w2075_,
		_w13058_
	);
	LUT2 #(
		.INIT('h8)
	) name11709 (
		_w13035_,
		_w13058_,
		_w13059_
	);
	LUT4 #(
		.INIT('h153f)
	) name11710 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w1952_,
		_w1961_,
		_w13060_
	);
	LUT4 #(
		.INIT('h153f)
	) name11711 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w1956_,
		_w1963_,
		_w13061_
	);
	LUT4 #(
		.INIT('h135f)
	) name11712 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w1950_,
		_w1967_,
		_w13062_
	);
	LUT4 #(
		.INIT('h153f)
	) name11713 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w1947_,
		_w1960_,
		_w13063_
	);
	LUT4 #(
		.INIT('h8000)
	) name11714 (
		_w13062_,
		_w13063_,
		_w13060_,
		_w13061_,
		_w13064_
	);
	LUT4 #(
		.INIT('h135f)
	) name11715 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w1957_,
		_w1949_,
		_w13065_
	);
	LUT4 #(
		.INIT('h153f)
	) name11716 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w1969_,
		_w1970_,
		_w13066_
	);
	LUT4 #(
		.INIT('h135f)
	) name11717 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w1954_,
		_w1964_,
		_w13067_
	);
	LUT4 #(
		.INIT('h153f)
	) name11718 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w1946_,
		_w1966_,
		_w13068_
	);
	LUT4 #(
		.INIT('h8000)
	) name11719 (
		_w13067_,
		_w13068_,
		_w13065_,
		_w13066_,
		_w13069_
	);
	LUT2 #(
		.INIT('h8)
	) name11720 (
		_w13064_,
		_w13069_,
		_w13070_
	);
	LUT2 #(
		.INIT('h2)
	) name11721 (
		_w8366_,
		_w13070_,
		_w13071_
	);
	LUT3 #(
		.INIT('h20)
	) name11722 (
		\buf2_reg[1]/NET0131 ,
		_w2060_,
		_w2047_,
		_w13072_
	);
	LUT3 #(
		.INIT('h80)
	) name11723 (
		\buf2_reg[17]/NET0131 ,
		_w2060_,
		_w2044_,
		_w13073_
	);
	LUT3 #(
		.INIT('ha8)
	) name11724 (
		_w2119_,
		_w13072_,
		_w13073_,
		_w13074_
	);
	LUT3 #(
		.INIT('h01)
	) name11725 (
		_w13059_,
		_w13071_,
		_w13074_,
		_w13075_
	);
	LUT4 #(
		.INIT('h08cc)
	) name11726 (
		\P3_EAX_reg[17]/NET0131 ,
		_w1945_,
		_w13057_,
		_w13075_,
		_w13076_
	);
	LUT2 #(
		.INIT('he)
	) name11727 (
		_w13056_,
		_w13076_,
		_w13077_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name11728 (
		\P3_EAX_reg[18]/NET0131 ,
		_w1945_,
		_w8341_,
		_w8367_,
		_w13078_
	);
	LUT4 #(
		.INIT('h070f)
	) name11729 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[18]/NET0131 ,
		_w8351_,
		_w13079_
	);
	LUT4 #(
		.INIT('h0888)
	) name11730 (
		_w2063_,
		_w2075_,
		_w8351_,
		_w8353_,
		_w13080_
	);
	LUT2 #(
		.INIT('h4)
	) name11731 (
		_w13079_,
		_w13080_,
		_w13081_
	);
	LUT4 #(
		.INIT('h5553)
	) name11732 (
		\P3_EAX_reg[18]/NET0131 ,
		\buf2_reg[18]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13082_
	);
	LUT3 #(
		.INIT('h08)
	) name11733 (
		_w2060_,
		_w2044_,
		_w13082_,
		_w13083_
	);
	LUT4 #(
		.INIT('h5553)
	) name11734 (
		\P3_EAX_reg[18]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13084_
	);
	LUT3 #(
		.INIT('h04)
	) name11735 (
		_w2060_,
		_w2047_,
		_w13084_,
		_w13085_
	);
	LUT4 #(
		.INIT('h135f)
	) name11736 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w1957_,
		_w1967_,
		_w13086_
	);
	LUT4 #(
		.INIT('h135f)
	) name11737 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w1952_,
		_w1949_,
		_w13087_
	);
	LUT4 #(
		.INIT('h135f)
	) name11738 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w1961_,
		_w1964_,
		_w13088_
	);
	LUT4 #(
		.INIT('h135f)
	) name11739 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w1954_,
		_w1950_,
		_w13089_
	);
	LUT4 #(
		.INIT('h8000)
	) name11740 (
		_w13088_,
		_w13089_,
		_w13086_,
		_w13087_,
		_w13090_
	);
	LUT4 #(
		.INIT('h153f)
	) name11741 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w1956_,
		_w1963_,
		_w13091_
	);
	LUT4 #(
		.INIT('h135f)
	) name11742 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w1966_,
		_w1970_,
		_w13092_
	);
	LUT4 #(
		.INIT('h153f)
	) name11743 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w1946_,
		_w1960_,
		_w13093_
	);
	LUT4 #(
		.INIT('h135f)
	) name11744 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w1947_,
		_w1969_,
		_w13094_
	);
	LUT4 #(
		.INIT('h8000)
	) name11745 (
		_w13093_,
		_w13094_,
		_w13091_,
		_w13092_,
		_w13095_
	);
	LUT2 #(
		.INIT('h8)
	) name11746 (
		_w13090_,
		_w13095_,
		_w13096_
	);
	LUT4 #(
		.INIT('h0031)
	) name11747 (
		_w8366_,
		_w13085_,
		_w13096_,
		_w13083_,
		_w13097_
	);
	LUT3 #(
		.INIT('h8a)
	) name11748 (
		_w1945_,
		_w13081_,
		_w13097_,
		_w13098_
	);
	LUT2 #(
		.INIT('he)
	) name11749 (
		_w13078_,
		_w13098_,
		_w13099_
	);
	LUT2 #(
		.INIT('h2)
	) name11750 (
		\P3_EAX_reg[19]/NET0131 ,
		_w8341_,
		_w13100_
	);
	LUT3 #(
		.INIT('h48)
	) name11751 (
		\P3_EAX_reg[19]/NET0131 ,
		_w8361_,
		_w8354_,
		_w13101_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11752 (
		\P3_EAX_reg[19]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w13102_
	);
	LUT4 #(
		.INIT('h135f)
	) name11753 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w1956_,
		_w1947_,
		_w13103_
	);
	LUT4 #(
		.INIT('h153f)
	) name11754 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w1946_,
		_w1950_,
		_w13104_
	);
	LUT4 #(
		.INIT('h153f)
	) name11755 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w1969_,
		_w1963_,
		_w13105_
	);
	LUT4 #(
		.INIT('h135f)
	) name11756 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w1966_,
		_w1967_,
		_w13106_
	);
	LUT4 #(
		.INIT('h8000)
	) name11757 (
		_w13105_,
		_w13106_,
		_w13103_,
		_w13104_,
		_w13107_
	);
	LUT4 #(
		.INIT('h135f)
	) name11758 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w1954_,
		_w1960_,
		_w13108_
	);
	LUT4 #(
		.INIT('h135f)
	) name11759 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w1957_,
		_w1949_,
		_w13109_
	);
	LUT4 #(
		.INIT('h135f)
	) name11760 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w1970_,
		_w1964_,
		_w13110_
	);
	LUT4 #(
		.INIT('h153f)
	) name11761 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w1952_,
		_w1961_,
		_w13111_
	);
	LUT4 #(
		.INIT('h8000)
	) name11762 (
		_w13110_,
		_w13111_,
		_w13108_,
		_w13109_,
		_w13112_
	);
	LUT2 #(
		.INIT('h8)
	) name11763 (
		_w13107_,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h2)
	) name11764 (
		_w8366_,
		_w13113_,
		_w13114_
	);
	LUT3 #(
		.INIT('h80)
	) name11765 (
		\buf2_reg[19]/NET0131 ,
		_w2060_,
		_w2044_,
		_w13115_
	);
	LUT3 #(
		.INIT('h20)
	) name11766 (
		\buf2_reg[3]/NET0131 ,
		_w2060_,
		_w2047_,
		_w13116_
	);
	LUT3 #(
		.INIT('ha8)
	) name11767 (
		_w2119_,
		_w13115_,
		_w13116_,
		_w13117_
	);
	LUT2 #(
		.INIT('h1)
	) name11768 (
		_w13114_,
		_w13117_,
		_w13118_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11769 (
		_w1945_,
		_w13102_,
		_w13101_,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('he)
	) name11770 (
		_w13100_,
		_w13119_,
		_w13120_
	);
	LUT4 #(
		.INIT('h5070)
	) name11771 (
		_w1945_,
		_w2121_,
		_w8341_,
		_w8367_,
		_w13121_
	);
	LUT3 #(
		.INIT('h48)
	) name11772 (
		\P3_EAX_reg[20]/NET0131 ,
		_w8361_,
		_w8355_,
		_w13122_
	);
	LUT4 #(
		.INIT('h5553)
	) name11773 (
		\P3_EAX_reg[20]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13123_
	);
	LUT3 #(
		.INIT('h04)
	) name11774 (
		_w2060_,
		_w2047_,
		_w13123_,
		_w13124_
	);
	LUT4 #(
		.INIT('h135f)
	) name11775 (
		\P3_InstQueue_reg[5][4]/NET0131 ,
		\P3_InstQueue_reg[6][4]/NET0131 ,
		_w1957_,
		_w1967_,
		_w13125_
	);
	LUT4 #(
		.INIT('h135f)
	) name11776 (
		\P3_InstQueue_reg[4][4]/NET0131 ,
		\P3_InstQueue_reg[9][4]/NET0131 ,
		_w1952_,
		_w1949_,
		_w13126_
	);
	LUT4 #(
		.INIT('h135f)
	) name11777 (
		\P3_InstQueue_reg[1][4]/NET0131 ,
		\P3_InstQueue_reg[8][4]/NET0131 ,
		_w1961_,
		_w1964_,
		_w13127_
	);
	LUT4 #(
		.INIT('h135f)
	) name11778 (
		\P3_InstQueue_reg[10][4]/NET0131 ,
		\P3_InstQueue_reg[11][4]/NET0131 ,
		_w1954_,
		_w1950_,
		_w13128_
	);
	LUT4 #(
		.INIT('h8000)
	) name11779 (
		_w13127_,
		_w13128_,
		_w13125_,
		_w13126_,
		_w13129_
	);
	LUT4 #(
		.INIT('h153f)
	) name11780 (
		\P3_InstQueue_reg[12][4]/NET0131 ,
		\P3_InstQueue_reg[13][4]/NET0131 ,
		_w1956_,
		_w1963_,
		_w13130_
	);
	LUT4 #(
		.INIT('h135f)
	) name11781 (
		\P3_InstQueue_reg[0][4]/NET0131 ,
		\P3_InstQueue_reg[2][4]/NET0131 ,
		_w1966_,
		_w1970_,
		_w13131_
	);
	LUT4 #(
		.INIT('h153f)
	) name11782 (
		\P3_InstQueue_reg[14][4]/NET0131 ,
		\P3_InstQueue_reg[7][4]/NET0131 ,
		_w1946_,
		_w1960_,
		_w13132_
	);
	LUT4 #(
		.INIT('h135f)
	) name11783 (
		\P3_InstQueue_reg[15][4]/NET0131 ,
		\P3_InstQueue_reg[3][4]/NET0131 ,
		_w1947_,
		_w1969_,
		_w13133_
	);
	LUT4 #(
		.INIT('h8000)
	) name11784 (
		_w13132_,
		_w13133_,
		_w13130_,
		_w13131_,
		_w13134_
	);
	LUT2 #(
		.INIT('h8)
	) name11785 (
		_w13129_,
		_w13134_,
		_w13135_
	);
	LUT4 #(
		.INIT('h8000)
	) name11786 (
		\buf2_reg[20]/NET0131 ,
		_w2060_,
		_w2044_,
		_w2119_,
		_w13136_
	);
	LUT4 #(
		.INIT('h000d)
	) name11787 (
		_w8366_,
		_w13135_,
		_w13124_,
		_w13136_,
		_w13137_
	);
	LUT3 #(
		.INIT('h8a)
	) name11788 (
		_w1945_,
		_w13122_,
		_w13137_,
		_w13138_
	);
	LUT3 #(
		.INIT('hf2)
	) name11789 (
		\P3_EAX_reg[20]/NET0131 ,
		_w13121_,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h2)
	) name11790 (
		\P3_EAX_reg[21]/NET0131 ,
		_w8341_,
		_w13140_
	);
	LUT3 #(
		.INIT('h48)
	) name11791 (
		\P3_EAX_reg[21]/NET0131 ,
		_w8361_,
		_w8356_,
		_w13141_
	);
	LUT4 #(
		.INIT('haaa8)
	) name11792 (
		\P3_EAX_reg[21]/NET0131 ,
		_w2120_,
		_w2121_,
		_w8367_,
		_w13142_
	);
	LUT4 #(
		.INIT('h135f)
	) name11793 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w1956_,
		_w1947_,
		_w13143_
	);
	LUT4 #(
		.INIT('h153f)
	) name11794 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w1946_,
		_w1950_,
		_w13144_
	);
	LUT4 #(
		.INIT('h153f)
	) name11795 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w1969_,
		_w1963_,
		_w13145_
	);
	LUT4 #(
		.INIT('h135f)
	) name11796 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w1966_,
		_w1967_,
		_w13146_
	);
	LUT4 #(
		.INIT('h8000)
	) name11797 (
		_w13145_,
		_w13146_,
		_w13143_,
		_w13144_,
		_w13147_
	);
	LUT4 #(
		.INIT('h135f)
	) name11798 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w1954_,
		_w1960_,
		_w13148_
	);
	LUT4 #(
		.INIT('h135f)
	) name11799 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w1957_,
		_w1949_,
		_w13149_
	);
	LUT4 #(
		.INIT('h135f)
	) name11800 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w1970_,
		_w1964_,
		_w13150_
	);
	LUT4 #(
		.INIT('h153f)
	) name11801 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w1952_,
		_w1961_,
		_w13151_
	);
	LUT4 #(
		.INIT('h8000)
	) name11802 (
		_w13150_,
		_w13151_,
		_w13148_,
		_w13149_,
		_w13152_
	);
	LUT2 #(
		.INIT('h8)
	) name11803 (
		_w13147_,
		_w13152_,
		_w13153_
	);
	LUT2 #(
		.INIT('h2)
	) name11804 (
		_w8366_,
		_w13153_,
		_w13154_
	);
	LUT3 #(
		.INIT('h80)
	) name11805 (
		\buf2_reg[21]/NET0131 ,
		_w2060_,
		_w2044_,
		_w13155_
	);
	LUT3 #(
		.INIT('h20)
	) name11806 (
		\buf2_reg[5]/NET0131 ,
		_w2060_,
		_w2047_,
		_w13156_
	);
	LUT3 #(
		.INIT('ha8)
	) name11807 (
		_w2119_,
		_w13155_,
		_w13156_,
		_w13157_
	);
	LUT2 #(
		.INIT('h1)
	) name11808 (
		_w13154_,
		_w13157_,
		_w13158_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11809 (
		_w1945_,
		_w13142_,
		_w13141_,
		_w13158_,
		_w13159_
	);
	LUT2 #(
		.INIT('he)
	) name11810 (
		_w13140_,
		_w13159_,
		_w13160_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name11811 (
		\P3_EAX_reg[22]/NET0131 ,
		_w1945_,
		_w8341_,
		_w8367_,
		_w13161_
	);
	LUT4 #(
		.INIT('h70f0)
	) name11812 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		_w8361_,
		_w8356_,
		_w13162_
	);
	LUT4 #(
		.INIT('h60c0)
	) name11813 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		_w8361_,
		_w8356_,
		_w13163_
	);
	LUT4 #(
		.INIT('h5553)
	) name11814 (
		\P3_EAX_reg[22]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13164_
	);
	LUT3 #(
		.INIT('h04)
	) name11815 (
		_w2060_,
		_w2047_,
		_w13164_,
		_w13165_
	);
	LUT4 #(
		.INIT('h135f)
	) name11816 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w1957_,
		_w1946_,
		_w13166_
	);
	LUT4 #(
		.INIT('h135f)
	) name11817 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w1947_,
		_w1964_,
		_w13167_
	);
	LUT4 #(
		.INIT('h153f)
	) name11818 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w1949_,
		_w1966_,
		_w13168_
	);
	LUT4 #(
		.INIT('h153f)
	) name11819 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w1969_,
		_w1961_,
		_w13169_
	);
	LUT4 #(
		.INIT('h8000)
	) name11820 (
		_w13168_,
		_w13169_,
		_w13166_,
		_w13167_,
		_w13170_
	);
	LUT4 #(
		.INIT('h135f)
	) name11821 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w1954_,
		_w1960_,
		_w13171_
	);
	LUT4 #(
		.INIT('h153f)
	) name11822 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w1952_,
		_w1956_,
		_w13172_
	);
	LUT4 #(
		.INIT('h135f)
	) name11823 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w1950_,
		_w1970_,
		_w13173_
	);
	LUT4 #(
		.INIT('h153f)
	) name11824 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w1967_,
		_w1963_,
		_w13174_
	);
	LUT4 #(
		.INIT('h8000)
	) name11825 (
		_w13173_,
		_w13174_,
		_w13171_,
		_w13172_,
		_w13175_
	);
	LUT2 #(
		.INIT('h8)
	) name11826 (
		_w13170_,
		_w13175_,
		_w13176_
	);
	LUT4 #(
		.INIT('h5553)
	) name11827 (
		\P3_EAX_reg[22]/NET0131 ,
		\buf2_reg[22]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13177_
	);
	LUT3 #(
		.INIT('h08)
	) name11828 (
		_w2060_,
		_w2044_,
		_w13177_,
		_w13178_
	);
	LUT4 #(
		.INIT('h000d)
	) name11829 (
		_w8366_,
		_w13176_,
		_w13178_,
		_w13165_,
		_w13179_
	);
	LUT3 #(
		.INIT('h8a)
	) name11830 (
		_w1945_,
		_w13163_,
		_w13179_,
		_w13180_
	);
	LUT2 #(
		.INIT('he)
	) name11831 (
		_w13161_,
		_w13180_,
		_w13181_
	);
	LUT2 #(
		.INIT('h2)
	) name11832 (
		\P3_EAX_reg[23]/NET0131 ,
		_w8341_,
		_w13182_
	);
	LUT3 #(
		.INIT('ha8)
	) name11833 (
		\P3_EAX_reg[23]/NET0131 ,
		_w8367_,
		_w13162_,
		_w13183_
	);
	LUT3 #(
		.INIT('h40)
	) name11834 (
		\P3_EAX_reg[23]/NET0131 ,
		_w2063_,
		_w2075_,
		_w13184_
	);
	LUT4 #(
		.INIT('h8000)
	) name11835 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		_w8356_,
		_w13184_,
		_w13185_
	);
	LUT3 #(
		.INIT('h02)
	) name11836 (
		\buf2_reg[7]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13186_
	);
	LUT4 #(
		.INIT('h5553)
	) name11837 (
		\P3_EAX_reg[23]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13187_
	);
	LUT3 #(
		.INIT('h04)
	) name11838 (
		_w2060_,
		_w2047_,
		_w13187_,
		_w13188_
	);
	LUT4 #(
		.INIT('h7888)
	) name11839 (
		_w8375_,
		_w8380_,
		_w8385_,
		_w8390_,
		_w13189_
	);
	LUT4 #(
		.INIT('h5553)
	) name11840 (
		\P3_EAX_reg[23]/NET0131 ,
		\buf2_reg[23]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13190_
	);
	LUT3 #(
		.INIT('h08)
	) name11841 (
		_w2060_,
		_w2044_,
		_w13190_,
		_w13191_
	);
	LUT4 #(
		.INIT('h0007)
	) name11842 (
		_w8366_,
		_w13189_,
		_w13191_,
		_w13188_,
		_w13192_
	);
	LUT2 #(
		.INIT('h4)
	) name11843 (
		_w13185_,
		_w13192_,
		_w13193_
	);
	LUT4 #(
		.INIT('hecee)
	) name11844 (
		_w1945_,
		_w13182_,
		_w13183_,
		_w13193_,
		_w13194_
	);
	LUT2 #(
		.INIT('h2)
	) name11845 (
		\P3_EAX_reg[24]/NET0131 ,
		_w8341_,
		_w13195_
	);
	LUT4 #(
		.INIT('h8000)
	) name11846 (
		\P3_EAX_reg[21]/NET0131 ,
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		_w8356_,
		_w13196_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name11847 (
		\P3_EAX_reg[24]/NET0131 ,
		_w8361_,
		_w8367_,
		_w13196_,
		_w13197_
	);
	LUT3 #(
		.INIT('h40)
	) name11848 (
		\P3_EAX_reg[24]/NET0131 ,
		_w2063_,
		_w2075_,
		_w13198_
	);
	LUT4 #(
		.INIT('h5553)
	) name11849 (
		\P3_EAX_reg[24]/NET0131 ,
		\buf2_reg[8]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13199_
	);
	LUT3 #(
		.INIT('h04)
	) name11850 (
		_w2060_,
		_w2047_,
		_w13199_,
		_w13200_
	);
	LUT2 #(
		.INIT('h9)
	) name11851 (
		_w8391_,
		_w8402_,
		_w13201_
	);
	LUT4 #(
		.INIT('h5553)
	) name11852 (
		\P3_EAX_reg[24]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w2105_,
		_w2116_,
		_w13202_
	);
	LUT3 #(
		.INIT('h08)
	) name11853 (
		_w2060_,
		_w2044_,
		_w13202_,
		_w13203_
	);
	LUT4 #(
		.INIT('h0007)
	) name11854 (
		_w8366_,
		_w13201_,
		_w13203_,
		_w13200_,
		_w13204_
	);
	LUT3 #(
		.INIT('h70)
	) name11855 (
		_w13196_,
		_w13198_,
		_w13204_,
		_w13205_
	);
	LUT4 #(
		.INIT('hecee)
	) name11856 (
		_w1945_,
		_w13195_,
		_w13197_,
		_w13205_,
		_w13206_
	);
	LUT2 #(
		.INIT('h2)
	) name11857 (
		\P3_EAX_reg[28]/NET0131 ,
		_w8341_,
		_w13207_
	);
	LUT3 #(
		.INIT('h40)
	) name11858 (
		\P3_EAX_reg[28]/NET0131 ,
		_w2063_,
		_w2075_,
		_w13208_
	);
	LUT3 #(
		.INIT('h2d)
	) name11859 (
		_w8426_,
		_w8437_,
		_w8867_,
		_w13209_
	);
	LUT2 #(
		.INIT('h8)
	) name11860 (
		_w8366_,
		_w13209_,
		_w13210_
	);
	LUT3 #(
		.INIT('h20)
	) name11861 (
		\buf2_reg[12]/NET0131 ,
		_w2060_,
		_w2047_,
		_w13211_
	);
	LUT3 #(
		.INIT('h80)
	) name11862 (
		\buf2_reg[28]/NET0131 ,
		_w2060_,
		_w2044_,
		_w13212_
	);
	LUT3 #(
		.INIT('ha8)
	) name11863 (
		_w2119_,
		_w13211_,
		_w13212_,
		_w13213_
	);
	LUT4 #(
		.INIT('h0007)
	) name11864 (
		_w8363_,
		_w13208_,
		_w13210_,
		_w13213_,
		_w13214_
	);
	LUT4 #(
		.INIT('h7500)
	) name11865 (
		\P3_EAX_reg[28]/NET0131 ,
		_w8364_,
		_w8892_,
		_w13214_,
		_w13215_
	);
	LUT3 #(
		.INIT('hce)
	) name11866 (
		_w1945_,
		_w13207_,
		_w13215_,
		_w13216_
	);
	LUT2 #(
		.INIT('h2)
	) name11867 (
		\P3_Flush_reg/NET0131 ,
		_w8341_,
		_w13217_
	);
	LUT3 #(
		.INIT('hf2)
	) name11868 (
		_w1945_,
		_w2183_,
		_w13217_,
		_w13218_
	);
	LUT2 #(
		.INIT('h2)
	) name11869 (
		\P2_EAX_reg[16]/NET0131 ,
		_w7767_,
		_w13219_
	);
	LUT3 #(
		.INIT('ha2)
	) name11870 (
		\P2_EAX_reg[16]/NET0131 ,
		_w7792_,
		_w9676_,
		_w13220_
	);
	LUT3 #(
		.INIT('h40)
	) name11871 (
		\P2_EAX_reg[16]/NET0131 ,
		_w7777_,
		_w7789_,
		_w13221_
	);
	LUT4 #(
		.INIT('h153f)
	) name11872 (
		\P2_InstQueue_reg[0][0]/NET0131 ,
		\P2_InstQueue_reg[11][0]/NET0131 ,
		_w1465_,
		_w1460_,
		_w13222_
	);
	LUT4 #(
		.INIT('h153f)
	) name11873 (
		\P2_InstQueue_reg[1][0]/NET0131 ,
		\P2_InstQueue_reg[3][0]/NET0131 ,
		_w1446_,
		_w1457_,
		_w13223_
	);
	LUT4 #(
		.INIT('h153f)
	) name11874 (
		\P2_InstQueue_reg[12][0]/NET0131 ,
		\P2_InstQueue_reg[6][0]/NET0131 ,
		_w1450_,
		_w1452_,
		_w13224_
	);
	LUT4 #(
		.INIT('h135f)
	) name11875 (
		\P2_InstQueue_reg[13][0]/NET0131 ,
		\P2_InstQueue_reg[4][0]/NET0131 ,
		_w1443_,
		_w1462_,
		_w13225_
	);
	LUT4 #(
		.INIT('h8000)
	) name11876 (
		_w13224_,
		_w13225_,
		_w13222_,
		_w13223_,
		_w13226_
	);
	LUT4 #(
		.INIT('h135f)
	) name11877 (
		\P2_InstQueue_reg[2][0]/NET0131 ,
		\P2_InstQueue_reg[9][0]/NET0131 ,
		_w1453_,
		_w1456_,
		_w13227_
	);
	LUT4 #(
		.INIT('h153f)
	) name11878 (
		\P2_InstQueue_reg[7][0]/NET0131 ,
		\P2_InstQueue_reg[8][0]/NET0131 ,
		_w1449_,
		_w1466_,
		_w13228_
	);
	LUT4 #(
		.INIT('h153f)
	) name11879 (
		\P2_InstQueue_reg[14][0]/NET0131 ,
		\P2_InstQueue_reg[15][0]/NET0131 ,
		_w1447_,
		_w1459_,
		_w13229_
	);
	LUT4 #(
		.INIT('h135f)
	) name11880 (
		\P2_InstQueue_reg[10][0]/NET0131 ,
		\P2_InstQueue_reg[5][0]/NET0131 ,
		_w1444_,
		_w1463_,
		_w13230_
	);
	LUT4 #(
		.INIT('h8000)
	) name11881 (
		_w13229_,
		_w13230_,
		_w13227_,
		_w13228_,
		_w13231_
	);
	LUT4 #(
		.INIT('h0111)
	) name11882 (
		_w1592_,
		_w1595_,
		_w13226_,
		_w13231_,
		_w13232_
	);
	LUT3 #(
		.INIT('h80)
	) name11883 (
		_w1549_,
		_w1553_,
		_w13232_,
		_w13233_
	);
	LUT3 #(
		.INIT('h08)
	) name11884 (
		_w1501_,
		_w1568_,
		_w9110_,
		_w13234_
	);
	LUT2 #(
		.INIT('h2)
	) name11885 (
		_w1565_,
		_w9115_,
		_w13235_
	);
	LUT4 #(
		.INIT('h1113)
	) name11886 (
		_w1606_,
		_w13233_,
		_w13234_,
		_w13235_,
		_w13236_
	);
	LUT2 #(
		.INIT('h4)
	) name11887 (
		_w13221_,
		_w13236_,
		_w13237_
	);
	LUT4 #(
		.INIT('hecee)
	) name11888 (
		_w1678_,
		_w13219_,
		_w13220_,
		_w13237_,
		_w13238_
	);
	LUT2 #(
		.INIT('h2)
	) name11889 (
		\P2_EAX_reg[17]/NET0131 ,
		_w7767_,
		_w13239_
	);
	LUT3 #(
		.INIT('h80)
	) name11890 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		_w7777_,
		_w13240_
	);
	LUT4 #(
		.INIT('h6c00)
	) name11891 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		_w7777_,
		_w7789_,
		_w13241_
	);
	LUT2 #(
		.INIT('h2)
	) name11892 (
		_w1565_,
		_w1606_,
		_w13242_
	);
	LUT4 #(
		.INIT('h0013)
	) name11893 (
		_w1604_,
		_w1642_,
		_w7790_,
		_w13242_,
		_w13243_
	);
	LUT2 #(
		.INIT('h8)
	) name11894 (
		_w1606_,
		_w7151_,
		_w13244_
	);
	LUT4 #(
		.INIT('h5054)
	) name11895 (
		\P2_EAX_reg[17]/NET0131 ,
		_w1592_,
		_w1605_,
		_w1601_,
		_w13245_
	);
	LUT4 #(
		.INIT('h0008)
	) name11896 (
		_w1501_,
		_w1568_,
		_w13245_,
		_w13244_,
		_w13246_
	);
	LUT4 #(
		.INIT('h135f)
	) name11897 (
		\P2_InstQueue_reg[13][1]/NET0131 ,
		\P2_InstQueue_reg[3][1]/NET0131 ,
		_w1443_,
		_w1446_,
		_w13247_
	);
	LUT4 #(
		.INIT('h135f)
	) name11898 (
		\P2_InstQueue_reg[7][1]/NET0131 ,
		\P2_InstQueue_reg[9][1]/NET0131 ,
		_w1466_,
		_w1456_,
		_w13248_
	);
	LUT4 #(
		.INIT('h153f)
	) name11899 (
		\P2_InstQueue_reg[12][1]/NET0131 ,
		\P2_InstQueue_reg[6][1]/NET0131 ,
		_w1450_,
		_w1452_,
		_w13249_
	);
	LUT4 #(
		.INIT('h153f)
	) name11900 (
		\P2_InstQueue_reg[11][1]/NET0131 ,
		\P2_InstQueue_reg[5][1]/NET0131 ,
		_w1463_,
		_w1465_,
		_w13250_
	);
	LUT4 #(
		.INIT('h8000)
	) name11901 (
		_w13249_,
		_w13250_,
		_w13247_,
		_w13248_,
		_w13251_
	);
	LUT4 #(
		.INIT('h153f)
	) name11902 (
		\P2_InstQueue_reg[15][1]/NET0131 ,
		\P2_InstQueue_reg[8][1]/NET0131 ,
		_w1449_,
		_w1447_,
		_w13252_
	);
	LUT4 #(
		.INIT('h153f)
	) name11903 (
		\P2_InstQueue_reg[0][1]/NET0131 ,
		\P2_InstQueue_reg[1][1]/NET0131 ,
		_w1457_,
		_w1460_,
		_w13253_
	);
	LUT4 #(
		.INIT('h135f)
	) name11904 (
		\P2_InstQueue_reg[2][1]/NET0131 ,
		\P2_InstQueue_reg[4][1]/NET0131 ,
		_w1453_,
		_w1462_,
		_w13254_
	);
	LUT4 #(
		.INIT('h135f)
	) name11905 (
		\P2_InstQueue_reg[10][1]/NET0131 ,
		\P2_InstQueue_reg[14][1]/NET0131 ,
		_w1444_,
		_w1459_,
		_w13255_
	);
	LUT4 #(
		.INIT('h8000)
	) name11906 (
		_w13254_,
		_w13255_,
		_w13252_,
		_w13253_,
		_w13256_
	);
	LUT4 #(
		.INIT('h0111)
	) name11907 (
		_w1592_,
		_w1595_,
		_w13251_,
		_w13256_,
		_w13257_
	);
	LUT3 #(
		.INIT('h80)
	) name11908 (
		_w1549_,
		_w1553_,
		_w13257_,
		_w13258_
	);
	LUT2 #(
		.INIT('h8)
	) name11909 (
		_w1565_,
		_w10396_,
		_w13259_
	);
	LUT3 #(
		.INIT('h01)
	) name11910 (
		_w13258_,
		_w13246_,
		_w13259_,
		_w13260_
	);
	LUT4 #(
		.INIT('h3100)
	) name11911 (
		\P2_EAX_reg[17]/NET0131 ,
		_w13241_,
		_w13243_,
		_w13260_,
		_w13261_
	);
	LUT3 #(
		.INIT('hce)
	) name11912 (
		_w1678_,
		_w13239_,
		_w13261_,
		_w13262_
	);
	LUT2 #(
		.INIT('h2)
	) name11913 (
		\P2_EAX_reg[18]/NET0131 ,
		_w7767_,
		_w13263_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11914 (
		\P2_EAX_reg[16]/NET0131 ,
		_w7777_,
		_w7778_,
		_w7789_,
		_w13264_
	);
	LUT4 #(
		.INIT('h0013)
	) name11915 (
		_w1604_,
		_w1642_,
		_w7790_,
		_w13264_,
		_w13265_
	);
	LUT2 #(
		.INIT('h8)
	) name11916 (
		_w13240_,
		_w13264_,
		_w13266_
	);
	LUT3 #(
		.INIT('hd1)
	) name11917 (
		\P2_EAX_reg[18]/NET0131 ,
		_w1606_,
		_w5482_,
		_w13267_
	);
	LUT3 #(
		.INIT('h08)
	) name11918 (
		_w1501_,
		_w1568_,
		_w13267_,
		_w13268_
	);
	LUT4 #(
		.INIT('h135f)
	) name11919 (
		\P2_InstQueue_reg[3][2]/NET0131 ,
		\P2_InstQueue_reg[9][2]/NET0131 ,
		_w1446_,
		_w1456_,
		_w13269_
	);
	LUT4 #(
		.INIT('h135f)
	) name11920 (
		\P2_InstQueue_reg[12][2]/NET0131 ,
		\P2_InstQueue_reg[7][2]/NET0131 ,
		_w1452_,
		_w1466_,
		_w13270_
	);
	LUT4 #(
		.INIT('h135f)
	) name11921 (
		\P2_InstQueue_reg[10][2]/NET0131 ,
		\P2_InstQueue_reg[5][2]/NET0131 ,
		_w1444_,
		_w1463_,
		_w13271_
	);
	LUT4 #(
		.INIT('h153f)
	) name11922 (
		\P2_InstQueue_reg[11][2]/NET0131 ,
		\P2_InstQueue_reg[4][2]/NET0131 ,
		_w1462_,
		_w1465_,
		_w13272_
	);
	LUT4 #(
		.INIT('h8000)
	) name11923 (
		_w13271_,
		_w13272_,
		_w13269_,
		_w13270_,
		_w13273_
	);
	LUT4 #(
		.INIT('h153f)
	) name11924 (
		\P2_InstQueue_reg[15][2]/NET0131 ,
		\P2_InstQueue_reg[8][2]/NET0131 ,
		_w1449_,
		_w1447_,
		_w13274_
	);
	LUT4 #(
		.INIT('h153f)
	) name11925 (
		\P2_InstQueue_reg[0][2]/NET0131 ,
		\P2_InstQueue_reg[13][2]/NET0131 ,
		_w1443_,
		_w1460_,
		_w13275_
	);
	LUT4 #(
		.INIT('h153f)
	) name11926 (
		\P2_InstQueue_reg[1][2]/NET0131 ,
		\P2_InstQueue_reg[2][2]/NET0131 ,
		_w1453_,
		_w1457_,
		_w13276_
	);
	LUT4 #(
		.INIT('h153f)
	) name11927 (
		\P2_InstQueue_reg[14][2]/NET0131 ,
		\P2_InstQueue_reg[6][2]/NET0131 ,
		_w1450_,
		_w1459_,
		_w13277_
	);
	LUT4 #(
		.INIT('h8000)
	) name11928 (
		_w13276_,
		_w13277_,
		_w13274_,
		_w13275_,
		_w13278_
	);
	LUT4 #(
		.INIT('h0111)
	) name11929 (
		_w1592_,
		_w1595_,
		_w13273_,
		_w13278_,
		_w13279_
	);
	LUT3 #(
		.INIT('h80)
	) name11930 (
		_w1549_,
		_w1553_,
		_w13279_,
		_w13280_
	);
	LUT3 #(
		.INIT('hd1)
	) name11931 (
		\P2_EAX_reg[18]/NET0131 ,
		_w1606_,
		_w5487_,
		_w13281_
	);
	LUT2 #(
		.INIT('h2)
	) name11932 (
		_w1565_,
		_w13281_,
		_w13282_
	);
	LUT3 #(
		.INIT('h01)
	) name11933 (
		_w13280_,
		_w13282_,
		_w13268_,
		_w13283_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11934 (
		\P2_EAX_reg[18]/NET0131 ,
		_w13265_,
		_w13266_,
		_w13283_,
		_w13284_
	);
	LUT3 #(
		.INIT('hce)
	) name11935 (
		_w1678_,
		_w13263_,
		_w13284_,
		_w13285_
	);
	LUT2 #(
		.INIT('h2)
	) name11936 (
		\P2_EAX_reg[19]/NET0131 ,
		_w7767_,
		_w13286_
	);
	LUT2 #(
		.INIT('h4)
	) name11937 (
		\P2_EAX_reg[19]/NET0131 ,
		_w7789_,
		_w13287_
	);
	LUT2 #(
		.INIT('h8)
	) name11938 (
		_w7779_,
		_w13287_,
		_w13288_
	);
	LUT3 #(
		.INIT('hd1)
	) name11939 (
		\P2_EAX_reg[19]/NET0131 ,
		_w1606_,
		_w3561_,
		_w13289_
	);
	LUT2 #(
		.INIT('h2)
	) name11940 (
		_w1565_,
		_w13289_,
		_w13290_
	);
	LUT4 #(
		.INIT('h135f)
	) name11941 (
		\P2_InstQueue_reg[3][3]/NET0131 ,
		\P2_InstQueue_reg[9][3]/NET0131 ,
		_w1446_,
		_w1456_,
		_w13291_
	);
	LUT4 #(
		.INIT('h135f)
	) name11942 (
		\P2_InstQueue_reg[12][3]/NET0131 ,
		\P2_InstQueue_reg[7][3]/NET0131 ,
		_w1452_,
		_w1466_,
		_w13292_
	);
	LUT4 #(
		.INIT('h135f)
	) name11943 (
		\P2_InstQueue_reg[10][3]/NET0131 ,
		\P2_InstQueue_reg[5][3]/NET0131 ,
		_w1444_,
		_w1463_,
		_w13293_
	);
	LUT4 #(
		.INIT('h153f)
	) name11944 (
		\P2_InstQueue_reg[11][3]/NET0131 ,
		\P2_InstQueue_reg[4][3]/NET0131 ,
		_w1462_,
		_w1465_,
		_w13294_
	);
	LUT4 #(
		.INIT('h8000)
	) name11945 (
		_w13293_,
		_w13294_,
		_w13291_,
		_w13292_,
		_w13295_
	);
	LUT4 #(
		.INIT('h153f)
	) name11946 (
		\P2_InstQueue_reg[15][3]/NET0131 ,
		\P2_InstQueue_reg[8][3]/NET0131 ,
		_w1449_,
		_w1447_,
		_w13296_
	);
	LUT4 #(
		.INIT('h153f)
	) name11947 (
		\P2_InstQueue_reg[0][3]/NET0131 ,
		\P2_InstQueue_reg[13][3]/NET0131 ,
		_w1443_,
		_w1460_,
		_w13297_
	);
	LUT4 #(
		.INIT('h153f)
	) name11948 (
		\P2_InstQueue_reg[1][3]/NET0131 ,
		\P2_InstQueue_reg[2][3]/NET0131 ,
		_w1453_,
		_w1457_,
		_w13298_
	);
	LUT4 #(
		.INIT('h153f)
	) name11949 (
		\P2_InstQueue_reg[14][3]/NET0131 ,
		\P2_InstQueue_reg[6][3]/NET0131 ,
		_w1450_,
		_w1459_,
		_w13299_
	);
	LUT4 #(
		.INIT('h8000)
	) name11950 (
		_w13298_,
		_w13299_,
		_w13296_,
		_w13297_,
		_w13300_
	);
	LUT4 #(
		.INIT('h0111)
	) name11951 (
		_w1592_,
		_w1595_,
		_w13295_,
		_w13300_,
		_w13301_
	);
	LUT3 #(
		.INIT('h80)
	) name11952 (
		_w1549_,
		_w1553_,
		_w13301_,
		_w13302_
	);
	LUT3 #(
		.INIT('hd1)
	) name11953 (
		\P2_EAX_reg[19]/NET0131 ,
		_w1606_,
		_w3556_,
		_w13303_
	);
	LUT3 #(
		.INIT('h08)
	) name11954 (
		_w1501_,
		_w1568_,
		_w13303_,
		_w13304_
	);
	LUT3 #(
		.INIT('h01)
	) name11955 (
		_w13302_,
		_w13304_,
		_w13290_,
		_w13305_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11956 (
		\P2_EAX_reg[19]/NET0131 ,
		_w13265_,
		_w13288_,
		_w13305_,
		_w13306_
	);
	LUT3 #(
		.INIT('hce)
	) name11957 (
		_w1678_,
		_w13286_,
		_w13306_,
		_w13307_
	);
	LUT4 #(
		.INIT('he0c0)
	) name11958 (
		_w1604_,
		_w1642_,
		_w1678_,
		_w7790_,
		_w13308_
	);
	LUT3 #(
		.INIT('ha2)
	) name11959 (
		\P2_EAX_reg[20]/NET0131 ,
		_w7767_,
		_w13308_,
		_w13309_
	);
	LUT4 #(
		.INIT('h8a88)
	) name11960 (
		\P2_EAX_reg[20]/NET0131 ,
		_w1607_,
		_w7780_,
		_w7789_,
		_w13310_
	);
	LUT3 #(
		.INIT('h40)
	) name11961 (
		\P2_EAX_reg[20]/NET0131 ,
		_w7780_,
		_w7789_,
		_w13311_
	);
	LUT4 #(
		.INIT('h153f)
	) name11962 (
		\P2_InstQueue_reg[1][4]/NET0131 ,
		\P2_InstQueue_reg[7][4]/NET0131 ,
		_w1466_,
		_w1457_,
		_w13312_
	);
	LUT4 #(
		.INIT('h135f)
	) name11963 (
		\P2_InstQueue_reg[11][4]/NET0131 ,
		\P2_InstQueue_reg[14][4]/NET0131 ,
		_w1465_,
		_w1459_,
		_w13313_
	);
	LUT4 #(
		.INIT('h135f)
	) name11964 (
		\P2_InstQueue_reg[10][4]/NET0131 ,
		\P2_InstQueue_reg[4][4]/NET0131 ,
		_w1444_,
		_w1462_,
		_w13314_
	);
	LUT4 #(
		.INIT('h135f)
	) name11965 (
		\P2_InstQueue_reg[13][4]/NET0131 ,
		\P2_InstQueue_reg[9][4]/NET0131 ,
		_w1443_,
		_w1456_,
		_w13315_
	);
	LUT4 #(
		.INIT('h8000)
	) name11966 (
		_w13314_,
		_w13315_,
		_w13312_,
		_w13313_,
		_w13316_
	);
	LUT4 #(
		.INIT('h153f)
	) name11967 (
		\P2_InstQueue_reg[2][4]/NET0131 ,
		\P2_InstQueue_reg[8][4]/NET0131 ,
		_w1449_,
		_w1453_,
		_w13317_
	);
	LUT4 #(
		.INIT('h135f)
	) name11968 (
		\P2_InstQueue_reg[3][4]/NET0131 ,
		\P2_InstQueue_reg[5][4]/NET0131 ,
		_w1446_,
		_w1463_,
		_w13318_
	);
	LUT4 #(
		.INIT('h135f)
	) name11969 (
		\P2_InstQueue_reg[12][4]/NET0131 ,
		\P2_InstQueue_reg[15][4]/NET0131 ,
		_w1452_,
		_w1447_,
		_w13319_
	);
	LUT4 #(
		.INIT('h153f)
	) name11970 (
		\P2_InstQueue_reg[0][4]/NET0131 ,
		\P2_InstQueue_reg[6][4]/NET0131 ,
		_w1450_,
		_w1460_,
		_w13320_
	);
	LUT4 #(
		.INIT('h8000)
	) name11971 (
		_w13319_,
		_w13320_,
		_w13317_,
		_w13318_,
		_w13321_
	);
	LUT4 #(
		.INIT('h0111)
	) name11972 (
		_w1592_,
		_w1595_,
		_w13316_,
		_w13321_,
		_w13322_
	);
	LUT3 #(
		.INIT('h80)
	) name11973 (
		_w1549_,
		_w1553_,
		_w13322_,
		_w13323_
	);
	LUT3 #(
		.INIT('h08)
	) name11974 (
		_w1501_,
		_w1568_,
		_w2267_,
		_w13324_
	);
	LUT2 #(
		.INIT('h2)
	) name11975 (
		_w1565_,
		_w2276_,
		_w13325_
	);
	LUT4 #(
		.INIT('h1113)
	) name11976 (
		_w1606_,
		_w13323_,
		_w13324_,
		_w13325_,
		_w13326_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name11977 (
		_w1678_,
		_w13310_,
		_w13311_,
		_w13326_,
		_w13327_
	);
	LUT2 #(
		.INIT('he)
	) name11978 (
		_w13309_,
		_w13327_,
		_w13328_
	);
	LUT2 #(
		.INIT('h2)
	) name11979 (
		\P2_EAX_reg[21]/NET0131 ,
		_w7767_,
		_w13329_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11980 (
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[21]/NET0131 ,
		_w7780_,
		_w7789_,
		_w13330_
	);
	LUT4 #(
		.INIT('h6c00)
	) name11981 (
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[21]/NET0131 ,
		_w7780_,
		_w7789_,
		_w13331_
	);
	LUT2 #(
		.INIT('h2)
	) name11982 (
		_w1565_,
		_w6502_,
		_w13332_
	);
	LUT3 #(
		.INIT('h08)
	) name11983 (
		_w1501_,
		_w1568_,
		_w6497_,
		_w13333_
	);
	LUT4 #(
		.INIT('h135f)
	) name11984 (
		\P2_InstQueue_reg[5][5]/NET0131 ,
		\P2_InstQueue_reg[9][5]/NET0131 ,
		_w1463_,
		_w1456_,
		_w13334_
	);
	LUT4 #(
		.INIT('h135f)
	) name11985 (
		\P2_InstQueue_reg[12][5]/NET0131 ,
		\P2_InstQueue_reg[7][5]/NET0131 ,
		_w1452_,
		_w1466_,
		_w13335_
	);
	LUT4 #(
		.INIT('h153f)
	) name11986 (
		\P2_InstQueue_reg[10][5]/NET0131 ,
		\P2_InstQueue_reg[8][5]/NET0131 ,
		_w1449_,
		_w1444_,
		_w13336_
	);
	LUT4 #(
		.INIT('h153f)
	) name11987 (
		\P2_InstQueue_reg[14][5]/NET0131 ,
		\P2_InstQueue_reg[4][5]/NET0131 ,
		_w1462_,
		_w1459_,
		_w13337_
	);
	LUT4 #(
		.INIT('h8000)
	) name11988 (
		_w13336_,
		_w13337_,
		_w13334_,
		_w13335_,
		_w13338_
	);
	LUT4 #(
		.INIT('h153f)
	) name11989 (
		\P2_InstQueue_reg[15][5]/NET0131 ,
		\P2_InstQueue_reg[3][5]/NET0131 ,
		_w1446_,
		_w1447_,
		_w13339_
	);
	LUT4 #(
		.INIT('h153f)
	) name11990 (
		\P2_InstQueue_reg[0][5]/NET0131 ,
		\P2_InstQueue_reg[13][5]/NET0131 ,
		_w1443_,
		_w1460_,
		_w13340_
	);
	LUT4 #(
		.INIT('h153f)
	) name11991 (
		\P2_InstQueue_reg[11][5]/NET0131 ,
		\P2_InstQueue_reg[2][5]/NET0131 ,
		_w1453_,
		_w1465_,
		_w13341_
	);
	LUT4 #(
		.INIT('h153f)
	) name11992 (
		\P2_InstQueue_reg[1][5]/NET0131 ,
		\P2_InstQueue_reg[6][5]/NET0131 ,
		_w1450_,
		_w1457_,
		_w13342_
	);
	LUT4 #(
		.INIT('h8000)
	) name11993 (
		_w13341_,
		_w13342_,
		_w13339_,
		_w13340_,
		_w13343_
	);
	LUT4 #(
		.INIT('h0111)
	) name11994 (
		_w1592_,
		_w1595_,
		_w13338_,
		_w13343_,
		_w13344_
	);
	LUT3 #(
		.INIT('h80)
	) name11995 (
		_w1549_,
		_w1553_,
		_w13344_,
		_w13345_
	);
	LUT4 #(
		.INIT('h0057)
	) name11996 (
		_w1606_,
		_w13332_,
		_w13333_,
		_w13345_,
		_w13346_
	);
	LUT4 #(
		.INIT('h0d00)
	) name11997 (
		\P2_EAX_reg[21]/NET0131 ,
		_w7792_,
		_w13331_,
		_w13346_,
		_w13347_
	);
	LUT3 #(
		.INIT('hce)
	) name11998 (
		_w1678_,
		_w13329_,
		_w13347_,
		_w13348_
	);
	LUT2 #(
		.INIT('h2)
	) name11999 (
		\P2_EAX_reg[22]/NET0131 ,
		_w7767_,
		_w13349_
	);
	LUT3 #(
		.INIT('ha2)
	) name12000 (
		\P2_EAX_reg[22]/NET0131 ,
		_w7792_,
		_w13330_,
		_w13350_
	);
	LUT2 #(
		.INIT('h4)
	) name12001 (
		\P2_EAX_reg[22]/NET0131 ,
		_w7789_,
		_w13351_
	);
	LUT4 #(
		.INIT('h8000)
	) name12002 (
		\P2_EAX_reg[20]/NET0131 ,
		\P2_EAX_reg[21]/NET0131 ,
		_w7780_,
		_w13351_,
		_w13352_
	);
	LUT4 #(
		.INIT('h135f)
	) name12003 (
		\P2_InstQueue_reg[2][6]/NET0131 ,
		\P2_InstQueue_reg[5][6]/NET0131 ,
		_w1453_,
		_w1463_,
		_w13353_
	);
	LUT4 #(
		.INIT('h153f)
	) name12004 (
		\P2_InstQueue_reg[0][6]/NET0131 ,
		\P2_InstQueue_reg[13][6]/NET0131 ,
		_w1443_,
		_w1460_,
		_w13354_
	);
	LUT4 #(
		.INIT('h153f)
	) name12005 (
		\P2_InstQueue_reg[12][6]/NET0131 ,
		\P2_InstQueue_reg[6][6]/NET0131 ,
		_w1450_,
		_w1452_,
		_w13355_
	);
	LUT4 #(
		.INIT('h153f)
	) name12006 (
		\P2_InstQueue_reg[1][6]/NET0131 ,
		\P2_InstQueue_reg[3][6]/NET0131 ,
		_w1446_,
		_w1457_,
		_w13356_
	);
	LUT4 #(
		.INIT('h8000)
	) name12007 (
		_w13355_,
		_w13356_,
		_w13353_,
		_w13354_,
		_w13357_
	);
	LUT4 #(
		.INIT('h153f)
	) name12008 (
		\P2_InstQueue_reg[11][6]/NET0131 ,
		\P2_InstQueue_reg[15][6]/NET0131 ,
		_w1447_,
		_w1465_,
		_w13358_
	);
	LUT4 #(
		.INIT('h153f)
	) name12009 (
		\P2_InstQueue_reg[14][6]/NET0131 ,
		\P2_InstQueue_reg[9][6]/NET0131 ,
		_w1456_,
		_w1459_,
		_w13359_
	);
	LUT4 #(
		.INIT('h153f)
	) name12010 (
		\P2_InstQueue_reg[4][6]/NET0131 ,
		\P2_InstQueue_reg[8][6]/NET0131 ,
		_w1449_,
		_w1462_,
		_w13360_
	);
	LUT4 #(
		.INIT('h135f)
	) name12011 (
		\P2_InstQueue_reg[10][6]/NET0131 ,
		\P2_InstQueue_reg[7][6]/NET0131 ,
		_w1444_,
		_w1466_,
		_w13361_
	);
	LUT4 #(
		.INIT('h8000)
	) name12012 (
		_w13360_,
		_w13361_,
		_w13358_,
		_w13359_,
		_w13362_
	);
	LUT4 #(
		.INIT('h0111)
	) name12013 (
		_w1592_,
		_w1595_,
		_w13357_,
		_w13362_,
		_w13363_
	);
	LUT3 #(
		.INIT('h80)
	) name12014 (
		_w1549_,
		_w1553_,
		_w13363_,
		_w13364_
	);
	LUT2 #(
		.INIT('h2)
	) name12015 (
		_w1565_,
		_w4977_,
		_w13365_
	);
	LUT3 #(
		.INIT('h08)
	) name12016 (
		_w1501_,
		_w1568_,
		_w4972_,
		_w13366_
	);
	LUT4 #(
		.INIT('h1113)
	) name12017 (
		_w1606_,
		_w13364_,
		_w13365_,
		_w13366_,
		_w13367_
	);
	LUT2 #(
		.INIT('h4)
	) name12018 (
		_w13352_,
		_w13367_,
		_w13368_
	);
	LUT4 #(
		.INIT('hecee)
	) name12019 (
		_w1678_,
		_w13349_,
		_w13350_,
		_w13368_,
		_w13369_
	);
	LUT2 #(
		.INIT('h2)
	) name12020 (
		\P2_EAX_reg[23]/NET0131 ,
		_w7767_,
		_w13370_
	);
	LUT3 #(
		.INIT('h60)
	) name12021 (
		\P2_EAX_reg[23]/NET0131 ,
		_w7782_,
		_w7789_,
		_w13371_
	);
	LUT3 #(
		.INIT('h08)
	) name12022 (
		_w1501_,
		_w1568_,
		_w2305_,
		_w13372_
	);
	LUT2 #(
		.INIT('h2)
	) name12023 (
		_w1565_,
		_w2295_,
		_w13373_
	);
	LUT4 #(
		.INIT('h7888)
	) name12024 (
		_w7799_,
		_w7804_,
		_w7809_,
		_w7814_,
		_w13374_
	);
	LUT2 #(
		.INIT('h8)
	) name12025 (
		_w1596_,
		_w13374_,
		_w13375_
	);
	LUT3 #(
		.INIT('h80)
	) name12026 (
		_w1549_,
		_w1553_,
		_w13375_,
		_w13376_
	);
	LUT4 #(
		.INIT('h0057)
	) name12027 (
		_w1606_,
		_w13372_,
		_w13373_,
		_w13376_,
		_w13377_
	);
	LUT3 #(
		.INIT('hd0)
	) name12028 (
		\P2_EAX_reg[23]/NET0131 ,
		_w7792_,
		_w13377_,
		_w13378_
	);
	LUT4 #(
		.INIT('hecee)
	) name12029 (
		_w1678_,
		_w13370_,
		_w13371_,
		_w13378_,
		_w13379_
	);
	LUT3 #(
		.INIT('ha2)
	) name12030 (
		\P2_EAX_reg[24]/NET0131 ,
		_w7767_,
		_w13308_,
		_w13380_
	);
	LUT3 #(
		.INIT('h48)
	) name12031 (
		\P2_EAX_reg[24]/NET0131 ,
		_w7789_,
		_w12546_,
		_w13381_
	);
	LUT3 #(
		.INIT('h54)
	) name12032 (
		_w1605_,
		_w9105_,
		_w9106_,
		_w13382_
	);
	LUT3 #(
		.INIT('h80)
	) name12033 (
		_w1501_,
		_w1568_,
		_w13382_,
		_w13383_
	);
	LUT3 #(
		.INIT('h54)
	) name12034 (
		_w1602_,
		_w10007_,
		_w13383_,
		_w13384_
	);
	LUT3 #(
		.INIT('h82)
	) name12035 (
		_w1596_,
		_w7815_,
		_w7826_,
		_w13385_
	);
	LUT3 #(
		.INIT('h80)
	) name12036 (
		_w1549_,
		_w1553_,
		_w13385_,
		_w13386_
	);
	LUT3 #(
		.INIT('h07)
	) name12037 (
		\P2_EAX_reg[24]/NET0131 ,
		_w1607_,
		_w13386_,
		_w13387_
	);
	LUT2 #(
		.INIT('h4)
	) name12038 (
		_w13384_,
		_w13387_,
		_w13388_
	);
	LUT4 #(
		.INIT('hecee)
	) name12039 (
		_w1678_,
		_w13380_,
		_w13381_,
		_w13388_,
		_w13389_
	);
	LUT3 #(
		.INIT('ha2)
	) name12040 (
		\P2_EAX_reg[28]/NET0131 ,
		_w7767_,
		_w13308_,
		_w13390_
	);
	LUT4 #(
		.INIT('h6a00)
	) name12041 (
		\P2_EAX_reg[28]/NET0131 ,
		_w7784_,
		_w7785_,
		_w7789_,
		_w13391_
	);
	LUT4 #(
		.INIT('h08a2)
	) name12042 (
		_w1596_,
		_w7850_,
		_w7861_,
		_w7872_,
		_w13392_
	);
	LUT2 #(
		.INIT('h8)
	) name12043 (
		_w1554_,
		_w13392_,
		_w13393_
	);
	LUT2 #(
		.INIT('h8)
	) name12044 (
		\P2_EAX_reg[28]/NET0131 ,
		_w1607_,
		_w13394_
	);
	LUT3 #(
		.INIT('h54)
	) name12045 (
		_w1605_,
		_w2261_,
		_w2262_,
		_w13395_
	);
	LUT3 #(
		.INIT('h80)
	) name12046 (
		_w1501_,
		_w1568_,
		_w13395_,
		_w13396_
	);
	LUT3 #(
		.INIT('h54)
	) name12047 (
		_w1602_,
		_w9452_,
		_w13396_,
		_w13397_
	);
	LUT3 #(
		.INIT('h01)
	) name12048 (
		_w13394_,
		_w13393_,
		_w13397_,
		_w13398_
	);
	LUT4 #(
		.INIT('hecee)
	) name12049 (
		_w1678_,
		_w13390_,
		_w13391_,
		_w13398_,
		_w13399_
	);
	LUT2 #(
		.INIT('h2)
	) name12050 (
		_w1867_,
		_w3471_,
		_w13400_
	);
	LUT4 #(
		.INIT('hec00)
	) name12051 (
		_w1725_,
		_w1795_,
		_w1802_,
		_w13400_,
		_w13401_
	);
	LUT4 #(
		.INIT('h0111)
	) name12052 (
		_w1842_,
		_w1845_,
		_w3162_,
		_w3167_,
		_w13402_
	);
	LUT4 #(
		.INIT('h4000)
	) name12053 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13402_,
		_w13403_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12054 (
		_w1933_,
		_w10601_,
		_w13403_,
		_w13401_,
		_w13404_
	);
	LUT3 #(
		.INIT('hf2)
	) name12055 (
		\P1_EAX_reg[0]/NET0131 ,
		_w10016_,
		_w13404_,
		_w13405_
	);
	LUT3 #(
		.INIT('h80)
	) name12056 (
		_w1750_,
		_w1813_,
		_w12514_,
		_w13406_
	);
	LUT4 #(
		.INIT('h0057)
	) name12057 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1863_,
		_w8992_,
		_w13406_,
		_w13407_
	);
	LUT4 #(
		.INIT('hb700)
	) name12058 (
		\P1_EBX_reg[25]/NET0131 ,
		_w1829_,
		_w8987_,
		_w13407_,
		_w13408_
	);
	LUT2 #(
		.INIT('h2)
	) name12059 (
		\P1_EBX_reg[25]/NET0131 ,
		_w9102_,
		_w13409_
	);
	LUT3 #(
		.INIT('hf2)
	) name12060 (
		_w1933_,
		_w13408_,
		_w13409_,
		_w13410_
	);
	LUT2 #(
		.INIT('h2)
	) name12061 (
		\P2_EBX_reg[25]/NET0131 ,
		_w7767_,
		_w13411_
	);
	LUT4 #(
		.INIT('hb030)
	) name12062 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1578_,
		_w8961_,
		_w8957_,
		_w13412_
	);
	LUT3 #(
		.INIT('h80)
	) name12063 (
		_w1503_,
		_w1549_,
		_w12551_,
		_w13413_
	);
	LUT2 #(
		.INIT('h4)
	) name12064 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1578_,
		_w13414_
	);
	LUT4 #(
		.INIT('h070f)
	) name12065 (
		\P2_EBX_reg[24]/NET0131 ,
		_w8957_,
		_w13413_,
		_w13414_,
		_w13415_
	);
	LUT4 #(
		.INIT('h08cc)
	) name12066 (
		\P2_EBX_reg[25]/NET0131 ,
		_w1678_,
		_w13412_,
		_w13415_,
		_w13416_
	);
	LUT2 #(
		.INIT('he)
	) name12067 (
		_w13411_,
		_w13416_,
		_w13417_
	);
	LUT4 #(
		.INIT('h2f00)
	) name12068 (
		\P2_Flush_reg/NET0131 ,
		_w1658_,
		_w1662_,
		_w1678_,
		_w13418_
	);
	LUT2 #(
		.INIT('h2)
	) name12069 (
		\P2_Flush_reg/NET0131 ,
		_w7767_,
		_w13419_
	);
	LUT2 #(
		.INIT('he)
	) name12070 (
		_w13418_,
		_w13419_,
		_w13420_
	);
	LUT4 #(
		.INIT('h2f00)
	) name12071 (
		\P1_Flush_reg/NET0131 ,
		_w1922_,
		_w1925_,
		_w1933_,
		_w13421_
	);
	LUT2 #(
		.INIT('h2)
	) name12072 (
		\P1_Flush_reg/NET0131 ,
		_w9102_,
		_w13422_
	);
	LUT2 #(
		.INIT('he)
	) name12073 (
		_w13421_,
		_w13422_,
		_w13423_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name12074 (
		_w1945_,
		_w2170_,
		_w2174_,
		_w2176_,
		_w13424_
	);
	LUT2 #(
		.INIT('h2)
	) name12075 (
		\P3_More_reg/NET0131 ,
		_w8341_,
		_w13425_
	);
	LUT2 #(
		.INIT('he)
	) name12076 (
		_w13424_,
		_w13425_,
		_w13426_
	);
	LUT3 #(
		.INIT('ha2)
	) name12077 (
		\P3_uWord_reg[11]/NET0131 ,
		_w8341_,
		_w9529_,
		_w13427_
	);
	LUT4 #(
		.INIT('h5551)
	) name12078 (
		_w8440_,
		_w9543_,
		_w9542_,
		_w12841_,
		_w13428_
	);
	LUT3 #(
		.INIT('hce)
	) name12079 (
		_w1945_,
		_w13427_,
		_w13428_,
		_w13429_
	);
	LUT4 #(
		.INIT('h40c0)
	) name12080 (
		\P1_EAX_reg[16]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9426_,
		_w13430_
	);
	LUT4 #(
		.INIT('h4080)
	) name12081 (
		\P1_EAX_reg[16]/NET0131 ,
		_w1804_,
		_w1826_,
		_w9426_,
		_w13431_
	);
	LUT2 #(
		.INIT('h2)
	) name12082 (
		_w1795_,
		_w3471_,
		_w13432_
	);
	LUT3 #(
		.INIT('h08)
	) name12083 (
		_w1725_,
		_w1802_,
		_w3500_,
		_w13433_
	);
	LUT4 #(
		.INIT('h135f)
	) name12084 (
		\P1_InstQueue_reg[15][0]/NET0131 ,
		\P1_InstQueue_reg[3][0]/NET0131 ,
		_w1698_,
		_w1688_,
		_w13434_
	);
	LUT4 #(
		.INIT('h153f)
	) name12085 (
		\P1_InstQueue_reg[5][0]/NET0131 ,
		\P1_InstQueue_reg[7][0]/NET0131 ,
		_w1689_,
		_w1709_,
		_w13435_
	);
	LUT4 #(
		.INIT('h135f)
	) name12086 (
		\P1_InstQueue_reg[11][0]/NET0131 ,
		\P1_InstQueue_reg[2][0]/NET0131 ,
		_w1712_,
		_w1706_,
		_w13436_
	);
	LUT4 #(
		.INIT('h135f)
	) name12087 (
		\P1_InstQueue_reg[4][0]/NET0131 ,
		\P1_InstQueue_reg[6][0]/NET0131 ,
		_w1692_,
		_w1702_,
		_w13437_
	);
	LUT4 #(
		.INIT('h8000)
	) name12088 (
		_w13436_,
		_w13437_,
		_w13434_,
		_w13435_,
		_w13438_
	);
	LUT4 #(
		.INIT('h153f)
	) name12089 (
		\P1_InstQueue_reg[12][0]/NET0131 ,
		\P1_InstQueue_reg[14][0]/NET0131 ,
		_w1696_,
		_w1703_,
		_w13439_
	);
	LUT4 #(
		.INIT('h153f)
	) name12090 (
		\P1_InstQueue_reg[10][0]/NET0131 ,
		\P1_InstQueue_reg[8][0]/NET0131 ,
		_w1691_,
		_w1708_,
		_w13440_
	);
	LUT4 #(
		.INIT('h135f)
	) name12091 (
		\P1_InstQueue_reg[13][0]/NET0131 ,
		\P1_InstQueue_reg[9][0]/NET0131 ,
		_w1694_,
		_w1711_,
		_w13441_
	);
	LUT4 #(
		.INIT('h153f)
	) name12092 (
		\P1_InstQueue_reg[0][0]/NET0131 ,
		\P1_InstQueue_reg[1][0]/NET0131 ,
		_w1699_,
		_w1705_,
		_w13442_
	);
	LUT4 #(
		.INIT('h8000)
	) name12093 (
		_w13441_,
		_w13442_,
		_w13439_,
		_w13440_,
		_w13443_
	);
	LUT4 #(
		.INIT('h0111)
	) name12094 (
		_w1842_,
		_w1845_,
		_w13438_,
		_w13443_,
		_w13444_
	);
	LUT4 #(
		.INIT('h4000)
	) name12095 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13444_,
		_w13445_
	);
	LUT4 #(
		.INIT('h0057)
	) name12096 (
		_w1867_,
		_w13432_,
		_w13433_,
		_w13445_,
		_w13446_
	);
	LUT4 #(
		.INIT('h7500)
	) name12097 (
		\P1_EAX_reg[16]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13446_,
		_w13447_
	);
	LUT2 #(
		.INIT('h2)
	) name12098 (
		\P1_EAX_reg[16]/NET0131 ,
		_w9102_,
		_w13448_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12099 (
		_w1933_,
		_w13431_,
		_w13447_,
		_w13448_,
		_w13449_
	);
	LUT2 #(
		.INIT('h2)
	) name12100 (
		\P1_EAX_reg[17]/NET0131 ,
		_w9102_,
		_w13450_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12101 (
		\P1_EAX_reg[17]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13430_,
		_w13451_
	);
	LUT3 #(
		.INIT('h40)
	) name12102 (
		\P1_EAX_reg[17]/NET0131 ,
		_w1804_,
		_w1826_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name12103 (
		_w9427_,
		_w13452_,
		_w13453_
	);
	LUT4 #(
		.INIT('h153f)
	) name12104 (
		\P1_InstQueue_reg[10][1]/NET0131 ,
		\P1_InstQueue_reg[3][1]/NET0131 ,
		_w1688_,
		_w1708_,
		_w13454_
	);
	LUT4 #(
		.INIT('h135f)
	) name12105 (
		\P1_InstQueue_reg[15][1]/NET0131 ,
		\P1_InstQueue_reg[8][1]/NET0131 ,
		_w1698_,
		_w1691_,
		_w13455_
	);
	LUT4 #(
		.INIT('h135f)
	) name12106 (
		\P1_InstQueue_reg[11][1]/NET0131 ,
		\P1_InstQueue_reg[2][1]/NET0131 ,
		_w1712_,
		_w1706_,
		_w13456_
	);
	LUT4 #(
		.INIT('h135f)
	) name12107 (
		\P1_InstQueue_reg[4][1]/NET0131 ,
		\P1_InstQueue_reg[6][1]/NET0131 ,
		_w1692_,
		_w1702_,
		_w13457_
	);
	LUT4 #(
		.INIT('h8000)
	) name12108 (
		_w13456_,
		_w13457_,
		_w13454_,
		_w13455_,
		_w13458_
	);
	LUT4 #(
		.INIT('h153f)
	) name12109 (
		\P1_InstQueue_reg[12][1]/NET0131 ,
		\P1_InstQueue_reg[14][1]/NET0131 ,
		_w1696_,
		_w1703_,
		_w13459_
	);
	LUT4 #(
		.INIT('h135f)
	) name12110 (
		\P1_InstQueue_reg[5][1]/NET0131 ,
		\P1_InstQueue_reg[9][1]/NET0131 ,
		_w1709_,
		_w1711_,
		_w13460_
	);
	LUT4 #(
		.INIT('h135f)
	) name12111 (
		\P1_InstQueue_reg[13][1]/NET0131 ,
		\P1_InstQueue_reg[7][1]/NET0131 ,
		_w1694_,
		_w1689_,
		_w13461_
	);
	LUT4 #(
		.INIT('h153f)
	) name12112 (
		\P1_InstQueue_reg[0][1]/NET0131 ,
		\P1_InstQueue_reg[1][1]/NET0131 ,
		_w1699_,
		_w1705_,
		_w13462_
	);
	LUT4 #(
		.INIT('h8000)
	) name12113 (
		_w13461_,
		_w13462_,
		_w13459_,
		_w13460_,
		_w13463_
	);
	LUT4 #(
		.INIT('h0111)
	) name12114 (
		_w1842_,
		_w1845_,
		_w13458_,
		_w13463_,
		_w13464_
	);
	LUT4 #(
		.INIT('h4000)
	) name12115 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13464_,
		_w13465_
	);
	LUT3 #(
		.INIT('h08)
	) name12116 (
		_w1725_,
		_w1802_,
		_w3493_,
		_w13466_
	);
	LUT2 #(
		.INIT('h2)
	) name12117 (
		_w1795_,
		_w3478_,
		_w13467_
	);
	LUT4 #(
		.INIT('h1113)
	) name12118 (
		_w1867_,
		_w13465_,
		_w13466_,
		_w13467_,
		_w13468_
	);
	LUT2 #(
		.INIT('h4)
	) name12119 (
		_w13453_,
		_w13468_,
		_w13469_
	);
	LUT4 #(
		.INIT('hecee)
	) name12120 (
		_w1933_,
		_w13450_,
		_w13451_,
		_w13469_,
		_w13470_
	);
	LUT2 #(
		.INIT('h2)
	) name12121 (
		\P1_More_reg/NET0131 ,
		_w9102_,
		_w13471_
	);
	LUT4 #(
		.INIT('hffb0)
	) name12122 (
		_w1912_,
		_w1918_,
		_w1933_,
		_w13471_,
		_w13472_
	);
	LUT2 #(
		.INIT('h2)
	) name12123 (
		\P1_EAX_reg[19]/NET0131 ,
		_w9102_,
		_w13473_
	);
	LUT2 #(
		.INIT('h2)
	) name12124 (
		_w1827_,
		_w9429_,
		_w13474_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12125 (
		\P1_EAX_reg[19]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13474_,
		_w13475_
	);
	LUT3 #(
		.INIT('h40)
	) name12126 (
		\P1_EAX_reg[19]/NET0131 ,
		_w1804_,
		_w1826_,
		_w13476_
	);
	LUT2 #(
		.INIT('h8)
	) name12127 (
		_w9429_,
		_w13476_,
		_w13477_
	);
	LUT4 #(
		.INIT('h153f)
	) name12128 (
		\P1_InstQueue_reg[10][3]/NET0131 ,
		\P1_InstQueue_reg[3][3]/NET0131 ,
		_w1688_,
		_w1708_,
		_w13478_
	);
	LUT4 #(
		.INIT('h135f)
	) name12129 (
		\P1_InstQueue_reg[5][3]/NET0131 ,
		\P1_InstQueue_reg[6][3]/NET0131 ,
		_w1709_,
		_w1702_,
		_w13479_
	);
	LUT4 #(
		.INIT('h153f)
	) name12130 (
		\P1_InstQueue_reg[2][3]/NET0131 ,
		\P1_InstQueue_reg[4][3]/NET0131 ,
		_w1692_,
		_w1706_,
		_w13480_
	);
	LUT4 #(
		.INIT('h153f)
	) name12131 (
		\P1_InstQueue_reg[11][3]/NET0131 ,
		\P1_InstQueue_reg[15][3]/NET0131 ,
		_w1698_,
		_w1712_,
		_w13481_
	);
	LUT4 #(
		.INIT('h8000)
	) name12132 (
		_w13480_,
		_w13481_,
		_w13478_,
		_w13479_,
		_w13482_
	);
	LUT4 #(
		.INIT('h153f)
	) name12133 (
		\P1_InstQueue_reg[12][3]/NET0131 ,
		\P1_InstQueue_reg[13][3]/NET0131 ,
		_w1694_,
		_w1703_,
		_w13483_
	);
	LUT4 #(
		.INIT('h135f)
	) name12134 (
		\P1_InstQueue_reg[8][3]/NET0131 ,
		\P1_InstQueue_reg[9][3]/NET0131 ,
		_w1691_,
		_w1711_,
		_w13484_
	);
	LUT4 #(
		.INIT('h135f)
	) name12135 (
		\P1_InstQueue_reg[14][3]/NET0131 ,
		\P1_InstQueue_reg[7][3]/NET0131 ,
		_w1696_,
		_w1689_,
		_w13485_
	);
	LUT4 #(
		.INIT('h153f)
	) name12136 (
		\P1_InstQueue_reg[0][3]/NET0131 ,
		\P1_InstQueue_reg[1][3]/NET0131 ,
		_w1699_,
		_w1705_,
		_w13486_
	);
	LUT4 #(
		.INIT('h8000)
	) name12137 (
		_w13485_,
		_w13486_,
		_w13483_,
		_w13484_,
		_w13487_
	);
	LUT4 #(
		.INIT('h0111)
	) name12138 (
		_w1842_,
		_w1845_,
		_w13482_,
		_w13487_,
		_w13488_
	);
	LUT4 #(
		.INIT('h4000)
	) name12139 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13488_,
		_w13489_
	);
	LUT3 #(
		.INIT('h08)
	) name12140 (
		_w1725_,
		_w1802_,
		_w3486_,
		_w13490_
	);
	LUT2 #(
		.INIT('h2)
	) name12141 (
		_w1795_,
		_w3428_,
		_w13491_
	);
	LUT4 #(
		.INIT('h1113)
	) name12142 (
		_w1867_,
		_w13489_,
		_w13490_,
		_w13491_,
		_w13492_
	);
	LUT2 #(
		.INIT('h4)
	) name12143 (
		_w13477_,
		_w13492_,
		_w13493_
	);
	LUT4 #(
		.INIT('hecee)
	) name12144 (
		_w1933_,
		_w13473_,
		_w13475_,
		_w13493_,
		_w13494_
	);
	LUT2 #(
		.INIT('h2)
	) name12145 (
		\P1_EAX_reg[18]/NET0131 ,
		_w9102_,
		_w13495_
	);
	LUT4 #(
		.INIT('haa8a)
	) name12146 (
		\P1_EAX_reg[18]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13474_,
		_w13496_
	);
	LUT3 #(
		.INIT('h80)
	) name12147 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		_w9426_,
		_w13497_
	);
	LUT3 #(
		.INIT('h20)
	) name12148 (
		_w1827_,
		_w9429_,
		_w13497_,
		_w13498_
	);
	LUT4 #(
		.INIT('h135f)
	) name12149 (
		\P1_InstQueue_reg[14][2]/NET0131 ,
		\P1_InstQueue_reg[1][2]/NET0131 ,
		_w1696_,
		_w1699_,
		_w13499_
	);
	LUT4 #(
		.INIT('h153f)
	) name12150 (
		\P1_InstQueue_reg[4][2]/NET0131 ,
		\P1_InstQueue_reg[8][2]/NET0131 ,
		_w1691_,
		_w1692_,
		_w13500_
	);
	LUT4 #(
		.INIT('h135f)
	) name12151 (
		\P1_InstQueue_reg[11][2]/NET0131 ,
		\P1_InstQueue_reg[6][2]/NET0131 ,
		_w1712_,
		_w1702_,
		_w13501_
	);
	LUT4 #(
		.INIT('h153f)
	) name12152 (
		\P1_InstQueue_reg[0][2]/NET0131 ,
		\P1_InstQueue_reg[3][2]/NET0131 ,
		_w1688_,
		_w1705_,
		_w13502_
	);
	LUT4 #(
		.INIT('h8000)
	) name12153 (
		_w13501_,
		_w13502_,
		_w13499_,
		_w13500_,
		_w13503_
	);
	LUT4 #(
		.INIT('h135f)
	) name12154 (
		\P1_InstQueue_reg[13][2]/NET0131 ,
		\P1_InstQueue_reg[9][2]/NET0131 ,
		_w1694_,
		_w1711_,
		_w13504_
	);
	LUT4 #(
		.INIT('h153f)
	) name12155 (
		\P1_InstQueue_reg[5][2]/NET0131 ,
		\P1_InstQueue_reg[7][2]/NET0131 ,
		_w1689_,
		_w1709_,
		_w13505_
	);
	LUT4 #(
		.INIT('h153f)
	) name12156 (
		\P1_InstQueue_reg[12][2]/NET0131 ,
		\P1_InstQueue_reg[15][2]/NET0131 ,
		_w1698_,
		_w1703_,
		_w13506_
	);
	LUT4 #(
		.INIT('h135f)
	) name12157 (
		\P1_InstQueue_reg[10][2]/NET0131 ,
		\P1_InstQueue_reg[2][2]/NET0131 ,
		_w1708_,
		_w1706_,
		_w13507_
	);
	LUT4 #(
		.INIT('h8000)
	) name12158 (
		_w13506_,
		_w13507_,
		_w13504_,
		_w13505_,
		_w13508_
	);
	LUT4 #(
		.INIT('h0111)
	) name12159 (
		_w1842_,
		_w1845_,
		_w13503_,
		_w13508_,
		_w13509_
	);
	LUT4 #(
		.INIT('h4000)
	) name12160 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13509_,
		_w13510_
	);
	LUT3 #(
		.INIT('h08)
	) name12161 (
		_w1725_,
		_w1802_,
		_w3489_,
		_w13511_
	);
	LUT2 #(
		.INIT('h2)
	) name12162 (
		_w1795_,
		_w3481_,
		_w13512_
	);
	LUT4 #(
		.INIT('h1113)
	) name12163 (
		_w1867_,
		_w13510_,
		_w13511_,
		_w13512_,
		_w13513_
	);
	LUT2 #(
		.INIT('h4)
	) name12164 (
		_w13498_,
		_w13513_,
		_w13514_
	);
	LUT4 #(
		.INIT('hecee)
	) name12165 (
		_w1933_,
		_w13495_,
		_w13496_,
		_w13514_,
		_w13515_
	);
	LUT2 #(
		.INIT('h2)
	) name12166 (
		\P1_EAX_reg[20]/NET0131 ,
		_w9102_,
		_w13516_
	);
	LUT3 #(
		.INIT('h48)
	) name12167 (
		\P1_EAX_reg[20]/NET0131 ,
		_w1827_,
		_w9430_,
		_w13517_
	);
	LUT2 #(
		.INIT('h2)
	) name12168 (
		_w1795_,
		_w3442_,
		_w13518_
	);
	LUT3 #(
		.INIT('h08)
	) name12169 (
		_w1725_,
		_w1802_,
		_w3496_,
		_w13519_
	);
	LUT4 #(
		.INIT('h153f)
	) name12170 (
		\P1_InstQueue_reg[12][4]/NET0131 ,
		\P1_InstQueue_reg[6][4]/NET0131 ,
		_w1702_,
		_w1703_,
		_w13520_
	);
	LUT4 #(
		.INIT('h153f)
	) name12171 (
		\P1_InstQueue_reg[10][4]/NET0131 ,
		\P1_InstQueue_reg[4][4]/NET0131 ,
		_w1692_,
		_w1708_,
		_w13521_
	);
	LUT4 #(
		.INIT('h153f)
	) name12172 (
		\P1_InstQueue_reg[11][4]/NET0131 ,
		\P1_InstQueue_reg[1][4]/NET0131 ,
		_w1699_,
		_w1712_,
		_w13522_
	);
	LUT4 #(
		.INIT('h153f)
	) name12173 (
		\P1_InstQueue_reg[0][4]/NET0131 ,
		\P1_InstQueue_reg[7][4]/NET0131 ,
		_w1689_,
		_w1705_,
		_w13523_
	);
	LUT4 #(
		.INIT('h8000)
	) name12174 (
		_w13522_,
		_w13523_,
		_w13520_,
		_w13521_,
		_w13524_
	);
	LUT4 #(
		.INIT('h135f)
	) name12175 (
		\P1_InstQueue_reg[14][4]/NET0131 ,
		\P1_InstQueue_reg[8][4]/NET0131 ,
		_w1696_,
		_w1691_,
		_w13525_
	);
	LUT4 #(
		.INIT('h135f)
	) name12176 (
		\P1_InstQueue_reg[15][4]/NET0131 ,
		\P1_InstQueue_reg[5][4]/NET0131 ,
		_w1698_,
		_w1709_,
		_w13526_
	);
	LUT4 #(
		.INIT('h135f)
	) name12177 (
		\P1_InstQueue_reg[13][4]/NET0131 ,
		\P1_InstQueue_reg[3][4]/NET0131 ,
		_w1694_,
		_w1688_,
		_w13527_
	);
	LUT4 #(
		.INIT('h153f)
	) name12178 (
		\P1_InstQueue_reg[2][4]/NET0131 ,
		\P1_InstQueue_reg[9][4]/NET0131 ,
		_w1711_,
		_w1706_,
		_w13528_
	);
	LUT4 #(
		.INIT('h8000)
	) name12179 (
		_w13527_,
		_w13528_,
		_w13525_,
		_w13526_,
		_w13529_
	);
	LUT4 #(
		.INIT('h0111)
	) name12180 (
		_w1842_,
		_w1845_,
		_w13524_,
		_w13529_,
		_w13530_
	);
	LUT4 #(
		.INIT('h4000)
	) name12181 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13530_,
		_w13531_
	);
	LUT4 #(
		.INIT('h0057)
	) name12182 (
		_w1867_,
		_w13518_,
		_w13519_,
		_w13531_,
		_w13532_
	);
	LUT4 #(
		.INIT('h7500)
	) name12183 (
		\P1_EAX_reg[20]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13532_,
		_w13533_
	);
	LUT4 #(
		.INIT('hecee)
	) name12184 (
		_w1933_,
		_w13516_,
		_w13517_,
		_w13533_,
		_w13534_
	);
	LUT2 #(
		.INIT('h2)
	) name12185 (
		\P1_EAX_reg[21]/NET0131 ,
		_w9102_,
		_w13535_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12186 (
		\P1_EAX_reg[20]/NET0131 ,
		\P1_EAX_reg[21]/NET0131 ,
		_w1827_,
		_w9430_,
		_w13536_
	);
	LUT3 #(
		.INIT('h08)
	) name12187 (
		_w1725_,
		_w1802_,
		_w3510_,
		_w13537_
	);
	LUT2 #(
		.INIT('h2)
	) name12188 (
		_w1795_,
		_w3452_,
		_w13538_
	);
	LUT4 #(
		.INIT('h135f)
	) name12189 (
		\P1_InstQueue_reg[14][5]/NET0131 ,
		\P1_InstQueue_reg[1][5]/NET0131 ,
		_w1696_,
		_w1699_,
		_w13539_
	);
	LUT4 #(
		.INIT('h153f)
	) name12190 (
		\P1_InstQueue_reg[11][5]/NET0131 ,
		\P1_InstQueue_reg[3][5]/NET0131 ,
		_w1688_,
		_w1712_,
		_w13540_
	);
	LUT4 #(
		.INIT('h135f)
	) name12191 (
		\P1_InstQueue_reg[15][5]/NET0131 ,
		\P1_InstQueue_reg[4][5]/NET0131 ,
		_w1698_,
		_w1692_,
		_w13541_
	);
	LUT4 #(
		.INIT('h153f)
	) name12192 (
		\P1_InstQueue_reg[0][5]/NET0131 ,
		\P1_InstQueue_reg[9][5]/NET0131 ,
		_w1711_,
		_w1705_,
		_w13542_
	);
	LUT4 #(
		.INIT('h8000)
	) name12193 (
		_w13541_,
		_w13542_,
		_w13539_,
		_w13540_,
		_w13543_
	);
	LUT4 #(
		.INIT('h135f)
	) name12194 (
		\P1_InstQueue_reg[13][5]/NET0131 ,
		\P1_InstQueue_reg[6][5]/NET0131 ,
		_w1694_,
		_w1702_,
		_w13544_
	);
	LUT4 #(
		.INIT('h153f)
	) name12195 (
		\P1_InstQueue_reg[5][5]/NET0131 ,
		\P1_InstQueue_reg[7][5]/NET0131 ,
		_w1689_,
		_w1709_,
		_w13545_
	);
	LUT4 #(
		.INIT('h135f)
	) name12196 (
		\P1_InstQueue_reg[10][5]/NET0131 ,
		\P1_InstQueue_reg[12][5]/NET0131 ,
		_w1708_,
		_w1703_,
		_w13546_
	);
	LUT4 #(
		.INIT('h153f)
	) name12197 (
		\P1_InstQueue_reg[2][5]/NET0131 ,
		\P1_InstQueue_reg[8][5]/NET0131 ,
		_w1691_,
		_w1706_,
		_w13547_
	);
	LUT4 #(
		.INIT('h8000)
	) name12198 (
		_w13546_,
		_w13547_,
		_w13544_,
		_w13545_,
		_w13548_
	);
	LUT4 #(
		.INIT('h0111)
	) name12199 (
		_w1842_,
		_w1845_,
		_w13543_,
		_w13548_,
		_w13549_
	);
	LUT4 #(
		.INIT('h4000)
	) name12200 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13549_,
		_w13550_
	);
	LUT4 #(
		.INIT('h0057)
	) name12201 (
		_w1867_,
		_w13537_,
		_w13538_,
		_w13550_,
		_w13551_
	);
	LUT4 #(
		.INIT('h7500)
	) name12202 (
		\P1_EAX_reg[21]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13551_,
		_w13552_
	);
	LUT4 #(
		.INIT('hecee)
	) name12203 (
		_w1933_,
		_w13535_,
		_w13536_,
		_w13552_,
		_w13553_
	);
	LUT2 #(
		.INIT('h2)
	) name12204 (
		\P1_EAX_reg[22]/NET0131 ,
		_w9102_,
		_w13554_
	);
	LUT4 #(
		.INIT('h4888)
	) name12205 (
		\P1_EAX_reg[22]/NET0131 ,
		_w1827_,
		_w9430_,
		_w9431_,
		_w13555_
	);
	LUT4 #(
		.INIT('h135f)
	) name12206 (
		\P1_InstQueue_reg[14][6]/NET0131 ,
		\P1_InstQueue_reg[1][6]/NET0131 ,
		_w1696_,
		_w1699_,
		_w13556_
	);
	LUT4 #(
		.INIT('h135f)
	) name12207 (
		\P1_InstQueue_reg[3][6]/NET0131 ,
		\P1_InstQueue_reg[4][6]/NET0131 ,
		_w1688_,
		_w1692_,
		_w13557_
	);
	LUT4 #(
		.INIT('h135f)
	) name12208 (
		\P1_InstQueue_reg[11][6]/NET0131 ,
		\P1_InstQueue_reg[6][6]/NET0131 ,
		_w1712_,
		_w1702_,
		_w13558_
	);
	LUT4 #(
		.INIT('h153f)
	) name12209 (
		\P1_InstQueue_reg[0][6]/NET0131 ,
		\P1_InstQueue_reg[9][6]/NET0131 ,
		_w1711_,
		_w1705_,
		_w13559_
	);
	LUT4 #(
		.INIT('h8000)
	) name12210 (
		_w13558_,
		_w13559_,
		_w13556_,
		_w13557_,
		_w13560_
	);
	LUT4 #(
		.INIT('h135f)
	) name12211 (
		\P1_InstQueue_reg[13][6]/NET0131 ,
		\P1_InstQueue_reg[7][6]/NET0131 ,
		_w1694_,
		_w1689_,
		_w13561_
	);
	LUT4 #(
		.INIT('h135f)
	) name12212 (
		\P1_InstQueue_reg[15][6]/NET0131 ,
		\P1_InstQueue_reg[5][6]/NET0131 ,
		_w1698_,
		_w1709_,
		_w13562_
	);
	LUT4 #(
		.INIT('h135f)
	) name12213 (
		\P1_InstQueue_reg[10][6]/NET0131 ,
		\P1_InstQueue_reg[12][6]/NET0131 ,
		_w1708_,
		_w1703_,
		_w13563_
	);
	LUT4 #(
		.INIT('h153f)
	) name12214 (
		\P1_InstQueue_reg[2][6]/NET0131 ,
		\P1_InstQueue_reg[8][6]/NET0131 ,
		_w1691_,
		_w1706_,
		_w13564_
	);
	LUT4 #(
		.INIT('h8000)
	) name12215 (
		_w13563_,
		_w13564_,
		_w13561_,
		_w13562_,
		_w13565_
	);
	LUT4 #(
		.INIT('h0111)
	) name12216 (
		_w1842_,
		_w1845_,
		_w13560_,
		_w13565_,
		_w13566_
	);
	LUT4 #(
		.INIT('h4000)
	) name12217 (
		_w1737_,
		_w1804_,
		_w1813_,
		_w13566_,
		_w13567_
	);
	LUT3 #(
		.INIT('h08)
	) name12218 (
		_w1725_,
		_w1802_,
		_w3503_,
		_w13568_
	);
	LUT2 #(
		.INIT('h2)
	) name12219 (
		_w1795_,
		_w3474_,
		_w13569_
	);
	LUT4 #(
		.INIT('h1113)
	) name12220 (
		_w1867_,
		_w13567_,
		_w13568_,
		_w13569_,
		_w13570_
	);
	LUT4 #(
		.INIT('h7500)
	) name12221 (
		\P1_EAX_reg[22]/NET0131 ,
		_w9436_,
		_w9437_,
		_w13570_,
		_w13571_
	);
	LUT4 #(
		.INIT('hecee)
	) name12222 (
		_w1933_,
		_w13554_,
		_w13555_,
		_w13571_,
		_w13572_
	);
	LUT2 #(
		.INIT('h2)
	) name12223 (
		\P2_More_reg/NET0131 ,
		_w7767_,
		_w13573_
	);
	LUT4 #(
		.INIT('hffb0)
	) name12224 (
		_w1665_,
		_w1669_,
		_w1678_,
		_w13573_,
		_w13574_
	);
	LUT2 #(
		.INIT('h1)
	) name12225 (
		\P2_ReadRequest_reg/NET0131 ,
		_w1656_,
		_w13575_
	);
	LUT4 #(
		.INIT('h1130)
	) name12226 (
		_w1501_,
		_w1565_,
		_w1566_,
		_w1568_,
		_w13576_
	);
	LUT3 #(
		.INIT('h8c)
	) name12227 (
		_w1603_,
		_w1678_,
		_w13576_,
		_w13577_
	);
	LUT3 #(
		.INIT('hc4)
	) name12228 (
		\P2_ReadRequest_reg/NET0131 ,
		_w2287_,
		_w12686_,
		_w13578_
	);
	LUT3 #(
		.INIT('h4f)
	) name12229 (
		_w13575_,
		_w13577_,
		_w13578_,
		_w13579_
	);
	LUT3 #(
		.INIT('hc8)
	) name12230 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		_w2215_,
		_w10611_,
		_w13580_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12231 (
		_w2033_,
		_w2038_,
		_w10611_,
		_w13580_,
		_w13581_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12232 (
		\P3_InstQueue_reg[0][3]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w13582_
	);
	LUT4 #(
		.INIT('h153f)
	) name12233 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10614_,
		_w10616_,
		_w13583_
	);
	LUT2 #(
		.INIT('h2)
	) name12234 (
		_w2199_,
		_w13583_,
		_w13584_
	);
	LUT3 #(
		.INIT('h02)
	) name12235 (
		\buf2_reg[3]/NET0131 ,
		_w10618_,
		_w10621_,
		_w13585_
	);
	LUT3 #(
		.INIT('h01)
	) name12236 (
		_w13582_,
		_w13584_,
		_w13585_,
		_w13586_
	);
	LUT2 #(
		.INIT('hb)
	) name12237 (
		_w13581_,
		_w13586_,
		_w13587_
	);
	LUT3 #(
		.INIT('hc8)
	) name12238 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		_w2215_,
		_w10611_,
		_w13588_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12239 (
		_w1959_,
		_w1972_,
		_w10611_,
		_w13588_,
		_w13589_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12240 (
		\P3_InstQueue_reg[0][6]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w13590_
	);
	LUT4 #(
		.INIT('h153f)
	) name12241 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10614_,
		_w10616_,
		_w13591_
	);
	LUT2 #(
		.INIT('h2)
	) name12242 (
		_w2199_,
		_w13591_,
		_w13592_
	);
	LUT3 #(
		.INIT('h02)
	) name12243 (
		\buf2_reg[6]/NET0131 ,
		_w10618_,
		_w10621_,
		_w13593_
	);
	LUT3 #(
		.INIT('h01)
	) name12244 (
		_w13590_,
		_w13592_,
		_w13593_,
		_w13594_
	);
	LUT2 #(
		.INIT('hb)
	) name12245 (
		_w13589_,
		_w13594_,
		_w13595_
	);
	LUT3 #(
		.INIT('hc8)
	) name12246 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		_w2215_,
		_w10630_,
		_w13596_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12247 (
		_w2033_,
		_w2038_,
		_w10630_,
		_w13596_,
		_w13597_
	);
	LUT4 #(
		.INIT('h222a)
	) name12248 (
		\P3_InstQueue_reg[10][3]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w13598_
	);
	LUT4 #(
		.INIT('h153f)
	) name12249 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10633_,
		_w10635_,
		_w13599_
	);
	LUT2 #(
		.INIT('h2)
	) name12250 (
		_w2199_,
		_w13599_,
		_w13600_
	);
	LUT3 #(
		.INIT('h20)
	) name12251 (
		\buf2_reg[3]/NET0131 ,
		_w10637_,
		_w10639_,
		_w13601_
	);
	LUT3 #(
		.INIT('h01)
	) name12252 (
		_w13598_,
		_w13600_,
		_w13601_,
		_w13602_
	);
	LUT2 #(
		.INIT('hb)
	) name12253 (
		_w13597_,
		_w13602_,
		_w13603_
	);
	LUT3 #(
		.INIT('hc8)
	) name12254 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		_w2215_,
		_w10630_,
		_w13604_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12255 (
		_w1959_,
		_w1972_,
		_w10630_,
		_w13604_,
		_w13605_
	);
	LUT4 #(
		.INIT('h222a)
	) name12256 (
		\P3_InstQueue_reg[10][6]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w13606_
	);
	LUT4 #(
		.INIT('h153f)
	) name12257 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10633_,
		_w10635_,
		_w13607_
	);
	LUT2 #(
		.INIT('h2)
	) name12258 (
		_w2199_,
		_w13607_,
		_w13608_
	);
	LUT3 #(
		.INIT('h20)
	) name12259 (
		\buf2_reg[6]/NET0131 ,
		_w10637_,
		_w10639_,
		_w13609_
	);
	LUT3 #(
		.INIT('h01)
	) name12260 (
		_w13606_,
		_w13608_,
		_w13609_,
		_w13610_
	);
	LUT2 #(
		.INIT('hb)
	) name12261 (
		_w13605_,
		_w13610_,
		_w13611_
	);
	LUT3 #(
		.INIT('hc8)
	) name12262 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		_w2215_,
		_w10646_,
		_w13612_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12263 (
		_w2033_,
		_w2038_,
		_w10646_,
		_w13612_,
		_w13613_
	);
	LUT3 #(
		.INIT('ha2)
	) name12264 (
		\P3_InstQueue_reg[11][3]/NET0131 ,
		_w10622_,
		_w10650_,
		_w13614_
	);
	LUT3 #(
		.INIT('hd8)
	) name12265 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w13615_
	);
	LUT3 #(
		.INIT('h80)
	) name12266 (
		_w2194_,
		_w10649_,
		_w13615_,
		_w13616_
	);
	LUT4 #(
		.INIT('h2000)
	) name12267 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w13617_
	);
	LUT4 #(
		.INIT('hce00)
	) name12268 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w13617_,
		_w13618_
	);
	LUT2 #(
		.INIT('h1)
	) name12269 (
		_w13616_,
		_w13618_,
		_w13619_
	);
	LUT2 #(
		.INIT('h4)
	) name12270 (
		_w13614_,
		_w13619_,
		_w13620_
	);
	LUT2 #(
		.INIT('hb)
	) name12271 (
		_w13613_,
		_w13620_,
		_w13621_
	);
	LUT3 #(
		.INIT('hc8)
	) name12272 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w2215_,
		_w10646_,
		_w13622_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12273 (
		_w1959_,
		_w1972_,
		_w10646_,
		_w13622_,
		_w13623_
	);
	LUT3 #(
		.INIT('ha2)
	) name12274 (
		\P3_InstQueue_reg[11][6]/NET0131 ,
		_w10622_,
		_w10650_,
		_w13624_
	);
	LUT3 #(
		.INIT('hd8)
	) name12275 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w13625_
	);
	LUT3 #(
		.INIT('h80)
	) name12276 (
		_w2194_,
		_w10649_,
		_w13625_,
		_w13626_
	);
	LUT4 #(
		.INIT('h2000)
	) name12277 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w13627_
	);
	LUT4 #(
		.INIT('hce00)
	) name12278 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w13627_,
		_w13628_
	);
	LUT2 #(
		.INIT('h1)
	) name12279 (
		_w13626_,
		_w13628_,
		_w13629_
	);
	LUT2 #(
		.INIT('h4)
	) name12280 (
		_w13624_,
		_w13629_,
		_w13630_
	);
	LUT2 #(
		.INIT('hb)
	) name12281 (
		_w13623_,
		_w13630_,
		_w13631_
	);
	LUT3 #(
		.INIT('hc8)
	) name12282 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		_w2215_,
		_w10659_,
		_w13632_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12283 (
		_w2033_,
		_w2038_,
		_w10659_,
		_w13632_,
		_w13633_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12284 (
		\P3_InstQueue_reg[12][3]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w13634_
	);
	LUT4 #(
		.INIT('h135f)
	) name12285 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10630_,
		_w10652_,
		_w13635_
	);
	LUT2 #(
		.INIT('h2)
	) name12286 (
		_w2199_,
		_w13635_,
		_w13636_
	);
	LUT3 #(
		.INIT('h02)
	) name12287 (
		\buf2_reg[3]/NET0131 ,
		_w10662_,
		_w10663_,
		_w13637_
	);
	LUT3 #(
		.INIT('h01)
	) name12288 (
		_w13634_,
		_w13636_,
		_w13637_,
		_w13638_
	);
	LUT2 #(
		.INIT('hb)
	) name12289 (
		_w13633_,
		_w13638_,
		_w13639_
	);
	LUT3 #(
		.INIT('hc8)
	) name12290 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w2215_,
		_w10659_,
		_w13640_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12291 (
		_w1959_,
		_w1972_,
		_w10659_,
		_w13640_,
		_w13641_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12292 (
		\P3_InstQueue_reg[12][6]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w13642_
	);
	LUT4 #(
		.INIT('h135f)
	) name12293 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10630_,
		_w10652_,
		_w13643_
	);
	LUT2 #(
		.INIT('h2)
	) name12294 (
		_w2199_,
		_w13643_,
		_w13644_
	);
	LUT3 #(
		.INIT('h02)
	) name12295 (
		\buf2_reg[6]/NET0131 ,
		_w10662_,
		_w10663_,
		_w13645_
	);
	LUT3 #(
		.INIT('h01)
	) name12296 (
		_w13642_,
		_w13644_,
		_w13645_,
		_w13646_
	);
	LUT2 #(
		.INIT('hb)
	) name12297 (
		_w13641_,
		_w13646_,
		_w13647_
	);
	LUT3 #(
		.INIT('hc8)
	) name12298 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w2215_,
		_w10614_,
		_w13648_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12299 (
		_w2033_,
		_w2038_,
		_w10614_,
		_w13648_,
		_w13649_
	);
	LUT2 #(
		.INIT('h4)
	) name12300 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w10672_,
		_w13650_
	);
	LUT2 #(
		.INIT('h1)
	) name12301 (
		\buf2_reg[3]/NET0131 ,
		_w10672_,
		_w13651_
	);
	LUT3 #(
		.INIT('h02)
	) name12302 (
		_w10674_,
		_w13651_,
		_w13650_,
		_w13652_
	);
	LUT3 #(
		.INIT('h80)
	) name12303 (
		_w2194_,
		_w10673_,
		_w13615_,
		_w13653_
	);
	LUT2 #(
		.INIT('h2)
	) name12304 (
		\P3_InstQueue_reg[13][3]/NET0131 ,
		_w10622_,
		_w13654_
	);
	LUT2 #(
		.INIT('h1)
	) name12305 (
		_w13653_,
		_w13654_,
		_w13655_
	);
	LUT2 #(
		.INIT('h4)
	) name12306 (
		_w13652_,
		_w13655_,
		_w13656_
	);
	LUT2 #(
		.INIT('hb)
	) name12307 (
		_w13649_,
		_w13656_,
		_w13657_
	);
	LUT3 #(
		.INIT('hc8)
	) name12308 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w2215_,
		_w10614_,
		_w13658_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12309 (
		_w1959_,
		_w1972_,
		_w10614_,
		_w13658_,
		_w13659_
	);
	LUT2 #(
		.INIT('h4)
	) name12310 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w10672_,
		_w13660_
	);
	LUT2 #(
		.INIT('h1)
	) name12311 (
		\buf2_reg[6]/NET0131 ,
		_w10672_,
		_w13661_
	);
	LUT3 #(
		.INIT('h02)
	) name12312 (
		_w10674_,
		_w13661_,
		_w13660_,
		_w13662_
	);
	LUT2 #(
		.INIT('h2)
	) name12313 (
		\P3_InstQueue_reg[13][6]/NET0131 ,
		_w10622_,
		_w13663_
	);
	LUT3 #(
		.INIT('h80)
	) name12314 (
		_w2194_,
		_w10673_,
		_w13625_,
		_w13664_
	);
	LUT2 #(
		.INIT('h1)
	) name12315 (
		_w13663_,
		_w13664_,
		_w13665_
	);
	LUT2 #(
		.INIT('h4)
	) name12316 (
		_w13662_,
		_w13665_,
		_w13666_
	);
	LUT2 #(
		.INIT('hb)
	) name12317 (
		_w13659_,
		_w13666_,
		_w13667_
	);
	LUT3 #(
		.INIT('hc8)
	) name12318 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w2215_,
		_w10616_,
		_w13668_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12319 (
		_w2033_,
		_w2038_,
		_w10616_,
		_w13668_,
		_w13669_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12320 (
		\P3_InstQueue_reg[14][3]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w13670_
	);
	LUT4 #(
		.INIT('h153f)
	) name12321 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10646_,
		_w10659_,
		_w13671_
	);
	LUT2 #(
		.INIT('h2)
	) name12322 (
		_w2199_,
		_w13671_,
		_w13672_
	);
	LUT3 #(
		.INIT('h02)
	) name12323 (
		\buf2_reg[3]/NET0131 ,
		_w10617_,
		_w10684_,
		_w13673_
	);
	LUT3 #(
		.INIT('h01)
	) name12324 (
		_w13670_,
		_w13672_,
		_w13673_,
		_w13674_
	);
	LUT2 #(
		.INIT('hb)
	) name12325 (
		_w13669_,
		_w13674_,
		_w13675_
	);
	LUT3 #(
		.INIT('hc8)
	) name12326 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w2215_,
		_w10616_,
		_w13676_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12327 (
		_w1959_,
		_w1972_,
		_w10616_,
		_w13676_,
		_w13677_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12328 (
		\P3_InstQueue_reg[14][6]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w13678_
	);
	LUT4 #(
		.INIT('h153f)
	) name12329 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10646_,
		_w10659_,
		_w13679_
	);
	LUT2 #(
		.INIT('h2)
	) name12330 (
		_w2199_,
		_w13679_,
		_w13680_
	);
	LUT3 #(
		.INIT('h02)
	) name12331 (
		\buf2_reg[6]/NET0131 ,
		_w10617_,
		_w10684_,
		_w13681_
	);
	LUT3 #(
		.INIT('h01)
	) name12332 (
		_w13678_,
		_w13680_,
		_w13681_,
		_w13682_
	);
	LUT2 #(
		.INIT('hb)
	) name12333 (
		_w13677_,
		_w13682_,
		_w13683_
	);
	LUT3 #(
		.INIT('hc8)
	) name12334 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w2215_,
		_w10620_,
		_w13684_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12335 (
		_w2033_,
		_w2038_,
		_w10620_,
		_w13684_,
		_w13685_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12336 (
		\P3_InstQueue_reg[15][3]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w13686_
	);
	LUT4 #(
		.INIT('h135f)
	) name12337 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10614_,
		_w10659_,
		_w13687_
	);
	LUT2 #(
		.INIT('h2)
	) name12338 (
		_w2199_,
		_w13687_,
		_w13688_
	);
	LUT3 #(
		.INIT('h02)
	) name12339 (
		\buf2_reg[3]/NET0131 ,
		_w10693_,
		_w10694_,
		_w13689_
	);
	LUT3 #(
		.INIT('h01)
	) name12340 (
		_w13686_,
		_w13688_,
		_w13689_,
		_w13690_
	);
	LUT2 #(
		.INIT('hb)
	) name12341 (
		_w13685_,
		_w13690_,
		_w13691_
	);
	LUT3 #(
		.INIT('hc8)
	) name12342 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w2215_,
		_w10620_,
		_w13692_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12343 (
		_w1959_,
		_w1972_,
		_w10620_,
		_w13692_,
		_w13693_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12344 (
		\P3_InstQueue_reg[15][6]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w13694_
	);
	LUT4 #(
		.INIT('h135f)
	) name12345 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10614_,
		_w10659_,
		_w13695_
	);
	LUT2 #(
		.INIT('h2)
	) name12346 (
		_w2199_,
		_w13695_,
		_w13696_
	);
	LUT3 #(
		.INIT('h02)
	) name12347 (
		\buf2_reg[6]/NET0131 ,
		_w10693_,
		_w10694_,
		_w13697_
	);
	LUT3 #(
		.INIT('h01)
	) name12348 (
		_w13694_,
		_w13696_,
		_w13697_,
		_w13698_
	);
	LUT2 #(
		.INIT('hb)
	) name12349 (
		_w13693_,
		_w13698_,
		_w13699_
	);
	LUT3 #(
		.INIT('hc8)
	) name12350 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w2215_,
		_w10701_,
		_w13700_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12351 (
		_w2033_,
		_w2038_,
		_w10701_,
		_w13700_,
		_w13701_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12352 (
		\P3_InstQueue_reg[1][3]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w13702_
	);
	LUT4 #(
		.INIT('h153f)
	) name12353 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10616_,
		_w10620_,
		_w13703_
	);
	LUT2 #(
		.INIT('h2)
	) name12354 (
		_w2199_,
		_w13703_,
		_w13704_
	);
	LUT3 #(
		.INIT('h02)
	) name12355 (
		\buf2_reg[3]/NET0131 ,
		_w10704_,
		_w10705_,
		_w13705_
	);
	LUT3 #(
		.INIT('h01)
	) name12356 (
		_w13702_,
		_w13704_,
		_w13705_,
		_w13706_
	);
	LUT2 #(
		.INIT('hb)
	) name12357 (
		_w13701_,
		_w13706_,
		_w13707_
	);
	LUT3 #(
		.INIT('hc8)
	) name12358 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w2215_,
		_w10701_,
		_w13708_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12359 (
		_w1959_,
		_w1972_,
		_w10701_,
		_w13708_,
		_w13709_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12360 (
		\P3_InstQueue_reg[1][6]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w13710_
	);
	LUT4 #(
		.INIT('h153f)
	) name12361 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10616_,
		_w10620_,
		_w13711_
	);
	LUT2 #(
		.INIT('h2)
	) name12362 (
		_w2199_,
		_w13711_,
		_w13712_
	);
	LUT3 #(
		.INIT('h02)
	) name12363 (
		\buf2_reg[6]/NET0131 ,
		_w10704_,
		_w10705_,
		_w13713_
	);
	LUT3 #(
		.INIT('h01)
	) name12364 (
		_w13710_,
		_w13712_,
		_w13713_,
		_w13714_
	);
	LUT2 #(
		.INIT('hb)
	) name12365 (
		_w13709_,
		_w13714_,
		_w13715_
	);
	LUT3 #(
		.INIT('hc8)
	) name12366 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w2215_,
		_w10713_,
		_w13716_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12367 (
		_w2033_,
		_w2038_,
		_w10713_,
		_w13716_,
		_w13717_
	);
	LUT4 #(
		.INIT('h222a)
	) name12368 (
		\P3_InstQueue_reg[2][3]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w13718_
	);
	LUT4 #(
		.INIT('h135f)
	) name12369 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10611_,
		_w10620_,
		_w13719_
	);
	LUT2 #(
		.INIT('h2)
	) name12370 (
		_w2199_,
		_w13719_,
		_w13720_
	);
	LUT3 #(
		.INIT('h20)
	) name12371 (
		\buf2_reg[3]/NET0131 ,
		_w10716_,
		_w10717_,
		_w13721_
	);
	LUT3 #(
		.INIT('h01)
	) name12372 (
		_w13718_,
		_w13720_,
		_w13721_,
		_w13722_
	);
	LUT2 #(
		.INIT('hb)
	) name12373 (
		_w13717_,
		_w13722_,
		_w13723_
	);
	LUT3 #(
		.INIT('hc8)
	) name12374 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w2215_,
		_w10713_,
		_w13724_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12375 (
		_w1959_,
		_w1972_,
		_w10713_,
		_w13724_,
		_w13725_
	);
	LUT4 #(
		.INIT('h222a)
	) name12376 (
		\P3_InstQueue_reg[2][6]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w13726_
	);
	LUT4 #(
		.INIT('h135f)
	) name12377 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10611_,
		_w10620_,
		_w13727_
	);
	LUT2 #(
		.INIT('h2)
	) name12378 (
		_w2199_,
		_w13727_,
		_w13728_
	);
	LUT3 #(
		.INIT('h20)
	) name12379 (
		\buf2_reg[6]/NET0131 ,
		_w10716_,
		_w10717_,
		_w13729_
	);
	LUT3 #(
		.INIT('h01)
	) name12380 (
		_w13726_,
		_w13728_,
		_w13729_,
		_w13730_
	);
	LUT2 #(
		.INIT('hb)
	) name12381 (
		_w13725_,
		_w13730_,
		_w13731_
	);
	LUT3 #(
		.INIT('hc8)
	) name12382 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w2215_,
		_w10724_,
		_w13732_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12383 (
		_w2033_,
		_w2038_,
		_w10724_,
		_w13732_,
		_w13733_
	);
	LUT4 #(
		.INIT('h222a)
	) name12384 (
		\P3_InstQueue_reg[3][3]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w13734_
	);
	LUT4 #(
		.INIT('h153f)
	) name12385 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10611_,
		_w10701_,
		_w13735_
	);
	LUT2 #(
		.INIT('h2)
	) name12386 (
		_w2199_,
		_w13735_,
		_w13736_
	);
	LUT3 #(
		.INIT('h08)
	) name12387 (
		\buf2_reg[3]/NET0131 ,
		_w10712_,
		_w10727_,
		_w13737_
	);
	LUT3 #(
		.INIT('h01)
	) name12388 (
		_w13734_,
		_w13736_,
		_w13737_,
		_w13738_
	);
	LUT2 #(
		.INIT('hb)
	) name12389 (
		_w13733_,
		_w13738_,
		_w13739_
	);
	LUT3 #(
		.INIT('hc8)
	) name12390 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w2215_,
		_w10724_,
		_w13740_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12391 (
		_w1959_,
		_w1972_,
		_w10724_,
		_w13740_,
		_w13741_
	);
	LUT4 #(
		.INIT('h222a)
	) name12392 (
		\P3_InstQueue_reg[3][6]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w13742_
	);
	LUT4 #(
		.INIT('h153f)
	) name12393 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10611_,
		_w10701_,
		_w13743_
	);
	LUT2 #(
		.INIT('h2)
	) name12394 (
		_w2199_,
		_w13743_,
		_w13744_
	);
	LUT3 #(
		.INIT('h08)
	) name12395 (
		\buf2_reg[6]/NET0131 ,
		_w10712_,
		_w10727_,
		_w13745_
	);
	LUT3 #(
		.INIT('h01)
	) name12396 (
		_w13742_,
		_w13744_,
		_w13745_,
		_w13746_
	);
	LUT2 #(
		.INIT('hb)
	) name12397 (
		_w13741_,
		_w13746_,
		_w13747_
	);
	LUT3 #(
		.INIT('hc8)
	) name12398 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w2215_,
		_w10734_,
		_w13748_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12399 (
		_w2033_,
		_w2038_,
		_w10734_,
		_w13748_,
		_w13749_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12400 (
		\P3_InstQueue_reg[4][3]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w13750_
	);
	LUT4 #(
		.INIT('h153f)
	) name12401 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10701_,
		_w10713_,
		_w13751_
	);
	LUT2 #(
		.INIT('h2)
	) name12402 (
		_w2199_,
		_w13751_,
		_w13752_
	);
	LUT3 #(
		.INIT('h02)
	) name12403 (
		\buf2_reg[3]/NET0131 ,
		_w10737_,
		_w10738_,
		_w13753_
	);
	LUT3 #(
		.INIT('h01)
	) name12404 (
		_w13750_,
		_w13752_,
		_w13753_,
		_w13754_
	);
	LUT2 #(
		.INIT('hb)
	) name12405 (
		_w13749_,
		_w13754_,
		_w13755_
	);
	LUT3 #(
		.INIT('hc8)
	) name12406 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w2215_,
		_w10734_,
		_w13756_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12407 (
		_w1959_,
		_w1972_,
		_w10734_,
		_w13756_,
		_w13757_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12408 (
		\P3_InstQueue_reg[4][6]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w13758_
	);
	LUT4 #(
		.INIT('h153f)
	) name12409 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10701_,
		_w10713_,
		_w13759_
	);
	LUT2 #(
		.INIT('h2)
	) name12410 (
		_w2199_,
		_w13759_,
		_w13760_
	);
	LUT3 #(
		.INIT('h02)
	) name12411 (
		\buf2_reg[6]/NET0131 ,
		_w10737_,
		_w10738_,
		_w13761_
	);
	LUT3 #(
		.INIT('h01)
	) name12412 (
		_w13758_,
		_w13760_,
		_w13761_,
		_w13762_
	);
	LUT2 #(
		.INIT('hb)
	) name12413 (
		_w13757_,
		_w13762_,
		_w13763_
	);
	LUT3 #(
		.INIT('hc8)
	) name12414 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w2215_,
		_w10745_,
		_w13764_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12415 (
		_w2033_,
		_w2038_,
		_w10745_,
		_w13764_,
		_w13765_
	);
	LUT2 #(
		.INIT('h4)
	) name12416 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w10748_,
		_w13766_
	);
	LUT2 #(
		.INIT('h1)
	) name12417 (
		\buf2_reg[3]/NET0131 ,
		_w10748_,
		_w13767_
	);
	LUT3 #(
		.INIT('h02)
	) name12418 (
		_w10750_,
		_w13767_,
		_w13766_,
		_w13768_
	);
	LUT3 #(
		.INIT('h80)
	) name12419 (
		_w2194_,
		_w10749_,
		_w13615_,
		_w13769_
	);
	LUT2 #(
		.INIT('h2)
	) name12420 (
		\P3_InstQueue_reg[5][3]/NET0131 ,
		_w10622_,
		_w13770_
	);
	LUT2 #(
		.INIT('h1)
	) name12421 (
		_w13769_,
		_w13770_,
		_w13771_
	);
	LUT2 #(
		.INIT('h4)
	) name12422 (
		_w13768_,
		_w13771_,
		_w13772_
	);
	LUT2 #(
		.INIT('hb)
	) name12423 (
		_w13765_,
		_w13772_,
		_w13773_
	);
	LUT3 #(
		.INIT('hc8)
	) name12424 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w2215_,
		_w10745_,
		_w13774_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12425 (
		_w1959_,
		_w1972_,
		_w10745_,
		_w13774_,
		_w13775_
	);
	LUT2 #(
		.INIT('h4)
	) name12426 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w10748_,
		_w13776_
	);
	LUT2 #(
		.INIT('h1)
	) name12427 (
		\buf2_reg[6]/NET0131 ,
		_w10748_,
		_w13777_
	);
	LUT3 #(
		.INIT('h02)
	) name12428 (
		_w10750_,
		_w13777_,
		_w13776_,
		_w13778_
	);
	LUT2 #(
		.INIT('h2)
	) name12429 (
		\P3_InstQueue_reg[5][6]/NET0131 ,
		_w10622_,
		_w13779_
	);
	LUT3 #(
		.INIT('h80)
	) name12430 (
		_w2194_,
		_w10749_,
		_w13625_,
		_w13780_
	);
	LUT2 #(
		.INIT('h1)
	) name12431 (
		_w13779_,
		_w13780_,
		_w13781_
	);
	LUT2 #(
		.INIT('h4)
	) name12432 (
		_w13778_,
		_w13781_,
		_w13782_
	);
	LUT2 #(
		.INIT('hb)
	) name12433 (
		_w13775_,
		_w13782_,
		_w13783_
	);
	LUT3 #(
		.INIT('hc8)
	) name12434 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w2215_,
		_w10758_,
		_w13784_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12435 (
		_w2033_,
		_w2038_,
		_w10758_,
		_w13784_,
		_w13785_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12436 (
		\P3_InstQueue_reg[6][3]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w13786_
	);
	LUT4 #(
		.INIT('h153f)
	) name12437 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10724_,
		_w10734_,
		_w13787_
	);
	LUT2 #(
		.INIT('h2)
	) name12438 (
		_w2199_,
		_w13787_,
		_w13788_
	);
	LUT3 #(
		.INIT('h02)
	) name12439 (
		\buf2_reg[3]/NET0131 ,
		_w10761_,
		_w10762_,
		_w13789_
	);
	LUT3 #(
		.INIT('h01)
	) name12440 (
		_w13786_,
		_w13788_,
		_w13789_,
		_w13790_
	);
	LUT2 #(
		.INIT('hb)
	) name12441 (
		_w13785_,
		_w13790_,
		_w13791_
	);
	LUT3 #(
		.INIT('hc8)
	) name12442 (
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w2215_,
		_w10758_,
		_w13792_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12443 (
		_w1959_,
		_w1972_,
		_w10758_,
		_w13792_,
		_w13793_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12444 (
		\P3_InstQueue_reg[6][6]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w13794_
	);
	LUT4 #(
		.INIT('h153f)
	) name12445 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10724_,
		_w10734_,
		_w13795_
	);
	LUT2 #(
		.INIT('h2)
	) name12446 (
		_w2199_,
		_w13795_,
		_w13796_
	);
	LUT3 #(
		.INIT('h02)
	) name12447 (
		\buf2_reg[6]/NET0131 ,
		_w10761_,
		_w10762_,
		_w13797_
	);
	LUT3 #(
		.INIT('h01)
	) name12448 (
		_w13794_,
		_w13796_,
		_w13797_,
		_w13798_
	);
	LUT2 #(
		.INIT('hb)
	) name12449 (
		_w13793_,
		_w13798_,
		_w13799_
	);
	LUT3 #(
		.INIT('hc8)
	) name12450 (
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w2215_,
		_w10633_,
		_w13800_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12451 (
		_w2033_,
		_w2038_,
		_w10633_,
		_w13800_,
		_w13801_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12452 (
		\P3_InstQueue_reg[7][3]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w13802_
	);
	LUT4 #(
		.INIT('h153f)
	) name12453 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10734_,
		_w10745_,
		_w13803_
	);
	LUT2 #(
		.INIT('h2)
	) name12454 (
		_w2199_,
		_w13803_,
		_w13804_
	);
	LUT3 #(
		.INIT('h02)
	) name12455 (
		\buf2_reg[3]/NET0131 ,
		_w10771_,
		_w10772_,
		_w13805_
	);
	LUT3 #(
		.INIT('h01)
	) name12456 (
		_w13802_,
		_w13804_,
		_w13805_,
		_w13806_
	);
	LUT2 #(
		.INIT('hb)
	) name12457 (
		_w13801_,
		_w13806_,
		_w13807_
	);
	LUT3 #(
		.INIT('hc8)
	) name12458 (
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w2215_,
		_w10633_,
		_w13808_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12459 (
		_w1959_,
		_w1972_,
		_w10633_,
		_w13808_,
		_w13809_
	);
	LUT4 #(
		.INIT('h2a22)
	) name12460 (
		\P3_InstQueue_reg[7][6]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w13810_
	);
	LUT4 #(
		.INIT('h153f)
	) name12461 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10734_,
		_w10745_,
		_w13811_
	);
	LUT2 #(
		.INIT('h2)
	) name12462 (
		_w2199_,
		_w13811_,
		_w13812_
	);
	LUT3 #(
		.INIT('h02)
	) name12463 (
		\buf2_reg[6]/NET0131 ,
		_w10771_,
		_w10772_,
		_w13813_
	);
	LUT3 #(
		.INIT('h01)
	) name12464 (
		_w13810_,
		_w13812_,
		_w13813_,
		_w13814_
	);
	LUT2 #(
		.INIT('hb)
	) name12465 (
		_w13809_,
		_w13814_,
		_w13815_
	);
	LUT3 #(
		.INIT('hc8)
	) name12466 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w2215_,
		_w10635_,
		_w13816_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12467 (
		_w2033_,
		_w2038_,
		_w10635_,
		_w13816_,
		_w13817_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12468 (
		\P3_InstQueue_reg[8][3]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w13818_
	);
	LUT4 #(
		.INIT('h153f)
	) name12469 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10745_,
		_w10758_,
		_w13819_
	);
	LUT2 #(
		.INIT('h2)
	) name12470 (
		_w2199_,
		_w13819_,
		_w13820_
	);
	LUT3 #(
		.INIT('h02)
	) name12471 (
		\buf2_reg[3]/NET0131 ,
		_w10636_,
		_w10781_,
		_w13821_
	);
	LUT3 #(
		.INIT('h01)
	) name12472 (
		_w13818_,
		_w13820_,
		_w13821_,
		_w13822_
	);
	LUT2 #(
		.INIT('hb)
	) name12473 (
		_w13817_,
		_w13822_,
		_w13823_
	);
	LUT3 #(
		.INIT('hc8)
	) name12474 (
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w2215_,
		_w10635_,
		_w13824_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12475 (
		_w1959_,
		_w1972_,
		_w10635_,
		_w13824_,
		_w13825_
	);
	LUT4 #(
		.INIT('h22a2)
	) name12476 (
		\P3_InstQueue_reg[8][6]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w13826_
	);
	LUT4 #(
		.INIT('h153f)
	) name12477 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10745_,
		_w10758_,
		_w13827_
	);
	LUT2 #(
		.INIT('h2)
	) name12478 (
		_w2199_,
		_w13827_,
		_w13828_
	);
	LUT3 #(
		.INIT('h02)
	) name12479 (
		\buf2_reg[6]/NET0131 ,
		_w10636_,
		_w10781_,
		_w13829_
	);
	LUT3 #(
		.INIT('h01)
	) name12480 (
		_w13826_,
		_w13828_,
		_w13829_,
		_w13830_
	);
	LUT2 #(
		.INIT('hb)
	) name12481 (
		_w13825_,
		_w13830_,
		_w13831_
	);
	LUT3 #(
		.INIT('hc8)
	) name12482 (
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w2215_,
		_w10652_,
		_w13832_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12483 (
		_w2033_,
		_w2038_,
		_w10652_,
		_w13832_,
		_w13833_
	);
	LUT4 #(
		.INIT('h135f)
	) name12484 (
		\buf2_reg[19]/NET0131 ,
		\buf2_reg[27]/NET0131 ,
		_w10633_,
		_w10758_,
		_w13834_
	);
	LUT4 #(
		.INIT('hef00)
	) name12485 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w13835_
	);
	LUT4 #(
		.INIT('h1000)
	) name12486 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w13836_
	);
	LUT4 #(
		.INIT('hddd0)
	) name12487 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w13835_,
		_w13836_,
		_w13837_
	);
	LUT4 #(
		.INIT('hcc08)
	) name12488 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w13834_,
		_w13837_,
		_w13838_
	);
	LUT3 #(
		.INIT('ha8)
	) name12489 (
		_w3055_,
		_w13835_,
		_w13836_,
		_w13839_
	);
	LUT2 #(
		.INIT('h2)
	) name12490 (
		\P3_InstQueue_reg[9][3]/NET0131 ,
		_w10622_,
		_w13840_
	);
	LUT2 #(
		.INIT('h1)
	) name12491 (
		_w13839_,
		_w13840_,
		_w13841_
	);
	LUT2 #(
		.INIT('h4)
	) name12492 (
		_w13838_,
		_w13841_,
		_w13842_
	);
	LUT2 #(
		.INIT('hb)
	) name12493 (
		_w13833_,
		_w13842_,
		_w13843_
	);
	LUT3 #(
		.INIT('hc8)
	) name12494 (
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w2215_,
		_w10652_,
		_w13844_
	);
	LUT4 #(
		.INIT('h7f00)
	) name12495 (
		_w1959_,
		_w1972_,
		_w10652_,
		_w13844_,
		_w13845_
	);
	LUT4 #(
		.INIT('h135f)
	) name12496 (
		\buf2_reg[22]/NET0131 ,
		\buf2_reg[30]/NET0131 ,
		_w10633_,
		_w10758_,
		_w13846_
	);
	LUT4 #(
		.INIT('hef00)
	) name12497 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w13847_
	);
	LUT4 #(
		.INIT('h1000)
	) name12498 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w13848_
	);
	LUT4 #(
		.INIT('hddd0)
	) name12499 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w13847_,
		_w13848_,
		_w13849_
	);
	LUT4 #(
		.INIT('hcc08)
	) name12500 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w13846_,
		_w13849_,
		_w13850_
	);
	LUT3 #(
		.INIT('ha8)
	) name12501 (
		_w3055_,
		_w13847_,
		_w13848_,
		_w13851_
	);
	LUT2 #(
		.INIT('h2)
	) name12502 (
		\P3_InstQueue_reg[9][6]/NET0131 ,
		_w10622_,
		_w13852_
	);
	LUT2 #(
		.INIT('h1)
	) name12503 (
		_w13851_,
		_w13852_,
		_w13853_
	);
	LUT2 #(
		.INIT('h4)
	) name12504 (
		_w13850_,
		_w13853_,
		_w13854_
	);
	LUT2 #(
		.INIT('hb)
	) name12505 (
		_w13845_,
		_w13854_,
		_w13855_
	);
	LUT4 #(
		.INIT('h000d)
	) name12506 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		_w7422_,
		_w8759_,
		_w8760_,
		_w13856_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12507 (
		\P3_PhyAddrPointer_reg[0]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w3054_,
		_w3056_,
		_w13857_
	);
	LUT3 #(
		.INIT('h2f)
	) name12508 (
		_w1945_,
		_w13856_,
		_w13857_,
		_w13858_
	);
	LUT4 #(
		.INIT('h00e4)
	) name12509 (
		_w2060_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w13859_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name12510 (
		\P3_ReadRequest_reg/NET0131 ,
		_w1945_,
		_w2108_,
		_w13859_,
		_w13860_
	);
	LUT3 #(
		.INIT('hc4)
	) name12511 (
		\P3_ReadRequest_reg/NET0131 ,
		_w9129_,
		_w12679_,
		_w13861_
	);
	LUT2 #(
		.INIT('hb)
	) name12512 (
		_w13860_,
		_w13861_,
		_w13862_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12513 (
		\P1_PhyAddrPointer_reg[0]/NET0131 ,
		_w1933_,
		_w7547_,
		_w3408_,
		_w13863_
	);
	LUT2 #(
		.INIT('h8)
	) name12514 (
		_w1810_,
		_w8802_,
		_w13864_
	);
	LUT4 #(
		.INIT('h1113)
	) name12515 (
		_w1933_,
		_w8808_,
		_w8805_,
		_w13864_,
		_w13865_
	);
	LUT2 #(
		.INIT('hb)
	) name12516 (
		_w13863_,
		_w13865_,
		_w13866_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name12517 (
		\P1_ReadRequest_reg/NET0131 ,
		_w1855_,
		_w1933_,
		_w4739_,
		_w13867_
	);
	LUT3 #(
		.INIT('hc4)
	) name12518 (
		\P1_ReadRequest_reg/NET0131 ,
		_w8459_,
		_w9470_,
		_w13868_
	);
	LUT2 #(
		.INIT('hb)
	) name12519 (
		_w13867_,
		_w13868_,
		_w13869_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12520 (
		\P2_PhyAddrPointer_reg[0]/NET0131 ,
		_w1678_,
		_w7642_,
		_w4441_,
		_w13870_
	);
	LUT2 #(
		.INIT('h8)
	) name12521 (
		_w1559_,
		_w8790_,
		_w13871_
	);
	LUT4 #(
		.INIT('h1113)
	) name12522 (
		_w1678_,
		_w8796_,
		_w8793_,
		_w13871_,
		_w13872_
	);
	LUT2 #(
		.INIT('hb)
	) name12523 (
		_w13870_,
		_w13872_,
		_w13873_
	);
	LUT4 #(
		.INIT('h2220)
	) name12524 (
		_w1559_,
		_w1661_,
		_w8819_,
		_w8820_,
		_w13874_
	);
	LUT4 #(
		.INIT('h000d)
	) name12525 (
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w7642_,
		_w8825_,
		_w13874_,
		_w13875_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12526 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w1679_,
		_w5747_,
		_w13876_
	);
	LUT4 #(
		.INIT('h3310)
	) name12527 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_PhyAddrPointer_reg[1]/NET0131 ,
		_w1679_,
		_w2283_,
		_w13877_
	);
	LUT3 #(
		.INIT('h01)
	) name12528 (
		_w8830_,
		_w13877_,
		_w13876_,
		_w13878_
	);
	LUT3 #(
		.INIT('h2f)
	) name12529 (
		_w1678_,
		_w13875_,
		_w13878_,
		_w13879_
	);
	LUT2 #(
		.INIT('h8)
	) name12530 (
		_w2171_,
		_w8775_,
		_w13880_
	);
	LUT3 #(
		.INIT('h0d)
	) name12531 (
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w7422_,
		_w8780_,
		_w13881_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12532 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w2194_,
		_w5783_,
		_w13882_
	);
	LUT4 #(
		.INIT('h3310)
	) name12533 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w13883_
	);
	LUT3 #(
		.INIT('h01)
	) name12534 (
		_w8784_,
		_w13883_,
		_w13882_,
		_w13884_
	);
	LUT4 #(
		.INIT('h8aff)
	) name12535 (
		_w1945_,
		_w13880_,
		_w13881_,
		_w13884_,
		_w13885_
	);
	LUT4 #(
		.INIT('h000d)
	) name12536 (
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w7547_,
		_w8843_,
		_w8845_,
		_w13886_
	);
	LUT4 #(
		.INIT('h80cc)
	) name12537 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w1939_,
		_w6383_,
		_w13887_
	);
	LUT4 #(
		.INIT('h3310)
	) name12538 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_PhyAddrPointer_reg[1]/NET0131 ,
		_w1939_,
		_w3407_,
		_w13888_
	);
	LUT3 #(
		.INIT('h01)
	) name12539 (
		_w8850_,
		_w13888_,
		_w13887_,
		_w13889_
	);
	LUT3 #(
		.INIT('h2f)
	) name12540 (
		_w1933_,
		_w13886_,
		_w13889_,
		_w13890_
	);
	LUT4 #(
		.INIT('h080a)
	) name12541 (
		\P1_Datao_reg[19]/NET0131 ,
		_w1725_,
		_w1797_,
		_w1802_,
		_w13891_
	);
	LUT3 #(
		.INIT('h6c)
	) name12542 (
		\P1_EAX_reg[18]/NET0131 ,
		\P1_EAX_reg[19]/NET0131 ,
		_w9483_,
		_w13892_
	);
	LUT3 #(
		.INIT('he2)
	) name12543 (
		\P1_Datao_reg[19]/NET0131 ,
		_w1859_,
		_w13892_,
		_w13893_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name12544 (
		_w1933_,
		_w12491_,
		_w13891_,
		_w13893_,
		_w13894_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12545 (
		\P1_Datao_reg[19]/NET0131 ,
		\P1_uWord_reg[3]/NET0131 ,
		_w1935_,
		_w9972_,
		_w13895_
	);
	LUT2 #(
		.INIT('hb)
	) name12546 (
		_w13894_,
		_w13895_,
		_w13896_
	);
	LUT4 #(
		.INIT('h0408)
	) name12547 (
		\P1_EAX_reg[23]/NET0131 ,
		_w1797_,
		_w1852_,
		_w9485_,
		_w13897_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name12548 (
		\P1_Datao_reg[23]/NET0131 ,
		_w1858_,
		_w1860_,
		_w13897_,
		_w13898_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12549 (
		\P1_Datao_reg[23]/NET0131 ,
		\P1_uWord_reg[7]/NET0131 ,
		_w1935_,
		_w9972_,
		_w13899_
	);
	LUT3 #(
		.INIT('h2f)
	) name12550 (
		_w1933_,
		_w13898_,
		_w13899_,
		_w13900_
	);
	LUT4 #(
		.INIT('h08aa)
	) name12551 (
		\datao[19]_pad ,
		_w1945_,
		_w2115_,
		_w9978_,
		_w13901_
	);
	LUT2 #(
		.INIT('h8)
	) name12552 (
		\P3_uWord_reg[3]/NET0131 ,
		_w9977_,
		_w13902_
	);
	LUT2 #(
		.INIT('h2)
	) name12553 (
		_w1945_,
		_w2111_,
		_w13903_
	);
	LUT2 #(
		.INIT('h6)
	) name12554 (
		\P3_EAX_reg[19]/NET0131 ,
		_w9538_,
		_w13904_
	);
	LUT4 #(
		.INIT('h0800)
	) name12555 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w13904_,
		_w13905_
	);
	LUT3 #(
		.INIT('h15)
	) name12556 (
		_w13902_,
		_w13903_,
		_w13905_,
		_w13906_
	);
	LUT2 #(
		.INIT('hb)
	) name12557 (
		_w13901_,
		_w13906_,
		_w13907_
	);
	LUT2 #(
		.INIT('h2)
	) name12558 (
		\datao[23]_pad ,
		_w2115_,
		_w13908_
	);
	LUT3 #(
		.INIT('h13)
	) name12559 (
		\P3_EAX_reg[22]/NET0131 ,
		\P3_EAX_reg[23]/NET0131 ,
		_w9539_,
		_w13909_
	);
	LUT4 #(
		.INIT('h0008)
	) name12560 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w9540_,
		_w13910_
	);
	LUT3 #(
		.INIT('h10)
	) name12561 (
		_w2111_,
		_w13909_,
		_w13910_,
		_w13911_
	);
	LUT4 #(
		.INIT('h5f13)
	) name12562 (
		\P3_uWord_reg[7]/NET0131 ,
		\datao[23]_pad ,
		_w9977_,
		_w9978_,
		_w13912_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name12563 (
		_w1945_,
		_w13908_,
		_w13911_,
		_w13912_,
		_w13913_
	);
	LUT3 #(
		.INIT('h6c)
	) name12564 (
		\P2_EAX_reg[18]/NET0131 ,
		\P2_EAX_reg[19]/NET0131 ,
		_w9458_,
		_w13914_
	);
	LUT3 #(
		.INIT('h20)
	) name12565 (
		_w1566_,
		_w1602_,
		_w13914_,
		_w13915_
	);
	LUT4 #(
		.INIT('h0200)
	) name12566 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w13914_,
		_w13916_
	);
	LUT4 #(
		.INIT('h0075)
	) name12567 (
		\P2_Datao_reg[19]/NET0131 ,
		_w1602_,
		_w1616_,
		_w13916_,
		_w13917_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12568 (
		\P2_Datao_reg[19]/NET0131 ,
		\P2_uWord_reg[3]/NET0131 ,
		_w9995_,
		_w9996_,
		_w13918_
	);
	LUT3 #(
		.INIT('h2f)
	) name12569 (
		_w1678_,
		_w13917_,
		_w13918_,
		_w13919_
	);
	LUT3 #(
		.INIT('h6a)
	) name12570 (
		\P2_EAX_reg[23]/NET0131 ,
		_w7781_,
		_w9459_,
		_w13920_
	);
	LUT3 #(
		.INIT('h80)
	) name12571 (
		_w1566_,
		_w1674_,
		_w13920_,
		_w13921_
	);
	LUT4 #(
		.INIT('h0075)
	) name12572 (
		\P2_Datao_reg[23]/NET0131 ,
		_w1602_,
		_w1616_,
		_w13921_,
		_w13922_
	);
	LUT4 #(
		.INIT('h3f15)
	) name12573 (
		\P2_Datao_reg[23]/NET0131 ,
		\P2_uWord_reg[7]/NET0131 ,
		_w9995_,
		_w9996_,
		_w13923_
	);
	LUT3 #(
		.INIT('h2f)
	) name12574 (
		_w1678_,
		_w13922_,
		_w13923_,
		_w13924_
	);
	LUT2 #(
		.INIT('h2)
	) name12575 (
		\P2_uWord_reg[3]/NET0131 ,
		_w7767_,
		_w13925_
	);
	LUT3 #(
		.INIT('h80)
	) name12576 (
		\P2_uWord_reg[3]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13926_
	);
	LUT3 #(
		.INIT('h0d)
	) name12577 (
		_w1606_,
		_w3561_,
		_w13926_,
		_w13927_
	);
	LUT2 #(
		.INIT('h2)
	) name12578 (
		_w1565_,
		_w13927_,
		_w13928_
	);
	LUT4 #(
		.INIT('haa02)
	) name12579 (
		\P2_uWord_reg[3]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w13929_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12580 (
		_w1678_,
		_w13915_,
		_w13928_,
		_w13929_,
		_w13930_
	);
	LUT2 #(
		.INIT('he)
	) name12581 (
		_w13925_,
		_w13930_,
		_w13931_
	);
	LUT2 #(
		.INIT('h2)
	) name12582 (
		\P2_uWord_reg[7]/NET0131 ,
		_w7767_,
		_w13932_
	);
	LUT3 #(
		.INIT('h80)
	) name12583 (
		\P2_uWord_reg[7]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w13933_
	);
	LUT3 #(
		.INIT('h0d)
	) name12584 (
		_w1606_,
		_w2295_,
		_w13933_,
		_w13934_
	);
	LUT2 #(
		.INIT('h2)
	) name12585 (
		_w1565_,
		_w13934_,
		_w13935_
	);
	LUT3 #(
		.INIT('h20)
	) name12586 (
		_w1566_,
		_w1602_,
		_w13920_,
		_w13936_
	);
	LUT4 #(
		.INIT('haa02)
	) name12587 (
		\P2_uWord_reg[7]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w13937_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12588 (
		_w1678_,
		_w13936_,
		_w13935_,
		_w13937_,
		_w13938_
	);
	LUT2 #(
		.INIT('he)
	) name12589 (
		_w13932_,
		_w13938_,
		_w13939_
	);
	LUT2 #(
		.INIT('h2)
	) name12590 (
		\P1_uWord_reg[3]/NET0131 ,
		_w9102_,
		_w13940_
	);
	LUT3 #(
		.INIT('h80)
	) name12591 (
		\P1_uWord_reg[3]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w13941_
	);
	LUT3 #(
		.INIT('h0d)
	) name12592 (
		_w1867_,
		_w3428_,
		_w13941_,
		_w13942_
	);
	LUT2 #(
		.INIT('h2)
	) name12593 (
		_w1795_,
		_w13942_,
		_w13943_
	);
	LUT4 #(
		.INIT('haa02)
	) name12594 (
		\P1_uWord_reg[3]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w13944_
	);
	LUT3 #(
		.INIT('h20)
	) name12595 (
		_w1797_,
		_w1852_,
		_w13892_,
		_w13945_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12596 (
		_w1933_,
		_w13944_,
		_w13943_,
		_w13945_,
		_w13946_
	);
	LUT2 #(
		.INIT('he)
	) name12597 (
		_w13940_,
		_w13946_,
		_w13947_
	);
	LUT2 #(
		.INIT('h2)
	) name12598 (
		\P1_uWord_reg[7]/NET0131 ,
		_w9102_,
		_w13948_
	);
	LUT4 #(
		.INIT('h000d)
	) name12599 (
		\P1_uWord_reg[7]/NET0131 ,
		_w9473_,
		_w12866_,
		_w13897_,
		_w13949_
	);
	LUT3 #(
		.INIT('hce)
	) name12600 (
		_w1933_,
		_w13948_,
		_w13949_,
		_w13950_
	);
	LUT4 #(
		.INIT('hccc4)
	) name12601 (
		_w1945_,
		_w8341_,
		_w8923_,
		_w8924_,
		_w13951_
	);
	LUT3 #(
		.INIT('h40)
	) name12602 (
		\P3_EBX_reg[0]/NET0131 ,
		_w2075_,
		_w2083_,
		_w13952_
	);
	LUT4 #(
		.INIT('h0080)
	) name12603 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2794_,
		_w13953_
	);
	LUT3 #(
		.INIT('ha8)
	) name12604 (
		_w1945_,
		_w13952_,
		_w13953_,
		_w13954_
	);
	LUT3 #(
		.INIT('hf2)
	) name12605 (
		\P3_EBX_reg[0]/NET0131 ,
		_w13951_,
		_w13954_,
		_w13955_
	);
	LUT3 #(
		.INIT('h02)
	) name12606 (
		\P3_EBX_reg[10]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13956_
	);
	LUT4 #(
		.INIT('h0080)
	) name12607 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10039_,
		_w13957_
	);
	LUT3 #(
		.INIT('h08)
	) name12608 (
		_w2075_,
		_w2083_,
		_w8909_,
		_w13958_
	);
	LUT4 #(
		.INIT('h4080)
	) name12609 (
		\P3_EBX_reg[10]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8908_,
		_w13959_
	);
	LUT2 #(
		.INIT('h1)
	) name12610 (
		_w13957_,
		_w13959_,
		_w13960_
	);
	LUT2 #(
		.INIT('h2)
	) name12611 (
		\P3_EBX_reg[10]/NET0131 ,
		_w8341_,
		_w13961_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12612 (
		_w1945_,
		_w13956_,
		_w13960_,
		_w13961_,
		_w13962_
	);
	LUT2 #(
		.INIT('h2)
	) name12613 (
		\P3_EBX_reg[11]/NET0131 ,
		_w8341_,
		_w13963_
	);
	LUT4 #(
		.INIT('haa02)
	) name12614 (
		\P3_EBX_reg[11]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13958_,
		_w13964_
	);
	LUT4 #(
		.INIT('h0080)
	) name12615 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10064_,
		_w13965_
	);
	LUT3 #(
		.INIT('h20)
	) name12616 (
		\P3_EBX_reg[10]/NET0131 ,
		\P3_EBX_reg[11]/NET0131 ,
		_w8908_,
		_w13966_
	);
	LUT3 #(
		.INIT('h80)
	) name12617 (
		_w2075_,
		_w2083_,
		_w13966_,
		_w13967_
	);
	LUT2 #(
		.INIT('h1)
	) name12618 (
		_w13965_,
		_w13967_,
		_w13968_
	);
	LUT4 #(
		.INIT('hecee)
	) name12619 (
		_w1945_,
		_w13963_,
		_w13964_,
		_w13968_,
		_w13969_
	);
	LUT3 #(
		.INIT('h02)
	) name12620 (
		\P3_EBX_reg[12]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13970_
	);
	LUT4 #(
		.INIT('h0080)
	) name12621 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10084_,
		_w13971_
	);
	LUT3 #(
		.INIT('h08)
	) name12622 (
		_w2075_,
		_w2083_,
		_w8911_,
		_w13972_
	);
	LUT4 #(
		.INIT('h4080)
	) name12623 (
		\P3_EBX_reg[12]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8910_,
		_w13973_
	);
	LUT2 #(
		.INIT('h1)
	) name12624 (
		_w13971_,
		_w13973_,
		_w13974_
	);
	LUT2 #(
		.INIT('h2)
	) name12625 (
		\P3_EBX_reg[12]/NET0131 ,
		_w8341_,
		_w13975_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12626 (
		_w1945_,
		_w13970_,
		_w13974_,
		_w13975_,
		_w13976_
	);
	LUT2 #(
		.INIT('h2)
	) name12627 (
		\P3_EBX_reg[13]/NET0131 ,
		_w8341_,
		_w13977_
	);
	LUT4 #(
		.INIT('haa02)
	) name12628 (
		\P3_EBX_reg[13]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13972_,
		_w13978_
	);
	LUT4 #(
		.INIT('h0080)
	) name12629 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10101_,
		_w13979_
	);
	LUT4 #(
		.INIT('h4000)
	) name12630 (
		\P3_EBX_reg[13]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8911_,
		_w13980_
	);
	LUT2 #(
		.INIT('h1)
	) name12631 (
		_w13979_,
		_w13980_,
		_w13981_
	);
	LUT4 #(
		.INIT('hecee)
	) name12632 (
		_w1945_,
		_w13977_,
		_w13978_,
		_w13981_,
		_w13982_
	);
	LUT4 #(
		.INIT('h4080)
	) name12633 (
		\P3_EBX_reg[14]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8912_,
		_w13983_
	);
	LUT4 #(
		.INIT('h0080)
	) name12634 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10118_,
		_w13984_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12635 (
		\P3_EBX_reg[14]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13984_,
		_w13985_
	);
	LUT2 #(
		.INIT('h2)
	) name12636 (
		\P3_EBX_reg[14]/NET0131 ,
		_w8341_,
		_w13986_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12637 (
		_w1945_,
		_w13983_,
		_w13985_,
		_w13986_,
		_w13987_
	);
	LUT4 #(
		.INIT('h4080)
	) name12638 (
		\P3_EBX_reg[15]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8913_,
		_w13988_
	);
	LUT4 #(
		.INIT('h0080)
	) name12639 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10136_,
		_w13989_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12640 (
		\P3_EBX_reg[15]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13989_,
		_w13990_
	);
	LUT2 #(
		.INIT('h2)
	) name12641 (
		\P3_EBX_reg[15]/NET0131 ,
		_w8341_,
		_w13991_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12642 (
		_w1945_,
		_w13988_,
		_w13990_,
		_w13991_,
		_w13992_
	);
	LUT4 #(
		.INIT('h4080)
	) name12643 (
		\P3_EBX_reg[16]/NET0131 ,
		_w2075_,
		_w2083_,
		_w8914_,
		_w13993_
	);
	LUT4 #(
		.INIT('h0080)
	) name12644 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13050_,
		_w13994_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12645 (
		\P3_EBX_reg[16]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13994_,
		_w13995_
	);
	LUT2 #(
		.INIT('h2)
	) name12646 (
		\P3_EBX_reg[16]/NET0131 ,
		_w8341_,
		_w13996_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12647 (
		_w1945_,
		_w13993_,
		_w13995_,
		_w13996_,
		_w13997_
	);
	LUT3 #(
		.INIT('h48)
	) name12648 (
		\P3_EBX_reg[17]/NET0131 ,
		_w2084_,
		_w8915_,
		_w13998_
	);
	LUT4 #(
		.INIT('h0080)
	) name12649 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13070_,
		_w13999_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12650 (
		\P3_EBX_reg[17]/NET0131 ,
		_w8923_,
		_w8924_,
		_w13999_,
		_w14000_
	);
	LUT2 #(
		.INIT('h2)
	) name12651 (
		\P3_EBX_reg[17]/NET0131 ,
		_w8341_,
		_w14001_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12652 (
		_w1945_,
		_w13998_,
		_w14000_,
		_w14001_,
		_w14002_
	);
	LUT2 #(
		.INIT('h2)
	) name12653 (
		\P3_EBX_reg[18]/NET0131 ,
		_w8341_,
		_w14003_
	);
	LUT4 #(
		.INIT('hf250)
	) name12654 (
		_w2084_,
		_w2070_,
		_w8923_,
		_w8916_,
		_w14004_
	);
	LUT4 #(
		.INIT('h0080)
	) name12655 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13096_,
		_w14005_
	);
	LUT3 #(
		.INIT('h40)
	) name12656 (
		\P3_EBX_reg[18]/NET0131 ,
		_w2075_,
		_w2083_,
		_w14006_
	);
	LUT3 #(
		.INIT('h13)
	) name12657 (
		_w8916_,
		_w14005_,
		_w14006_,
		_w14007_
	);
	LUT4 #(
		.INIT('h08cc)
	) name12658 (
		\P3_EBX_reg[18]/NET0131 ,
		_w1945_,
		_w14004_,
		_w14007_,
		_w14008_
	);
	LUT2 #(
		.INIT('he)
	) name12659 (
		_w14003_,
		_w14008_,
		_w14009_
	);
	LUT3 #(
		.INIT('h48)
	) name12660 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2084_,
		_w8917_,
		_w14010_
	);
	LUT4 #(
		.INIT('h0080)
	) name12661 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13113_,
		_w14011_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12662 (
		\P3_EBX_reg[19]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14011_,
		_w14012_
	);
	LUT2 #(
		.INIT('h2)
	) name12663 (
		\P3_EBX_reg[19]/NET0131 ,
		_w8341_,
		_w14013_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12664 (
		_w1945_,
		_w14010_,
		_w14012_,
		_w14013_,
		_w14014_
	);
	LUT3 #(
		.INIT('h02)
	) name12665 (
		\P3_EBX_reg[1]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14015_
	);
	LUT3 #(
		.INIT('h80)
	) name12666 (
		_w2075_,
		_w2083_,
		_w12004_,
		_w14016_
	);
	LUT4 #(
		.INIT('h0080)
	) name12667 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2783_,
		_w14017_
	);
	LUT2 #(
		.INIT('h1)
	) name12668 (
		_w14016_,
		_w14017_,
		_w14018_
	);
	LUT2 #(
		.INIT('h2)
	) name12669 (
		\P3_EBX_reg[1]/NET0131 ,
		_w8341_,
		_w14019_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12670 (
		_w1945_,
		_w14015_,
		_w14018_,
		_w14019_,
		_w14020_
	);
	LUT3 #(
		.INIT('h80)
	) name12671 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		_w8917_,
		_w14021_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12672 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		_w2084_,
		_w8917_,
		_w14022_
	);
	LUT4 #(
		.INIT('h0080)
	) name12673 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13135_,
		_w14023_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12674 (
		\P3_EBX_reg[20]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14023_,
		_w14024_
	);
	LUT2 #(
		.INIT('h2)
	) name12675 (
		\P3_EBX_reg[20]/NET0131 ,
		_w8341_,
		_w14025_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12676 (
		_w1945_,
		_w14022_,
		_w14024_,
		_w14025_,
		_w14026_
	);
	LUT4 #(
		.INIT('h8000)
	) name12677 (
		\P3_EBX_reg[19]/NET0131 ,
		\P3_EBX_reg[20]/NET0131 ,
		\P3_EBX_reg[21]/NET0131 ,
		_w8917_,
		_w14027_
	);
	LUT4 #(
		.INIT('h0080)
	) name12678 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13153_,
		_w14028_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12679 (
		\P3_EBX_reg[21]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14028_,
		_w14029_
	);
	LUT4 #(
		.INIT('hb700)
	) name12680 (
		\P3_EBX_reg[21]/NET0131 ,
		_w2084_,
		_w14021_,
		_w14029_,
		_w14030_
	);
	LUT2 #(
		.INIT('h2)
	) name12681 (
		\P3_EBX_reg[21]/NET0131 ,
		_w8341_,
		_w14031_
	);
	LUT3 #(
		.INIT('hf2)
	) name12682 (
		_w1945_,
		_w14030_,
		_w14031_,
		_w14032_
	);
	LUT4 #(
		.INIT('h0080)
	) name12683 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13176_,
		_w14033_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12684 (
		\P3_EBX_reg[22]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14033_,
		_w14034_
	);
	LUT4 #(
		.INIT('hb700)
	) name12685 (
		\P3_EBX_reg[22]/NET0131 ,
		_w2084_,
		_w14027_,
		_w14034_,
		_w14035_
	);
	LUT2 #(
		.INIT('h2)
	) name12686 (
		\P3_EBX_reg[22]/NET0131 ,
		_w8341_,
		_w14036_
	);
	LUT3 #(
		.INIT('hf2)
	) name12687 (
		_w1945_,
		_w14035_,
		_w14036_,
		_w14037_
	);
	LUT2 #(
		.INIT('h2)
	) name12688 (
		\P3_EBX_reg[23]/NET0131 ,
		_w8341_,
		_w14038_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name12689 (
		\P3_EBX_reg[19]/NET0131 ,
		_w2084_,
		_w8917_,
		_w8918_,
		_w14039_
	);
	LUT4 #(
		.INIT('hec00)
	) name12690 (
		\P3_EBX_reg[22]/NET0131 ,
		\P3_EBX_reg[23]/NET0131 ,
		_w14027_,
		_w14039_,
		_w14040_
	);
	LUT4 #(
		.INIT('h8000)
	) name12691 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13189_,
		_w14041_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12692 (
		\P3_EBX_reg[23]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14041_,
		_w14042_
	);
	LUT4 #(
		.INIT('hecee)
	) name12693 (
		_w1945_,
		_w14038_,
		_w14040_,
		_w14042_,
		_w14043_
	);
	LUT4 #(
		.INIT('h8000)
	) name12694 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w13201_,
		_w14044_
	);
	LUT4 #(
		.INIT('h00fd)
	) name12695 (
		\P3_EBX_reg[24]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14044_,
		_w14045_
	);
	LUT4 #(
		.INIT('hb700)
	) name12696 (
		\P3_EBX_reg[24]/NET0131 ,
		_w2084_,
		_w8919_,
		_w14045_,
		_w14046_
	);
	LUT2 #(
		.INIT('h2)
	) name12697 (
		\P3_EBX_reg[24]/NET0131 ,
		_w8341_,
		_w14047_
	);
	LUT3 #(
		.INIT('hf2)
	) name12698 (
		_w1945_,
		_w14046_,
		_w14047_,
		_w14048_
	);
	LUT2 #(
		.INIT('h2)
	) name12699 (
		\P3_EBX_reg[28]/NET0131 ,
		_w8341_,
		_w14049_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name12700 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2084_,
		_w8925_,
		_w10254_,
		_w14050_
	);
	LUT2 #(
		.INIT('h8)
	) name12701 (
		_w8923_,
		_w13209_,
		_w14051_
	);
	LUT3 #(
		.INIT('h40)
	) name12702 (
		\P3_EBX_reg[28]/NET0131 ,
		_w2075_,
		_w2083_,
		_w14052_
	);
	LUT3 #(
		.INIT('h13)
	) name12703 (
		_w10254_,
		_w14051_,
		_w14052_,
		_w14053_
	);
	LUT4 #(
		.INIT('hecee)
	) name12704 (
		_w1945_,
		_w14049_,
		_w14050_,
		_w14053_,
		_w14054_
	);
	LUT3 #(
		.INIT('h02)
	) name12705 (
		\P3_EBX_reg[2]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14055_
	);
	LUT4 #(
		.INIT('h0080)
	) name12706 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2769_,
		_w14056_
	);
	LUT3 #(
		.INIT('h78)
	) name12707 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		_w14057_
	);
	LUT3 #(
		.INIT('h80)
	) name12708 (
		_w2075_,
		_w2083_,
		_w14057_,
		_w14058_
	);
	LUT2 #(
		.INIT('h1)
	) name12709 (
		_w14056_,
		_w14058_,
		_w14059_
	);
	LUT2 #(
		.INIT('h2)
	) name12710 (
		\P3_EBX_reg[2]/NET0131 ,
		_w8341_,
		_w14060_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12711 (
		_w1945_,
		_w14055_,
		_w14059_,
		_w14060_,
		_w14061_
	);
	LUT3 #(
		.INIT('h02)
	) name12712 (
		\P3_EBX_reg[3]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14062_
	);
	LUT4 #(
		.INIT('h0080)
	) name12713 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2809_,
		_w14063_
	);
	LUT4 #(
		.INIT('h7f80)
	) name12714 (
		\P3_EBX_reg[0]/NET0131 ,
		\P3_EBX_reg[1]/NET0131 ,
		\P3_EBX_reg[2]/NET0131 ,
		\P3_EBX_reg[3]/NET0131 ,
		_w14064_
	);
	LUT3 #(
		.INIT('h80)
	) name12715 (
		_w2075_,
		_w2083_,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h1)
	) name12716 (
		_w14063_,
		_w14065_,
		_w14066_
	);
	LUT2 #(
		.INIT('h2)
	) name12717 (
		\P3_EBX_reg[3]/NET0131 ,
		_w8341_,
		_w14067_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12718 (
		_w1945_,
		_w14062_,
		_w14066_,
		_w14067_,
		_w14068_
	);
	LUT3 #(
		.INIT('h02)
	) name12719 (
		\P3_EBX_reg[4]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14069_
	);
	LUT4 #(
		.INIT('h0080)
	) name12720 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2824_,
		_w14070_
	);
	LUT2 #(
		.INIT('h6)
	) name12721 (
		\P3_EBX_reg[4]/NET0131 ,
		_w8906_,
		_w14071_
	);
	LUT3 #(
		.INIT('h80)
	) name12722 (
		_w2075_,
		_w2083_,
		_w14071_,
		_w14072_
	);
	LUT2 #(
		.INIT('h1)
	) name12723 (
		_w14070_,
		_w14072_,
		_w14073_
	);
	LUT2 #(
		.INIT('h2)
	) name12724 (
		\P3_EBX_reg[4]/NET0131 ,
		_w8341_,
		_w14074_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12725 (
		_w1945_,
		_w14069_,
		_w14073_,
		_w14074_,
		_w14075_
	);
	LUT3 #(
		.INIT('h02)
	) name12726 (
		\P3_EBX_reg[5]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14076_
	);
	LUT4 #(
		.INIT('h0080)
	) name12727 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2855_,
		_w14077_
	);
	LUT3 #(
		.INIT('h6c)
	) name12728 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		_w8906_,
		_w14078_
	);
	LUT3 #(
		.INIT('h80)
	) name12729 (
		_w2075_,
		_w2083_,
		_w14078_,
		_w14079_
	);
	LUT2 #(
		.INIT('h1)
	) name12730 (
		_w14077_,
		_w14079_,
		_w14080_
	);
	LUT2 #(
		.INIT('h2)
	) name12731 (
		\P3_EBX_reg[5]/NET0131 ,
		_w8341_,
		_w14081_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12732 (
		_w1945_,
		_w14076_,
		_w14080_,
		_w14081_,
		_w14082_
	);
	LUT3 #(
		.INIT('h02)
	) name12733 (
		\P3_EBX_reg[6]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14083_
	);
	LUT4 #(
		.INIT('h0080)
	) name12734 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2842_,
		_w14084_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12735 (
		\P3_EBX_reg[4]/NET0131 ,
		\P3_EBX_reg[5]/NET0131 ,
		\P3_EBX_reg[6]/NET0131 ,
		_w8906_,
		_w14085_
	);
	LUT3 #(
		.INIT('h80)
	) name12736 (
		_w2075_,
		_w2083_,
		_w14085_,
		_w14086_
	);
	LUT2 #(
		.INIT('h1)
	) name12737 (
		_w14084_,
		_w14086_,
		_w14087_
	);
	LUT2 #(
		.INIT('h2)
	) name12738 (
		\P3_EBX_reg[6]/NET0131 ,
		_w8341_,
		_w14088_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12739 (
		_w1945_,
		_w14083_,
		_w14087_,
		_w14088_,
		_w14089_
	);
	LUT3 #(
		.INIT('h02)
	) name12740 (
		\P3_EBX_reg[7]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14090_
	);
	LUT4 #(
		.INIT('h0080)
	) name12741 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w2755_,
		_w14091_
	);
	LUT2 #(
		.INIT('h6)
	) name12742 (
		\P3_EBX_reg[7]/NET0131 ,
		_w8907_,
		_w14092_
	);
	LUT3 #(
		.INIT('h80)
	) name12743 (
		_w2075_,
		_w2083_,
		_w14092_,
		_w14093_
	);
	LUT2 #(
		.INIT('h1)
	) name12744 (
		_w14091_,
		_w14093_,
		_w14094_
	);
	LUT2 #(
		.INIT('h2)
	) name12745 (
		\P3_EBX_reg[7]/NET0131 ,
		_w8341_,
		_w14095_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12746 (
		_w1945_,
		_w14090_,
		_w14094_,
		_w14095_,
		_w14096_
	);
	LUT3 #(
		.INIT('h02)
	) name12747 (
		\P3_EBX_reg[8]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14097_
	);
	LUT4 #(
		.INIT('h0080)
	) name12748 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10221_,
		_w14098_
	);
	LUT3 #(
		.INIT('h6c)
	) name12749 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		_w8907_,
		_w14099_
	);
	LUT3 #(
		.INIT('h80)
	) name12750 (
		_w2075_,
		_w2083_,
		_w14099_,
		_w14100_
	);
	LUT2 #(
		.INIT('h1)
	) name12751 (
		_w14098_,
		_w14100_,
		_w14101_
	);
	LUT2 #(
		.INIT('h2)
	) name12752 (
		\P3_EBX_reg[8]/NET0131 ,
		_w8341_,
		_w14102_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12753 (
		_w1945_,
		_w14097_,
		_w14101_,
		_w14102_,
		_w14103_
	);
	LUT3 #(
		.INIT('h02)
	) name12754 (
		\P3_EBX_reg[9]/NET0131 ,
		_w8923_,
		_w8924_,
		_w14104_
	);
	LUT4 #(
		.INIT('h0080)
	) name12755 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w10238_,
		_w14105_
	);
	LUT4 #(
		.INIT('h78f0)
	) name12756 (
		\P3_EBX_reg[7]/NET0131 ,
		\P3_EBX_reg[8]/NET0131 ,
		\P3_EBX_reg[9]/NET0131 ,
		_w8907_,
		_w14106_
	);
	LUT3 #(
		.INIT('h80)
	) name12757 (
		_w2075_,
		_w2083_,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h1)
	) name12758 (
		_w14105_,
		_w14107_,
		_w14108_
	);
	LUT2 #(
		.INIT('h2)
	) name12759 (
		\P3_EBX_reg[9]/NET0131 ,
		_w8341_,
		_w14109_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12760 (
		_w1945_,
		_w14104_,
		_w14108_,
		_w14109_,
		_w14110_
	);
	LUT4 #(
		.INIT('h3700)
	) name12761 (
		_w1863_,
		_w1933_,
		_w8992_,
		_w9102_,
		_w14111_
	);
	LUT3 #(
		.INIT('h40)
	) name12762 (
		\P1_EBX_reg[0]/NET0131 ,
		_w1826_,
		_w1828_,
		_w14112_
	);
	LUT3 #(
		.INIT('h80)
	) name12763 (
		_w1750_,
		_w1813_,
		_w13402_,
		_w14113_
	);
	LUT3 #(
		.INIT('ha8)
	) name12764 (
		_w1933_,
		_w14112_,
		_w14113_,
		_w14114_
	);
	LUT3 #(
		.INIT('hf2)
	) name12765 (
		\P1_EBX_reg[0]/NET0131 ,
		_w14111_,
		_w14114_,
		_w14115_
	);
	LUT3 #(
		.INIT('ha8)
	) name12766 (
		\P1_EBX_reg[10]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14116_
	);
	LUT3 #(
		.INIT('h80)
	) name12767 (
		_w1750_,
		_w1813_,
		_w10439_,
		_w14117_
	);
	LUT2 #(
		.INIT('h6)
	) name12768 (
		\P1_EBX_reg[10]/NET0131 ,
		_w8975_,
		_w14118_
	);
	LUT3 #(
		.INIT('h80)
	) name12769 (
		_w1826_,
		_w1828_,
		_w14118_,
		_w14119_
	);
	LUT2 #(
		.INIT('h1)
	) name12770 (
		_w14117_,
		_w14119_,
		_w14120_
	);
	LUT2 #(
		.INIT('h2)
	) name12771 (
		\P1_EBX_reg[10]/NET0131 ,
		_w9102_,
		_w14121_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12772 (
		_w1933_,
		_w14116_,
		_w14120_,
		_w14121_,
		_w14122_
	);
	LUT3 #(
		.INIT('ha8)
	) name12773 (
		\P1_EBX_reg[11]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14123_
	);
	LUT3 #(
		.INIT('h80)
	) name12774 (
		_w1750_,
		_w1813_,
		_w10519_,
		_w14124_
	);
	LUT3 #(
		.INIT('h08)
	) name12775 (
		_w1826_,
		_w1828_,
		_w8977_,
		_w14125_
	);
	LUT4 #(
		.INIT('h4080)
	) name12776 (
		\P1_EBX_reg[11]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8976_,
		_w14126_
	);
	LUT2 #(
		.INIT('h1)
	) name12777 (
		_w14124_,
		_w14126_,
		_w14127_
	);
	LUT2 #(
		.INIT('h2)
	) name12778 (
		\P1_EBX_reg[11]/NET0131 ,
		_w9102_,
		_w14128_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12779 (
		_w1933_,
		_w14123_,
		_w14127_,
		_w14128_,
		_w14129_
	);
	LUT2 #(
		.INIT('h2)
	) name12780 (
		\P1_EBX_reg[12]/NET0131 ,
		_w9102_,
		_w14130_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12781 (
		\P1_EBX_reg[12]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14125_,
		_w14131_
	);
	LUT3 #(
		.INIT('h80)
	) name12782 (
		_w1750_,
		_w1813_,
		_w10589_,
		_w14132_
	);
	LUT4 #(
		.INIT('h4000)
	) name12783 (
		\P1_EBX_reg[12]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8977_,
		_w14133_
	);
	LUT2 #(
		.INIT('h1)
	) name12784 (
		_w14132_,
		_w14133_,
		_w14134_
	);
	LUT4 #(
		.INIT('hecee)
	) name12785 (
		_w1933_,
		_w14130_,
		_w14131_,
		_w14134_,
		_w14135_
	);
	LUT3 #(
		.INIT('h08)
	) name12786 (
		_w1826_,
		_w1828_,
		_w8979_,
		_w14136_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12787 (
		\P1_EBX_reg[14]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14136_,
		_w14137_
	);
	LUT3 #(
		.INIT('h80)
	) name12788 (
		_w1750_,
		_w1813_,
		_w10551_,
		_w14138_
	);
	LUT4 #(
		.INIT('h4000)
	) name12789 (
		\P1_EBX_reg[14]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8979_,
		_w14139_
	);
	LUT2 #(
		.INIT('h1)
	) name12790 (
		_w14138_,
		_w14139_,
		_w14140_
	);
	LUT2 #(
		.INIT('h2)
	) name12791 (
		\P1_EBX_reg[14]/NET0131 ,
		_w9102_,
		_w14141_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12792 (
		_w1933_,
		_w14137_,
		_w14140_,
		_w14141_,
		_w14142_
	);
	LUT4 #(
		.INIT('h4080)
	) name12793 (
		\P1_EBX_reg[13]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8978_,
		_w14143_
	);
	LUT3 #(
		.INIT('h80)
	) name12794 (
		_w1750_,
		_w1813_,
		_w10569_,
		_w14144_
	);
	LUT4 #(
		.INIT('h0057)
	) name12795 (
		\P1_EBX_reg[13]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14144_,
		_w14145_
	);
	LUT2 #(
		.INIT('h2)
	) name12796 (
		\P1_EBX_reg[13]/NET0131 ,
		_w9102_,
		_w14146_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12797 (
		_w1933_,
		_w14143_,
		_w14145_,
		_w14146_,
		_w14147_
	);
	LUT4 #(
		.INIT('h4080)
	) name12798 (
		\P1_EBX_reg[15]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8980_,
		_w14148_
	);
	LUT3 #(
		.INIT('h80)
	) name12799 (
		_w1750_,
		_w1813_,
		_w9734_,
		_w14149_
	);
	LUT4 #(
		.INIT('h0057)
	) name12800 (
		\P1_EBX_reg[15]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14149_,
		_w14150_
	);
	LUT2 #(
		.INIT('h2)
	) name12801 (
		\P1_EBX_reg[15]/NET0131 ,
		_w9102_,
		_w14151_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12802 (
		_w1933_,
		_w14148_,
		_w14150_,
		_w14151_,
		_w14152_
	);
	LUT4 #(
		.INIT('h4080)
	) name12803 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1826_,
		_w1828_,
		_w8981_,
		_w14153_
	);
	LUT3 #(
		.INIT('h80)
	) name12804 (
		_w1750_,
		_w1813_,
		_w13444_,
		_w14154_
	);
	LUT4 #(
		.INIT('h0057)
	) name12805 (
		\P1_EBX_reg[16]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14154_,
		_w14155_
	);
	LUT2 #(
		.INIT('h2)
	) name12806 (
		\P1_EBX_reg[16]/NET0131 ,
		_w9102_,
		_w14156_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12807 (
		_w1933_,
		_w14153_,
		_w14155_,
		_w14156_,
		_w14157_
	);
	LUT3 #(
		.INIT('h48)
	) name12808 (
		\P1_EBX_reg[17]/NET0131 ,
		_w1829_,
		_w8982_,
		_w14158_
	);
	LUT3 #(
		.INIT('h80)
	) name12809 (
		_w1750_,
		_w1813_,
		_w13464_,
		_w14159_
	);
	LUT4 #(
		.INIT('h0057)
	) name12810 (
		\P1_EBX_reg[17]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h2)
	) name12811 (
		\P1_EBX_reg[17]/NET0131 ,
		_w9102_,
		_w14161_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12812 (
		_w1933_,
		_w14158_,
		_w14160_,
		_w14161_,
		_w14162_
	);
	LUT3 #(
		.INIT('h4c)
	) name12813 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1829_,
		_w8984_,
		_w14163_
	);
	LUT3 #(
		.INIT('h48)
	) name12814 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1829_,
		_w8984_,
		_w14164_
	);
	LUT3 #(
		.INIT('h80)
	) name12815 (
		_w1750_,
		_w1813_,
		_w13488_,
		_w14165_
	);
	LUT4 #(
		.INIT('h0057)
	) name12816 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14165_,
		_w14166_
	);
	LUT2 #(
		.INIT('h2)
	) name12817 (
		\P1_EBX_reg[19]/NET0131 ,
		_w9102_,
		_w14167_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12818 (
		_w1933_,
		_w14164_,
		_w14166_,
		_w14167_,
		_w14168_
	);
	LUT3 #(
		.INIT('h48)
	) name12819 (
		\P1_EBX_reg[18]/NET0131 ,
		_w1829_,
		_w8983_,
		_w14169_
	);
	LUT3 #(
		.INIT('h80)
	) name12820 (
		_w1750_,
		_w1813_,
		_w13509_,
		_w14170_
	);
	LUT4 #(
		.INIT('h0057)
	) name12821 (
		\P1_EBX_reg[18]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14170_,
		_w14171_
	);
	LUT2 #(
		.INIT('h2)
	) name12822 (
		\P1_EBX_reg[18]/NET0131 ,
		_w9102_,
		_w14172_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12823 (
		_w1933_,
		_w14169_,
		_w14171_,
		_w14172_,
		_w14173_
	);
	LUT3 #(
		.INIT('ha8)
	) name12824 (
		\P1_EBX_reg[1]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14174_
	);
	LUT3 #(
		.INIT('h80)
	) name12825 (
		_w1750_,
		_w1813_,
		_w10604_,
		_w14175_
	);
	LUT3 #(
		.INIT('h80)
	) name12826 (
		_w1826_,
		_w1828_,
		_w10947_,
		_w14176_
	);
	LUT2 #(
		.INIT('h1)
	) name12827 (
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT2 #(
		.INIT('h2)
	) name12828 (
		\P1_EBX_reg[1]/NET0131 ,
		_w9102_,
		_w14178_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12829 (
		_w1933_,
		_w14174_,
		_w14177_,
		_w14178_,
		_w14179_
	);
	LUT2 #(
		.INIT('h2)
	) name12830 (
		\P1_EBX_reg[20]/NET0131 ,
		_w9102_,
		_w14180_
	);
	LUT3 #(
		.INIT('h80)
	) name12831 (
		_w1750_,
		_w1813_,
		_w13530_,
		_w14181_
	);
	LUT3 #(
		.INIT('h40)
	) name12832 (
		\P1_EBX_reg[20]/NET0131 ,
		_w1826_,
		_w1828_,
		_w14182_
	);
	LUT4 #(
		.INIT('h070f)
	) name12833 (
		\P1_EBX_reg[19]/NET0131 ,
		_w8984_,
		_w14181_,
		_w14182_,
		_w14183_
	);
	LUT4 #(
		.INIT('h5d00)
	) name12834 (
		\P1_EBX_reg[20]/NET0131 ,
		_w8993_,
		_w14163_,
		_w14183_,
		_w14184_
	);
	LUT3 #(
		.INIT('hce)
	) name12835 (
		_w1933_,
		_w14180_,
		_w14184_,
		_w14185_
	);
	LUT3 #(
		.INIT('h80)
	) name12836 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		_w8984_,
		_w14186_
	);
	LUT4 #(
		.INIT('h8000)
	) name12837 (
		\P1_EBX_reg[19]/NET0131 ,
		\P1_EBX_reg[20]/NET0131 ,
		\P1_EBX_reg[21]/NET0131 ,
		_w8984_,
		_w14187_
	);
	LUT3 #(
		.INIT('h80)
	) name12838 (
		_w1750_,
		_w1813_,
		_w13549_,
		_w14188_
	);
	LUT4 #(
		.INIT('h0057)
	) name12839 (
		\P1_EBX_reg[21]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14188_,
		_w14189_
	);
	LUT4 #(
		.INIT('hb700)
	) name12840 (
		\P1_EBX_reg[21]/NET0131 ,
		_w1829_,
		_w14186_,
		_w14189_,
		_w14190_
	);
	LUT2 #(
		.INIT('h2)
	) name12841 (
		\P1_EBX_reg[21]/NET0131 ,
		_w9102_,
		_w14191_
	);
	LUT3 #(
		.INIT('hf2)
	) name12842 (
		_w1933_,
		_w14190_,
		_w14191_,
		_w14192_
	);
	LUT3 #(
		.INIT('h80)
	) name12843 (
		_w1750_,
		_w1813_,
		_w13566_,
		_w14193_
	);
	LUT4 #(
		.INIT('h0057)
	) name12844 (
		\P1_EBX_reg[22]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14193_,
		_w14194_
	);
	LUT4 #(
		.INIT('hb700)
	) name12845 (
		\P1_EBX_reg[22]/NET0131 ,
		_w1829_,
		_w14187_,
		_w14194_,
		_w14195_
	);
	LUT2 #(
		.INIT('h2)
	) name12846 (
		\P1_EBX_reg[22]/NET0131 ,
		_w9102_,
		_w14196_
	);
	LUT3 #(
		.INIT('hf2)
	) name12847 (
		_w1933_,
		_w14195_,
		_w14196_,
		_w14197_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name12848 (
		\P1_EBX_reg[19]/NET0131 ,
		_w1829_,
		_w8984_,
		_w8985_,
		_w14198_
	);
	LUT4 #(
		.INIT('hec00)
	) name12849 (
		\P1_EBX_reg[22]/NET0131 ,
		\P1_EBX_reg[23]/NET0131 ,
		_w14187_,
		_w14198_,
		_w14199_
	);
	LUT3 #(
		.INIT('h80)
	) name12850 (
		_w1750_,
		_w1813_,
		_w12864_,
		_w14200_
	);
	LUT4 #(
		.INIT('h0057)
	) name12851 (
		\P1_EBX_reg[23]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14200_,
		_w14201_
	);
	LUT2 #(
		.INIT('h2)
	) name12852 (
		\P1_EBX_reg[23]/NET0131 ,
		_w9102_,
		_w14202_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12853 (
		_w1933_,
		_w14199_,
		_w14201_,
		_w14202_,
		_w14203_
	);
	LUT3 #(
		.INIT('h80)
	) name12854 (
		_w1750_,
		_w1813_,
		_w12901_,
		_w14204_
	);
	LUT4 #(
		.INIT('h0057)
	) name12855 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14204_,
		_w14205_
	);
	LUT4 #(
		.INIT('hb700)
	) name12856 (
		\P1_EBX_reg[24]/NET0131 ,
		_w1829_,
		_w8986_,
		_w14205_,
		_w14206_
	);
	LUT2 #(
		.INIT('h2)
	) name12857 (
		\P1_EBX_reg[24]/NET0131 ,
		_w9102_,
		_w14207_
	);
	LUT3 #(
		.INIT('hf2)
	) name12858 (
		_w1933_,
		_w14206_,
		_w14207_,
		_w14208_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12859 (
		\P2_EBX_reg[0]/NET0131 ,
		_w1678_,
		_w7767_,
		_w8961_,
		_w14209_
	);
	LUT2 #(
		.INIT('h4)
	) name12860 (
		\P2_EBX_reg[0]/NET0131 ,
		_w1578_,
		_w14210_
	);
	LUT3 #(
		.INIT('h80)
	) name12861 (
		_w1503_,
		_w1549_,
		_w10248_,
		_w14211_
	);
	LUT3 #(
		.INIT('ha8)
	) name12862 (
		_w1678_,
		_w14210_,
		_w14211_,
		_w14212_
	);
	LUT2 #(
		.INIT('he)
	) name12863 (
		_w14209_,
		_w14212_,
		_w14213_
	);
	LUT3 #(
		.INIT('h80)
	) name12864 (
		_w1503_,
		_w1549_,
		_w10289_,
		_w14214_
	);
	LUT2 #(
		.INIT('h2)
	) name12865 (
		_w1578_,
		_w8947_,
		_w14215_
	);
	LUT3 #(
		.INIT('h48)
	) name12866 (
		\P2_EBX_reg[10]/NET0131 ,
		_w1578_,
		_w8946_,
		_w14216_
	);
	LUT4 #(
		.INIT('h000d)
	) name12867 (
		\P2_EBX_reg[10]/NET0131 ,
		_w8961_,
		_w14214_,
		_w14216_,
		_w14217_
	);
	LUT2 #(
		.INIT('h2)
	) name12868 (
		\P2_EBX_reg[10]/NET0131 ,
		_w7767_,
		_w14218_
	);
	LUT3 #(
		.INIT('hf2)
	) name12869 (
		_w1678_,
		_w14217_,
		_w14218_,
		_w14219_
	);
	LUT3 #(
		.INIT('ha2)
	) name12870 (
		\P2_EBX_reg[11]/NET0131 ,
		_w8961_,
		_w14215_,
		_w14220_
	);
	LUT3 #(
		.INIT('h80)
	) name12871 (
		_w1503_,
		_w1549_,
		_w10306_,
		_w14221_
	);
	LUT3 #(
		.INIT('h40)
	) name12872 (
		\P2_EBX_reg[11]/NET0131 ,
		_w1578_,
		_w8947_,
		_w14222_
	);
	LUT2 #(
		.INIT('h1)
	) name12873 (
		_w14221_,
		_w14222_,
		_w14223_
	);
	LUT2 #(
		.INIT('h2)
	) name12874 (
		\P2_EBX_reg[11]/NET0131 ,
		_w7767_,
		_w14224_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12875 (
		_w1678_,
		_w14220_,
		_w14223_,
		_w14224_,
		_w14225_
	);
	LUT2 #(
		.INIT('h2)
	) name12876 (
		_w1578_,
		_w8949_,
		_w14226_
	);
	LUT3 #(
		.INIT('h48)
	) name12877 (
		\P2_EBX_reg[12]/NET0131 ,
		_w1578_,
		_w8948_,
		_w14227_
	);
	LUT3 #(
		.INIT('h80)
	) name12878 (
		_w1503_,
		_w1549_,
		_w10326_,
		_w14228_
	);
	LUT4 #(
		.INIT('h000d)
	) name12879 (
		\P2_EBX_reg[12]/NET0131 ,
		_w8961_,
		_w14228_,
		_w14227_,
		_w14229_
	);
	LUT2 #(
		.INIT('h2)
	) name12880 (
		\P2_EBX_reg[12]/NET0131 ,
		_w7767_,
		_w14230_
	);
	LUT3 #(
		.INIT('hf2)
	) name12881 (
		_w1678_,
		_w14229_,
		_w14230_,
		_w14231_
	);
	LUT3 #(
		.INIT('ha2)
	) name12882 (
		\P2_EBX_reg[13]/NET0131 ,
		_w8961_,
		_w14226_,
		_w14232_
	);
	LUT3 #(
		.INIT('h80)
	) name12883 (
		_w1503_,
		_w1549_,
		_w10371_,
		_w14233_
	);
	LUT3 #(
		.INIT('h40)
	) name12884 (
		\P2_EBX_reg[13]/NET0131 ,
		_w1578_,
		_w8949_,
		_w14234_
	);
	LUT2 #(
		.INIT('h1)
	) name12885 (
		_w14233_,
		_w14234_,
		_w14235_
	);
	LUT2 #(
		.INIT('h2)
	) name12886 (
		\P2_EBX_reg[13]/NET0131 ,
		_w7767_,
		_w14236_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12887 (
		_w1678_,
		_w14232_,
		_w14235_,
		_w14236_,
		_w14237_
	);
	LUT3 #(
		.INIT('h13)
	) name12888 (
		\P2_EBX_reg[13]/NET0131 ,
		\P2_EBX_reg[14]/NET0131 ,
		_w8949_,
		_w14238_
	);
	LUT3 #(
		.INIT('h02)
	) name12889 (
		_w1578_,
		_w8951_,
		_w14238_,
		_w14239_
	);
	LUT3 #(
		.INIT('h80)
	) name12890 (
		_w1503_,
		_w1549_,
		_w10390_,
		_w14240_
	);
	LUT4 #(
		.INIT('h000d)
	) name12891 (
		\P2_EBX_reg[14]/NET0131 ,
		_w8961_,
		_w14240_,
		_w14239_,
		_w14241_
	);
	LUT2 #(
		.INIT('h2)
	) name12892 (
		\P2_EBX_reg[14]/NET0131 ,
		_w7767_,
		_w14242_
	);
	LUT3 #(
		.INIT('hf2)
	) name12893 (
		_w1678_,
		_w14241_,
		_w14242_,
		_w14243_
	);
	LUT3 #(
		.INIT('h48)
	) name12894 (
		\P2_EBX_reg[15]/NET0131 ,
		_w1578_,
		_w8951_,
		_w14244_
	);
	LUT3 #(
		.INIT('h80)
	) name12895 (
		_w1503_,
		_w1549_,
		_w9688_,
		_w14245_
	);
	LUT4 #(
		.INIT('h000d)
	) name12896 (
		\P2_EBX_reg[15]/NET0131 ,
		_w8961_,
		_w14245_,
		_w14244_,
		_w14246_
	);
	LUT2 #(
		.INIT('h2)
	) name12897 (
		\P2_EBX_reg[15]/NET0131 ,
		_w7767_,
		_w14247_
	);
	LUT3 #(
		.INIT('hf2)
	) name12898 (
		_w1678_,
		_w14246_,
		_w14247_,
		_w14248_
	);
	LUT3 #(
		.INIT('h48)
	) name12899 (
		\P2_EBX_reg[16]/NET0131 ,
		_w1578_,
		_w8952_,
		_w14249_
	);
	LUT3 #(
		.INIT('h80)
	) name12900 (
		_w1503_,
		_w1549_,
		_w13232_,
		_w14250_
	);
	LUT4 #(
		.INIT('h000d)
	) name12901 (
		\P2_EBX_reg[16]/NET0131 ,
		_w8961_,
		_w14250_,
		_w14249_,
		_w14251_
	);
	LUT2 #(
		.INIT('h2)
	) name12902 (
		\P2_EBX_reg[16]/NET0131 ,
		_w7767_,
		_w14252_
	);
	LUT3 #(
		.INIT('hf2)
	) name12903 (
		_w1678_,
		_w14251_,
		_w14252_,
		_w14253_
	);
	LUT2 #(
		.INIT('h2)
	) name12904 (
		\P1_EBX_reg[28]/NET0131 ,
		_w9102_,
		_w14254_
	);
	LUT4 #(
		.INIT('h8000)
	) name12905 (
		\P1_EBX_reg[25]/NET0131 ,
		\P1_EBX_reg[26]/NET0131 ,
		\P1_EBX_reg[27]/NET0131 ,
		_w8987_,
		_w14255_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name12906 (
		\P1_EBX_reg[28]/NET0131 ,
		_w1829_,
		_w8993_,
		_w14255_,
		_w14256_
	);
	LUT2 #(
		.INIT('h8)
	) name12907 (
		_w1814_,
		_w13021_,
		_w14257_
	);
	LUT3 #(
		.INIT('h40)
	) name12908 (
		\P1_EBX_reg[28]/NET0131 ,
		_w1826_,
		_w1828_,
		_w14258_
	);
	LUT3 #(
		.INIT('h13)
	) name12909 (
		_w14255_,
		_w14257_,
		_w14258_,
		_w14259_
	);
	LUT4 #(
		.INIT('hecee)
	) name12910 (
		_w1933_,
		_w14254_,
		_w14256_,
		_w14259_,
		_w14260_
	);
	LUT3 #(
		.INIT('h4c)
	) name12911 (
		\P2_EBX_reg[17]/NET0131 ,
		_w1578_,
		_w8953_,
		_w14261_
	);
	LUT3 #(
		.INIT('h48)
	) name12912 (
		\P2_EBX_reg[17]/NET0131 ,
		_w1578_,
		_w8953_,
		_w14262_
	);
	LUT3 #(
		.INIT('h80)
	) name12913 (
		_w1503_,
		_w1549_,
		_w13257_,
		_w14263_
	);
	LUT4 #(
		.INIT('h000d)
	) name12914 (
		\P2_EBX_reg[17]/NET0131 ,
		_w8961_,
		_w14263_,
		_w14262_,
		_w14264_
	);
	LUT2 #(
		.INIT('h2)
	) name12915 (
		\P2_EBX_reg[17]/NET0131 ,
		_w7767_,
		_w14265_
	);
	LUT3 #(
		.INIT('hf2)
	) name12916 (
		_w1678_,
		_w14264_,
		_w14265_,
		_w14266_
	);
	LUT2 #(
		.INIT('h2)
	) name12917 (
		\P2_EBX_reg[18]/NET0131 ,
		_w7767_,
		_w14267_
	);
	LUT3 #(
		.INIT('ha2)
	) name12918 (
		\P2_EBX_reg[18]/NET0131 ,
		_w8961_,
		_w14261_,
		_w14268_
	);
	LUT3 #(
		.INIT('h80)
	) name12919 (
		_w1503_,
		_w1549_,
		_w13279_,
		_w14269_
	);
	LUT4 #(
		.INIT('h2000)
	) name12920 (
		\P2_EBX_reg[17]/NET0131 ,
		\P2_EBX_reg[18]/NET0131 ,
		_w1578_,
		_w8953_,
		_w14270_
	);
	LUT2 #(
		.INIT('h1)
	) name12921 (
		_w14269_,
		_w14270_,
		_w14271_
	);
	LUT4 #(
		.INIT('hecee)
	) name12922 (
		_w1678_,
		_w14267_,
		_w14268_,
		_w14271_,
		_w14272_
	);
	LUT4 #(
		.INIT('h4888)
	) name12923 (
		\P2_EBX_reg[19]/NET0131 ,
		_w1578_,
		_w8953_,
		_w8954_,
		_w14273_
	);
	LUT3 #(
		.INIT('h80)
	) name12924 (
		_w1503_,
		_w1549_,
		_w13301_,
		_w14274_
	);
	LUT4 #(
		.INIT('h000d)
	) name12925 (
		\P2_EBX_reg[19]/NET0131 ,
		_w8961_,
		_w14274_,
		_w14273_,
		_w14275_
	);
	LUT2 #(
		.INIT('h2)
	) name12926 (
		\P2_EBX_reg[19]/NET0131 ,
		_w7767_,
		_w14276_
	);
	LUT3 #(
		.INIT('hf2)
	) name12927 (
		_w1678_,
		_w14275_,
		_w14276_,
		_w14277_
	);
	LUT3 #(
		.INIT('h80)
	) name12928 (
		_w1503_,
		_w1549_,
		_w10398_,
		_w14278_
	);
	LUT2 #(
		.INIT('h8)
	) name12929 (
		_w1578_,
		_w11358_,
		_w14279_
	);
	LUT4 #(
		.INIT('h000d)
	) name12930 (
		\P2_EBX_reg[1]/NET0131 ,
		_w8961_,
		_w14278_,
		_w14279_,
		_w14280_
	);
	LUT2 #(
		.INIT('h2)
	) name12931 (
		\P2_EBX_reg[1]/NET0131 ,
		_w7767_,
		_w14281_
	);
	LUT3 #(
		.INIT('hf2)
	) name12932 (
		_w1678_,
		_w14280_,
		_w14281_,
		_w14282_
	);
	LUT4 #(
		.INIT('h8000)
	) name12933 (
		\P2_EBX_reg[19]/NET0131 ,
		\P2_EBX_reg[20]/NET0131 ,
		_w8953_,
		_w8954_,
		_w14283_
	);
	LUT3 #(
		.INIT('h48)
	) name12934 (
		\P2_EBX_reg[20]/NET0131 ,
		_w1578_,
		_w8955_,
		_w14284_
	);
	LUT3 #(
		.INIT('h80)
	) name12935 (
		_w1503_,
		_w1549_,
		_w13322_,
		_w14285_
	);
	LUT3 #(
		.INIT('h0d)
	) name12936 (
		\P2_EBX_reg[20]/NET0131 ,
		_w8961_,
		_w14285_,
		_w14286_
	);
	LUT2 #(
		.INIT('h2)
	) name12937 (
		\P2_EBX_reg[20]/NET0131 ,
		_w7767_,
		_w14287_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12938 (
		_w1678_,
		_w14284_,
		_w14286_,
		_w14287_,
		_w14288_
	);
	LUT3 #(
		.INIT('h48)
	) name12939 (
		\P2_EBX_reg[21]/NET0131 ,
		_w1578_,
		_w14283_,
		_w14289_
	);
	LUT3 #(
		.INIT('h80)
	) name12940 (
		_w1503_,
		_w1549_,
		_w13344_,
		_w14290_
	);
	LUT3 #(
		.INIT('h0d)
	) name12941 (
		\P2_EBX_reg[21]/NET0131 ,
		_w8961_,
		_w14290_,
		_w14291_
	);
	LUT2 #(
		.INIT('h2)
	) name12942 (
		\P2_EBX_reg[21]/NET0131 ,
		_w7767_,
		_w14292_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12943 (
		_w1678_,
		_w14289_,
		_w14291_,
		_w14292_,
		_w14293_
	);
	LUT4 #(
		.INIT('h60c0)
	) name12944 (
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		_w1578_,
		_w14283_,
		_w14294_
	);
	LUT3 #(
		.INIT('h80)
	) name12945 (
		_w1503_,
		_w1549_,
		_w13363_,
		_w14295_
	);
	LUT3 #(
		.INIT('h0d)
	) name12946 (
		\P2_EBX_reg[22]/NET0131 ,
		_w8961_,
		_w14295_,
		_w14296_
	);
	LUT2 #(
		.INIT('h2)
	) name12947 (
		\P2_EBX_reg[22]/NET0131 ,
		_w7767_,
		_w14297_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12948 (
		_w1678_,
		_w14294_,
		_w14296_,
		_w14297_,
		_w14298_
	);
	LUT4 #(
		.INIT('h070f)
	) name12949 (
		\P2_EBX_reg[21]/NET0131 ,
		\P2_EBX_reg[22]/NET0131 ,
		\P2_EBX_reg[23]/NET0131 ,
		_w14283_,
		_w14299_
	);
	LUT2 #(
		.INIT('h2)
	) name12950 (
		_w1578_,
		_w8957_,
		_w14300_
	);
	LUT3 #(
		.INIT('h80)
	) name12951 (
		_w1503_,
		_w1549_,
		_w13375_,
		_w14301_
	);
	LUT3 #(
		.INIT('h0d)
	) name12952 (
		\P2_EBX_reg[23]/NET0131 ,
		_w8961_,
		_w14301_,
		_w14302_
	);
	LUT4 #(
		.INIT('h20aa)
	) name12953 (
		_w1678_,
		_w14299_,
		_w14300_,
		_w14302_,
		_w14303_
	);
	LUT2 #(
		.INIT('h2)
	) name12954 (
		\P2_EBX_reg[23]/NET0131 ,
		_w7767_,
		_w14304_
	);
	LUT2 #(
		.INIT('he)
	) name12955 (
		_w14303_,
		_w14304_,
		_w14305_
	);
	LUT3 #(
		.INIT('h48)
	) name12956 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1578_,
		_w8957_,
		_w14306_
	);
	LUT4 #(
		.INIT('h002a)
	) name12957 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1503_,
		_w1549_,
		_w1578_,
		_w14307_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name12958 (
		\P2_EBX_reg[24]/NET0131 ,
		_w1596_,
		_w7815_,
		_w7826_,
		_w14308_
	);
	LUT3 #(
		.INIT('h08)
	) name12959 (
		_w1503_,
		_w1549_,
		_w14308_,
		_w14309_
	);
	LUT2 #(
		.INIT('h1)
	) name12960 (
		_w14307_,
		_w14309_,
		_w14310_
	);
	LUT2 #(
		.INIT('h2)
	) name12961 (
		\P2_EBX_reg[24]/NET0131 ,
		_w7767_,
		_w14311_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12962 (
		_w1678_,
		_w14306_,
		_w14310_,
		_w14311_,
		_w14312_
	);
	LUT3 #(
		.INIT('ha8)
	) name12963 (
		\P1_EBX_reg[2]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14313_
	);
	LUT3 #(
		.INIT('h80)
	) name12964 (
		_w1750_,
		_w1813_,
		_w10017_,
		_w14314_
	);
	LUT3 #(
		.INIT('h78)
	) name12965 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		_w14315_
	);
	LUT3 #(
		.INIT('h80)
	) name12966 (
		_w1826_,
		_w1828_,
		_w14315_,
		_w14316_
	);
	LUT2 #(
		.INIT('h1)
	) name12967 (
		_w14314_,
		_w14316_,
		_w14317_
	);
	LUT2 #(
		.INIT('h2)
	) name12968 (
		\P1_EBX_reg[2]/NET0131 ,
		_w9102_,
		_w14318_
	);
	LUT4 #(
		.INIT('hff8a)
	) name12969 (
		_w1933_,
		_w14313_,
		_w14317_,
		_w14318_,
		_w14319_
	);
	LUT4 #(
		.INIT('h31f5)
	) name12970 (
		\P2_EBX_reg[28]/NET0131 ,
		_w1550_,
		_w8961_,
		_w13392_,
		_w14320_
	);
	LUT4 #(
		.INIT('hb700)
	) name12971 (
		\P2_EBX_reg[28]/NET0131 ,
		_w1578_,
		_w8960_,
		_w14320_,
		_w14321_
	);
	LUT2 #(
		.INIT('h2)
	) name12972 (
		\P2_EBX_reg[28]/NET0131 ,
		_w7767_,
		_w14322_
	);
	LUT3 #(
		.INIT('hf2)
	) name12973 (
		_w1678_,
		_w14321_,
		_w14322_,
		_w14323_
	);
	LUT3 #(
		.INIT('h80)
	) name12974 (
		_w1503_,
		_w1549_,
		_w10406_,
		_w14324_
	);
	LUT3 #(
		.INIT('h78)
	) name12975 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		_w14325_
	);
	LUT2 #(
		.INIT('h8)
	) name12976 (
		_w1578_,
		_w14325_,
		_w14326_
	);
	LUT4 #(
		.INIT('h000d)
	) name12977 (
		\P2_EBX_reg[2]/NET0131 ,
		_w8961_,
		_w14324_,
		_w14326_,
		_w14327_
	);
	LUT2 #(
		.INIT('h2)
	) name12978 (
		\P2_EBX_reg[2]/NET0131 ,
		_w7767_,
		_w14328_
	);
	LUT3 #(
		.INIT('hf2)
	) name12979 (
		_w1678_,
		_w14327_,
		_w14328_,
		_w14329_
	);
	LUT3 #(
		.INIT('h80)
	) name12980 (
		_w1503_,
		_w1549_,
		_w10414_,
		_w14330_
	);
	LUT4 #(
		.INIT('h7f80)
	) name12981 (
		\P2_EBX_reg[0]/NET0131 ,
		\P2_EBX_reg[1]/NET0131 ,
		\P2_EBX_reg[2]/NET0131 ,
		\P2_EBX_reg[3]/NET0131 ,
		_w14331_
	);
	LUT2 #(
		.INIT('h8)
	) name12982 (
		_w1578_,
		_w14331_,
		_w14332_
	);
	LUT4 #(
		.INIT('h000d)
	) name12983 (
		\P2_EBX_reg[3]/NET0131 ,
		_w8961_,
		_w14330_,
		_w14332_,
		_w14333_
	);
	LUT2 #(
		.INIT('h2)
	) name12984 (
		\P2_EBX_reg[3]/NET0131 ,
		_w7767_,
		_w14334_
	);
	LUT3 #(
		.INIT('hf2)
	) name12985 (
		_w1678_,
		_w14333_,
		_w14334_,
		_w14335_
	);
	LUT3 #(
		.INIT('h80)
	) name12986 (
		_w1503_,
		_w1549_,
		_w10422_,
		_w14336_
	);
	LUT2 #(
		.INIT('h6)
	) name12987 (
		\P2_EBX_reg[4]/NET0131 ,
		_w8944_,
		_w14337_
	);
	LUT2 #(
		.INIT('h8)
	) name12988 (
		_w1578_,
		_w14337_,
		_w14338_
	);
	LUT4 #(
		.INIT('h000d)
	) name12989 (
		\P2_EBX_reg[4]/NET0131 ,
		_w8961_,
		_w14336_,
		_w14338_,
		_w14339_
	);
	LUT2 #(
		.INIT('h2)
	) name12990 (
		\P2_EBX_reg[4]/NET0131 ,
		_w7767_,
		_w14340_
	);
	LUT3 #(
		.INIT('hf2)
	) name12991 (
		_w1678_,
		_w14339_,
		_w14340_,
		_w14341_
	);
	LUT3 #(
		.INIT('h80)
	) name12992 (
		_w1503_,
		_w1549_,
		_w10448_,
		_w14342_
	);
	LUT3 #(
		.INIT('h6c)
	) name12993 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		_w8944_,
		_w14343_
	);
	LUT2 #(
		.INIT('h8)
	) name12994 (
		_w1578_,
		_w14343_,
		_w14344_
	);
	LUT4 #(
		.INIT('h000d)
	) name12995 (
		\P2_EBX_reg[5]/NET0131 ,
		_w8961_,
		_w14342_,
		_w14344_,
		_w14345_
	);
	LUT2 #(
		.INIT('h2)
	) name12996 (
		\P2_EBX_reg[5]/NET0131 ,
		_w7767_,
		_w14346_
	);
	LUT3 #(
		.INIT('hf2)
	) name12997 (
		_w1678_,
		_w14345_,
		_w14346_,
		_w14347_
	);
	LUT3 #(
		.INIT('ha8)
	) name12998 (
		\P1_EBX_reg[3]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14348_
	);
	LUT3 #(
		.INIT('h80)
	) name12999 (
		_w1750_,
		_w1813_,
		_w10045_,
		_w14349_
	);
	LUT4 #(
		.INIT('h7f80)
	) name13000 (
		\P1_EBX_reg[0]/NET0131 ,
		\P1_EBX_reg[1]/NET0131 ,
		\P1_EBX_reg[2]/NET0131 ,
		\P1_EBX_reg[3]/NET0131 ,
		_w14350_
	);
	LUT3 #(
		.INIT('h80)
	) name13001 (
		_w1826_,
		_w1828_,
		_w14350_,
		_w14351_
	);
	LUT2 #(
		.INIT('h1)
	) name13002 (
		_w14349_,
		_w14351_,
		_w14352_
	);
	LUT2 #(
		.INIT('h2)
	) name13003 (
		\P1_EBX_reg[3]/NET0131 ,
		_w9102_,
		_w14353_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13004 (
		_w1933_,
		_w14348_,
		_w14352_,
		_w14353_,
		_w14354_
	);
	LUT3 #(
		.INIT('h80)
	) name13005 (
		_w1503_,
		_w1549_,
		_w10456_,
		_w14355_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13006 (
		\P2_EBX_reg[4]/NET0131 ,
		\P2_EBX_reg[5]/NET0131 ,
		\P2_EBX_reg[6]/NET0131 ,
		_w8944_,
		_w14356_
	);
	LUT2 #(
		.INIT('h8)
	) name13007 (
		_w1578_,
		_w14356_,
		_w14357_
	);
	LUT4 #(
		.INIT('h000d)
	) name13008 (
		\P2_EBX_reg[6]/NET0131 ,
		_w8961_,
		_w14355_,
		_w14357_,
		_w14358_
	);
	LUT2 #(
		.INIT('h2)
	) name13009 (
		\P2_EBX_reg[6]/NET0131 ,
		_w7767_,
		_w14359_
	);
	LUT3 #(
		.INIT('hf2)
	) name13010 (
		_w1678_,
		_w14358_,
		_w14359_,
		_w14360_
	);
	LUT2 #(
		.INIT('h2)
	) name13011 (
		_w1596_,
		_w4214_,
		_w14361_
	);
	LUT3 #(
		.INIT('h80)
	) name13012 (
		_w1503_,
		_w1549_,
		_w14361_,
		_w14362_
	);
	LUT2 #(
		.INIT('h6)
	) name13013 (
		\P2_EBX_reg[7]/NET0131 ,
		_w8945_,
		_w14363_
	);
	LUT2 #(
		.INIT('h8)
	) name13014 (
		_w1578_,
		_w14363_,
		_w14364_
	);
	LUT4 #(
		.INIT('h000d)
	) name13015 (
		\P2_EBX_reg[7]/NET0131 ,
		_w8961_,
		_w14362_,
		_w14364_,
		_w14365_
	);
	LUT2 #(
		.INIT('h2)
	) name13016 (
		\P2_EBX_reg[7]/NET0131 ,
		_w7767_,
		_w14366_
	);
	LUT3 #(
		.INIT('hf2)
	) name13017 (
		_w1678_,
		_w14365_,
		_w14366_,
		_w14367_
	);
	LUT3 #(
		.INIT('h80)
	) name13018 (
		_w1503_,
		_w1549_,
		_w10474_,
		_w14368_
	);
	LUT3 #(
		.INIT('h6c)
	) name13019 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		_w8945_,
		_w14369_
	);
	LUT2 #(
		.INIT('h8)
	) name13020 (
		_w1578_,
		_w14369_,
		_w14370_
	);
	LUT4 #(
		.INIT('h000d)
	) name13021 (
		\P2_EBX_reg[8]/NET0131 ,
		_w8961_,
		_w14368_,
		_w14370_,
		_w14371_
	);
	LUT2 #(
		.INIT('h2)
	) name13022 (
		\P2_EBX_reg[8]/NET0131 ,
		_w7767_,
		_w14372_
	);
	LUT3 #(
		.INIT('hf2)
	) name13023 (
		_w1678_,
		_w14371_,
		_w14372_,
		_w14373_
	);
	LUT3 #(
		.INIT('h80)
	) name13024 (
		_w1503_,
		_w1549_,
		_w10497_,
		_w14374_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13025 (
		\P2_EBX_reg[7]/NET0131 ,
		\P2_EBX_reg[8]/NET0131 ,
		\P2_EBX_reg[9]/NET0131 ,
		_w8945_,
		_w14375_
	);
	LUT2 #(
		.INIT('h8)
	) name13026 (
		_w1578_,
		_w14375_,
		_w14376_
	);
	LUT4 #(
		.INIT('h000d)
	) name13027 (
		\P2_EBX_reg[9]/NET0131 ,
		_w8961_,
		_w14374_,
		_w14376_,
		_w14377_
	);
	LUT2 #(
		.INIT('h2)
	) name13028 (
		\P2_EBX_reg[9]/NET0131 ,
		_w7767_,
		_w14378_
	);
	LUT3 #(
		.INIT('hf2)
	) name13029 (
		_w1678_,
		_w14377_,
		_w14378_,
		_w14379_
	);
	LUT3 #(
		.INIT('ha8)
	) name13030 (
		\P1_EBX_reg[4]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14380_
	);
	LUT3 #(
		.INIT('h80)
	) name13031 (
		_w1750_,
		_w1813_,
		_w10141_,
		_w14381_
	);
	LUT2 #(
		.INIT('h6)
	) name13032 (
		\P1_EBX_reg[4]/NET0131 ,
		_w8973_,
		_w14382_
	);
	LUT3 #(
		.INIT('h80)
	) name13033 (
		_w1826_,
		_w1828_,
		_w14382_,
		_w14383_
	);
	LUT2 #(
		.INIT('h1)
	) name13034 (
		_w14381_,
		_w14383_,
		_w14384_
	);
	LUT2 #(
		.INIT('h2)
	) name13035 (
		\P1_EBX_reg[4]/NET0131 ,
		_w9102_,
		_w14385_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13036 (
		_w1933_,
		_w14380_,
		_w14384_,
		_w14385_,
		_w14386_
	);
	LUT3 #(
		.INIT('ha8)
	) name13037 (
		\P1_EBX_reg[5]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14387_
	);
	LUT3 #(
		.INIT('h80)
	) name13038 (
		_w1750_,
		_w1813_,
		_w10159_,
		_w14388_
	);
	LUT3 #(
		.INIT('h6c)
	) name13039 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		_w8973_,
		_w14389_
	);
	LUT3 #(
		.INIT('h80)
	) name13040 (
		_w1826_,
		_w1828_,
		_w14389_,
		_w14390_
	);
	LUT2 #(
		.INIT('h1)
	) name13041 (
		_w14388_,
		_w14390_,
		_w14391_
	);
	LUT2 #(
		.INIT('h2)
	) name13042 (
		\P1_EBX_reg[5]/NET0131 ,
		_w9102_,
		_w14392_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13043 (
		_w1933_,
		_w14387_,
		_w14391_,
		_w14392_,
		_w14393_
	);
	LUT3 #(
		.INIT('ha8)
	) name13044 (
		\P1_EBX_reg[6]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14394_
	);
	LUT3 #(
		.INIT('h80)
	) name13045 (
		_w1750_,
		_w1813_,
		_w10332_,
		_w14395_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13046 (
		\P1_EBX_reg[4]/NET0131 ,
		\P1_EBX_reg[5]/NET0131 ,
		\P1_EBX_reg[6]/NET0131 ,
		_w8973_,
		_w14396_
	);
	LUT3 #(
		.INIT('h80)
	) name13047 (
		_w1826_,
		_w1828_,
		_w14396_,
		_w14397_
	);
	LUT2 #(
		.INIT('h1)
	) name13048 (
		_w14395_,
		_w14397_,
		_w14398_
	);
	LUT2 #(
		.INIT('h2)
	) name13049 (
		\P1_EBX_reg[6]/NET0131 ,
		_w9102_,
		_w14399_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13050 (
		_w1933_,
		_w14394_,
		_w14398_,
		_w14399_,
		_w14400_
	);
	LUT3 #(
		.INIT('ha8)
	) name13051 (
		\P1_EBX_reg[7]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14401_
	);
	LUT3 #(
		.INIT('h80)
	) name13052 (
		_w1750_,
		_w1813_,
		_w10179_,
		_w14402_
	);
	LUT2 #(
		.INIT('h6)
	) name13053 (
		\P1_EBX_reg[7]/NET0131 ,
		_w8974_,
		_w14403_
	);
	LUT3 #(
		.INIT('h80)
	) name13054 (
		_w1826_,
		_w1828_,
		_w14403_,
		_w14404_
	);
	LUT2 #(
		.INIT('h1)
	) name13055 (
		_w14402_,
		_w14404_,
		_w14405_
	);
	LUT2 #(
		.INIT('h2)
	) name13056 (
		\P1_EBX_reg[7]/NET0131 ,
		_w9102_,
		_w14406_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13057 (
		_w1933_,
		_w14401_,
		_w14405_,
		_w14406_,
		_w14407_
	);
	LUT3 #(
		.INIT('ha8)
	) name13058 (
		\P1_EBX_reg[8]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14408_
	);
	LUT3 #(
		.INIT('h80)
	) name13059 (
		_w1750_,
		_w1813_,
		_w10269_,
		_w14409_
	);
	LUT3 #(
		.INIT('h6c)
	) name13060 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		_w8974_,
		_w14410_
	);
	LUT3 #(
		.INIT('h80)
	) name13061 (
		_w1826_,
		_w1828_,
		_w14410_,
		_w14411_
	);
	LUT2 #(
		.INIT('h1)
	) name13062 (
		_w14409_,
		_w14411_,
		_w14412_
	);
	LUT2 #(
		.INIT('h2)
	) name13063 (
		\P1_EBX_reg[8]/NET0131 ,
		_w9102_,
		_w14413_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13064 (
		_w1933_,
		_w14408_,
		_w14412_,
		_w14413_,
		_w14414_
	);
	LUT3 #(
		.INIT('ha8)
	) name13065 (
		\P1_EBX_reg[9]/NET0131 ,
		_w1863_,
		_w8992_,
		_w14415_
	);
	LUT3 #(
		.INIT('h80)
	) name13066 (
		_w1750_,
		_w1813_,
		_w10350_,
		_w14416_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13067 (
		\P1_EBX_reg[7]/NET0131 ,
		\P1_EBX_reg[8]/NET0131 ,
		\P1_EBX_reg[9]/NET0131 ,
		_w8974_,
		_w14417_
	);
	LUT3 #(
		.INIT('h80)
	) name13068 (
		_w1826_,
		_w1828_,
		_w14417_,
		_w14418_
	);
	LUT2 #(
		.INIT('h1)
	) name13069 (
		_w14416_,
		_w14418_,
		_w14419_
	);
	LUT2 #(
		.INIT('h2)
	) name13070 (
		\P1_EBX_reg[9]/NET0131 ,
		_w9102_,
		_w14420_
	);
	LUT4 #(
		.INIT('hff8a)
	) name13071 (
		_w1933_,
		_w14415_,
		_w14419_,
		_w14420_,
		_w14421_
	);
	LUT2 #(
		.INIT('h2)
	) name13072 (
		\P3_uWord_reg[3]/NET0131 ,
		_w8341_,
		_w14422_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13073 (
		\P3_uWord_reg[3]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14423_
	);
	LUT3 #(
		.INIT('h04)
	) name13074 (
		_w2060_,
		_w2047_,
		_w14423_,
		_w14424_
	);
	LUT3 #(
		.INIT('ha2)
	) name13075 (
		\P3_uWord_reg[3]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14425_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13076 (
		_w1945_,
		_w13905_,
		_w14424_,
		_w14425_,
		_w14426_
	);
	LUT2 #(
		.INIT('he)
	) name13077 (
		_w14422_,
		_w14426_,
		_w14427_
	);
	LUT3 #(
		.INIT('ha2)
	) name13078 (
		\P3_uWord_reg[7]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14428_
	);
	LUT3 #(
		.INIT('h40)
	) name13079 (
		_w2060_,
		_w2047_,
		_w13186_,
		_w14429_
	);
	LUT4 #(
		.INIT('haa20)
	) name13080 (
		_w1945_,
		_w13909_,
		_w13910_,
		_w14429_,
		_w14430_
	);
	LUT2 #(
		.INIT('he)
	) name13081 (
		_w14428_,
		_w14430_,
		_w14431_
	);
	LUT4 #(
		.INIT('haa02)
	) name13082 (
		_w1945_,
		_w2044_,
		_w2047_,
		_w2105_,
		_w14432_
	);
	LUT4 #(
		.INIT('heece)
	) name13083 (
		\P3_CodeFetch_reg/NET0131 ,
		_w2195_,
		_w8341_,
		_w14432_,
		_w14433_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13084 (
		\P2_CodeFetch_reg/NET0131 ,
		_w1678_,
		_w7767_,
		_w9788_,
		_w14434_
	);
	LUT2 #(
		.INIT('he)
	) name13085 (
		_w1682_,
		_w14434_,
		_w14435_
	);
	LUT2 #(
		.INIT('h2)
	) name13086 (
		\datao[30]_pad ,
		_w2115_,
		_w14436_
	);
	LUT4 #(
		.INIT('h8000)
	) name13087 (
		\P3_EAX_reg[28]/NET0131 ,
		\P3_EAX_reg[29]/NET0131 ,
		_w8362_,
		_w9541_,
		_w14437_
	);
	LUT3 #(
		.INIT('h48)
	) name13088 (
		\P3_EAX_reg[30]/NET0131 ,
		_w9543_,
		_w14437_,
		_w14438_
	);
	LUT4 #(
		.INIT('h1020)
	) name13089 (
		\P3_EAX_reg[30]/NET0131 ,
		_w2111_,
		_w9543_,
		_w14437_,
		_w14439_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13090 (
		\P3_uWord_reg[14]/NET0131 ,
		\datao[30]_pad ,
		_w9977_,
		_w9978_,
		_w14440_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13091 (
		_w1945_,
		_w14436_,
		_w14439_,
		_w14440_,
		_w14441_
	);
	LUT3 #(
		.INIT('h8a)
	) name13092 (
		\P2_Datao_reg[30]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14442_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13093 (
		\P2_EAX_reg[28]/NET0131 ,
		\P2_EAX_reg[29]/NET0131 ,
		\P2_EAX_reg[30]/NET0131 ,
		_w9461_,
		_w14443_
	);
	LUT2 #(
		.INIT('h8)
	) name13094 (
		_w1675_,
		_w14443_,
		_w14444_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13095 (
		\P2_Datao_reg[30]/NET0131 ,
		\P2_uWord_reg[14]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14445_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13096 (
		_w1678_,
		_w14442_,
		_w14444_,
		_w14445_,
		_w14446_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		_w1858_,
		_w1933_,
		_w14447_
	);
	LUT3 #(
		.INIT('h80)
	) name13098 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w9487_,
		_w14448_
	);
	LUT3 #(
		.INIT('h48)
	) name13099 (
		\P1_EAX_reg[30]/NET0131 ,
		_w9471_,
		_w14448_,
		_w14449_
	);
	LUT4 #(
		.INIT('h4080)
	) name13100 (
		\P1_EAX_reg[30]/NET0131 ,
		_w9471_,
		_w14447_,
		_w14448_,
		_w14450_
	);
	LUT2 #(
		.INIT('h8)
	) name13101 (
		\P1_uWord_reg[14]/NET0131 ,
		_w1935_,
		_w14451_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13102 (
		\P1_Datao_reg[30]/NET0131 ,
		_w1860_,
		_w1933_,
		_w9972_,
		_w14452_
	);
	LUT3 #(
		.INIT('hfe)
	) name13103 (
		_w14451_,
		_w14450_,
		_w14452_,
		_w14453_
	);
	LUT2 #(
		.INIT('h8)
	) name13104 (
		\P1_CodeFetch_reg/NET0131 ,
		_w1933_,
		_w14454_
	);
	LUT3 #(
		.INIT('h31)
	) name13105 (
		\P1_CodeFetch_reg/NET0131 ,
		_w1941_,
		_w9102_,
		_w14455_
	);
	LUT3 #(
		.INIT('h4f)
	) name13106 (
		_w10808_,
		_w14454_,
		_w14455_,
		_w14456_
	);
	LUT2 #(
		.INIT('h2)
	) name13107 (
		\P1_uWord_reg[0]/NET0131 ,
		_w9102_,
		_w14457_
	);
	LUT3 #(
		.INIT('h80)
	) name13108 (
		\P1_uWord_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14458_
	);
	LUT3 #(
		.INIT('h0d)
	) name13109 (
		_w1867_,
		_w3471_,
		_w14458_,
		_w14459_
	);
	LUT2 #(
		.INIT('h2)
	) name13110 (
		_w1795_,
		_w14459_,
		_w14460_
	);
	LUT3 #(
		.INIT('ha6)
	) name13111 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9482_,
		_w14461_
	);
	LUT3 #(
		.INIT('h20)
	) name13112 (
		_w1797_,
		_w1852_,
		_w14461_,
		_w14462_
	);
	LUT4 #(
		.INIT('haa02)
	) name13113 (
		\P1_uWord_reg[0]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14463_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13114 (
		_w1933_,
		_w14462_,
		_w14460_,
		_w14463_,
		_w14464_
	);
	LUT2 #(
		.INIT('he)
	) name13115 (
		_w14457_,
		_w14464_,
		_w14465_
	);
	LUT2 #(
		.INIT('h2)
	) name13116 (
		\P2_uWord_reg[0]/NET0131 ,
		_w7767_,
		_w14466_
	);
	LUT3 #(
		.INIT('h80)
	) name13117 (
		\P2_uWord_reg[0]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w14467_
	);
	LUT3 #(
		.INIT('h0d)
	) name13118 (
		_w1606_,
		_w9115_,
		_w14467_,
		_w14468_
	);
	LUT2 #(
		.INIT('h2)
	) name13119 (
		_w1565_,
		_w14468_,
		_w14469_
	);
	LUT4 #(
		.INIT('haa02)
	) name13120 (
		\P2_uWord_reg[0]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w14470_
	);
	LUT3 #(
		.INIT('ha6)
	) name13121 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9457_,
		_w14471_
	);
	LUT3 #(
		.INIT('h20)
	) name13122 (
		_w1566_,
		_w1602_,
		_w14471_,
		_w14472_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13123 (
		_w1678_,
		_w14469_,
		_w14470_,
		_w14472_,
		_w14473_
	);
	LUT2 #(
		.INIT('he)
	) name13124 (
		_w14466_,
		_w14473_,
		_w14474_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13125 (
		\P2_uWord_reg[10]/NET0131 ,
		_w1678_,
		_w7767_,
		_w9467_,
		_w14475_
	);
	LUT2 #(
		.INIT('h8)
	) name13126 (
		_w1565_,
		_w9522_,
		_w14476_
	);
	LUT3 #(
		.INIT('h48)
	) name13127 (
		\P2_EAX_reg[26]/NET0131 ,
		_w1566_,
		_w9460_,
		_w14477_
	);
	LUT3 #(
		.INIT('ha8)
	) name13128 (
		_w10009_,
		_w14476_,
		_w14477_,
		_w14478_
	);
	LUT2 #(
		.INIT('he)
	) name13129 (
		_w14475_,
		_w14478_,
		_w14479_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13130 (
		\P1_uWord_reg[10]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14480_
	);
	LUT3 #(
		.INIT('h02)
	) name13131 (
		_w1795_,
		_w1861_,
		_w3449_,
		_w14481_
	);
	LUT3 #(
		.INIT('h48)
	) name13132 (
		\P1_EAX_reg[26]/NET0131 ,
		_w1797_,
		_w12846_,
		_w14482_
	);
	LUT3 #(
		.INIT('ha8)
	) name13133 (
		_w9489_,
		_w14481_,
		_w14482_,
		_w14483_
	);
	LUT2 #(
		.INIT('he)
	) name13134 (
		_w14480_,
		_w14483_,
		_w14484_
	);
	LUT2 #(
		.INIT('h2)
	) name13135 (
		\P2_uWord_reg[14]/NET0131 ,
		_w7767_,
		_w14485_
	);
	LUT2 #(
		.INIT('h8)
	) name13136 (
		_w9465_,
		_w14443_,
		_w14486_
	);
	LUT3 #(
		.INIT('h31)
	) name13137 (
		\P2_uWord_reg[14]/NET0131 ,
		_w8939_,
		_w9467_,
		_w14487_
	);
	LUT4 #(
		.INIT('hecee)
	) name13138 (
		_w1678_,
		_w14485_,
		_w14486_,
		_w14487_,
		_w14488_
	);
	LUT2 #(
		.INIT('h2)
	) name13139 (
		\P2_uWord_reg[1]/NET0131 ,
		_w7767_,
		_w14489_
	);
	LUT3 #(
		.INIT('h80)
	) name13140 (
		\P2_uWord_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w14490_
	);
	LUT3 #(
		.INIT('h0d)
	) name13141 (
		_w1606_,
		_w7156_,
		_w14490_,
		_w14491_
	);
	LUT2 #(
		.INIT('h2)
	) name13142 (
		_w1565_,
		_w14491_,
		_w14492_
	);
	LUT4 #(
		.INIT('haa02)
	) name13143 (
		\P2_uWord_reg[1]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w14493_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name13144 (
		\P2_EAX_reg[16]/NET0131 ,
		\P2_EAX_reg[17]/NET0131 ,
		\P2_EAX_reg[31]/NET0131 ,
		_w9457_,
		_w14494_
	);
	LUT3 #(
		.INIT('h20)
	) name13145 (
		_w1566_,
		_w1602_,
		_w14494_,
		_w14495_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13146 (
		_w1678_,
		_w14492_,
		_w14493_,
		_w14495_,
		_w14496_
	);
	LUT2 #(
		.INIT('he)
	) name13147 (
		_w14489_,
		_w14496_,
		_w14497_
	);
	LUT2 #(
		.INIT('h2)
	) name13148 (
		\P2_uWord_reg[2]/NET0131 ,
		_w7767_,
		_w14498_
	);
	LUT3 #(
		.INIT('h80)
	) name13149 (
		\P2_uWord_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w14499_
	);
	LUT3 #(
		.INIT('h0d)
	) name13150 (
		_w1606_,
		_w5487_,
		_w14499_,
		_w14500_
	);
	LUT2 #(
		.INIT('h2)
	) name13151 (
		_w1565_,
		_w14500_,
		_w14501_
	);
	LUT4 #(
		.INIT('haa02)
	) name13152 (
		\P2_uWord_reg[2]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w14502_
	);
	LUT2 #(
		.INIT('h6)
	) name13153 (
		\P2_EAX_reg[18]/NET0131 ,
		_w9458_,
		_w14503_
	);
	LUT3 #(
		.INIT('h20)
	) name13154 (
		_w1566_,
		_w1602_,
		_w14503_,
		_w14504_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13155 (
		_w1678_,
		_w14501_,
		_w14502_,
		_w14504_,
		_w14505_
	);
	LUT2 #(
		.INIT('he)
	) name13156 (
		_w14498_,
		_w14505_,
		_w14506_
	);
	LUT2 #(
		.INIT('h2)
	) name13157 (
		\P1_uWord_reg[13]/NET0131 ,
		_w9102_,
		_w14507_
	);
	LUT3 #(
		.INIT('h6c)
	) name13158 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		_w9487_,
		_w14508_
	);
	LUT2 #(
		.INIT('h8)
	) name13159 (
		_w9471_,
		_w14508_,
		_w14509_
	);
	LUT3 #(
		.INIT('h0d)
	) name13160 (
		\P1_uWord_reg[13]/NET0131 ,
		_w9473_,
		_w9660_,
		_w14510_
	);
	LUT4 #(
		.INIT('hecee)
	) name13161 (
		_w1933_,
		_w14507_,
		_w14509_,
		_w14510_,
		_w14511_
	);
	LUT2 #(
		.INIT('h2)
	) name13162 (
		\P2_uWord_reg[5]/NET0131 ,
		_w7767_,
		_w14512_
	);
	LUT3 #(
		.INIT('h80)
	) name13163 (
		\P2_uWord_reg[5]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w14513_
	);
	LUT3 #(
		.INIT('h0d)
	) name13164 (
		_w1606_,
		_w6502_,
		_w14513_,
		_w14514_
	);
	LUT2 #(
		.INIT('h2)
	) name13165 (
		_w1565_,
		_w14514_,
		_w14515_
	);
	LUT4 #(
		.INIT('haa02)
	) name13166 (
		\P2_uWord_reg[5]/NET0131 ,
		_w1565_,
		_w1566_,
		_w1602_,
		_w14516_
	);
	LUT4 #(
		.INIT('h0408)
	) name13167 (
		\P2_EAX_reg[21]/NET0131 ,
		_w1566_,
		_w1602_,
		_w9459_,
		_w14517_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13168 (
		_w1678_,
		_w14515_,
		_w14516_,
		_w14517_,
		_w14518_
	);
	LUT2 #(
		.INIT('he)
	) name13169 (
		_w14512_,
		_w14518_,
		_w14519_
	);
	LUT2 #(
		.INIT('h2)
	) name13170 (
		\P1_uWord_reg[14]/NET0131 ,
		_w9102_,
		_w14520_
	);
	LUT3 #(
		.INIT('h08)
	) name13171 (
		_w1795_,
		_w1867_,
		_w3457_,
		_w14521_
	);
	LUT3 #(
		.INIT('h0d)
	) name13172 (
		\P1_uWord_reg[14]/NET0131 ,
		_w9473_,
		_w14521_,
		_w14522_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name13173 (
		_w1933_,
		_w14449_,
		_w14520_,
		_w14522_,
		_w14523_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13174 (
		\P2_uWord_reg[6]/NET0131 ,
		_w1678_,
		_w7767_,
		_w9467_,
		_w14524_
	);
	LUT3 #(
		.INIT('h6c)
	) name13175 (
		\P2_EAX_reg[21]/NET0131 ,
		\P2_EAX_reg[22]/NET0131 ,
		_w9459_,
		_w14525_
	);
	LUT4 #(
		.INIT('h135f)
	) name13176 (
		_w1565_,
		_w1566_,
		_w12977_,
		_w14525_,
		_w14526_
	);
	LUT2 #(
		.INIT('h2)
	) name13177 (
		_w10009_,
		_w14526_,
		_w14527_
	);
	LUT2 #(
		.INIT('he)
	) name13178 (
		_w14524_,
		_w14527_,
		_w14528_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13179 (
		\P1_uWord_reg[1]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14529_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name13180 (
		\P1_EAX_reg[16]/NET0131 ,
		\P1_EAX_reg[17]/NET0131 ,
		\P1_EAX_reg[31]/NET0131 ,
		_w9482_,
		_w14530_
	);
	LUT3 #(
		.INIT('h20)
	) name13181 (
		_w1797_,
		_w1852_,
		_w14530_,
		_w14531_
	);
	LUT3 #(
		.INIT('h08)
	) name13182 (
		_w1795_,
		_w1867_,
		_w3478_,
		_w14532_
	);
	LUT3 #(
		.INIT('ha8)
	) name13183 (
		_w1933_,
		_w14531_,
		_w14532_,
		_w14533_
	);
	LUT2 #(
		.INIT('he)
	) name13184 (
		_w14529_,
		_w14533_,
		_w14534_
	);
	LUT2 #(
		.INIT('h2)
	) name13185 (
		\P1_uWord_reg[2]/NET0131 ,
		_w9102_,
		_w14535_
	);
	LUT3 #(
		.INIT('h80)
	) name13186 (
		\P1_uWord_reg[2]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14536_
	);
	LUT3 #(
		.INIT('h0d)
	) name13187 (
		_w1867_,
		_w3481_,
		_w14536_,
		_w14537_
	);
	LUT2 #(
		.INIT('h2)
	) name13188 (
		_w1795_,
		_w14537_,
		_w14538_
	);
	LUT4 #(
		.INIT('haa02)
	) name13189 (
		\P1_uWord_reg[2]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14539_
	);
	LUT2 #(
		.INIT('h6)
	) name13190 (
		\P1_EAX_reg[18]/NET0131 ,
		_w9483_,
		_w14540_
	);
	LUT3 #(
		.INIT('h20)
	) name13191 (
		_w1797_,
		_w1852_,
		_w14540_,
		_w14541_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13192 (
		_w1933_,
		_w14539_,
		_w14538_,
		_w14541_,
		_w14542_
	);
	LUT2 #(
		.INIT('he)
	) name13193 (
		_w14535_,
		_w14542_,
		_w14543_
	);
	LUT2 #(
		.INIT('h2)
	) name13194 (
		\P2_uWord_reg[9]/NET0131 ,
		_w7767_,
		_w14544_
	);
	LUT2 #(
		.INIT('h1)
	) name13195 (
		\P2_EAX_reg[25]/NET0131 ,
		_w9990_,
		_w14545_
	);
	LUT3 #(
		.INIT('h02)
	) name13196 (
		_w1566_,
		_w1602_,
		_w9460_,
		_w14546_
	);
	LUT2 #(
		.INIT('h4)
	) name13197 (
		_w14545_,
		_w14546_,
		_w14547_
	);
	LUT2 #(
		.INIT('h8)
	) name13198 (
		_w1565_,
		_w10485_,
		_w14548_
	);
	LUT3 #(
		.INIT('h0d)
	) name13199 (
		\P2_uWord_reg[9]/NET0131 ,
		_w9467_,
		_w14548_,
		_w14549_
	);
	LUT4 #(
		.INIT('hecee)
	) name13200 (
		_w1678_,
		_w14544_,
		_w14547_,
		_w14549_,
		_w14550_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13201 (
		\P1_uWord_reg[5]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14551_
	);
	LUT2 #(
		.INIT('h1)
	) name13202 (
		\P1_EAX_reg[21]/NET0131 ,
		_w12492_,
		_w14552_
	);
	LUT4 #(
		.INIT('h0002)
	) name13203 (
		_w1797_,
		_w1852_,
		_w9484_,
		_w14552_,
		_w14553_
	);
	LUT3 #(
		.INIT('h08)
	) name13204 (
		_w1795_,
		_w1867_,
		_w3452_,
		_w14554_
	);
	LUT3 #(
		.INIT('ha8)
	) name13205 (
		_w1933_,
		_w14553_,
		_w14554_,
		_w14555_
	);
	LUT2 #(
		.INIT('he)
	) name13206 (
		_w14551_,
		_w14555_,
		_w14556_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13207 (
		\P1_uWord_reg[6]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14557_
	);
	LUT3 #(
		.INIT('h08)
	) name13208 (
		_w1795_,
		_w1867_,
		_w3474_,
		_w14558_
	);
	LUT4 #(
		.INIT('h0408)
	) name13209 (
		\P1_EAX_reg[22]/NET0131 ,
		_w1797_,
		_w1852_,
		_w9484_,
		_w14559_
	);
	LUT3 #(
		.INIT('ha8)
	) name13210 (
		_w1933_,
		_w14558_,
		_w14559_,
		_w14560_
	);
	LUT2 #(
		.INIT('he)
	) name13211 (
		_w14557_,
		_w14560_,
		_w14561_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13212 (
		\P1_uWord_reg[9]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14562_
	);
	LUT3 #(
		.INIT('h48)
	) name13213 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1797_,
		_w9486_,
		_w14563_
	);
	LUT3 #(
		.INIT('h02)
	) name13214 (
		_w1795_,
		_w1861_,
		_w3445_,
		_w14564_
	);
	LUT3 #(
		.INIT('ha8)
	) name13215 (
		_w9489_,
		_w14563_,
		_w14564_,
		_w14565_
	);
	LUT2 #(
		.INIT('he)
	) name13216 (
		_w14562_,
		_w14565_,
		_w14566_
	);
	LUT2 #(
		.INIT('h2)
	) name13217 (
		\P3_uWord_reg[0]/NET0131 ,
		_w8341_,
		_w14567_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13218 (
		\P3_uWord_reg[0]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14568_
	);
	LUT3 #(
		.INIT('h04)
	) name13219 (
		_w2060_,
		_w2047_,
		_w14568_,
		_w14569_
	);
	LUT3 #(
		.INIT('ha2)
	) name13220 (
		\P3_uWord_reg[0]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14570_
	);
	LUT3 #(
		.INIT('ha6)
	) name13221 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w9537_,
		_w14571_
	);
	LUT4 #(
		.INIT('h0800)
	) name13222 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w14571_,
		_w14572_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13223 (
		_w1945_,
		_w14569_,
		_w14570_,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('he)
	) name13224 (
		_w14567_,
		_w14573_,
		_w14574_
	);
	LUT3 #(
		.INIT('ha2)
	) name13225 (
		\P3_uWord_reg[10]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14575_
	);
	LUT4 #(
		.INIT('h0020)
	) name13226 (
		\buf2_reg[10]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2116_,
		_w14576_
	);
	LUT4 #(
		.INIT('h4080)
	) name13227 (
		\P3_EAX_reg[26]/NET0131 ,
		_w2060_,
		_w2047_,
		_w9541_,
		_w14577_
	);
	LUT3 #(
		.INIT('ha8)
	) name13228 (
		_w10595_,
		_w14576_,
		_w14577_,
		_w14578_
	);
	LUT2 #(
		.INIT('he)
	) name13229 (
		_w14575_,
		_w14578_,
		_w14579_
	);
	LUT2 #(
		.INIT('h2)
	) name13230 (
		\P3_uWord_reg[13]/NET0131 ,
		_w8341_,
		_w14580_
	);
	LUT3 #(
		.INIT('h48)
	) name13231 (
		\P3_EAX_reg[29]/NET0131 ,
		_w9543_,
		_w9544_,
		_w14581_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13232 (
		\P3_uWord_reg[13]/NET0131 ,
		_w2047_,
		_w2105_,
		_w9528_,
		_w14582_
	);
	LUT3 #(
		.INIT('h02)
	) name13233 (
		\buf2_reg[13]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14583_
	);
	LUT3 #(
		.INIT('h40)
	) name13234 (
		_w2060_,
		_w2047_,
		_w14583_,
		_w14584_
	);
	LUT2 #(
		.INIT('h1)
	) name13235 (
		_w14582_,
		_w14584_,
		_w14585_
	);
	LUT4 #(
		.INIT('hecee)
	) name13236 (
		_w1945_,
		_w14580_,
		_w14581_,
		_w14585_,
		_w14586_
	);
	LUT2 #(
		.INIT('h2)
	) name13237 (
		\P3_uWord_reg[14]/NET0131 ,
		_w8341_,
		_w14587_
	);
	LUT4 #(
		.INIT('haaa2)
	) name13238 (
		\P3_uWord_reg[14]/NET0131 ,
		_w2047_,
		_w2105_,
		_w9528_,
		_w14588_
	);
	LUT4 #(
		.INIT('h2000)
	) name13239 (
		\buf2_reg[14]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2119_,
		_w14589_
	);
	LUT2 #(
		.INIT('h1)
	) name13240 (
		_w14588_,
		_w14589_,
		_w14590_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name13241 (
		_w1945_,
		_w14438_,
		_w14587_,
		_w14590_,
		_w14591_
	);
	LUT2 #(
		.INIT('h2)
	) name13242 (
		\P3_uWord_reg[1]/NET0131 ,
		_w8341_,
		_w14592_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13243 (
		\P3_uWord_reg[1]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14593_
	);
	LUT3 #(
		.INIT('h04)
	) name13244 (
		_w2060_,
		_w2047_,
		_w14593_,
		_w14594_
	);
	LUT3 #(
		.INIT('ha2)
	) name13245 (
		\P3_uWord_reg[1]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14595_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name13246 (
		\P3_EAX_reg[16]/NET0131 ,
		\P3_EAX_reg[17]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w9537_,
		_w14596_
	);
	LUT4 #(
		.INIT('h0800)
	) name13247 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w14596_,
		_w14597_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13248 (
		_w1945_,
		_w14594_,
		_w14595_,
		_w14597_,
		_w14598_
	);
	LUT2 #(
		.INIT('he)
	) name13249 (
		_w14592_,
		_w14598_,
		_w14599_
	);
	LUT2 #(
		.INIT('h2)
	) name13250 (
		\P3_uWord_reg[2]/NET0131 ,
		_w8341_,
		_w14600_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13251 (
		\P3_uWord_reg[2]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14601_
	);
	LUT3 #(
		.INIT('h04)
	) name13252 (
		_w2060_,
		_w2047_,
		_w14601_,
		_w14602_
	);
	LUT3 #(
		.INIT('ha2)
	) name13253 (
		\P3_uWord_reg[2]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14603_
	);
	LUT4 #(
		.INIT('haa6a)
	) name13254 (
		\P3_EAX_reg[18]/NET0131 ,
		\P3_EAX_reg[31]/NET0131 ,
		_w8352_,
		_w9537_,
		_w14604_
	);
	LUT4 #(
		.INIT('h0800)
	) name13255 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w14604_,
		_w14605_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13256 (
		_w1945_,
		_w14602_,
		_w14603_,
		_w14605_,
		_w14606_
	);
	LUT2 #(
		.INIT('he)
	) name13257 (
		_w14600_,
		_w14606_,
		_w14607_
	);
	LUT2 #(
		.INIT('h2)
	) name13258 (
		\P3_uWord_reg[5]/NET0131 ,
		_w8341_,
		_w14608_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13259 (
		\P3_uWord_reg[5]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14609_
	);
	LUT3 #(
		.INIT('h04)
	) name13260 (
		_w2060_,
		_w2047_,
		_w14609_,
		_w14610_
	);
	LUT3 #(
		.INIT('ha2)
	) name13261 (
		\P3_uWord_reg[5]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14611_
	);
	LUT4 #(
		.INIT('h78f0)
	) name13262 (
		\P3_EAX_reg[19]/NET0131 ,
		\P3_EAX_reg[20]/NET0131 ,
		\P3_EAX_reg[21]/NET0131 ,
		_w9538_,
		_w14612_
	);
	LUT4 #(
		.INIT('h0800)
	) name13263 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w14612_,
		_w14613_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13264 (
		_w1945_,
		_w14610_,
		_w14611_,
		_w14613_,
		_w14614_
	);
	LUT2 #(
		.INIT('he)
	) name13265 (
		_w14608_,
		_w14614_,
		_w14615_
	);
	LUT2 #(
		.INIT('h2)
	) name13266 (
		\P3_uWord_reg[6]/NET0131 ,
		_w8341_,
		_w14616_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13267 (
		\P3_uWord_reg[6]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14617_
	);
	LUT3 #(
		.INIT('h04)
	) name13268 (
		_w2060_,
		_w2047_,
		_w14617_,
		_w14618_
	);
	LUT3 #(
		.INIT('ha2)
	) name13269 (
		\P3_uWord_reg[6]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14619_
	);
	LUT2 #(
		.INIT('h6)
	) name13270 (
		\P3_EAX_reg[22]/NET0131 ,
		_w9539_,
		_w14620_
	);
	LUT4 #(
		.INIT('h0800)
	) name13271 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w14620_,
		_w14621_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13272 (
		_w1945_,
		_w14618_,
		_w14619_,
		_w14621_,
		_w14622_
	);
	LUT2 #(
		.INIT('he)
	) name13273 (
		_w14616_,
		_w14622_,
		_w14623_
	);
	LUT3 #(
		.INIT('ha2)
	) name13274 (
		\P3_uWord_reg[9]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14624_
	);
	LUT4 #(
		.INIT('h1333)
	) name13275 (
		\P3_EAX_reg[24]/NET0131 ,
		\P3_EAX_reg[25]/NET0131 ,
		_w8357_,
		_w9539_,
		_w14625_
	);
	LUT4 #(
		.INIT('h0008)
	) name13276 (
		_w2060_,
		_w2047_,
		_w2105_,
		_w9541_,
		_w14626_
	);
	LUT3 #(
		.INIT('h02)
	) name13277 (
		\buf2_reg[9]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14627_
	);
	LUT3 #(
		.INIT('h40)
	) name13278 (
		_w2060_,
		_w2047_,
		_w14627_,
		_w14628_
	);
	LUT4 #(
		.INIT('haa20)
	) name13279 (
		_w1945_,
		_w14625_,
		_w14626_,
		_w14628_,
		_w14629_
	);
	LUT2 #(
		.INIT('he)
	) name13280 (
		_w14624_,
		_w14629_,
		_w14630_
	);
	LUT3 #(
		.INIT('h80)
	) name13281 (
		\P1_lWord_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14631_
	);
	LUT3 #(
		.INIT('h0d)
	) name13282 (
		_w1867_,
		_w3471_,
		_w14631_,
		_w14632_
	);
	LUT2 #(
		.INIT('h2)
	) name13283 (
		_w1795_,
		_w14632_,
		_w14633_
	);
	LUT4 #(
		.INIT('haa02)
	) name13284 (
		\P1_lWord_reg[0]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14634_
	);
	LUT3 #(
		.INIT('h08)
	) name13285 (
		\P1_EAX_reg[0]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14635_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13286 (
		_w1933_,
		_w14634_,
		_w14633_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h2)
	) name13287 (
		\P1_lWord_reg[0]/NET0131 ,
		_w9102_,
		_w14637_
	);
	LUT2 #(
		.INIT('he)
	) name13288 (
		_w14636_,
		_w14637_,
		_w14638_
	);
	LUT3 #(
		.INIT('h80)
	) name13289 (
		\P1_lWord_reg[10]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14639_
	);
	LUT3 #(
		.INIT('h0d)
	) name13290 (
		_w1867_,
		_w3449_,
		_w14639_,
		_w14640_
	);
	LUT2 #(
		.INIT('h2)
	) name13291 (
		_w1795_,
		_w14640_,
		_w14641_
	);
	LUT4 #(
		.INIT('haa02)
	) name13292 (
		\P1_lWord_reg[10]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14642_
	);
	LUT3 #(
		.INIT('h08)
	) name13293 (
		\P1_EAX_reg[10]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14643_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13294 (
		_w1933_,
		_w14642_,
		_w14641_,
		_w14643_,
		_w14644_
	);
	LUT2 #(
		.INIT('h2)
	) name13295 (
		\P1_lWord_reg[10]/NET0131 ,
		_w9102_,
		_w14645_
	);
	LUT2 #(
		.INIT('he)
	) name13296 (
		_w14644_,
		_w14645_,
		_w14646_
	);
	LUT3 #(
		.INIT('h80)
	) name13297 (
		\P1_lWord_reg[11]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14647_
	);
	LUT3 #(
		.INIT('h0d)
	) name13298 (
		_w1867_,
		_w3431_,
		_w14647_,
		_w14648_
	);
	LUT2 #(
		.INIT('h2)
	) name13299 (
		_w1795_,
		_w14648_,
		_w14649_
	);
	LUT4 #(
		.INIT('haa02)
	) name13300 (
		\P1_lWord_reg[11]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14650_
	);
	LUT3 #(
		.INIT('h08)
	) name13301 (
		\P1_EAX_reg[11]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14651_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13302 (
		_w1933_,
		_w14650_,
		_w14649_,
		_w14651_,
		_w14652_
	);
	LUT2 #(
		.INIT('h2)
	) name13303 (
		\P1_lWord_reg[11]/NET0131 ,
		_w9102_,
		_w14653_
	);
	LUT2 #(
		.INIT('he)
	) name13304 (
		_w14652_,
		_w14653_,
		_w14654_
	);
	LUT3 #(
		.INIT('h80)
	) name13305 (
		\P1_lWord_reg[12]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w14655_
	);
	LUT3 #(
		.INIT('h0d)
	) name13306 (
		_w1867_,
		_w3464_,
		_w14655_,
		_w14656_
	);
	LUT2 #(
		.INIT('h2)
	) name13307 (
		_w1795_,
		_w14656_,
		_w14657_
	);
	LUT4 #(
		.INIT('haa02)
	) name13308 (
		\P1_lWord_reg[12]/NET0131 ,
		_w1795_,
		_w1797_,
		_w1852_,
		_w14658_
	);
	LUT3 #(
		.INIT('h08)
	) name13309 (
		\P1_EAX_reg[12]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14659_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13310 (
		_w1933_,
		_w14658_,
		_w14657_,
		_w14659_,
		_w14660_
	);
	LUT2 #(
		.INIT('h2)
	) name13311 (
		\P1_lWord_reg[12]/NET0131 ,
		_w9102_,
		_w14661_
	);
	LUT2 #(
		.INIT('he)
	) name13312 (
		_w14660_,
		_w14661_,
		_w14662_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13313 (
		\P1_lWord_reg[13]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14663_
	);
	LUT3 #(
		.INIT('h08)
	) name13314 (
		\P1_EAX_reg[13]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14664_
	);
	LUT3 #(
		.INIT('ha8)
	) name13315 (
		_w1933_,
		_w9660_,
		_w14664_,
		_w14665_
	);
	LUT2 #(
		.INIT('he)
	) name13316 (
		_w14663_,
		_w14665_,
		_w14666_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13317 (
		\P1_lWord_reg[14]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14667_
	);
	LUT3 #(
		.INIT('h08)
	) name13318 (
		\P1_EAX_reg[14]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14668_
	);
	LUT3 #(
		.INIT('ha8)
	) name13319 (
		_w1933_,
		_w14521_,
		_w14668_,
		_w14669_
	);
	LUT2 #(
		.INIT('he)
	) name13320 (
		_w14667_,
		_w14669_,
		_w14670_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13321 (
		\P1_lWord_reg[15]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14671_
	);
	LUT2 #(
		.INIT('h8)
	) name13322 (
		\P1_EAX_reg[15]/NET0131 ,
		_w1797_,
		_w14672_
	);
	LUT3 #(
		.INIT('h02)
	) name13323 (
		_w1795_,
		_w1861_,
		_w3460_,
		_w14673_
	);
	LUT3 #(
		.INIT('ha8)
	) name13324 (
		_w9489_,
		_w14672_,
		_w14673_,
		_w14674_
	);
	LUT2 #(
		.INIT('he)
	) name13325 (
		_w14671_,
		_w14674_,
		_w14675_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13326 (
		\P1_lWord_reg[1]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14676_
	);
	LUT3 #(
		.INIT('h08)
	) name13327 (
		\P1_EAX_reg[1]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14677_
	);
	LUT3 #(
		.INIT('ha8)
	) name13328 (
		_w1933_,
		_w14532_,
		_w14677_,
		_w14678_
	);
	LUT2 #(
		.INIT('he)
	) name13329 (
		_w14676_,
		_w14678_,
		_w14679_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13330 (
		\P1_lWord_reg[3]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14680_
	);
	LUT3 #(
		.INIT('h08)
	) name13331 (
		\P1_EAX_reg[3]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14681_
	);
	LUT3 #(
		.INIT('h08)
	) name13332 (
		_w1795_,
		_w1867_,
		_w3428_,
		_w14682_
	);
	LUT3 #(
		.INIT('ha8)
	) name13333 (
		_w1933_,
		_w14681_,
		_w14682_,
		_w14683_
	);
	LUT2 #(
		.INIT('he)
	) name13334 (
		_w14680_,
		_w14683_,
		_w14684_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13335 (
		\P1_lWord_reg[2]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14685_
	);
	LUT3 #(
		.INIT('h08)
	) name13336 (
		\P1_EAX_reg[2]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14686_
	);
	LUT3 #(
		.INIT('h08)
	) name13337 (
		_w1795_,
		_w1867_,
		_w3481_,
		_w14687_
	);
	LUT3 #(
		.INIT('ha8)
	) name13338 (
		_w1933_,
		_w14686_,
		_w14687_,
		_w14688_
	);
	LUT2 #(
		.INIT('he)
	) name13339 (
		_w14685_,
		_w14688_,
		_w14689_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13340 (
		\P1_lWord_reg[4]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14690_
	);
	LUT3 #(
		.INIT('h08)
	) name13341 (
		\P1_EAX_reg[4]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14691_
	);
	LUT3 #(
		.INIT('ha8)
	) name13342 (
		_w1933_,
		_w12529_,
		_w14691_,
		_w14692_
	);
	LUT2 #(
		.INIT('he)
	) name13343 (
		_w14690_,
		_w14692_,
		_w14693_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13344 (
		\P1_lWord_reg[5]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14694_
	);
	LUT3 #(
		.INIT('h08)
	) name13345 (
		\P1_EAX_reg[5]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14695_
	);
	LUT3 #(
		.INIT('ha8)
	) name13346 (
		_w1933_,
		_w14554_,
		_w14695_,
		_w14696_
	);
	LUT2 #(
		.INIT('he)
	) name13347 (
		_w14694_,
		_w14696_,
		_w14697_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13348 (
		\P1_lWord_reg[6]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14698_
	);
	LUT3 #(
		.INIT('h08)
	) name13349 (
		\P1_EAX_reg[6]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14699_
	);
	LUT3 #(
		.INIT('ha8)
	) name13350 (
		_w1933_,
		_w14558_,
		_w14699_,
		_w14700_
	);
	LUT2 #(
		.INIT('he)
	) name13351 (
		_w14698_,
		_w14700_,
		_w14701_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13352 (
		\P1_lWord_reg[7]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14702_
	);
	LUT3 #(
		.INIT('h08)
	) name13353 (
		\P1_EAX_reg[7]/NET0131 ,
		_w1797_,
		_w1852_,
		_w14703_
	);
	LUT3 #(
		.INIT('ha8)
	) name13354 (
		_w1933_,
		_w12866_,
		_w14703_,
		_w14704_
	);
	LUT2 #(
		.INIT('he)
	) name13355 (
		_w14702_,
		_w14704_,
		_w14705_
	);
	LUT2 #(
		.INIT('h8)
	) name13356 (
		\P1_EAX_reg[8]/NET0131 ,
		_w1797_,
		_w14706_
	);
	LUT3 #(
		.INIT('h54)
	) name13357 (
		_w1852_,
		_w10013_,
		_w14706_,
		_w14707_
	);
	LUT2 #(
		.INIT('h2)
	) name13358 (
		\P1_lWord_reg[8]/NET0131 ,
		_w9473_,
		_w14708_
	);
	LUT2 #(
		.INIT('h2)
	) name13359 (
		\P1_lWord_reg[8]/NET0131 ,
		_w9102_,
		_w14709_
	);
	LUT4 #(
		.INIT('hffa8)
	) name13360 (
		_w1933_,
		_w14707_,
		_w14708_,
		_w14709_,
		_w14710_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13361 (
		\P1_lWord_reg[9]/NET0131 ,
		_w1933_,
		_w9102_,
		_w9473_,
		_w14711_
	);
	LUT2 #(
		.INIT('h8)
	) name13362 (
		\P1_EAX_reg[9]/NET0131 ,
		_w1797_,
		_w14712_
	);
	LUT3 #(
		.INIT('ha8)
	) name13363 (
		_w9489_,
		_w14564_,
		_w14712_,
		_w14713_
	);
	LUT2 #(
		.INIT('he)
	) name13364 (
		_w14711_,
		_w14713_,
		_w14714_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13365 (
		\P3_EAX_reg[12]/NET0131 ,
		\datao[12]_pad ,
		_w1945_,
		_w2115_,
		_w14715_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13366 (
		\P3_lWord_reg[12]/NET0131 ,
		\datao[12]_pad ,
		_w9977_,
		_w9978_,
		_w14716_
	);
	LUT2 #(
		.INIT('hb)
	) name13367 (
		_w14715_,
		_w14716_,
		_w14717_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13368 (
		\P3_EAX_reg[13]/NET0131 ,
		\datao[13]_pad ,
		_w1945_,
		_w2115_,
		_w14718_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13369 (
		\P3_lWord_reg[13]/NET0131 ,
		\datao[13]_pad ,
		_w9977_,
		_w9978_,
		_w14719_
	);
	LUT2 #(
		.INIT('hb)
	) name13370 (
		_w14718_,
		_w14719_,
		_w14720_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13371 (
		\P3_EAX_reg[14]/NET0131 ,
		\datao[14]_pad ,
		_w1945_,
		_w2115_,
		_w14721_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13372 (
		\P3_lWord_reg[14]/NET0131 ,
		\datao[14]_pad ,
		_w9977_,
		_w9978_,
		_w14722_
	);
	LUT2 #(
		.INIT('hb)
	) name13373 (
		_w14721_,
		_w14722_,
		_w14723_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13374 (
		\P3_EAX_reg[2]/NET0131 ,
		\datao[2]_pad ,
		_w1945_,
		_w2115_,
		_w14724_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13375 (
		\P3_lWord_reg[2]/NET0131 ,
		\datao[2]_pad ,
		_w9977_,
		_w9978_,
		_w14725_
	);
	LUT2 #(
		.INIT('hb)
	) name13376 (
		_w14724_,
		_w14725_,
		_w14726_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13377 (
		\P3_EAX_reg[3]/NET0131 ,
		\datao[3]_pad ,
		_w1945_,
		_w2115_,
		_w14727_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13378 (
		\P3_lWord_reg[3]/NET0131 ,
		\datao[3]_pad ,
		_w9977_,
		_w9978_,
		_w14728_
	);
	LUT2 #(
		.INIT('hb)
	) name13379 (
		_w14727_,
		_w14728_,
		_w14729_
	);
	LUT3 #(
		.INIT('h10)
	) name13380 (
		\P2_EAX_reg[0]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14730_
	);
	LUT4 #(
		.INIT('hba00)
	) name13381 (
		\P2_Datao_reg[0]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14731_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13382 (
		\P2_Datao_reg[0]/NET0131 ,
		\P2_lWord_reg[0]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14732_
	);
	LUT3 #(
		.INIT('h4f)
	) name13383 (
		_w14730_,
		_w14731_,
		_w14732_,
		_w14733_
	);
	LUT3 #(
		.INIT('h10)
	) name13384 (
		\P2_EAX_reg[10]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14734_
	);
	LUT4 #(
		.INIT('hba00)
	) name13385 (
		\P2_Datao_reg[10]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14735_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13386 (
		\P2_Datao_reg[10]/NET0131 ,
		\P2_lWord_reg[10]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14736_
	);
	LUT3 #(
		.INIT('h4f)
	) name13387 (
		_w14734_,
		_w14735_,
		_w14736_,
		_w14737_
	);
	LUT3 #(
		.INIT('h10)
	) name13388 (
		\P2_EAX_reg[11]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14738_
	);
	LUT4 #(
		.INIT('hba00)
	) name13389 (
		\P2_Datao_reg[11]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14739_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13390 (
		\P2_Datao_reg[11]/NET0131 ,
		\P2_lWord_reg[11]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14740_
	);
	LUT3 #(
		.INIT('h4f)
	) name13391 (
		_w14738_,
		_w14739_,
		_w14740_,
		_w14741_
	);
	LUT3 #(
		.INIT('h10)
	) name13392 (
		\P2_EAX_reg[12]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14742_
	);
	LUT4 #(
		.INIT('hba00)
	) name13393 (
		\P2_Datao_reg[12]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14743_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13394 (
		\P2_Datao_reg[12]/NET0131 ,
		\P2_lWord_reg[12]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14744_
	);
	LUT3 #(
		.INIT('h4f)
	) name13395 (
		_w14742_,
		_w14743_,
		_w14744_,
		_w14745_
	);
	LUT4 #(
		.INIT('hca00)
	) name13396 (
		\P1_Datao_reg[2]/NET0131 ,
		\P1_EAX_reg[2]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14746_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13397 (
		\P1_Datao_reg[2]/NET0131 ,
		\P1_lWord_reg[2]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14747_
	);
	LUT2 #(
		.INIT('hb)
	) name13398 (
		_w14746_,
		_w14747_,
		_w14748_
	);
	LUT3 #(
		.INIT('h10)
	) name13399 (
		\P2_EAX_reg[5]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14749_
	);
	LUT4 #(
		.INIT('hba00)
	) name13400 (
		\P2_Datao_reg[5]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14750_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13401 (
		\P2_Datao_reg[5]/NET0131 ,
		\P2_lWord_reg[5]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14751_
	);
	LUT3 #(
		.INIT('h4f)
	) name13402 (
		_w14749_,
		_w14750_,
		_w14751_,
		_w14752_
	);
	LUT3 #(
		.INIT('h10)
	) name13403 (
		\P2_EAX_reg[7]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14753_
	);
	LUT4 #(
		.INIT('hba00)
	) name13404 (
		\P2_Datao_reg[7]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14754_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13405 (
		\P2_Datao_reg[7]/NET0131 ,
		\P2_lWord_reg[7]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14755_
	);
	LUT3 #(
		.INIT('h4f)
	) name13406 (
		_w14753_,
		_w14754_,
		_w14755_,
		_w14756_
	);
	LUT3 #(
		.INIT('h10)
	) name13407 (
		\P2_EAX_reg[8]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14757_
	);
	LUT4 #(
		.INIT('hba00)
	) name13408 (
		\P2_Datao_reg[8]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w14758_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13409 (
		\P2_Datao_reg[8]/NET0131 ,
		\P2_lWord_reg[8]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14759_
	);
	LUT3 #(
		.INIT('h4f)
	) name13410 (
		_w14757_,
		_w14758_,
		_w14759_,
		_w14760_
	);
	LUT4 #(
		.INIT('hca00)
	) name13411 (
		\P1_Datao_reg[4]/NET0131 ,
		\P1_EAX_reg[4]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14761_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13412 (
		\P1_Datao_reg[4]/NET0131 ,
		\P1_lWord_reg[4]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14762_
	);
	LUT2 #(
		.INIT('hb)
	) name13413 (
		_w14761_,
		_w14762_,
		_w14763_
	);
	LUT4 #(
		.INIT('hca00)
	) name13414 (
		\P1_Datao_reg[6]/NET0131 ,
		\P1_EAX_reg[6]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14764_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13415 (
		\P1_Datao_reg[6]/NET0131 ,
		\P1_lWord_reg[6]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14765_
	);
	LUT2 #(
		.INIT('hb)
	) name13416 (
		_w14764_,
		_w14765_,
		_w14766_
	);
	LUT4 #(
		.INIT('hca00)
	) name13417 (
		\P1_Datao_reg[8]/NET0131 ,
		\P1_EAX_reg[8]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14767_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13418 (
		\P1_Datao_reg[8]/NET0131 ,
		\P1_lWord_reg[8]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14768_
	);
	LUT2 #(
		.INIT('hb)
	) name13419 (
		_w14767_,
		_w14768_,
		_w14769_
	);
	LUT4 #(
		.INIT('hca00)
	) name13420 (
		\P1_Datao_reg[14]/NET0131 ,
		\P1_EAX_reg[14]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14770_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13421 (
		\P1_Datao_reg[14]/NET0131 ,
		\P1_lWord_reg[14]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14771_
	);
	LUT2 #(
		.INIT('hb)
	) name13422 (
		_w14770_,
		_w14771_,
		_w14772_
	);
	LUT4 #(
		.INIT('hca00)
	) name13423 (
		\P1_Datao_reg[15]/NET0131 ,
		\P1_EAX_reg[15]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14773_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13424 (
		\P1_Datao_reg[15]/NET0131 ,
		\P1_lWord_reg[15]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14774_
	);
	LUT2 #(
		.INIT('hb)
	) name13425 (
		_w14773_,
		_w14774_,
		_w14775_
	);
	LUT4 #(
		.INIT('h080a)
	) name13426 (
		\P1_Datao_reg[18]/NET0131 ,
		_w1725_,
		_w1797_,
		_w1802_,
		_w14776_
	);
	LUT3 #(
		.INIT('he2)
	) name13427 (
		\P1_Datao_reg[18]/NET0131 ,
		_w1859_,
		_w14540_,
		_w14777_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name13428 (
		_w1933_,
		_w12491_,
		_w14776_,
		_w14777_,
		_w14778_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13429 (
		\P1_Datao_reg[18]/NET0131 ,
		\P1_uWord_reg[2]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14779_
	);
	LUT2 #(
		.INIT('hb)
	) name13430 (
		_w14778_,
		_w14779_,
		_w14780_
	);
	LUT4 #(
		.INIT('h0200)
	) name13431 (
		_w1797_,
		_w1852_,
		_w1858_,
		_w14530_,
		_w14781_
	);
	LUT4 #(
		.INIT('hf020)
	) name13432 (
		\P1_Datao_reg[17]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14781_,
		_w14782_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13433 (
		\P1_Datao_reg[17]/NET0131 ,
		\P1_uWord_reg[1]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14783_
	);
	LUT2 #(
		.INIT('hb)
	) name13434 (
		_w14782_,
		_w14783_,
		_w14784_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13435 (
		\P1_Datao_reg[21]/NET0131 ,
		_w1858_,
		_w1860_,
		_w14553_,
		_w14785_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13436 (
		\P1_Datao_reg[21]/NET0131 ,
		\P1_uWord_reg[5]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14786_
	);
	LUT3 #(
		.INIT('h2f)
	) name13437 (
		_w1933_,
		_w14785_,
		_w14786_,
		_w14787_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13438 (
		\P1_Datao_reg[22]/NET0131 ,
		_w1860_,
		_w1933_,
		_w9972_,
		_w14788_
	);
	LUT2 #(
		.INIT('h8)
	) name13439 (
		\P1_uWord_reg[6]/NET0131 ,
		_w1935_,
		_w14789_
	);
	LUT3 #(
		.INIT('h07)
	) name13440 (
		_w14447_,
		_w14559_,
		_w14789_,
		_w14790_
	);
	LUT2 #(
		.INIT('hb)
	) name13441 (
		_w14788_,
		_w14790_,
		_w14791_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13442 (
		\datao[16]_pad ,
		_w2111_,
		_w2115_,
		_w14572_,
		_w14792_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13443 (
		\P3_uWord_reg[0]/NET0131 ,
		\datao[16]_pad ,
		_w9977_,
		_w9978_,
		_w14793_
	);
	LUT3 #(
		.INIT('h2f)
	) name13444 (
		_w1945_,
		_w14792_,
		_w14793_,
		_w14794_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13445 (
		\datao[17]_pad ,
		_w1945_,
		_w2115_,
		_w9978_,
		_w14795_
	);
	LUT2 #(
		.INIT('h8)
	) name13446 (
		\P3_uWord_reg[1]/NET0131 ,
		_w9977_,
		_w14796_
	);
	LUT3 #(
		.INIT('h07)
	) name13447 (
		_w13903_,
		_w14597_,
		_w14796_,
		_w14797_
	);
	LUT2 #(
		.INIT('hb)
	) name13448 (
		_w14795_,
		_w14797_,
		_w14798_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13449 (
		\datao[18]_pad ,
		_w2111_,
		_w2115_,
		_w14605_,
		_w14799_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13450 (
		\P3_uWord_reg[2]/NET0131 ,
		\datao[18]_pad ,
		_w9977_,
		_w9978_,
		_w14800_
	);
	LUT3 #(
		.INIT('h2f)
	) name13451 (
		_w1945_,
		_w14799_,
		_w14800_,
		_w14801_
	);
	LUT4 #(
		.INIT('h4080)
	) name13452 (
		\P1_EAX_reg[25]/NET0131 ,
		_w1797_,
		_w1859_,
		_w9486_,
		_w14802_
	);
	LUT4 #(
		.INIT('hf020)
	) name13453 (
		\P1_Datao_reg[25]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14802_,
		_w14803_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13454 (
		\P1_Datao_reg[25]/NET0131 ,
		\P1_uWord_reg[9]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14804_
	);
	LUT2 #(
		.INIT('hb)
	) name13455 (
		_w14803_,
		_w14804_,
		_w14805_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13456 (
		\datao[21]_pad ,
		_w2111_,
		_w2115_,
		_w14613_,
		_w14806_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13457 (
		\P3_uWord_reg[5]/NET0131 ,
		\datao[21]_pad ,
		_w9977_,
		_w9978_,
		_w14807_
	);
	LUT3 #(
		.INIT('h2f)
	) name13458 (
		_w1945_,
		_w14806_,
		_w14807_,
		_w14808_
	);
	LUT4 #(
		.INIT('h4080)
	) name13459 (
		\P1_EAX_reg[26]/NET0131 ,
		_w1797_,
		_w1859_,
		_w12846_,
		_w14809_
	);
	LUT4 #(
		.INIT('hf020)
	) name13460 (
		\P1_Datao_reg[26]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14809_,
		_w14810_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13461 (
		\P1_Datao_reg[26]/NET0131 ,
		\P1_uWord_reg[10]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14811_
	);
	LUT2 #(
		.INIT('hb)
	) name13462 (
		_w14810_,
		_w14811_,
		_w14812_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name13463 (
		\datao[22]_pad ,
		_w2111_,
		_w2115_,
		_w14621_,
		_w14813_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13464 (
		\P3_uWord_reg[6]/NET0131 ,
		\datao[22]_pad ,
		_w9977_,
		_w9978_,
		_w14814_
	);
	LUT3 #(
		.INIT('h2f)
	) name13465 (
		_w1945_,
		_w14813_,
		_w14814_,
		_w14815_
	);
	LUT2 #(
		.INIT('h2)
	) name13466 (
		\datao[25]_pad ,
		_w2115_,
		_w14816_
	);
	LUT3 #(
		.INIT('h10)
	) name13467 (
		_w2111_,
		_w14625_,
		_w14626_,
		_w14817_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13468 (
		\P3_uWord_reg[9]/NET0131 ,
		\datao[25]_pad ,
		_w9977_,
		_w9978_,
		_w14818_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13469 (
		_w1945_,
		_w14816_,
		_w14817_,
		_w14818_,
		_w14819_
	);
	LUT2 #(
		.INIT('h4)
	) name13470 (
		_w2105_,
		_w13903_,
		_w14820_
	);
	LUT2 #(
		.INIT('h8)
	) name13471 (
		_w14577_,
		_w14820_,
		_w14821_
	);
	LUT2 #(
		.INIT('h8)
	) name13472 (
		\P3_uWord_reg[10]/NET0131 ,
		_w9977_,
		_w14822_
	);
	LUT4 #(
		.INIT('h08aa)
	) name13473 (
		\datao[26]_pad ,
		_w1945_,
		_w2115_,
		_w9978_,
		_w14823_
	);
	LUT3 #(
		.INIT('hfe)
	) name13474 (
		_w14822_,
		_w14823_,
		_w14821_,
		_w14824_
	);
	LUT2 #(
		.INIT('h2)
	) name13475 (
		\datao[29]_pad ,
		_w2115_,
		_w14825_
	);
	LUT4 #(
		.INIT('h1020)
	) name13476 (
		\P3_EAX_reg[29]/NET0131 ,
		_w2111_,
		_w9543_,
		_w9544_,
		_w14826_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13477 (
		\P3_uWord_reg[13]/NET0131 ,
		\datao[29]_pad ,
		_w9977_,
		_w9978_,
		_w14827_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13478 (
		_w1945_,
		_w14825_,
		_w14826_,
		_w14827_,
		_w14828_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name13479 (
		\P1_Datao_reg[29]/NET0131 ,
		_w1860_,
		_w1931_,
		_w14508_,
		_w14829_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13480 (
		\P1_Datao_reg[29]/NET0131 ,
		\P1_uWord_reg[13]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14830_
	);
	LUT3 #(
		.INIT('h2f)
	) name13481 (
		_w1933_,
		_w14829_,
		_w14830_,
		_w14831_
	);
	LUT4 #(
		.INIT('h0200)
	) name13482 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w14471_,
		_w14832_
	);
	LUT4 #(
		.INIT('h0075)
	) name13483 (
		\P2_Datao_reg[16]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14832_,
		_w14833_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13484 (
		\P2_Datao_reg[16]/NET0131 ,
		\P2_uWord_reg[0]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14834_
	);
	LUT3 #(
		.INIT('h2f)
	) name13485 (
		_w1678_,
		_w14833_,
		_w14834_,
		_w14835_
	);
	LUT4 #(
		.INIT('h0200)
	) name13486 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w14494_,
		_w14836_
	);
	LUT4 #(
		.INIT('h0075)
	) name13487 (
		\P2_Datao_reg[17]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14836_,
		_w14837_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13488 (
		\P2_Datao_reg[17]/NET0131 ,
		\P2_uWord_reg[1]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14838_
	);
	LUT3 #(
		.INIT('h2f)
	) name13489 (
		_w1678_,
		_w14837_,
		_w14838_,
		_w14839_
	);
	LUT4 #(
		.INIT('h0200)
	) name13490 (
		_w1566_,
		_w1602_,
		_w1611_,
		_w14503_,
		_w14840_
	);
	LUT4 #(
		.INIT('h0075)
	) name13491 (
		\P2_Datao_reg[18]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14840_,
		_w14841_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13492 (
		\P2_Datao_reg[18]/NET0131 ,
		\P2_uWord_reg[2]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14842_
	);
	LUT3 #(
		.INIT('h2f)
	) name13493 (
		_w1678_,
		_w14841_,
		_w14842_,
		_w14843_
	);
	LUT3 #(
		.INIT('h8a)
	) name13494 (
		\P2_Datao_reg[21]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14844_
	);
	LUT2 #(
		.INIT('h4)
	) name13495 (
		_w1611_,
		_w14517_,
		_w14845_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13496 (
		\P2_Datao_reg[21]/NET0131 ,
		\P2_uWord_reg[5]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14846_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13497 (
		_w1678_,
		_w14844_,
		_w14845_,
		_w14846_,
		_w14847_
	);
	LUT4 #(
		.INIT('h0903)
	) name13498 (
		\P2_EAX_reg[21]/NET0131 ,
		\P2_EAX_reg[22]/NET0131 ,
		_w1611_,
		_w9459_,
		_w14848_
	);
	LUT4 #(
		.INIT('h5445)
	) name13499 (
		\P2_Datao_reg[22]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w14849_
	);
	LUT4 #(
		.INIT('h0002)
	) name13500 (
		_w1566_,
		_w1602_,
		_w14848_,
		_w14849_,
		_w14850_
	);
	LUT4 #(
		.INIT('h005d)
	) name13501 (
		\P2_Datao_reg[22]/NET0131 ,
		_w4927_,
		_w9989_,
		_w14850_,
		_w14851_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13502 (
		\P2_Datao_reg[22]/NET0131 ,
		\P2_uWord_reg[6]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14852_
	);
	LUT3 #(
		.INIT('h2f)
	) name13503 (
		_w1678_,
		_w14851_,
		_w14852_,
		_w14853_
	);
	LUT3 #(
		.INIT('h8a)
	) name13504 (
		\P2_Datao_reg[25]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14854_
	);
	LUT3 #(
		.INIT('h10)
	) name13505 (
		_w1611_,
		_w14545_,
		_w14546_,
		_w14855_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13506 (
		\P2_Datao_reg[25]/NET0131 ,
		\P2_uWord_reg[9]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14856_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13507 (
		_w1678_,
		_w14854_,
		_w14855_,
		_w14856_,
		_w14857_
	);
	LUT4 #(
		.INIT('h4f00)
	) name13508 (
		_w1602_,
		_w1616_,
		_w1678_,
		_w9996_,
		_w14858_
	);
	LUT2 #(
		.INIT('h8)
	) name13509 (
		\P2_uWord_reg[10]/NET0131 ,
		_w9995_,
		_w14859_
	);
	LUT4 #(
		.INIT('h0d00)
	) name13510 (
		_w1592_,
		_w1601_,
		_w1611_,
		_w1678_,
		_w14860_
	);
	LUT4 #(
		.INIT('h4800)
	) name13511 (
		\P2_EAX_reg[26]/NET0131 ,
		_w1566_,
		_w9460_,
		_w14860_,
		_w14861_
	);
	LUT2 #(
		.INIT('h1)
	) name13512 (
		_w14859_,
		_w14861_,
		_w14862_
	);
	LUT3 #(
		.INIT('h2f)
	) name13513 (
		\P2_Datao_reg[26]/NET0131 ,
		_w14858_,
		_w14862_,
		_w14863_
	);
	LUT3 #(
		.INIT('h8a)
	) name13514 (
		\P2_Datao_reg[29]/NET0131 ,
		_w1602_,
		_w1616_,
		_w14864_
	);
	LUT3 #(
		.INIT('h60)
	) name13515 (
		\P2_EAX_reg[29]/NET0131 ,
		_w9462_,
		_w9465_,
		_w14865_
	);
	LUT4 #(
		.INIT('h1200)
	) name13516 (
		\P2_EAX_reg[29]/NET0131 ,
		_w1611_,
		_w9462_,
		_w9465_,
		_w14866_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13517 (
		\P2_Datao_reg[29]/NET0131 ,
		\P2_uWord_reg[13]/NET0131 ,
		_w9995_,
		_w9996_,
		_w14867_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name13518 (
		_w1678_,
		_w14864_,
		_w14866_,
		_w14867_,
		_w14868_
	);
	LUT4 #(
		.INIT('h0200)
	) name13519 (
		_w1797_,
		_w1852_,
		_w1858_,
		_w14461_,
		_w14869_
	);
	LUT4 #(
		.INIT('hf020)
	) name13520 (
		\P1_Datao_reg[16]/NET0131 ,
		_w1860_,
		_w1933_,
		_w14869_,
		_w14870_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13521 (
		\P1_Datao_reg[16]/NET0131 ,
		\P1_uWord_reg[0]/NET0131 ,
		_w1935_,
		_w9972_,
		_w14871_
	);
	LUT2 #(
		.INIT('hb)
	) name13522 (
		_w14870_,
		_w14871_,
		_w14872_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13523 (
		\P3_lWord_reg[0]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14873_
	);
	LUT3 #(
		.INIT('h04)
	) name13524 (
		_w2060_,
		_w2047_,
		_w14873_,
		_w14874_
	);
	LUT4 #(
		.INIT('h0080)
	) name13525 (
		\P3_EAX_reg[0]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14875_
	);
	LUT3 #(
		.INIT('ha2)
	) name13526 (
		\P3_lWord_reg[0]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14876_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13527 (
		_w1945_,
		_w14875_,
		_w14874_,
		_w14876_,
		_w14877_
	);
	LUT2 #(
		.INIT('h2)
	) name13528 (
		\P3_lWord_reg[0]/NET0131 ,
		_w8341_,
		_w14878_
	);
	LUT2 #(
		.INIT('he)
	) name13529 (
		_w14877_,
		_w14878_,
		_w14879_
	);
	LUT3 #(
		.INIT('ha2)
	) name13530 (
		\P3_lWord_reg[10]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14880_
	);
	LUT4 #(
		.INIT('h0080)
	) name13531 (
		\P3_EAX_reg[10]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14881_
	);
	LUT4 #(
		.INIT('h2000)
	) name13532 (
		\buf2_reg[10]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2119_,
		_w14882_
	);
	LUT3 #(
		.INIT('ha8)
	) name13533 (
		_w1945_,
		_w14881_,
		_w14882_,
		_w14883_
	);
	LUT2 #(
		.INIT('he)
	) name13534 (
		_w14880_,
		_w14883_,
		_w14884_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13535 (
		\P3_lWord_reg[11]/NET0131 ,
		\buf2_reg[11]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14885_
	);
	LUT3 #(
		.INIT('h04)
	) name13536 (
		_w2060_,
		_w2047_,
		_w14885_,
		_w14886_
	);
	LUT4 #(
		.INIT('h0080)
	) name13537 (
		\P3_EAX_reg[11]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14887_
	);
	LUT3 #(
		.INIT('ha2)
	) name13538 (
		\P3_lWord_reg[11]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14888_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13539 (
		_w1945_,
		_w14887_,
		_w14886_,
		_w14888_,
		_w14889_
	);
	LUT2 #(
		.INIT('h2)
	) name13540 (
		\P3_lWord_reg[11]/NET0131 ,
		_w8341_,
		_w14890_
	);
	LUT2 #(
		.INIT('he)
	) name13541 (
		_w14889_,
		_w14890_,
		_w14891_
	);
	LUT3 #(
		.INIT('ha2)
	) name13542 (
		\P3_lWord_reg[12]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14892_
	);
	LUT4 #(
		.INIT('h0080)
	) name13543 (
		\P3_EAX_reg[12]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14893_
	);
	LUT3 #(
		.INIT('ha8)
	) name13544 (
		_w1945_,
		_w9532_,
		_w14893_,
		_w14894_
	);
	LUT2 #(
		.INIT('he)
	) name13545 (
		_w14892_,
		_w14894_,
		_w14895_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13546 (
		\P3_lWord_reg[13]/NET0131 ,
		\buf2_reg[13]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14896_
	);
	LUT3 #(
		.INIT('h04)
	) name13547 (
		_w2060_,
		_w2047_,
		_w14896_,
		_w14897_
	);
	LUT4 #(
		.INIT('h0080)
	) name13548 (
		\P3_EAX_reg[13]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14898_
	);
	LUT3 #(
		.INIT('ha2)
	) name13549 (
		\P3_lWord_reg[13]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14899_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13550 (
		_w1945_,
		_w14898_,
		_w14897_,
		_w14899_,
		_w14900_
	);
	LUT2 #(
		.INIT('h2)
	) name13551 (
		\P3_lWord_reg[13]/NET0131 ,
		_w8341_,
		_w14901_
	);
	LUT2 #(
		.INIT('he)
	) name13552 (
		_w14900_,
		_w14901_,
		_w14902_
	);
	LUT3 #(
		.INIT('ha2)
	) name13553 (
		\P3_lWord_reg[14]/NET0131 ,
		_w8341_,
		_w9529_,
		_w14903_
	);
	LUT4 #(
		.INIT('h0080)
	) name13554 (
		\P3_EAX_reg[14]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14904_
	);
	LUT3 #(
		.INIT('ha8)
	) name13555 (
		_w1945_,
		_w14589_,
		_w14904_,
		_w14905_
	);
	LUT2 #(
		.INIT('he)
	) name13556 (
		_w14903_,
		_w14905_,
		_w14906_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13557 (
		\P3_lWord_reg[15]/NET0131 ,
		\buf2_reg[15]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14907_
	);
	LUT3 #(
		.INIT('h04)
	) name13558 (
		_w2060_,
		_w2047_,
		_w14907_,
		_w14908_
	);
	LUT4 #(
		.INIT('h0080)
	) name13559 (
		\P3_EAX_reg[15]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14909_
	);
	LUT3 #(
		.INIT('ha2)
	) name13560 (
		\P3_lWord_reg[15]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14910_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13561 (
		_w1945_,
		_w14909_,
		_w14908_,
		_w14910_,
		_w14911_
	);
	LUT2 #(
		.INIT('h2)
	) name13562 (
		\P3_lWord_reg[15]/NET0131 ,
		_w8341_,
		_w14912_
	);
	LUT2 #(
		.INIT('he)
	) name13563 (
		_w14911_,
		_w14912_,
		_w14913_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13564 (
		\P3_lWord_reg[1]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14914_
	);
	LUT3 #(
		.INIT('h04)
	) name13565 (
		_w2060_,
		_w2047_,
		_w14914_,
		_w14915_
	);
	LUT4 #(
		.INIT('h0080)
	) name13566 (
		\P3_EAX_reg[1]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14916_
	);
	LUT3 #(
		.INIT('ha2)
	) name13567 (
		\P3_lWord_reg[1]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14917_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13568 (
		_w1945_,
		_w14916_,
		_w14915_,
		_w14917_,
		_w14918_
	);
	LUT2 #(
		.INIT('h2)
	) name13569 (
		\P3_lWord_reg[1]/NET0131 ,
		_w8341_,
		_w14919_
	);
	LUT2 #(
		.INIT('he)
	) name13570 (
		_w14918_,
		_w14919_,
		_w14920_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13571 (
		\P3_lWord_reg[2]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14921_
	);
	LUT3 #(
		.INIT('h04)
	) name13572 (
		_w2060_,
		_w2047_,
		_w14921_,
		_w14922_
	);
	LUT4 #(
		.INIT('h0080)
	) name13573 (
		\P3_EAX_reg[2]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14923_
	);
	LUT3 #(
		.INIT('ha2)
	) name13574 (
		\P3_lWord_reg[2]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14924_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13575 (
		_w1945_,
		_w14923_,
		_w14922_,
		_w14924_,
		_w14925_
	);
	LUT2 #(
		.INIT('h2)
	) name13576 (
		\P3_lWord_reg[2]/NET0131 ,
		_w8341_,
		_w14926_
	);
	LUT2 #(
		.INIT('he)
	) name13577 (
		_w14925_,
		_w14926_,
		_w14927_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13578 (
		\P3_lWord_reg[3]/NET0131 ,
		\buf2_reg[3]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14928_
	);
	LUT3 #(
		.INIT('h04)
	) name13579 (
		_w2060_,
		_w2047_,
		_w14928_,
		_w14929_
	);
	LUT4 #(
		.INIT('h0080)
	) name13580 (
		\P3_EAX_reg[3]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14930_
	);
	LUT3 #(
		.INIT('ha2)
	) name13581 (
		\P3_lWord_reg[3]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14931_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13582 (
		_w1945_,
		_w14930_,
		_w14929_,
		_w14931_,
		_w14932_
	);
	LUT2 #(
		.INIT('h2)
	) name13583 (
		\P3_lWord_reg[3]/NET0131 ,
		_w8341_,
		_w14933_
	);
	LUT2 #(
		.INIT('he)
	) name13584 (
		_w14932_,
		_w14933_,
		_w14934_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13585 (
		\P3_lWord_reg[4]/NET0131 ,
		\buf2_reg[4]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14935_
	);
	LUT3 #(
		.INIT('h04)
	) name13586 (
		_w2060_,
		_w2047_,
		_w14935_,
		_w14936_
	);
	LUT4 #(
		.INIT('h0080)
	) name13587 (
		\P3_EAX_reg[4]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14937_
	);
	LUT3 #(
		.INIT('ha2)
	) name13588 (
		\P3_lWord_reg[4]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14938_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13589 (
		_w1945_,
		_w14937_,
		_w14936_,
		_w14938_,
		_w14939_
	);
	LUT2 #(
		.INIT('h2)
	) name13590 (
		\P3_lWord_reg[4]/NET0131 ,
		_w8341_,
		_w14940_
	);
	LUT2 #(
		.INIT('he)
	) name13591 (
		_w14939_,
		_w14940_,
		_w14941_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13592 (
		\P3_lWord_reg[5]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14942_
	);
	LUT3 #(
		.INIT('h04)
	) name13593 (
		_w2060_,
		_w2047_,
		_w14942_,
		_w14943_
	);
	LUT4 #(
		.INIT('h0080)
	) name13594 (
		\P3_EAX_reg[5]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14944_
	);
	LUT3 #(
		.INIT('ha2)
	) name13595 (
		\P3_lWord_reg[5]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14945_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13596 (
		_w1945_,
		_w14944_,
		_w14943_,
		_w14945_,
		_w14946_
	);
	LUT2 #(
		.INIT('h2)
	) name13597 (
		\P3_lWord_reg[5]/NET0131 ,
		_w8341_,
		_w14947_
	);
	LUT2 #(
		.INIT('he)
	) name13598 (
		_w14946_,
		_w14947_,
		_w14948_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13599 (
		\P3_lWord_reg[6]/NET0131 ,
		\buf2_reg[6]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14949_
	);
	LUT3 #(
		.INIT('h04)
	) name13600 (
		_w2060_,
		_w2047_,
		_w14949_,
		_w14950_
	);
	LUT4 #(
		.INIT('h0080)
	) name13601 (
		\P3_EAX_reg[6]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14951_
	);
	LUT3 #(
		.INIT('ha2)
	) name13602 (
		\P3_lWord_reg[6]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14952_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13603 (
		_w1945_,
		_w14951_,
		_w14950_,
		_w14952_,
		_w14953_
	);
	LUT2 #(
		.INIT('h2)
	) name13604 (
		\P3_lWord_reg[6]/NET0131 ,
		_w8341_,
		_w14954_
	);
	LUT2 #(
		.INIT('he)
	) name13605 (
		_w14953_,
		_w14954_,
		_w14955_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13606 (
		\P3_lWord_reg[7]/NET0131 ,
		\buf2_reg[7]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14956_
	);
	LUT3 #(
		.INIT('h04)
	) name13607 (
		_w2060_,
		_w2047_,
		_w14956_,
		_w14957_
	);
	LUT4 #(
		.INIT('h0080)
	) name13608 (
		\P3_EAX_reg[7]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14958_
	);
	LUT3 #(
		.INIT('ha2)
	) name13609 (
		\P3_lWord_reg[7]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14959_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13610 (
		_w1945_,
		_w14958_,
		_w14957_,
		_w14959_,
		_w14960_
	);
	LUT2 #(
		.INIT('h2)
	) name13611 (
		\P3_lWord_reg[7]/NET0131 ,
		_w8341_,
		_w14961_
	);
	LUT2 #(
		.INIT('he)
	) name13612 (
		_w14960_,
		_w14961_,
		_w14962_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13613 (
		\P3_lWord_reg[8]/NET0131 ,
		\buf2_reg[8]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14963_
	);
	LUT3 #(
		.INIT('h04)
	) name13614 (
		_w2060_,
		_w2047_,
		_w14963_,
		_w14964_
	);
	LUT3 #(
		.INIT('ha2)
	) name13615 (
		\P3_lWord_reg[8]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14965_
	);
	LUT4 #(
		.INIT('h0080)
	) name13616 (
		\P3_EAX_reg[8]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14966_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13617 (
		_w1945_,
		_w14965_,
		_w14964_,
		_w14966_,
		_w14967_
	);
	LUT2 #(
		.INIT('h2)
	) name13618 (
		\P3_lWord_reg[8]/NET0131 ,
		_w8341_,
		_w14968_
	);
	LUT2 #(
		.INIT('he)
	) name13619 (
		_w14967_,
		_w14968_,
		_w14969_
	);
	LUT4 #(
		.INIT('h55f3)
	) name13620 (
		\P3_lWord_reg[9]/NET0131 ,
		\buf2_reg[9]/NET0131 ,
		_w2105_,
		_w2116_,
		_w14970_
	);
	LUT3 #(
		.INIT('h04)
	) name13621 (
		_w2060_,
		_w2047_,
		_w14970_,
		_w14971_
	);
	LUT4 #(
		.INIT('h0080)
	) name13622 (
		\P3_EAX_reg[9]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w14972_
	);
	LUT3 #(
		.INIT('ha2)
	) name13623 (
		\P3_lWord_reg[9]/NET0131 ,
		_w2047_,
		_w2105_,
		_w14973_
	);
	LUT4 #(
		.INIT('haaa8)
	) name13624 (
		_w1945_,
		_w14972_,
		_w14971_,
		_w14973_,
		_w14974_
	);
	LUT2 #(
		.INIT('h2)
	) name13625 (
		\P3_lWord_reg[9]/NET0131 ,
		_w8341_,
		_w14975_
	);
	LUT2 #(
		.INIT('he)
	) name13626 (
		_w14974_,
		_w14975_,
		_w14976_
	);
	LUT3 #(
		.INIT('hc8)
	) name13627 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		_w2215_,
		_w10611_,
		_w14977_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13628 (
		_w2011_,
		_w2016_,
		_w10611_,
		_w14977_,
		_w14978_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13629 (
		\P3_InstQueue_reg[0][2]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w14979_
	);
	LUT4 #(
		.INIT('h153f)
	) name13630 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10614_,
		_w10616_,
		_w14980_
	);
	LUT2 #(
		.INIT('h2)
	) name13631 (
		_w2199_,
		_w14980_,
		_w14981_
	);
	LUT3 #(
		.INIT('h02)
	) name13632 (
		\buf2_reg[2]/NET0131 ,
		_w10618_,
		_w10621_,
		_w14982_
	);
	LUT3 #(
		.INIT('h01)
	) name13633 (
		_w14979_,
		_w14981_,
		_w14982_,
		_w14983_
	);
	LUT2 #(
		.INIT('hb)
	) name13634 (
		_w14978_,
		_w14983_,
		_w14984_
	);
	LUT3 #(
		.INIT('hc8)
	) name13635 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		_w2215_,
		_w10630_,
		_w14985_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13636 (
		_w2011_,
		_w2016_,
		_w10630_,
		_w14985_,
		_w14986_
	);
	LUT4 #(
		.INIT('h222a)
	) name13637 (
		\P3_InstQueue_reg[10][2]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w14987_
	);
	LUT4 #(
		.INIT('h153f)
	) name13638 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10633_,
		_w10635_,
		_w14988_
	);
	LUT2 #(
		.INIT('h2)
	) name13639 (
		_w2199_,
		_w14988_,
		_w14989_
	);
	LUT3 #(
		.INIT('h20)
	) name13640 (
		\buf2_reg[2]/NET0131 ,
		_w10637_,
		_w10639_,
		_w14990_
	);
	LUT3 #(
		.INIT('h01)
	) name13641 (
		_w14987_,
		_w14989_,
		_w14990_,
		_w14991_
	);
	LUT2 #(
		.INIT('hb)
	) name13642 (
		_w14986_,
		_w14991_,
		_w14992_
	);
	LUT3 #(
		.INIT('hc8)
	) name13643 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w2215_,
		_w10646_,
		_w14993_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13644 (
		_w2011_,
		_w2016_,
		_w10646_,
		_w14993_,
		_w14994_
	);
	LUT3 #(
		.INIT('ha2)
	) name13645 (
		\P3_InstQueue_reg[11][2]/NET0131 ,
		_w10622_,
		_w10650_,
		_w14995_
	);
	LUT3 #(
		.INIT('hd8)
	) name13646 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w14996_
	);
	LUT3 #(
		.INIT('h80)
	) name13647 (
		_w2194_,
		_w10649_,
		_w14996_,
		_w14997_
	);
	LUT4 #(
		.INIT('h2000)
	) name13648 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w14998_
	);
	LUT4 #(
		.INIT('hce00)
	) name13649 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w14998_,
		_w14999_
	);
	LUT2 #(
		.INIT('h1)
	) name13650 (
		_w14997_,
		_w14999_,
		_w15000_
	);
	LUT2 #(
		.INIT('h4)
	) name13651 (
		_w14995_,
		_w15000_,
		_w15001_
	);
	LUT2 #(
		.INIT('hb)
	) name13652 (
		_w14994_,
		_w15001_,
		_w15002_
	);
	LUT3 #(
		.INIT('hc8)
	) name13653 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w2215_,
		_w10659_,
		_w15003_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13654 (
		_w2011_,
		_w2016_,
		_w10659_,
		_w15003_,
		_w15004_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13655 (
		\P3_InstQueue_reg[12][2]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w15005_
	);
	LUT4 #(
		.INIT('h135f)
	) name13656 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10630_,
		_w10652_,
		_w15006_
	);
	LUT2 #(
		.INIT('h2)
	) name13657 (
		_w2199_,
		_w15006_,
		_w15007_
	);
	LUT3 #(
		.INIT('h02)
	) name13658 (
		\buf2_reg[2]/NET0131 ,
		_w10662_,
		_w10663_,
		_w15008_
	);
	LUT3 #(
		.INIT('h01)
	) name13659 (
		_w15005_,
		_w15007_,
		_w15008_,
		_w15009_
	);
	LUT2 #(
		.INIT('hb)
	) name13660 (
		_w15004_,
		_w15009_,
		_w15010_
	);
	LUT3 #(
		.INIT('hc8)
	) name13661 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w2215_,
		_w10614_,
		_w15011_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13662 (
		_w2011_,
		_w2016_,
		_w10614_,
		_w15011_,
		_w15012_
	);
	LUT2 #(
		.INIT('h4)
	) name13663 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w10672_,
		_w15013_
	);
	LUT2 #(
		.INIT('h1)
	) name13664 (
		\buf2_reg[2]/NET0131 ,
		_w10672_,
		_w15014_
	);
	LUT3 #(
		.INIT('h02)
	) name13665 (
		_w10674_,
		_w15014_,
		_w15013_,
		_w15015_
	);
	LUT2 #(
		.INIT('h2)
	) name13666 (
		\P3_InstQueue_reg[13][2]/NET0131 ,
		_w10622_,
		_w15016_
	);
	LUT3 #(
		.INIT('h80)
	) name13667 (
		_w2194_,
		_w10673_,
		_w14996_,
		_w15017_
	);
	LUT2 #(
		.INIT('h1)
	) name13668 (
		_w15016_,
		_w15017_,
		_w15018_
	);
	LUT2 #(
		.INIT('h4)
	) name13669 (
		_w15015_,
		_w15018_,
		_w15019_
	);
	LUT2 #(
		.INIT('hb)
	) name13670 (
		_w15012_,
		_w15019_,
		_w15020_
	);
	LUT3 #(
		.INIT('hc8)
	) name13671 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w2215_,
		_w10616_,
		_w15021_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13672 (
		_w2011_,
		_w2016_,
		_w10616_,
		_w15021_,
		_w15022_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name13673 (
		\P3_InstQueue_reg[14][2]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w15023_
	);
	LUT4 #(
		.INIT('h153f)
	) name13674 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10646_,
		_w10659_,
		_w15024_
	);
	LUT2 #(
		.INIT('h2)
	) name13675 (
		_w2199_,
		_w15024_,
		_w15025_
	);
	LUT3 #(
		.INIT('h02)
	) name13676 (
		\buf2_reg[2]/NET0131 ,
		_w10617_,
		_w10684_,
		_w15026_
	);
	LUT3 #(
		.INIT('h01)
	) name13677 (
		_w15023_,
		_w15025_,
		_w15026_,
		_w15027_
	);
	LUT2 #(
		.INIT('hb)
	) name13678 (
		_w15022_,
		_w15027_,
		_w15028_
	);
	LUT3 #(
		.INIT('hc8)
	) name13679 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w2215_,
		_w10620_,
		_w15029_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13680 (
		_w2011_,
		_w2016_,
		_w10620_,
		_w15029_,
		_w15030_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13681 (
		\P3_InstQueue_reg[15][2]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w15031_
	);
	LUT4 #(
		.INIT('h135f)
	) name13682 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10614_,
		_w10659_,
		_w15032_
	);
	LUT2 #(
		.INIT('h2)
	) name13683 (
		_w2199_,
		_w15032_,
		_w15033_
	);
	LUT3 #(
		.INIT('h02)
	) name13684 (
		\buf2_reg[2]/NET0131 ,
		_w10693_,
		_w10694_,
		_w15034_
	);
	LUT3 #(
		.INIT('h01)
	) name13685 (
		_w15031_,
		_w15033_,
		_w15034_,
		_w15035_
	);
	LUT2 #(
		.INIT('hb)
	) name13686 (
		_w15030_,
		_w15035_,
		_w15036_
	);
	LUT3 #(
		.INIT('hc8)
	) name13687 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w2215_,
		_w10701_,
		_w15037_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13688 (
		_w2011_,
		_w2016_,
		_w10701_,
		_w15037_,
		_w15038_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13689 (
		\P3_InstQueue_reg[1][2]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w15039_
	);
	LUT4 #(
		.INIT('h153f)
	) name13690 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10616_,
		_w10620_,
		_w15040_
	);
	LUT2 #(
		.INIT('h2)
	) name13691 (
		_w2199_,
		_w15040_,
		_w15041_
	);
	LUT3 #(
		.INIT('h02)
	) name13692 (
		\buf2_reg[2]/NET0131 ,
		_w10704_,
		_w10705_,
		_w15042_
	);
	LUT3 #(
		.INIT('h01)
	) name13693 (
		_w15039_,
		_w15041_,
		_w15042_,
		_w15043_
	);
	LUT2 #(
		.INIT('hb)
	) name13694 (
		_w15038_,
		_w15043_,
		_w15044_
	);
	LUT3 #(
		.INIT('hc8)
	) name13695 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w2215_,
		_w10713_,
		_w15045_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13696 (
		_w2011_,
		_w2016_,
		_w10713_,
		_w15045_,
		_w15046_
	);
	LUT4 #(
		.INIT('h222a)
	) name13697 (
		\P3_InstQueue_reg[2][2]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w15047_
	);
	LUT4 #(
		.INIT('h135f)
	) name13698 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10611_,
		_w10620_,
		_w15048_
	);
	LUT2 #(
		.INIT('h2)
	) name13699 (
		_w2199_,
		_w15048_,
		_w15049_
	);
	LUT3 #(
		.INIT('h20)
	) name13700 (
		\buf2_reg[2]/NET0131 ,
		_w10716_,
		_w10717_,
		_w15050_
	);
	LUT3 #(
		.INIT('h01)
	) name13701 (
		_w15047_,
		_w15049_,
		_w15050_,
		_w15051_
	);
	LUT2 #(
		.INIT('hb)
	) name13702 (
		_w15046_,
		_w15051_,
		_w15052_
	);
	LUT3 #(
		.INIT('hc8)
	) name13703 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w2215_,
		_w10724_,
		_w15053_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13704 (
		_w2011_,
		_w2016_,
		_w10724_,
		_w15053_,
		_w15054_
	);
	LUT4 #(
		.INIT('h222a)
	) name13705 (
		\P3_InstQueue_reg[3][2]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w15055_
	);
	LUT4 #(
		.INIT('h153f)
	) name13706 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10611_,
		_w10701_,
		_w15056_
	);
	LUT2 #(
		.INIT('h2)
	) name13707 (
		_w2199_,
		_w15056_,
		_w15057_
	);
	LUT3 #(
		.INIT('h08)
	) name13708 (
		\buf2_reg[2]/NET0131 ,
		_w10712_,
		_w10727_,
		_w15058_
	);
	LUT3 #(
		.INIT('h01)
	) name13709 (
		_w15055_,
		_w15057_,
		_w15058_,
		_w15059_
	);
	LUT2 #(
		.INIT('hb)
	) name13710 (
		_w15054_,
		_w15059_,
		_w15060_
	);
	LUT3 #(
		.INIT('hc8)
	) name13711 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w2215_,
		_w10734_,
		_w15061_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13712 (
		_w2011_,
		_w2016_,
		_w10734_,
		_w15061_,
		_w15062_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13713 (
		\P3_InstQueue_reg[4][2]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w15063_
	);
	LUT4 #(
		.INIT('h153f)
	) name13714 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10701_,
		_w10713_,
		_w15064_
	);
	LUT2 #(
		.INIT('h2)
	) name13715 (
		_w2199_,
		_w15064_,
		_w15065_
	);
	LUT3 #(
		.INIT('h02)
	) name13716 (
		\buf2_reg[2]/NET0131 ,
		_w10737_,
		_w10738_,
		_w15066_
	);
	LUT3 #(
		.INIT('h01)
	) name13717 (
		_w15063_,
		_w15065_,
		_w15066_,
		_w15067_
	);
	LUT2 #(
		.INIT('hb)
	) name13718 (
		_w15062_,
		_w15067_,
		_w15068_
	);
	LUT3 #(
		.INIT('hc8)
	) name13719 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w2215_,
		_w10745_,
		_w15069_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13720 (
		_w2011_,
		_w2016_,
		_w10745_,
		_w15069_,
		_w15070_
	);
	LUT2 #(
		.INIT('h4)
	) name13721 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w10748_,
		_w15071_
	);
	LUT2 #(
		.INIT('h1)
	) name13722 (
		\buf2_reg[2]/NET0131 ,
		_w10748_,
		_w15072_
	);
	LUT3 #(
		.INIT('h02)
	) name13723 (
		_w10750_,
		_w15072_,
		_w15071_,
		_w15073_
	);
	LUT2 #(
		.INIT('h2)
	) name13724 (
		\P3_InstQueue_reg[5][2]/NET0131 ,
		_w10622_,
		_w15074_
	);
	LUT3 #(
		.INIT('h80)
	) name13725 (
		_w2194_,
		_w10749_,
		_w14996_,
		_w15075_
	);
	LUT2 #(
		.INIT('h1)
	) name13726 (
		_w15074_,
		_w15075_,
		_w15076_
	);
	LUT2 #(
		.INIT('h4)
	) name13727 (
		_w15073_,
		_w15076_,
		_w15077_
	);
	LUT2 #(
		.INIT('hb)
	) name13728 (
		_w15070_,
		_w15077_,
		_w15078_
	);
	LUT3 #(
		.INIT('hc8)
	) name13729 (
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w2215_,
		_w10758_,
		_w15079_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13730 (
		_w2011_,
		_w2016_,
		_w10758_,
		_w15079_,
		_w15080_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13731 (
		\P3_InstQueue_reg[6][2]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w15081_
	);
	LUT4 #(
		.INIT('h153f)
	) name13732 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10724_,
		_w10734_,
		_w15082_
	);
	LUT2 #(
		.INIT('h2)
	) name13733 (
		_w2199_,
		_w15082_,
		_w15083_
	);
	LUT3 #(
		.INIT('h02)
	) name13734 (
		\buf2_reg[2]/NET0131 ,
		_w10761_,
		_w10762_,
		_w15084_
	);
	LUT3 #(
		.INIT('h01)
	) name13735 (
		_w15081_,
		_w15083_,
		_w15084_,
		_w15085_
	);
	LUT2 #(
		.INIT('hb)
	) name13736 (
		_w15080_,
		_w15085_,
		_w15086_
	);
	LUT3 #(
		.INIT('hc8)
	) name13737 (
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w2215_,
		_w10633_,
		_w15087_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13738 (
		_w2011_,
		_w2016_,
		_w10633_,
		_w15087_,
		_w15088_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13739 (
		\P3_InstQueue_reg[7][2]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w15089_
	);
	LUT4 #(
		.INIT('h153f)
	) name13740 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10734_,
		_w10745_,
		_w15090_
	);
	LUT2 #(
		.INIT('h2)
	) name13741 (
		_w2199_,
		_w15090_,
		_w15091_
	);
	LUT3 #(
		.INIT('h02)
	) name13742 (
		\buf2_reg[2]/NET0131 ,
		_w10771_,
		_w10772_,
		_w15092_
	);
	LUT3 #(
		.INIT('h01)
	) name13743 (
		_w15089_,
		_w15091_,
		_w15092_,
		_w15093_
	);
	LUT2 #(
		.INIT('hb)
	) name13744 (
		_w15088_,
		_w15093_,
		_w15094_
	);
	LUT3 #(
		.INIT('hc8)
	) name13745 (
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w2215_,
		_w10635_,
		_w15095_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13746 (
		_w2011_,
		_w2016_,
		_w10635_,
		_w15095_,
		_w15096_
	);
	LUT4 #(
		.INIT('h22a2)
	) name13747 (
		\P3_InstQueue_reg[8][2]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w15097_
	);
	LUT4 #(
		.INIT('h153f)
	) name13748 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10745_,
		_w10758_,
		_w15098_
	);
	LUT2 #(
		.INIT('h2)
	) name13749 (
		_w2199_,
		_w15098_,
		_w15099_
	);
	LUT3 #(
		.INIT('h02)
	) name13750 (
		\buf2_reg[2]/NET0131 ,
		_w10636_,
		_w10781_,
		_w15100_
	);
	LUT3 #(
		.INIT('h01)
	) name13751 (
		_w15097_,
		_w15099_,
		_w15100_,
		_w15101_
	);
	LUT2 #(
		.INIT('hb)
	) name13752 (
		_w15096_,
		_w15101_,
		_w15102_
	);
	LUT3 #(
		.INIT('hc8)
	) name13753 (
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w2215_,
		_w10652_,
		_w15103_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13754 (
		_w2011_,
		_w2016_,
		_w10652_,
		_w15103_,
		_w15104_
	);
	LUT4 #(
		.INIT('h135f)
	) name13755 (
		\buf2_reg[18]/NET0131 ,
		\buf2_reg[26]/NET0131 ,
		_w10633_,
		_w10758_,
		_w15105_
	);
	LUT4 #(
		.INIT('hef00)
	) name13756 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w15106_
	);
	LUT4 #(
		.INIT('h1000)
	) name13757 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[2]/NET0131 ,
		_w15107_
	);
	LUT4 #(
		.INIT('hddd0)
	) name13758 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w15106_,
		_w15107_,
		_w15108_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13759 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w15105_,
		_w15108_,
		_w15109_
	);
	LUT3 #(
		.INIT('ha8)
	) name13760 (
		_w3055_,
		_w15106_,
		_w15107_,
		_w15110_
	);
	LUT2 #(
		.INIT('h2)
	) name13761 (
		\P3_InstQueue_reg[9][2]/NET0131 ,
		_w10622_,
		_w15111_
	);
	LUT2 #(
		.INIT('h1)
	) name13762 (
		_w15110_,
		_w15111_,
		_w15112_
	);
	LUT2 #(
		.INIT('h4)
	) name13763 (
		_w15109_,
		_w15112_,
		_w15113_
	);
	LUT2 #(
		.INIT('hb)
	) name13764 (
		_w15104_,
		_w15113_,
		_w15114_
	);
	LUT4 #(
		.INIT('hca00)
	) name13765 (
		\P1_Datao_reg[1]/NET0131 ,
		\P1_EAX_reg[1]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15115_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13766 (
		\P1_Datao_reg[1]/NET0131 ,
		\P1_lWord_reg[1]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15116_
	);
	LUT2 #(
		.INIT('hb)
	) name13767 (
		_w15115_,
		_w15116_,
		_w15117_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13768 (
		\P3_EAX_reg[0]/NET0131 ,
		\datao[0]_pad ,
		_w1945_,
		_w2115_,
		_w15118_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13769 (
		\P3_lWord_reg[0]/NET0131 ,
		\datao[0]_pad ,
		_w9977_,
		_w9978_,
		_w15119_
	);
	LUT2 #(
		.INIT('hb)
	) name13770 (
		_w15118_,
		_w15119_,
		_w15120_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13771 (
		\P3_EAX_reg[10]/NET0131 ,
		\datao[10]_pad ,
		_w1945_,
		_w2115_,
		_w15121_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13772 (
		\P3_lWord_reg[10]/NET0131 ,
		\datao[10]_pad ,
		_w9977_,
		_w9978_,
		_w15122_
	);
	LUT2 #(
		.INIT('hb)
	) name13773 (
		_w15121_,
		_w15122_,
		_w15123_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13774 (
		\P3_EAX_reg[11]/NET0131 ,
		\datao[11]_pad ,
		_w1945_,
		_w2115_,
		_w15124_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13775 (
		\P3_lWord_reg[11]/NET0131 ,
		\datao[11]_pad ,
		_w9977_,
		_w9978_,
		_w15125_
	);
	LUT2 #(
		.INIT('hb)
	) name13776 (
		_w15124_,
		_w15125_,
		_w15126_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13777 (
		\P3_EAX_reg[15]/NET0131 ,
		\datao[15]_pad ,
		_w1945_,
		_w2115_,
		_w15127_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13778 (
		\P3_lWord_reg[15]/NET0131 ,
		\datao[15]_pad ,
		_w9977_,
		_w9978_,
		_w15128_
	);
	LUT2 #(
		.INIT('hb)
	) name13779 (
		_w15127_,
		_w15128_,
		_w15129_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13780 (
		\P3_EAX_reg[1]/NET0131 ,
		\datao[1]_pad ,
		_w1945_,
		_w2115_,
		_w15130_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13781 (
		\P3_lWord_reg[1]/NET0131 ,
		\datao[1]_pad ,
		_w9977_,
		_w9978_,
		_w15131_
	);
	LUT2 #(
		.INIT('hb)
	) name13782 (
		_w15130_,
		_w15131_,
		_w15132_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13783 (
		\P3_EAX_reg[4]/NET0131 ,
		\datao[4]_pad ,
		_w1945_,
		_w2115_,
		_w15133_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13784 (
		\P3_lWord_reg[4]/NET0131 ,
		\datao[4]_pad ,
		_w9977_,
		_w9978_,
		_w15134_
	);
	LUT2 #(
		.INIT('hb)
	) name13785 (
		_w15133_,
		_w15134_,
		_w15135_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13786 (
		\P3_EAX_reg[5]/NET0131 ,
		\datao[5]_pad ,
		_w1945_,
		_w2115_,
		_w15136_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13787 (
		\P3_lWord_reg[5]/NET0131 ,
		\datao[5]_pad ,
		_w9977_,
		_w9978_,
		_w15137_
	);
	LUT2 #(
		.INIT('hb)
	) name13788 (
		_w15136_,
		_w15137_,
		_w15138_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13789 (
		\P3_EAX_reg[6]/NET0131 ,
		\datao[6]_pad ,
		_w1945_,
		_w2115_,
		_w15139_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13790 (
		\P3_lWord_reg[6]/NET0131 ,
		\datao[6]_pad ,
		_w9977_,
		_w9978_,
		_w15140_
	);
	LUT2 #(
		.INIT('hb)
	) name13791 (
		_w15139_,
		_w15140_,
		_w15141_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13792 (
		\P3_EAX_reg[7]/NET0131 ,
		\datao[7]_pad ,
		_w1945_,
		_w2115_,
		_w15142_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13793 (
		\P3_lWord_reg[7]/NET0131 ,
		\datao[7]_pad ,
		_w9977_,
		_w9978_,
		_w15143_
	);
	LUT2 #(
		.INIT('hb)
	) name13794 (
		_w15142_,
		_w15143_,
		_w15144_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13795 (
		\P3_EAX_reg[8]/NET0131 ,
		\datao[8]_pad ,
		_w1945_,
		_w2115_,
		_w15145_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13796 (
		\P3_lWord_reg[8]/NET0131 ,
		\datao[8]_pad ,
		_w9977_,
		_w9978_,
		_w15146_
	);
	LUT2 #(
		.INIT('hb)
	) name13797 (
		_w15145_,
		_w15146_,
		_w15147_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name13798 (
		\P3_EAX_reg[9]/NET0131 ,
		\datao[9]_pad ,
		_w1945_,
		_w2115_,
		_w15148_
	);
	LUT4 #(
		.INIT('h5f13)
	) name13799 (
		\P3_lWord_reg[9]/NET0131 ,
		\datao[9]_pad ,
		_w9977_,
		_w9978_,
		_w15149_
	);
	LUT2 #(
		.INIT('hb)
	) name13800 (
		_w15148_,
		_w15149_,
		_w15150_
	);
	LUT3 #(
		.INIT('h10)
	) name13801 (
		\P2_EAX_reg[13]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15151_
	);
	LUT4 #(
		.INIT('hba00)
	) name13802 (
		\P2_Datao_reg[13]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15152_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13803 (
		\P2_Datao_reg[13]/NET0131 ,
		\P2_lWord_reg[13]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15153_
	);
	LUT3 #(
		.INIT('h4f)
	) name13804 (
		_w15151_,
		_w15152_,
		_w15153_,
		_w15154_
	);
	LUT3 #(
		.INIT('h10)
	) name13805 (
		\P2_EAX_reg[14]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15155_
	);
	LUT4 #(
		.INIT('hba00)
	) name13806 (
		\P2_Datao_reg[14]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15156_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13807 (
		\P2_Datao_reg[14]/NET0131 ,
		\P2_lWord_reg[14]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15157_
	);
	LUT3 #(
		.INIT('h4f)
	) name13808 (
		_w15155_,
		_w15156_,
		_w15157_,
		_w15158_
	);
	LUT3 #(
		.INIT('h10)
	) name13809 (
		\P2_EAX_reg[15]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15159_
	);
	LUT4 #(
		.INIT('hba00)
	) name13810 (
		\P2_Datao_reg[15]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15160_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13811 (
		\P2_Datao_reg[15]/NET0131 ,
		\P2_lWord_reg[15]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15161_
	);
	LUT3 #(
		.INIT('h4f)
	) name13812 (
		_w15159_,
		_w15160_,
		_w15161_,
		_w15162_
	);
	LUT3 #(
		.INIT('h10)
	) name13813 (
		\P2_EAX_reg[1]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15163_
	);
	LUT4 #(
		.INIT('hba00)
	) name13814 (
		\P2_Datao_reg[1]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15164_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13815 (
		\P2_Datao_reg[1]/NET0131 ,
		\P2_lWord_reg[1]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15165_
	);
	LUT3 #(
		.INIT('h4f)
	) name13816 (
		_w15163_,
		_w15164_,
		_w15165_,
		_w15166_
	);
	LUT3 #(
		.INIT('h10)
	) name13817 (
		\P2_EAX_reg[2]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15167_
	);
	LUT4 #(
		.INIT('hba00)
	) name13818 (
		\P2_Datao_reg[2]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15168_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13819 (
		\P2_Datao_reg[2]/NET0131 ,
		\P2_lWord_reg[2]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15169_
	);
	LUT3 #(
		.INIT('h4f)
	) name13820 (
		_w15167_,
		_w15168_,
		_w15169_,
		_w15170_
	);
	LUT3 #(
		.INIT('h10)
	) name13821 (
		\P2_EAX_reg[3]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15171_
	);
	LUT4 #(
		.INIT('hba00)
	) name13822 (
		\P2_Datao_reg[3]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15172_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13823 (
		\P2_Datao_reg[3]/NET0131 ,
		\P2_lWord_reg[3]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15173_
	);
	LUT3 #(
		.INIT('h4f)
	) name13824 (
		_w15171_,
		_w15172_,
		_w15173_,
		_w15174_
	);
	LUT3 #(
		.INIT('h10)
	) name13825 (
		\P2_EAX_reg[4]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15175_
	);
	LUT4 #(
		.INIT('hba00)
	) name13826 (
		\P2_Datao_reg[4]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15176_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13827 (
		\P2_Datao_reg[4]/NET0131 ,
		\P2_lWord_reg[4]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15177_
	);
	LUT3 #(
		.INIT('h4f)
	) name13828 (
		_w15175_,
		_w15176_,
		_w15177_,
		_w15178_
	);
	LUT3 #(
		.INIT('h10)
	) name13829 (
		\P2_EAX_reg[6]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15179_
	);
	LUT4 #(
		.INIT('hba00)
	) name13830 (
		\P2_Datao_reg[6]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15180_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13831 (
		\P2_Datao_reg[6]/NET0131 ,
		\P2_lWord_reg[6]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15181_
	);
	LUT3 #(
		.INIT('h4f)
	) name13832 (
		_w15179_,
		_w15180_,
		_w15181_,
		_w15182_
	);
	LUT3 #(
		.INIT('h10)
	) name13833 (
		\P2_EAX_reg[9]/NET0131 ,
		_w1602_,
		_w1616_,
		_w15183_
	);
	LUT4 #(
		.INIT('hba00)
	) name13834 (
		\P2_Datao_reg[9]/NET0131 ,
		_w1602_,
		_w1616_,
		_w1678_,
		_w15184_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13835 (
		\P2_Datao_reg[9]/NET0131 ,
		\P2_lWord_reg[9]/NET0131 ,
		_w9995_,
		_w9996_,
		_w15185_
	);
	LUT3 #(
		.INIT('h4f)
	) name13836 (
		_w15183_,
		_w15184_,
		_w15185_,
		_w15186_
	);
	LUT4 #(
		.INIT('hca00)
	) name13837 (
		\P1_Datao_reg[3]/NET0131 ,
		\P1_EAX_reg[3]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15187_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13838 (
		\P1_Datao_reg[3]/NET0131 ,
		\P1_lWord_reg[3]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15188_
	);
	LUT2 #(
		.INIT('hb)
	) name13839 (
		_w15187_,
		_w15188_,
		_w15189_
	);
	LUT4 #(
		.INIT('hca00)
	) name13840 (
		\P1_Datao_reg[5]/NET0131 ,
		\P1_EAX_reg[5]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15190_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13841 (
		\P1_Datao_reg[5]/NET0131 ,
		\P1_lWord_reg[5]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15191_
	);
	LUT2 #(
		.INIT('hb)
	) name13842 (
		_w15190_,
		_w15191_,
		_w15192_
	);
	LUT4 #(
		.INIT('hca00)
	) name13843 (
		\P1_Datao_reg[7]/NET0131 ,
		\P1_EAX_reg[7]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15193_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13844 (
		\P1_Datao_reg[7]/NET0131 ,
		\P1_lWord_reg[7]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15194_
	);
	LUT2 #(
		.INIT('hb)
	) name13845 (
		_w15193_,
		_w15194_,
		_w15195_
	);
	LUT4 #(
		.INIT('hca00)
	) name13846 (
		\P1_Datao_reg[9]/NET0131 ,
		\P1_EAX_reg[9]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15196_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13847 (
		\P1_Datao_reg[9]/NET0131 ,
		\P1_lWord_reg[9]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15197_
	);
	LUT2 #(
		.INIT('hb)
	) name13848 (
		_w15196_,
		_w15197_,
		_w15198_
	);
	LUT4 #(
		.INIT('hca00)
	) name13849 (
		\P1_Datao_reg[0]/NET0131 ,
		\P1_EAX_reg[0]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15199_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13850 (
		\P1_Datao_reg[0]/NET0131 ,
		\P1_lWord_reg[0]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15200_
	);
	LUT2 #(
		.INIT('hb)
	) name13851 (
		_w15199_,
		_w15200_,
		_w15201_
	);
	LUT4 #(
		.INIT('hca00)
	) name13852 (
		\P1_Datao_reg[10]/NET0131 ,
		\P1_EAX_reg[10]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15202_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13853 (
		\P1_Datao_reg[10]/NET0131 ,
		\P1_lWord_reg[10]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15203_
	);
	LUT2 #(
		.INIT('hb)
	) name13854 (
		_w15202_,
		_w15203_,
		_w15204_
	);
	LUT4 #(
		.INIT('hca00)
	) name13855 (
		\P1_Datao_reg[11]/NET0131 ,
		\P1_EAX_reg[11]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15205_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13856 (
		\P1_Datao_reg[11]/NET0131 ,
		\P1_lWord_reg[11]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15206_
	);
	LUT2 #(
		.INIT('hb)
	) name13857 (
		_w15205_,
		_w15206_,
		_w15207_
	);
	LUT4 #(
		.INIT('hca00)
	) name13858 (
		\P1_Datao_reg[12]/NET0131 ,
		\P1_EAX_reg[12]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15208_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13859 (
		\P1_Datao_reg[12]/NET0131 ,
		\P1_lWord_reg[12]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15209_
	);
	LUT2 #(
		.INIT('hb)
	) name13860 (
		_w15208_,
		_w15209_,
		_w15210_
	);
	LUT4 #(
		.INIT('hca00)
	) name13861 (
		\P1_Datao_reg[13]/NET0131 ,
		\P1_EAX_reg[13]/NET0131 ,
		_w1860_,
		_w1933_,
		_w15211_
	);
	LUT4 #(
		.INIT('h3f15)
	) name13862 (
		\P1_Datao_reg[13]/NET0131 ,
		\P1_lWord_reg[13]/NET0131 ,
		_w1935_,
		_w9972_,
		_w15212_
	);
	LUT2 #(
		.INIT('hb)
	) name13863 (
		_w15211_,
		_w15212_,
		_w15213_
	);
	LUT2 #(
		.INIT('he)
	) name13864 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w15214_
	);
	LUT3 #(
		.INIT('he0)
	) name13865 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15215_
	);
	LUT4 #(
		.INIT('he000)
	) name13866 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15216_
	);
	LUT3 #(
		.INIT('h80)
	) name13867 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w15216_,
		_w15217_
	);
	LUT4 #(
		.INIT('h8000)
	) name13868 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w15216_,
		_w15218_
	);
	LUT3 #(
		.INIT('h80)
	) name13869 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w15218_,
		_w15219_
	);
	LUT4 #(
		.INIT('h8000)
	) name13870 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w15218_,
		_w15220_
	);
	LUT3 #(
		.INIT('h80)
	) name13871 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w15220_,
		_w15221_
	);
	LUT4 #(
		.INIT('h8000)
	) name13872 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w15220_,
		_w15222_
	);
	LUT3 #(
		.INIT('h80)
	) name13873 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w15222_,
		_w15223_
	);
	LUT4 #(
		.INIT('h8000)
	) name13874 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w15222_,
		_w15224_
	);
	LUT3 #(
		.INIT('h80)
	) name13875 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w15224_,
		_w15225_
	);
	LUT4 #(
		.INIT('h8000)
	) name13876 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w12026_,
		_w15224_,
		_w15226_
	);
	LUT3 #(
		.INIT('h80)
	) name13877 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w15226_,
		_w15227_
	);
	LUT4 #(
		.INIT('h8000)
	) name13878 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w15226_,
		_w15228_
	);
	LUT3 #(
		.INIT('h80)
	) name13879 (
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w15228_,
		_w15229_
	);
	LUT4 #(
		.INIT('h8000)
	) name13880 (
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w12192_,
		_w15228_,
		_w15230_
	);
	LUT3 #(
		.INIT('h80)
	) name13881 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w15230_,
		_w15231_
	);
	LUT4 #(
		.INIT('h60c0)
	) name13882 (
		\P3_rEIP_reg[29]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w2110_,
		_w15230_,
		_w15232_
	);
	LUT3 #(
		.INIT('h8a)
	) name13883 (
		\P3_Address_reg[28]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15233_
	);
	LUT2 #(
		.INIT('h8)
	) name13884 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15234_
	);
	LUT4 #(
		.INIT('h8000)
	) name13885 (
		_w11923_,
		_w12026_,
		_w12069_,
		_w15234_,
		_w15235_
	);
	LUT4 #(
		.INIT('h1555)
	) name13886 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w12119_,
		_w12192_,
		_w15235_,
		_w15236_
	);
	LUT3 #(
		.INIT('h40)
	) name13887 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w15237_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13888 (
		_w12120_,
		_w12193_,
		_w15234_,
		_w15237_,
		_w15238_
	);
	LUT3 #(
		.INIT('h45)
	) name13889 (
		_w15233_,
		_w15236_,
		_w15238_,
		_w15239_
	);
	LUT2 #(
		.INIT('hb)
	) name13890 (
		_w15232_,
		_w15239_,
		_w15240_
	);
	LUT2 #(
		.INIT('he)
	) name13891 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w15241_
	);
	LUT3 #(
		.INIT('he0)
	) name13892 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15242_
	);
	LUT4 #(
		.INIT('he000)
	) name13893 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15243_
	);
	LUT3 #(
		.INIT('h80)
	) name13894 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15243_,
		_w15244_
	);
	LUT4 #(
		.INIT('h8000)
	) name13895 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w9769_,
		_w15243_,
		_w15245_
	);
	LUT3 #(
		.INIT('h80)
	) name13896 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15245_,
		_w15246_
	);
	LUT4 #(
		.INIT('h8000)
	) name13897 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15245_,
		_w15247_
	);
	LUT3 #(
		.INIT('h80)
	) name13898 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w15247_,
		_w15248_
	);
	LUT4 #(
		.INIT('h8000)
	) name13899 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9777_,
		_w15247_,
		_w15249_
	);
	LUT3 #(
		.INIT('h80)
	) name13900 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w15249_,
		_w15250_
	);
	LUT4 #(
		.INIT('h8000)
	) name13901 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w15249_,
		_w15251_
	);
	LUT3 #(
		.INIT('h80)
	) name13902 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w15251_,
		_w15252_
	);
	LUT4 #(
		.INIT('h8000)
	) name13903 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w15251_,
		_w15253_
	);
	LUT3 #(
		.INIT('h80)
	) name13904 (
		\P2_rEIP_reg[25]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w15253_,
		_w15254_
	);
	LUT4 #(
		.INIT('h8000)
	) name13905 (
		\P2_rEIP_reg[25]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w15253_,
		_w15255_
	);
	LUT3 #(
		.INIT('h80)
	) name13906 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w15255_,
		_w15256_
	);
	LUT4 #(
		.INIT('h8000)
	) name13907 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w15255_,
		_w15257_
	);
	LUT3 #(
		.INIT('h8a)
	) name13908 (
		\P2_Address_reg[28]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15258_
	);
	LUT2 #(
		.INIT('h8)
	) name13909 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15259_
	);
	LUT3 #(
		.INIT('h80)
	) name13910 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9782_,
		_w15259_,
		_w15260_
	);
	LUT4 #(
		.INIT('h8000)
	) name13911 (
		\P2_rEIP_reg[26]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w9782_,
		_w15259_,
		_w15261_
	);
	LUT3 #(
		.INIT('h40)
	) name13912 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w15262_
	);
	LUT4 #(
		.INIT('h60c0)
	) name13913 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w15262_,
		_w15261_,
		_w15263_
	);
	LUT2 #(
		.INIT('h1)
	) name13914 (
		_w15258_,
		_w15263_,
		_w15264_
	);
	LUT4 #(
		.INIT('h48ff)
	) name13915 (
		\P2_rEIP_reg[30]/NET0131 ,
		_w1609_,
		_w15256_,
		_w15264_,
		_w15265_
	);
	LUT2 #(
		.INIT('he)
	) name13916 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w15266_
	);
	LUT3 #(
		.INIT('he0)
	) name13917 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15267_
	);
	LUT4 #(
		.INIT('he000)
	) name13918 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15268_
	);
	LUT3 #(
		.INIT('h80)
	) name13919 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15268_,
		_w15269_
	);
	LUT4 #(
		.INIT('h8000)
	) name13920 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w15268_,
		_w15270_
	);
	LUT3 #(
		.INIT('h80)
	) name13921 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w15270_,
		_w15271_
	);
	LUT4 #(
		.INIT('h8000)
	) name13922 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15270_,
		_w15272_
	);
	LUT3 #(
		.INIT('h80)
	) name13923 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w15272_,
		_w15273_
	);
	LUT4 #(
		.INIT('h8000)
	) name13924 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w15272_,
		_w15274_
	);
	LUT3 #(
		.INIT('h80)
	) name13925 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w15274_,
		_w15275_
	);
	LUT4 #(
		.INIT('h8000)
	) name13926 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w15274_,
		_w15276_
	);
	LUT3 #(
		.INIT('h80)
	) name13927 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w15276_,
		_w15277_
	);
	LUT4 #(
		.INIT('h8000)
	) name13928 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		_w15276_,
		_w15278_
	);
	LUT3 #(
		.INIT('h80)
	) name13929 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w11107_,
		_w15278_,
		_w15279_
	);
	LUT4 #(
		.INIT('h8000)
	) name13930 (
		\P1_rEIP_reg[26]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w11107_,
		_w15278_,
		_w15280_
	);
	LUT3 #(
		.INIT('h80)
	) name13931 (
		\P1_rEIP_reg[28]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w15280_,
		_w15281_
	);
	LUT4 #(
		.INIT('h8000)
	) name13932 (
		\P1_rEIP_reg[28]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w15280_,
		_w15282_
	);
	LUT3 #(
		.INIT('hb0)
	) name13933 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[28]_pad ,
		_w15283_
	);
	LUT2 #(
		.INIT('h8)
	) name13934 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15284_
	);
	LUT3 #(
		.INIT('h80)
	) name13935 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w11159_,
		_w15284_,
		_w15285_
	);
	LUT4 #(
		.INIT('h8000)
	) name13936 (
		\P1_rEIP_reg[27]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w11159_,
		_w15284_,
		_w15286_
	);
	LUT3 #(
		.INIT('h40)
	) name13937 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w15287_
	);
	LUT4 #(
		.INIT('h2133)
	) name13938 (
		\P1_rEIP_reg[29]/NET0131 ,
		_w15283_,
		_w15286_,
		_w15287_,
		_w15288_
	);
	LUT4 #(
		.INIT('h48ff)
	) name13939 (
		\P1_rEIP_reg[30]/NET0131 ,
		_w1856_,
		_w15281_,
		_w15288_,
		_w15289_
	);
	LUT4 #(
		.INIT('h1050)
	) name13940 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2230_,
		_w2232_,
		_w15290_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name13941 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w15291_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name13942 (
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3544_,
		_w15290_,
		_w15291_,
		_w15292_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13943 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3407_,
		_w3535_,
		_w15293_
	);
	LUT3 #(
		.INIT('h54)
	) name13944 (
		_w2248_,
		_w4953_,
		_w15293_,
		_w15294_
	);
	LUT2 #(
		.INIT('h2)
	) name13945 (
		_w3535_,
		_w4953_,
		_w15295_
	);
	LUT3 #(
		.INIT('h07)
	) name13946 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15296_
	);
	LUT3 #(
		.INIT('h70)
	) name13947 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w15296_,
		_w15297_
	);
	LUT3 #(
		.INIT('h45)
	) name13948 (
		_w3579_,
		_w15295_,
		_w15297_,
		_w15298_
	);
	LUT3 #(
		.INIT('hba)
	) name13949 (
		_w15292_,
		_w15294_,
		_w15298_,
		_w15299_
	);
	LUT4 #(
		.INIT('h1050)
	) name13950 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2216_,
		_w2221_,
		_w15300_
	);
	LUT4 #(
		.INIT('hfd94)
	) name13951 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w15301_
	);
	LUT3 #(
		.INIT('h8a)
	) name13952 (
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15300_,
		_w15301_,
		_w15302_
	);
	LUT4 #(
		.INIT('hcc08)
	) name13953 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3055_,
		_w10615_,
		_w15303_
	);
	LUT3 #(
		.INIT('h54)
	) name13954 (
		_w2215_,
		_w6349_,
		_w15303_,
		_w15304_
	);
	LUT3 #(
		.INIT('h8c)
	) name13955 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w6349_,
		_w15305_
	);
	LUT3 #(
		.INIT('h13)
	) name13956 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2194_,
		_w15306_
	);
	LUT3 #(
		.INIT('h45)
	) name13957 (
		_w10619_,
		_w15305_,
		_w15306_,
		_w15307_
	);
	LUT3 #(
		.INIT('hba)
	) name13958 (
		_w15302_,
		_w15304_,
		_w15307_,
		_w15308_
	);
	LUT3 #(
		.INIT('hc8)
	) name13959 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		_w2215_,
		_w10611_,
		_w15309_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13960 (
		_w1999_,
		_w2004_,
		_w10611_,
		_w15309_,
		_w15310_
	);
	LUT4 #(
		.INIT('h20aa)
	) name13961 (
		\P3_InstQueue_reg[0][5]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w15311_
	);
	LUT4 #(
		.INIT('h153f)
	) name13962 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10614_,
		_w10616_,
		_w15312_
	);
	LUT2 #(
		.INIT('h2)
	) name13963 (
		_w2199_,
		_w15312_,
		_w15313_
	);
	LUT3 #(
		.INIT('h02)
	) name13964 (
		\buf2_reg[5]/NET0131 ,
		_w10618_,
		_w10621_,
		_w15314_
	);
	LUT3 #(
		.INIT('h01)
	) name13965 (
		_w15311_,
		_w15313_,
		_w15314_,
		_w15315_
	);
	LUT2 #(
		.INIT('hb)
	) name13966 (
		_w15310_,
		_w15315_,
		_w15316_
	);
	LUT3 #(
		.INIT('hc8)
	) name13967 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		_w2215_,
		_w10630_,
		_w15317_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13968 (
		_w1999_,
		_w2004_,
		_w10630_,
		_w15317_,
		_w15318_
	);
	LUT4 #(
		.INIT('h222a)
	) name13969 (
		\P3_InstQueue_reg[10][5]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w15319_
	);
	LUT4 #(
		.INIT('h153f)
	) name13970 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10633_,
		_w10635_,
		_w15320_
	);
	LUT2 #(
		.INIT('h2)
	) name13971 (
		_w2199_,
		_w15320_,
		_w15321_
	);
	LUT3 #(
		.INIT('h20)
	) name13972 (
		\buf2_reg[5]/NET0131 ,
		_w10637_,
		_w10639_,
		_w15322_
	);
	LUT3 #(
		.INIT('h01)
	) name13973 (
		_w15319_,
		_w15321_,
		_w15322_,
		_w15323_
	);
	LUT2 #(
		.INIT('hb)
	) name13974 (
		_w15318_,
		_w15323_,
		_w15324_
	);
	LUT3 #(
		.INIT('hc8)
	) name13975 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w2215_,
		_w10646_,
		_w15325_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13976 (
		_w1999_,
		_w2004_,
		_w10646_,
		_w15325_,
		_w15326_
	);
	LUT3 #(
		.INIT('ha2)
	) name13977 (
		\P3_InstQueue_reg[11][5]/NET0131 ,
		_w10622_,
		_w10650_,
		_w15327_
	);
	LUT3 #(
		.INIT('hd8)
	) name13978 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w15328_
	);
	LUT3 #(
		.INIT('h80)
	) name13979 (
		_w2194_,
		_w10649_,
		_w15328_,
		_w15329_
	);
	LUT4 #(
		.INIT('h2000)
	) name13980 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w15330_
	);
	LUT4 #(
		.INIT('hce00)
	) name13981 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w15330_,
		_w15331_
	);
	LUT2 #(
		.INIT('h1)
	) name13982 (
		_w15329_,
		_w15331_,
		_w15332_
	);
	LUT2 #(
		.INIT('h4)
	) name13983 (
		_w15327_,
		_w15332_,
		_w15333_
	);
	LUT2 #(
		.INIT('hb)
	) name13984 (
		_w15326_,
		_w15333_,
		_w15334_
	);
	LUT3 #(
		.INIT('hc8)
	) name13985 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w2215_,
		_w10659_,
		_w15335_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13986 (
		_w1999_,
		_w2004_,
		_w10659_,
		_w15335_,
		_w15336_
	);
	LUT4 #(
		.INIT('h2a22)
	) name13987 (
		\P3_InstQueue_reg[12][5]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w15337_
	);
	LUT4 #(
		.INIT('h135f)
	) name13988 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10630_,
		_w10652_,
		_w15338_
	);
	LUT2 #(
		.INIT('h2)
	) name13989 (
		_w2199_,
		_w15338_,
		_w15339_
	);
	LUT3 #(
		.INIT('h02)
	) name13990 (
		\buf2_reg[5]/NET0131 ,
		_w10662_,
		_w10663_,
		_w15340_
	);
	LUT3 #(
		.INIT('h01)
	) name13991 (
		_w15337_,
		_w15339_,
		_w15340_,
		_w15341_
	);
	LUT2 #(
		.INIT('hb)
	) name13992 (
		_w15336_,
		_w15341_,
		_w15342_
	);
	LUT3 #(
		.INIT('hc8)
	) name13993 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w2215_,
		_w10614_,
		_w15343_
	);
	LUT4 #(
		.INIT('h7f00)
	) name13994 (
		_w1999_,
		_w2004_,
		_w10614_,
		_w15343_,
		_w15344_
	);
	LUT2 #(
		.INIT('h4)
	) name13995 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w10672_,
		_w15345_
	);
	LUT2 #(
		.INIT('h1)
	) name13996 (
		\buf2_reg[5]/NET0131 ,
		_w10672_,
		_w15346_
	);
	LUT3 #(
		.INIT('h02)
	) name13997 (
		_w10674_,
		_w15346_,
		_w15345_,
		_w15347_
	);
	LUT2 #(
		.INIT('h2)
	) name13998 (
		\P3_InstQueue_reg[13][5]/NET0131 ,
		_w10622_,
		_w15348_
	);
	LUT3 #(
		.INIT('h80)
	) name13999 (
		_w2194_,
		_w10673_,
		_w15328_,
		_w15349_
	);
	LUT2 #(
		.INIT('h1)
	) name14000 (
		_w15348_,
		_w15349_,
		_w15350_
	);
	LUT2 #(
		.INIT('h4)
	) name14001 (
		_w15347_,
		_w15350_,
		_w15351_
	);
	LUT2 #(
		.INIT('hb)
	) name14002 (
		_w15344_,
		_w15351_,
		_w15352_
	);
	LUT3 #(
		.INIT('hc8)
	) name14003 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w2215_,
		_w10616_,
		_w15353_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14004 (
		_w1999_,
		_w2004_,
		_w10616_,
		_w15353_,
		_w15354_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name14005 (
		\P3_InstQueue_reg[14][5]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w15355_
	);
	LUT4 #(
		.INIT('h153f)
	) name14006 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10646_,
		_w10659_,
		_w15356_
	);
	LUT2 #(
		.INIT('h2)
	) name14007 (
		_w2199_,
		_w15356_,
		_w15357_
	);
	LUT3 #(
		.INIT('h02)
	) name14008 (
		\buf2_reg[5]/NET0131 ,
		_w10617_,
		_w10684_,
		_w15358_
	);
	LUT3 #(
		.INIT('h01)
	) name14009 (
		_w15355_,
		_w15357_,
		_w15358_,
		_w15359_
	);
	LUT2 #(
		.INIT('hb)
	) name14010 (
		_w15354_,
		_w15359_,
		_w15360_
	);
	LUT3 #(
		.INIT('hc8)
	) name14011 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w2215_,
		_w10620_,
		_w15361_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14012 (
		_w1999_,
		_w2004_,
		_w10620_,
		_w15361_,
		_w15362_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14013 (
		\P3_InstQueue_reg[15][5]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w15363_
	);
	LUT4 #(
		.INIT('h135f)
	) name14014 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10614_,
		_w10659_,
		_w15364_
	);
	LUT2 #(
		.INIT('h2)
	) name14015 (
		_w2199_,
		_w15364_,
		_w15365_
	);
	LUT3 #(
		.INIT('h02)
	) name14016 (
		\buf2_reg[5]/NET0131 ,
		_w10693_,
		_w10694_,
		_w15366_
	);
	LUT3 #(
		.INIT('h01)
	) name14017 (
		_w15363_,
		_w15365_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('hb)
	) name14018 (
		_w15362_,
		_w15367_,
		_w15368_
	);
	LUT3 #(
		.INIT('hc8)
	) name14019 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w2215_,
		_w10701_,
		_w15369_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14020 (
		_w1999_,
		_w2004_,
		_w10701_,
		_w15369_,
		_w15370_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14021 (
		\P3_InstQueue_reg[1][5]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w15371_
	);
	LUT4 #(
		.INIT('h153f)
	) name14022 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10616_,
		_w10620_,
		_w15372_
	);
	LUT2 #(
		.INIT('h2)
	) name14023 (
		_w2199_,
		_w15372_,
		_w15373_
	);
	LUT3 #(
		.INIT('h02)
	) name14024 (
		\buf2_reg[5]/NET0131 ,
		_w10704_,
		_w10705_,
		_w15374_
	);
	LUT3 #(
		.INIT('h01)
	) name14025 (
		_w15371_,
		_w15373_,
		_w15374_,
		_w15375_
	);
	LUT2 #(
		.INIT('hb)
	) name14026 (
		_w15370_,
		_w15375_,
		_w15376_
	);
	LUT3 #(
		.INIT('hc8)
	) name14027 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w2215_,
		_w10713_,
		_w15377_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14028 (
		_w1999_,
		_w2004_,
		_w10713_,
		_w15377_,
		_w15378_
	);
	LUT4 #(
		.INIT('h222a)
	) name14029 (
		\P3_InstQueue_reg[2][5]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w15379_
	);
	LUT4 #(
		.INIT('h135f)
	) name14030 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10611_,
		_w10620_,
		_w15380_
	);
	LUT2 #(
		.INIT('h2)
	) name14031 (
		_w2199_,
		_w15380_,
		_w15381_
	);
	LUT3 #(
		.INIT('h20)
	) name14032 (
		\buf2_reg[5]/NET0131 ,
		_w10716_,
		_w10717_,
		_w15382_
	);
	LUT3 #(
		.INIT('h01)
	) name14033 (
		_w15379_,
		_w15381_,
		_w15382_,
		_w15383_
	);
	LUT2 #(
		.INIT('hb)
	) name14034 (
		_w15378_,
		_w15383_,
		_w15384_
	);
	LUT3 #(
		.INIT('hc8)
	) name14035 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w2215_,
		_w10724_,
		_w15385_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14036 (
		_w1999_,
		_w2004_,
		_w10724_,
		_w15385_,
		_w15386_
	);
	LUT4 #(
		.INIT('h222a)
	) name14037 (
		\P3_InstQueue_reg[3][5]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w15387_
	);
	LUT4 #(
		.INIT('h153f)
	) name14038 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10611_,
		_w10701_,
		_w15388_
	);
	LUT2 #(
		.INIT('h2)
	) name14039 (
		_w2199_,
		_w15388_,
		_w15389_
	);
	LUT3 #(
		.INIT('h08)
	) name14040 (
		\buf2_reg[5]/NET0131 ,
		_w10712_,
		_w10727_,
		_w15390_
	);
	LUT3 #(
		.INIT('h01)
	) name14041 (
		_w15387_,
		_w15389_,
		_w15390_,
		_w15391_
	);
	LUT2 #(
		.INIT('hb)
	) name14042 (
		_w15386_,
		_w15391_,
		_w15392_
	);
	LUT3 #(
		.INIT('hc8)
	) name14043 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w2215_,
		_w10734_,
		_w15393_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14044 (
		_w1999_,
		_w2004_,
		_w10734_,
		_w15393_,
		_w15394_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14045 (
		\P3_InstQueue_reg[4][5]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w15395_
	);
	LUT4 #(
		.INIT('h153f)
	) name14046 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10701_,
		_w10713_,
		_w15396_
	);
	LUT2 #(
		.INIT('h2)
	) name14047 (
		_w2199_,
		_w15396_,
		_w15397_
	);
	LUT3 #(
		.INIT('h02)
	) name14048 (
		\buf2_reg[5]/NET0131 ,
		_w10737_,
		_w10738_,
		_w15398_
	);
	LUT3 #(
		.INIT('h01)
	) name14049 (
		_w15395_,
		_w15397_,
		_w15398_,
		_w15399_
	);
	LUT2 #(
		.INIT('hb)
	) name14050 (
		_w15394_,
		_w15399_,
		_w15400_
	);
	LUT3 #(
		.INIT('hc8)
	) name14051 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w2215_,
		_w10745_,
		_w15401_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14052 (
		_w1999_,
		_w2004_,
		_w10745_,
		_w15401_,
		_w15402_
	);
	LUT2 #(
		.INIT('h4)
	) name14053 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w10748_,
		_w15403_
	);
	LUT2 #(
		.INIT('h1)
	) name14054 (
		\buf2_reg[5]/NET0131 ,
		_w10748_,
		_w15404_
	);
	LUT3 #(
		.INIT('h02)
	) name14055 (
		_w10750_,
		_w15404_,
		_w15403_,
		_w15405_
	);
	LUT2 #(
		.INIT('h2)
	) name14056 (
		\P3_InstQueue_reg[5][5]/NET0131 ,
		_w10622_,
		_w15406_
	);
	LUT3 #(
		.INIT('h80)
	) name14057 (
		_w2194_,
		_w10749_,
		_w15328_,
		_w15407_
	);
	LUT2 #(
		.INIT('h1)
	) name14058 (
		_w15406_,
		_w15407_,
		_w15408_
	);
	LUT2 #(
		.INIT('h4)
	) name14059 (
		_w15405_,
		_w15408_,
		_w15409_
	);
	LUT2 #(
		.INIT('hb)
	) name14060 (
		_w15402_,
		_w15409_,
		_w15410_
	);
	LUT3 #(
		.INIT('hc8)
	) name14061 (
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w2215_,
		_w10758_,
		_w15411_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14062 (
		_w1999_,
		_w2004_,
		_w10758_,
		_w15411_,
		_w15412_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14063 (
		\P3_InstQueue_reg[6][5]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w15413_
	);
	LUT4 #(
		.INIT('h153f)
	) name14064 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10724_,
		_w10734_,
		_w15414_
	);
	LUT2 #(
		.INIT('h2)
	) name14065 (
		_w2199_,
		_w15414_,
		_w15415_
	);
	LUT3 #(
		.INIT('h02)
	) name14066 (
		\buf2_reg[5]/NET0131 ,
		_w10761_,
		_w10762_,
		_w15416_
	);
	LUT3 #(
		.INIT('h01)
	) name14067 (
		_w15413_,
		_w15415_,
		_w15416_,
		_w15417_
	);
	LUT2 #(
		.INIT('hb)
	) name14068 (
		_w15412_,
		_w15417_,
		_w15418_
	);
	LUT3 #(
		.INIT('hc8)
	) name14069 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w2215_,
		_w10633_,
		_w15419_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14070 (
		_w1999_,
		_w2004_,
		_w10633_,
		_w15419_,
		_w15420_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14071 (
		\P3_InstQueue_reg[7][5]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w15421_
	);
	LUT4 #(
		.INIT('h153f)
	) name14072 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10734_,
		_w10745_,
		_w15422_
	);
	LUT2 #(
		.INIT('h2)
	) name14073 (
		_w2199_,
		_w15422_,
		_w15423_
	);
	LUT3 #(
		.INIT('h02)
	) name14074 (
		\buf2_reg[5]/NET0131 ,
		_w10771_,
		_w10772_,
		_w15424_
	);
	LUT3 #(
		.INIT('h01)
	) name14075 (
		_w15421_,
		_w15423_,
		_w15424_,
		_w15425_
	);
	LUT2 #(
		.INIT('hb)
	) name14076 (
		_w15420_,
		_w15425_,
		_w15426_
	);
	LUT3 #(
		.INIT('hc8)
	) name14077 (
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w2215_,
		_w10635_,
		_w15427_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14078 (
		_w1999_,
		_w2004_,
		_w10635_,
		_w15427_,
		_w15428_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14079 (
		\P3_InstQueue_reg[8][5]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w15429_
	);
	LUT4 #(
		.INIT('h153f)
	) name14080 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10745_,
		_w10758_,
		_w15430_
	);
	LUT2 #(
		.INIT('h2)
	) name14081 (
		_w2199_,
		_w15430_,
		_w15431_
	);
	LUT3 #(
		.INIT('h02)
	) name14082 (
		\buf2_reg[5]/NET0131 ,
		_w10636_,
		_w10781_,
		_w15432_
	);
	LUT3 #(
		.INIT('h01)
	) name14083 (
		_w15429_,
		_w15431_,
		_w15432_,
		_w15433_
	);
	LUT2 #(
		.INIT('hb)
	) name14084 (
		_w15428_,
		_w15433_,
		_w15434_
	);
	LUT3 #(
		.INIT('hc8)
	) name14085 (
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w2215_,
		_w10652_,
		_w15435_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14086 (
		_w1999_,
		_w2004_,
		_w10652_,
		_w15435_,
		_w15436_
	);
	LUT4 #(
		.INIT('h135f)
	) name14087 (
		\buf2_reg[21]/NET0131 ,
		\buf2_reg[29]/NET0131 ,
		_w10633_,
		_w10758_,
		_w15437_
	);
	LUT4 #(
		.INIT('hef00)
	) name14088 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w15438_
	);
	LUT4 #(
		.INIT('h1000)
	) name14089 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[5]/NET0131 ,
		_w15439_
	);
	LUT4 #(
		.INIT('hddd0)
	) name14090 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w15438_,
		_w15439_,
		_w15440_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14091 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w15437_,
		_w15440_,
		_w15441_
	);
	LUT3 #(
		.INIT('ha8)
	) name14092 (
		_w3055_,
		_w15438_,
		_w15439_,
		_w15442_
	);
	LUT2 #(
		.INIT('h2)
	) name14093 (
		\P3_InstQueue_reg[9][5]/NET0131 ,
		_w10622_,
		_w15443_
	);
	LUT2 #(
		.INIT('h1)
	) name14094 (
		_w15442_,
		_w15443_,
		_w15444_
	);
	LUT2 #(
		.INIT('h4)
	) name14095 (
		_w15441_,
		_w15444_,
		_w15445_
	);
	LUT2 #(
		.INIT('hb)
	) name14096 (
		_w15436_,
		_w15445_,
		_w15446_
	);
	LUT4 #(
		.INIT('h1050)
	) name14097 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueRd_Addr_reg[2]/NET0131 ,
		_w2205_,
		_w2207_,
		_w15447_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name14098 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w15448_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14099 (
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w12455_,
		_w15447_,
		_w15448_,
		_w15449_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name14100 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2270_,
		_w2283_,
		_w15450_
	);
	LUT3 #(
		.INIT('h54)
	) name14101 (
		_w2246_,
		_w2298_,
		_w15450_,
		_w15451_
	);
	LUT2 #(
		.INIT('h2)
	) name14102 (
		_w2270_,
		_w2298_,
		_w15452_
	);
	LUT3 #(
		.INIT('h07)
	) name14103 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		_w15453_
	);
	LUT3 #(
		.INIT('h70)
	) name14104 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w15453_,
		_w15454_
	);
	LUT3 #(
		.INIT('h45)
	) name14105 (
		_w2321_,
		_w15452_,
		_w15454_,
		_w15455_
	);
	LUT3 #(
		.INIT('hba)
	) name14106 (
		_w15449_,
		_w15451_,
		_w15455_,
		_w15456_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14107 (
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w2110_,
		_w15225_,
		_w15457_
	);
	LUT3 #(
		.INIT('h8a)
	) name14108 (
		\P3_Address_reg[16]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15458_
	);
	LUT3 #(
		.INIT('h80)
	) name14109 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w11871_,
		_w15234_,
		_w15459_
	);
	LUT4 #(
		.INIT('h8000)
	) name14110 (
		\P3_rEIP_reg[14]/NET0131 ,
		\P3_rEIP_reg[15]/NET0131 ,
		_w11871_,
		_w15234_,
		_w15460_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14111 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w15237_,
		_w15460_,
		_w15461_
	);
	LUT2 #(
		.INIT('h1)
	) name14112 (
		_w15458_,
		_w15461_,
		_w15462_
	);
	LUT2 #(
		.INIT('hb)
	) name14113 (
		_w15457_,
		_w15462_,
		_w15463_
	);
	LUT4 #(
		.INIT('h4888)
	) name14114 (
		\P2_rEIP_reg[18]/NET0131 ,
		_w1609_,
		_w9776_,
		_w15248_,
		_w15464_
	);
	LUT3 #(
		.INIT('h8a)
	) name14115 (
		\P2_Address_reg[16]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15465_
	);
	LUT3 #(
		.INIT('h13)
	) name14116 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15466_
	);
	LUT2 #(
		.INIT('h2)
	) name14117 (
		_w15262_,
		_w15466_,
		_w15467_
	);
	LUT4 #(
		.INIT('h040f)
	) name14118 (
		_w11261_,
		_w15259_,
		_w15465_,
		_w15467_,
		_w15468_
	);
	LUT2 #(
		.INIT('hb)
	) name14119 (
		_w15464_,
		_w15468_,
		_w15469_
	);
	LUT3 #(
		.INIT('h48)
	) name14120 (
		\P1_rEIP_reg[18]/NET0131 ,
		_w1856_,
		_w15278_,
		_w15470_
	);
	LUT3 #(
		.INIT('hb0)
	) name14121 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[16]_pad ,
		_w15471_
	);
	LUT3 #(
		.INIT('h13)
	) name14122 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15472_
	);
	LUT2 #(
		.INIT('h2)
	) name14123 (
		_w15287_,
		_w15472_,
		_w15473_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14124 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w10858_,
		_w15284_,
		_w15473_,
		_w15474_
	);
	LUT2 #(
		.INIT('h1)
	) name14125 (
		_w15471_,
		_w15474_,
		_w15475_
	);
	LUT2 #(
		.INIT('hb)
	) name14126 (
		_w15470_,
		_w15475_,
		_w15476_
	);
	LUT4 #(
		.INIT('h7f80)
	) name14127 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15477_
	);
	LUT4 #(
		.INIT('hc03f)
	) name14128 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15478_
	);
	LUT4 #(
		.INIT('he00f)
	) name14129 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15479_
	);
	LUT4 #(
		.INIT('h0008)
	) name14130 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3611_,
		_w15479_,
		_w15480_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14131 (
		\P1_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3544_,
		_w15290_,
		_w15291_,
		_w15481_
	);
	LUT2 #(
		.INIT('h8)
	) name14132 (
		_w2248_,
		_w15477_,
		_w15482_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14133 (
		\P1_DataWidth_reg[1]/NET0131 ,
		_w1939_,
		_w3407_,
		_w15478_,
		_w15483_
	);
	LUT2 #(
		.INIT('h1)
	) name14134 (
		_w15482_,
		_w15483_,
		_w15484_
	);
	LUT3 #(
		.INIT('hef)
	) name14135 (
		_w15480_,
		_w15481_,
		_w15484_,
		_w15485_
	);
	LUT4 #(
		.INIT('h7f80)
	) name14136 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15486_
	);
	LUT4 #(
		.INIT('hc03f)
	) name14137 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15487_
	);
	LUT4 #(
		.INIT('he00f)
	) name14138 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15488_
	);
	LUT4 #(
		.INIT('h0008)
	) name14139 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w10659_,
		_w15488_,
		_w15489_
	);
	LUT3 #(
		.INIT('h8a)
	) name14140 (
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15300_,
		_w15301_,
		_w15490_
	);
	LUT2 #(
		.INIT('h8)
	) name14141 (
		_w2215_,
		_w15486_,
		_w15491_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14142 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w15487_,
		_w15492_
	);
	LUT2 #(
		.INIT('h1)
	) name14143 (
		_w15491_,
		_w15492_,
		_w15493_
	);
	LUT3 #(
		.INIT('hef)
	) name14144 (
		_w15489_,
		_w15490_,
		_w15493_,
		_w15494_
	);
	LUT4 #(
		.INIT('h807f)
	) name14145 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15495_
	);
	LUT4 #(
		.INIT('hc03f)
	) name14146 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15496_
	);
	LUT4 #(
		.INIT('he00f)
	) name14147 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w15497_
	);
	LUT4 #(
		.INIT('h0008)
	) name14148 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2376_,
		_w15497_,
		_w15498_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name14149 (
		\P2_InstQueueWr_Addr_reg[3]/NET0131 ,
		_w12455_,
		_w15447_,
		_w15448_,
		_w15499_
	);
	LUT2 #(
		.INIT('h2)
	) name14150 (
		_w2246_,
		_w15495_,
		_w15500_
	);
	LUT4 #(
		.INIT('h00f4)
	) name14151 (
		\P2_DataWidth_reg[1]/NET0131 ,
		_w1679_,
		_w2283_,
		_w15496_,
		_w15501_
	);
	LUT2 #(
		.INIT('h1)
	) name14152 (
		_w15500_,
		_w15501_,
		_w15502_
	);
	LUT3 #(
		.INIT('hef)
	) name14153 (
		_w15498_,
		_w15499_,
		_w15502_,
		_w15503_
	);
	LUT3 #(
		.INIT('h8a)
	) name14154 (
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w15290_,
		_w15291_,
		_w15504_
	);
	LUT2 #(
		.INIT('h4)
	) name14155 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2248_,
		_w15505_
	);
	LUT4 #(
		.INIT('h4c00)
	) name14156 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1939_,
		_w3544_,
		_w15506_
	);
	LUT3 #(
		.INIT('h13)
	) name14157 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P1_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2248_,
		_w15507_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14158 (
		_w6378_,
		_w15505_,
		_w15506_,
		_w15507_,
		_w15508_
	);
	LUT2 #(
		.INIT('he)
	) name14159 (
		_w15504_,
		_w15508_,
		_w15509_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name14160 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2199_,
		_w15300_,
		_w15301_,
		_w15510_
	);
	LUT4 #(
		.INIT('h3310)
	) name14161 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2194_,
		_w3055_,
		_w15511_
	);
	LUT2 #(
		.INIT('h2)
	) name14162 (
		_w2215_,
		_w10638_,
		_w15512_
	);
	LUT2 #(
		.INIT('h1)
	) name14163 (
		_w15511_,
		_w15512_,
		_w15513_
	);
	LUT2 #(
		.INIT('hb)
	) name14164 (
		_w15510_,
		_w15513_,
		_w15514_
	);
	LUT3 #(
		.INIT('h8a)
	) name14165 (
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w15447_,
		_w15448_,
		_w15515_
	);
	LUT2 #(
		.INIT('h4)
	) name14166 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2246_,
		_w15516_
	);
	LUT4 #(
		.INIT('h4c00)
	) name14167 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w1679_,
		_w12455_,
		_w15517_
	);
	LUT3 #(
		.INIT('h13)
	) name14168 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		\P2_InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2246_,
		_w15518_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14169 (
		_w5746_,
		_w15516_,
		_w15517_,
		_w15518_,
		_w15519_
	);
	LUT2 #(
		.INIT('he)
	) name14170 (
		_w15515_,
		_w15519_,
		_w15520_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14171 (
		\P1_State2_reg[0]/NET0131 ,
		\P1_State2_reg[1]/NET0131 ,
		\P1_State2_reg[2]/NET0131 ,
		\P1_State2_reg[3]/NET0131 ,
		_w15521_
	);
	LUT2 #(
		.INIT('h2)
	) name14172 (
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15521_,
		_w15522_
	);
	LUT2 #(
		.INIT('h1)
	) name14173 (
		\P1_Flush_reg/NET0131 ,
		\P1_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15523_
	);
	LUT4 #(
		.INIT('h002a)
	) name14174 (
		_w2230_,
		_w2231_,
		_w2232_,
		_w15523_,
		_w15524_
	);
	LUT3 #(
		.INIT('hfe)
	) name14175 (
		_w15505_,
		_w15524_,
		_w15522_,
		_w15525_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14176 (
		\P3_State2_reg[0]/NET0131 ,
		\P3_State2_reg[1]/NET0131 ,
		\P3_State2_reg[2]/NET0131 ,
		\P3_State2_reg[3]/NET0131 ,
		_w15526_
	);
	LUT2 #(
		.INIT('h2)
	) name14177 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15526_,
		_w15527_
	);
	LUT2 #(
		.INIT('h4)
	) name14178 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w2215_,
		_w15528_
	);
	LUT2 #(
		.INIT('h1)
	) name14179 (
		\P3_Flush_reg/NET0131 ,
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15529_
	);
	LUT4 #(
		.INIT('h002a)
	) name14180 (
		_w2216_,
		_w2220_,
		_w2221_,
		_w15529_,
		_w15530_
	);
	LUT3 #(
		.INIT('hfe)
	) name14181 (
		_w15528_,
		_w15530_,
		_w15527_,
		_w15531_
	);
	LUT3 #(
		.INIT('hc8)
	) name14182 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		_w2215_,
		_w10611_,
		_w15532_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14183 (
		_w2054_,
		_w2059_,
		_w10611_,
		_w15532_,
		_w15533_
	);
	LUT4 #(
		.INIT('h20aa)
	) name14184 (
		\P3_InstQueue_reg[0][1]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w15534_
	);
	LUT4 #(
		.INIT('h153f)
	) name14185 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10614_,
		_w10616_,
		_w15535_
	);
	LUT2 #(
		.INIT('h2)
	) name14186 (
		_w2199_,
		_w15535_,
		_w15536_
	);
	LUT3 #(
		.INIT('h02)
	) name14187 (
		\buf2_reg[1]/NET0131 ,
		_w10618_,
		_w10621_,
		_w15537_
	);
	LUT3 #(
		.INIT('h01)
	) name14188 (
		_w15534_,
		_w15536_,
		_w15537_,
		_w15538_
	);
	LUT2 #(
		.INIT('hb)
	) name14189 (
		_w15533_,
		_w15538_,
		_w15539_
	);
	LUT3 #(
		.INIT('hc8)
	) name14190 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		_w2215_,
		_w10630_,
		_w15540_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14191 (
		_w2054_,
		_w2059_,
		_w10630_,
		_w15540_,
		_w15541_
	);
	LUT4 #(
		.INIT('h222a)
	) name14192 (
		\P3_InstQueue_reg[10][1]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w15542_
	);
	LUT4 #(
		.INIT('h153f)
	) name14193 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10633_,
		_w10635_,
		_w15543_
	);
	LUT2 #(
		.INIT('h2)
	) name14194 (
		_w2199_,
		_w15543_,
		_w15544_
	);
	LUT3 #(
		.INIT('h20)
	) name14195 (
		\buf2_reg[1]/NET0131 ,
		_w10637_,
		_w10639_,
		_w15545_
	);
	LUT3 #(
		.INIT('h01)
	) name14196 (
		_w15542_,
		_w15544_,
		_w15545_,
		_w15546_
	);
	LUT2 #(
		.INIT('hb)
	) name14197 (
		_w15541_,
		_w15546_,
		_w15547_
	);
	LUT3 #(
		.INIT('hc8)
	) name14198 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w2215_,
		_w10646_,
		_w15548_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14199 (
		_w2022_,
		_w2027_,
		_w10646_,
		_w15548_,
		_w15549_
	);
	LUT3 #(
		.INIT('ha2)
	) name14200 (
		\P3_InstQueue_reg[11][0]/NET0131 ,
		_w10622_,
		_w10650_,
		_w15550_
	);
	LUT3 #(
		.INIT('hd8)
	) name14201 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w15551_
	);
	LUT3 #(
		.INIT('h80)
	) name14202 (
		_w2194_,
		_w10649_,
		_w15551_,
		_w15552_
	);
	LUT4 #(
		.INIT('h2000)
	) name14203 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w15553_
	);
	LUT4 #(
		.INIT('hce00)
	) name14204 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w15553_,
		_w15554_
	);
	LUT2 #(
		.INIT('h1)
	) name14205 (
		_w15552_,
		_w15554_,
		_w15555_
	);
	LUT2 #(
		.INIT('h4)
	) name14206 (
		_w15550_,
		_w15555_,
		_w15556_
	);
	LUT2 #(
		.INIT('hb)
	) name14207 (
		_w15549_,
		_w15556_,
		_w15557_
	);
	LUT3 #(
		.INIT('hc8)
	) name14208 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w2215_,
		_w10646_,
		_w15558_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14209 (
		_w2054_,
		_w2059_,
		_w10646_,
		_w15558_,
		_w15559_
	);
	LUT3 #(
		.INIT('ha2)
	) name14210 (
		\P3_InstQueue_reg[11][1]/NET0131 ,
		_w10622_,
		_w10650_,
		_w15560_
	);
	LUT3 #(
		.INIT('hd8)
	) name14211 (
		\P3_InstQueueWr_Addr_reg[0]/NET0131 ,
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w15561_
	);
	LUT3 #(
		.INIT('h80)
	) name14212 (
		_w2194_,
		_w10649_,
		_w15561_,
		_w15562_
	);
	LUT4 #(
		.INIT('h2000)
	) name14213 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w15563_
	);
	LUT4 #(
		.INIT('hce00)
	) name14214 (
		_w2194_,
		_w3055_,
		_w10649_,
		_w15563_,
		_w15564_
	);
	LUT2 #(
		.INIT('h1)
	) name14215 (
		_w15562_,
		_w15564_,
		_w15565_
	);
	LUT2 #(
		.INIT('h4)
	) name14216 (
		_w15560_,
		_w15565_,
		_w15566_
	);
	LUT2 #(
		.INIT('hb)
	) name14217 (
		_w15559_,
		_w15566_,
		_w15567_
	);
	LUT3 #(
		.INIT('hc8)
	) name14218 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w2215_,
		_w10659_,
		_w15568_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14219 (
		_w2054_,
		_w2059_,
		_w10659_,
		_w15568_,
		_w15569_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14220 (
		\P3_InstQueue_reg[12][1]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w15570_
	);
	LUT4 #(
		.INIT('h135f)
	) name14221 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10630_,
		_w10652_,
		_w15571_
	);
	LUT2 #(
		.INIT('h2)
	) name14222 (
		_w2199_,
		_w15571_,
		_w15572_
	);
	LUT3 #(
		.INIT('h02)
	) name14223 (
		\buf2_reg[1]/NET0131 ,
		_w10662_,
		_w10663_,
		_w15573_
	);
	LUT3 #(
		.INIT('h01)
	) name14224 (
		_w15570_,
		_w15572_,
		_w15573_,
		_w15574_
	);
	LUT2 #(
		.INIT('hb)
	) name14225 (
		_w15569_,
		_w15574_,
		_w15575_
	);
	LUT3 #(
		.INIT('hc8)
	) name14226 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w2215_,
		_w10614_,
		_w15576_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14227 (
		_w2054_,
		_w2059_,
		_w10614_,
		_w15576_,
		_w15577_
	);
	LUT2 #(
		.INIT('h4)
	) name14228 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w10672_,
		_w15578_
	);
	LUT2 #(
		.INIT('h1)
	) name14229 (
		\buf2_reg[1]/NET0131 ,
		_w10672_,
		_w15579_
	);
	LUT3 #(
		.INIT('h02)
	) name14230 (
		_w10674_,
		_w15579_,
		_w15578_,
		_w15580_
	);
	LUT2 #(
		.INIT('h2)
	) name14231 (
		\P3_InstQueue_reg[13][1]/NET0131 ,
		_w10622_,
		_w15581_
	);
	LUT3 #(
		.INIT('h80)
	) name14232 (
		_w2194_,
		_w10673_,
		_w15561_,
		_w15582_
	);
	LUT2 #(
		.INIT('h1)
	) name14233 (
		_w15581_,
		_w15582_,
		_w15583_
	);
	LUT2 #(
		.INIT('h4)
	) name14234 (
		_w15580_,
		_w15583_,
		_w15584_
	);
	LUT2 #(
		.INIT('hb)
	) name14235 (
		_w15577_,
		_w15584_,
		_w15585_
	);
	LUT3 #(
		.INIT('hc8)
	) name14236 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		_w2215_,
		_w10616_,
		_w15586_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14237 (
		_w2054_,
		_w2059_,
		_w10616_,
		_w15586_,
		_w15587_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name14238 (
		\P3_InstQueue_reg[14][1]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w15588_
	);
	LUT4 #(
		.INIT('h153f)
	) name14239 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10646_,
		_w10659_,
		_w15589_
	);
	LUT2 #(
		.INIT('h2)
	) name14240 (
		_w2199_,
		_w15589_,
		_w15590_
	);
	LUT3 #(
		.INIT('h02)
	) name14241 (
		\buf2_reg[1]/NET0131 ,
		_w10617_,
		_w10684_,
		_w15591_
	);
	LUT3 #(
		.INIT('h01)
	) name14242 (
		_w15588_,
		_w15590_,
		_w15591_,
		_w15592_
	);
	LUT2 #(
		.INIT('hb)
	) name14243 (
		_w15587_,
		_w15592_,
		_w15593_
	);
	LUT3 #(
		.INIT('hc8)
	) name14244 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w2215_,
		_w10620_,
		_w15594_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14245 (
		_w2054_,
		_w2059_,
		_w10620_,
		_w15594_,
		_w15595_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14246 (
		\P3_InstQueue_reg[15][1]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w15596_
	);
	LUT4 #(
		.INIT('h135f)
	) name14247 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10614_,
		_w10659_,
		_w15597_
	);
	LUT2 #(
		.INIT('h2)
	) name14248 (
		_w2199_,
		_w15597_,
		_w15598_
	);
	LUT3 #(
		.INIT('h02)
	) name14249 (
		\buf2_reg[1]/NET0131 ,
		_w10693_,
		_w10694_,
		_w15599_
	);
	LUT3 #(
		.INIT('h01)
	) name14250 (
		_w15596_,
		_w15598_,
		_w15599_,
		_w15600_
	);
	LUT2 #(
		.INIT('hb)
	) name14251 (
		_w15595_,
		_w15600_,
		_w15601_
	);
	LUT3 #(
		.INIT('hc8)
	) name14252 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w2215_,
		_w10701_,
		_w15602_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14253 (
		_w2054_,
		_w2059_,
		_w10701_,
		_w15602_,
		_w15603_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14254 (
		\P3_InstQueue_reg[1][1]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w15604_
	);
	LUT4 #(
		.INIT('h153f)
	) name14255 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10616_,
		_w10620_,
		_w15605_
	);
	LUT2 #(
		.INIT('h2)
	) name14256 (
		_w2199_,
		_w15605_,
		_w15606_
	);
	LUT3 #(
		.INIT('h02)
	) name14257 (
		\buf2_reg[1]/NET0131 ,
		_w10704_,
		_w10705_,
		_w15607_
	);
	LUT3 #(
		.INIT('h01)
	) name14258 (
		_w15604_,
		_w15606_,
		_w15607_,
		_w15608_
	);
	LUT2 #(
		.INIT('hb)
	) name14259 (
		_w15603_,
		_w15608_,
		_w15609_
	);
	LUT3 #(
		.INIT('hc8)
	) name14260 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w2215_,
		_w10713_,
		_w15610_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14261 (
		_w2054_,
		_w2059_,
		_w10713_,
		_w15610_,
		_w15611_
	);
	LUT4 #(
		.INIT('h222a)
	) name14262 (
		\P3_InstQueue_reg[2][1]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w15612_
	);
	LUT4 #(
		.INIT('h135f)
	) name14263 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10611_,
		_w10620_,
		_w15613_
	);
	LUT2 #(
		.INIT('h2)
	) name14264 (
		_w2199_,
		_w15613_,
		_w15614_
	);
	LUT3 #(
		.INIT('h20)
	) name14265 (
		\buf2_reg[1]/NET0131 ,
		_w10716_,
		_w10717_,
		_w15615_
	);
	LUT3 #(
		.INIT('h01)
	) name14266 (
		_w15612_,
		_w15614_,
		_w15615_,
		_w15616_
	);
	LUT2 #(
		.INIT('hb)
	) name14267 (
		_w15611_,
		_w15616_,
		_w15617_
	);
	LUT3 #(
		.INIT('hc8)
	) name14268 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w2215_,
		_w10724_,
		_w15618_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14269 (
		_w2022_,
		_w2027_,
		_w10724_,
		_w15618_,
		_w15619_
	);
	LUT4 #(
		.INIT('h222a)
	) name14270 (
		\P3_InstQueue_reg[3][0]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w15620_
	);
	LUT4 #(
		.INIT('h153f)
	) name14271 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10611_,
		_w10701_,
		_w15621_
	);
	LUT2 #(
		.INIT('h2)
	) name14272 (
		_w2199_,
		_w15621_,
		_w15622_
	);
	LUT3 #(
		.INIT('h08)
	) name14273 (
		\buf2_reg[0]/NET0131 ,
		_w10712_,
		_w10727_,
		_w15623_
	);
	LUT3 #(
		.INIT('h01)
	) name14274 (
		_w15620_,
		_w15622_,
		_w15623_,
		_w15624_
	);
	LUT2 #(
		.INIT('hb)
	) name14275 (
		_w15619_,
		_w15624_,
		_w15625_
	);
	LUT3 #(
		.INIT('hc8)
	) name14276 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w2215_,
		_w10724_,
		_w15626_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14277 (
		_w2054_,
		_w2059_,
		_w10724_,
		_w15626_,
		_w15627_
	);
	LUT4 #(
		.INIT('h222a)
	) name14278 (
		\P3_InstQueue_reg[3][1]/NET0131 ,
		_w10622_,
		_w10712_,
		_w10727_,
		_w15628_
	);
	LUT4 #(
		.INIT('h153f)
	) name14279 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10611_,
		_w10701_,
		_w15629_
	);
	LUT2 #(
		.INIT('h2)
	) name14280 (
		_w2199_,
		_w15629_,
		_w15630_
	);
	LUT3 #(
		.INIT('h08)
	) name14281 (
		\buf2_reg[1]/NET0131 ,
		_w10712_,
		_w10727_,
		_w15631_
	);
	LUT3 #(
		.INIT('h01)
	) name14282 (
		_w15628_,
		_w15630_,
		_w15631_,
		_w15632_
	);
	LUT2 #(
		.INIT('hb)
	) name14283 (
		_w15627_,
		_w15632_,
		_w15633_
	);
	LUT3 #(
		.INIT('hc8)
	) name14284 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w2215_,
		_w10734_,
		_w15634_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14285 (
		_w2054_,
		_w2059_,
		_w10734_,
		_w15634_,
		_w15635_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14286 (
		\P3_InstQueue_reg[4][1]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w15636_
	);
	LUT4 #(
		.INIT('h153f)
	) name14287 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10701_,
		_w10713_,
		_w15637_
	);
	LUT2 #(
		.INIT('h2)
	) name14288 (
		_w2199_,
		_w15637_,
		_w15638_
	);
	LUT3 #(
		.INIT('h02)
	) name14289 (
		\buf2_reg[1]/NET0131 ,
		_w10737_,
		_w10738_,
		_w15639_
	);
	LUT3 #(
		.INIT('h01)
	) name14290 (
		_w15636_,
		_w15638_,
		_w15639_,
		_w15640_
	);
	LUT2 #(
		.INIT('hb)
	) name14291 (
		_w15635_,
		_w15640_,
		_w15641_
	);
	LUT3 #(
		.INIT('hc8)
	) name14292 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w2215_,
		_w10745_,
		_w15642_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14293 (
		_w2054_,
		_w2059_,
		_w10745_,
		_w15642_,
		_w15643_
	);
	LUT2 #(
		.INIT('h4)
	) name14294 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w10748_,
		_w15644_
	);
	LUT2 #(
		.INIT('h1)
	) name14295 (
		\buf2_reg[1]/NET0131 ,
		_w10748_,
		_w15645_
	);
	LUT3 #(
		.INIT('h02)
	) name14296 (
		_w10750_,
		_w15645_,
		_w15644_,
		_w15646_
	);
	LUT2 #(
		.INIT('h2)
	) name14297 (
		\P3_InstQueue_reg[5][1]/NET0131 ,
		_w10622_,
		_w15647_
	);
	LUT3 #(
		.INIT('h80)
	) name14298 (
		_w2194_,
		_w10749_,
		_w15561_,
		_w15648_
	);
	LUT2 #(
		.INIT('h1)
	) name14299 (
		_w15647_,
		_w15648_,
		_w15649_
	);
	LUT2 #(
		.INIT('h4)
	) name14300 (
		_w15646_,
		_w15649_,
		_w15650_
	);
	LUT2 #(
		.INIT('hb)
	) name14301 (
		_w15643_,
		_w15650_,
		_w15651_
	);
	LUT3 #(
		.INIT('hc8)
	) name14302 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w2215_,
		_w10758_,
		_w15652_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14303 (
		_w2054_,
		_w2059_,
		_w10758_,
		_w15652_,
		_w15653_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14304 (
		\P3_InstQueue_reg[6][1]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w15654_
	);
	LUT4 #(
		.INIT('h153f)
	) name14305 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10724_,
		_w10734_,
		_w15655_
	);
	LUT2 #(
		.INIT('h2)
	) name14306 (
		_w2199_,
		_w15655_,
		_w15656_
	);
	LUT3 #(
		.INIT('h02)
	) name14307 (
		\buf2_reg[1]/NET0131 ,
		_w10761_,
		_w10762_,
		_w15657_
	);
	LUT3 #(
		.INIT('h01)
	) name14308 (
		_w15654_,
		_w15656_,
		_w15657_,
		_w15658_
	);
	LUT2 #(
		.INIT('hb)
	) name14309 (
		_w15653_,
		_w15658_,
		_w15659_
	);
	LUT3 #(
		.INIT('hc8)
	) name14310 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w2215_,
		_w10633_,
		_w15660_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14311 (
		_w2022_,
		_w2027_,
		_w10633_,
		_w15660_,
		_w15661_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14312 (
		\P3_InstQueue_reg[7][0]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w15662_
	);
	LUT4 #(
		.INIT('h153f)
	) name14313 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10734_,
		_w10745_,
		_w15663_
	);
	LUT2 #(
		.INIT('h2)
	) name14314 (
		_w2199_,
		_w15663_,
		_w15664_
	);
	LUT3 #(
		.INIT('h02)
	) name14315 (
		\buf2_reg[0]/NET0131 ,
		_w10771_,
		_w10772_,
		_w15665_
	);
	LUT3 #(
		.INIT('h01)
	) name14316 (
		_w15662_,
		_w15664_,
		_w15665_,
		_w15666_
	);
	LUT2 #(
		.INIT('hb)
	) name14317 (
		_w15661_,
		_w15666_,
		_w15667_
	);
	LUT3 #(
		.INIT('hc8)
	) name14318 (
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w2215_,
		_w10633_,
		_w15668_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14319 (
		_w2054_,
		_w2059_,
		_w10633_,
		_w15668_,
		_w15669_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14320 (
		\P3_InstQueue_reg[7][1]/NET0131 ,
		_w10622_,
		_w10771_,
		_w10772_,
		_w15670_
	);
	LUT4 #(
		.INIT('h153f)
	) name14321 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10734_,
		_w10745_,
		_w15671_
	);
	LUT2 #(
		.INIT('h2)
	) name14322 (
		_w2199_,
		_w15671_,
		_w15672_
	);
	LUT3 #(
		.INIT('h02)
	) name14323 (
		\buf2_reg[1]/NET0131 ,
		_w10771_,
		_w10772_,
		_w15673_
	);
	LUT3 #(
		.INIT('h01)
	) name14324 (
		_w15670_,
		_w15672_,
		_w15673_,
		_w15674_
	);
	LUT2 #(
		.INIT('hb)
	) name14325 (
		_w15669_,
		_w15674_,
		_w15675_
	);
	LUT3 #(
		.INIT('hc8)
	) name14326 (
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w2215_,
		_w10635_,
		_w15676_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14327 (
		_w2054_,
		_w2059_,
		_w10635_,
		_w15676_,
		_w15677_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14328 (
		\P3_InstQueue_reg[8][1]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w15678_
	);
	LUT4 #(
		.INIT('h153f)
	) name14329 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10745_,
		_w10758_,
		_w15679_
	);
	LUT2 #(
		.INIT('h2)
	) name14330 (
		_w2199_,
		_w15679_,
		_w15680_
	);
	LUT3 #(
		.INIT('h02)
	) name14331 (
		\buf2_reg[1]/NET0131 ,
		_w10636_,
		_w10781_,
		_w15681_
	);
	LUT3 #(
		.INIT('h01)
	) name14332 (
		_w15678_,
		_w15680_,
		_w15681_,
		_w15682_
	);
	LUT2 #(
		.INIT('hb)
	) name14333 (
		_w15677_,
		_w15682_,
		_w15683_
	);
	LUT3 #(
		.INIT('hc8)
	) name14334 (
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w2215_,
		_w10652_,
		_w15684_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14335 (
		_w2054_,
		_w2059_,
		_w10652_,
		_w15684_,
		_w15685_
	);
	LUT4 #(
		.INIT('h135f)
	) name14336 (
		\buf2_reg[17]/NET0131 ,
		\buf2_reg[25]/NET0131 ,
		_w10633_,
		_w10758_,
		_w15686_
	);
	LUT4 #(
		.INIT('hef00)
	) name14337 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w15687_
	);
	LUT4 #(
		.INIT('h1000)
	) name14338 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[1]/NET0131 ,
		_w15688_
	);
	LUT4 #(
		.INIT('hddd0)
	) name14339 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w15687_,
		_w15688_,
		_w15689_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14340 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w15686_,
		_w15689_,
		_w15690_
	);
	LUT3 #(
		.INIT('ha8)
	) name14341 (
		_w3055_,
		_w15687_,
		_w15688_,
		_w15691_
	);
	LUT2 #(
		.INIT('h2)
	) name14342 (
		\P3_InstQueue_reg[9][1]/NET0131 ,
		_w10622_,
		_w15692_
	);
	LUT2 #(
		.INIT('h1)
	) name14343 (
		_w15691_,
		_w15692_,
		_w15693_
	);
	LUT2 #(
		.INIT('h4)
	) name14344 (
		_w15690_,
		_w15693_,
		_w15694_
	);
	LUT2 #(
		.INIT('hb)
	) name14345 (
		_w15685_,
		_w15694_,
		_w15695_
	);
	LUT4 #(
		.INIT('hfd80)
	) name14346 (
		\P2_State2_reg[0]/NET0131 ,
		\P2_State2_reg[1]/NET0131 ,
		\P2_State2_reg[2]/NET0131 ,
		\P2_State2_reg[3]/NET0131 ,
		_w15696_
	);
	LUT2 #(
		.INIT('h2)
	) name14347 (
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15696_,
		_w15697_
	);
	LUT2 #(
		.INIT('h1)
	) name14348 (
		\P2_Flush_reg/NET0131 ,
		\P2_InstQueueWr_Addr_reg[0]/NET0131 ,
		_w15698_
	);
	LUT4 #(
		.INIT('h002a)
	) name14349 (
		_w2205_,
		_w2206_,
		_w2207_,
		_w15698_,
		_w15699_
	);
	LUT3 #(
		.INIT('hfe)
	) name14350 (
		_w15516_,
		_w15699_,
		_w15697_,
		_w15700_
	);
	LUT4 #(
		.INIT('h8000)
	) name14351 (
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w15228_,
		_w15701_
	);
	LUT3 #(
		.INIT('h8a)
	) name14352 (
		\P3_Address_reg[24]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15702_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14353 (
		\P3_rEIP_reg[25]/NET0131 ,
		_w12118_,
		_w15235_,
		_w15237_,
		_w15703_
	);
	LUT2 #(
		.INIT('h1)
	) name14354 (
		_w15702_,
		_w15703_,
		_w15704_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14355 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w2110_,
		_w15229_,
		_w15704_,
		_w15705_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14356 (
		\P2_rEIP_reg[25]/NET0131 ,
		\P2_rEIP_reg[26]/NET0131 ,
		_w1609_,
		_w15253_,
		_w15706_
	);
	LUT3 #(
		.INIT('h8a)
	) name14357 (
		\P2_Address_reg[24]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15707_
	);
	LUT4 #(
		.INIT('h8000)
	) name14358 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w9780_,
		_w15259_,
		_w15708_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14359 (
		\P2_rEIP_reg[25]/NET0131 ,
		_w9781_,
		_w15262_,
		_w15259_,
		_w15709_
	);
	LUT2 #(
		.INIT('h1)
	) name14360 (
		_w15707_,
		_w15709_,
		_w15710_
	);
	LUT2 #(
		.INIT('hb)
	) name14361 (
		_w15706_,
		_w15710_,
		_w15711_
	);
	LUT3 #(
		.INIT('h13)
	) name14362 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15712_
	);
	LUT2 #(
		.INIT('h2)
	) name14363 (
		_w15287_,
		_w15712_,
		_w15713_
	);
	LUT4 #(
		.INIT('h1f00)
	) name14364 (
		_w11104_,
		_w11108_,
		_w15284_,
		_w15713_,
		_w15714_
	);
	LUT3 #(
		.INIT('hb0)
	) name14365 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[24]_pad ,
		_w15715_
	);
	LUT4 #(
		.INIT('h4888)
	) name14366 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w1856_,
		_w11107_,
		_w15278_,
		_w15716_
	);
	LUT2 #(
		.INIT('h1)
	) name14367 (
		_w15715_,
		_w15716_,
		_w15717_
	);
	LUT2 #(
		.INIT('hb)
	) name14368 (
		_w15714_,
		_w15717_,
		_w15718_
	);
	LUT3 #(
		.INIT('h8a)
	) name14369 (
		\P3_Address_reg[12]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15719_
	);
	LUT3 #(
		.INIT('h80)
	) name14370 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w11806_,
		_w15234_,
		_w15720_
	);
	LUT4 #(
		.INIT('h8000)
	) name14371 (
		\P3_rEIP_reg[11]/NET0131 ,
		\P3_rEIP_reg[12]/NET0131 ,
		_w11806_,
		_w15234_,
		_w15721_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14372 (
		\P3_rEIP_reg[13]/NET0131 ,
		_w15237_,
		_w15719_,
		_w15721_,
		_w15722_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14373 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w2110_,
		_w15223_,
		_w15722_,
		_w15723_
	);
	LUT4 #(
		.INIT('h8000)
	) name14374 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[13]/NET0131 ,
		_w15247_,
		_w15724_
	);
	LUT3 #(
		.INIT('h8a)
	) name14375 (
		\P2_Address_reg[12]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15725_
	);
	LUT3 #(
		.INIT('h80)
	) name14376 (
		_w9770_,
		_w9772_,
		_w15259_,
		_w15726_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14377 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w15262_,
		_w15725_,
		_w15726_,
		_w15727_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14378 (
		\P2_rEIP_reg[14]/NET0131 ,
		_w1609_,
		_w15724_,
		_w15727_,
		_w15728_
	);
	LUT3 #(
		.INIT('h48)
	) name14379 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w1856_,
		_w15275_,
		_w15729_
	);
	LUT3 #(
		.INIT('hb0)
	) name14380 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[12]_pad ,
		_w15730_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14381 (
		\P1_rEIP_reg[13]/NET0131 ,
		_w10813_,
		_w15284_,
		_w15287_,
		_w15731_
	);
	LUT2 #(
		.INIT('h1)
	) name14382 (
		_w15730_,
		_w15731_,
		_w15732_
	);
	LUT2 #(
		.INIT('hb)
	) name14383 (
		_w15729_,
		_w15732_,
		_w15733_
	);
	LUT3 #(
		.INIT('hc8)
	) name14384 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		_w2215_,
		_w10611_,
		_w15734_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14385 (
		_w2022_,
		_w2027_,
		_w10611_,
		_w15734_,
		_w15735_
	);
	LUT4 #(
		.INIT('h20aa)
	) name14386 (
		\P3_InstQueue_reg[0][0]/NET0131 ,
		_w10618_,
		_w10621_,
		_w10622_,
		_w15736_
	);
	LUT4 #(
		.INIT('h153f)
	) name14387 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10614_,
		_w10616_,
		_w15737_
	);
	LUT2 #(
		.INIT('h2)
	) name14388 (
		_w2199_,
		_w15737_,
		_w15738_
	);
	LUT3 #(
		.INIT('h02)
	) name14389 (
		\buf2_reg[0]/NET0131 ,
		_w10618_,
		_w10621_,
		_w15739_
	);
	LUT3 #(
		.INIT('h01)
	) name14390 (
		_w15736_,
		_w15738_,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('hb)
	) name14391 (
		_w15735_,
		_w15740_,
		_w15741_
	);
	LUT3 #(
		.INIT('hc8)
	) name14392 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		_w2215_,
		_w10630_,
		_w15742_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14393 (
		_w2022_,
		_w2027_,
		_w10630_,
		_w15742_,
		_w15743_
	);
	LUT4 #(
		.INIT('h222a)
	) name14394 (
		\P3_InstQueue_reg[10][0]/NET0131 ,
		_w10622_,
		_w10637_,
		_w10639_,
		_w15744_
	);
	LUT4 #(
		.INIT('h153f)
	) name14395 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10633_,
		_w10635_,
		_w15745_
	);
	LUT2 #(
		.INIT('h2)
	) name14396 (
		_w2199_,
		_w15745_,
		_w15746_
	);
	LUT3 #(
		.INIT('h20)
	) name14397 (
		\buf2_reg[0]/NET0131 ,
		_w10637_,
		_w10639_,
		_w15747_
	);
	LUT3 #(
		.INIT('h01)
	) name14398 (
		_w15744_,
		_w15746_,
		_w15747_,
		_w15748_
	);
	LUT2 #(
		.INIT('hb)
	) name14399 (
		_w15743_,
		_w15748_,
		_w15749_
	);
	LUT3 #(
		.INIT('hc8)
	) name14400 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w2215_,
		_w10659_,
		_w15750_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14401 (
		_w2022_,
		_w2027_,
		_w10659_,
		_w15750_,
		_w15751_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14402 (
		\P3_InstQueue_reg[12][0]/NET0131 ,
		_w10622_,
		_w10662_,
		_w10663_,
		_w15752_
	);
	LUT4 #(
		.INIT('h135f)
	) name14403 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10630_,
		_w10652_,
		_w15753_
	);
	LUT2 #(
		.INIT('h2)
	) name14404 (
		_w2199_,
		_w15753_,
		_w15754_
	);
	LUT3 #(
		.INIT('h02)
	) name14405 (
		\buf2_reg[0]/NET0131 ,
		_w10662_,
		_w10663_,
		_w15755_
	);
	LUT3 #(
		.INIT('h01)
	) name14406 (
		_w15752_,
		_w15754_,
		_w15755_,
		_w15756_
	);
	LUT2 #(
		.INIT('hb)
	) name14407 (
		_w15751_,
		_w15756_,
		_w15757_
	);
	LUT3 #(
		.INIT('hc8)
	) name14408 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w2215_,
		_w10614_,
		_w15758_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14409 (
		_w2022_,
		_w2027_,
		_w10614_,
		_w15758_,
		_w15759_
	);
	LUT2 #(
		.INIT('h4)
	) name14410 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w10672_,
		_w15760_
	);
	LUT2 #(
		.INIT('h1)
	) name14411 (
		\buf2_reg[0]/NET0131 ,
		_w10672_,
		_w15761_
	);
	LUT3 #(
		.INIT('h02)
	) name14412 (
		_w10674_,
		_w15761_,
		_w15760_,
		_w15762_
	);
	LUT2 #(
		.INIT('h2)
	) name14413 (
		\P3_InstQueue_reg[13][0]/NET0131 ,
		_w10622_,
		_w15763_
	);
	LUT3 #(
		.INIT('h80)
	) name14414 (
		_w2194_,
		_w10673_,
		_w15551_,
		_w15764_
	);
	LUT2 #(
		.INIT('h1)
	) name14415 (
		_w15763_,
		_w15764_,
		_w15765_
	);
	LUT2 #(
		.INIT('h4)
	) name14416 (
		_w15762_,
		_w15765_,
		_w15766_
	);
	LUT2 #(
		.INIT('hb)
	) name14417 (
		_w15759_,
		_w15766_,
		_w15767_
	);
	LUT3 #(
		.INIT('hc8)
	) name14418 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w2215_,
		_w10616_,
		_w15768_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14419 (
		_w2022_,
		_w2027_,
		_w10616_,
		_w15768_,
		_w15769_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name14420 (
		\P3_InstQueue_reg[14][0]/NET0131 ,
		_w10617_,
		_w10622_,
		_w10684_,
		_w15770_
	);
	LUT4 #(
		.INIT('h153f)
	) name14421 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10646_,
		_w10659_,
		_w15771_
	);
	LUT2 #(
		.INIT('h2)
	) name14422 (
		_w2199_,
		_w15771_,
		_w15772_
	);
	LUT3 #(
		.INIT('h02)
	) name14423 (
		\buf2_reg[0]/NET0131 ,
		_w10617_,
		_w10684_,
		_w15773_
	);
	LUT3 #(
		.INIT('h01)
	) name14424 (
		_w15770_,
		_w15772_,
		_w15773_,
		_w15774_
	);
	LUT2 #(
		.INIT('hb)
	) name14425 (
		_w15769_,
		_w15774_,
		_w15775_
	);
	LUT3 #(
		.INIT('hc8)
	) name14426 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w2215_,
		_w10620_,
		_w15776_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14427 (
		_w2022_,
		_w2027_,
		_w10620_,
		_w15776_,
		_w15777_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14428 (
		\P3_InstQueue_reg[15][0]/NET0131 ,
		_w10622_,
		_w10693_,
		_w10694_,
		_w15778_
	);
	LUT4 #(
		.INIT('h135f)
	) name14429 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10614_,
		_w10659_,
		_w15779_
	);
	LUT2 #(
		.INIT('h2)
	) name14430 (
		_w2199_,
		_w15779_,
		_w15780_
	);
	LUT3 #(
		.INIT('h02)
	) name14431 (
		\buf2_reg[0]/NET0131 ,
		_w10693_,
		_w10694_,
		_w15781_
	);
	LUT3 #(
		.INIT('h01)
	) name14432 (
		_w15778_,
		_w15780_,
		_w15781_,
		_w15782_
	);
	LUT2 #(
		.INIT('hb)
	) name14433 (
		_w15777_,
		_w15782_,
		_w15783_
	);
	LUT3 #(
		.INIT('hc8)
	) name14434 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w2215_,
		_w10701_,
		_w15784_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14435 (
		_w2022_,
		_w2027_,
		_w10701_,
		_w15784_,
		_w15785_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14436 (
		\P3_InstQueue_reg[1][0]/NET0131 ,
		_w10622_,
		_w10704_,
		_w10705_,
		_w15786_
	);
	LUT4 #(
		.INIT('h153f)
	) name14437 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10616_,
		_w10620_,
		_w15787_
	);
	LUT2 #(
		.INIT('h2)
	) name14438 (
		_w2199_,
		_w15787_,
		_w15788_
	);
	LUT3 #(
		.INIT('h02)
	) name14439 (
		\buf2_reg[0]/NET0131 ,
		_w10704_,
		_w10705_,
		_w15789_
	);
	LUT3 #(
		.INIT('h01)
	) name14440 (
		_w15786_,
		_w15788_,
		_w15789_,
		_w15790_
	);
	LUT2 #(
		.INIT('hb)
	) name14441 (
		_w15785_,
		_w15790_,
		_w15791_
	);
	LUT3 #(
		.INIT('hc8)
	) name14442 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w2215_,
		_w10713_,
		_w15792_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14443 (
		_w2022_,
		_w2027_,
		_w10713_,
		_w15792_,
		_w15793_
	);
	LUT4 #(
		.INIT('h222a)
	) name14444 (
		\P3_InstQueue_reg[2][0]/NET0131 ,
		_w10622_,
		_w10716_,
		_w10717_,
		_w15794_
	);
	LUT4 #(
		.INIT('h135f)
	) name14445 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10611_,
		_w10620_,
		_w15795_
	);
	LUT2 #(
		.INIT('h2)
	) name14446 (
		_w2199_,
		_w15795_,
		_w15796_
	);
	LUT3 #(
		.INIT('h20)
	) name14447 (
		\buf2_reg[0]/NET0131 ,
		_w10716_,
		_w10717_,
		_w15797_
	);
	LUT3 #(
		.INIT('h01)
	) name14448 (
		_w15794_,
		_w15796_,
		_w15797_,
		_w15798_
	);
	LUT2 #(
		.INIT('hb)
	) name14449 (
		_w15793_,
		_w15798_,
		_w15799_
	);
	LUT3 #(
		.INIT('hc8)
	) name14450 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w2215_,
		_w10734_,
		_w15800_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14451 (
		_w2022_,
		_w2027_,
		_w10734_,
		_w15800_,
		_w15801_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14452 (
		\P3_InstQueue_reg[4][0]/NET0131 ,
		_w10622_,
		_w10737_,
		_w10738_,
		_w15802_
	);
	LUT4 #(
		.INIT('h153f)
	) name14453 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10701_,
		_w10713_,
		_w15803_
	);
	LUT2 #(
		.INIT('h2)
	) name14454 (
		_w2199_,
		_w15803_,
		_w15804_
	);
	LUT3 #(
		.INIT('h02)
	) name14455 (
		\buf2_reg[0]/NET0131 ,
		_w10737_,
		_w10738_,
		_w15805_
	);
	LUT3 #(
		.INIT('h01)
	) name14456 (
		_w15802_,
		_w15804_,
		_w15805_,
		_w15806_
	);
	LUT2 #(
		.INIT('hb)
	) name14457 (
		_w15801_,
		_w15806_,
		_w15807_
	);
	LUT3 #(
		.INIT('hc8)
	) name14458 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w2215_,
		_w10745_,
		_w15808_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14459 (
		_w2022_,
		_w2027_,
		_w10745_,
		_w15808_,
		_w15809_
	);
	LUT2 #(
		.INIT('h4)
	) name14460 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w10748_,
		_w15810_
	);
	LUT2 #(
		.INIT('h1)
	) name14461 (
		\buf2_reg[0]/NET0131 ,
		_w10748_,
		_w15811_
	);
	LUT3 #(
		.INIT('h02)
	) name14462 (
		_w10750_,
		_w15811_,
		_w15810_,
		_w15812_
	);
	LUT2 #(
		.INIT('h2)
	) name14463 (
		\P3_InstQueue_reg[5][0]/NET0131 ,
		_w10622_,
		_w15813_
	);
	LUT3 #(
		.INIT('h80)
	) name14464 (
		_w2194_,
		_w10749_,
		_w15551_,
		_w15814_
	);
	LUT2 #(
		.INIT('h1)
	) name14465 (
		_w15813_,
		_w15814_,
		_w15815_
	);
	LUT2 #(
		.INIT('h4)
	) name14466 (
		_w15812_,
		_w15815_,
		_w15816_
	);
	LUT2 #(
		.INIT('hb)
	) name14467 (
		_w15809_,
		_w15816_,
		_w15817_
	);
	LUT3 #(
		.INIT('hc8)
	) name14468 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w2215_,
		_w10758_,
		_w15818_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14469 (
		_w2022_,
		_w2027_,
		_w10758_,
		_w15818_,
		_w15819_
	);
	LUT4 #(
		.INIT('h2a22)
	) name14470 (
		\P3_InstQueue_reg[6][0]/NET0131 ,
		_w10622_,
		_w10761_,
		_w10762_,
		_w15820_
	);
	LUT4 #(
		.INIT('h153f)
	) name14471 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10724_,
		_w10734_,
		_w15821_
	);
	LUT2 #(
		.INIT('h2)
	) name14472 (
		_w2199_,
		_w15821_,
		_w15822_
	);
	LUT3 #(
		.INIT('h02)
	) name14473 (
		\buf2_reg[0]/NET0131 ,
		_w10761_,
		_w10762_,
		_w15823_
	);
	LUT3 #(
		.INIT('h01)
	) name14474 (
		_w15820_,
		_w15822_,
		_w15823_,
		_w15824_
	);
	LUT2 #(
		.INIT('hb)
	) name14475 (
		_w15819_,
		_w15824_,
		_w15825_
	);
	LUT3 #(
		.INIT('hc8)
	) name14476 (
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w2215_,
		_w10635_,
		_w15826_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14477 (
		_w2022_,
		_w2027_,
		_w10635_,
		_w15826_,
		_w15827_
	);
	LUT4 #(
		.INIT('h22a2)
	) name14478 (
		\P3_InstQueue_reg[8][0]/NET0131 ,
		_w10622_,
		_w10636_,
		_w10781_,
		_w15828_
	);
	LUT4 #(
		.INIT('h153f)
	) name14479 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10745_,
		_w10758_,
		_w15829_
	);
	LUT2 #(
		.INIT('h2)
	) name14480 (
		_w2199_,
		_w15829_,
		_w15830_
	);
	LUT3 #(
		.INIT('h02)
	) name14481 (
		\buf2_reg[0]/NET0131 ,
		_w10636_,
		_w10781_,
		_w15831_
	);
	LUT3 #(
		.INIT('h01)
	) name14482 (
		_w15828_,
		_w15830_,
		_w15831_,
		_w15832_
	);
	LUT2 #(
		.INIT('hb)
	) name14483 (
		_w15827_,
		_w15832_,
		_w15833_
	);
	LUT3 #(
		.INIT('hc8)
	) name14484 (
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w2215_,
		_w10652_,
		_w15834_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14485 (
		_w2022_,
		_w2027_,
		_w10652_,
		_w15834_,
		_w15835_
	);
	LUT4 #(
		.INIT('h135f)
	) name14486 (
		\buf2_reg[16]/NET0131 ,
		\buf2_reg[24]/NET0131 ,
		_w10633_,
		_w10758_,
		_w15836_
	);
	LUT4 #(
		.INIT('hef00)
	) name14487 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w15837_
	);
	LUT4 #(
		.INIT('h1000)
	) name14488 (
		\P3_InstQueueWr_Addr_reg[1]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[2]/NET0131 ,
		\P3_InstQueueWr_Addr_reg[3]/NET0131 ,
		\buf2_reg[0]/NET0131 ,
		_w15838_
	);
	LUT4 #(
		.INIT('hddd0)
	) name14489 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w10772_,
		_w15837_,
		_w15838_,
		_w15839_
	);
	LUT4 #(
		.INIT('hcc08)
	) name14490 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w15836_,
		_w15839_,
		_w15840_
	);
	LUT3 #(
		.INIT('ha8)
	) name14491 (
		_w3055_,
		_w15837_,
		_w15838_,
		_w15841_
	);
	LUT2 #(
		.INIT('h2)
	) name14492 (
		\P3_InstQueue_reg[9][0]/NET0131 ,
		_w10622_,
		_w15842_
	);
	LUT2 #(
		.INIT('h1)
	) name14493 (
		_w15841_,
		_w15842_,
		_w15843_
	);
	LUT2 #(
		.INIT('h4)
	) name14494 (
		_w15840_,
		_w15843_,
		_w15844_
	);
	LUT2 #(
		.INIT('hb)
	) name14495 (
		_w15835_,
		_w15844_,
		_w15845_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14496 (
		\P3_rEIP_reg[21]/NET0131 ,
		\P3_rEIP_reg[22]/NET0131 ,
		_w2110_,
		_w15226_,
		_w15846_
	);
	LUT3 #(
		.INIT('h8a)
	) name14497 (
		\P3_Address_reg[20]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15847_
	);
	LUT3 #(
		.INIT('h80)
	) name14498 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w12026_,
		_w15460_,
		_w15848_
	);
	LUT4 #(
		.INIT('h8000)
	) name14499 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[21]/NET0131 ,
		_w12026_,
		_w15460_,
		_w15849_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14500 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w15237_,
		_w15847_,
		_w15848_,
		_w15850_
	);
	LUT2 #(
		.INIT('hb)
	) name14501 (
		_w15846_,
		_w15850_,
		_w15851_
	);
	LUT3 #(
		.INIT('h8a)
	) name14502 (
		\P2_Address_reg[20]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15852_
	);
	LUT4 #(
		.INIT('h8000)
	) name14503 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w9778_,
		_w15259_,
		_w15853_
	);
	LUT4 #(
		.INIT('h1333)
	) name14504 (
		\P2_rEIP_reg[20]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w9778_,
		_w15259_,
		_w15854_
	);
	LUT4 #(
		.INIT('h3331)
	) name14505 (
		_w15262_,
		_w15852_,
		_w15854_,
		_w15853_,
		_w15855_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14506 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w1609_,
		_w15251_,
		_w15855_,
		_w15856_
	);
	LUT3 #(
		.INIT('h80)
	) name14507 (
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w15278_,
		_w15857_
	);
	LUT4 #(
		.INIT('h8000)
	) name14508 (
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		\P1_rEIP_reg[20]/NET0131 ,
		_w15278_,
		_w15858_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14509 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w1856_,
		_w15858_,
		_w15859_
	);
	LUT3 #(
		.INIT('hb0)
	) name14510 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[20]_pad ,
		_w15860_
	);
	LUT4 #(
		.INIT('h8000)
	) name14511 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10858_,
		_w15284_,
		_w15861_
	);
	LUT3 #(
		.INIT('h80)
	) name14512 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w10973_,
		_w15861_,
		_w15862_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14513 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w10973_,
		_w15287_,
		_w15861_,
		_w15863_
	);
	LUT2 #(
		.INIT('h1)
	) name14514 (
		_w15860_,
		_w15863_,
		_w15864_
	);
	LUT2 #(
		.INIT('hb)
	) name14515 (
		_w15859_,
		_w15864_,
		_w15865_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14516 (
		\P3_rEIP_reg[10]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w2110_,
		_w15220_,
		_w15866_
	);
	LUT3 #(
		.INIT('h8a)
	) name14517 (
		\P3_Address_reg[8]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15867_
	);
	LUT4 #(
		.INIT('h9300)
	) name14518 (
		\P3_rEIP_reg[8]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w11804_,
		_w15234_,
		_w15868_
	);
	LUT3 #(
		.INIT('h07)
	) name14519 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		\P3_rEIP_reg[9]/NET0131 ,
		_w15869_
	);
	LUT2 #(
		.INIT('h2)
	) name14520 (
		_w15237_,
		_w15869_,
		_w15870_
	);
	LUT3 #(
		.INIT('h45)
	) name14521 (
		_w15867_,
		_w15868_,
		_w15870_,
		_w15871_
	);
	LUT2 #(
		.INIT('hb)
	) name14522 (
		_w15866_,
		_w15871_,
		_w15872_
	);
	LUT3 #(
		.INIT('h8a)
	) name14523 (
		\P2_Address_reg[8]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15873_
	);
	LUT3 #(
		.INIT('h07)
	) name14524 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w15874_
	);
	LUT2 #(
		.INIT('h2)
	) name14525 (
		_w15262_,
		_w15874_,
		_w15875_
	);
	LUT4 #(
		.INIT('h040f)
	) name14526 (
		_w11783_,
		_w15259_,
		_w15873_,
		_w15875_,
		_w15876_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14527 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w1609_,
		_w15246_,
		_w15876_,
		_w15877_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14528 (
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w1856_,
		_w15272_,
		_w15878_
	);
	LUT3 #(
		.INIT('hb0)
	) name14529 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[8]_pad ,
		_w15879_
	);
	LUT4 #(
		.INIT('h8000)
	) name14530 (
		\P1_rEIP_reg[5]/NET0131 ,
		\P1_rEIP_reg[6]/NET0131 ,
		_w10810_,
		_w15284_,
		_w15880_
	);
	LUT3 #(
		.INIT('h80)
	) name14531 (
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15880_,
		_w15881_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14532 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w15287_,
		_w15879_,
		_w15881_,
		_w15882_
	);
	LUT2 #(
		.INIT('hb)
	) name14533 (
		_w15878_,
		_w15882_,
		_w15883_
	);
	LUT3 #(
		.INIT('h48)
	) name14534 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w2110_,
		_w15218_,
		_w15884_
	);
	LUT3 #(
		.INIT('h8a)
	) name14535 (
		\P3_Address_reg[4]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15885_
	);
	LUT3 #(
		.INIT('h80)
	) name14536 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15886_
	);
	LUT4 #(
		.INIT('h8000)
	) name14537 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w15887_
	);
	LUT4 #(
		.INIT('h070f)
	) name14538 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		\P3_rEIP_reg[5]/NET0131 ,
		_w15887_,
		_w15888_
	);
	LUT3 #(
		.INIT('h80)
	) name14539 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w11803_,
		_w15234_,
		_w15889_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14540 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w11803_,
		_w15234_,
		_w15237_,
		_w15890_
	);
	LUT3 #(
		.INIT('h45)
	) name14541 (
		_w15885_,
		_w15888_,
		_w15890_,
		_w15891_
	);
	LUT2 #(
		.INIT('hb)
	) name14542 (
		_w15884_,
		_w15891_,
		_w15892_
	);
	LUT4 #(
		.INIT('h8000)
	) name14543 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w15243_,
		_w15893_
	);
	LUT3 #(
		.INIT('h48)
	) name14544 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w1609_,
		_w15893_,
		_w15894_
	);
	LUT3 #(
		.INIT('h8a)
	) name14545 (
		\P2_Address_reg[4]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15895_
	);
	LUT3 #(
		.INIT('h80)
	) name14546 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15896_
	);
	LUT4 #(
		.INIT('h8000)
	) name14547 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15897_
	);
	LUT3 #(
		.INIT('h80)
	) name14548 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15897_,
		_w15898_
	);
	LUT4 #(
		.INIT('h8000)
	) name14549 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		\P2_rEIP_reg[5]/NET0131 ,
		_w15897_,
		_w15899_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14550 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w15262_,
		_w15895_,
		_w15898_,
		_w15900_
	);
	LUT2 #(
		.INIT('hb)
	) name14551 (
		_w15894_,
		_w15900_,
		_w15901_
	);
	LUT3 #(
		.INIT('h48)
	) name14552 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w1856_,
		_w15270_,
		_w15902_
	);
	LUT3 #(
		.INIT('hb0)
	) name14553 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[4]_pad ,
		_w15903_
	);
	LUT3 #(
		.INIT('h80)
	) name14554 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15904_
	);
	LUT4 #(
		.INIT('h8000)
	) name14555 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		\P1_rEIP_reg[2]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15905_
	);
	LUT3 #(
		.INIT('h80)
	) name14556 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15905_,
		_w15906_
	);
	LUT4 #(
		.INIT('h8000)
	) name14557 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		\P1_rEIP_reg[5]/NET0131 ,
		_w15905_,
		_w15907_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14558 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w15287_,
		_w15903_,
		_w15906_,
		_w15908_
	);
	LUT2 #(
		.INIT('hb)
	) name14559 (
		_w15902_,
		_w15908_,
		_w15909_
	);
	LUT3 #(
		.INIT('hb0)
	) name14560 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[15]_pad ,
		_w15910_
	);
	LUT3 #(
		.INIT('h80)
	) name14561 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10814_,
		_w15284_,
		_w15911_
	);
	LUT4 #(
		.INIT('h8000)
	) name14562 (
		\P1_rEIP_reg[14]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w10814_,
		_w15284_,
		_w15912_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14563 (
		\P1_rEIP_reg[16]/NET0131 ,
		_w15287_,
		_w15910_,
		_w15912_,
		_w15913_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14564 (
		\P1_rEIP_reg[17]/NET0131 ,
		_w1856_,
		_w15277_,
		_w15913_,
		_w15914_
	);
	LUT3 #(
		.INIT('h8a)
	) name14565 (
		\P3_Address_reg[15]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15915_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14566 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w15237_,
		_w15460_,
		_w15915_,
		_w15916_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14567 (
		\P3_rEIP_reg[17]/NET0131 ,
		_w2110_,
		_w15225_,
		_w15916_,
		_w15917_
	);
	LUT3 #(
		.INIT('h8a)
	) name14568 (
		\P3_Address_reg[27]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15918_
	);
	LUT3 #(
		.INIT('h80)
	) name14569 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w12119_,
		_w15235_,
		_w15919_
	);
	LUT4 #(
		.INIT('h8000)
	) name14570 (
		\P3_rEIP_reg[26]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w12119_,
		_w15235_,
		_w15920_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14571 (
		_w12119_,
		_w12192_,
		_w15235_,
		_w15237_,
		_w15921_
	);
	LUT4 #(
		.INIT('h0133)
	) name14572 (
		\P3_rEIP_reg[28]/NET0131 ,
		_w15918_,
		_w15920_,
		_w15921_,
		_w15922_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14573 (
		\P3_rEIP_reg[29]/NET0131 ,
		_w2110_,
		_w15230_,
		_w15922_,
		_w15923_
	);
	LUT4 #(
		.INIT('h8000)
	) name14574 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w9775_,
		_w15247_,
		_w15924_
	);
	LUT4 #(
		.INIT('h4888)
	) name14575 (
		\P2_rEIP_reg[17]/NET0131 ,
		_w1609_,
		_w9775_,
		_w15248_,
		_w15925_
	);
	LUT3 #(
		.INIT('h8a)
	) name14576 (
		\P2_Address_reg[15]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15926_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14577 (
		\P2_rEIP_reg[16]/NET0131 ,
		_w9774_,
		_w15262_,
		_w15726_,
		_w15927_
	);
	LUT2 #(
		.INIT('h1)
	) name14578 (
		_w15926_,
		_w15927_,
		_w15928_
	);
	LUT2 #(
		.INIT('hb)
	) name14579 (
		_w15925_,
		_w15928_,
		_w15929_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14580 (
		\P2_rEIP_reg[28]/NET0131 ,
		\P2_rEIP_reg[29]/NET0131 ,
		_w1609_,
		_w15255_,
		_w15930_
	);
	LUT3 #(
		.INIT('h8a)
	) name14581 (
		\P2_Address_reg[27]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15931_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14582 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w15262_,
		_w15261_,
		_w15931_,
		_w15932_
	);
	LUT2 #(
		.INIT('hb)
	) name14583 (
		_w15930_,
		_w15932_,
		_w15933_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14584 (
		\P1_rEIP_reg[28]/NET0131 ,
		\P1_rEIP_reg[29]/NET0131 ,
		_w1856_,
		_w15280_,
		_w15934_
	);
	LUT3 #(
		.INIT('hb0)
	) name14585 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[27]_pad ,
		_w15935_
	);
	LUT4 #(
		.INIT('h009f)
	) name14586 (
		\P1_rEIP_reg[28]/NET0131 ,
		_w15285_,
		_w15287_,
		_w15935_,
		_w15936_
	);
	LUT2 #(
		.INIT('hb)
	) name14587 (
		_w15934_,
		_w15936_,
		_w15937_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14588 (
		\P3_rEIP_reg[24]/NET0131 ,
		\P3_rEIP_reg[25]/NET0131 ,
		_w2110_,
		_w15228_,
		_w15938_
	);
	LUT3 #(
		.INIT('h8a)
	) name14589 (
		\P3_Address_reg[23]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15939_
	);
	LUT4 #(
		.INIT('h6c00)
	) name14590 (
		\P3_rEIP_reg[23]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w15235_,
		_w15237_,
		_w15940_
	);
	LUT2 #(
		.INIT('h1)
	) name14591 (
		_w15939_,
		_w15940_,
		_w15941_
	);
	LUT2 #(
		.INIT('hb)
	) name14592 (
		_w15938_,
		_w15941_,
		_w15942_
	);
	LUT3 #(
		.INIT('h8a)
	) name14593 (
		\P2_Address_reg[23]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15943_
	);
	LUT4 #(
		.INIT('h1333)
	) name14594 (
		\P2_rEIP_reg[23]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w9780_,
		_w15259_,
		_w15944_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name14595 (
		_w15262_,
		_w15708_,
		_w15943_,
		_w15944_,
		_w15945_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14596 (
		\P2_rEIP_reg[25]/NET0131 ,
		_w1609_,
		_w15253_,
		_w15945_,
		_w15946_
	);
	LUT3 #(
		.INIT('h2a)
	) name14597 (
		_w1856_,
		_w11107_,
		_w15278_,
		_w15947_
	);
	LUT4 #(
		.INIT('hea00)
	) name14598 (
		\P1_rEIP_reg[25]/NET0131 ,
		_w11105_,
		_w15858_,
		_w15947_,
		_w15948_
	);
	LUT3 #(
		.INIT('hb0)
	) name14599 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[23]_pad ,
		_w15949_
	);
	LUT3 #(
		.INIT('h80)
	) name14600 (
		_w10973_,
		_w11024_,
		_w15861_,
		_w15950_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14601 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w15287_,
		_w15949_,
		_w15950_,
		_w15951_
	);
	LUT2 #(
		.INIT('hb)
	) name14602 (
		_w15948_,
		_w15951_,
		_w15952_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14603 (
		\P3_rEIP_reg[12]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w2110_,
		_w15222_,
		_w15953_
	);
	LUT3 #(
		.INIT('h8a)
	) name14604 (
		\P3_Address_reg[11]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15954_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14605 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w15237_,
		_w15720_,
		_w15954_,
		_w15955_
	);
	LUT2 #(
		.INIT('hb)
	) name14606 (
		_w15953_,
		_w15955_,
		_w15956_
	);
	LUT3 #(
		.INIT('h8a)
	) name14607 (
		\P2_Address_reg[11]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15957_
	);
	LUT4 #(
		.INIT('h9500)
	) name14608 (
		\P2_rEIP_reg[12]/NET0131 ,
		_w9771_,
		_w9770_,
		_w15259_,
		_w15958_
	);
	LUT3 #(
		.INIT('h13)
	) name14609 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w15959_
	);
	LUT2 #(
		.INIT('h2)
	) name14610 (
		_w15262_,
		_w15959_,
		_w15960_
	);
	LUT3 #(
		.INIT('h45)
	) name14611 (
		_w15957_,
		_w15958_,
		_w15960_,
		_w15961_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14612 (
		\P2_rEIP_reg[13]/NET0131 ,
		_w1609_,
		_w15248_,
		_w15961_,
		_w15962_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14613 (
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w1856_,
		_w15274_,
		_w15963_
	);
	LUT3 #(
		.INIT('hb0)
	) name14614 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[11]_pad ,
		_w15964_
	);
	LUT4 #(
		.INIT('h9300)
	) name14615 (
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		_w10812_,
		_w15284_,
		_w15965_
	);
	LUT3 #(
		.INIT('h13)
	) name14616 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[12]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w15966_
	);
	LUT2 #(
		.INIT('h2)
	) name14617 (
		_w15287_,
		_w15966_,
		_w15967_
	);
	LUT3 #(
		.INIT('h45)
	) name14618 (
		_w15964_,
		_w15965_,
		_w15967_,
		_w15968_
	);
	LUT2 #(
		.INIT('hb)
	) name14619 (
		_w15963_,
		_w15968_,
		_w15969_
	);
	LUT3 #(
		.INIT('h48)
	) name14620 (
		\P3_rEIP_reg[5]/NET0131 ,
		_w2110_,
		_w15217_,
		_w15970_
	);
	LUT3 #(
		.INIT('h8a)
	) name14621 (
		\P3_Address_reg[3]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15971_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14622 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w15237_,
		_w15887_,
		_w15972_
	);
	LUT2 #(
		.INIT('h1)
	) name14623 (
		_w15971_,
		_w15972_,
		_w15973_
	);
	LUT2 #(
		.INIT('hb)
	) name14624 (
		_w15970_,
		_w15973_,
		_w15974_
	);
	LUT3 #(
		.INIT('h48)
	) name14625 (
		\P2_rEIP_reg[5]/NET0131 ,
		_w1609_,
		_w15244_,
		_w15975_
	);
	LUT3 #(
		.INIT('h8a)
	) name14626 (
		\P2_Address_reg[3]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15976_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14627 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w15262_,
		_w15897_,
		_w15977_
	);
	LUT2 #(
		.INIT('h1)
	) name14628 (
		_w15976_,
		_w15977_,
		_w15978_
	);
	LUT2 #(
		.INIT('hb)
	) name14629 (
		_w15975_,
		_w15978_,
		_w15979_
	);
	LUT3 #(
		.INIT('h48)
	) name14630 (
		\P1_rEIP_reg[5]/NET0131 ,
		_w1856_,
		_w15269_,
		_w15980_
	);
	LUT3 #(
		.INIT('hb0)
	) name14631 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[3]_pad ,
		_w15981_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14632 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w15287_,
		_w15905_,
		_w15982_
	);
	LUT2 #(
		.INIT('h1)
	) name14633 (
		_w15981_,
		_w15982_,
		_w15983_
	);
	LUT2 #(
		.INIT('hb)
	) name14634 (
		_w15980_,
		_w15983_,
		_w15984_
	);
	LUT3 #(
		.INIT('h48)
	) name14635 (
		\P3_rEIP_reg[21]/NET0131 ,
		_w2110_,
		_w15226_,
		_w15985_
	);
	LUT3 #(
		.INIT('h8a)
	) name14636 (
		\P3_Address_reg[19]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w15986_
	);
	LUT4 #(
		.INIT('h8000)
	) name14637 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11923_,
		_w11970_,
		_w15234_,
		_w15987_
	);
	LUT4 #(
		.INIT('h70f0)
	) name14638 (
		\P3_rEIP_reg[16]/NET0131 ,
		_w12026_,
		_w15237_,
		_w15460_,
		_w15988_
	);
	LUT4 #(
		.INIT('h0133)
	) name14639 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w15986_,
		_w15987_,
		_w15988_,
		_w15989_
	);
	LUT2 #(
		.INIT('hb)
	) name14640 (
		_w15985_,
		_w15989_,
		_w15990_
	);
	LUT3 #(
		.INIT('h8a)
	) name14641 (
		\P2_Address_reg[19]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w15991_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14642 (
		\P2_rEIP_reg[20]/NET0131 ,
		_w9778_,
		_w15262_,
		_w15259_,
		_w15992_
	);
	LUT2 #(
		.INIT('h1)
	) name14643 (
		_w15991_,
		_w15992_,
		_w15993_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14644 (
		\P2_rEIP_reg[21]/NET0131 ,
		_w1609_,
		_w15250_,
		_w15993_,
		_w15994_
	);
	LUT3 #(
		.INIT('h48)
	) name14645 (
		\P1_rEIP_reg[21]/NET0131 ,
		_w1856_,
		_w15858_,
		_w15995_
	);
	LUT3 #(
		.INIT('hb0)
	) name14646 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[19]_pad ,
		_w15996_
	);
	LUT3 #(
		.INIT('h15)
	) name14647 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w10923_,
		_w15284_,
		_w15997_
	);
	LUT3 #(
		.INIT('h4c)
	) name14648 (
		_w10973_,
		_w15287_,
		_w15861_,
		_w15998_
	);
	LUT3 #(
		.INIT('h45)
	) name14649 (
		_w15996_,
		_w15997_,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('hb)
	) name14650 (
		_w15995_,
		_w15999_,
		_w16000_
	);
	LUT3 #(
		.INIT('h48)
	) name14651 (
		\P3_rEIP_reg[9]/NET0131 ,
		_w2110_,
		_w15220_,
		_w16001_
	);
	LUT3 #(
		.INIT('h8a)
	) name14652 (
		\P3_Address_reg[7]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16002_
	);
	LUT3 #(
		.INIT('h07)
	) name14653 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		\P3_rEIP_reg[8]/NET0131 ,
		_w16003_
	);
	LUT2 #(
		.INIT('h2)
	) name14654 (
		_w15237_,
		_w16003_,
		_w16004_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14655 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w11804_,
		_w15234_,
		_w16004_,
		_w16005_
	);
	LUT2 #(
		.INIT('h1)
	) name14656 (
		_w16002_,
		_w16005_,
		_w16006_
	);
	LUT2 #(
		.INIT('hb)
	) name14657 (
		_w16001_,
		_w16006_,
		_w16007_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14658 (
		\P2_rEIP_reg[8]/NET0131 ,
		\P2_rEIP_reg[9]/NET0131 ,
		_w1609_,
		_w15245_,
		_w16008_
	);
	LUT3 #(
		.INIT('h8a)
	) name14659 (
		\P2_Address_reg[7]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16009_
	);
	LUT4 #(
		.INIT('h9500)
	) name14660 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w9768_,
		_w9769_,
		_w15259_,
		_w16010_
	);
	LUT3 #(
		.INIT('h07)
	) name14661 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w16011_
	);
	LUT2 #(
		.INIT('h2)
	) name14662 (
		_w15262_,
		_w16011_,
		_w16012_
	);
	LUT3 #(
		.INIT('h45)
	) name14663 (
		_w16009_,
		_w16010_,
		_w16012_,
		_w16013_
	);
	LUT2 #(
		.INIT('hb)
	) name14664 (
		_w16008_,
		_w16013_,
		_w16014_
	);
	LUT3 #(
		.INIT('h48)
	) name14665 (
		\P1_rEIP_reg[9]/NET0131 ,
		_w1856_,
		_w15272_,
		_w16015_
	);
	LUT3 #(
		.INIT('hb0)
	) name14666 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[7]_pad ,
		_w16016_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14667 (
		\P1_rEIP_reg[7]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w15287_,
		_w15880_,
		_w16017_
	);
	LUT2 #(
		.INIT('h1)
	) name14668 (
		_w16016_,
		_w16017_,
		_w16018_
	);
	LUT2 #(
		.INIT('hb)
	) name14669 (
		_w16015_,
		_w16018_,
		_w16019_
	);
	LUT4 #(
		.INIT('h0040)
	) name14670 (
		\P1_D_C_n_reg/NET0131 ,
		\P1_M_IO_n_reg/NET0131 ,
		\P1_W_R_n_reg/NET0131 ,
		\ast1_pad ,
		_w16020_
	);
	LUT4 #(
		.INIT('h0001)
	) name14671 (
		\P1_BE_n_reg[0]/NET0131 ,
		\P1_BE_n_reg[1]/NET0131 ,
		\P1_BE_n_reg[2]/NET0131 ,
		\P1_BE_n_reg[3]/NET0131 ,
		_w16021_
	);
	LUT2 #(
		.INIT('h8)
	) name14672 (
		_w16020_,
		_w16021_,
		_w16022_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14673 (
		\address1[29]_pad ,
		_w3419_,
		_w3424_,
		_w16022_,
		_w16023_
	);
	LUT4 #(
		.INIT('hd5ff)
	) name14674 (
		\address1[29]_pad ,
		_w3419_,
		_w3424_,
		_w16022_,
		_w16024_
	);
	LUT4 #(
		.INIT('h1000)
	) name14675 (
		\P2_BE_n_reg[3]/NET0131 ,
		\P2_D_C_n_reg/NET0131 ,
		\P2_M_IO_n_reg/NET0131 ,
		\P2_W_R_n_reg/NET0131 ,
		_w16025_
	);
	LUT4 #(
		.INIT('h0001)
	) name14676 (
		\P2_ADS_n_reg/NET0131 ,
		\P2_BE_n_reg[0]/NET0131 ,
		\P2_BE_n_reg[1]/NET0131 ,
		\P2_BE_n_reg[2]/NET0131 ,
		_w16026_
	);
	LUT2 #(
		.INIT('h8)
	) name14677 (
		_w16025_,
		_w16026_,
		_w16027_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14678 (
		\P2_Address_reg[29]/NET0131 ,
		_w2255_,
		_w2260_,
		_w16027_,
		_w16028_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14679 (
		\P2_Datao_reg[16]/NET0131 ,
		\buf1_reg[16]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16029_
	);
	LUT2 #(
		.INIT('h8)
	) name14680 (
		\P1_Datao_reg[16]/NET0131 ,
		_w16023_,
		_w16030_
	);
	LUT2 #(
		.INIT('he)
	) name14681 (
		_w16029_,
		_w16030_,
		_w16031_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14682 (
		\P2_Datao_reg[27]/NET0131 ,
		\buf1_reg[27]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16032_
	);
	LUT2 #(
		.INIT('h8)
	) name14683 (
		\P1_Datao_reg[27]/NET0131 ,
		_w16023_,
		_w16033_
	);
	LUT2 #(
		.INIT('he)
	) name14684 (
		_w16032_,
		_w16033_,
		_w16034_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14685 (
		\P2_Datao_reg[3]/NET0131 ,
		\buf1_reg[3]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16035_
	);
	LUT2 #(
		.INIT('h8)
	) name14686 (
		\P1_Datao_reg[3]/NET0131 ,
		_w16023_,
		_w16036_
	);
	LUT2 #(
		.INIT('he)
	) name14687 (
		_w16035_,
		_w16036_,
		_w16037_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14688 (
		\P2_Datao_reg[14]/NET0131 ,
		\buf1_reg[14]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16038_
	);
	LUT2 #(
		.INIT('h8)
	) name14689 (
		\P1_Datao_reg[14]/NET0131 ,
		_w16023_,
		_w16039_
	);
	LUT2 #(
		.INIT('he)
	) name14690 (
		_w16038_,
		_w16039_,
		_w16040_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14691 (
		\P2_Datao_reg[30]/NET0131 ,
		\buf1_reg[30]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16041_
	);
	LUT2 #(
		.INIT('h8)
	) name14692 (
		\P1_Datao_reg[30]/NET0131 ,
		_w16023_,
		_w16042_
	);
	LUT2 #(
		.INIT('he)
	) name14693 (
		_w16041_,
		_w16042_,
		_w16043_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14694 (
		\P2_Datao_reg[25]/NET0131 ,
		\buf1_reg[25]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16044_
	);
	LUT2 #(
		.INIT('h8)
	) name14695 (
		\P1_Datao_reg[25]/NET0131 ,
		_w16023_,
		_w16045_
	);
	LUT2 #(
		.INIT('he)
	) name14696 (
		_w16044_,
		_w16045_,
		_w16046_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14697 (
		\P2_Datao_reg[26]/NET0131 ,
		\buf1_reg[26]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16047_
	);
	LUT2 #(
		.INIT('h8)
	) name14698 (
		\P1_Datao_reg[26]/NET0131 ,
		_w16023_,
		_w16048_
	);
	LUT2 #(
		.INIT('he)
	) name14699 (
		_w16047_,
		_w16048_,
		_w16049_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14700 (
		\P2_Datao_reg[15]/NET0131 ,
		\buf1_reg[15]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16050_
	);
	LUT2 #(
		.INIT('h8)
	) name14701 (
		\P1_Datao_reg[15]/NET0131 ,
		_w16023_,
		_w16051_
	);
	LUT2 #(
		.INIT('he)
	) name14702 (
		_w16050_,
		_w16051_,
		_w16052_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14703 (
		\P2_Datao_reg[19]/NET0131 ,
		\buf1_reg[19]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16053_
	);
	LUT2 #(
		.INIT('h8)
	) name14704 (
		\P1_Datao_reg[19]/NET0131 ,
		_w16023_,
		_w16054_
	);
	LUT2 #(
		.INIT('he)
	) name14705 (
		_w16053_,
		_w16054_,
		_w16055_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14706 (
		\P2_Datao_reg[0]/NET0131 ,
		\buf1_reg[0]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16056_
	);
	LUT2 #(
		.INIT('h8)
	) name14707 (
		\P1_Datao_reg[0]/NET0131 ,
		_w16023_,
		_w16057_
	);
	LUT2 #(
		.INIT('he)
	) name14708 (
		_w16056_,
		_w16057_,
		_w16058_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14709 (
		\P2_Datao_reg[10]/NET0131 ,
		\buf1_reg[10]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16059_
	);
	LUT2 #(
		.INIT('h8)
	) name14710 (
		\P1_Datao_reg[10]/NET0131 ,
		_w16023_,
		_w16060_
	);
	LUT2 #(
		.INIT('he)
	) name14711 (
		_w16059_,
		_w16060_,
		_w16061_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14712 (
		\P2_Datao_reg[11]/NET0131 ,
		\buf1_reg[11]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16062_
	);
	LUT2 #(
		.INIT('h8)
	) name14713 (
		\P1_Datao_reg[11]/NET0131 ,
		_w16023_,
		_w16063_
	);
	LUT2 #(
		.INIT('he)
	) name14714 (
		_w16062_,
		_w16063_,
		_w16064_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14715 (
		\P2_Datao_reg[12]/NET0131 ,
		\buf1_reg[12]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16065_
	);
	LUT2 #(
		.INIT('h8)
	) name14716 (
		\P1_Datao_reg[12]/NET0131 ,
		_w16023_,
		_w16066_
	);
	LUT2 #(
		.INIT('he)
	) name14717 (
		_w16065_,
		_w16066_,
		_w16067_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14718 (
		\P2_Datao_reg[13]/NET0131 ,
		\buf1_reg[13]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16068_
	);
	LUT2 #(
		.INIT('h8)
	) name14719 (
		\P1_Datao_reg[13]/NET0131 ,
		_w16023_,
		_w16069_
	);
	LUT2 #(
		.INIT('he)
	) name14720 (
		_w16068_,
		_w16069_,
		_w16070_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14721 (
		\P2_Datao_reg[17]/NET0131 ,
		\buf1_reg[17]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16071_
	);
	LUT2 #(
		.INIT('h8)
	) name14722 (
		\P1_Datao_reg[17]/NET0131 ,
		_w16023_,
		_w16072_
	);
	LUT2 #(
		.INIT('he)
	) name14723 (
		_w16071_,
		_w16072_,
		_w16073_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14724 (
		\P2_Datao_reg[1]/NET0131 ,
		\buf1_reg[1]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16074_
	);
	LUT2 #(
		.INIT('h8)
	) name14725 (
		\P1_Datao_reg[1]/NET0131 ,
		_w16023_,
		_w16075_
	);
	LUT2 #(
		.INIT('he)
	) name14726 (
		_w16074_,
		_w16075_,
		_w16076_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14727 (
		\P2_Datao_reg[20]/NET0131 ,
		\buf1_reg[20]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16077_
	);
	LUT2 #(
		.INIT('h8)
	) name14728 (
		\P1_Datao_reg[20]/NET0131 ,
		_w16023_,
		_w16078_
	);
	LUT2 #(
		.INIT('he)
	) name14729 (
		_w16077_,
		_w16078_,
		_w16079_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14730 (
		\P2_Datao_reg[21]/NET0131 ,
		\buf1_reg[21]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16080_
	);
	LUT2 #(
		.INIT('h8)
	) name14731 (
		\P1_Datao_reg[21]/NET0131 ,
		_w16023_,
		_w16081_
	);
	LUT2 #(
		.INIT('he)
	) name14732 (
		_w16080_,
		_w16081_,
		_w16082_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14733 (
		\P2_Datao_reg[22]/NET0131 ,
		\buf1_reg[22]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16083_
	);
	LUT2 #(
		.INIT('h8)
	) name14734 (
		\P1_Datao_reg[22]/NET0131 ,
		_w16023_,
		_w16084_
	);
	LUT2 #(
		.INIT('he)
	) name14735 (
		_w16083_,
		_w16084_,
		_w16085_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14736 (
		\P2_Datao_reg[23]/NET0131 ,
		\buf1_reg[23]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16086_
	);
	LUT2 #(
		.INIT('h8)
	) name14737 (
		\P1_Datao_reg[23]/NET0131 ,
		_w16023_,
		_w16087_
	);
	LUT2 #(
		.INIT('he)
	) name14738 (
		_w16086_,
		_w16087_,
		_w16088_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14739 (
		\P2_Datao_reg[24]/NET0131 ,
		\buf1_reg[24]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16089_
	);
	LUT2 #(
		.INIT('h8)
	) name14740 (
		\P1_Datao_reg[24]/NET0131 ,
		_w16023_,
		_w16090_
	);
	LUT2 #(
		.INIT('he)
	) name14741 (
		_w16089_,
		_w16090_,
		_w16091_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14742 (
		\P2_Datao_reg[28]/NET0131 ,
		\buf1_reg[28]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16092_
	);
	LUT2 #(
		.INIT('h8)
	) name14743 (
		\P1_Datao_reg[28]/NET0131 ,
		_w16023_,
		_w16093_
	);
	LUT2 #(
		.INIT('he)
	) name14744 (
		_w16092_,
		_w16093_,
		_w16094_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14745 (
		\P2_Datao_reg[2]/NET0131 ,
		\buf1_reg[2]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16095_
	);
	LUT2 #(
		.INIT('h8)
	) name14746 (
		\P1_Datao_reg[2]/NET0131 ,
		_w16023_,
		_w16096_
	);
	LUT2 #(
		.INIT('he)
	) name14747 (
		_w16095_,
		_w16096_,
		_w16097_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14748 (
		\P2_Datao_reg[4]/NET0131 ,
		\buf1_reg[4]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16098_
	);
	LUT2 #(
		.INIT('h8)
	) name14749 (
		\P1_Datao_reg[4]/NET0131 ,
		_w16023_,
		_w16099_
	);
	LUT2 #(
		.INIT('he)
	) name14750 (
		_w16098_,
		_w16099_,
		_w16100_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14751 (
		\P2_Datao_reg[6]/NET0131 ,
		\buf1_reg[6]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16101_
	);
	LUT2 #(
		.INIT('h8)
	) name14752 (
		\P1_Datao_reg[6]/NET0131 ,
		_w16023_,
		_w16102_
	);
	LUT2 #(
		.INIT('he)
	) name14753 (
		_w16101_,
		_w16102_,
		_w16103_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14754 (
		\P2_Datao_reg[9]/NET0131 ,
		\buf1_reg[9]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16104_
	);
	LUT2 #(
		.INIT('h8)
	) name14755 (
		\P1_Datao_reg[9]/NET0131 ,
		_w16023_,
		_w16105_
	);
	LUT2 #(
		.INIT('he)
	) name14756 (
		_w16104_,
		_w16105_,
		_w16106_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14757 (
		\P2_Datao_reg[29]/NET0131 ,
		\buf1_reg[29]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16107_
	);
	LUT2 #(
		.INIT('h8)
	) name14758 (
		\P1_Datao_reg[29]/NET0131 ,
		_w16023_,
		_w16108_
	);
	LUT2 #(
		.INIT('he)
	) name14759 (
		_w16107_,
		_w16108_,
		_w16109_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14760 (
		\P2_Datao_reg[18]/NET0131 ,
		\buf1_reg[18]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16110_
	);
	LUT2 #(
		.INIT('h8)
	) name14761 (
		\P1_Datao_reg[18]/NET0131 ,
		_w16023_,
		_w16111_
	);
	LUT2 #(
		.INIT('he)
	) name14762 (
		_w16110_,
		_w16111_,
		_w16112_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14763 (
		\P2_Datao_reg[7]/NET0131 ,
		\buf1_reg[7]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16113_
	);
	LUT2 #(
		.INIT('h8)
	) name14764 (
		\P1_Datao_reg[7]/NET0131 ,
		_w16023_,
		_w16114_
	);
	LUT2 #(
		.INIT('he)
	) name14765 (
		_w16113_,
		_w16114_,
		_w16115_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14766 (
		\P2_Datao_reg[8]/NET0131 ,
		\buf1_reg[8]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16116_
	);
	LUT2 #(
		.INIT('h8)
	) name14767 (
		\P1_Datao_reg[8]/NET0131 ,
		_w16023_,
		_w16117_
	);
	LUT2 #(
		.INIT('he)
	) name14768 (
		_w16116_,
		_w16117_,
		_w16118_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name14769 (
		\P2_Datao_reg[5]/NET0131 ,
		\buf1_reg[5]/NET0131 ,
		_w16023_,
		_w16028_,
		_w16119_
	);
	LUT2 #(
		.INIT('h8)
	) name14770 (
		\P1_Datao_reg[5]/NET0131 ,
		_w16023_,
		_w16120_
	);
	LUT2 #(
		.INIT('he)
	) name14771 (
		_w16119_,
		_w16120_,
		_w16121_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14772 (
		\P3_rEIP_reg[15]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w2110_,
		_w15224_,
		_w16122_
	);
	LUT3 #(
		.INIT('h8a)
	) name14773 (
		\P3_Address_reg[14]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16123_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14774 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w15237_,
		_w15459_,
		_w16123_,
		_w16124_
	);
	LUT2 #(
		.INIT('hb)
	) name14775 (
		_w16122_,
		_w16124_,
		_w16125_
	);
	LUT4 #(
		.INIT('h070f)
	) name14776 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w15724_,
		_w16126_
	);
	LUT2 #(
		.INIT('h2)
	) name14777 (
		_w1609_,
		_w15924_,
		_w16127_
	);
	LUT3 #(
		.INIT('h8a)
	) name14778 (
		\P2_Address_reg[14]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16128_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14779 (
		\P2_rEIP_reg[15]/NET0131 ,
		_w9773_,
		_w15262_,
		_w15726_,
		_w16129_
	);
	LUT2 #(
		.INIT('h1)
	) name14780 (
		_w16128_,
		_w16129_,
		_w16130_
	);
	LUT3 #(
		.INIT('h4f)
	) name14781 (
		_w16126_,
		_w16127_,
		_w16130_,
		_w16131_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14782 (
		\P1_rEIP_reg[15]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w1856_,
		_w15276_,
		_w16132_
	);
	LUT3 #(
		.INIT('hb0)
	) name14783 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[14]_pad ,
		_w16133_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14784 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w15287_,
		_w15911_,
		_w16133_,
		_w16134_
	);
	LUT2 #(
		.INIT('hb)
	) name14785 (
		_w16132_,
		_w16134_,
		_w16135_
	);
	LUT3 #(
		.INIT('h48)
	) name14786 (
		\P1_rEIP_reg[28]/NET0131 ,
		_w1856_,
		_w15280_,
		_w16136_
	);
	LUT3 #(
		.INIT('hb0)
	) name14787 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[26]_pad ,
		_w16137_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14788 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w11159_,
		_w15284_,
		_w15287_,
		_w16138_
	);
	LUT2 #(
		.INIT('h1)
	) name14789 (
		_w16137_,
		_w16138_,
		_w16139_
	);
	LUT2 #(
		.INIT('hb)
	) name14790 (
		_w16136_,
		_w16139_,
		_w16140_
	);
	LUT3 #(
		.INIT('h13)
	) name14791 (
		\P3_rEIP_reg[27]/NET0131 ,
		\P3_rEIP_reg[28]/NET0131 ,
		_w15701_,
		_w16141_
	);
	LUT2 #(
		.INIT('h2)
	) name14792 (
		_w2110_,
		_w15230_,
		_w16142_
	);
	LUT3 #(
		.INIT('h8a)
	) name14793 (
		\P3_Address_reg[26]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16143_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14794 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w15237_,
		_w15919_,
		_w16143_,
		_w16144_
	);
	LUT3 #(
		.INIT('h4f)
	) name14795 (
		_w16141_,
		_w16142_,
		_w16144_,
		_w16145_
	);
	LUT3 #(
		.INIT('h8a)
	) name14796 (
		\P2_Address_reg[26]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16146_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14797 (
		\P2_rEIP_reg[27]/NET0131 ,
		_w15262_,
		_w15260_,
		_w16146_,
		_w16147_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14798 (
		\P2_rEIP_reg[28]/NET0131 ,
		_w1609_,
		_w15255_,
		_w16147_,
		_w16148_
	);
	LUT3 #(
		.INIT('h8a)
	) name14799 (
		\P3_Address_reg[22]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16149_
	);
	LUT4 #(
		.INIT('h009f)
	) name14800 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w15235_,
		_w15237_,
		_w16149_,
		_w16150_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14801 (
		\P3_rEIP_reg[24]/NET0131 ,
		_w2110_,
		_w15228_,
		_w16150_,
		_w16151_
	);
	LUT3 #(
		.INIT('h8a)
	) name14802 (
		\P2_Address_reg[22]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16152_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14803 (
		\P2_rEIP_reg[23]/NET0131 ,
		_w9780_,
		_w15262_,
		_w15259_,
		_w16153_
	);
	LUT2 #(
		.INIT('h1)
	) name14804 (
		_w16152_,
		_w16153_,
		_w16154_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14805 (
		\P2_rEIP_reg[24]/NET0131 ,
		_w1609_,
		_w15252_,
		_w16154_,
		_w16155_
	);
	LUT4 #(
		.INIT('h4888)
	) name14806 (
		\P1_rEIP_reg[24]/NET0131 ,
		_w1856_,
		_w11024_,
		_w15858_,
		_w16156_
	);
	LUT3 #(
		.INIT('hb0)
	) name14807 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[22]_pad ,
		_w16157_
	);
	LUT4 #(
		.INIT('h8000)
	) name14808 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w10973_,
		_w15861_,
		_w16158_
	);
	LUT4 #(
		.INIT('h70f0)
	) name14809 (
		_w10973_,
		_w11024_,
		_w15287_,
		_w15861_,
		_w16159_
	);
	LUT4 #(
		.INIT('h0133)
	) name14810 (
		\P1_rEIP_reg[23]/NET0131 ,
		_w16157_,
		_w16158_,
		_w16159_,
		_w16160_
	);
	LUT2 #(
		.INIT('hb)
	) name14811 (
		_w16156_,
		_w16160_,
		_w16161_
	);
	LUT3 #(
		.INIT('h48)
	) name14812 (
		\P3_rEIP_reg[12]/NET0131 ,
		_w2110_,
		_w15222_,
		_w16162_
	);
	LUT3 #(
		.INIT('h8a)
	) name14813 (
		\P3_Address_reg[10]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16163_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14814 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w11806_,
		_w15234_,
		_w15237_,
		_w16164_
	);
	LUT2 #(
		.INIT('h1)
	) name14815 (
		_w16163_,
		_w16164_,
		_w16165_
	);
	LUT2 #(
		.INIT('hb)
	) name14816 (
		_w16162_,
		_w16165_,
		_w16166_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14817 (
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[12]/NET0131 ,
		_w1609_,
		_w15247_,
		_w16167_
	);
	LUT3 #(
		.INIT('h8a)
	) name14818 (
		\P2_Address_reg[10]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16168_
	);
	LUT4 #(
		.INIT('h9300)
	) name14819 (
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		_w9770_,
		_w15259_,
		_w16169_
	);
	LUT3 #(
		.INIT('h13)
	) name14820 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[11]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16170_
	);
	LUT2 #(
		.INIT('h2)
	) name14821 (
		_w15262_,
		_w16170_,
		_w16171_
	);
	LUT3 #(
		.INIT('h45)
	) name14822 (
		_w16168_,
		_w16169_,
		_w16171_,
		_w16172_
	);
	LUT2 #(
		.INIT('hb)
	) name14823 (
		_w16167_,
		_w16172_,
		_w16173_
	);
	LUT3 #(
		.INIT('h48)
	) name14824 (
		\P1_rEIP_reg[12]/NET0131 ,
		_w1856_,
		_w15274_,
		_w16174_
	);
	LUT3 #(
		.INIT('hb0)
	) name14825 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[10]_pad ,
		_w16175_
	);
	LUT3 #(
		.INIT('h13)
	) name14826 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w16176_
	);
	LUT2 #(
		.INIT('h2)
	) name14827 (
		_w15287_,
		_w16176_,
		_w16177_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14828 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w10812_,
		_w15284_,
		_w16177_,
		_w16178_
	);
	LUT2 #(
		.INIT('h1)
	) name14829 (
		_w16175_,
		_w16178_,
		_w16179_
	);
	LUT2 #(
		.INIT('hb)
	) name14830 (
		_w16174_,
		_w16179_,
		_w16180_
	);
	LUT2 #(
		.INIT('hb)
	) name14831 (
		_w16023_,
		_w16028_,
		_w16181_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14832 (
		\P3_rEIP_reg[3]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w2110_,
		_w15216_,
		_w16182_
	);
	LUT3 #(
		.INIT('h8a)
	) name14833 (
		\P3_Address_reg[2]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16183_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14834 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w15237_,
		_w15887_,
		_w16183_,
		_w16184_
	);
	LUT2 #(
		.INIT('hb)
	) name14835 (
		_w16182_,
		_w16184_,
		_w16185_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14836 (
		\P2_rEIP_reg[3]/NET0131 ,
		\P2_rEIP_reg[4]/NET0131 ,
		_w1609_,
		_w15243_,
		_w16186_
	);
	LUT3 #(
		.INIT('h8a)
	) name14837 (
		\P2_Address_reg[2]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16187_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14838 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w15262_,
		_w15897_,
		_w16187_,
		_w16188_
	);
	LUT2 #(
		.INIT('hb)
	) name14839 (
		_w16186_,
		_w16188_,
		_w16189_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14840 (
		\P1_rEIP_reg[3]/NET0131 ,
		\P1_rEIP_reg[4]/NET0131 ,
		_w1856_,
		_w15268_,
		_w16190_
	);
	LUT3 #(
		.INIT('hb0)
	) name14841 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[2]_pad ,
		_w16191_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14842 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w15287_,
		_w15905_,
		_w16191_,
		_w16192_
	);
	LUT2 #(
		.INIT('hb)
	) name14843 (
		_w16190_,
		_w16192_,
		_w16193_
	);
	LUT4 #(
		.INIT('h1555)
	) name14844 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w11923_,
		_w11970_,
		_w15234_,
		_w16194_
	);
	LUT3 #(
		.INIT('h02)
	) name14845 (
		_w15237_,
		_w15987_,
		_w16194_,
		_w16195_
	);
	LUT3 #(
		.INIT('h8a)
	) name14846 (
		\P3_Address_reg[18]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16196_
	);
	LUT4 #(
		.INIT('h4888)
	) name14847 (
		\P3_rEIP_reg[20]/NET0131 ,
		_w2110_,
		_w12025_,
		_w15225_,
		_w16197_
	);
	LUT3 #(
		.INIT('hfe)
	) name14848 (
		_w16196_,
		_w16197_,
		_w16195_,
		_w16198_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14849 (
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w1609_,
		_w15249_,
		_w16199_
	);
	LUT3 #(
		.INIT('h8a)
	) name14850 (
		\P2_Address_reg[18]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16200_
	);
	LUT3 #(
		.INIT('h13)
	) name14851 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16201_
	);
	LUT2 #(
		.INIT('h2)
	) name14852 (
		_w15262_,
		_w16201_,
		_w16202_
	);
	LUT4 #(
		.INIT('h040f)
	) name14853 (
		_w11316_,
		_w15259_,
		_w16200_,
		_w16202_,
		_w16203_
	);
	LUT2 #(
		.INIT('hb)
	) name14854 (
		_w16199_,
		_w16203_,
		_w16204_
	);
	LUT3 #(
		.INIT('h48)
	) name14855 (
		\P1_rEIP_reg[20]/NET0131 ,
		_w1856_,
		_w15857_,
		_w16205_
	);
	LUT3 #(
		.INIT('hb0)
	) name14856 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[18]_pad ,
		_w16206_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14857 (
		\P1_rEIP_reg[19]/NET0131 ,
		_w10908_,
		_w15284_,
		_w15287_,
		_w16207_
	);
	LUT2 #(
		.INIT('h1)
	) name14858 (
		_w16206_,
		_w16207_,
		_w16208_
	);
	LUT2 #(
		.INIT('hb)
	) name14859 (
		_w16205_,
		_w16208_,
		_w16209_
	);
	LUT3 #(
		.INIT('h8a)
	) name14860 (
		\P3_Address_reg[6]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16210_
	);
	LUT4 #(
		.INIT('h8000)
	) name14861 (
		\P3_rEIP_reg[5]/NET0131 ,
		\P3_rEIP_reg[6]/NET0131 ,
		_w11803_,
		_w15234_,
		_w16211_
	);
	LUT4 #(
		.INIT('h0b07)
	) name14862 (
		\P3_rEIP_reg[7]/NET0131 ,
		_w15237_,
		_w16210_,
		_w16211_,
		_w16212_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14863 (
		\P3_rEIP_reg[8]/NET0131 ,
		_w2110_,
		_w15219_,
		_w16212_,
		_w16213_
	);
	LUT3 #(
		.INIT('h48)
	) name14864 (
		\P2_rEIP_reg[8]/NET0131 ,
		_w1609_,
		_w15245_,
		_w16214_
	);
	LUT3 #(
		.INIT('h8a)
	) name14865 (
		\P2_Address_reg[6]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16215_
	);
	LUT3 #(
		.INIT('h07)
	) name14866 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w16216_
	);
	LUT2 #(
		.INIT('h2)
	) name14867 (
		_w15262_,
		_w16216_,
		_w16217_
	);
	LUT4 #(
		.INIT('h040f)
	) name14868 (
		_w11730_,
		_w15259_,
		_w16215_,
		_w16217_,
		_w16218_
	);
	LUT2 #(
		.INIT('hb)
	) name14869 (
		_w16214_,
		_w16218_,
		_w16219_
	);
	LUT3 #(
		.INIT('hb0)
	) name14870 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[6]_pad ,
		_w16220_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14871 (
		\P1_rEIP_reg[7]/NET0131 ,
		_w15287_,
		_w15880_,
		_w16220_,
		_w16221_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14872 (
		\P1_rEIP_reg[8]/NET0131 ,
		_w1856_,
		_w15271_,
		_w16221_,
		_w16222_
	);
	LUT3 #(
		.INIT('h8a)
	) name14873 (
		\P3_Address_reg[25]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16223_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14874 (
		\P3_rEIP_reg[26]/NET0131 ,
		_w12119_,
		_w15235_,
		_w15237_,
		_w16224_
	);
	LUT2 #(
		.INIT('h1)
	) name14875 (
		_w16223_,
		_w16224_,
		_w16225_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14876 (
		\P3_rEIP_reg[27]/NET0131 ,
		_w2110_,
		_w15701_,
		_w16225_,
		_w16226_
	);
	LUT3 #(
		.INIT('h8a)
	) name14877 (
		\P2_Address_reg[25]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16227_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14878 (
		\P2_rEIP_reg[26]/NET0131 ,
		_w9782_,
		_w15262_,
		_w15259_,
		_w16228_
	);
	LUT2 #(
		.INIT('h1)
	) name14879 (
		_w16227_,
		_w16228_,
		_w16229_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14880 (
		\P2_rEIP_reg[27]/NET0131 ,
		_w1609_,
		_w15254_,
		_w16229_,
		_w16230_
	);
	LUT3 #(
		.INIT('h48)
	) name14881 (
		\P1_rEIP_reg[27]/NET0131 ,
		_w1856_,
		_w15279_,
		_w16231_
	);
	LUT3 #(
		.INIT('hb0)
	) name14882 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[25]_pad ,
		_w16232_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14883 (
		\P1_rEIP_reg[26]/NET0131 ,
		_w11108_,
		_w15284_,
		_w15287_,
		_w16233_
	);
	LUT2 #(
		.INIT('h1)
	) name14884 (
		_w16232_,
		_w16233_,
		_w16234_
	);
	LUT2 #(
		.INIT('hb)
	) name14885 (
		_w16231_,
		_w16234_,
		_w16235_
	);
	LUT3 #(
		.INIT('h8a)
	) name14886 (
		\P3_Address_reg[29]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16236_
	);
	LUT4 #(
		.INIT('h9500)
	) name14887 (
		\P3_rEIP_reg[30]/NET0131 ,
		_w12120_,
		_w12193_,
		_w15234_,
		_w16237_
	);
	LUT3 #(
		.INIT('h13)
	) name14888 (
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w16238_
	);
	LUT2 #(
		.INIT('h2)
	) name14889 (
		_w15237_,
		_w16238_,
		_w16239_
	);
	LUT3 #(
		.INIT('h45)
	) name14890 (
		_w16236_,
		_w16237_,
		_w16239_,
		_w16240_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14891 (
		\P3_rEIP_reg[31]/NET0131 ,
		_w2110_,
		_w15231_,
		_w16240_,
		_w16241_
	);
	LUT3 #(
		.INIT('h8a)
	) name14892 (
		\P2_Address_reg[29]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16242_
	);
	LUT4 #(
		.INIT('h9300)
	) name14893 (
		\P2_rEIP_reg[29]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w9784_,
		_w15259_,
		_w16243_
	);
	LUT3 #(
		.INIT('h13)
	) name14894 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16244_
	);
	LUT2 #(
		.INIT('h2)
	) name14895 (
		_w15262_,
		_w16244_,
		_w16245_
	);
	LUT3 #(
		.INIT('h45)
	) name14896 (
		_w16242_,
		_w16243_,
		_w16245_,
		_w16246_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14897 (
		\P2_rEIP_reg[31]/NET0131 ,
		_w1609_,
		_w15257_,
		_w16246_,
		_w16247_
	);
	LUT3 #(
		.INIT('h48)
	) name14898 (
		\P1_rEIP_reg[31]/NET0131 ,
		_w1856_,
		_w15282_,
		_w16248_
	);
	LUT3 #(
		.INIT('hb0)
	) name14899 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[29]_pad ,
		_w16249_
	);
	LUT4 #(
		.INIT('h6c00)
	) name14900 (
		\P1_rEIP_reg[29]/NET0131 ,
		\P1_rEIP_reg[30]/NET0131 ,
		_w15286_,
		_w15287_,
		_w16250_
	);
	LUT2 #(
		.INIT('h1)
	) name14901 (
		_w16249_,
		_w16250_,
		_w16251_
	);
	LUT2 #(
		.INIT('hb)
	) name14902 (
		_w16248_,
		_w16251_,
		_w16252_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name14903 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		hold_pad,
		_w16253_
	);
	LUT3 #(
		.INIT('h80)
	) name14904 (
		\P2_State_reg[1]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16254_
	);
	LUT2 #(
		.INIT('h2)
	) name14905 (
		\P2_RequestPending_reg/NET0131 ,
		hold_pad,
		_w16255_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14906 (
		\P2_State_reg[0]/NET0131 ,
		_w16254_,
		_w16253_,
		_w16255_,
		_w16256_
	);
	LUT4 #(
		.INIT('h8000)
	) name14907 (
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16257_
	);
	LUT2 #(
		.INIT('h2)
	) name14908 (
		_w1611_,
		_w16257_,
		_w16258_
	);
	LUT2 #(
		.INIT('hb)
	) name14909 (
		_w16256_,
		_w16258_,
		_w16259_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name14910 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		hold_pad,
		_w16260_
	);
	LUT3 #(
		.INIT('h80)
	) name14911 (
		\P3_State_reg[1]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16261_
	);
	LUT2 #(
		.INIT('h2)
	) name14912 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		_w16262_
	);
	LUT4 #(
		.INIT('haaa8)
	) name14913 (
		\P3_State_reg[0]/NET0131 ,
		_w16261_,
		_w16260_,
		_w16262_,
		_w16263_
	);
	LUT4 #(
		.INIT('h8000)
	) name14914 (
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16264_
	);
	LUT2 #(
		.INIT('h2)
	) name14915 (
		_w2111_,
		_w16264_,
		_w16265_
	);
	LUT2 #(
		.INIT('hb)
	) name14916 (
		_w16263_,
		_w16265_,
		_w16266_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name14917 (
		\P1_State_reg[2]/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16267_
	);
	LUT3 #(
		.INIT('hc8)
	) name14918 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16268_
	);
	LUT4 #(
		.INIT('h0888)
	) name14919 (
		\P1_RequestPending_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		hold_pad,
		_w16269_
	);
	LUT4 #(
		.INIT('hdfdd)
	) name14920 (
		_w1858_,
		_w16269_,
		_w16267_,
		_w16268_,
		_w16270_
	);
	LUT3 #(
		.INIT('h2a)
	) name14921 (
		\P2_State_reg[0]/NET0131 ,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16271_
	);
	LUT3 #(
		.INIT('h8c)
	) name14922 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		na_pad,
		_w16272_
	);
	LUT3 #(
		.INIT('h02)
	) name14923 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16273_
	);
	LUT4 #(
		.INIT('h00ab)
	) name14924 (
		hold_pad,
		_w16271_,
		_w16272_,
		_w16273_,
		_w16274_
	);
	LUT3 #(
		.INIT('h31)
	) name14925 (
		\P2_RequestPending_reg/NET0131 ,
		_w15262_,
		_w16274_,
		_w16275_
	);
	LUT4 #(
		.INIT('hcc04)
	) name14926 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16276_
	);
	LUT2 #(
		.INIT('h4)
	) name14927 (
		_w16262_,
		_w16276_,
		_w16277_
	);
	LUT4 #(
		.INIT('h0222)
	) name14928 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16278_
	);
	LUT3 #(
		.INIT('ha2)
	) name14929 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16278_,
		_w16279_
	);
	LUT4 #(
		.INIT('h3331)
	) name14930 (
		\P3_RequestPending_reg/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		hold_pad,
		na_pad,
		_w16280_
	);
	LUT2 #(
		.INIT('h2)
	) name14931 (
		\P3_State_reg[2]/NET0131 ,
		_w16280_,
		_w16281_
	);
	LUT3 #(
		.INIT('hab)
	) name14932 (
		_w16277_,
		_w16279_,
		_w16281_,
		_w16282_
	);
	LUT3 #(
		.INIT('h02)
	) name14933 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16283_
	);
	LUT3 #(
		.INIT('h2a)
	) name14934 (
		\P1_State_reg[0]/NET0131 ,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16284_
	);
	LUT3 #(
		.INIT('h8c)
	) name14935 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		na_pad,
		_w16285_
	);
	LUT4 #(
		.INIT('h2223)
	) name14936 (
		hold_pad,
		_w16283_,
		_w16284_,
		_w16285_,
		_w16286_
	);
	LUT3 #(
		.INIT('h31)
	) name14937 (
		\P1_RequestPending_reg/NET0131 ,
		_w15287_,
		_w16286_,
		_w16287_
	);
	LUT3 #(
		.INIT('h48)
	) name14938 (
		\P3_rEIP_reg[15]/NET0131 ,
		_w2110_,
		_w15224_,
		_w16288_
	);
	LUT3 #(
		.INIT('h8a)
	) name14939 (
		\P3_Address_reg[13]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16289_
	);
	LUT3 #(
		.INIT('h13)
	) name14940 (
		\P3_rEIP_reg[13]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w15721_,
		_w16290_
	);
	LUT4 #(
		.INIT('h7f00)
	) name14941 (
		\P3_rEIP_reg[14]/NET0131 ,
		_w11871_,
		_w15234_,
		_w15237_,
		_w16291_
	);
	LUT3 #(
		.INIT('h45)
	) name14942 (
		_w16289_,
		_w16290_,
		_w16291_,
		_w16292_
	);
	LUT2 #(
		.INIT('hb)
	) name14943 (
		_w16288_,
		_w16292_,
		_w16293_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14944 (
		\P2_rEIP_reg[14]/NET0131 ,
		\P2_rEIP_reg[15]/NET0131 ,
		_w1609_,
		_w15724_,
		_w16294_
	);
	LUT3 #(
		.INIT('h8a)
	) name14945 (
		\P2_Address_reg[13]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16295_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14946 (
		\P2_rEIP_reg[13]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w15262_,
		_w15726_,
		_w16296_
	);
	LUT2 #(
		.INIT('h1)
	) name14947 (
		_w16295_,
		_w16296_,
		_w16297_
	);
	LUT2 #(
		.INIT('hb)
	) name14948 (
		_w16294_,
		_w16297_,
		_w16298_
	);
	LUT3 #(
		.INIT('h48)
	) name14949 (
		\P1_rEIP_reg[15]/NET0131 ,
		_w1856_,
		_w15276_,
		_w16299_
	);
	LUT3 #(
		.INIT('hb0)
	) name14950 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[13]_pad ,
		_w16300_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14951 (
		\P1_rEIP_reg[14]/NET0131 ,
		_w10814_,
		_w15284_,
		_w15287_,
		_w16301_
	);
	LUT2 #(
		.INIT('h1)
	) name14952 (
		_w16300_,
		_w16301_,
		_w16302_
	);
	LUT2 #(
		.INIT('hb)
	) name14953 (
		_w16299_,
		_w16302_,
		_w16303_
	);
	LUT3 #(
		.INIT('h48)
	) name14954 (
		\P2_rEIP_reg[11]/NET0131 ,
		_w1609_,
		_w15247_,
		_w16304_
	);
	LUT3 #(
		.INIT('h8a)
	) name14955 (
		\P2_Address_reg[9]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16305_
	);
	LUT3 #(
		.INIT('h13)
	) name14956 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[10]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16306_
	);
	LUT2 #(
		.INIT('h2)
	) name14957 (
		_w15262_,
		_w16306_,
		_w16307_
	);
	LUT4 #(
		.INIT('h6f00)
	) name14958 (
		\P2_rEIP_reg[10]/NET0131 ,
		_w9770_,
		_w15259_,
		_w16307_,
		_w16308_
	);
	LUT2 #(
		.INIT('h1)
	) name14959 (
		_w16305_,
		_w16308_,
		_w16309_
	);
	LUT2 #(
		.INIT('hb)
	) name14960 (
		_w16304_,
		_w16309_,
		_w16310_
	);
	LUT3 #(
		.INIT('h48)
	) name14961 (
		\P3_rEIP_reg[11]/NET0131 ,
		_w2110_,
		_w15221_,
		_w16311_
	);
	LUT3 #(
		.INIT('h8a)
	) name14962 (
		\P3_Address_reg[9]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16312_
	);
	LUT4 #(
		.INIT('h6a00)
	) name14963 (
		\P3_rEIP_reg[10]/NET0131 ,
		_w11805_,
		_w15234_,
		_w15237_,
		_w16313_
	);
	LUT2 #(
		.INIT('h1)
	) name14964 (
		_w16312_,
		_w16313_,
		_w16314_
	);
	LUT2 #(
		.INIT('hb)
	) name14965 (
		_w16311_,
		_w16314_,
		_w16315_
	);
	LUT3 #(
		.INIT('hb0)
	) name14966 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[9]_pad ,
		_w16316_
	);
	LUT3 #(
		.INIT('h13)
	) name14967 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[10]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w16317_
	);
	LUT2 #(
		.INIT('h2)
	) name14968 (
		_w15287_,
		_w16317_,
		_w16318_
	);
	LUT4 #(
		.INIT('h040f)
	) name14969 (
		_w12370_,
		_w15284_,
		_w16316_,
		_w16318_,
		_w16319_
	);
	LUT4 #(
		.INIT('h48ff)
	) name14970 (
		\P1_rEIP_reg[11]/NET0131 ,
		_w1856_,
		_w15273_,
		_w16319_,
		_w16320_
	);
	LUT3 #(
		.INIT('h48)
	) name14971 (
		\P3_rEIP_reg[23]/NET0131 ,
		_w2110_,
		_w15227_,
		_w16321_
	);
	LUT3 #(
		.INIT('h8a)
	) name14972 (
		\P3_Address_reg[21]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16322_
	);
	LUT4 #(
		.INIT('h3020)
	) name14973 (
		\P3_rEIP_reg[22]/NET0131 ,
		_w15235_,
		_w15237_,
		_w15849_,
		_w16323_
	);
	LUT2 #(
		.INIT('h1)
	) name14974 (
		_w16322_,
		_w16323_,
		_w16324_
	);
	LUT2 #(
		.INIT('hb)
	) name14975 (
		_w16321_,
		_w16324_,
		_w16325_
	);
	LUT4 #(
		.INIT('h60c0)
	) name14976 (
		\P2_rEIP_reg[22]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w1609_,
		_w15251_,
		_w16326_
	);
	LUT3 #(
		.INIT('h8a)
	) name14977 (
		\P2_Address_reg[21]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16327_
	);
	LUT4 #(
		.INIT('h60a0)
	) name14978 (
		\P2_rEIP_reg[22]/NET0131 ,
		_w9779_,
		_w15262_,
		_w15259_,
		_w16328_
	);
	LUT2 #(
		.INIT('h1)
	) name14979 (
		_w16327_,
		_w16328_,
		_w16329_
	);
	LUT2 #(
		.INIT('hb)
	) name14980 (
		_w16326_,
		_w16329_,
		_w16330_
	);
	LUT4 #(
		.INIT('h070f)
	) name14981 (
		\P1_rEIP_reg[21]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		\P1_rEIP_reg[23]/NET0131 ,
		_w15858_,
		_w16331_
	);
	LUT3 #(
		.INIT('h2a)
	) name14982 (
		_w1856_,
		_w11024_,
		_w15858_,
		_w16332_
	);
	LUT3 #(
		.INIT('hb0)
	) name14983 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[21]_pad ,
		_w16333_
	);
	LUT4 #(
		.INIT('h00b7)
	) name14984 (
		\P1_rEIP_reg[22]/NET0131 ,
		_w15287_,
		_w15862_,
		_w16333_,
		_w16334_
	);
	LUT3 #(
		.INIT('h4f)
	) name14985 (
		_w16331_,
		_w16332_,
		_w16334_,
		_w16335_
	);
	LUT3 #(
		.INIT('h08)
	) name14986 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16336_
	);
	LUT4 #(
		.INIT('he000)
	) name14987 (
		\P2_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready12_reg/NET0131 ,
		\ready21_reg/NET0131 ,
		_w16337_
	);
	LUT4 #(
		.INIT('h5444)
	) name14988 (
		na_pad,
		_w1610_,
		_w16336_,
		_w16337_,
		_w16338_
	);
	LUT3 #(
		.INIT('h0e)
	) name14989 (
		\P2_RequestPending_reg/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16339_
	);
	LUT2 #(
		.INIT('h8)
	) name14990 (
		\P2_State_reg[0]/NET0131 ,
		hold_pad,
		_w16340_
	);
	LUT2 #(
		.INIT('h8)
	) name14991 (
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16341_
	);
	LUT4 #(
		.INIT('h8acf)
	) name14992 (
		_w16271_,
		_w16339_,
		_w16340_,
		_w16341_,
		_w16342_
	);
	LUT2 #(
		.INIT('hb)
	) name14993 (
		_w16338_,
		_w16342_,
		_w16343_
	);
	LUT3 #(
		.INIT('h08)
	) name14994 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16344_
	);
	LUT2 #(
		.INIT('h1)
	) name14995 (
		\P3_RequestPending_reg/NET0131 ,
		hold_pad,
		_w16345_
	);
	LUT3 #(
		.INIT('h40)
	) name14996 (
		na_pad,
		\ready22_reg/NET0131 ,
		\ready2_pad ,
		_w16346_
	);
	LUT3 #(
		.INIT('h20)
	) name14997 (
		_w16344_,
		_w16345_,
		_w16346_,
		_w16347_
	);
	LUT2 #(
		.INIT('h8)
	) name14998 (
		hold_pad,
		_w16276_,
		_w16348_
	);
	LUT3 #(
		.INIT('h45)
	) name14999 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		na_pad,
		_w16349_
	);
	LUT3 #(
		.INIT('ha8)
	) name15000 (
		\P3_State_reg[2]/NET0131 ,
		_w16261_,
		_w16349_,
		_w16350_
	);
	LUT3 #(
		.INIT('hfe)
	) name15001 (
		_w16348_,
		_w16350_,
		_w16347_,
		_w16351_
	);
	LUT3 #(
		.INIT('h08)
	) name15002 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16352_
	);
	LUT4 #(
		.INIT('he000)
	) name15003 (
		\P1_RequestPending_reg/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16353_
	);
	LUT4 #(
		.INIT('h5444)
	) name15004 (
		na_pad,
		_w1857_,
		_w16352_,
		_w16353_,
		_w16354_
	);
	LUT2 #(
		.INIT('h2)
	) name15005 (
		\P1_RequestPending_reg/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16355_
	);
	LUT3 #(
		.INIT('h20)
	) name15006 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		hold_pad,
		_w16356_
	);
	LUT4 #(
		.INIT('h0222)
	) name15007 (
		\P1_State_reg[0]/NET0131 ,
		hold_pad,
		\ready11_reg/NET0131 ,
		\ready1_pad ,
		_w16357_
	);
	LUT2 #(
		.INIT('h8)
	) name15008 (
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16358_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name15009 (
		_w16355_,
		_w16356_,
		_w16357_,
		_w16358_,
		_w16359_
	);
	LUT2 #(
		.INIT('hb)
	) name15010 (
		_w16354_,
		_w16359_,
		_w16360_
	);
	LUT2 #(
		.INIT('h7)
	) name15011 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16361_
	);
	LUT4 #(
		.INIT('h7010)
	) name15012 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16362_
	);
	LUT3 #(
		.INIT('h01)
	) name15013 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16363_
	);
	LUT3 #(
		.INIT('h80)
	) name15014 (
		\P2_ByteEnable_reg[2]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16364_
	);
	LUT3 #(
		.INIT('hfe)
	) name15015 (
		_w16363_,
		_w16362_,
		_w16364_,
		_w16365_
	);
	LUT2 #(
		.INIT('h7)
	) name15016 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16366_
	);
	LUT4 #(
		.INIT('h7000)
	) name15017 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16367_
	);
	LUT3 #(
		.INIT('h80)
	) name15018 (
		\P1_ByteEnable_reg[2]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16368_
	);
	LUT4 #(
		.INIT('h0013)
	) name15019 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16369_
	);
	LUT3 #(
		.INIT('hfe)
	) name15020 (
		_w16368_,
		_w16367_,
		_w16369_,
		_w16370_
	);
	LUT2 #(
		.INIT('h7)
	) name15021 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16371_
	);
	LUT4 #(
		.INIT('h7010)
	) name15022 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16372_
	);
	LUT3 #(
		.INIT('h01)
	) name15023 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16373_
	);
	LUT3 #(
		.INIT('h80)
	) name15024 (
		\P3_ByteEnable_reg[2]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16374_
	);
	LUT3 #(
		.INIT('hfe)
	) name15025 (
		_w16373_,
		_w16372_,
		_w16374_,
		_w16375_
	);
	LUT3 #(
		.INIT('h01)
	) name15026 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		_w16376_
	);
	LUT4 #(
		.INIT('h407f)
	) name15027 (
		\P3_ByteEnable_reg[1]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16377_
	);
	LUT2 #(
		.INIT('hb)
	) name15028 (
		_w16376_,
		_w16377_,
		_w16378_
	);
	LUT3 #(
		.INIT('h01)
	) name15029 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		_w16379_
	);
	LUT4 #(
		.INIT('h407f)
	) name15030 (
		\P1_ByteEnable_reg[1]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16380_
	);
	LUT2 #(
		.INIT('hb)
	) name15031 (
		_w16379_,
		_w16380_,
		_w16381_
	);
	LUT3 #(
		.INIT('h01)
	) name15032 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		_w16382_
	);
	LUT4 #(
		.INIT('h407f)
	) name15033 (
		\P2_ByteEnable_reg[1]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16383_
	);
	LUT2 #(
		.INIT('hb)
	) name15034 (
		_w16382_,
		_w16383_,
		_w16384_
	);
	LUT3 #(
		.INIT('h48)
	) name15035 (
		\P3_rEIP_reg[3]/NET0131 ,
		_w2110_,
		_w15216_,
		_w16385_
	);
	LUT3 #(
		.INIT('h8a)
	) name15036 (
		\P3_Address_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16386_
	);
	LUT4 #(
		.INIT('h00b7)
	) name15037 (
		\P3_rEIP_reg[2]/NET0131 ,
		_w15237_,
		_w15886_,
		_w16386_,
		_w16387_
	);
	LUT2 #(
		.INIT('hb)
	) name15038 (
		_w16385_,
		_w16387_,
		_w16388_
	);
	LUT3 #(
		.INIT('h48)
	) name15039 (
		\P2_rEIP_reg[3]/NET0131 ,
		_w1609_,
		_w15243_,
		_w16389_
	);
	LUT3 #(
		.INIT('h8a)
	) name15040 (
		\P2_Address_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16390_
	);
	LUT4 #(
		.INIT('h00b7)
	) name15041 (
		\P2_rEIP_reg[2]/NET0131 ,
		_w15262_,
		_w15896_,
		_w16390_,
		_w16391_
	);
	LUT2 #(
		.INIT('hb)
	) name15042 (
		_w16389_,
		_w16391_,
		_w16392_
	);
	LUT3 #(
		.INIT('h48)
	) name15043 (
		\P1_rEIP_reg[3]/NET0131 ,
		_w1856_,
		_w15268_,
		_w16393_
	);
	LUT3 #(
		.INIT('hb0)
	) name15044 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[1]_pad ,
		_w16394_
	);
	LUT4 #(
		.INIT('h00b7)
	) name15045 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w15287_,
		_w15904_,
		_w16394_,
		_w16395_
	);
	LUT2 #(
		.INIT('hb)
	) name15046 (
		_w16393_,
		_w16395_,
		_w16396_
	);
	LUT4 #(
		.INIT('h4888)
	) name15047 (
		\P3_rEIP_reg[19]/NET0131 ,
		_w2110_,
		_w11970_,
		_w15225_,
		_w16397_
	);
	LUT3 #(
		.INIT('h8a)
	) name15048 (
		\P3_Address_reg[17]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16398_
	);
	LUT4 #(
		.INIT('h070f)
	) name15049 (
		\P3_rEIP_reg[16]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w15460_,
		_w16399_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15050 (
		_w11923_,
		_w11970_,
		_w15234_,
		_w15237_,
		_w16400_
	);
	LUT3 #(
		.INIT('h45)
	) name15051 (
		_w16398_,
		_w16399_,
		_w16400_,
		_w16401_
	);
	LUT2 #(
		.INIT('hb)
	) name15052 (
		_w16397_,
		_w16401_,
		_w16402_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15053 (
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w1856_,
		_w15278_,
		_w16403_
	);
	LUT3 #(
		.INIT('hb0)
	) name15054 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[17]_pad ,
		_w16404_
	);
	LUT4 #(
		.INIT('h9300)
	) name15055 (
		\P1_rEIP_reg[17]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		_w10858_,
		_w15284_,
		_w16405_
	);
	LUT3 #(
		.INIT('h13)
	) name15056 (
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[18]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w16406_
	);
	LUT2 #(
		.INIT('h2)
	) name15057 (
		_w15287_,
		_w16406_,
		_w16407_
	);
	LUT3 #(
		.INIT('h45)
	) name15058 (
		_w16404_,
		_w16405_,
		_w16407_,
		_w16408_
	);
	LUT2 #(
		.INIT('hb)
	) name15059 (
		_w16403_,
		_w16408_,
		_w16409_
	);
	LUT3 #(
		.INIT('h8a)
	) name15060 (
		\P2_Address_reg[17]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16410_
	);
	LUT3 #(
		.INIT('h13)
	) name15061 (
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[18]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16411_
	);
	LUT2 #(
		.INIT('h2)
	) name15062 (
		_w15262_,
		_w16411_,
		_w16412_
	);
	LUT4 #(
		.INIT('h040f)
	) name15063 (
		_w11302_,
		_w15259_,
		_w16410_,
		_w16412_,
		_w16413_
	);
	LUT4 #(
		.INIT('h48ff)
	) name15064 (
		\P2_rEIP_reg[19]/NET0131 ,
		_w1609_,
		_w15249_,
		_w16413_,
		_w16414_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15065 (
		\P3_rEIP_reg[6]/NET0131 ,
		\P3_rEIP_reg[7]/NET0131 ,
		_w2110_,
		_w15218_,
		_w16415_
	);
	LUT3 #(
		.INIT('h8a)
	) name15066 (
		\P3_Address_reg[5]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16416_
	);
	LUT4 #(
		.INIT('h00b7)
	) name15067 (
		\P3_rEIP_reg[6]/NET0131 ,
		_w15237_,
		_w15889_,
		_w16416_,
		_w16417_
	);
	LUT2 #(
		.INIT('hb)
	) name15068 (
		_w16415_,
		_w16417_,
		_w16418_
	);
	LUT3 #(
		.INIT('h13)
	) name15069 (
		\P2_rEIP_reg[6]/NET0131 ,
		\P2_rEIP_reg[7]/NET0131 ,
		_w15893_,
		_w16419_
	);
	LUT2 #(
		.INIT('h2)
	) name15070 (
		_w1609_,
		_w15245_,
		_w16420_
	);
	LUT3 #(
		.INIT('h8a)
	) name15071 (
		\P2_Address_reg[5]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16421_
	);
	LUT4 #(
		.INIT('h00b7)
	) name15072 (
		\P2_rEIP_reg[6]/NET0131 ,
		_w15262_,
		_w15899_,
		_w16421_,
		_w16422_
	);
	LUT3 #(
		.INIT('h4f)
	) name15073 (
		_w16419_,
		_w16420_,
		_w16422_,
		_w16423_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15074 (
		\P1_rEIP_reg[6]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w1856_,
		_w15270_,
		_w16424_
	);
	LUT3 #(
		.INIT('hb0)
	) name15075 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[5]_pad ,
		_w16425_
	);
	LUT4 #(
		.INIT('h0c08)
	) name15076 (
		\P1_rEIP_reg[6]/NET0131 ,
		_w15287_,
		_w15880_,
		_w15907_,
		_w16426_
	);
	LUT3 #(
		.INIT('hfe)
	) name15077 (
		_w16425_,
		_w16424_,
		_w16426_,
		_w16427_
	);
	LUT3 #(
		.INIT('h80)
	) name15078 (
		\P1_ByteEnable_reg[3]/NET0131 ,
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		_w16428_
	);
	LUT4 #(
		.INIT('h0133)
	) name15079 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_rEIP_reg[0]/NET0131 ,
		\P1_rEIP_reg[1]/NET0131 ,
		_w16429_
	);
	LUT2 #(
		.INIT('he)
	) name15080 (
		_w16428_,
		_w16429_,
		_w16430_
	);
	LUT3 #(
		.INIT('h80)
	) name15081 (
		\P3_ByteEnable_reg[3]/NET0131 ,
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		_w16431_
	);
	LUT4 #(
		.INIT('h0133)
	) name15082 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		_w16432_
	);
	LUT2 #(
		.INIT('he)
	) name15083 (
		_w16431_,
		_w16432_,
		_w16433_
	);
	LUT3 #(
		.INIT('h80)
	) name15084 (
		\P2_ByteEnable_reg[3]/NET0131 ,
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		_w16434_
	);
	LUT4 #(
		.INIT('h0133)
	) name15085 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		_w16435_
	);
	LUT2 #(
		.INIT('he)
	) name15086 (
		_w16434_,
		_w16435_,
		_w16436_
	);
	LUT3 #(
		.INIT('h48)
	) name15087 (
		\P1_rEIP_reg[2]/NET0131 ,
		_w1856_,
		_w15267_,
		_w16437_
	);
	LUT3 #(
		.INIT('hb0)
	) name15088 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\address1[0]_pad ,
		_w16438_
	);
	LUT4 #(
		.INIT('h009f)
	) name15089 (
		\P1_rEIP_reg[1]/NET0131 ,
		_w15284_,
		_w15287_,
		_w16438_,
		_w16439_
	);
	LUT2 #(
		.INIT('hb)
	) name15090 (
		_w16437_,
		_w16439_,
		_w16440_
	);
	LUT4 #(
		.INIT('h28a0)
	) name15091 (
		\P2_State_reg[2]/NET0131 ,
		\P2_rEIP_reg[0]/NET0131 ,
		\P2_rEIP_reg[1]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w16441_
	);
	LUT4 #(
		.INIT('h00eb)
	) name15092 (
		\P2_State_reg[2]/NET0131 ,
		\P2_rEIP_reg[2]/NET0131 ,
		_w15242_,
		_w16441_,
		_w16442_
	);
	LUT3 #(
		.INIT('h2e)
	) name15093 (
		\P2_Address_reg[0]/NET0131 ,
		_w1608_,
		_w16442_,
		_w16443_
	);
	LUT4 #(
		.INIT('h28a0)
	) name15094 (
		\P3_State_reg[2]/NET0131 ,
		\P3_rEIP_reg[0]/NET0131 ,
		\P3_rEIP_reg[1]/NET0131 ,
		\P3_rEIP_reg[31]/NET0131 ,
		_w16444_
	);
	LUT4 #(
		.INIT('h00eb)
	) name15095 (
		\P3_State_reg[2]/NET0131 ,
		\P3_rEIP_reg[2]/NET0131 ,
		_w15215_,
		_w16444_,
		_w16445_
	);
	LUT3 #(
		.INIT('h2e)
	) name15096 (
		\P3_Address_reg[0]/NET0131 ,
		_w2109_,
		_w16445_,
		_w16446_
	);
	LUT3 #(
		.INIT('h40)
	) name15097 (
		\P2_Address_reg[29]/NET0131 ,
		_w16025_,
		_w16026_,
		_w16447_
	);
	LUT3 #(
		.INIT('hbf)
	) name15098 (
		\P2_Address_reg[29]/NET0131 ,
		_w16025_,
		_w16026_,
		_w16448_
	);
	LUT4 #(
		.INIT('h0010)
	) name15099 (
		\ast2_pad ,
		dc_pad,
		mio_pad,
		wr_pad,
		_w16449_
	);
	LUT4 #(
		.INIT('h0001)
	) name15100 (
		\P3_BE_n_reg[0]/NET0131 ,
		\P3_BE_n_reg[1]/NET0131 ,
		\P3_BE_n_reg[2]/NET0131 ,
		\P3_BE_n_reg[3]/NET0131 ,
		_w16450_
	);
	LUT2 #(
		.INIT('h8)
	) name15101 (
		_w16449_,
		_w16450_,
		_w16451_
	);
	LUT2 #(
		.INIT('hb)
	) name15102 (
		_w16447_,
		_w16451_,
		_w16452_
	);
	LUT4 #(
		.INIT('h5414)
	) name15103 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16453_
	);
	LUT4 #(
		.INIT('h0018)
	) name15104 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16454_
	);
	LUT2 #(
		.INIT('h1)
	) name15105 (
		_w16453_,
		_w16454_,
		_w16455_
	);
	LUT4 #(
		.INIT('h0018)
	) name15106 (
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16456_
	);
	LUT4 #(
		.INIT('h5414)
	) name15107 (
		\P2_DataWidth_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16457_
	);
	LUT2 #(
		.INIT('h1)
	) name15108 (
		_w16456_,
		_w16457_,
		_w16458_
	);
	LUT4 #(
		.INIT('h0018)
	) name15109 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		\bs16_pad ,
		_w16459_
	);
	LUT4 #(
		.INIT('h5414)
	) name15110 (
		\P1_DataWidth_reg[1]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16460_
	);
	LUT2 #(
		.INIT('h1)
	) name15111 (
		_w16459_,
		_w16460_,
		_w16461_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15112 (
		\P1_BE_n_reg[2]/NET0131 ,
		\P1_ByteEnable_reg[2]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16462_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15113 (
		\P1_BE_n_reg[3]/NET0131 ,
		\P1_ByteEnable_reg[3]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16463_
	);
	LUT4 #(
		.INIT('hbb19)
	) name15114 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		\ast2_pad ,
		_w16464_
	);
	LUT4 #(
		.INIT('ha828)
	) name15115 (
		\P3_DataWidth_reg[0]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		_w16465_
	);
	LUT2 #(
		.INIT('he)
	) name15116 (
		_w16454_,
		_w16465_,
		_w16466_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15117 (
		\P2_BE_n_reg[0]/NET0131 ,
		\P2_ByteEnable_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16467_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15118 (
		\P2_BE_n_reg[3]/NET0131 ,
		\P2_ByteEnable_reg[3]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16468_
	);
	LUT4 #(
		.INIT('ha828)
	) name15119 (
		\P2_DataWidth_reg[0]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16469_
	);
	LUT2 #(
		.INIT('he)
	) name15120 (
		_w16456_,
		_w16469_,
		_w16470_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15121 (
		\P3_BE_n_reg[3]/NET0131 ,
		\P3_ByteEnable_reg[3]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16471_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15122 (
		\P3_BE_n_reg[1]/NET0131 ,
		\P3_ByteEnable_reg[1]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16472_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15123 (
		\P3_BE_n_reg[2]/NET0131 ,
		\P3_ByteEnable_reg[2]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16473_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15124 (
		\P3_BE_n_reg[0]/NET0131 ,
		\P3_ByteEnable_reg[0]/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16474_
	);
	LUT4 #(
		.INIT('hbb19)
	) name15125 (
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		\ast1_pad ,
		_w16475_
	);
	LUT4 #(
		.INIT('h8bcb)
	) name15126 (
		\P2_ADS_n_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16476_
	);
	LUT4 #(
		.INIT('hef20)
	) name15127 (
		\P3_MemoryFetch_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		mio_pad,
		_w16477_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15128 (
		\P3_ReadRequest_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		wr_pad,
		_w16478_
	);
	LUT4 #(
		.INIT('ha828)
	) name15129 (
		\P1_DataWidth_reg[0]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16479_
	);
	LUT2 #(
		.INIT('he)
	) name15130 (
		_w16459_,
		_w16479_,
		_w16480_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15131 (
		\P1_M_IO_n_reg/NET0131 ,
		\P1_MemoryFetch_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16481_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15132 (
		\P2_BE_n_reg[2]/NET0131 ,
		\P2_ByteEnable_reg[2]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16482_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15133 (
		\P2_ReadRequest_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_W_R_n_reg/NET0131 ,
		_w16483_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15134 (
		\P2_BE_n_reg[1]/NET0131 ,
		\P2_ByteEnable_reg[1]/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16484_
	);
	LUT4 #(
		.INIT('hdf10)
	) name15135 (
		\P1_ReadRequest_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_W_R_n_reg/NET0131 ,
		_w16485_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15136 (
		\P1_BE_n_reg[0]/NET0131 ,
		\P1_ByteEnable_reg[0]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16486_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15137 (
		\P2_M_IO_n_reg/NET0131 ,
		\P2_MemoryFetch_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16487_
	);
	LUT4 #(
		.INIT('hacaa)
	) name15138 (
		\P1_BE_n_reg[1]/NET0131 ,
		\P1_ByteEnable_reg[1]/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16488_
	);
	LUT4 #(
		.INIT('h00ba)
	) name15139 (
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		\P3_State_reg[2]/NET0131 ,
		dc_pad,
		_w16489_
	);
	LUT3 #(
		.INIT('h20)
	) name15140 (
		\P3_CodeFetch_reg/NET0131 ,
		\P3_State_reg[0]/NET0131 ,
		\P3_State_reg[1]/NET0131 ,
		_w16490_
	);
	LUT2 #(
		.INIT('h1)
	) name15141 (
		_w16489_,
		_w16490_,
		_w16491_
	);
	LUT4 #(
		.INIT('h4544)
	) name15142 (
		\P2_D_C_n_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		\P2_State_reg[2]/NET0131 ,
		_w16492_
	);
	LUT3 #(
		.INIT('h20)
	) name15143 (
		\P2_CodeFetch_reg/NET0131 ,
		\P2_State_reg[0]/NET0131 ,
		\P2_State_reg[1]/NET0131 ,
		_w16493_
	);
	LUT2 #(
		.INIT('h1)
	) name15144 (
		_w16492_,
		_w16493_,
		_w16494_
	);
	LUT4 #(
		.INIT('h4544)
	) name15145 (
		\P1_D_C_n_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		\P1_State_reg[2]/NET0131 ,
		_w16495_
	);
	LUT3 #(
		.INIT('h20)
	) name15146 (
		\P1_CodeFetch_reg/NET0131 ,
		\P1_State_reg[0]/NET0131 ,
		\P1_State_reg[1]/NET0131 ,
		_w16496_
	);
	LUT2 #(
		.INIT('h1)
	) name15147 (
		_w16495_,
		_w16496_,
		_w16497_
	);
	LUT3 #(
		.INIT('h02)
	) name15148 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16498_
	);
	LUT4 #(
		.INIT('haa20)
	) name15149 (
		_w2171_,
		_w8663_,
		_w8666_,
		_w16498_,
		_w16499_
	);
	LUT4 #(
		.INIT('he000)
	) name15150 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w2987_,
		_w16500_
	);
	LUT4 #(
		.INIT('h004f)
	) name15151 (
		_w2073_,
		_w2086_,
		_w2869_,
		_w16500_,
		_w16501_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15152 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16502_
	);
	LUT2 #(
		.INIT('h4)
	) name15153 (
		_w2117_,
		_w4052_,
		_w16503_
	);
	LUT3 #(
		.INIT('h10)
	) name15154 (
		_w16502_,
		_w16503_,
		_w16501_,
		_w16504_
	);
	LUT2 #(
		.INIT('h4)
	) name15155 (
		_w8669_,
		_w16504_,
		_w16505_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15156 (
		\P3_InstAddrPointer_reg[10]/NET0131 ,
		\P3_rEIP_reg[10]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16506_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15157 (
		_w1945_,
		_w16499_,
		_w16505_,
		_w16506_,
		_w16507_
	);
	LUT4 #(
		.INIT('h7774)
	) name15158 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2173_,
		_w6977_,
		_w6974_,
		_w16508_
	);
	LUT2 #(
		.INIT('h2)
	) name15159 (
		_w2171_,
		_w16508_,
		_w16509_
	);
	LUT4 #(
		.INIT('he000)
	) name15160 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w6981_,
		_w16510_
	);
	LUT3 #(
		.INIT('h0e)
	) name15161 (
		_w2071_,
		_w2087_,
		_w4082_,
		_w16511_
	);
	LUT4 #(
		.INIT('h0002)
	) name15162 (
		_w2126_,
		_w2127_,
		_w2175_,
		_w16511_,
		_w16512_
	);
	LUT3 #(
		.INIT('hb0)
	) name15163 (
		_w2073_,
		_w2086_,
		_w2731_,
		_w16513_
	);
	LUT4 #(
		.INIT('h0020)
	) name15164 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w2060_,
		_w2047_,
		_w2105_,
		_w16514_
	);
	LUT3 #(
		.INIT('hc4)
	) name15165 (
		_w2117_,
		_w6975_,
		_w16514_,
		_w16515_
	);
	LUT4 #(
		.INIT('h0031)
	) name15166 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		_w16513_,
		_w16512_,
		_w16515_,
		_w16516_
	);
	LUT2 #(
		.INIT('h4)
	) name15167 (
		_w16510_,
		_w16516_,
		_w16517_
	);
	LUT3 #(
		.INIT('hb0)
	) name15168 (
		_w6982_,
		_w6983_,
		_w16517_,
		_w16518_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15169 (
		\P3_InstAddrPointer_reg[29]/NET0131 ,
		\P3_rEIP_reg[29]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16519_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15170 (
		_w1945_,
		_w16509_,
		_w16518_,
		_w16519_,
		_w16520_
	);
	LUT3 #(
		.INIT('h08)
	) name15171 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16521_
	);
	LUT4 #(
		.INIT('h004f)
	) name15172 (
		_w7363_,
		_w7364_,
		_w7366_,
		_w16521_,
		_w16522_
	);
	LUT2 #(
		.INIT('h8)
	) name15173 (
		_w1640_,
		_w6899_,
		_w16523_
	);
	LUT4 #(
		.INIT('h004f)
	) name15174 (
		_w1571_,
		_w1583_,
		_w4345_,
		_w16523_,
		_w16524_
	);
	LUT3 #(
		.INIT('h2a)
	) name15175 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		_w1614_,
		_w1668_,
		_w16525_
	);
	LUT2 #(
		.INIT('h4)
	) name15176 (
		_w1617_,
		_w4256_,
		_w16526_
	);
	LUT3 #(
		.INIT('h10)
	) name15177 (
		_w16525_,
		_w16526_,
		_w16524_,
		_w16527_
	);
	LUT3 #(
		.INIT('hb0)
	) name15178 (
		_w7369_,
		_w7370_,
		_w16527_,
		_w16528_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15179 (
		_w1559_,
		_w1678_,
		_w16522_,
		_w16528_,
		_w16529_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15180 (
		\P2_InstAddrPointer_reg[20]/NET0131 ,
		\P2_rEIP_reg[20]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16530_
	);
	LUT2 #(
		.INIT('hb)
	) name15181 (
		_w16529_,
		_w16530_,
		_w16531_
	);
	LUT3 #(
		.INIT('h08)
	) name15182 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16532_
	);
	LUT4 #(
		.INIT('haa20)
	) name15183 (
		_w1559_,
		_w5703_,
		_w5709_,
		_w16532_,
		_w16533_
	);
	LUT2 #(
		.INIT('h2)
	) name15184 (
		_w1640_,
		_w5719_,
		_w16534_
	);
	LUT3 #(
		.INIT('h0b)
	) name15185 (
		_w1571_,
		_w1583_,
		_w5702_,
		_w16535_
	);
	LUT2 #(
		.INIT('h4)
	) name15186 (
		_w1617_,
		_w5708_,
		_w16536_
	);
	LUT3 #(
		.INIT('h2a)
	) name15187 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		_w1614_,
		_w1668_,
		_w16537_
	);
	LUT4 #(
		.INIT('h0001)
	) name15188 (
		_w16535_,
		_w16536_,
		_w16537_,
		_w16534_,
		_w16538_
	);
	LUT4 #(
		.INIT('h7d00)
	) name15189 (
		_w1659_,
		_w5718_,
		_w5719_,
		_w16538_,
		_w16539_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15190 (
		\P2_InstAddrPointer_reg[31]/NET0131 ,
		\P2_rEIP_reg[31]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16540_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15191 (
		_w1678_,
		_w16533_,
		_w16539_,
		_w16540_,
		_w16541_
	);
	LUT3 #(
		.INIT('h02)
	) name15192 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16542_
	);
	LUT4 #(
		.INIT('haa20)
	) name15193 (
		_w2171_,
		_w7956_,
		_w7959_,
		_w16542_,
		_w16543_
	);
	LUT4 #(
		.INIT('he000)
	) name15194 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7962_,
		_w16544_
	);
	LUT3 #(
		.INIT('h0b)
	) name15195 (
		_w2117_,
		_w5358_,
		_w16544_,
		_w16545_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15196 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16546_
	);
	LUT3 #(
		.INIT('hb0)
	) name15197 (
		_w2073_,
		_w2086_,
		_w2883_,
		_w16547_
	);
	LUT3 #(
		.INIT('h10)
	) name15198 (
		_w16546_,
		_w16547_,
		_w16545_,
		_w16548_
	);
	LUT2 #(
		.INIT('h4)
	) name15199 (
		_w7965_,
		_w16548_,
		_w16549_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15200 (
		\P3_InstAddrPointer_reg[13]/NET0131 ,
		\P3_rEIP_reg[13]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16550_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15201 (
		_w1945_,
		_w16543_,
		_w16549_,
		_w16550_,
		_w16551_
	);
	LUT3 #(
		.INIT('h08)
	) name15202 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16552_
	);
	LUT4 #(
		.INIT('haa20)
	) name15203 (
		_w1559_,
		_w7653_,
		_w7655_,
		_w16552_,
		_w16553_
	);
	LUT2 #(
		.INIT('h8)
	) name15204 (
		_w1640_,
		_w4873_,
		_w16554_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15205 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		_w1614_,
		_w1668_,
		_w16554_,
		_w16555_
	);
	LUT3 #(
		.INIT('hb0)
	) name15206 (
		_w1571_,
		_w1583_,
		_w4346_,
		_w16556_
	);
	LUT2 #(
		.INIT('h4)
	) name15207 (
		_w1617_,
		_w4898_,
		_w16557_
	);
	LUT3 #(
		.INIT('h10)
	) name15208 (
		_w16556_,
		_w16557_,
		_w16555_,
		_w16558_
	);
	LUT2 #(
		.INIT('h4)
	) name15209 (
		_w7658_,
		_w16558_,
		_w16559_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15210 (
		\P2_InstAddrPointer_reg[19]/NET0131 ,
		\P2_rEIP_reg[19]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16560_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15211 (
		_w1678_,
		_w16553_,
		_w16559_,
		_w16560_,
		_w16561_
	);
	LUT3 #(
		.INIT('h02)
	) name15212 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16562_
	);
	LUT4 #(
		.INIT('haa20)
	) name15213 (
		_w2171_,
		_w6338_,
		_w6343_,
		_w16562_,
		_w16563_
	);
	LUT4 #(
		.INIT('he000)
	) name15214 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3041_,
		_w16564_
	);
	LUT2 #(
		.INIT('h1)
	) name15215 (
		_w2117_,
		_w2978_,
		_w16565_
	);
	LUT3 #(
		.INIT('hb0)
	) name15216 (
		_w2073_,
		_w2086_,
		_w2743_,
		_w16566_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15217 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16567_
	);
	LUT4 #(
		.INIT('h0001)
	) name15218 (
		_w16566_,
		_w16567_,
		_w16565_,
		_w16564_,
		_w16568_
	);
	LUT2 #(
		.INIT('h4)
	) name15219 (
		_w6346_,
		_w16568_,
		_w16569_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15220 (
		\P3_InstAddrPointer_reg[30]/NET0131 ,
		\P3_rEIP_reg[30]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16570_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15221 (
		_w1945_,
		_w16563_,
		_w16569_,
		_w16570_,
		_w16571_
	);
	LUT3 #(
		.INIT('h08)
	) name15222 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16572_
	);
	LUT4 #(
		.INIT('haa20)
	) name15223 (
		_w1559_,
		_w6313_,
		_w6318_,
		_w16572_,
		_w16573_
	);
	LUT4 #(
		.INIT('h80c0)
	) name15224 (
		_w1555_,
		_w1614_,
		_w1668_,
		_w6321_,
		_w16574_
	);
	LUT2 #(
		.INIT('h2)
	) name15225 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		_w16574_,
		_w16575_
	);
	LUT3 #(
		.INIT('h40)
	) name15226 (
		_w1555_,
		_w1596_,
		_w6321_,
		_w16576_
	);
	LUT2 #(
		.INIT('h4)
	) name15227 (
		_w1617_,
		_w6314_,
		_w16577_
	);
	LUT3 #(
		.INIT('hb0)
	) name15228 (
		_w1571_,
		_w1583_,
		_w5699_,
		_w16578_
	);
	LUT3 #(
		.INIT('h01)
	) name15229 (
		_w16577_,
		_w16578_,
		_w16576_,
		_w16579_
	);
	LUT2 #(
		.INIT('h4)
	) name15230 (
		_w16575_,
		_w16579_,
		_w16580_
	);
	LUT3 #(
		.INIT('hb0)
	) name15231 (
		_w6323_,
		_w6324_,
		_w16580_,
		_w16581_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15232 (
		\P2_InstAddrPointer_reg[30]/NET0131 ,
		\P2_rEIP_reg[30]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16582_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15233 (
		_w1678_,
		_w16573_,
		_w16581_,
		_w16582_,
		_w16583_
	);
	LUT2 #(
		.INIT('h6)
	) name15234 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w3029_,
		_w16584_
	);
	LUT4 #(
		.INIT('h007f)
	) name15235 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w3025_,
		_w3027_,
		_w16584_,
		_w16585_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name15236 (
		_w2181_,
		_w2708_,
		_w3025_,
		_w3027_,
		_w16586_
	);
	LUT2 #(
		.INIT('h4)
	) name15237 (
		_w16585_,
		_w16586_,
		_w16587_
	);
	LUT4 #(
		.INIT('h7f00)
	) name15238 (
		_w2874_,
		_w2884_,
		_w2897_,
		_w2913_,
		_w16588_
	);
	LUT3 #(
		.INIT('h01)
	) name15239 (
		_w2755_,
		_w6929_,
		_w16588_,
		_w16589_
	);
	LUT2 #(
		.INIT('h2)
	) name15240 (
		_w2967_,
		_w2960_,
		_w16590_
	);
	LUT4 #(
		.INIT('h1115)
	) name15241 (
		_w2173_,
		_w2755_,
		_w4058_,
		_w16590_,
		_w16591_
	);
	LUT3 #(
		.INIT('h20)
	) name15242 (
		_w2171_,
		_w16589_,
		_w16591_,
		_w16592_
	);
	LUT4 #(
		.INIT('he000)
	) name15243 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w16584_,
		_w16593_
	);
	LUT2 #(
		.INIT('h1)
	) name15244 (
		_w2117_,
		_w2967_,
		_w16594_
	);
	LUT3 #(
		.INIT('hb0)
	) name15245 (
		_w2073_,
		_w2086_,
		_w2913_,
		_w16595_
	);
	LUT4 #(
		.INIT('h000d)
	) name15246 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		_w7103_,
		_w16594_,
		_w16595_,
		_w16596_
	);
	LUT2 #(
		.INIT('h4)
	) name15247 (
		_w16593_,
		_w16596_,
		_w16597_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15248 (
		_w1945_,
		_w16592_,
		_w16587_,
		_w16597_,
		_w16598_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15249 (
		\P3_InstAddrPointer_reg[19]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16599_
	);
	LUT2 #(
		.INIT('hb)
	) name15250 (
		_w16598_,
		_w16599_,
		_w16600_
	);
	LUT3 #(
		.INIT('h01)
	) name15251 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16601_
	);
	LUT3 #(
		.INIT('h04)
	) name15252 (
		_w2060_,
		_w2041_,
		_w16601_,
		_w16602_
	);
	LUT4 #(
		.INIT('hab00)
	) name15253 (
		_w2173_,
		_w8009_,
		_w8012_,
		_w16602_,
		_w16603_
	);
	LUT4 #(
		.INIT('he000)
	) name15254 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w8015_,
		_w16604_
	);
	LUT3 #(
		.INIT('h0b)
	) name15255 (
		_w2117_,
		_w8008_,
		_w16604_,
		_w16605_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15256 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16606_
	);
	LUT3 #(
		.INIT('hb0)
	) name15257 (
		_w2073_,
		_w2086_,
		_w2896_,
		_w16607_
	);
	LUT3 #(
		.INIT('h10)
	) name15258 (
		_w16606_,
		_w16607_,
		_w16605_,
		_w16608_
	);
	LUT2 #(
		.INIT('h4)
	) name15259 (
		_w8016_,
		_w16608_,
		_w16609_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15260 (
		\P3_InstAddrPointer_reg[18]/NET0131 ,
		\P3_rEIP_reg[18]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16610_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15261 (
		_w1945_,
		_w16603_,
		_w16609_,
		_w16610_,
		_w16611_
	);
	LUT3 #(
		.INIT('h02)
	) name15262 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16612_
	);
	LUT4 #(
		.INIT('haa20)
	) name15263 (
		_w2171_,
		_w7975_,
		_w7978_,
		_w16612_,
		_w16613_
	);
	LUT4 #(
		.INIT('he000)
	) name15264 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3023_,
		_w16614_
	);
	LUT4 #(
		.INIT('h004f)
	) name15265 (
		_w2073_,
		_w2086_,
		_w2881_,
		_w16614_,
		_w16615_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15266 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16616_
	);
	LUT2 #(
		.INIT('h4)
	) name15267 (
		_w2117_,
		_w2949_,
		_w16617_
	);
	LUT4 #(
		.INIT('h0100)
	) name15268 (
		_w7980_,
		_w16616_,
		_w16617_,
		_w16615_,
		_w16618_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15269 (
		\P3_InstAddrPointer_reg[14]/NET0131 ,
		\P3_rEIP_reg[14]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16619_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15270 (
		_w1945_,
		_w16613_,
		_w16618_,
		_w16619_,
		_w16620_
	);
	LUT3 #(
		.INIT('h02)
	) name15271 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16621_
	);
	LUT4 #(
		.INIT('haa20)
	) name15272 (
		_w2171_,
		_w7505_,
		_w7506_,
		_w16621_,
		_w16622_
	);
	LUT4 #(
		.INIT('he000)
	) name15273 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7509_,
		_w16623_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15274 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16624_
	);
	LUT2 #(
		.INIT('h4)
	) name15275 (
		_w2117_,
		_w2969_,
		_w16625_
	);
	LUT3 #(
		.INIT('hb0)
	) name15276 (
		_w2073_,
		_w2086_,
		_w2911_,
		_w16626_
	);
	LUT4 #(
		.INIT('h0001)
	) name15277 (
		_w16623_,
		_w16625_,
		_w16626_,
		_w16624_,
		_w16627_
	);
	LUT4 #(
		.INIT('hfd00)
	) name15278 (
		_w2181_,
		_w4090_,
		_w7510_,
		_w16627_,
		_w16628_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15279 (
		\P3_InstAddrPointer_reg[26]/NET0131 ,
		\P3_rEIP_reg[26]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16629_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15280 (
		_w1945_,
		_w16622_,
		_w16628_,
		_w16629_,
		_w16630_
	);
	LUT3 #(
		.INIT('h08)
	) name15281 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16631_
	);
	LUT3 #(
		.INIT('h93)
	) name15282 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w3081_,
		_w16632_
	);
	LUT3 #(
		.INIT('h80)
	) name15283 (
		\P1_InstAddrPointer_reg[29]/NET0131 ,
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		_w3319_,
		_w16633_
	);
	LUT4 #(
		.INIT('he000)
	) name15284 (
		_w4445_,
		_w4447_,
		_w4453_,
		_w16633_,
		_w16634_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name15285 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w3080_,
		_w3322_,
		_w16635_
	);
	LUT4 #(
		.INIT('h1551)
	) name15286 (
		_w1916_,
		_w3101_,
		_w16634_,
		_w16635_,
		_w16636_
	);
	LUT4 #(
		.INIT('heb00)
	) name15287 (
		_w3101_,
		_w3265_,
		_w16632_,
		_w16636_,
		_w16637_
	);
	LUT4 #(
		.INIT('h8000)
	) name15288 (
		_w3392_,
		_w4481_,
		_w4483_,
		_w7019_,
		_w16638_
	);
	LUT4 #(
		.INIT('h9333)
	) name15289 (
		\P1_InstAddrPointer_reg[30]/NET0131 ,
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w3322_,
		_w3387_,
		_w16639_
	);
	LUT2 #(
		.INIT('h2)
	) name15290 (
		_w1847_,
		_w16639_,
		_w16640_
	);
	LUT3 #(
		.INIT('h0b)
	) name15291 (
		_w1816_,
		_w1831_,
		_w16632_,
		_w16641_
	);
	LUT2 #(
		.INIT('h4)
	) name15292 (
		_w1862_,
		_w16635_,
		_w16642_
	);
	LUT2 #(
		.INIT('h1)
	) name15293 (
		_w1867_,
		_w4710_,
		_w16643_
	);
	LUT4 #(
		.INIT('haa2a)
	) name15294 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		_w1914_,
		_w8833_,
		_w16643_,
		_w16644_
	);
	LUT4 #(
		.INIT('h0001)
	) name15295 (
		_w16642_,
		_w16641_,
		_w16640_,
		_w16644_,
		_w16645_
	);
	LUT4 #(
		.INIT('h7d00)
	) name15296 (
		_w1924_,
		_w16638_,
		_w16639_,
		_w16645_,
		_w16646_
	);
	LUT4 #(
		.INIT('h5700)
	) name15297 (
		_w1810_,
		_w16631_,
		_w16637_,
		_w16646_,
		_w16647_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15298 (
		\P1_InstAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16648_
	);
	LUT3 #(
		.INIT('h2f)
	) name15299 (
		_w1933_,
		_w16647_,
		_w16648_,
		_w16649_
	);
	LUT3 #(
		.INIT('h08)
	) name15300 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16650_
	);
	LUT3 #(
		.INIT('h40)
	) name15301 (
		_w1833_,
		_w1846_,
		_w3388_,
		_w16651_
	);
	LUT3 #(
		.INIT('h2a)
	) name15302 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		_w1922_,
		_w4037_,
		_w16652_
	);
	LUT3 #(
		.INIT('hb0)
	) name15303 (
		_w1816_,
		_w1831_,
		_w3260_,
		_w16653_
	);
	LUT2 #(
		.INIT('h4)
	) name15304 (
		_w1862_,
		_w3314_,
		_w16654_
	);
	LUT4 #(
		.INIT('h0001)
	) name15305 (
		_w16652_,
		_w16653_,
		_w16654_,
		_w16651_,
		_w16655_
	);
	LUT4 #(
		.INIT('hd700)
	) name15306 (
		_w1924_,
		_w3388_,
		_w7020_,
		_w16655_,
		_w16656_
	);
	LUT4 #(
		.INIT('h5700)
	) name15307 (
		_w1810_,
		_w7017_,
		_w16650_,
		_w16656_,
		_w16657_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15308 (
		\P1_InstAddrPointer_reg[27]/NET0131 ,
		\P1_rEIP_reg[27]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16658_
	);
	LUT3 #(
		.INIT('h2f)
	) name15309 (
		_w1933_,
		_w16657_,
		_w16658_,
		_w16659_
	);
	LUT3 #(
		.INIT('h02)
	) name15310 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16660_
	);
	LUT4 #(
		.INIT('h1405)
	) name15311 (
		_w2755_,
		_w2886_,
		_w2889_,
		_w4751_,
		_w16661_
	);
	LUT4 #(
		.INIT('h8222)
	) name15312 (
		_w2755_,
		_w5360_,
		_w5357_,
		_w5359_,
		_w16662_
	);
	LUT2 #(
		.INIT('h1)
	) name15313 (
		_w2173_,
		_w16662_,
		_w16663_
	);
	LUT4 #(
		.INIT('h8a88)
	) name15314 (
		_w2171_,
		_w16660_,
		_w16661_,
		_w16663_,
		_w16664_
	);
	LUT3 #(
		.INIT('h28)
	) name15315 (
		_w2181_,
		_w3025_,
		_w3027_,
		_w16665_
	);
	LUT4 #(
		.INIT('he000)
	) name15316 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3027_,
		_w16666_
	);
	LUT4 #(
		.INIT('h004f)
	) name15317 (
		_w2073_,
		_w2086_,
		_w2889_,
		_w16666_,
		_w16667_
	);
	LUT2 #(
		.INIT('h4)
	) name15318 (
		_w2117_,
		_w5360_,
		_w16668_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15319 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16669_
	);
	LUT3 #(
		.INIT('h10)
	) name15320 (
		_w16668_,
		_w16669_,
		_w16667_,
		_w16670_
	);
	LUT2 #(
		.INIT('h4)
	) name15321 (
		_w16665_,
		_w16670_,
		_w16671_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15322 (
		\P3_InstAddrPointer_reg[17]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16672_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15323 (
		_w1945_,
		_w16664_,
		_w16671_,
		_w16672_,
		_w16673_
	);
	LUT3 #(
		.INIT('h02)
	) name15324 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16674_
	);
	LUT4 #(
		.INIT('h004f)
	) name15325 (
		_w6931_,
		_w6932_,
		_w6934_,
		_w16674_,
		_w16675_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name15326 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w2060_,
		_w2044_,
		_w2047_,
		_w16676_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name15327 (
		_w2108_,
		_w2115_,
		_w2116_,
		_w16676_,
		_w16677_
	);
	LUT4 #(
		.INIT('hf111)
	) name15328 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3033_,
		_w16678_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name15329 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		_w4785_,
		_w16677_,
		_w16678_,
		_w16679_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name15330 (
		_w2108_,
		_w2115_,
		_w2116_,
		_w16676_,
		_w16680_
	);
	LUT3 #(
		.INIT('hc8)
	) name15331 (
		_w2064_,
		_w2971_,
		_w16680_,
		_w16681_
	);
	LUT4 #(
		.INIT('he000)
	) name15332 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w6926_,
		_w16682_
	);
	LUT4 #(
		.INIT('h004f)
	) name15333 (
		_w2073_,
		_w2086_,
		_w2906_,
		_w16682_,
		_w16683_
	);
	LUT3 #(
		.INIT('h10)
	) name15334 (
		_w16681_,
		_w16679_,
		_w16683_,
		_w16684_
	);
	LUT4 #(
		.INIT('h3100)
	) name15335 (
		_w2171_,
		_w6927_,
		_w16675_,
		_w16684_,
		_w16685_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15336 (
		\P3_InstAddrPointer_reg[23]/NET0131 ,
		\P3_rEIP_reg[23]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16686_
	);
	LUT3 #(
		.INIT('h2f)
	) name15337 (
		_w1945_,
		_w16685_,
		_w16686_,
		_w16687_
	);
	LUT4 #(
		.INIT('h3f35)
	) name15338 (
		\P3_EBX_reg[27]/NET0131 ,
		_w8438_,
		_w8923_,
		_w8924_,
		_w16688_
	);
	LUT4 #(
		.INIT('hb700)
	) name15339 (
		\P3_EBX_reg[27]/NET0131 ,
		_w2084_,
		_w10253_,
		_w16688_,
		_w16689_
	);
	LUT2 #(
		.INIT('h2)
	) name15340 (
		\P3_EBX_reg[27]/NET0131 ,
		_w8341_,
		_w16690_
	);
	LUT3 #(
		.INIT('hf2)
	) name15341 (
		_w1945_,
		_w16689_,
		_w16690_,
		_w16691_
	);
	LUT4 #(
		.INIT('h4744)
	) name15342 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w1661_,
		_w8218_,
		_w8219_,
		_w16692_
	);
	LUT2 #(
		.INIT('h8)
	) name15343 (
		_w1640_,
		_w4411_,
		_w16693_
	);
	LUT3 #(
		.INIT('h0b)
	) name15344 (
		_w1617_,
		_w4240_,
		_w16693_,
		_w16694_
	);
	LUT3 #(
		.INIT('hb0)
	) name15345 (
		_w1571_,
		_w1583_,
		_w4328_,
		_w16695_
	);
	LUT3 #(
		.INIT('h2a)
	) name15346 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		_w1658_,
		_w4844_,
		_w16696_
	);
	LUT3 #(
		.INIT('h10)
	) name15347 (
		_w16695_,
		_w16696_,
		_w16694_,
		_w16697_
	);
	LUT2 #(
		.INIT('h4)
	) name15348 (
		_w8224_,
		_w16697_,
		_w16698_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15349 (
		_w1559_,
		_w1678_,
		_w16692_,
		_w16698_,
		_w16699_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15350 (
		\P2_InstAddrPointer_reg[14]/NET0131 ,
		\P2_rEIP_reg[14]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16700_
	);
	LUT2 #(
		.INIT('hb)
	) name15351 (
		_w16699_,
		_w16700_,
		_w16701_
	);
	LUT3 #(
		.INIT('h02)
	) name15352 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16702_
	);
	LUT4 #(
		.INIT('haa20)
	) name15353 (
		_w2171_,
		_w7457_,
		_w7459_,
		_w16702_,
		_w16703_
	);
	LUT4 #(
		.INIT('he000)
	) name15354 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7462_,
		_w16704_
	);
	LUT3 #(
		.INIT('hb0)
	) name15355 (
		_w2073_,
		_w2086_,
		_w2900_,
		_w16705_
	);
	LUT2 #(
		.INIT('h4)
	) name15356 (
		_w2117_,
		_w2965_,
		_w16706_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15357 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16707_
	);
	LUT4 #(
		.INIT('h0001)
	) name15358 (
		_w16704_,
		_w16706_,
		_w16707_,
		_w16705_,
		_w16708_
	);
	LUT3 #(
		.INIT('hb0)
	) name15359 (
		_w7464_,
		_w7465_,
		_w16708_,
		_w16709_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15360 (
		\P3_InstAddrPointer_reg[20]/NET0131 ,
		\P3_rEIP_reg[20]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16710_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15361 (
		_w1945_,
		_w16703_,
		_w16709_,
		_w16710_,
		_w16711_
	);
	LUT3 #(
		.INIT('h08)
	) name15362 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16712_
	);
	LUT4 #(
		.INIT('haa20)
	) name15363 (
		_w1810_,
		_w8731_,
		_w8733_,
		_w16712_,
		_w16713_
	);
	LUT2 #(
		.INIT('h1)
	) name15364 (
		_w1833_,
		_w3357_,
		_w16714_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15365 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16714_,
		_w16715_
	);
	LUT2 #(
		.INIT('h4)
	) name15366 (
		_w1862_,
		_w3267_,
		_w16716_
	);
	LUT3 #(
		.INIT('h40)
	) name15367 (
		_w1833_,
		_w1846_,
		_w8735_,
		_w16717_
	);
	LUT4 #(
		.INIT('h004f)
	) name15368 (
		_w1816_,
		_w1831_,
		_w3211_,
		_w16717_,
		_w16718_
	);
	LUT4 #(
		.INIT('h0100)
	) name15369 (
		_w8736_,
		_w16715_,
		_w16716_,
		_w16718_,
		_w16719_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15370 (
		\P1_InstAddrPointer_reg[9]/NET0131 ,
		\P1_rEIP_reg[9]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16720_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15371 (
		_w1933_,
		_w16713_,
		_w16719_,
		_w16720_,
		_w16721_
	);
	LUT3 #(
		.INIT('h08)
	) name15372 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16722_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15373 (
		\P2_InstAddrPointer_reg[26]/NET0131 ,
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w1640_,
		_w4424_,
		_w16723_
	);
	LUT4 #(
		.INIT('h1033)
	) name15374 (
		_w1602_,
		_w1606_,
		_w1616_,
		_w6440_,
		_w16724_
	);
	LUT3 #(
		.INIT('h04)
	) name15375 (
		_w1625_,
		_w1643_,
		_w1667_,
		_w16725_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15376 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		_w6446_,
		_w16724_,
		_w16725_,
		_w16726_
	);
	LUT3 #(
		.INIT('hb0)
	) name15377 (
		_w1571_,
		_w1583_,
		_w4363_,
		_w16727_
	);
	LUT4 #(
		.INIT('h40cc)
	) name15378 (
		_w1602_,
		_w1606_,
		_w1616_,
		_w6440_,
		_w16728_
	);
	LUT3 #(
		.INIT('hc8)
	) name15379 (
		_w1563_,
		_w4274_,
		_w16728_,
		_w16729_
	);
	LUT4 #(
		.INIT('h0001)
	) name15380 (
		_w16723_,
		_w16727_,
		_w16729_,
		_w16726_,
		_w16730_
	);
	LUT4 #(
		.INIT('hd700)
	) name15381 (
		_w1659_,
		_w4426_,
		_w5716_,
		_w16730_,
		_w16731_
	);
	LUT4 #(
		.INIT('h5700)
	) name15382 (
		_w1559_,
		_w6873_,
		_w16722_,
		_w16731_,
		_w16732_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15383 (
		\P2_InstAddrPointer_reg[27]/NET0131 ,
		\P2_rEIP_reg[27]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16733_
	);
	LUT3 #(
		.INIT('h2f)
	) name15384 (
		_w1678_,
		_w16732_,
		_w16733_,
		_w16734_
	);
	LUT3 #(
		.INIT('h02)
	) name15385 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16735_
	);
	LUT3 #(
		.INIT('ha8)
	) name15386 (
		_w2171_,
		_w7991_,
		_w16735_,
		_w16736_
	);
	LUT3 #(
		.INIT('he0)
	) name15387 (
		_w2071_,
		_w2087_,
		_w7993_,
		_w16737_
	);
	LUT4 #(
		.INIT('h0002)
	) name15388 (
		_w2126_,
		_w2127_,
		_w2175_,
		_w16737_,
		_w16738_
	);
	LUT3 #(
		.INIT('hb0)
	) name15389 (
		_w2073_,
		_w2086_,
		_w2886_,
		_w16739_
	);
	LUT4 #(
		.INIT('he000)
	) name15390 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7993_,
		_w16740_
	);
	LUT3 #(
		.INIT('h0b)
	) name15391 (
		_w2117_,
		_w2955_,
		_w16740_,
		_w16741_
	);
	LUT4 #(
		.INIT('h0d00)
	) name15392 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		_w16738_,
		_w16739_,
		_w16741_,
		_w16742_
	);
	LUT2 #(
		.INIT('h4)
	) name15393 (
		_w7996_,
		_w16742_,
		_w16743_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15394 (
		\P3_InstAddrPointer_reg[16]/NET0131 ,
		\P3_rEIP_reg[16]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16744_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15395 (
		_w1945_,
		_w16736_,
		_w16743_,
		_w16744_,
		_w16745_
	);
	LUT3 #(
		.INIT('h02)
	) name15396 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16746_
	);
	LUT4 #(
		.INIT('haa20)
	) name15397 (
		_w2171_,
		_w6951_,
		_w6952_,
		_w16746_,
		_w16747_
	);
	LUT4 #(
		.INIT('he000)
	) name15398 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w3042_,
		_w16748_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15399 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16749_
	);
	LUT3 #(
		.INIT('hb0)
	) name15400 (
		_w2073_,
		_w2086_,
		_w2728_,
		_w16750_
	);
	LUT2 #(
		.INIT('h4)
	) name15401 (
		_w2117_,
		_w2975_,
		_w16751_
	);
	LUT4 #(
		.INIT('h0001)
	) name15402 (
		_w16750_,
		_w16751_,
		_w16749_,
		_w16748_,
		_w16752_
	);
	LUT4 #(
		.INIT('hd700)
	) name15403 (
		_w2181_,
		_w3042_,
		_w6948_,
		_w16752_,
		_w16753_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15404 (
		\P3_InstAddrPointer_reg[27]/NET0131 ,
		\P3_rEIP_reg[27]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16754_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15405 (
		_w1945_,
		_w16747_,
		_w16753_,
		_w16754_,
		_w16755_
	);
	LUT3 #(
		.INIT('h08)
	) name15406 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16756_
	);
	LUT4 #(
		.INIT('haa20)
	) name15407 (
		_w1559_,
		_w6889_,
		_w6892_,
		_w16756_,
		_w16757_
	);
	LUT3 #(
		.INIT('h54)
	) name15408 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w1592_,
		_w1595_,
		_w16758_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15409 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w16758_,
		_w16759_
	);
	LUT3 #(
		.INIT('h60)
	) name15410 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4425_,
		_w16759_,
		_w16760_
	);
	LUT3 #(
		.INIT('h2a)
	) name15411 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		_w4844_,
		_w5429_,
		_w16761_
	);
	LUT2 #(
		.INIT('h4)
	) name15412 (
		_w1617_,
		_w6890_,
		_w16762_
	);
	LUT3 #(
		.INIT('hb0)
	) name15413 (
		_w1571_,
		_w1583_,
		_w4365_,
		_w16763_
	);
	LUT4 #(
		.INIT('h0001)
	) name15414 (
		_w16762_,
		_w16760_,
		_w16763_,
		_w16761_,
		_w16764_
	);
	LUT4 #(
		.INIT('hd700)
	) name15415 (
		_w1659_,
		_w6895_,
		_w6905_,
		_w16764_,
		_w16765_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15416 (
		\P2_InstAddrPointer_reg[28]/NET0131 ,
		\P2_rEIP_reg[28]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16766_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15417 (
		_w1678_,
		_w16757_,
		_w16765_,
		_w16766_,
		_w16767_
	);
	LUT3 #(
		.INIT('h08)
	) name15418 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16768_
	);
	LUT4 #(
		.INIT('haa20)
	) name15419 (
		_w1810_,
		_w8154_,
		_w8157_,
		_w16768_,
		_w16769_
	);
	LUT3 #(
		.INIT('h2a)
	) name15420 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		_w1922_,
		_w4037_,
		_w16770_
	);
	LUT3 #(
		.INIT('h40)
	) name15421 (
		_w1833_,
		_w1846_,
		_w3380_,
		_w16771_
	);
	LUT2 #(
		.INIT('h4)
	) name15422 (
		_w1862_,
		_w3317_,
		_w16772_
	);
	LUT3 #(
		.INIT('hb0)
	) name15423 (
		_w1816_,
		_w1831_,
		_w3240_,
		_w16773_
	);
	LUT4 #(
		.INIT('h0001)
	) name15424 (
		_w16772_,
		_w16773_,
		_w16771_,
		_w16770_,
		_w16774_
	);
	LUT3 #(
		.INIT('hb0)
	) name15425 (
		_w8160_,
		_w8161_,
		_w16774_,
		_w16775_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15426 (
		\P1_InstAddrPointer_reg[25]/NET0131 ,
		\P1_rEIP_reg[25]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16776_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15427 (
		_w1933_,
		_w16769_,
		_w16775_,
		_w16776_,
		_w16777_
	);
	LUT3 #(
		.INIT('h08)
	) name15428 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16778_
	);
	LUT4 #(
		.INIT('haa20)
	) name15429 (
		_w1559_,
		_w8236_,
		_w8238_,
		_w16778_,
		_w16779_
	);
	LUT2 #(
		.INIT('h8)
	) name15430 (
		_w1640_,
		_w6898_,
		_w16780_
	);
	LUT3 #(
		.INIT('h0b)
	) name15431 (
		_w1617_,
		_w8233_,
		_w16780_,
		_w16781_
	);
	LUT3 #(
		.INIT('h2a)
	) name15432 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		_w1614_,
		_w1668_,
		_w16782_
	);
	LUT3 #(
		.INIT('hb0)
	) name15433 (
		_w1571_,
		_w1583_,
		_w4336_,
		_w16783_
	);
	LUT3 #(
		.INIT('h10)
	) name15434 (
		_w16782_,
		_w16783_,
		_w16781_,
		_w16784_
	);
	LUT2 #(
		.INIT('h4)
	) name15435 (
		_w8241_,
		_w16784_,
		_w16785_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15436 (
		\P2_InstAddrPointer_reg[16]/NET0131 ,
		\P2_rEIP_reg[16]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16786_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15437 (
		_w1678_,
		_w16779_,
		_w16785_,
		_w16786_,
		_w16787_
	);
	LUT4 #(
		.INIT('h4447)
	) name15438 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2173_,
		_w7487_,
		_w7488_,
		_w16788_
	);
	LUT4 #(
		.INIT('he000)
	) name15439 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7490_,
		_w16789_
	);
	LUT3 #(
		.INIT('h0b)
	) name15440 (
		_w2117_,
		_w4061_,
		_w16789_,
		_w16790_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15441 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16791_
	);
	LUT3 #(
		.INIT('hb0)
	) name15442 (
		_w2073_,
		_w2086_,
		_w2905_,
		_w16792_
	);
	LUT3 #(
		.INIT('h10)
	) name15443 (
		_w16791_,
		_w16792_,
		_w16790_,
		_w16793_
	);
	LUT4 #(
		.INIT('h1f00)
	) name15444 (
		_w7490_,
		_w7491_,
		_w7492_,
		_w16793_,
		_w16794_
	);
	LUT4 #(
		.INIT('h08aa)
	) name15445 (
		_w1945_,
		_w2171_,
		_w16788_,
		_w16794_,
		_w16795_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15446 (
		\P3_InstAddrPointer_reg[24]/NET0131 ,
		\P3_rEIP_reg[24]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16796_
	);
	LUT2 #(
		.INIT('hb)
	) name15447 (
		_w16795_,
		_w16796_,
		_w16797_
	);
	LUT3 #(
		.INIT('h08)
	) name15448 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16798_
	);
	LUT4 #(
		.INIT('h002f)
	) name15449 (
		_w3101_,
		_w7522_,
		_w7523_,
		_w16798_,
		_w16799_
	);
	LUT2 #(
		.INIT('h4)
	) name15450 (
		_w1862_,
		_w3300_,
		_w16800_
	);
	LUT3 #(
		.INIT('ha2)
	) name15451 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16801_
	);
	LUT3 #(
		.INIT('h40)
	) name15452 (
		_w1833_,
		_w1846_,
		_w3362_,
		_w16802_
	);
	LUT4 #(
		.INIT('h004f)
	) name15453 (
		_w1816_,
		_w1831_,
		_w3216_,
		_w16802_,
		_w16803_
	);
	LUT4 #(
		.INIT('h0100)
	) name15454 (
		_w7525_,
		_w16801_,
		_w16800_,
		_w16803_,
		_w16804_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15455 (
		_w1810_,
		_w1933_,
		_w16799_,
		_w16804_,
		_w16805_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15456 (
		\P1_InstAddrPointer_reg[11]/NET0131 ,
		\P1_rEIP_reg[11]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16806_
	);
	LUT2 #(
		.INIT('hb)
	) name15457 (
		_w16805_,
		_w16806_,
		_w16807_
	);
	LUT4 #(
		.INIT('h7774)
	) name15458 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w1916_,
		_w7033_,
		_w7031_,
		_w16808_
	);
	LUT4 #(
		.INIT('h1020)
	) name15459 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w1833_,
		_w1846_,
		_w3387_,
		_w16809_
	);
	LUT3 #(
		.INIT('h2a)
	) name15460 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		_w1922_,
		_w4037_,
		_w16810_
	);
	LUT2 #(
		.INIT('h4)
	) name15461 (
		_w1862_,
		_w7030_,
		_w16811_
	);
	LUT3 #(
		.INIT('hb0)
	) name15462 (
		_w1816_,
		_w1831_,
		_w3258_,
		_w16812_
	);
	LUT4 #(
		.INIT('h0001)
	) name15463 (
		_w16811_,
		_w16812_,
		_w16809_,
		_w16810_,
		_w16813_
	);
	LUT4 #(
		.INIT('h3100)
	) name15464 (
		_w1810_,
		_w7036_,
		_w16808_,
		_w16813_,
		_w16814_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15465 (
		\P1_InstAddrPointer_reg[28]/NET0131 ,
		\P1_rEIP_reg[28]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16815_
	);
	LUT3 #(
		.INIT('h2f)
	) name15466 (
		_w1933_,
		_w16814_,
		_w16815_,
		_w16816_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15467 (
		\P3_EBX_reg[25]/NET0131 ,
		\P3_EBX_reg[26]/NET0131 ,
		_w2084_,
		_w8920_,
		_w16817_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name15468 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2098_,
		_w8414_,
		_w8425_,
		_w16818_
	);
	LUT3 #(
		.INIT('h2a)
	) name15469 (
		\P3_EBX_reg[26]/NET0131 ,
		_w2075_,
		_w2083_,
		_w16819_
	);
	LUT3 #(
		.INIT('h8d)
	) name15470 (
		_w2071_,
		_w16818_,
		_w16819_,
		_w16820_
	);
	LUT2 #(
		.INIT('h2)
	) name15471 (
		\P3_EBX_reg[26]/NET0131 ,
		_w8341_,
		_w16821_
	);
	LUT4 #(
		.INIT('hff8a)
	) name15472 (
		_w1945_,
		_w16817_,
		_w16820_,
		_w16821_,
		_w16822_
	);
	LUT3 #(
		.INIT('h08)
	) name15473 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16823_
	);
	LUT2 #(
		.INIT('h8)
	) name15474 (
		_w1640_,
		_w4913_,
		_w16824_
	);
	LUT2 #(
		.INIT('h4)
	) name15475 (
		_w1617_,
		_w7394_,
		_w16825_
	);
	LUT3 #(
		.INIT('hb0)
	) name15476 (
		_w1571_,
		_w1583_,
		_w4356_,
		_w16826_
	);
	LUT3 #(
		.INIT('h2a)
	) name15477 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		_w1658_,
		_w4844_,
		_w16827_
	);
	LUT4 #(
		.INIT('h0001)
	) name15478 (
		_w16826_,
		_w16824_,
		_w16827_,
		_w16825_,
		_w16828_
	);
	LUT4 #(
		.INIT('hd700)
	) name15479 (
		_w1659_,
		_w4913_,
		_w7400_,
		_w16828_,
		_w16829_
	);
	LUT4 #(
		.INIT('h5700)
	) name15480 (
		_w1559_,
		_w7398_,
		_w16823_,
		_w16829_,
		_w16830_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15481 (
		\P2_InstAddrPointer_reg[24]/NET0131 ,
		\P2_rEIP_reg[24]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16831_
	);
	LUT3 #(
		.INIT('h2f)
	) name15482 (
		_w1678_,
		_w16830_,
		_w16831_,
		_w16832_
	);
	LUT3 #(
		.INIT('h08)
	) name15483 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16833_
	);
	LUT4 #(
		.INIT('haa20)
	) name15484 (
		_w1810_,
		_w8071_,
		_w8072_,
		_w16833_,
		_w16834_
	);
	LUT3 #(
		.INIT('ha2)
	) name15485 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16835_
	);
	LUT2 #(
		.INIT('h4)
	) name15486 (
		_w1862_,
		_w3302_,
		_w16836_
	);
	LUT3 #(
		.INIT('h40)
	) name15487 (
		_w1833_,
		_w1846_,
		_w8074_,
		_w16837_
	);
	LUT4 #(
		.INIT('h004f)
	) name15488 (
		_w1816_,
		_w1831_,
		_w3219_,
		_w16837_,
		_w16838_
	);
	LUT3 #(
		.INIT('h10)
	) name15489 (
		_w16836_,
		_w16835_,
		_w16838_,
		_w16839_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15490 (
		_w1933_,
		_w8076_,
		_w16834_,
		_w16839_,
		_w16840_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15491 (
		\P1_InstAddrPointer_reg[13]/NET0131 ,
		\P1_rEIP_reg[13]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16841_
	);
	LUT2 #(
		.INIT('hb)
	) name15492 (
		_w16840_,
		_w16841_,
		_w16842_
	);
	LUT3 #(
		.INIT('h08)
	) name15493 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16843_
	);
	LUT4 #(
		.INIT('haa20)
	) name15494 (
		_w1810_,
		_w7541_,
		_w7543_,
		_w16843_,
		_w16844_
	);
	LUT2 #(
		.INIT('h1)
	) name15495 (
		_w1833_,
		_w3367_,
		_w16845_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15496 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16845_,
		_w16846_
	);
	LUT2 #(
		.INIT('h4)
	) name15497 (
		_w1862_,
		_w7539_,
		_w16847_
	);
	LUT3 #(
		.INIT('h40)
	) name15498 (
		_w1833_,
		_w1846_,
		_w4026_,
		_w16848_
	);
	LUT4 #(
		.INIT('h004f)
	) name15499 (
		_w1816_,
		_w1831_,
		_w3243_,
		_w16848_,
		_w16849_
	);
	LUT3 #(
		.INIT('h10)
	) name15500 (
		_w16846_,
		_w16847_,
		_w16849_,
		_w16850_
	);
	LUT2 #(
		.INIT('h4)
	) name15501 (
		_w7546_,
		_w16850_,
		_w16851_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15502 (
		\P1_InstAddrPointer_reg[15]/NET0131 ,
		\P1_rEIP_reg[15]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16852_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15503 (
		_w1933_,
		_w16844_,
		_w16851_,
		_w16852_,
		_w16853_
	);
	LUT3 #(
		.INIT('h82)
	) name15504 (
		_w1846_,
		_w9050_,
		_w9061_,
		_w16854_
	);
	LUT2 #(
		.INIT('h8)
	) name15505 (
		_w1814_,
		_w16854_,
		_w16855_
	);
	LUT3 #(
		.INIT('ha8)
	) name15506 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1863_,
		_w8992_,
		_w16856_
	);
	LUT2 #(
		.INIT('h1)
	) name15507 (
		_w16855_,
		_w16856_,
		_w16857_
	);
	LUT4 #(
		.INIT('hb700)
	) name15508 (
		\P1_EBX_reg[27]/NET0131 ,
		_w1829_,
		_w8988_,
		_w16857_,
		_w16858_
	);
	LUT2 #(
		.INIT('h2)
	) name15509 (
		\P1_EBX_reg[27]/NET0131 ,
		_w9102_,
		_w16859_
	);
	LUT3 #(
		.INIT('hf2)
	) name15510 (
		_w1933_,
		_w16858_,
		_w16859_,
		_w16860_
	);
	LUT3 #(
		.INIT('h08)
	) name15511 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16861_
	);
	LUT4 #(
		.INIT('haa20)
	) name15512 (
		_w1559_,
		_w8250_,
		_w8251_,
		_w16861_,
		_w16862_
	);
	LUT3 #(
		.INIT('h65)
	) name15513 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w1605_,
		_w4247_,
		_w16863_
	);
	LUT2 #(
		.INIT('h4)
	) name15514 (
		_w1602_,
		_w16863_,
		_w16864_
	);
	LUT3 #(
		.INIT('h08)
	) name15515 (
		_w1501_,
		_w1568_,
		_w16864_,
		_w16865_
	);
	LUT4 #(
		.INIT('haa8a)
	) name15516 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		_w6446_,
		_w16725_,
		_w16865_,
		_w16866_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15517 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w5424_,
		_w16867_
	);
	LUT2 #(
		.INIT('h8)
	) name15518 (
		_w4413_,
		_w16867_,
		_w16868_
	);
	LUT3 #(
		.INIT('hb0)
	) name15519 (
		_w1571_,
		_w1583_,
		_w4340_,
		_w16869_
	);
	LUT2 #(
		.INIT('h8)
	) name15520 (
		_w1563_,
		_w4251_,
		_w16870_
	);
	LUT4 #(
		.INIT('h0031)
	) name15521 (
		_w1604_,
		_w1602_,
		_w1616_,
		_w16863_,
		_w16871_
	);
	LUT2 #(
		.INIT('h1)
	) name15522 (
		_w16870_,
		_w16871_,
		_w16872_
	);
	LUT4 #(
		.INIT('h0100)
	) name15523 (
		_w16866_,
		_w16869_,
		_w16868_,
		_w16872_,
		_w16873_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name15524 (
		_w1678_,
		_w8255_,
		_w16862_,
		_w16873_,
		_w16874_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15525 (
		\P2_InstAddrPointer_reg[17]/NET0131 ,
		\P2_rEIP_reg[17]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16875_
	);
	LUT2 #(
		.INIT('hb)
	) name15526 (
		_w16874_,
		_w16875_,
		_w16876_
	);
	LUT3 #(
		.INIT('h13)
	) name15527 (
		\P1_EBX_reg[29]/NET0131 ,
		\P1_EBX_reg[30]/NET0131 ,
		_w10523_,
		_w16877_
	);
	LUT2 #(
		.INIT('h2)
	) name15528 (
		_w1829_,
		_w8991_,
		_w16878_
	);
	LUT4 #(
		.INIT('h8008)
	) name15529 (
		_w1814_,
		_w1846_,
		_w9096_,
		_w9085_,
		_w16879_
	);
	LUT3 #(
		.INIT('ha8)
	) name15530 (
		\P1_EBX_reg[30]/NET0131 ,
		_w1863_,
		_w8992_,
		_w16880_
	);
	LUT2 #(
		.INIT('h1)
	) name15531 (
		_w16879_,
		_w16880_,
		_w16881_
	);
	LUT4 #(
		.INIT('h20aa)
	) name15532 (
		_w1933_,
		_w16877_,
		_w16878_,
		_w16881_,
		_w16882_
	);
	LUT2 #(
		.INIT('h2)
	) name15533 (
		\P1_EBX_reg[30]/NET0131 ,
		_w9102_,
		_w16883_
	);
	LUT2 #(
		.INIT('he)
	) name15534 (
		_w16882_,
		_w16883_,
		_w16884_
	);
	LUT2 #(
		.INIT('h2)
	) name15535 (
		\P1_EAX_reg[27]/NET0131 ,
		_w9102_,
		_w16885_
	);
	LUT4 #(
		.INIT('h4888)
	) name15536 (
		\P1_EAX_reg[27]/NET0131 ,
		_w1827_,
		_w9434_,
		_w9476_,
		_w16886_
	);
	LUT3 #(
		.INIT('hd1)
	) name15537 (
		\P1_EAX_reg[27]/NET0131 ,
		_w1867_,
		_w3431_,
		_w16887_
	);
	LUT2 #(
		.INIT('h2)
	) name15538 (
		_w1795_,
		_w16887_,
		_w16888_
	);
	LUT3 #(
		.INIT('hd1)
	) name15539 (
		\P1_EAX_reg[27]/NET0131 ,
		_w1867_,
		_w3526_,
		_w16889_
	);
	LUT3 #(
		.INIT('h08)
	) name15540 (
		_w1725_,
		_w1802_,
		_w16889_,
		_w16890_
	);
	LUT4 #(
		.INIT('h0007)
	) name15541 (
		_w1832_,
		_w16854_,
		_w16888_,
		_w16890_,
		_w16891_
	);
	LUT3 #(
		.INIT('hd0)
	) name15542 (
		\P1_EAX_reg[27]/NET0131 ,
		_w9437_,
		_w16891_,
		_w16892_
	);
	LUT4 #(
		.INIT('hecee)
	) name15543 (
		_w1933_,
		_w16885_,
		_w16886_,
		_w16892_,
		_w16893_
	);
	LUT3 #(
		.INIT('h08)
	) name15544 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w1592_,
		_w1660_,
		_w16894_
	);
	LUT4 #(
		.INIT('h004f)
	) name15545 (
		_w6844_,
		_w6847_,
		_w6851_,
		_w16894_,
		_w16895_
	);
	LUT2 #(
		.INIT('h4)
	) name15546 (
		_w1596_,
		_w4419_,
		_w16896_
	);
	LUT3 #(
		.INIT('h04)
	) name15547 (
		_w1555_,
		_w4912_,
		_w16896_,
		_w16897_
	);
	LUT2 #(
		.INIT('h4)
	) name15548 (
		_w1617_,
		_w6848_,
		_w16898_
	);
	LUT3 #(
		.INIT('h2a)
	) name15549 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		_w1658_,
		_w4844_,
		_w16899_
	);
	LUT3 #(
		.INIT('hb0)
	) name15550 (
		_w1571_,
		_w1583_,
		_w4354_,
		_w16900_
	);
	LUT4 #(
		.INIT('h0001)
	) name15551 (
		_w16899_,
		_w16900_,
		_w16898_,
		_w16897_,
		_w16901_
	);
	LUT2 #(
		.INIT('h4)
	) name15552 (
		_w6854_,
		_w16901_,
		_w16902_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15553 (
		_w1559_,
		_w1678_,
		_w16895_,
		_w16902_,
		_w16903_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15554 (
		\P2_InstAddrPointer_reg[23]/NET0131 ,
		\P2_rEIP_reg[23]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16904_
	);
	LUT2 #(
		.INIT('hb)
	) name15555 (
		_w16903_,
		_w16904_,
		_w16905_
	);
	LUT3 #(
		.INIT('h08)
	) name15556 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16906_
	);
	LUT4 #(
		.INIT('haa20)
	) name15557 (
		_w1810_,
		_w8087_,
		_w8088_,
		_w16906_,
		_w16907_
	);
	LUT2 #(
		.INIT('h4)
	) name15558 (
		_w1862_,
		_w8085_,
		_w16908_
	);
	LUT3 #(
		.INIT('ha2)
	) name15559 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16909_
	);
	LUT3 #(
		.INIT('h40)
	) name15560 (
		_w1833_,
		_w1846_,
		_w3369_,
		_w16910_
	);
	LUT4 #(
		.INIT('h004f)
	) name15561 (
		_w1816_,
		_w1831_,
		_w3254_,
		_w16910_,
		_w16911_
	);
	LUT3 #(
		.INIT('h10)
	) name15562 (
		_w16909_,
		_w16908_,
		_w16911_,
		_w16912_
	);
	LUT2 #(
		.INIT('h4)
	) name15563 (
		_w8090_,
		_w16912_,
		_w16913_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15564 (
		\P1_InstAddrPointer_reg[14]/NET0131 ,
		\P1_rEIP_reg[14]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16914_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15565 (
		_w1933_,
		_w16907_,
		_w16913_,
		_w16914_,
		_w16915_
	);
	LUT3 #(
		.INIT('h08)
	) name15566 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16916_
	);
	LUT4 #(
		.INIT('haa20)
	) name15567 (
		_w1810_,
		_w8137_,
		_w8139_,
		_w16916_,
		_w16917_
	);
	LUT2 #(
		.INIT('h8)
	) name15568 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w4739_,
		_w16918_
	);
	LUT3 #(
		.INIT('hc4)
	) name15569 (
		_w1862_,
		_w3308_,
		_w16918_,
		_w16919_
	);
	LUT3 #(
		.INIT('h40)
	) name15570 (
		_w1833_,
		_w1846_,
		_w8141_,
		_w16920_
	);
	LUT3 #(
		.INIT('hb0)
	) name15571 (
		_w1816_,
		_w1831_,
		_w3235_,
		_w16921_
	);
	LUT3 #(
		.INIT('ha2)
	) name15572 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16922_
	);
	LUT4 #(
		.INIT('h0001)
	) name15573 (
		_w16921_,
		_w16919_,
		_w16922_,
		_w16920_,
		_w16923_
	);
	LUT3 #(
		.INIT('hb0)
	) name15574 (
		_w8142_,
		_w8143_,
		_w16923_,
		_w16924_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15575 (
		\P1_InstAddrPointer_reg[21]/NET0131 ,
		\P1_rEIP_reg[21]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16925_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15576 (
		_w1933_,
		_w16917_,
		_w16924_,
		_w16925_,
		_w16926_
	);
	LUT4 #(
		.INIT('h4447)
	) name15577 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w1661_,
		_w7929_,
		_w7930_,
		_w16927_
	);
	LUT3 #(
		.INIT('h01)
	) name15578 (
		_w1592_,
		_w1595_,
		_w4403_,
		_w16928_
	);
	LUT4 #(
		.INIT('h00c8)
	) name15579 (
		_w1503_,
		_w1549_,
		_w1553_,
		_w16928_,
		_w16929_
	);
	LUT2 #(
		.INIT('h8)
	) name15580 (
		_w1596_,
		_w16929_,
		_w16930_
	);
	LUT4 #(
		.INIT('h004f)
	) name15581 (
		_w1571_,
		_w1583_,
		_w4315_,
		_w16930_,
		_w16931_
	);
	LUT2 #(
		.INIT('h4)
	) name15582 (
		_w1617_,
		_w4223_,
		_w16932_
	);
	LUT3 #(
		.INIT('h07)
	) name15583 (
		_w1605_,
		_w1656_,
		_w16929_,
		_w16933_
	);
	LUT3 #(
		.INIT('h2a)
	) name15584 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		_w4926_,
		_w16933_,
		_w16934_
	);
	LUT4 #(
		.INIT('h0100)
	) name15585 (
		_w7933_,
		_w16932_,
		_w16934_,
		_w16931_,
		_w16935_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15586 (
		_w1559_,
		_w1678_,
		_w16927_,
		_w16935_,
		_w16936_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15587 (
		\P2_InstAddrPointer_reg[8]/NET0131 ,
		\P2_rEIP_reg[8]/NET0131 ,
		_w2286_,
		_w4441_,
		_w16937_
	);
	LUT2 #(
		.INIT('hb)
	) name15588 (
		_w16936_,
		_w16937_,
		_w16938_
	);
	LUT3 #(
		.INIT('h08)
	) name15589 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16939_
	);
	LUT4 #(
		.INIT('h004f)
	) name15590 (
		_w7591_,
		_w7592_,
		_w7593_,
		_w16939_,
		_w16940_
	);
	LUT3 #(
		.INIT('ha2)
	) name15591 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w4037_,
		_w4741_,
		_w16941_
	);
	LUT3 #(
		.INIT('h40)
	) name15592 (
		_w1833_,
		_w1846_,
		_w3382_,
		_w16942_
	);
	LUT3 #(
		.INIT('h80)
	) name15593 (
		_w1805_,
		_w1806_,
		_w3313_,
		_w16943_
	);
	LUT3 #(
		.INIT('h9a)
	) name15594 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		_w1861_,
		_w3230_,
		_w16944_
	);
	LUT4 #(
		.INIT('h010f)
	) name15595 (
		_w1855_,
		_w1860_,
		_w16943_,
		_w16944_,
		_w16945_
	);
	LUT4 #(
		.INIT('h4f00)
	) name15596 (
		_w1816_,
		_w1831_,
		_w3237_,
		_w16945_,
		_w16946_
	);
	LUT3 #(
		.INIT('h10)
	) name15597 (
		_w16941_,
		_w16942_,
		_w16946_,
		_w16947_
	);
	LUT4 #(
		.INIT('hd700)
	) name15598 (
		_w1924_,
		_w3377_,
		_w3382_,
		_w16947_,
		_w16948_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15599 (
		_w1810_,
		_w1933_,
		_w16940_,
		_w16948_,
		_w16949_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15600 (
		\P1_InstAddrPointer_reg[22]/NET0131 ,
		\P1_rEIP_reg[22]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16950_
	);
	LUT2 #(
		.INIT('hb)
	) name15601 (
		_w16949_,
		_w16950_,
		_w16951_
	);
	LUT3 #(
		.INIT('h02)
	) name15602 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16952_
	);
	LUT4 #(
		.INIT('h002f)
	) name15603 (
		_w2755_,
		_w7425_,
		_w7426_,
		_w16952_,
		_w16953_
	);
	LUT2 #(
		.INIT('h2)
	) name15604 (
		_w2171_,
		_w16953_,
		_w16954_
	);
	LUT4 #(
		.INIT('he000)
	) name15605 (
		_w2071_,
		_w2087_,
		_w2098_,
		_w7420_,
		_w16955_
	);
	LUT3 #(
		.INIT('h0b)
	) name15606 (
		_w2117_,
		_w2950_,
		_w16955_,
		_w16956_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15607 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		_w2126_,
		_w2127_,
		_w2175_,
		_w16957_
	);
	LUT3 #(
		.INIT('hb0)
	) name15608 (
		_w2073_,
		_w2086_,
		_w2876_,
		_w16958_
	);
	LUT3 #(
		.INIT('h10)
	) name15609 (
		_w16957_,
		_w16958_,
		_w16956_,
		_w16959_
	);
	LUT3 #(
		.INIT('hb0)
	) name15610 (
		_w7419_,
		_w7421_,
		_w16959_,
		_w16960_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15611 (
		\P3_InstAddrPointer_reg[11]/NET0131 ,
		\P3_rEIP_reg[11]/NET0131 ,
		_w3054_,
		_w3056_,
		_w16961_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15612 (
		_w1945_,
		_w16954_,
		_w16960_,
		_w16961_,
		_w16962_
	);
	LUT4 #(
		.INIT('h8000)
	) name15613 (
		_w2069_,
		_w2070_,
		_w2098_,
		_w12537_,
		_w16963_
	);
	LUT4 #(
		.INIT('h00fd)
	) name15614 (
		\P3_EBX_reg[25]/NET0131 ,
		_w8923_,
		_w8924_,
		_w16963_,
		_w16964_
	);
	LUT4 #(
		.INIT('hb700)
	) name15615 (
		\P3_EBX_reg[25]/NET0131 ,
		_w2084_,
		_w8920_,
		_w16964_,
		_w16965_
	);
	LUT2 #(
		.INIT('h2)
	) name15616 (
		\P3_EBX_reg[25]/NET0131 ,
		_w8341_,
		_w16966_
	);
	LUT3 #(
		.INIT('hf2)
	) name15617 (
		_w1945_,
		_w16965_,
		_w16966_,
		_w16967_
	);
	LUT3 #(
		.INIT('h08)
	) name15618 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16968_
	);
	LUT4 #(
		.INIT('haa20)
	) name15619 (
		_w1810_,
		_w7559_,
		_w7561_,
		_w16968_,
		_w16969_
	);
	LUT2 #(
		.INIT('h4)
	) name15620 (
		_w1862_,
		_w4450_,
		_w16970_
	);
	LUT3 #(
		.INIT('ha2)
	) name15621 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16971_
	);
	LUT3 #(
		.INIT('h40)
	) name15622 (
		_w1833_,
		_w1846_,
		_w3374_,
		_w16972_
	);
	LUT4 #(
		.INIT('h004f)
	) name15623 (
		_w1816_,
		_w1831_,
		_w3250_,
		_w16972_,
		_w16973_
	);
	LUT3 #(
		.INIT('h10)
	) name15624 (
		_w16971_,
		_w16970_,
		_w16973_,
		_w16974_
	);
	LUT3 #(
		.INIT('hb0)
	) name15625 (
		_w7563_,
		_w7564_,
		_w16974_,
		_w16975_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15626 (
		\P1_InstAddrPointer_reg[19]/NET0131 ,
		\P1_rEIP_reg[19]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16976_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15627 (
		_w1933_,
		_w16969_,
		_w16975_,
		_w16976_,
		_w16977_
	);
	LUT3 #(
		.INIT('h08)
	) name15628 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16978_
	);
	LUT3 #(
		.INIT('ha8)
	) name15629 (
		_w1810_,
		_w8102_,
		_w16978_,
		_w16979_
	);
	LUT2 #(
		.INIT('h4)
	) name15630 (
		_w1862_,
		_w3297_,
		_w16980_
	);
	LUT3 #(
		.INIT('ha2)
	) name15631 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		_w1914_,
		_w1868_,
		_w16981_
	);
	LUT3 #(
		.INIT('h40)
	) name15632 (
		_w1833_,
		_w1846_,
		_w3368_,
		_w16982_
	);
	LUT4 #(
		.INIT('h004f)
	) name15633 (
		_w1816_,
		_w1831_,
		_w3246_,
		_w16982_,
		_w16983_
	);
	LUT3 #(
		.INIT('h10)
	) name15634 (
		_w16981_,
		_w16980_,
		_w16983_,
		_w16984_
	);
	LUT2 #(
		.INIT('h4)
	) name15635 (
		_w8103_,
		_w16984_,
		_w16985_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15636 (
		\P1_InstAddrPointer_reg[16]/NET0131 ,
		\P1_rEIP_reg[16]/NET0131 ,
		_w3406_,
		_w3408_,
		_w16986_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15637 (
		_w1933_,
		_w16979_,
		_w16985_,
		_w16986_,
		_w16987_
	);
	LUT3 #(
		.INIT('h08)
	) name15638 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w1842_,
		_w1915_,
		_w16988_
	);
	LUT4 #(
		.INIT('h028a)
	) name15639 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w1809_,
		_w1810_,
		_w1846_,
		_w16989_
	);
	LUT4 #(
		.INIT('h007d)
	) name15640 (
		_w1924_,
		_w16638_,
		_w16639_,
		_w16989_,
		_w16990_
	);
	LUT4 #(
		.INIT('h5700)
	) name15641 (
		_w1810_,
		_w16637_,
		_w16988_,
		_w16990_,
		_w16991_
	);
	LUT3 #(
		.INIT('h60)
	) name15642 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w6376_,
		_w6378_,
		_w16992_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15643 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		\P1_rEIP_reg[31]/NET0131 ,
		_w3406_,
		_w6383_,
		_w16993_
	);
	LUT4 #(
		.INIT('hb700)
	) name15644 (
		\P1_PhyAddrPointer_reg[31]/NET0131 ,
		_w2310_,
		_w6381_,
		_w16993_,
		_w16994_
	);
	LUT2 #(
		.INIT('h4)
	) name15645 (
		_w16992_,
		_w16994_,
		_w16995_
	);
	LUT3 #(
		.INIT('h2f)
	) name15646 (
		_w1933_,
		_w16991_,
		_w16995_,
		_w16996_
	);
	LUT3 #(
		.INIT('h02)
	) name15647 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2103_,
		_w2172_,
		_w16997_
	);
	LUT4 #(
		.INIT('haa20)
	) name15648 (
		_w2171_,
		_w16661_,
		_w16663_,
		_w16997_,
		_w16998_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name15649 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w16999_
	);
	LUT4 #(
		.INIT('h00d7)
	) name15650 (
		_w2181_,
		_w3025_,
		_w3027_,
		_w16999_,
		_w17000_
	);
	LUT3 #(
		.INIT('h02)
	) name15651 (
		_w3055_,
		_w8018_,
		_w11938_,
		_w17001_
	);
	LUT3 #(
		.INIT('h15)
	) name15652 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w5765_,
		_w7447_,
		_w17002_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name15653 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		_w2194_,
		_w5766_,
		_w6938_,
		_w17003_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15654 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_rEIP_reg[17]/NET0131 ,
		_w3054_,
		_w5783_,
		_w17004_
	);
	LUT3 #(
		.INIT('hb0)
	) name15655 (
		_w17002_,
		_w17003_,
		_w17004_,
		_w17005_
	);
	LUT2 #(
		.INIT('h4)
	) name15656 (
		_w17001_,
		_w17005_,
		_w17006_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15657 (
		_w1945_,
		_w16998_,
		_w17000_,
		_w17006_,
		_w17007_
	);
	LUT3 #(
		.INIT('h08)
	) name15658 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w1842_,
		_w1915_,
		_w17008_
	);
	LUT3 #(
		.INIT('ha8)
	) name15659 (
		_w1810_,
		_w8716_,
		_w17008_,
		_w17009_
	);
	LUT2 #(
		.INIT('h1)
	) name15660 (
		_w1833_,
		_w3347_,
		_w17010_
	);
	LUT4 #(
		.INIT('haaa2)
	) name15661 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		_w1914_,
		_w1868_,
		_w17010_,
		_w17011_
	);
	LUT2 #(
		.INIT('h4)
	) name15662 (
		_w1862_,
		_w3269_,
		_w17012_
	);
	LUT3 #(
		.INIT('h40)
	) name15663 (
		_w1833_,
		_w1846_,
		_w3348_,
		_w17013_
	);
	LUT4 #(
		.INIT('h004f)
	) name15664 (
		_w1816_,
		_w1831_,
		_w3102_,
		_w17013_,
		_w17014_
	);
	LUT4 #(
		.INIT('h0100)
	) name15665 (
		_w8720_,
		_w17012_,
		_w17011_,
		_w17014_,
		_w17015_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15666 (
		\P1_InstAddrPointer_reg[7]/NET0131 ,
		\P1_rEIP_reg[7]/NET0131 ,
		_w3406_,
		_w3408_,
		_w17016_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15667 (
		_w1933_,
		_w17009_,
		_w17015_,
		_w17016_,
		_w17017_
	);
	LUT2 #(
		.INIT('h2)
	) name15668 (
		\P2_EBX_reg[30]/NET0131 ,
		_w7767_,
		_w17018_
	);
	LUT2 #(
		.INIT('h2)
	) name15669 (
		\P2_EBX_reg[30]/NET0131 ,
		_w8961_,
		_w17019_
	);
	LUT4 #(
		.INIT('h8008)
	) name15670 (
		_w1550_,
		_w1596_,
		_w7885_,
		_w7896_,
		_w17020_
	);
	LUT2 #(
		.INIT('h1)
	) name15671 (
		_w17019_,
		_w17020_,
		_w17021_
	);
	LUT4 #(
		.INIT('hb700)
	) name15672 (
		\P2_EBX_reg[30]/NET0131 ,
		_w1578_,
		_w8966_,
		_w17021_,
		_w17022_
	);
	LUT3 #(
		.INIT('hce)
	) name15673 (
		_w1678_,
		_w17018_,
		_w17022_,
		_w17023_
	);
	LUT4 #(
		.INIT('h8000)
	) name15674 (
		\P1_EAX_reg[28]/NET0131 ,
		\P1_EAX_reg[29]/NET0131 ,
		\P1_EAX_reg[30]/NET0131 ,
		_w9655_,
		_w17024_
	);
	LUT3 #(
		.INIT('h48)
	) name15675 (
		\P1_EAX_reg[30]/NET0131 ,
		_w1827_,
		_w9656_,
		_w17025_
	);
	LUT4 #(
		.INIT('h8008)
	) name15676 (
		_w1832_,
		_w1846_,
		_w9096_,
		_w9085_,
		_w17026_
	);
	LUT2 #(
		.INIT('h2)
	) name15677 (
		_w1795_,
		_w3457_,
		_w17027_
	);
	LUT3 #(
		.INIT('h08)
	) name15678 (
		_w1725_,
		_w1802_,
		_w4506_,
		_w17028_
	);
	LUT3 #(
		.INIT('ha8)
	) name15679 (
		_w1867_,
		_w17027_,
		_w17028_,
		_w17029_
	);
	LUT4 #(
		.INIT('h0075)
	) name15680 (
		\P1_EAX_reg[30]/NET0131 ,
		_w9436_,
		_w9437_,
		_w17029_,
		_w17030_
	);
	LUT2 #(
		.INIT('h4)
	) name15681 (
		_w17026_,
		_w17030_,
		_w17031_
	);
	LUT2 #(
		.INIT('h2)
	) name15682 (
		\P1_EAX_reg[30]/NET0131 ,
		_w9102_,
		_w17032_
	);
	LUT4 #(
		.INIT('hff8a)
	) name15683 (
		_w1933_,
		_w17025_,
		_w17031_,
		_w17032_,
		_w17033_
	);
	LUT4 #(
		.INIT('h4447)
	) name15684 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w1916_,
		_w8174_,
		_w8176_,
		_w17034_
	);
	LUT2 #(
		.INIT('h4)
	) name15685 (
		_w1862_,
		_w3268_,
		_w17035_
	);
	LUT3 #(
		.INIT('ha2)
	) name15686 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		_w1914_,
		_w1868_,
		_w17036_
	);
	LUT3 #(
		.INIT('h40)
	) name15687 (
		_w1833_,
		_w1846_,
		_w3358_,
		_w17037_
	);
	LUT4 #(
		.INIT('h004f)
	) name15688 (
		_w1816_,
		_w1831_,
		_w3210_,
		_w17037_,
		_w17038_
	);
	LUT4 #(
		.INIT('h0100)
	) name15689 (
		_w8178_,
		_w17036_,
		_w17035_,
		_w17038_,
		_w17039_
	);
	LUT4 #(
		.INIT('h08cc)
	) name15690 (
		_w1810_,
		_w1933_,
		_w17034_,
		_w17039_,
		_w17040_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15691 (
		\P1_InstAddrPointer_reg[8]/NET0131 ,
		\P1_rEIP_reg[8]/NET0131 ,
		_w3406_,
		_w3408_,
		_w17041_
	);
	LUT2 #(
		.INIT('hb)
	) name15692 (
		_w17040_,
		_w17041_,
		_w17042_
	);
	LUT2 #(
		.INIT('h2)
	) name15693 (
		\P2_uWord_reg[13]/NET0131 ,
		_w7767_,
		_w17043_
	);
	LUT2 #(
		.INIT('h8)
	) name15694 (
		_w1565_,
		_w10359_,
		_w17044_
	);
	LUT3 #(
		.INIT('h0d)
	) name15695 (
		\P2_uWord_reg[13]/NET0131 ,
		_w9467_,
		_w17044_,
		_w17045_
	);
	LUT4 #(
		.INIT('hf8fa)
	) name15696 (
		_w1678_,
		_w14865_,
		_w17043_,
		_w17045_,
		_w17046_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name15697 (
		\P2_EAX_reg[7]/NET0131 ,
		_w1678_,
		_w7767_,
		_w7792_,
		_w17047_
	);
	LUT3 #(
		.INIT('h80)
	) name15698 (
		_w1549_,
		_w1553_,
		_w14361_,
		_w17048_
	);
	LUT2 #(
		.INIT('h6)
	) name15699 (
		\P2_EAX_reg[7]/NET0131 ,
		_w7770_,
		_w17049_
	);
	LUT2 #(
		.INIT('h8)
	) name15700 (
		_w7789_,
		_w17049_,
		_w17050_
	);
	LUT4 #(
		.INIT('h000b)
	) name15701 (
		_w2295_,
		_w8812_,
		_w17048_,
		_w17050_,
		_w17051_
	);
	LUT2 #(
		.INIT('h2)
	) name15702 (
		_w1678_,
		_w17051_,
		_w17052_
	);
	LUT2 #(
		.INIT('he)
	) name15703 (
		_w17047_,
		_w17052_,
		_w17053_
	);
	LUT3 #(
		.INIT('h6a)
	) name15704 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2098_,
		_w2984_,
		_w17054_
	);
	LUT3 #(
		.INIT('he0)
	) name15705 (
		_w2071_,
		_w2087_,
		_w17054_,
		_w17055_
	);
	LUT3 #(
		.INIT('h01)
	) name15706 (
		_w9354_,
		_w9358_,
		_w17055_,
		_w17056_
	);
	LUT3 #(
		.INIT('hb0)
	) name15707 (
		_w2073_,
		_w2086_,
		_w2825_,
		_w17057_
	);
	LUT4 #(
		.INIT('h0002)
	) name15708 (
		_w2122_,
		_w2125_,
		_w2174_,
		_w2175_,
		_w17058_
	);
	LUT4 #(
		.INIT('hed45)
	) name15709 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		_w2117_,
		_w2713_,
		_w17058_,
		_w17059_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name15710 (
		_w1945_,
		_w17057_,
		_w17056_,
		_w17059_,
		_w17060_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15711 (
		\P3_InstAddrPointer_reg[4]/NET0131 ,
		\P3_rEIP_reg[4]/NET0131 ,
		_w3054_,
		_w3056_,
		_w17061_
	);
	LUT2 #(
		.INIT('hb)
	) name15712 (
		_w17060_,
		_w17061_,
		_w17062_
	);
	LUT3 #(
		.INIT('h02)
	) name15713 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2103_,
		_w2172_,
		_w17063_
	);
	LUT4 #(
		.INIT('haa20)
	) name15714 (
		_w2171_,
		_w16589_,
		_w16591_,
		_w17063_,
		_w17064_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name15715 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w2060_,
		_w2041_,
		_w2098_,
		_w17065_
	);
	LUT3 #(
		.INIT('h0b)
	) name15716 (
		_w16585_,
		_w16586_,
		_w17065_,
		_w17066_
	);
	LUT4 #(
		.INIT('h5051)
	) name15717 (
		\P3_DataWidth_reg[1]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w7467_,
		_w8019_,
		_w17067_
	);
	LUT4 #(
		.INIT('h78f0)
	) name15718 (
		\P3_PhyAddrPointer_reg[17]/NET0131 ,
		\P3_PhyAddrPointer_reg[18]/NET0131 ,
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w5766_,
		_w17068_
	);
	LUT3 #(
		.INIT('hc4)
	) name15719 (
		\P3_DataWidth_reg[1]/NET0131 ,
		_w2194_,
		_w17068_,
		_w17069_
	);
	LUT4 #(
		.INIT('h0c08)
	) name15720 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		_w3055_,
		_w7467_,
		_w8019_,
		_w17070_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15721 (
		\P3_PhyAddrPointer_reg[19]/NET0131 ,
		\P3_rEIP_reg[19]/NET0131 ,
		_w3054_,
		_w5783_,
		_w17071_
	);
	LUT4 #(
		.INIT('h4500)
	) name15722 (
		_w17070_,
		_w17067_,
		_w17069_,
		_w17071_,
		_w17072_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15723 (
		_w1945_,
		_w17064_,
		_w17066_,
		_w17072_,
		_w17073_
	);
	LUT2 #(
		.INIT('h2)
	) name15724 (
		\P1_EAX_reg[31]/NET0131 ,
		_w9102_,
		_w17074_
	);
	LUT4 #(
		.INIT('h8000)
	) name15725 (
		_w1725_,
		_w1802_,
		_w1867_,
		_w3425_,
		_w17075_
	);
	LUT4 #(
		.INIT('h007f)
	) name15726 (
		_w1832_,
		_w9085_,
		_w9097_,
		_w17075_,
		_w17076_
	);
	LUT4 #(
		.INIT('h7500)
	) name15727 (
		\P1_EAX_reg[31]/NET0131 ,
		_w9436_,
		_w9437_,
		_w17076_,
		_w17077_
	);
	LUT4 #(
		.INIT('hb700)
	) name15728 (
		\P1_EAX_reg[31]/NET0131 ,
		_w1827_,
		_w17024_,
		_w17077_,
		_w17078_
	);
	LUT3 #(
		.INIT('hce)
	) name15729 (
		_w1933_,
		_w17074_,
		_w17078_,
		_w17079_
	);
	LUT3 #(
		.INIT('h08)
	) name15730 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w1592_,
		_w1660_,
		_w17080_
	);
	LUT4 #(
		.INIT('haa20)
	) name15731 (
		_w1559_,
		_w7904_,
		_w7906_,
		_w17080_,
		_w17081_
	);
	LUT2 #(
		.INIT('h8)
	) name15732 (
		_w1640_,
		_w4418_,
		_w17082_
	);
	LUT4 #(
		.INIT('h00d5)
	) name15733 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		_w1614_,
		_w1668_,
		_w17082_,
		_w17083_
	);
	LUT2 #(
		.INIT('h4)
	) name15734 (
		_w1617_,
		_w4261_,
		_w17084_
	);
	LUT3 #(
		.INIT('hb0)
	) name15735 (
		_w1571_,
		_w1583_,
		_w4349_,
		_w17085_
	);
	LUT3 #(
		.INIT('h10)
	) name15736 (
		_w17084_,
		_w17085_,
		_w17083_,
		_w17086_
	);
	LUT2 #(
		.INIT('h4)
	) name15737 (
		_w7909_,
		_w17086_,
		_w17087_
	);
	LUT4 #(
		.INIT('h3f15)
	) name15738 (
		\P2_InstAddrPointer_reg[21]/NET0131 ,
		\P2_rEIP_reg[21]/NET0131 ,
		_w2286_,
		_w4441_,
		_w17088_
	);
	LUT4 #(
		.INIT('h8aff)
	) name15739 (
		_w1678_,
		_w17081_,
		_w17087_,
		_w17088_,
		_w17089_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \address2[0]_pad  = _w1352_ ;
	assign \address2[10]_pad  = _w1355_ ;
	assign \address2[11]_pad  = _w1358_ ;
	assign \address2[12]_pad  = _w1361_ ;
	assign \address2[13]_pad  = _w1364_ ;
	assign \address2[14]_pad  = _w1367_ ;
	assign \address2[15]_pad  = _w1370_ ;
	assign \address2[16]_pad  = _w1373_ ;
	assign \address2[17]_pad  = _w1376_ ;
	assign \address2[18]_pad  = _w1379_ ;
	assign \address2[19]_pad  = _w1382_ ;
	assign \address2[1]_pad  = _w1385_ ;
	assign \address2[20]_pad  = _w1388_ ;
	assign \address2[21]_pad  = _w1391_ ;
	assign \address2[22]_pad  = _w1394_ ;
	assign \address2[23]_pad  = _w1397_ ;
	assign \address2[24]_pad  = _w1400_ ;
	assign \address2[25]_pad  = _w1403_ ;
	assign \address2[26]_pad  = _w1406_ ;
	assign \address2[27]_pad  = _w1409_ ;
	assign \address2[28]_pad  = _w1412_ ;
	assign \address2[29]_pad  = _w1415_ ;
	assign \address2[2]_pad  = _w1418_ ;
	assign \address2[3]_pad  = _w1421_ ;
	assign \address2[4]_pad  = _w1424_ ;
	assign \address2[5]_pad  = _w1427_ ;
	assign \address2[6]_pad  = _w1430_ ;
	assign \address2[7]_pad  = _w1433_ ;
	assign \address2[8]_pad  = _w1436_ ;
	assign \address2[9]_pad  = _w1439_ ;
	assign \g133468/_2_  = _w1687_ ;
	assign \g133469/_2_  = _w1944_ ;
	assign \g133470/_2_  = _w2198_ ;
	assign \g133475/_0_  = _w2203_ ;
	assign \g133476/_2_  = _w2214_ ;
	assign \g133515/_0_  = _w2217_ ;
	assign \g133516/_0_  = _w2228_ ;
	assign \g133517/_0_  = _w2239_ ;
	assign \g133518/_0_  = _w2245_ ;
	assign \g133523/_0_  = _w2247_ ;
	assign \g133524/_0_  = _w2249_ ;
	assign \g133528/_0_  = _w2292_ ;
	assign \g133529/_0_  = _w2309_ ;
	assign \g133531/_0_  = _w2314_ ;
	assign \g133532/_0_  = _w2335_ ;
	assign \g133533/_0_  = _w2345_ ;
	assign \g133534/_0_  = _w2359_ ;
	assign \g133535/_0_  = _w2372_ ;
	assign \g133536/_0_  = _w2388_ ;
	assign \g133537/_0_  = _w2398_ ;
	assign \g133538/_0_  = _w2413_ ;
	assign \g133539/_0_  = _w2423_ ;
	assign \g133540/_0_  = _w2437_ ;
	assign \g133541/_0_  = _w2447_ ;
	assign \g133542/_0_  = _w2462_ ;
	assign \g133543/_0_  = _w2472_ ;
	assign \g133544/_0_  = _w2485_ ;
	assign \g133545/_0_  = _w2498_ ;
	assign \g133546/_0_  = _w2514_ ;
	assign \g133547/_0_  = _w2524_ ;
	assign \g133548/_0_  = _w2540_ ;
	assign \g133549/_0_  = _w2550_ ;
	assign \g133550/_0_  = _w2566_ ;
	assign \g133551/_0_  = _w2576_ ;
	assign \g133552/_0_  = _w2592_ ;
	assign \g133553/_0_  = _w2602_ ;
	assign \g133554/_0_  = _w2618_ ;
	assign \g133555/_0_  = _w2628_ ;
	assign \g133556/_0_  = _w2643_ ;
	assign \g133557/_0_  = _w2653_ ;
	assign \g133558/_0_  = _w2667_ ;
	assign \g133559/_0_  = _w2677_ ;
	assign \g133560/_0_  = _w2691_ ;
	assign \g133561/_0_  = _w2701_ ;
	assign \g133566/_0_  = _w3058_ ;
	assign \g133619/_0_  = _w3410_ ;
	assign \g133659/_0_  = _w3549_ ;
	assign \g133660/_0_  = _w3571_ ;
	assign \g133662/_0_  = _w3591_ ;
	assign \g133663/_0_  = _w3607_ ;
	assign \g133664/_0_  = _w3622_ ;
	assign \g133665/_0_  = _w3636_ ;
	assign \g133666/_0_  = _w3649_ ;
	assign \g133667/_0_  = _w3663_ ;
	assign \g133668/_0_  = _w3678_ ;
	assign \g133669/_0_  = _w3694_ ;
	assign \g133670/_0_  = _w3708_ ;
	assign \g133671/_0_  = _w3723_ ;
	assign \g133672/_0_  = _w3738_ ;
	assign \g133673/_0_  = _w3753_ ;
	assign \g133674/_0_  = _w3767_ ;
	assign \g133675/_0_  = _w3780_ ;
	assign \g133676/_0_  = _w3793_ ;
	assign \g133677/_0_  = _w3806_ ;
	assign \g133678/_0_  = _w3819_ ;
	assign \g133679/_0_  = _w3832_ ;
	assign \g133680/_0_  = _w3845_ ;
	assign \g133681/_0_  = _w3858_ ;
	assign \g133682/_0_  = _w3871_ ;
	assign \g133683/_0_  = _w3884_ ;
	assign \g133684/_0_  = _w3897_ ;
	assign \g133685/_0_  = _w3910_ ;
	assign \g133686/_0_  = _w3923_ ;
	assign \g133687/_0_  = _w3936_ ;
	assign \g133688/_0_  = _w3949_ ;
	assign \g133689/_0_  = _w3962_ ;
	assign \g133690/_0_  = _w3975_ ;
	assign \g133691/_0_  = _w3988_ ;
	assign \g133694/_0_  = _w4043_ ;
	assign \g133697/_0_  = _w4103_ ;
	assign \g133702/_0_  = _w4443_ ;
	assign \g133703/_0_  = _w4499_ ;
	assign \g133756/_0_  = _w4519_ ;
	assign \g133792/_0_  = _w4531_ ;
	assign \g133793/_0_  = _w4543_ ;
	assign \g133794/_0_  = _w4555_ ;
	assign \g133796/_0_  = _w4567_ ;
	assign \g133797/_0_  = _w4579_ ;
	assign \g133798/_0_  = _w4591_ ;
	assign \g133799/_0_  = _w4603_ ;
	assign \g133800/_0_  = _w4615_ ;
	assign \g133801/_0_  = _w4627_ ;
	assign \g133802/_0_  = _w4639_ ;
	assign \g133803/_0_  = _w4651_ ;
	assign \g133804/_0_  = _w4663_ ;
	assign \g133806/_0_  = _w4675_ ;
	assign \g133807/_0_  = _w4687_ ;
	assign \g133808/_0_  = _w4699_ ;
	assign \g133812/_0_  = _w4719_ ;
	assign \g133813/_0_  = _w4749_ ;
	assign \g133814/_0_  = _w4770_ ;
	assign \g133817/_0_  = _w4793_ ;
	assign \g133821/_0_  = _w4853_ ;
	assign \g133824/_0_  = _w4894_ ;
	assign \g133826/_0_  = _w4933_ ;
	assign \g133828/_0_  = _w4952_ ;
	assign \g133864/_0_  = _w4965_ ;
	assign \g133865/_0_  = _w4987_ ;
	assign \g133867/_0_  = _w4998_ ;
	assign \g133868/_0_  = _w5009_ ;
	assign \g133869/_0_  = _w5020_ ;
	assign \g133871/_0_  = _w5031_ ;
	assign \g133872/_0_  = _w5042_ ;
	assign \g133873/_0_  = _w5053_ ;
	assign \g133874/_0_  = _w5064_ ;
	assign \g133875/_0_  = _w5075_ ;
	assign \g133876/_0_  = _w5086_ ;
	assign \g133877/_0_  = _w5097_ ;
	assign \g133878/_0_  = _w5108_ ;
	assign \g133879/_0_  = _w5119_ ;
	assign \g133881/_0_  = _w5130_ ;
	assign \g133882/_0_  = _w5141_ ;
	assign \g133883/_0_  = _w5152_ ;
	assign \g133884/_0_  = _w5165_ ;
	assign \g133885/_0_  = _w5178_ ;
	assign \g133886/_0_  = _w5191_ ;
	assign \g133887/_0_  = _w5204_ ;
	assign \g133888/_0_  = _w5217_ ;
	assign \g133889/_0_  = _w5230_ ;
	assign \g133890/_0_  = _w5243_ ;
	assign \g133891/_0_  = _w5256_ ;
	assign \g133892/_0_  = _w5269_ ;
	assign \g133893/_0_  = _w5282_ ;
	assign \g133894/_0_  = _w5295_ ;
	assign \g133895/_0_  = _w5308_ ;
	assign \g133896/_0_  = _w5321_ ;
	assign \g133897/_0_  = _w5334_ ;
	assign \g133898/_0_  = _w5347_ ;
	assign \g133910/_0_  = _w5379_ ;
	assign \g133911/_0_  = _w5400_ ;
	assign \g133912/_0_  = _w5415_ ;
	assign \g133915/_0_  = _w5434_ ;
	assign \g133917/_0_  = _w5449_ ;
	assign \g133929/_0_  = _w5475_ ;
	assign \g134014/_0_  = _w5497_ ;
	assign \g134040/_0_  = _w5510_ ;
	assign \g134041/_0_  = _w5523_ ;
	assign \g134042/_0_  = _w5536_ ;
	assign \g134043/_0_  = _w5549_ ;
	assign \g134044/_0_  = _w5562_ ;
	assign \g134045/_0_  = _w5575_ ;
	assign \g134046/_0_  = _w5588_ ;
	assign \g134047/_0_  = _w5601_ ;
	assign \g134048/_0_  = _w5614_ ;
	assign \g134049/_0_  = _w5627_ ;
	assign \g134050/_0_  = _w5640_ ;
	assign \g134051/_0_  = _w5653_ ;
	assign \g134052/_0_  = _w5666_ ;
	assign \g134053/_0_  = _w5679_ ;
	assign \g134054/_0_  = _w5692_ ;
	assign \g134056/_0_  = _w5751_ ;
	assign \g134059/_0_  = _w5787_ ;
	assign \g134064/_0_  = _w5814_ ;
	assign \g134067/_0_  = _w5832_ ;
	assign \g134068/_0_  = _w5850_ ;
	assign \g134069/_0_  = _w5863_ ;
	assign \g134070/_0_  = _w5884_ ;
	assign \g134071/_0_  = _w5904_ ;
	assign \g134073/_0_  = _w5919_ ;
	assign \g134076/_0_  = _w5939_ ;
	assign \g134131/_0_  = _w5951_ ;
	assign \g134132/_0_  = _w5964_ ;
	assign \g134156/_0_  = _w5975_ ;
	assign \g134157/_0_  = _w5987_ ;
	assign \g134158/_0_  = _w5998_ ;
	assign \g134159/_0_  = _w6010_ ;
	assign \g134163/_0_  = _w6021_ ;
	assign \g134164/_0_  = _w6033_ ;
	assign \g134165/_0_  = _w6044_ ;
	assign \g134166/_0_  = _w6056_ ;
	assign \g134167/_0_  = _w6067_ ;
	assign \g134168/_0_  = _w6079_ ;
	assign \g134169/_0_  = _w6090_ ;
	assign \g134170/_0_  = _w6102_ ;
	assign \g134171/_0_  = _w6113_ ;
	assign \g134172/_0_  = _w6125_ ;
	assign \g134173/_0_  = _w6136_ ;
	assign \g134174/_0_  = _w6148_ ;
	assign \g134176/_0_  = _w6159_ ;
	assign \g134177/_0_  = _w6171_ ;
	assign \g134178/_0_  = _w6182_ ;
	assign \g134179/_0_  = _w6194_ ;
	assign \g134181/_0_  = _w6205_ ;
	assign \g134183/_0_  = _w6217_ ;
	assign \g134184/_0_  = _w6228_ ;
	assign \g134185/_0_  = _w6240_ ;
	assign \g134186/_0_  = _w6251_ ;
	assign \g134187/_0_  = _w6263_ ;
	assign \g134188/_0_  = _w6274_ ;
	assign \g134189/_0_  = _w6286_ ;
	assign \g134190/_0_  = _w6297_ ;
	assign \g134191/_0_  = _w6309_ ;
	assign \g134194/_0_  = _w6331_ ;
	assign \g134202/_0_  = _w6354_ ;
	assign \g134207/_0_  = _w6386_ ;
	assign \g134214/_0_  = _w6402_ ;
	assign \g134216/_0_  = _w6430_ ;
	assign \g134226/_0_  = _w6454_ ;
	assign \g134228/_0_  = _w6479_ ;
	assign \g134360/_0_  = _w6490_ ;
	assign \g134383/_0_  = _w6512_ ;
	assign \g134412/_0_  = _w6521_ ;
	assign \g134413/_0_  = _w6530_ ;
	assign \g134419/_0_  = _w6539_ ;
	assign \g134420/_0_  = _w6548_ ;
	assign \g134421/_0_  = _w6557_ ;
	assign \g134422/_0_  = _w6566_ ;
	assign \g134423/_0_  = _w6575_ ;
	assign \g134424/_0_  = _w6584_ ;
	assign \g134426/_0_  = _w6593_ ;
	assign \g134429/_0_  = _w6602_ ;
	assign \g134431/_0_  = _w6611_ ;
	assign \g134433/_0_  = _w6620_ ;
	assign \g134434/_0_  = _w6629_ ;
	assign \g134435/_0_  = _w6638_ ;
	assign \g134436/_0_  = _w6647_ ;
	assign \g134438/_0_  = _w6660_ ;
	assign \g134439/_0_  = _w6673_ ;
	assign \g134441/_0_  = _w6686_ ;
	assign \g134442/_0_  = _w6699_ ;
	assign \g134443/_0_  = _w6712_ ;
	assign \g134445/_0_  = _w6725_ ;
	assign \g134446/_0_  = _w6738_ ;
	assign \g134447/_0_  = _w6751_ ;
	assign \g134448/_0_  = _w6764_ ;
	assign \g134449/_0_  = _w6777_ ;
	assign \g134450/_0_  = _w6790_ ;
	assign \g134451/_0_  = _w6803_ ;
	assign \g134453/_0_  = _w6816_ ;
	assign \g134454/_0_  = _w6829_ ;
	assign \g134455/_0_  = _w6842_ ;
	assign \g134457/_0_  = _w6865_ ;
	assign \g134458/_0_  = _w6881_ ;
	assign \g134459/_0_  = _w6912_ ;
	assign \g134460/_0_  = _w6924_ ;
	assign \g134469/_0_  = _w6947_ ;
	assign \g134470/_0_  = _w6962_ ;
	assign \g134471/_0_  = _w6972_ ;
	assign \g134472/_0_  = _w6991_ ;
	assign \g134479/_0_  = _w7006_ ;
	assign \g134480/_0_  = _w7029_ ;
	assign \g134481/_0_  = _w7046_ ;
	assign \g134482/_0_  = _w7058_ ;
	assign \g134490/_0_  = _w7080_ ;
	assign \g134491/_0_  = _w7095_ ;
	assign \g134496/_0_  = _w7108_ ;
	assign \g134506/_0_  = _w7125_ ;
	assign \g134508/_0_  = _w7144_ ;
	assign \g134579/_0_  = _w7166_ ;
	assign \g134603/_0_  = _w7179_ ;
	assign \g134604/_0_  = _w7192_ ;
	assign \g134605/_0_  = _w7205_ ;
	assign \g134606/_0_  = _w7218_ ;
	assign \g134607/_0_  = _w7231_ ;
	assign \g134608/_0_  = _w7244_ ;
	assign \g134609/_0_  = _w7257_ ;
	assign \g134610/_0_  = _w7270_ ;
	assign \g134611/_0_  = _w7283_ ;
	assign \g134612/_0_  = _w7296_ ;
	assign \g134613/_0_  = _w7309_ ;
	assign \g134614/_0_  = _w7322_ ;
	assign \g134615/_0_  = _w7335_ ;
	assign \g134616/_0_  = _w7348_ ;
	assign \g134617/_0_  = _w7361_ ;
	assign \g134618/_0_  = _w7378_ ;
	assign \g134619/_0_  = _w7392_ ;
	assign \g134620/_0_  = _w7408_ ;
	assign \g134621/_0_  = _w7418_ ;
	assign \g134632/_0_  = _w7436_ ;
	assign \g134633/_0_  = _w7453_ ;
	assign \g134636/_0_  = _w7476_ ;
	assign \g134637/_0_  = _w7486_ ;
	assign \g134638/_0_  = _w7503_ ;
	assign \g134639/_0_  = _w7520_ ;
	assign \g134645/_0_  = _w7538_ ;
	assign \g134646/_0_  = _w7557_ ;
	assign \g134648/_0_  = _w7578_ ;
	assign \g134649/_0_  = _w7589_ ;
	assign \g134650/_0_  = _w7602_ ;
	assign \g134651/_0_  = _w7612_ ;
	assign \g134652/_0_  = _w7625_ ;
	assign \g134656/_0_  = _w7640_ ;
	assign \g134657/_0_  = _w7650_ ;
	assign \g134658/_0_  = _w7666_ ;
	assign \g134664/_0_  = _w7683_ ;
	assign \g134665/_0_  = _w7698_ ;
	assign \g134671/_0_  = _w7719_ ;
	assign \g134672/_0_  = _w7734_ ;
	assign \g134686/_0_  = _w7750_ ;
	assign \g134687/_0_  = _w7765_ ;
	assign \g134735/_0_  = _w7901_ ;
	assign \g134908/_0_  = _w7917_ ;
	assign \g134909/_0_  = _w7927_ ;
	assign \g134910/_0_  = _w7943_ ;
	assign \g134920/_0_  = _w7954_ ;
	assign \g134921/_0_  = _w7973_ ;
	assign \g134922/_0_  = _w7988_ ;
	assign \g134923/_0_  = _w8007_ ;
	assign \g134925/_0_  = _w8024_ ;
	assign \g134926/_0_  = _w8036_ ;
	assign \g134928/_0_  = _w8048_ ;
	assign \g134929/_0_  = _w8060_ ;
	assign \g134933/_0_  = _w8069_ ;
	assign \g134934/_0_  = _w8083_ ;
	assign \g134935/_0_  = _w8098_ ;
	assign \g134936/_0_  = _w8115_ ;
	assign \g134937/_0_  = _w8124_ ;
	assign \g134938/_0_  = _w8135_ ;
	assign \g134940/_0_  = _w8152_ ;
	assign \g134941/_0_  = _w8171_ ;
	assign \g134943/_0_  = _w8189_ ;
	assign \g134945/_0_  = _w8200_ ;
	assign \g134946/_0_  = _w8215_ ;
	assign \g134947/_0_  = _w8231_ ;
	assign \g134948/_0_  = _w8248_ ;
	assign \g134949/_0_  = _w8264_ ;
	assign \g134950/_0_  = _w8275_ ;
	assign \g134959/_0_  = _w8298_ ;
	assign \g134960/_0_  = _w8316_ ;
	assign \g134961/_0_  = _w8339_ ;
	assign \g134979/_0_  = _w8443_ ;
	assign \g134980/_0_  = _w8458_ ;
	assign \g135054/_0_  = _w8465_ ;
	assign \g135061/_0_  = _w8475_ ;
	assign \g135072/_0_  = _w8481_ ;
	assign \g135100/_0_  = _w8487_ ;
	assign \g135127/_0_  = _w8497_ ;
	assign \g135128/_0_  = _w8507_ ;
	assign \g135129/_0_  = _w8517_ ;
	assign \g135130/_0_  = _w8527_ ;
	assign \g135132/_0_  = _w8537_ ;
	assign \g135133/_0_  = _w8547_ ;
	assign \g135134/_0_  = _w8557_ ;
	assign \g135135/_0_  = _w8567_ ;
	assign \g135136/_0_  = _w8577_ ;
	assign \g135137/_0_  = _w8587_ ;
	assign \g135138/_0_  = _w8597_ ;
	assign \g135139/_0_  = _w8607_ ;
	assign \g135140/_0_  = _w8617_ ;
	assign \g135141/_0_  = _w8627_ ;
	assign \g135142/_0_  = _w8637_ ;
	assign \g135145/_0_  = _w8649_ ;
	assign \g135146/_0_  = _w8661_ ;
	assign \g135151/_0_  = _w8678_ ;
	assign \g135154/_0_  = _w8689_ ;
	assign \g135155/_0_  = _w8700_ ;
	assign \g135158/_0_  = _w8712_ ;
	assign \g135163/_0_  = _w8729_ ;
	assign \g135164/_0_  = _w8745_ ;
	assign \g135165/_0_  = _w8756_ ;
	assign \g135192/_0_  = _w8767_ ;
	assign \g135197/_0_  = _w8786_ ;
	assign \g135217/_0_  = _w8798_ ;
	assign \g135225/_0_  = _w8810_ ;
	assign \g135231/_0_  = _w8832_ ;
	assign \g135272/_0_  = _w8852_ ;
	assign \g135290/_0_  = _w8895_ ;
	assign \g135291/_0_  = _w8905_ ;
	assign \g135293/_0_  = _w8931_ ;
	assign \g135294/_0_  = _w8943_ ;
	assign \g135295/_0_  = _w8965_ ;
	assign \g135296/_0_  = _w8972_ ;
	assign \g135297/_0_  = _w9104_ ;
	assign \g135412/_0_  = _w9125_ ;
	assign \g135437/_0_  = _w9132_ ;
	assign \g135438/_0_  = _w9137_ ;
	assign \g135443/_0_  = _w9150_ ;
	assign \g135444/_0_  = _w9163_ ;
	assign \g135445/_0_  = _w9176_ ;
	assign \g135446/_0_  = _w9189_ ;
	assign \g135447/_0_  = _w9202_ ;
	assign \g135448/_0_  = _w9215_ ;
	assign \g135449/_0_  = _w9228_ ;
	assign \g135450/_0_  = _w9241_ ;
	assign \g135451/_0_  = _w9254_ ;
	assign \g135452/_0_  = _w9267_ ;
	assign \g135454/_0_  = _w9280_ ;
	assign \g135455/_0_  = _w9293_ ;
	assign \g135456/_0_  = _w9306_ ;
	assign \g135457/_0_  = _w9319_ ;
	assign \g135458/_0_  = _w9332_ ;
	assign \g135463/_0_  = _w9344_ ;
	assign \g135466/_0_  = _w9349_ ;
	assign \g135473/_0_  = _w9369_ ;
	assign \g135481/_0_  = _w9381_ ;
	assign \g135497/_0_  = _w9387_ ;
	assign \g135503/_0_  = _w9393_ ;
	assign \g135505/_0_  = _w9398_ ;
	assign \g135506/_0_  = _w9403_ ;
	assign \g135557/_0_  = _w9410_ ;
	assign \g135558/_0_  = _w9416_ ;
	assign \g135569/_0_  = _w9447_ ;
	assign \g135570/_0_  = _w9469_ ;
	assign \g135571/_0_  = _w9491_ ;
	assign \g135572/_0_  = _w9503_ ;
	assign \g135573/_0_  = _w9511_ ;
	assign \g135575/_0_  = _w9527_ ;
	assign \g135578/_0_  = _w9546_ ;
	assign \g135754/_0_  = _w9560_ ;
	assign \g135755/_0_  = _w9571_ ;
	assign \g135756/_0_  = _w9581_ ;
	assign \g135767/_0_  = _w9594_ ;
	assign \g135768/_0_  = _w9607_ ;
	assign \g135769/_0_  = _w9619_ ;
	assign \g135777/_0_  = _w9631_ ;
	assign \g135778/_0_  = _w9643_ ;
	assign \g135779/_0_  = _w9653_ ;
	assign \g135872/_0_  = _w9664_ ;
	assign \g135873/_0_  = _w9675_ ;
	assign \g135875/_0_  = _w9696_ ;
	assign \g135877/_0_  = _w9707_ ;
	assign \g135878/_0_  = _w9712_ ;
	assign \g135879/_0_  = _w9718_ ;
	assign \g135880/_0_  = _w9738_ ;
	assign \g136087/_0_  = _w9750_ ;
	assign \g136118/_0_  = _w9802_ ;
	assign \g136119/_0_  = _w9813_ ;
	assign \g136120/_0_  = _w9824_ ;
	assign \g136121/_0_  = _w9835_ ;
	assign \g136122/_0_  = _w9846_ ;
	assign \g136123/_0_  = _w9857_ ;
	assign \g136124/_0_  = _w9868_ ;
	assign \g136125/_0_  = _w9879_ ;
	assign \g136126/_0_  = _w9890_ ;
	assign \g136127/_0_  = _w9901_ ;
	assign \g136128/_0_  = _w9912_ ;
	assign \g136129/_0_  = _w9923_ ;
	assign \g136130/_0_  = _w9934_ ;
	assign \g136131/_0_  = _w9945_ ;
	assign \g136132/_0_  = _w9956_ ;
	assign \g136133/_0_  = _w9967_ ;
	assign \g136172/_0_  = _w9974_ ;
	assign \g136173/_0_  = _w9980_ ;
	assign \g136174/_0_  = _w9984_ ;
	assign \g136175/_0_  = _w9988_ ;
	assign \g136177/_0_  = _w9998_ ;
	assign \g136178/_0_  = _w10002_ ;
	assign \g136242/_0_  = _w10011_ ;
	assign \g136243/_0_  = _w10015_ ;
	assign \g136244/_0_  = _w10024_ ;
	assign \g136246/_0_  = _w10044_ ;
	assign \g136248/_0_  = _w10052_ ;
	assign \g136249/_0_  = _w10070_ ;
	assign \g136250/_0_  = _w10088_ ;
	assign \g136251/_0_  = _w10105_ ;
	assign \g136252/_0_  = _w10121_ ;
	assign \g136253/_0_  = _w10139_ ;
	assign \g136254/_0_  = _w10147_ ;
	assign \g136255/_0_  = _w10157_ ;
	assign \g136256/_0_  = _w10165_ ;
	assign \g136257/_0_  = _w10171_ ;
	assign \g136258/_0_  = _w10177_ ;
	assign \g136259/_0_  = _w10185_ ;
	assign \g136260/_0_  = _w10191_ ;
	assign \g136261/_0_  = _w10197_ ;
	assign \g136262/_0_  = _w10203_ ;
	assign \g136263/_0_  = _w10209_ ;
	assign \g136264/_0_  = _w10226_ ;
	assign \g136265/_0_  = _w10243_ ;
	assign \g136266/_0_  = _w10251_ ;
	assign \g136267/_0_  = _w10258_ ;
	assign \g136268/_0_  = _w10276_ ;
	assign \g136269/_0_  = _w10294_ ;
	assign \g136270/_0_  = _w10312_ ;
	assign \g136271/_0_  = _w10330_ ;
	assign \g136272/_0_  = _w10338_ ;
	assign \g136273/_0_  = _w10356_ ;
	assign \g136274/_0_  = _w10375_ ;
	assign \g136275/_0_  = _w10394_ ;
	assign \g136276/_0_  = _w10404_ ;
	assign \g136277/_0_  = _w10412_ ;
	assign \g136279/_0_  = _w10420_ ;
	assign \g136280/_0_  = _w10428_ ;
	assign \g136281/_0_  = _w10446_ ;
	assign \g136282/_0_  = _w10454_ ;
	assign \g136283/_0_  = _w10462_ ;
	assign \g136285/_0_  = _w10480_ ;
	assign \g136286/_0_  = _w10502_ ;
	assign \g136287/_0_  = _w10522_ ;
	assign \g136288/_0_  = _w10529_ ;
	assign \g136289/_0_  = _w10535_ ;
	assign \g136290/_0_  = _w10555_ ;
	assign \g136291/_0_  = _w10573_ ;
	assign \g136292/_0_  = _w10593_ ;
	assign \g136293/_0_  = _w10599_ ;
	assign \g136295/_0_  = _w10610_ ;
	assign \g136467/_0_  = _w10628_ ;
	assign \g136468/_0_  = _w10645_ ;
	assign \g136469/_0_  = _w10658_ ;
	assign \g136470/_0_  = _w10669_ ;
	assign \g136472/_0_  = _w10681_ ;
	assign \g136473/_0_  = _w10690_ ;
	assign \g136474/_0_  = _w10700_ ;
	assign \g136476/_0_  = _w10711_ ;
	assign \g136479/_0_  = _w10723_ ;
	assign \g136480/_0_  = _w10733_ ;
	assign \g136481/_0_  = _w10744_ ;
	assign \g136482/_0_  = _w10757_ ;
	assign \g136483/_0_  = _w10768_ ;
	assign \g136484/_0_  = _w10778_ ;
	assign \g136485/_0_  = _w10787_ ;
	assign \g136486/_0_  = _w10799_ ;
	assign \g136528/_0_  = _w10833_ ;
	assign \g136529/_0_  = _w10851_ ;
	assign \g136530/_0_  = _w10873_ ;
	assign \g136531/_0_  = _w10897_ ;
	assign \g136532/_0_  = _w10917_ ;
	assign \g136533/_0_  = _w10942_ ;
	assign \g136534/_0_  = _w10962_ ;
	assign \g136535/_0_  = _w10980_ ;
	assign \g136536/_0_  = _w11000_ ;
	assign \g136537/_0_  = _w11018_ ;
	assign \g136538/_0_  = _w11040_ ;
	assign \g136539/_0_  = _w11058_ ;
	assign \g136540/_0_  = _w11077_ ;
	assign \g136541/_0_  = _w11096_ ;
	assign \g136542/_0_  = _w11116_ ;
	assign \g136543/_0_  = _w11133_ ;
	assign \g136544/_0_  = _w11151_ ;
	assign \g136545/_0_  = _w11173_ ;
	assign \g136546/_0_  = _w11193_ ;
	assign \g136547/_0_  = _w11213_ ;
	assign \g136548/_0_  = _w11233_ ;
	assign \g136549/_0_  = _w11254_ ;
	assign \g136550/_0_  = _w11276_ ;
	assign \g136551/_0_  = _w11292_ ;
	assign \g136552/_0_  = _w11310_ ;
	assign \g136553/_0_  = _w11329_ ;
	assign \g136554/_0_  = _w11352_ ;
	assign \g136555/_0_  = _w11372_ ;
	assign \g136556/_0_  = _w11390_ ;
	assign \g136557/_0_  = _w11407_ ;
	assign \g136558/_0_  = _w11427_ ;
	assign \g136559/_0_  = _w11444_ ;
	assign \g136560/_0_  = _w11461_ ;
	assign \g136561/_0_  = _w11477_ ;
	assign \g136562/_0_  = _w11492_ ;
	assign \g136563/_0_  = _w11512_ ;
	assign \g136564/_0_  = _w11527_ ;
	assign \g136565/_0_  = _w11543_ ;
	assign \g136566/_0_  = _w11561_ ;
	assign \g136567/_0_  = _w11581_ ;
	assign \g136568/_0_  = _w11596_ ;
	assign \g136570/_0_  = _w11615_ ;
	assign \g136571/_0_  = _w11633_ ;
	assign \g136572/_0_  = _w11653_ ;
	assign \g136573/_0_  = _w11670_ ;
	assign \g136574/_0_  = _w11688_ ;
	assign \g136575/_0_  = _w11706_ ;
	assign \g136576/_0_  = _w11725_ ;
	assign \g136577/_0_  = _w11742_ ;
	assign \g136578/_0_  = _w11760_ ;
	assign \g136579/_0_  = _w11777_ ;
	assign \g136580/_0_  = _w11795_ ;
	assign \g136582/_0_  = _w11823_ ;
	assign \g136583/_0_  = _w11843_ ;
	assign \g136584/_0_  = _w11860_ ;
	assign \g136585/_0_  = _w11879_ ;
	assign \g136586/_0_  = _w11897_ ;
	assign \g136587/_0_  = _w11916_ ;
	assign \g136588/_0_  = _w11936_ ;
	assign \g136589/_0_  = _w11960_ ;
	assign \g136590/_0_  = _w11979_ ;
	assign \g136591/_0_  = _w11999_ ;
	assign \g136592/_0_  = _w12019_ ;
	assign \g136593/_0_  = _w12040_ ;
	assign \g136594/_0_  = _w12058_ ;
	assign \g136595/_0_  = _w12077_ ;
	assign \g136596/_0_  = _w12095_ ;
	assign \g136597/_0_  = _w12113_ ;
	assign \g136598/_0_  = _w12135_ ;
	assign \g136599/_0_  = _w12151_ ;
	assign \g136600/_0_  = _w12171_ ;
	assign \g136601/_0_  = _w12189_ ;
	assign \g136602/_0_  = _w12211_ ;
	assign \g136603/_0_  = _w12232_ ;
	assign \g136604/_0_  = _w12253_ ;
	assign \g136605/_0_  = _w12273_ ;
	assign \g136606/_0_  = _w12293_ ;
	assign \g136607/_0_  = _w12311_ ;
	assign \g136609/_0_  = _w12328_ ;
	assign \g136610/_0_  = _w12345_ ;
	assign \g136611/_0_  = _w12363_ ;
	assign \g136616/_0_  = _w12382_ ;
	assign \g136617/_0_  = _w12401_ ;
	assign \g136618/_0_  = _w12420_ ;
	assign \g136619/_0_  = _w12439_ ;
	assign \g136626/_0_  = _w12447_ ;
	assign \g136628/_0_  = _w12458_ ;
	assign \g136646/_0_  = _w12466_ ;
	assign \g136649/_0_  = _w12474_ ;
	assign \g136662/_0_  = _w12481_ ;
	assign \g136666/_0_  = _w12489_ ;
	assign \g136695/_0_  = _w12497_ ;
	assign \g136696/_0_  = _w12502_ ;
	assign \g136699/_0_  = _w12509_ ;
	assign \g136762/_0_  = _w12518_ ;
	assign \g136763/_0_  = _w12526_ ;
	assign \g136764/_0_  = _w12531_ ;
	assign \g136765/_0_  = _w12544_ ;
	assign \g136768/_0_  = _w12558_ ;
	assign \g136769/_0_  = _w12564_ ;
	assign \g137051/_0_  = _w12570_ ;
	assign \g137052/_0_  = _w12576_ ;
	assign \g137053/_0_  = _w12585_ ;
	assign \g137054/_0_  = _w12591_ ;
	assign \g137055/_0_  = _w12601_ ;
	assign \g137056/_0_  = _w12607_ ;
	assign \g137057/_0_  = _w12614_ ;
	assign \g137060/_0_  = _w12620_ ;
	assign \g137061/_0_  = _w12626_ ;
	assign \g137063/_0_  = _w12632_ ;
	assign \g137064/_0_  = _w12638_ ;
	assign \g137065/_0_  = _w12648_ ;
	assign \g137067/_0_  = _w12654_ ;
	assign \g137069/_0_  = _w12661_ ;
	assign \g137072/_0_  = _w12667_ ;
	assign \g137073/_0_  = _w12677_ ;
	assign \g137075/_0_  = _w12681_ ;
	assign \g137111/_0_  = _w12684_ ;
	assign \g137122/_0_  = _w12688_ ;
	assign \g137133/_0_  = _w12695_ ;
	assign \g137134/_0_  = _w12711_ ;
	assign \g137135/_0_  = _w12728_ ;
	assign \g137136/_0_  = _w12747_ ;
	assign \g137137/_0_  = _w12764_ ;
	assign \g137138/_0_  = _w12781_ ;
	assign \g137144/_0_  = _w12790_ ;
	assign \g137145/_0_  = _w12807_ ;
	assign \g137146/_0_  = _w12826_ ;
	assign \g137149/_0_  = _w12839_ ;
	assign \g137234/_0_  = _w12844_ ;
	assign \g137237/_0_  = _w12851_ ;
	assign \g137238/_0_  = _w12858_ ;
	assign \g137294/_0_  = _w12869_ ;
	assign \g137295/_0_  = _w12877_ ;
	assign \g137296/_0_  = _w12885_ ;
	assign \g137297/_0_  = _w12894_ ;
	assign \g137298/_0_  = _w12907_ ;
	assign \g137299/_0_  = _w12915_ ;
	assign \g137300/_0_  = _w12923_ ;
	assign \g137301/_0_  = _w12931_ ;
	assign \g137302/_0_  = _w12935_ ;
	assign \g137303/_0_  = _w12943_ ;
	assign \g137304/_0_  = _w12951_ ;
	assign \g137305/_0_  = _w12959_ ;
	assign \g137306/_0_  = _w12967_ ;
	assign \g137307/_0_  = _w12975_ ;
	assign \g137308/_0_  = _w12984_ ;
	assign \g137309/_0_  = _w12992_ ;
	assign \g137310/_0_  = _w13000_ ;
	assign \g137311/_0_  = _w13008_ ;
	assign \g137312/_0_  = _w13013_ ;
	assign \g137313/_0_  = _w13017_ ;
	assign \g137314/_0_  = _w13028_ ;
	assign \g137315/_0_  = _w13032_ ;
	assign \g137316/_0_  = _w13055_ ;
	assign \g137317/_0_  = _w13077_ ;
	assign \g137318/_0_  = _w13099_ ;
	assign \g137319/_0_  = _w13120_ ;
	assign \g137320/_0_  = _w13139_ ;
	assign \g137321/_0_  = _w13160_ ;
	assign \g137322/_0_  = _w13181_ ;
	assign \g137323/_0_  = _w13194_ ;
	assign \g137324/_0_  = _w13206_ ;
	assign \g137325/_0_  = _w13216_ ;
	assign \g137327/_0_  = _w13218_ ;
	assign \g137328/_0_  = _w13238_ ;
	assign \g137329/_0_  = _w13262_ ;
	assign \g137330/_0_  = _w13285_ ;
	assign \g137331/_0_  = _w13307_ ;
	assign \g137332/_0_  = _w13328_ ;
	assign \g137333/_0_  = _w13348_ ;
	assign \g137334/_0_  = _w13369_ ;
	assign \g137335/_0_  = _w13379_ ;
	assign \g137336/_0_  = _w13389_ ;
	assign \g137337/_0_  = _w13399_ ;
	assign \g137338/_0_  = _w13405_ ;
	assign \g137339/_0_  = _w13410_ ;
	assign \g137340/_0_  = _w13417_ ;
	assign \g137341/_0_  = _w13420_ ;
	assign \g137342/_0_  = _w13423_ ;
	assign \g137343/_0_  = _w13426_ ;
	assign \g137344/_0_  = _w13429_ ;
	assign \g137345/_0_  = _w13449_ ;
	assign \g137346/_0_  = _w13470_ ;
	assign \g137347/_0_  = _w13472_ ;
	assign \g137349/_0_  = _w13494_ ;
	assign \g137350/_0_  = _w13515_ ;
	assign \g137351/_0_  = _w13534_ ;
	assign \g137352/_0_  = _w13553_ ;
	assign \g137353/_0_  = _w13572_ ;
	assign \g137354/_0_  = _w13574_ ;
	assign \g137448/_0_  = _w13579_ ;
	assign \g137483/_0_  = _w13587_ ;
	assign \g137484/_0_  = _w13595_ ;
	assign \g137485/_0_  = _w13603_ ;
	assign \g137486/_0_  = _w13611_ ;
	assign \g137487/_0_  = _w13621_ ;
	assign \g137488/_0_  = _w13631_ ;
	assign \g137491/_0_  = _w13639_ ;
	assign \g137492/_0_  = _w13647_ ;
	assign \g137493/_0_  = _w13657_ ;
	assign \g137494/_0_  = _w13667_ ;
	assign \g137495/_0_  = _w13675_ ;
	assign \g137496/_0_  = _w13683_ ;
	assign \g137497/_0_  = _w13691_ ;
	assign \g137499/_0_  = _w13699_ ;
	assign \g137501/_0_  = _w13707_ ;
	assign \g137502/_0_  = _w13715_ ;
	assign \g137503/_0_  = _w13723_ ;
	assign \g137504/_0_  = _w13731_ ;
	assign \g137505/_0_  = _w13739_ ;
	assign \g137506/_0_  = _w13747_ ;
	assign \g137507/_0_  = _w13755_ ;
	assign \g137508/_0_  = _w13763_ ;
	assign \g137509/_0_  = _w13773_ ;
	assign \g137511/_0_  = _w13783_ ;
	assign \g137512/_0_  = _w13791_ ;
	assign \g137513/_0_  = _w13799_ ;
	assign \g137514/_0_  = _w13807_ ;
	assign \g137515/_0_  = _w13815_ ;
	assign \g137516/_0_  = _w13823_ ;
	assign \g137517/_0_  = _w13831_ ;
	assign \g137519/_0_  = _w13843_ ;
	assign \g137520/_0_  = _w13855_ ;
	assign \g137521/_0_  = _w13858_ ;
	assign \g137524/_0_  = _w13862_ ;
	assign \g137541/_0_  = _w13866_ ;
	assign \g137547/_0_  = _w13869_ ;
	assign \g137554/_0_  = _w13873_ ;
	assign \g137559/_0_  = _w13879_ ;
	assign \g137566/_0_  = _w13885_ ;
	assign \g137571/_0_  = _w13890_ ;
	assign \g137778/_0_  = _w13896_ ;
	assign \g137782/_0_  = _w13900_ ;
	assign \g137783/_0_  = _w13907_ ;
	assign \g137784/_0_  = _w13913_ ;
	assign \g137785/_0_  = _w13919_ ;
	assign \g137786/_0_  = _w13924_ ;
	assign \g137820/_0_  = _w13931_ ;
	assign \g137821/_0_  = _w13939_ ;
	assign \g137822/_0_  = _w13947_ ;
	assign \g137823/_0_  = _w13950_ ;
	assign \g137824/_0_  = _w13955_ ;
	assign \g137825/_0_  = _w13962_ ;
	assign \g137826/_0_  = _w13969_ ;
	assign \g137827/_0_  = _w13976_ ;
	assign \g137828/_0_  = _w13982_ ;
	assign \g137829/_0_  = _w13987_ ;
	assign \g137830/_0_  = _w13992_ ;
	assign \g137831/_0_  = _w13997_ ;
	assign \g137832/_0_  = _w14002_ ;
	assign \g137833/_0_  = _w14009_ ;
	assign \g137834/_0_  = _w14014_ ;
	assign \g137835/_0_  = _w14020_ ;
	assign \g137836/_0_  = _w14026_ ;
	assign \g137837/_0_  = _w14032_ ;
	assign \g137838/_0_  = _w14037_ ;
	assign \g137839/_0_  = _w14043_ ;
	assign \g137840/_0_  = _w14048_ ;
	assign \g137841/_0_  = _w14054_ ;
	assign \g137842/_0_  = _w14061_ ;
	assign \g137843/_0_  = _w14068_ ;
	assign \g137844/_0_  = _w14075_ ;
	assign \g137845/_0_  = _w14082_ ;
	assign \g137846/_0_  = _w14089_ ;
	assign \g137847/_0_  = _w14096_ ;
	assign \g137848/_0_  = _w14103_ ;
	assign \g137849/_0_  = _w14110_ ;
	assign \g137850/_0_  = _w14115_ ;
	assign \g137851/_0_  = _w14122_ ;
	assign \g137852/_0_  = _w14129_ ;
	assign \g137853/_0_  = _w14135_ ;
	assign \g137854/_0_  = _w14142_ ;
	assign \g137855/_0_  = _w14147_ ;
	assign \g137856/_0_  = _w14152_ ;
	assign \g137857/_0_  = _w14157_ ;
	assign \g137858/_0_  = _w14162_ ;
	assign \g137859/_0_  = _w14168_ ;
	assign \g137860/_0_  = _w14173_ ;
	assign \g137861/_0_  = _w14179_ ;
	assign \g137862/_0_  = _w14185_ ;
	assign \g137863/_0_  = _w14192_ ;
	assign \g137864/_0_  = _w14197_ ;
	assign \g137865/_0_  = _w14203_ ;
	assign \g137866/_0_  = _w14208_ ;
	assign \g137867/_0_  = _w14213_ ;
	assign \g137868/_0_  = _w14219_ ;
	assign \g137869/_0_  = _w14225_ ;
	assign \g137870/_0_  = _w14231_ ;
	assign \g137871/_0_  = _w14237_ ;
	assign \g137872/_0_  = _w14243_ ;
	assign \g137873/_0_  = _w14248_ ;
	assign \g137874/_0_  = _w14253_ ;
	assign \g137875/_0_  = _w14260_ ;
	assign \g137876/_0_  = _w14266_ ;
	assign \g137877/_0_  = _w14272_ ;
	assign \g137878/_0_  = _w14277_ ;
	assign \g137879/_0_  = _w14282_ ;
	assign \g137880/_0_  = _w14288_ ;
	assign \g137881/_0_  = _w14293_ ;
	assign \g137882/_0_  = _w14298_ ;
	assign \g137883/_0_  = _w14305_ ;
	assign \g137884/_0_  = _w14312_ ;
	assign \g137885/_0_  = _w14319_ ;
	assign \g137886/_0_  = _w14323_ ;
	assign \g137887/_0_  = _w14329_ ;
	assign \g137888/_0_  = _w14335_ ;
	assign \g137889/_0_  = _w14341_ ;
	assign \g137890/_0_  = _w14347_ ;
	assign \g137891/_0_  = _w14354_ ;
	assign \g137892/_0_  = _w14360_ ;
	assign \g137893/_0_  = _w14367_ ;
	assign \g137894/_0_  = _w14373_ ;
	assign \g137895/_0_  = _w14379_ ;
	assign \g137896/_0_  = _w14386_ ;
	assign \g137897/_0_  = _w14393_ ;
	assign \g137898/_0_  = _w14400_ ;
	assign \g137899/_0_  = _w14407_ ;
	assign \g137900/_0_  = _w14414_ ;
	assign \g137901/_0_  = _w14421_ ;
	assign \g137902/_0_  = _w14427_ ;
	assign \g137903/_0_  = _w14431_ ;
	assign \g138338/_0_  = _w14433_ ;
	assign \g138340/_0_  = _w14435_ ;
	assign \g138341/_0_  = _w14441_ ;
	assign \g138346/_0_  = _w14446_ ;
	assign \g138347/_0_  = _w14453_ ;
	assign \g138375/_0_  = _w14456_ ;
	assign \g138395/_0_  = _w14465_ ;
	assign \g138396/_0_  = _w14474_ ;
	assign \g138397/_0_  = _w14479_ ;
	assign \g138398/_0_  = _w14484_ ;
	assign \g138400/_0_  = _w14488_ ;
	assign \g138401/_0_  = _w14497_ ;
	assign \g138402/_0_  = _w14506_ ;
	assign \g138403/_0_  = _w14511_ ;
	assign \g138404/_0_  = _w14519_ ;
	assign \g138405/_0_  = _w14523_ ;
	assign \g138406/_0_  = _w14528_ ;
	assign \g138407/_0_  = _w14534_ ;
	assign \g138408/_0_  = _w14543_ ;
	assign \g138409/_0_  = _w14550_ ;
	assign \g138410/_0_  = _w14556_ ;
	assign \g138411/_0_  = _w14561_ ;
	assign \g138412/_0_  = _w14566_ ;
	assign \g138419/_0_  = _w14574_ ;
	assign \g138420/_0_  = _w14579_ ;
	assign \g138421/_0_  = _w14586_ ;
	assign \g138422/_0_  = _w14591_ ;
	assign \g138423/_0_  = _w14599_ ;
	assign \g138424/_0_  = _w14607_ ;
	assign \g138425/_0_  = _w14615_ ;
	assign \g138426/_0_  = _w14623_ ;
	assign \g138427/_0_  = _w14630_ ;
	assign \g138428/_0_  = _w14638_ ;
	assign \g138429/_0_  = _w14646_ ;
	assign \g138430/_0_  = _w14654_ ;
	assign \g138431/_0_  = _w14662_ ;
	assign \g138432/_0_  = _w14666_ ;
	assign \g138433/_0_  = _w14670_ ;
	assign \g138434/_0_  = _w14675_ ;
	assign \g138435/_0_  = _w14679_ ;
	assign \g138436/_0_  = _w14684_ ;
	assign \g138437/_0_  = _w14689_ ;
	assign \g138438/_0_  = _w14693_ ;
	assign \g138439/_0_  = _w14697_ ;
	assign \g138440/_0_  = _w14701_ ;
	assign \g138441/_0_  = _w14705_ ;
	assign \g138442/_0_  = _w14710_ ;
	assign \g138443/_0_  = _w14714_ ;
	assign \g138908/_0_  = _w14717_ ;
	assign \g138909/_0_  = _w14720_ ;
	assign \g138910/_0_  = _w14723_ ;
	assign \g138914/_0_  = _w14726_ ;
	assign \g138915/_0_  = _w14729_ ;
	assign \g138917/_0_  = _w14733_ ;
	assign \g138918/_0_  = _w14737_ ;
	assign \g138919/_0_  = _w14741_ ;
	assign \g138920/_0_  = _w14745_ ;
	assign \g138921/_0_  = _w14748_ ;
	assign \g138925/_0_  = _w14752_ ;
	assign \g138926/_0_  = _w14756_ ;
	assign \g138927/_0_  = _w14760_ ;
	assign \g138930/_0_  = _w14763_ ;
	assign \g138931/_0_  = _w14766_ ;
	assign \g138932/_0_  = _w14769_ ;
	assign \g138960/_0_  = _w14772_ ;
	assign \g138962/_0_  = _w14775_ ;
	assign \g139037/_0_  = _w14780_ ;
	assign \g139038/_0_  = _w14784_ ;
	assign \g139040/_0_  = _w14787_ ;
	assign \g139043/_0_  = _w14791_ ;
	assign \g139044/_0_  = _w14794_ ;
	assign \g139045/_0_  = _w14798_ ;
	assign \g139046/_0_  = _w14801_ ;
	assign \g139047/_0_  = _w14805_ ;
	assign \g139048/_0_  = _w14808_ ;
	assign \g139049/_0_  = _w14812_ ;
	assign \g139050/_0_  = _w14815_ ;
	assign \g139051/_0_  = _w14819_ ;
	assign \g139053/_0_  = _w14824_ ;
	assign \g139054/_0_  = _w14828_ ;
	assign \g139055/_0_  = _w14831_ ;
	assign \g139056/_0_  = _w14835_ ;
	assign \g139057/_0_  = _w14839_ ;
	assign \g139058/_0_  = _w14843_ ;
	assign \g139059/_0_  = _w14847_ ;
	assign \g139060/_0_  = _w14853_ ;
	assign \g139062/_0_  = _w14857_ ;
	assign \g139063/_0_  = _w14863_ ;
	assign \g139064/_0_  = _w14868_ ;
	assign \g139099/_0_  = _w14872_ ;
	assign \g139126/_0_  = _w14879_ ;
	assign \g139127/_0_  = _w14884_ ;
	assign \g139128/_0_  = _w14891_ ;
	assign \g139129/_0_  = _w14895_ ;
	assign \g139130/_0_  = _w14902_ ;
	assign \g139131/_0_  = _w14906_ ;
	assign \g139132/_0_  = _w14913_ ;
	assign \g139133/_0_  = _w14920_ ;
	assign \g139134/_0_  = _w14927_ ;
	assign \g139135/_0_  = _w14934_ ;
	assign \g139136/_0_  = _w14941_ ;
	assign \g139137/_0_  = _w14948_ ;
	assign \g139138/_0_  = _w14955_ ;
	assign \g139139/_0_  = _w14962_ ;
	assign \g139140/_0_  = _w14969_ ;
	assign \g139141/_0_  = _w14976_ ;
	assign \g139260/_0_  = _w14984_ ;
	assign \g139263/_0_  = _w14992_ ;
	assign \g139267/_0_  = _w15002_ ;
	assign \g139270/_0_  = _w15010_ ;
	assign \g139273/_0_  = _w15020_ ;
	assign \g139276/_0_  = _w15028_ ;
	assign \g139279/_0_  = _w15036_ ;
	assign \g139283/_0_  = _w15044_ ;
	assign \g139286/_0_  = _w15052_ ;
	assign \g139289/_0_  = _w15060_ ;
	assign \g139292/_0_  = _w15068_ ;
	assign \g139295/_0_  = _w15078_ ;
	assign \g139298/_0_  = _w15086_ ;
	assign \g139302/_0_  = _w15094_ ;
	assign \g139305/_0_  = _w15102_ ;
	assign \g139309/_0_  = _w15114_ ;
	assign \g139871/_0_  = _w15117_ ;
	assign \g139872/_0_  = _w15120_ ;
	assign \g139873/_0_  = _w15123_ ;
	assign \g139874/_0_  = _w15126_ ;
	assign \g139875/_0_  = _w15129_ ;
	assign \g139876/_0_  = _w15132_ ;
	assign \g139877/_0_  = _w15135_ ;
	assign \g139878/_0_  = _w15138_ ;
	assign \g139879/_0_  = _w15141_ ;
	assign \g139880/_0_  = _w15144_ ;
	assign \g139881/_0_  = _w15147_ ;
	assign \g139882/_0_  = _w15150_ ;
	assign \g139883/_0_  = _w15154_ ;
	assign \g139884/_0_  = _w15158_ ;
	assign \g139885/_0_  = _w15162_ ;
	assign \g139886/_0_  = _w15166_ ;
	assign \g139887/_0_  = _w15170_ ;
	assign \g139888/_0_  = _w15174_ ;
	assign \g139889/_0_  = _w15178_ ;
	assign \g139890/_0_  = _w15182_ ;
	assign \g139891/_0_  = _w15186_ ;
	assign \g139892/_0_  = _w15189_ ;
	assign \g139893/_0_  = _w15192_ ;
	assign \g139895/_0_  = _w15195_ ;
	assign \g139896/_0_  = _w15198_ ;
	assign \g139899/_0_  = _w15201_ ;
	assign \g139901/_0_  = _w15204_ ;
	assign \g139902/_0_  = _w15207_ ;
	assign \g139903/_0_  = _w15210_ ;
	assign \g139904/_0_  = _w15213_ ;
	assign \g140285/_0_  = _w15240_ ;
	assign \g140288/_0_  = _w15265_ ;
	assign \g140329/_0_  = _w15289_ ;
	assign \g140774/_0_  = _w15299_ ;
	assign \g140832/_0_  = _w15308_ ;
	assign \g140834/_0_  = _w15316_ ;
	assign \g140836/_0_  = _w15324_ ;
	assign \g140838/_0_  = _w15334_ ;
	assign \g140840/_0_  = _w15342_ ;
	assign \g140842/_0_  = _w15352_ ;
	assign \g140844/_0_  = _w15360_ ;
	assign \g140846/_0_  = _w15368_ ;
	assign \g140847/_0_  = _w15376_ ;
	assign \g140848/_0_  = _w15384_ ;
	assign \g140850/_0_  = _w15392_ ;
	assign \g140851/_0_  = _w15400_ ;
	assign \g140852/_0_  = _w15410_ ;
	assign \g140853/_0_  = _w15418_ ;
	assign \g140855/_0_  = _w15426_ ;
	assign \g140857/_0_  = _w15434_ ;
	assign \g140861/_0_  = _w15446_ ;
	assign \g140923/_0_  = _w15456_ ;
	assign \g141178/_0_  = _w15463_ ;
	assign \g141179/_0_  = _w15469_ ;
	assign \g141180/_0_  = _w15476_ ;
	assign \g141480/_0_  = _w15485_ ;
	assign \g141495/_0_  = _w15494_ ;
	assign \g141497/_0_  = _w15503_ ;
	assign \g141562/_0_  = _w15509_ ;
	assign \g141563/_0_  = _w15514_ ;
	assign \g141564/_0_  = _w15520_ ;
	assign \g141589/_0_  = _w15525_ ;
	assign \g141617/_0_  = _w15531_ ;
	assign \g141618/_0_  = _w15539_ ;
	assign \g141621/_0_  = _w15547_ ;
	assign \g141625/_0_  = _w15557_ ;
	assign \g141626/_0_  = _w15567_ ;
	assign \g141630/_0_  = _w15575_ ;
	assign \g141634/_0_  = _w15585_ ;
	assign \g141638/_0_  = _w15593_ ;
	assign \g141642/_0_  = _w15601_ ;
	assign \g141646/_0_  = _w15609_ ;
	assign \g141649/_0_  = _w15617_ ;
	assign \g141651/_0_  = _w15625_ ;
	assign \g141652/_0_  = _w15633_ ;
	assign \g141655/_0_  = _w15641_ ;
	assign \g141658/_0_  = _w15651_ ;
	assign \g141661/_0_  = _w15659_ ;
	assign \g141663/_0_  = _w15667_ ;
	assign \g141664/_0_  = _w15675_ ;
	assign \g141667/_0_  = _w15683_ ;
	assign \g141671/_0_  = _w15695_ ;
	assign \g141706/_0_  = _w15700_ ;
	assign \g141976/_0_  = _w15705_ ;
	assign \g141977/_0_  = _w15711_ ;
	assign \g141994/_0_  = _w15718_ ;
	assign \g142246/_0_  = _w15723_ ;
	assign \g142247/_0_  = _w15728_ ;
	assign \g142253/_0_  = _w15733_ ;
	assign \g142689/_0_  = _w15741_ ;
	assign \g142693/_0_  = _w15749_ ;
	assign \g142701/_0_  = _w15757_ ;
	assign \g142704/_0_  = _w15767_ ;
	assign \g142707/_0_  = _w15775_ ;
	assign \g142710/_0_  = _w15783_ ;
	assign \g142713/_0_  = _w15791_ ;
	assign \g142714/_0_  = _w15799_ ;
	assign \g142717/_0_  = _w15807_ ;
	assign \g142720/_0_  = _w15817_ ;
	assign \g142723/_0_  = _w15825_ ;
	assign \g142727/_0_  = _w15833_ ;
	assign \g142734/_0_  = _w15845_ ;
	assign \g143080/_0_  = _w15851_ ;
	assign \g143081/_0_  = _w15856_ ;
	assign \g143083/_0_  = _w15865_ ;
	assign \g143149/_0_  = _w15872_ ;
	assign \g143150/_0_  = _w15877_ ;
	assign \g143153/_0_  = _w15883_ ;
	assign \g143752/_0_  = _w15892_ ;
	assign \g143753/_0_  = _w15901_ ;
	assign \g143759/_0_  = _w15909_ ;
	assign \g144242/_0_  = _w15914_ ;
	assign \g144243/_0_  = _w15917_ ;
	assign \g144244/_0_  = _w15923_ ;
	assign \g144245/_0_  = _w15929_ ;
	assign \g144246/_0_  = _w15933_ ;
	assign \g144249/_0_  = _w15937_ ;
	assign \g145699/_0_  = _w15942_ ;
	assign \g145700/_0_  = _w15946_ ;
	assign \g145702/_0_  = _w15952_ ;
	assign \g145756/_0_  = _w15956_ ;
	assign \g145757/_0_  = _w15962_ ;
	assign \g145758/_0_  = _w15969_ ;
	assign \g146850/_0_  = _w15974_ ;
	assign \g146851/_0_  = _w15979_ ;
	assign \g146864/_0_  = _w15984_ ;
	assign \g147277/_0_  = _w15990_ ;
	assign \g147278/_0_  = _w15994_ ;
	assign \g147279/_0_  = _w16000_ ;
	assign \g147304/_0_  = _w16007_ ;
	assign \g147305/_0_  = _w16014_ ;
	assign \g147306/_0_  = _w16019_ ;
	assign \g147338/_3_  = _w16031_ ;
	assign \g147339/_3_  = _w16034_ ;
	assign \g147340/_3_  = _w16037_ ;
	assign \g147341/_3_  = _w16040_ ;
	assign \g147342/_3_  = _w16043_ ;
	assign \g147343/_3_  = _w16046_ ;
	assign \g147344/_3_  = _w16049_ ;
	assign \g147345/_3_  = _w16052_ ;
	assign \g147346/_3_  = _w16055_ ;
	assign \g147347/_3_  = _w16058_ ;
	assign \g147348/_3_  = _w16061_ ;
	assign \g147349/_3_  = _w16064_ ;
	assign \g147350/_3_  = _w16067_ ;
	assign \g147351/_3_  = _w16070_ ;
	assign \g147352/_3_  = _w16073_ ;
	assign \g147353/_3_  = _w16076_ ;
	assign \g147354/_3_  = _w16079_ ;
	assign \g147355/_3_  = _w16082_ ;
	assign \g147356/_3_  = _w16085_ ;
	assign \g147357/_3_  = _w16088_ ;
	assign \g147358/_3_  = _w16091_ ;
	assign \g147359/_3_  = _w16094_ ;
	assign \g147360/_3_  = _w16097_ ;
	assign \g147362/_3_  = _w16100_ ;
	assign \g147363/_3_  = _w16103_ ;
	assign \g147364/_3_  = _w16106_ ;
	assign \g147365/_3_  = _w16109_ ;
	assign \g147366/_3_  = _w16112_ ;
	assign \g147367/_3_  = _w16115_ ;
	assign \g147368/_3_  = _w16118_ ;
	assign \g147369/_3_  = _w16121_ ;
	assign \g148630/_0_  = _w16125_ ;
	assign \g148631/_0_  = _w16131_ ;
	assign \g148676/_0_  = _w16135_ ;
	assign \g148785/_0_  = _w16140_ ;
	assign \g148788/_0_  = _w16145_ ;
	assign \g148789/_0_  = _w16148_ ;
	assign \g148834/_0_  = _w16151_ ;
	assign \g148836/_0_  = _w16155_ ;
	assign \g148838/_0_  = _w16161_ ;
	assign \g149836/_0_  = _w16166_ ;
	assign \g149837/_0_  = _w16173_ ;
	assign \g149838/_0_  = _w16180_ ;
	assign \g150142/_0_  = _w16181_ ;
	assign \g152366/_0_  = _w16185_ ;
	assign \g152367/_0_  = _w16189_ ;
	assign \g152368/_0_  = _w16193_ ;
	assign \g152426/_0_  = _w16198_ ;
	assign \g152427/_0_  = _w16204_ ;
	assign \g152428/_0_  = _w16209_ ;
	assign \g152586/_0_  = _w16213_ ;
	assign \g152587/_0_  = _w16219_ ;
	assign \g152588/_0_  = _w16222_ ;
	assign \g153217/_0_  = _w16024_ ;
	assign \g154117/_0_  = _w16226_ ;
	assign \g154118/_0_  = _w16230_ ;
	assign \g154130/_0_  = _w16235_ ;
	assign \g154269/_0_  = _w16241_ ;
	assign \g154270/_0_  = _w16247_ ;
	assign \g154284/_0_  = _w16252_ ;
	assign \g154682/_0_  = _w16259_ ;
	assign \g155004/_0_  = _w16266_ ;
	assign \g155020/_0_  = _w16270_ ;
	assign \g155121/_0_  = _w16275_ ;
	assign \g155124/_0_  = _w16282_ ;
	assign \g155126/_0_  = _w16287_ ;
	assign \g155228/_0_  = _w16293_ ;
	assign \g155229/_0_  = _w16298_ ;
	assign \g155230/_0_  = _w16303_ ;
	assign \g155326/_0_  = _w16310_ ;
	assign \g155327/_0_  = _w16315_ ;
	assign \g155330/_0_  = _w16320_ ;
	assign \g155353/_0_  = _w16325_ ;
	assign \g155354/_0_  = _w16330_ ;
	assign \g155356/_0_  = _w16335_ ;
	assign \g155602/_0_  = _w16343_ ;
	assign \g155633/_0_  = _w16351_ ;
	assign \g155634/_0_  = _w16360_ ;
	assign \g155699/_0_  = _w16365_ ;
	assign \g155708/_0_  = _w16370_ ;
	assign \g155715/_0_  = _w16375_ ;
	assign \g156008/_0_  = _w16378_ ;
	assign \g156013/_0_  = _w16381_ ;
	assign \g156019/_0_  = _w16384_ ;
	assign \g156352/_0_  = _w16388_ ;
	assign \g156353/_0_  = _w16392_ ;
	assign \g156356/_0_  = _w16396_ ;
	assign \g156359/_0_  = _w16402_ ;
	assign \g156360/_0_  = _w16409_ ;
	assign \g156361/_0_  = _w16414_ ;
	assign \g156464/_0_  = _w16418_ ;
	assign \g156465/_0_  = _w16423_ ;
	assign \g156469/_0_  = _w16427_ ;
	assign \g156777/_0_  = _w16430_ ;
	assign \g156778/_0_  = _w16433_ ;
	assign \g156789/_0_  = _w16436_ ;
	assign \g158956/_0_  = _w16440_ ;
	assign \g158957/_0_  = _w16443_ ;
	assign \g158966/_0_  = _w16446_ ;
	assign \g159429/_1_  = _w16371_ ;
	assign \g159477/_1_  = _w16361_ ;
	assign \g159500/_1_  = _w16366_ ;
	assign \g159681/_0_  = _w16452_ ;
	assign \g159890/_0_  = _w16455_ ;
	assign \g159950/_0_  = _w16458_ ;
	assign \g160246/_0_  = _w16461_ ;
	assign \g160846/_0_  = _w16462_ ;
	assign \g160860/_0_  = _w16463_ ;
	assign \g160961/_0_  = _w16464_ ;
	assign \g160987/_0_  = _w16466_ ;
	assign \g161000/_0_  = _w16467_ ;
	assign \g161005/_0_  = _w16468_ ;
	assign \g161042/_0_  = _w16470_ ;
	assign \g161119/_0_  = _w16471_ ;
	assign \g161143/_0_  = _w16472_ ;
	assign \g161150/_0_  = _w16473_ ;
	assign \g161172/_0_  = _w16474_ ;
	assign \g161207/_0_  = _w16475_ ;
	assign \g161315/_0_  = _w16476_ ;
	assign \g161332/_0_  = _w16477_ ;
	assign \g161421/_0_  = _w16478_ ;
	assign \g161492/_0_  = _w16480_ ;
	assign \g161541/_0_  = _w16481_ ;
	assign \g161623/_0_  = _w16482_ ;
	assign \g161655/_0_  = _w16483_ ;
	assign \g161678/_0_  = _w16484_ ;
	assign \g161709/_0_  = _w16485_ ;
	assign \g161737/_0_  = _w16486_ ;
	assign \g161751/_0_  = _w16487_ ;
	assign \g161756/_0_  = _w16488_ ;
	assign \g162016/_0_  = _w16491_ ;
	assign \g162020/_0_  = _w16494_ ;
	assign \g162024/_0_  = _w16497_ ;
	assign \g163326/_0_  = _w16448_ ;
	assign \g163326/_3_  = _w16447_ ;
	assign \g174072/_1_  = _w15241_ ;
	assign \g174360/_1_  = _w15214_ ;
	assign \g174391/_0_  = _w15266_ ;
	assign \g180307/_0_  = _w16507_ ;
	assign \g180335/_0_  = _w16520_ ;
	assign \g180369/_0_  = _w16531_ ;
	assign \g180385/_0_  = _w16541_ ;
	assign \g180395/_0_  = _w16551_ ;
	assign \g180442/_0_  = _w16561_ ;
	assign \g180453/_0_  = _w16571_ ;
	assign \g180524/_0_  = _w16583_ ;
	assign \g180586/_0_  = _w16600_ ;
	assign \g180596/_0_  = _w16611_ ;
	assign \g180606/_0_  = _w16620_ ;
	assign \g180654/_0_  = _w16630_ ;
	assign \g180715/_0_  = _w16649_ ;
	assign \g180805/_0_  = _w16659_ ;
	assign \g180836/_0_  = _w16673_ ;
	assign \g180929/_0_  = _w16687_ ;
	assign \g180944/_0_  = _w16691_ ;
	assign \g180975/_0_  = _w16701_ ;
	assign \g181036/_0_  = _w16711_ ;
	assign \g181072/_0_  = _w16721_ ;
	assign \g181083/_0_  = _w16734_ ;
	assign \g181093/_0_  = _w16745_ ;
	assign \g181127/_0_  = _w16755_ ;
	assign \g181137/_0_  = _w16767_ ;
	assign \g181150/_0_  = _w16777_ ;
	assign \g181160/_0_  = _w16787_ ;
	assign \g181180/_0_  = _w16797_ ;
	assign \g181191/_0_  = _w16807_ ;
	assign \g181238/_0_  = _w16816_ ;
	assign \g181262/_0_  = _w16822_ ;
	assign \g181270/_0_  = _w16832_ ;
	assign \g181280/_0_  = _w16842_ ;
	assign \g181315/_0_  = _w16853_ ;
	assign \g181366/_0_  = _w16860_ ;
	assign \g181385/_0_  = _w16876_ ;
	assign \g181458/_0_  = _w16884_ ;
	assign \g181464/_0_  = _w16893_ ;
	assign \g181478/_0_  = _w16905_ ;
	assign \g181522/_0_  = _w16915_ ;
	assign \g181537/_0_  = _w16926_ ;
	assign \g181584/_0_  = _w16938_ ;
	assign \g181669/_0_  = _w16951_ ;
	assign \g181681/_0_  = _w16962_ ;
	assign \g181719/_0_  = _w16967_ ;
	assign \g181778/_0_  = _w16977_ ;
	assign \g181840/_0_  = _w16987_ ;
	assign \g181936/_0_  = _w16996_ ;
	assign \g181986/_0_  = _w17007_ ;
	assign \g182000/_0_  = _w17017_ ;
	assign \g182083/_0_  = _w17023_ ;
	assign \g182179/_0_  = _w17033_ ;
	assign \g182201/_0_  = _w17042_ ;
	assign \g182227/_0_  = _w17046_ ;
	assign \g182316/_0_  = _w17053_ ;
	assign \g182358/_0_  = _w17062_ ;
	assign \g182473/_0_  = _w17073_ ;
	assign \g182678/_0_  = _w17079_ ;
	assign \g53/_0_  = _w17089_ ;
endmodule;