module top (\ahb_mst0_hsizeo_reg[0]/NET0131 , \ahb_mst0_hsizeo_reg[1]/NET0131 , \ahb_mst0_hsizeo_reg[2]/NET0131 , \ahb_mst0_m0_m1_diff_tx_reg/NET0131 , \ahb_mst0_mx_cmd_st_reg[0]/NET0131 , \ahb_mst0_mx_cmd_st_reg[1]/NET0131 , \ahb_mst0_mx_dtp_reg/NET0131 , \ahb_mst1_mx_cmd_st_reg[0]/NET0131 , \ahb_mst1_mx_cmd_st_reg[1]/NET0131 , \ahb_mst1_mx_dtp_reg/NET0131 , \ahb_slv_br_st_reg[0]/NET0131 , \ahb_slv_br_st_reg[1]/NET0131 , \ahb_slv_br_st_reg[2]/NET0131 , \ahb_slv_slv_ad_d1o_reg[2]/NET0131 , \ahb_slv_slv_ad_d1o_reg[3]/NET0131 , \ahb_slv_slv_ad_d1o_reg[4]/NET0131 , \ahb_slv_slv_ad_d1o_reg[5]/NET0131 , \ahb_slv_slv_ad_d1o_reg[6]/NET0131 , \ahb_slv_slv_ad_d1o_reg[7]/NET0131 , \ahb_slv_slv_ad_d1o_reg[8]/NET0131 , \ahb_slv_slv_br_req_reg/NET0131 , \ahb_slv_slv_pt_d1o_reg[0]/NET0131 , \ahb_slv_slv_pt_d1o_reg[1]/NET0131 , \ahb_slv_slv_pt_d1o_reg[2]/NET0131 , \ahb_slv_slv_pt_d1o_reg[3]/NET0131 , \ahb_slv_slv_sz_d1o_reg[0]/NET0131 , \ahb_slv_slv_sz_d1o_reg[1]/NET0131 , \ahb_slv_slv_sz_d1o_reg[2]/NET0131 , \ahb_slv_slv_wr_d1o_reg/NET0131 , \ch_sel_arb_ch_sel_reg[0]/P0000_reg_syn_2 , \ch_sel_arb_ch_sel_reg[1]/P0000_reg_syn_2 , \ch_sel_arb_ch_sel_reg[2]/P0000_reg_syn_2 , \ch_sel_arb_chcsr_reg_reg[10]/NET0131 , \ch_sel_arb_chcsr_reg_reg[11]/NET0131 , \ch_sel_arb_chcsr_reg_reg[12]/NET0131 , \ch_sel_arb_chcsr_reg_reg[13]/NET0131 , \ch_sel_arb_chcsr_reg_reg[15]/NET0131 , \ch_sel_arb_chcsr_reg_reg[16]/NET0131 , \ch_sel_arb_chcsr_reg_reg[17]/NET0131 , \ch_sel_arb_chcsr_reg_reg[18]/NET0131 , \ch_sel_arb_chcsr_reg_reg[19]/NET0131 , \ch_sel_arb_chcsr_reg_reg[1]/NET0131 , \ch_sel_arb_chcsr_reg_reg[20]/NET0131 , \ch_sel_arb_chcsr_reg_reg[2]/NET0131 , \ch_sel_arb_chcsr_reg_reg[3]/NET0131 , \ch_sel_arb_chcsr_reg_reg[4]/NET0131 , \ch_sel_arb_chcsr_reg_reg[5]/NET0131 , \ch_sel_arb_chcsr_reg_reg[6]/NET0131 , \ch_sel_arb_chcsr_reg_reg[8]/NET0131 , \ch_sel_arb_chcsr_reg_reg[9]/NET0131 , \ch_sel_arb_req_reg/NET0131 , \ch_sel_de_stup_d1_reg/NET0131 , \ch_sel_dma_reqd1_reg[0]/NET0131 , \ch_sel_dma_reqd1_reg[1]/NET0131 , \ch_sel_dma_reqd1_reg[2]/NET0131 , \ch_sel_dma_reqd1_reg[3]/NET0131 , \ch_sel_dma_reqd1_reg[4]/NET0131 , \ch_sel_dma_reqd1_reg[5]/NET0131 , \ch_sel_dma_reqd1_reg[6]/NET0131 , \ch_sel_dma_reqd1_reg[7]/NET0131 , \ch_sel_dma_reqd2_reg[0]/NET0131 , \ch_sel_dma_reqd2_reg[1]/P0001 , \ch_sel_dma_reqd2_reg[2]/P0001 , \ch_sel_dma_reqd2_reg[3]/P0001 , \ch_sel_dma_reqd2_reg[4]/NET0131 , \ch_sel_dma_reqd2_reg[5]/NET0131 , \ch_sel_dma_reqd2_reg[6]/NET0131 , \ch_sel_dma_reqd2_reg[7]/NET0131 , \ch_sel_dma_rrarb0_state_reg[0]/NET0131 , \ch_sel_dma_rrarb0_state_reg[1]/NET0131 , \ch_sel_dma_rrarb0_state_reg[2]/NET0131 , \ch_sel_dma_rrarb1_state_reg[0]/NET0131 , \ch_sel_dma_rrarb1_state_reg[1]/NET0131 , \ch_sel_dma_rrarb1_state_reg[2]/NET0131 , \ch_sel_dma_rrarb2_state_reg[0]/NET0131 , \ch_sel_dma_rrarb2_state_reg[1]/NET0131 , \ch_sel_dma_rrarb2_state_reg[2]/NET0131 , \ch_sel_dma_rrarb3_state_reg[0]/NET0131 , \ch_sel_dma_rrarb3_state_reg[1]/NET0131 , \ch_sel_dma_rrarb3_state_reg[2]/NET0131 , \ch_sel_fix_pri_sel_reg[0]/NET0131 , \ch_sel_fix_pri_sel_reg[1]/NET0131 , \ch_sel_vld_req_any_d1_reg/NET0131 , \ctl_rf_abt_reg[0]/NET0131 , \ctl_rf_abt_reg[1]/NET0131 , \ctl_rf_abt_reg[2]/NET0131 , \ctl_rf_abt_reg[3]/NET0131 , \ctl_rf_abt_reg[4]/NET0131 , \ctl_rf_abt_reg[5]/NET0131 , \ctl_rf_abt_reg[6]/NET0131 , \ctl_rf_abt_reg[7]/NET0131 , \ctl_rf_be_d1_reg[0]/P0001 , \ctl_rf_be_d1_reg[1]/P0001 , \ctl_rf_be_d1_reg[2]/P0001 , \ctl_rf_be_d1_reg[3]/P0001 , \ctl_rf_c0_rf_autold_reg/NET0131 , \ctl_rf_c0_rf_ch_en_reg/NET0131 , \ctl_rf_c0_rf_chabt_reg/NET0131 , \ctl_rf_c0_rf_chdad_reg[0]/NET0131 , \ctl_rf_c0_rf_chdad_reg[10]/P0002 , \ctl_rf_c0_rf_chdad_reg[11]/NET0131 , \ctl_rf_c0_rf_chdad_reg[12]/NET0131 , \ctl_rf_c0_rf_chdad_reg[13]/P0002 , \ctl_rf_c0_rf_chdad_reg[14]/NET0131 , \ctl_rf_c0_rf_chdad_reg[15]/NET0131 , \ctl_rf_c0_rf_chdad_reg[16]/NET0131 , \ctl_rf_c0_rf_chdad_reg[17]/NET0131 , \ctl_rf_c0_rf_chdad_reg[18]/NET0131 , \ctl_rf_c0_rf_chdad_reg[19]/NET0131 , \ctl_rf_c0_rf_chdad_reg[1]/NET0131 , \ctl_rf_c0_rf_chdad_reg[20]/P0002 , \ctl_rf_c0_rf_chdad_reg[21]/P0002 , \ctl_rf_c0_rf_chdad_reg[22]/P0002 , \ctl_rf_c0_rf_chdad_reg[23]/P0002 , \ctl_rf_c0_rf_chdad_reg[24]/P0002 , \ctl_rf_c0_rf_chdad_reg[25]/P0002 , \ctl_rf_c0_rf_chdad_reg[26]/P0002 , \ctl_rf_c0_rf_chdad_reg[27]/P0002 , \ctl_rf_c0_rf_chdad_reg[28]/P0002 , \ctl_rf_c0_rf_chdad_reg[29]/P0002 , \ctl_rf_c0_rf_chdad_reg[2]/NET0131 , \ctl_rf_c0_rf_chdad_reg[30]/P0002 , \ctl_rf_c0_rf_chdad_reg[31]/P0002 , \ctl_rf_c0_rf_chdad_reg[3]/P0002 , \ctl_rf_c0_rf_chdad_reg[4]/P0002 , \ctl_rf_c0_rf_chdad_reg[5]/P0002 , \ctl_rf_c0_rf_chdad_reg[6]/P0002 , \ctl_rf_c0_rf_chdad_reg[7]/P0002 , \ctl_rf_c0_rf_chdad_reg[8]/NET0131 , \ctl_rf_c0_rf_chdad_reg[9]/P0002 , \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c0_rf_chllp_on_reg/NET0131 , \ctl_rf_c0_rf_chllp_reg[0]/P0002 , \ctl_rf_c0_rf_chllp_reg[10]/NET0131 , \ctl_rf_c0_rf_chllp_reg[11]/NET0131 , \ctl_rf_c0_rf_chllp_reg[12]/NET0131 , \ctl_rf_c0_rf_chllp_reg[13]/NET0131 , \ctl_rf_c0_rf_chllp_reg[14]/NET0131 , \ctl_rf_c0_rf_chllp_reg[15]/NET0131 , \ctl_rf_c0_rf_chllp_reg[16]/NET0131 , \ctl_rf_c0_rf_chllp_reg[17]/NET0131 , \ctl_rf_c0_rf_chllp_reg[18]/NET0131 , \ctl_rf_c0_rf_chllp_reg[19]/NET0131 , \ctl_rf_c0_rf_chllp_reg[1]/P0002 , \ctl_rf_c0_rf_chllp_reg[20]/NET0131 , \ctl_rf_c0_rf_chllp_reg[21]/NET0131 , \ctl_rf_c0_rf_chllp_reg[22]/NET0131 , \ctl_rf_c0_rf_chllp_reg[23]/NET0131 , \ctl_rf_c0_rf_chllp_reg[24]/NET0131 , \ctl_rf_c0_rf_chllp_reg[25]/NET0131 , \ctl_rf_c0_rf_chllp_reg[26]/NET0131 , \ctl_rf_c0_rf_chllp_reg[27]/NET0131 , \ctl_rf_c0_rf_chllp_reg[28]/NET0131 , \ctl_rf_c0_rf_chllp_reg[29]/NET0131 , \ctl_rf_c0_rf_chllp_reg[2]/NET0131 , \ctl_rf_c0_rf_chllp_reg[30]/NET0131 , \ctl_rf_c0_rf_chllp_reg[31]/NET0131 , \ctl_rf_c0_rf_chllp_reg[3]/NET0131 , \ctl_rf_c0_rf_chllp_reg[4]/NET0131 , \ctl_rf_c0_rf_chllp_reg[5]/NET0131 , \ctl_rf_c0_rf_chllp_reg[6]/NET0131 , \ctl_rf_c0_rf_chllp_reg[7]/NET0131 , \ctl_rf_c0_rf_chllp_reg[8]/NET0131 , \ctl_rf_c0_rf_chllp_reg[9]/NET0131 , \ctl_rf_c0_rf_chllpen_reg/NET0131 , \ctl_rf_c0_rf_chpri_reg[0]/NET0131 , \ctl_rf_c0_rf_chpri_reg[1]/NET0131 , \ctl_rf_c0_rf_chsad_reg[0]/NET0131 , \ctl_rf_c0_rf_chsad_reg[10]/NET0131 , \ctl_rf_c0_rf_chsad_reg[11]/P0002 , \ctl_rf_c0_rf_chsad_reg[12]/P0002 , \ctl_rf_c0_rf_chsad_reg[13]/NET0131 , \ctl_rf_c0_rf_chsad_reg[14]/P0002 , \ctl_rf_c0_rf_chsad_reg[15]/P0002 , \ctl_rf_c0_rf_chsad_reg[16]/NET0131 , \ctl_rf_c0_rf_chsad_reg[17]/NET0131 , \ctl_rf_c0_rf_chsad_reg[18]/NET0131 , \ctl_rf_c0_rf_chsad_reg[19]/NET0131 , \ctl_rf_c0_rf_chsad_reg[1]/NET0131 , \ctl_rf_c0_rf_chsad_reg[20]/NET0131 , \ctl_rf_c0_rf_chsad_reg[21]/NET0131 , \ctl_rf_c0_rf_chsad_reg[22]/NET0131 , \ctl_rf_c0_rf_chsad_reg[23]/NET0131 , \ctl_rf_c0_rf_chsad_reg[24]/NET0131 , \ctl_rf_c0_rf_chsad_reg[25]/P0002 , \ctl_rf_c0_rf_chsad_reg[26]/P0002 , \ctl_rf_c0_rf_chsad_reg[27]/P0002 , \ctl_rf_c0_rf_chsad_reg[28]/P0002 , \ctl_rf_c0_rf_chsad_reg[29]/P0002 , \ctl_rf_c0_rf_chsad_reg[2]/NET0131 , \ctl_rf_c0_rf_chsad_reg[30]/P0002 , \ctl_rf_c0_rf_chsad_reg[31]/NET0131 , \ctl_rf_c0_rf_chsad_reg[3]/NET0131 , \ctl_rf_c0_rf_chsad_reg[4]/NET0131 , \ctl_rf_c0_rf_chsad_reg[5]/NET0131 , \ctl_rf_c0_rf_chsad_reg[6]/NET0131 , \ctl_rf_c0_rf_chsad_reg[7]/NET0131 , \ctl_rf_c0_rf_chsad_reg[8]/P0002 , \ctl_rf_c0_rf_chsad_reg[9]/NET0131 , \ctl_rf_c0_rf_chtsz_reg[0]/P0002 , \ctl_rf_c0_rf_chtsz_reg[10]/P0002 , \ctl_rf_c0_rf_chtsz_reg[11]/P0002 , \ctl_rf_c0_rf_chtsz_reg[1]/P0002 , \ctl_rf_c0_rf_chtsz_reg[2]/P0002 , \ctl_rf_c0_rf_chtsz_reg[3]/P0002 , \ctl_rf_c0_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c0_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c0_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c0_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c0_rf_chtsz_reg[8]/P0002 , \ctl_rf_c0_rf_chtsz_reg[9]/P0002 , \ctl_rf_c0_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c0_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c0_rf_dreqmode_reg/NET0131 , \ctl_rf_c0_rf_dst_sel_reg/NET0131 , \ctl_rf_c0_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c0_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c0_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c0_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c0_rf_int_err_msk_reg/NET0131 , \ctl_rf_c0_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c0_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c0_rf_mode_reg/NET0131 , \ctl_rf_c0_rf_prot1_reg/NET0131 , \ctl_rf_c0_rf_prot2_reg/NET0131 , \ctl_rf_c0_rf_prot3_reg/NET0131 , \ctl_rf_c0_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c0_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c0_rf_src_sel_reg/NET0131 , \ctl_rf_c0_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c0_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c0_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c0_rf_swidth_reg[0]/NET0131 , \ctl_rf_c0_rf_swidth_reg[1]/NET0131 , \ctl_rf_c0_rf_swidth_reg[2]/NET0131 , \ctl_rf_c0brbs_reg[16]/NET0131 , \ctl_rf_c0brbs_reg[17]/NET0131 , \ctl_rf_c0brbs_reg[18]/NET0131 , \ctl_rf_c0brbs_reg[19]/NET0131 , \ctl_rf_c0brbs_reg[20]/NET0131 , \ctl_rf_c0brbs_reg[21]/NET0131 , \ctl_rf_c0brbs_reg[22]/NET0131 , \ctl_rf_c0brbs_reg[23]/NET0131 , \ctl_rf_c0brbs_reg[24]/NET0131 , \ctl_rf_c0brbs_reg[25]/NET0131 , \ctl_rf_c0brbs_reg[26]/NET0131 , \ctl_rf_c0brbs_reg[27]/NET0131 , \ctl_rf_c0brbs_reg[28]/NET0131 , \ctl_rf_c0brbs_reg[29]/NET0131 , \ctl_rf_c0brbs_reg[30]/NET0131 , \ctl_rf_c0brbs_reg[31]/NET0131 , \ctl_rf_c0dmabs_reg[16]/NET0131 , \ctl_rf_c0dmabs_reg[17]/NET0131 , \ctl_rf_c0dmabs_reg[18]/NET0131 , \ctl_rf_c0dmabs_reg[19]/NET0131 , \ctl_rf_c0dmabs_reg[20]/NET0131 , \ctl_rf_c0dmabs_reg[21]/NET0131 , \ctl_rf_c0dmabs_reg[22]/NET0131 , \ctl_rf_c0dmabs_reg[23]/NET0131 , \ctl_rf_c0dmabs_reg[24]/NET0131 , \ctl_rf_c0dmabs_reg[25]/NET0131 , \ctl_rf_c0dmabs_reg[26]/NET0131 , \ctl_rf_c0dmabs_reg[27]/NET0131 , \ctl_rf_c0dmabs_reg[28]/NET0131 , \ctl_rf_c0dmabs_reg[29]/NET0131 , \ctl_rf_c0dmabs_reg[30]/NET0131 , \ctl_rf_c0dmabs_reg[31]/NET0131 , \ctl_rf_c1_rf_autold_reg/NET0131 , \ctl_rf_c1_rf_ch_en_reg/NET0131 , \ctl_rf_c1_rf_chabt_reg/NET0131 , \ctl_rf_c1_rf_chdad_reg[0]/NET0131 , \ctl_rf_c1_rf_chdad_reg[10]/NET0131 , \ctl_rf_c1_rf_chdad_reg[11]/P0002 , \ctl_rf_c1_rf_chdad_reg[12]/NET0131 , \ctl_rf_c1_rf_chdad_reg[13]/NET0131 , \ctl_rf_c1_rf_chdad_reg[14]/NET0131 , \ctl_rf_c1_rf_chdad_reg[15]/NET0131 , \ctl_rf_c1_rf_chdad_reg[16]/NET0131 , \ctl_rf_c1_rf_chdad_reg[17]/NET0131 , \ctl_rf_c1_rf_chdad_reg[18]/NET0131 , \ctl_rf_c1_rf_chdad_reg[19]/NET0131 , \ctl_rf_c1_rf_chdad_reg[1]/NET0131 , \ctl_rf_c1_rf_chdad_reg[20]/P0002 , \ctl_rf_c1_rf_chdad_reg[21]/P0002 , \ctl_rf_c1_rf_chdad_reg[22]/P0002 , \ctl_rf_c1_rf_chdad_reg[23]/P0002 , \ctl_rf_c1_rf_chdad_reg[24]/P0002 , \ctl_rf_c1_rf_chdad_reg[25]/P0002 , \ctl_rf_c1_rf_chdad_reg[26]/P0002 , \ctl_rf_c1_rf_chdad_reg[27]/P0002 , \ctl_rf_c1_rf_chdad_reg[28]/P0002 , \ctl_rf_c1_rf_chdad_reg[29]/P0002 , \ctl_rf_c1_rf_chdad_reg[2]/NET0131 , \ctl_rf_c1_rf_chdad_reg[30]/P0002 , \ctl_rf_c1_rf_chdad_reg[31]/P0002 , \ctl_rf_c1_rf_chdad_reg[3]/P0002 , \ctl_rf_c1_rf_chdad_reg[4]/P0002 , \ctl_rf_c1_rf_chdad_reg[5]/P0002 , \ctl_rf_c1_rf_chdad_reg[6]/P0002 , \ctl_rf_c1_rf_chdad_reg[7]/P0002 , \ctl_rf_c1_rf_chdad_reg[8]/NET0131 , \ctl_rf_c1_rf_chdad_reg[9]/P0002 , \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c1_rf_chllp_on_reg/NET0131 , \ctl_rf_c1_rf_chllp_reg[0]/P0002 , \ctl_rf_c1_rf_chllp_reg[10]/NET0131 , \ctl_rf_c1_rf_chllp_reg[11]/NET0131 , \ctl_rf_c1_rf_chllp_reg[12]/NET0131 , \ctl_rf_c1_rf_chllp_reg[13]/NET0131 , \ctl_rf_c1_rf_chllp_reg[14]/NET0131 , \ctl_rf_c1_rf_chllp_reg[15]/NET0131 , \ctl_rf_c1_rf_chllp_reg[16]/NET0131 , \ctl_rf_c1_rf_chllp_reg[17]/NET0131 , \ctl_rf_c1_rf_chllp_reg[18]/NET0131 , \ctl_rf_c1_rf_chllp_reg[19]/NET0131 , \ctl_rf_c1_rf_chllp_reg[1]/P0002 , \ctl_rf_c1_rf_chllp_reg[20]/NET0131 , \ctl_rf_c1_rf_chllp_reg[21]/NET0131 , \ctl_rf_c1_rf_chllp_reg[22]/NET0131 , \ctl_rf_c1_rf_chllp_reg[23]/NET0131 , \ctl_rf_c1_rf_chllp_reg[24]/NET0131 , \ctl_rf_c1_rf_chllp_reg[25]/NET0131 , \ctl_rf_c1_rf_chllp_reg[26]/NET0131 , \ctl_rf_c1_rf_chllp_reg[27]/NET0131 , \ctl_rf_c1_rf_chllp_reg[28]/NET0131 , \ctl_rf_c1_rf_chllp_reg[29]/NET0131 , \ctl_rf_c1_rf_chllp_reg[2]/NET0131 , \ctl_rf_c1_rf_chllp_reg[30]/NET0131 , \ctl_rf_c1_rf_chllp_reg[31]/NET0131 , \ctl_rf_c1_rf_chllp_reg[3]/NET0131 , \ctl_rf_c1_rf_chllp_reg[4]/NET0131 , \ctl_rf_c1_rf_chllp_reg[5]/NET0131 , \ctl_rf_c1_rf_chllp_reg[6]/NET0131 , \ctl_rf_c1_rf_chllp_reg[7]/NET0131 , \ctl_rf_c1_rf_chllp_reg[8]/NET0131 , \ctl_rf_c1_rf_chllp_reg[9]/NET0131 , \ctl_rf_c1_rf_chllpen_reg/NET0131 , \ctl_rf_c1_rf_chpri_reg[0]/NET0131 , \ctl_rf_c1_rf_chpri_reg[1]/NET0131 , \ctl_rf_c1_rf_chsad_reg[0]/NET0131 , \ctl_rf_c1_rf_chsad_reg[10]/P0002 , \ctl_rf_c1_rf_chsad_reg[11]/NET0131 , \ctl_rf_c1_rf_chsad_reg[12]/P0002 , \ctl_rf_c1_rf_chsad_reg[13]/P0002 , \ctl_rf_c1_rf_chsad_reg[14]/P0002 , \ctl_rf_c1_rf_chsad_reg[15]/P0002 , \ctl_rf_c1_rf_chsad_reg[16]/NET0131 , \ctl_rf_c1_rf_chsad_reg[17]/NET0131 , \ctl_rf_c1_rf_chsad_reg[18]/NET0131 , \ctl_rf_c1_rf_chsad_reg[19]/NET0131 , \ctl_rf_c1_rf_chsad_reg[1]/NET0131 , \ctl_rf_c1_rf_chsad_reg[20]/NET0131 , \ctl_rf_c1_rf_chsad_reg[21]/NET0131 , \ctl_rf_c1_rf_chsad_reg[22]/NET0131 , \ctl_rf_c1_rf_chsad_reg[23]/NET0131 , \ctl_rf_c1_rf_chsad_reg[24]/NET0131 , \ctl_rf_c1_rf_chsad_reg[25]/P0002 , \ctl_rf_c1_rf_chsad_reg[26]/P0002 , \ctl_rf_c1_rf_chsad_reg[27]/P0002 , \ctl_rf_c1_rf_chsad_reg[28]/P0002 , \ctl_rf_c1_rf_chsad_reg[29]/P0002 , \ctl_rf_c1_rf_chsad_reg[2]/NET0131 , \ctl_rf_c1_rf_chsad_reg[30]/P0002 , \ctl_rf_c1_rf_chsad_reg[31]/NET0131 , \ctl_rf_c1_rf_chsad_reg[3]/NET0131 , \ctl_rf_c1_rf_chsad_reg[4]/NET0131 , \ctl_rf_c1_rf_chsad_reg[5]/NET0131 , \ctl_rf_c1_rf_chsad_reg[6]/NET0131 , \ctl_rf_c1_rf_chsad_reg[7]/NET0131 , \ctl_rf_c1_rf_chsad_reg[8]/P0002 , \ctl_rf_c1_rf_chsad_reg[9]/NET0131 , \ctl_rf_c1_rf_chtsz_reg[0]/P0002 , \ctl_rf_c1_rf_chtsz_reg[10]/P0002 , \ctl_rf_c1_rf_chtsz_reg[11]/P0002 , \ctl_rf_c1_rf_chtsz_reg[1]/P0002 , \ctl_rf_c1_rf_chtsz_reg[2]/P0002 , \ctl_rf_c1_rf_chtsz_reg[3]/P0002 , \ctl_rf_c1_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c1_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c1_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c1_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c1_rf_chtsz_reg[8]/P0002 , \ctl_rf_c1_rf_chtsz_reg[9]/P0002 , \ctl_rf_c1_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c1_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c1_rf_dreqmode_reg/NET0131 , \ctl_rf_c1_rf_dst_sel_reg/NET0131 , \ctl_rf_c1_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c1_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c1_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c1_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c1_rf_int_err_msk_reg/NET0131 , \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c1_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c1_rf_mode_reg/NET0131 , \ctl_rf_c1_rf_prot1_reg/NET0131 , \ctl_rf_c1_rf_prot2_reg/NET0131 , \ctl_rf_c1_rf_prot3_reg/NET0131 , \ctl_rf_c1_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c1_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c1_rf_src_sel_reg/NET0131 , \ctl_rf_c1_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c1_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c1_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c1_rf_swidth_reg[0]/NET0131 , \ctl_rf_c1_rf_swidth_reg[1]/NET0131 , \ctl_rf_c1_rf_swidth_reg[2]/NET0131 , \ctl_rf_c1brbs_reg[16]/NET0131 , \ctl_rf_c1brbs_reg[17]/NET0131 , \ctl_rf_c1brbs_reg[18]/NET0131 , \ctl_rf_c1brbs_reg[19]/NET0131 , \ctl_rf_c1brbs_reg[20]/NET0131 , \ctl_rf_c1brbs_reg[21]/NET0131 , \ctl_rf_c1brbs_reg[22]/NET0131 , \ctl_rf_c1brbs_reg[23]/NET0131 , \ctl_rf_c1brbs_reg[24]/NET0131 , \ctl_rf_c1brbs_reg[25]/NET0131 , \ctl_rf_c1brbs_reg[26]/NET0131 , \ctl_rf_c1brbs_reg[27]/NET0131 , \ctl_rf_c1brbs_reg[28]/NET0131 , \ctl_rf_c1brbs_reg[29]/NET0131 , \ctl_rf_c1brbs_reg[30]/NET0131 , \ctl_rf_c1brbs_reg[31]/NET0131 , \ctl_rf_c1dmabs_reg[16]/NET0131 , \ctl_rf_c1dmabs_reg[17]/NET0131 , \ctl_rf_c1dmabs_reg[18]/NET0131 , \ctl_rf_c1dmabs_reg[19]/NET0131 , \ctl_rf_c1dmabs_reg[20]/NET0131 , \ctl_rf_c1dmabs_reg[21]/NET0131 , \ctl_rf_c1dmabs_reg[22]/NET0131 , \ctl_rf_c1dmabs_reg[23]/NET0131 , \ctl_rf_c1dmabs_reg[24]/NET0131 , \ctl_rf_c1dmabs_reg[25]/NET0131 , \ctl_rf_c1dmabs_reg[26]/NET0131 , \ctl_rf_c1dmabs_reg[27]/NET0131 , \ctl_rf_c1dmabs_reg[28]/NET0131 , \ctl_rf_c1dmabs_reg[29]/NET0131 , \ctl_rf_c1dmabs_reg[30]/NET0131 , \ctl_rf_c1dmabs_reg[31]/NET0131 , \ctl_rf_c2_rf_autold_reg/NET0131 , \ctl_rf_c2_rf_ch_en_reg/NET0131 , \ctl_rf_c2_rf_chabt_reg/NET0131 , \ctl_rf_c2_rf_chdad_reg[0]/NET0131 , \ctl_rf_c2_rf_chdad_reg[10]/P0002 , \ctl_rf_c2_rf_chdad_reg[11]/P0002 , \ctl_rf_c2_rf_chdad_reg[12]/P0002 , \ctl_rf_c2_rf_chdad_reg[13]/P0002 , \ctl_rf_c2_rf_chdad_reg[14]/P0002 , \ctl_rf_c2_rf_chdad_reg[15]/P0002 , \ctl_rf_c2_rf_chdad_reg[16]/NET0131 , \ctl_rf_c2_rf_chdad_reg[17]/NET0131 , \ctl_rf_c2_rf_chdad_reg[18]/NET0131 , \ctl_rf_c2_rf_chdad_reg[19]/NET0131 , \ctl_rf_c2_rf_chdad_reg[1]/NET0131 , \ctl_rf_c2_rf_chdad_reg[20]/P0002 , \ctl_rf_c2_rf_chdad_reg[21]/P0002 , \ctl_rf_c2_rf_chdad_reg[22]/P0002 , \ctl_rf_c2_rf_chdad_reg[23]/P0002 , \ctl_rf_c2_rf_chdad_reg[24]/P0002 , \ctl_rf_c2_rf_chdad_reg[25]/P0002 , \ctl_rf_c2_rf_chdad_reg[26]/P0002 , \ctl_rf_c2_rf_chdad_reg[27]/P0002 , \ctl_rf_c2_rf_chdad_reg[28]/P0002 , \ctl_rf_c2_rf_chdad_reg[29]/P0002 , \ctl_rf_c2_rf_chdad_reg[2]/NET0131 , \ctl_rf_c2_rf_chdad_reg[30]/P0002 , \ctl_rf_c2_rf_chdad_reg[31]/P0002 , \ctl_rf_c2_rf_chdad_reg[3]/P0002 , \ctl_rf_c2_rf_chdad_reg[4]/P0002 , \ctl_rf_c2_rf_chdad_reg[5]/P0002 , \ctl_rf_c2_rf_chdad_reg[6]/P0002 , \ctl_rf_c2_rf_chdad_reg[7]/P0002 , \ctl_rf_c2_rf_chdad_reg[8]/NET0131 , \ctl_rf_c2_rf_chdad_reg[9]/P0002 , \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c2_rf_chllp_on_reg/NET0131 , \ctl_rf_c2_rf_chllp_reg[0]/P0002 , \ctl_rf_c2_rf_chllp_reg[10]/NET0131 , \ctl_rf_c2_rf_chllp_reg[11]/NET0131 , \ctl_rf_c2_rf_chllp_reg[12]/NET0131 , \ctl_rf_c2_rf_chllp_reg[13]/NET0131 , \ctl_rf_c2_rf_chllp_reg[14]/NET0131 , \ctl_rf_c2_rf_chllp_reg[15]/NET0131 , \ctl_rf_c2_rf_chllp_reg[16]/NET0131 , \ctl_rf_c2_rf_chllp_reg[17]/NET0131 , \ctl_rf_c2_rf_chllp_reg[18]/NET0131 , \ctl_rf_c2_rf_chllp_reg[19]/NET0131 , \ctl_rf_c2_rf_chllp_reg[1]/P0002 , \ctl_rf_c2_rf_chllp_reg[20]/NET0131 , \ctl_rf_c2_rf_chllp_reg[21]/NET0131 , \ctl_rf_c2_rf_chllp_reg[22]/NET0131 , \ctl_rf_c2_rf_chllp_reg[23]/NET0131 , \ctl_rf_c2_rf_chllp_reg[24]/NET0131 , \ctl_rf_c2_rf_chllp_reg[25]/NET0131 , \ctl_rf_c2_rf_chllp_reg[26]/NET0131 , \ctl_rf_c2_rf_chllp_reg[27]/NET0131 , \ctl_rf_c2_rf_chllp_reg[28]/NET0131 , \ctl_rf_c2_rf_chllp_reg[29]/NET0131 , \ctl_rf_c2_rf_chllp_reg[2]/NET0131 , \ctl_rf_c2_rf_chllp_reg[30]/NET0131 , \ctl_rf_c2_rf_chllp_reg[31]/NET0131 , \ctl_rf_c2_rf_chllp_reg[3]/NET0131 , \ctl_rf_c2_rf_chllp_reg[4]/NET0131 , \ctl_rf_c2_rf_chllp_reg[5]/NET0131 , \ctl_rf_c2_rf_chllp_reg[6]/NET0131 , \ctl_rf_c2_rf_chllp_reg[7]/NET0131 , \ctl_rf_c2_rf_chllp_reg[8]/NET0131 , \ctl_rf_c2_rf_chllp_reg[9]/NET0131 , \ctl_rf_c2_rf_chllpen_reg/NET0131 , \ctl_rf_c2_rf_chpri_reg[0]/NET0131 , \ctl_rf_c2_rf_chpri_reg[1]/NET0131 , \ctl_rf_c2_rf_chsad_reg[0]/NET0131 , \ctl_rf_c2_rf_chsad_reg[10]/NET0131 , \ctl_rf_c2_rf_chsad_reg[11]/NET0131 , \ctl_rf_c2_rf_chsad_reg[12]/NET0131 , \ctl_rf_c2_rf_chsad_reg[13]/NET0131 , \ctl_rf_c2_rf_chsad_reg[14]/NET0131 , \ctl_rf_c2_rf_chsad_reg[15]/NET0131 , \ctl_rf_c2_rf_chsad_reg[16]/NET0131 , \ctl_rf_c2_rf_chsad_reg[17]/NET0131 , \ctl_rf_c2_rf_chsad_reg[18]/NET0131 , \ctl_rf_c2_rf_chsad_reg[19]/NET0131 , \ctl_rf_c2_rf_chsad_reg[1]/NET0131 , \ctl_rf_c2_rf_chsad_reg[20]/NET0131 , \ctl_rf_c2_rf_chsad_reg[21]/NET0131 , \ctl_rf_c2_rf_chsad_reg[22]/NET0131 , \ctl_rf_c2_rf_chsad_reg[23]/NET0131 , \ctl_rf_c2_rf_chsad_reg[24]/NET0131 , \ctl_rf_c2_rf_chsad_reg[25]/P0002 , \ctl_rf_c2_rf_chsad_reg[26]/P0002 , \ctl_rf_c2_rf_chsad_reg[27]/P0002 , \ctl_rf_c2_rf_chsad_reg[28]/P0002 , \ctl_rf_c2_rf_chsad_reg[29]/P0002 , \ctl_rf_c2_rf_chsad_reg[2]/NET0131 , \ctl_rf_c2_rf_chsad_reg[30]/P0002 , \ctl_rf_c2_rf_chsad_reg[31]/NET0131 , \ctl_rf_c2_rf_chsad_reg[3]/NET0131 , \ctl_rf_c2_rf_chsad_reg[4]/NET0131 , \ctl_rf_c2_rf_chsad_reg[5]/NET0131 , \ctl_rf_c2_rf_chsad_reg[6]/NET0131 , \ctl_rf_c2_rf_chsad_reg[7]/NET0131 , \ctl_rf_c2_rf_chsad_reg[8]/P0002 , \ctl_rf_c2_rf_chsad_reg[9]/NET0131 , \ctl_rf_c2_rf_chtsz_reg[0]/P0002 , \ctl_rf_c2_rf_chtsz_reg[10]/P0002 , \ctl_rf_c2_rf_chtsz_reg[11]/P0002 , \ctl_rf_c2_rf_chtsz_reg[1]/P0002 , \ctl_rf_c2_rf_chtsz_reg[2]/P0002 , \ctl_rf_c2_rf_chtsz_reg[3]/P0002 , \ctl_rf_c2_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c2_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c2_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c2_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c2_rf_chtsz_reg[8]/P0002 , \ctl_rf_c2_rf_chtsz_reg[9]/P0002 , \ctl_rf_c2_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c2_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c2_rf_dreqmode_reg/NET0131 , \ctl_rf_c2_rf_dst_sel_reg/NET0131 , \ctl_rf_c2_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c2_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c2_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c2_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c2_rf_int_err_msk_reg/NET0131 , \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c2_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c2_rf_mode_reg/NET0131 , \ctl_rf_c2_rf_prot1_reg/NET0131 , \ctl_rf_c2_rf_prot2_reg/NET0131 , \ctl_rf_c2_rf_prot3_reg/NET0131 , \ctl_rf_c2_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c2_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c2_rf_src_sel_reg/NET0131 , \ctl_rf_c2_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c2_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c2_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c2_rf_swidth_reg[0]/NET0131 , \ctl_rf_c2_rf_swidth_reg[1]/NET0131 , \ctl_rf_c2_rf_swidth_reg[2]/NET0131 , \ctl_rf_c2brbs_reg[16]/NET0131 , \ctl_rf_c2brbs_reg[17]/NET0131 , \ctl_rf_c2brbs_reg[18]/NET0131 , \ctl_rf_c2brbs_reg[19]/NET0131 , \ctl_rf_c2brbs_reg[20]/NET0131 , \ctl_rf_c2brbs_reg[21]/NET0131 , \ctl_rf_c2brbs_reg[22]/NET0131 , \ctl_rf_c2brbs_reg[23]/NET0131 , \ctl_rf_c2brbs_reg[24]/NET0131 , \ctl_rf_c2brbs_reg[25]/NET0131 , \ctl_rf_c2brbs_reg[26]/NET0131 , \ctl_rf_c2brbs_reg[27]/NET0131 , \ctl_rf_c2brbs_reg[28]/NET0131 , \ctl_rf_c2brbs_reg[29]/NET0131 , \ctl_rf_c2brbs_reg[30]/NET0131 , \ctl_rf_c2brbs_reg[31]/NET0131 , \ctl_rf_c2dmabs_reg[16]/NET0131 , \ctl_rf_c2dmabs_reg[17]/NET0131 , \ctl_rf_c2dmabs_reg[18]/NET0131 , \ctl_rf_c2dmabs_reg[19]/NET0131 , \ctl_rf_c2dmabs_reg[20]/NET0131 , \ctl_rf_c2dmabs_reg[21]/NET0131 , \ctl_rf_c2dmabs_reg[22]/NET0131 , \ctl_rf_c2dmabs_reg[23]/NET0131 , \ctl_rf_c2dmabs_reg[24]/NET0131 , \ctl_rf_c2dmabs_reg[25]/NET0131 , \ctl_rf_c2dmabs_reg[26]/NET0131 , \ctl_rf_c2dmabs_reg[27]/NET0131 , \ctl_rf_c2dmabs_reg[28]/NET0131 , \ctl_rf_c2dmabs_reg[29]/NET0131 , \ctl_rf_c2dmabs_reg[30]/NET0131 , \ctl_rf_c2dmabs_reg[31]/NET0131 , \ctl_rf_c3_rf_autold_reg/NET0131 , \ctl_rf_c3_rf_ch_en_reg/NET0131 , \ctl_rf_c3_rf_chabt_reg/NET0131 , \ctl_rf_c3_rf_chdad_reg[0]/NET0131 , \ctl_rf_c3_rf_chdad_reg[10]/NET0131 , \ctl_rf_c3_rf_chdad_reg[11]/NET0131 , \ctl_rf_c3_rf_chdad_reg[12]/NET0131 , \ctl_rf_c3_rf_chdad_reg[13]/P0002 , \ctl_rf_c3_rf_chdad_reg[14]/P0002 , \ctl_rf_c3_rf_chdad_reg[15]/NET0131 , \ctl_rf_c3_rf_chdad_reg[16]/NET0131 , \ctl_rf_c3_rf_chdad_reg[17]/NET0131 , \ctl_rf_c3_rf_chdad_reg[18]/NET0131 , \ctl_rf_c3_rf_chdad_reg[19]/NET0131 , \ctl_rf_c3_rf_chdad_reg[1]/NET0131 , \ctl_rf_c3_rf_chdad_reg[20]/P0002 , \ctl_rf_c3_rf_chdad_reg[21]/P0002 , \ctl_rf_c3_rf_chdad_reg[22]/P0002 , \ctl_rf_c3_rf_chdad_reg[23]/P0002 , \ctl_rf_c3_rf_chdad_reg[24]/P0002 , \ctl_rf_c3_rf_chdad_reg[25]/P0002 , \ctl_rf_c3_rf_chdad_reg[26]/P0002 , \ctl_rf_c3_rf_chdad_reg[27]/P0002 , \ctl_rf_c3_rf_chdad_reg[28]/P0002 , \ctl_rf_c3_rf_chdad_reg[29]/P0002 , \ctl_rf_c3_rf_chdad_reg[2]/NET0131 , \ctl_rf_c3_rf_chdad_reg[30]/P0002 , \ctl_rf_c3_rf_chdad_reg[31]/P0002 , \ctl_rf_c3_rf_chdad_reg[3]/P0002 , \ctl_rf_c3_rf_chdad_reg[4]/P0002 , \ctl_rf_c3_rf_chdad_reg[5]/P0002 , \ctl_rf_c3_rf_chdad_reg[6]/P0002 , \ctl_rf_c3_rf_chdad_reg[7]/P0002 , \ctl_rf_c3_rf_chdad_reg[8]/NET0131 , \ctl_rf_c3_rf_chdad_reg[9]/P0002 , \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c3_rf_chllp_on_reg/NET0131 , \ctl_rf_c3_rf_chllp_reg[0]/P0002 , \ctl_rf_c3_rf_chllp_reg[10]/NET0131 , \ctl_rf_c3_rf_chllp_reg[11]/NET0131 , \ctl_rf_c3_rf_chllp_reg[12]/NET0131 , \ctl_rf_c3_rf_chllp_reg[13]/NET0131 , \ctl_rf_c3_rf_chllp_reg[14]/NET0131 , \ctl_rf_c3_rf_chllp_reg[15]/NET0131 , \ctl_rf_c3_rf_chllp_reg[16]/NET0131 , \ctl_rf_c3_rf_chllp_reg[17]/NET0131 , \ctl_rf_c3_rf_chllp_reg[18]/NET0131 , \ctl_rf_c3_rf_chllp_reg[19]/NET0131 , \ctl_rf_c3_rf_chllp_reg[1]/P0002 , \ctl_rf_c3_rf_chllp_reg[20]/NET0131 , \ctl_rf_c3_rf_chllp_reg[21]/NET0131 , \ctl_rf_c3_rf_chllp_reg[22]/NET0131 , \ctl_rf_c3_rf_chllp_reg[23]/NET0131 , \ctl_rf_c3_rf_chllp_reg[24]/NET0131 , \ctl_rf_c3_rf_chllp_reg[25]/NET0131 , \ctl_rf_c3_rf_chllp_reg[26]/NET0131 , \ctl_rf_c3_rf_chllp_reg[27]/NET0131 , \ctl_rf_c3_rf_chllp_reg[28]/NET0131 , \ctl_rf_c3_rf_chllp_reg[29]/NET0131 , \ctl_rf_c3_rf_chllp_reg[2]/NET0131 , \ctl_rf_c3_rf_chllp_reg[30]/NET0131 , \ctl_rf_c3_rf_chllp_reg[31]/NET0131 , \ctl_rf_c3_rf_chllp_reg[3]/NET0131 , \ctl_rf_c3_rf_chllp_reg[4]/NET0131 , \ctl_rf_c3_rf_chllp_reg[5]/NET0131 , \ctl_rf_c3_rf_chllp_reg[6]/NET0131 , \ctl_rf_c3_rf_chllp_reg[7]/NET0131 , \ctl_rf_c3_rf_chllp_reg[8]/NET0131 , \ctl_rf_c3_rf_chllp_reg[9]/NET0131 , \ctl_rf_c3_rf_chllpen_reg/NET0131 , \ctl_rf_c3_rf_chpri_reg[0]/NET0131 , \ctl_rf_c3_rf_chpri_reg[1]/NET0131 , \ctl_rf_c3_rf_chsad_reg[0]/NET0131 , \ctl_rf_c3_rf_chsad_reg[10]/P0002 , \ctl_rf_c3_rf_chsad_reg[11]/P0002 , \ctl_rf_c3_rf_chsad_reg[12]/P0002 , \ctl_rf_c3_rf_chsad_reg[13]/NET0131 , \ctl_rf_c3_rf_chsad_reg[14]/NET0131 , \ctl_rf_c3_rf_chsad_reg[15]/P0002 , \ctl_rf_c3_rf_chsad_reg[16]/NET0131 , \ctl_rf_c3_rf_chsad_reg[17]/NET0131 , \ctl_rf_c3_rf_chsad_reg[18]/NET0131 , \ctl_rf_c3_rf_chsad_reg[19]/NET0131 , \ctl_rf_c3_rf_chsad_reg[1]/NET0131 , \ctl_rf_c3_rf_chsad_reg[20]/NET0131 , \ctl_rf_c3_rf_chsad_reg[21]/NET0131 , \ctl_rf_c3_rf_chsad_reg[22]/NET0131 , \ctl_rf_c3_rf_chsad_reg[23]/NET0131 , \ctl_rf_c3_rf_chsad_reg[24]/NET0131 , \ctl_rf_c3_rf_chsad_reg[25]/P0002 , \ctl_rf_c3_rf_chsad_reg[26]/P0002 , \ctl_rf_c3_rf_chsad_reg[27]/P0002 , \ctl_rf_c3_rf_chsad_reg[28]/P0002 , \ctl_rf_c3_rf_chsad_reg[29]/P0002 , \ctl_rf_c3_rf_chsad_reg[2]/NET0131 , \ctl_rf_c3_rf_chsad_reg[30]/P0002 , \ctl_rf_c3_rf_chsad_reg[31]/NET0131 , \ctl_rf_c3_rf_chsad_reg[3]/NET0131 , \ctl_rf_c3_rf_chsad_reg[4]/NET0131 , \ctl_rf_c3_rf_chsad_reg[5]/NET0131 , \ctl_rf_c3_rf_chsad_reg[6]/NET0131 , \ctl_rf_c3_rf_chsad_reg[7]/NET0131 , \ctl_rf_c3_rf_chsad_reg[8]/P0002 , \ctl_rf_c3_rf_chsad_reg[9]/NET0131 , \ctl_rf_c3_rf_chtsz_reg[0]/P0002 , \ctl_rf_c3_rf_chtsz_reg[10]/P0002 , \ctl_rf_c3_rf_chtsz_reg[11]/P0002 , \ctl_rf_c3_rf_chtsz_reg[1]/P0002 , \ctl_rf_c3_rf_chtsz_reg[2]/P0002 , \ctl_rf_c3_rf_chtsz_reg[3]/P0002 , \ctl_rf_c3_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c3_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c3_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c3_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c3_rf_chtsz_reg[8]/P0002 , \ctl_rf_c3_rf_chtsz_reg[9]/P0002 , \ctl_rf_c3_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c3_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c3_rf_dreqmode_reg/NET0131 , \ctl_rf_c3_rf_dst_sel_reg/NET0131 , \ctl_rf_c3_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c3_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c3_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c3_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c3_rf_int_err_msk_reg/NET0131 , \ctl_rf_c3_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c3_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c3_rf_mode_reg/NET0131 , \ctl_rf_c3_rf_prot1_reg/NET0131 , \ctl_rf_c3_rf_prot2_reg/NET0131 , \ctl_rf_c3_rf_prot3_reg/NET0131 , \ctl_rf_c3_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c3_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c3_rf_src_sel_reg/NET0131 , \ctl_rf_c3_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c3_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c3_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c3_rf_swidth_reg[0]/NET0131 , \ctl_rf_c3_rf_swidth_reg[1]/NET0131 , \ctl_rf_c3_rf_swidth_reg[2]/NET0131 , \ctl_rf_c3brbs_reg[16]/NET0131 , \ctl_rf_c3brbs_reg[17]/NET0131 , \ctl_rf_c3brbs_reg[18]/NET0131 , \ctl_rf_c3brbs_reg[19]/NET0131 , \ctl_rf_c3brbs_reg[20]/NET0131 , \ctl_rf_c3brbs_reg[21]/NET0131 , \ctl_rf_c3brbs_reg[22]/NET0131 , \ctl_rf_c3brbs_reg[23]/NET0131 , \ctl_rf_c3brbs_reg[24]/NET0131 , \ctl_rf_c3brbs_reg[25]/NET0131 , \ctl_rf_c3brbs_reg[26]/NET0131 , \ctl_rf_c3brbs_reg[27]/NET0131 , \ctl_rf_c3brbs_reg[28]/NET0131 , \ctl_rf_c3brbs_reg[29]/NET0131 , \ctl_rf_c3brbs_reg[30]/NET0131 , \ctl_rf_c3brbs_reg[31]/NET0131 , \ctl_rf_c3dmabs_reg[16]/NET0131 , \ctl_rf_c3dmabs_reg[17]/NET0131 , \ctl_rf_c3dmabs_reg[18]/NET0131 , \ctl_rf_c3dmabs_reg[19]/NET0131 , \ctl_rf_c3dmabs_reg[20]/NET0131 , \ctl_rf_c3dmabs_reg[21]/NET0131 , \ctl_rf_c3dmabs_reg[22]/NET0131 , \ctl_rf_c3dmabs_reg[23]/NET0131 , \ctl_rf_c3dmabs_reg[24]/NET0131 , \ctl_rf_c3dmabs_reg[25]/NET0131 , \ctl_rf_c3dmabs_reg[26]/NET0131 , \ctl_rf_c3dmabs_reg[27]/NET0131 , \ctl_rf_c3dmabs_reg[28]/NET0131 , \ctl_rf_c3dmabs_reg[29]/NET0131 , \ctl_rf_c3dmabs_reg[30]/NET0131 , \ctl_rf_c3dmabs_reg[31]/NET0131 , \ctl_rf_c4_rf_autold_reg/NET0131 , \ctl_rf_c4_rf_ch_en_reg/NET0131 , \ctl_rf_c4_rf_chabt_reg/NET0131 , \ctl_rf_c4_rf_chdad_reg[0]/NET0131 , \ctl_rf_c4_rf_chdad_reg[10]/P0002 , \ctl_rf_c4_rf_chdad_reg[11]/P0002 , \ctl_rf_c4_rf_chdad_reg[12]/P0002 , \ctl_rf_c4_rf_chdad_reg[13]/P0002 , \ctl_rf_c4_rf_chdad_reg[14]/P0002 , \ctl_rf_c4_rf_chdad_reg[15]/P0002 , \ctl_rf_c4_rf_chdad_reg[16]/NET0131 , \ctl_rf_c4_rf_chdad_reg[17]/NET0131 , \ctl_rf_c4_rf_chdad_reg[18]/NET0131 , \ctl_rf_c4_rf_chdad_reg[19]/NET0131 , \ctl_rf_c4_rf_chdad_reg[1]/NET0131 , \ctl_rf_c4_rf_chdad_reg[20]/P0002 , \ctl_rf_c4_rf_chdad_reg[21]/P0002 , \ctl_rf_c4_rf_chdad_reg[22]/P0002 , \ctl_rf_c4_rf_chdad_reg[23]/P0002 , \ctl_rf_c4_rf_chdad_reg[24]/P0002 , \ctl_rf_c4_rf_chdad_reg[25]/P0002 , \ctl_rf_c4_rf_chdad_reg[26]/P0002 , \ctl_rf_c4_rf_chdad_reg[27]/P0002 , \ctl_rf_c4_rf_chdad_reg[28]/P0002 , \ctl_rf_c4_rf_chdad_reg[29]/P0002 , \ctl_rf_c4_rf_chdad_reg[2]/NET0131 , \ctl_rf_c4_rf_chdad_reg[30]/P0002 , \ctl_rf_c4_rf_chdad_reg[31]/P0002 , \ctl_rf_c4_rf_chdad_reg[3]/P0002 , \ctl_rf_c4_rf_chdad_reg[4]/P0002 , \ctl_rf_c4_rf_chdad_reg[5]/P0002 , \ctl_rf_c4_rf_chdad_reg[6]/P0002 , \ctl_rf_c4_rf_chdad_reg[7]/P0002 , \ctl_rf_c4_rf_chdad_reg[8]/NET0131 , \ctl_rf_c4_rf_chdad_reg[9]/P0002 , \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c4_rf_chllp_on_reg/NET0131 , \ctl_rf_c4_rf_chllp_reg[0]/P0002 , \ctl_rf_c4_rf_chllp_reg[10]/NET0131 , \ctl_rf_c4_rf_chllp_reg[11]/NET0131 , \ctl_rf_c4_rf_chllp_reg[12]/NET0131 , \ctl_rf_c4_rf_chllp_reg[13]/NET0131 , \ctl_rf_c4_rf_chllp_reg[14]/NET0131 , \ctl_rf_c4_rf_chllp_reg[15]/NET0131 , \ctl_rf_c4_rf_chllp_reg[16]/NET0131 , \ctl_rf_c4_rf_chllp_reg[17]/NET0131 , \ctl_rf_c4_rf_chllp_reg[18]/NET0131 , \ctl_rf_c4_rf_chllp_reg[19]/NET0131 , \ctl_rf_c4_rf_chllp_reg[1]/P0002 , \ctl_rf_c4_rf_chllp_reg[20]/NET0131 , \ctl_rf_c4_rf_chllp_reg[21]/NET0131 , \ctl_rf_c4_rf_chllp_reg[22]/NET0131 , \ctl_rf_c4_rf_chllp_reg[23]/NET0131 , \ctl_rf_c4_rf_chllp_reg[24]/NET0131 , \ctl_rf_c4_rf_chllp_reg[25]/NET0131 , \ctl_rf_c4_rf_chllp_reg[26]/NET0131 , \ctl_rf_c4_rf_chllp_reg[27]/NET0131 , \ctl_rf_c4_rf_chllp_reg[28]/NET0131 , \ctl_rf_c4_rf_chllp_reg[29]/NET0131 , \ctl_rf_c4_rf_chllp_reg[2]/NET0131 , \ctl_rf_c4_rf_chllp_reg[30]/NET0131 , \ctl_rf_c4_rf_chllp_reg[31]/NET0131 , \ctl_rf_c4_rf_chllp_reg[3]/NET0131 , \ctl_rf_c4_rf_chllp_reg[4]/NET0131 , \ctl_rf_c4_rf_chllp_reg[5]/NET0131 , \ctl_rf_c4_rf_chllp_reg[6]/NET0131 , \ctl_rf_c4_rf_chllp_reg[7]/NET0131 , \ctl_rf_c4_rf_chllp_reg[8]/NET0131 , \ctl_rf_c4_rf_chllp_reg[9]/NET0131 , \ctl_rf_c4_rf_chllpen_reg/NET0131 , \ctl_rf_c4_rf_chpri_reg[0]/NET0131 , \ctl_rf_c4_rf_chpri_reg[1]/NET0131 , \ctl_rf_c4_rf_chsad_reg[0]/NET0131 , \ctl_rf_c4_rf_chsad_reg[10]/NET0131 , \ctl_rf_c4_rf_chsad_reg[11]/NET0131 , \ctl_rf_c4_rf_chsad_reg[12]/NET0131 , \ctl_rf_c4_rf_chsad_reg[13]/NET0131 , \ctl_rf_c4_rf_chsad_reg[14]/NET0131 , \ctl_rf_c4_rf_chsad_reg[15]/NET0131 , \ctl_rf_c4_rf_chsad_reg[16]/NET0131 , \ctl_rf_c4_rf_chsad_reg[17]/NET0131 , \ctl_rf_c4_rf_chsad_reg[18]/NET0131 , \ctl_rf_c4_rf_chsad_reg[19]/NET0131 , \ctl_rf_c4_rf_chsad_reg[1]/NET0131 , \ctl_rf_c4_rf_chsad_reg[20]/NET0131 , \ctl_rf_c4_rf_chsad_reg[21]/NET0131 , \ctl_rf_c4_rf_chsad_reg[22]/NET0131 , \ctl_rf_c4_rf_chsad_reg[23]/NET0131 , \ctl_rf_c4_rf_chsad_reg[24]/NET0131 , \ctl_rf_c4_rf_chsad_reg[25]/P0002 , \ctl_rf_c4_rf_chsad_reg[26]/P0002 , \ctl_rf_c4_rf_chsad_reg[27]/P0002 , \ctl_rf_c4_rf_chsad_reg[28]/P0002 , \ctl_rf_c4_rf_chsad_reg[29]/P0002 , \ctl_rf_c4_rf_chsad_reg[2]/NET0131 , \ctl_rf_c4_rf_chsad_reg[30]/P0002 , \ctl_rf_c4_rf_chsad_reg[31]/NET0131 , \ctl_rf_c4_rf_chsad_reg[3]/NET0131 , \ctl_rf_c4_rf_chsad_reg[4]/NET0131 , \ctl_rf_c4_rf_chsad_reg[5]/NET0131 , \ctl_rf_c4_rf_chsad_reg[6]/NET0131 , \ctl_rf_c4_rf_chsad_reg[7]/NET0131 , \ctl_rf_c4_rf_chsad_reg[8]/P0002 , \ctl_rf_c4_rf_chsad_reg[9]/NET0131 , \ctl_rf_c4_rf_chtsz_reg[0]/P0002 , \ctl_rf_c4_rf_chtsz_reg[10]/P0002 , \ctl_rf_c4_rf_chtsz_reg[11]/P0002 , \ctl_rf_c4_rf_chtsz_reg[1]/P0002 , \ctl_rf_c4_rf_chtsz_reg[2]/P0002 , \ctl_rf_c4_rf_chtsz_reg[3]/P0002 , \ctl_rf_c4_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c4_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c4_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c4_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c4_rf_chtsz_reg[8]/P0002 , \ctl_rf_c4_rf_chtsz_reg[9]/P0002 , \ctl_rf_c4_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c4_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c4_rf_dreqmode_reg/NET0131 , \ctl_rf_c4_rf_dst_sel_reg/NET0131 , \ctl_rf_c4_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c4_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c4_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c4_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c4_rf_int_err_msk_reg/NET0131 , \ctl_rf_c4_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c4_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c4_rf_mode_reg/NET0131 , \ctl_rf_c4_rf_prot1_reg/NET0131 , \ctl_rf_c4_rf_prot2_reg/NET0131 , \ctl_rf_c4_rf_prot3_reg/NET0131 , \ctl_rf_c4_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c4_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c4_rf_src_sel_reg/NET0131 , \ctl_rf_c4_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c4_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c4_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c4_rf_swidth_reg[0]/NET0131 , \ctl_rf_c4_rf_swidth_reg[1]/NET0131 , \ctl_rf_c4_rf_swidth_reg[2]/NET0131 , \ctl_rf_c4brbs_reg[16]/NET0131 , \ctl_rf_c4brbs_reg[17]/NET0131 , \ctl_rf_c4brbs_reg[18]/NET0131 , \ctl_rf_c4brbs_reg[19]/NET0131 , \ctl_rf_c4brbs_reg[20]/NET0131 , \ctl_rf_c4brbs_reg[21]/NET0131 , \ctl_rf_c4brbs_reg[22]/NET0131 , \ctl_rf_c4brbs_reg[23]/NET0131 , \ctl_rf_c4brbs_reg[24]/NET0131 , \ctl_rf_c4brbs_reg[25]/NET0131 , \ctl_rf_c4brbs_reg[26]/NET0131 , \ctl_rf_c4brbs_reg[27]/NET0131 , \ctl_rf_c4brbs_reg[28]/NET0131 , \ctl_rf_c4brbs_reg[29]/NET0131 , \ctl_rf_c4brbs_reg[30]/NET0131 , \ctl_rf_c4brbs_reg[31]/NET0131 , \ctl_rf_c4dmabs_reg[16]/NET0131 , \ctl_rf_c4dmabs_reg[17]/NET0131 , \ctl_rf_c4dmabs_reg[18]/NET0131 , \ctl_rf_c4dmabs_reg[19]/NET0131 , \ctl_rf_c4dmabs_reg[20]/NET0131 , \ctl_rf_c4dmabs_reg[21]/NET0131 , \ctl_rf_c4dmabs_reg[22]/NET0131 , \ctl_rf_c4dmabs_reg[23]/NET0131 , \ctl_rf_c4dmabs_reg[24]/NET0131 , \ctl_rf_c4dmabs_reg[25]/NET0131 , \ctl_rf_c4dmabs_reg[26]/NET0131 , \ctl_rf_c4dmabs_reg[27]/NET0131 , \ctl_rf_c4dmabs_reg[28]/NET0131 , \ctl_rf_c4dmabs_reg[29]/NET0131 , \ctl_rf_c4dmabs_reg[30]/NET0131 , \ctl_rf_c4dmabs_reg[31]/NET0131 , \ctl_rf_c5_rf_autold_reg/NET0131 , \ctl_rf_c5_rf_ch_en_reg/NET0131 , \ctl_rf_c5_rf_chabt_reg/NET0131 , \ctl_rf_c5_rf_chdad_reg[0]/NET0131 , \ctl_rf_c5_rf_chdad_reg[10]/P0002 , \ctl_rf_c5_rf_chdad_reg[11]/P0002 , \ctl_rf_c5_rf_chdad_reg[12]/P0002 , \ctl_rf_c5_rf_chdad_reg[13]/NET0131 , \ctl_rf_c5_rf_chdad_reg[14]/P0002 , \ctl_rf_c5_rf_chdad_reg[15]/P0002 , \ctl_rf_c5_rf_chdad_reg[16]/NET0131 , \ctl_rf_c5_rf_chdad_reg[17]/NET0131 , \ctl_rf_c5_rf_chdad_reg[18]/NET0131 , \ctl_rf_c5_rf_chdad_reg[19]/NET0131 , \ctl_rf_c5_rf_chdad_reg[1]/NET0131 , \ctl_rf_c5_rf_chdad_reg[20]/P0002 , \ctl_rf_c5_rf_chdad_reg[21]/P0002 , \ctl_rf_c5_rf_chdad_reg[22]/P0002 , \ctl_rf_c5_rf_chdad_reg[23]/P0002 , \ctl_rf_c5_rf_chdad_reg[24]/P0002 , \ctl_rf_c5_rf_chdad_reg[25]/P0002 , \ctl_rf_c5_rf_chdad_reg[26]/P0002 , \ctl_rf_c5_rf_chdad_reg[27]/P0002 , \ctl_rf_c5_rf_chdad_reg[28]/P0002 , \ctl_rf_c5_rf_chdad_reg[29]/P0002 , \ctl_rf_c5_rf_chdad_reg[2]/NET0131 , \ctl_rf_c5_rf_chdad_reg[30]/P0002 , \ctl_rf_c5_rf_chdad_reg[31]/P0002 , \ctl_rf_c5_rf_chdad_reg[3]/P0002 , \ctl_rf_c5_rf_chdad_reg[4]/P0002 , \ctl_rf_c5_rf_chdad_reg[5]/P0002 , \ctl_rf_c5_rf_chdad_reg[6]/P0002 , \ctl_rf_c5_rf_chdad_reg[7]/P0002 , \ctl_rf_c5_rf_chdad_reg[8]/NET0131 , \ctl_rf_c5_rf_chdad_reg[9]/P0002 , \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c5_rf_chllp_on_reg/NET0131 , \ctl_rf_c5_rf_chllp_reg[0]/P0002 , \ctl_rf_c5_rf_chllp_reg[10]/NET0131 , \ctl_rf_c5_rf_chllp_reg[11]/NET0131 , \ctl_rf_c5_rf_chllp_reg[12]/NET0131 , \ctl_rf_c5_rf_chllp_reg[13]/NET0131 , \ctl_rf_c5_rf_chllp_reg[14]/NET0131 , \ctl_rf_c5_rf_chllp_reg[15]/NET0131 , \ctl_rf_c5_rf_chllp_reg[16]/NET0131 , \ctl_rf_c5_rf_chllp_reg[17]/NET0131 , \ctl_rf_c5_rf_chllp_reg[18]/NET0131 , \ctl_rf_c5_rf_chllp_reg[19]/NET0131 , \ctl_rf_c5_rf_chllp_reg[1]/P0002 , \ctl_rf_c5_rf_chllp_reg[20]/NET0131 , \ctl_rf_c5_rf_chllp_reg[21]/NET0131 , \ctl_rf_c5_rf_chllp_reg[22]/NET0131 , \ctl_rf_c5_rf_chllp_reg[23]/NET0131 , \ctl_rf_c5_rf_chllp_reg[24]/NET0131 , \ctl_rf_c5_rf_chllp_reg[25]/NET0131 , \ctl_rf_c5_rf_chllp_reg[26]/NET0131 , \ctl_rf_c5_rf_chllp_reg[27]/NET0131 , \ctl_rf_c5_rf_chllp_reg[28]/NET0131 , \ctl_rf_c5_rf_chllp_reg[29]/NET0131 , \ctl_rf_c5_rf_chllp_reg[2]/NET0131 , \ctl_rf_c5_rf_chllp_reg[30]/NET0131 , \ctl_rf_c5_rf_chllp_reg[31]/NET0131 , \ctl_rf_c5_rf_chllp_reg[3]/NET0131 , \ctl_rf_c5_rf_chllp_reg[4]/NET0131 , \ctl_rf_c5_rf_chllp_reg[5]/NET0131 , \ctl_rf_c5_rf_chllp_reg[6]/NET0131 , \ctl_rf_c5_rf_chllp_reg[7]/NET0131 , \ctl_rf_c5_rf_chllp_reg[8]/NET0131 , \ctl_rf_c5_rf_chllp_reg[9]/NET0131 , \ctl_rf_c5_rf_chllpen_reg/NET0131 , \ctl_rf_c5_rf_chpri_reg[0]/NET0131 , \ctl_rf_c5_rf_chpri_reg[1]/NET0131 , \ctl_rf_c5_rf_chsad_reg[0]/NET0131 , \ctl_rf_c5_rf_chsad_reg[10]/NET0131 , \ctl_rf_c5_rf_chsad_reg[11]/NET0131 , \ctl_rf_c5_rf_chsad_reg[12]/NET0131 , \ctl_rf_c5_rf_chsad_reg[13]/P0002 , \ctl_rf_c5_rf_chsad_reg[14]/NET0131 , \ctl_rf_c5_rf_chsad_reg[15]/NET0131 , \ctl_rf_c5_rf_chsad_reg[16]/NET0131 , \ctl_rf_c5_rf_chsad_reg[17]/NET0131 , \ctl_rf_c5_rf_chsad_reg[18]/NET0131 , \ctl_rf_c5_rf_chsad_reg[19]/NET0131 , \ctl_rf_c5_rf_chsad_reg[1]/NET0131 , \ctl_rf_c5_rf_chsad_reg[20]/NET0131 , \ctl_rf_c5_rf_chsad_reg[21]/NET0131 , \ctl_rf_c5_rf_chsad_reg[22]/NET0131 , \ctl_rf_c5_rf_chsad_reg[23]/NET0131 , \ctl_rf_c5_rf_chsad_reg[24]/NET0131 , \ctl_rf_c5_rf_chsad_reg[25]/P0002 , \ctl_rf_c5_rf_chsad_reg[26]/P0002 , \ctl_rf_c5_rf_chsad_reg[27]/P0002 , \ctl_rf_c5_rf_chsad_reg[28]/P0002 , \ctl_rf_c5_rf_chsad_reg[29]/P0002 , \ctl_rf_c5_rf_chsad_reg[2]/NET0131 , \ctl_rf_c5_rf_chsad_reg[30]/P0002 , \ctl_rf_c5_rf_chsad_reg[31]/NET0131 , \ctl_rf_c5_rf_chsad_reg[3]/NET0131 , \ctl_rf_c5_rf_chsad_reg[4]/NET0131 , \ctl_rf_c5_rf_chsad_reg[5]/NET0131 , \ctl_rf_c5_rf_chsad_reg[6]/NET0131 , \ctl_rf_c5_rf_chsad_reg[7]/NET0131 , \ctl_rf_c5_rf_chsad_reg[8]/P0002 , \ctl_rf_c5_rf_chsad_reg[9]/NET0131 , \ctl_rf_c5_rf_chtsz_reg[0]/P0002 , \ctl_rf_c5_rf_chtsz_reg[10]/P0002 , \ctl_rf_c5_rf_chtsz_reg[11]/P0002 , \ctl_rf_c5_rf_chtsz_reg[1]/P0002 , \ctl_rf_c5_rf_chtsz_reg[2]/P0002 , \ctl_rf_c5_rf_chtsz_reg[3]/P0002 , \ctl_rf_c5_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c5_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c5_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c5_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c5_rf_chtsz_reg[8]/P0002 , \ctl_rf_c5_rf_chtsz_reg[9]/P0002 , \ctl_rf_c5_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c5_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c5_rf_dreqmode_reg/NET0131 , \ctl_rf_c5_rf_dst_sel_reg/NET0131 , \ctl_rf_c5_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c5_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c5_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c5_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c5_rf_int_err_msk_reg/NET0131 , \ctl_rf_c5_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c5_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c5_rf_mode_reg/NET0131 , \ctl_rf_c5_rf_prot1_reg/NET0131 , \ctl_rf_c5_rf_prot2_reg/NET0131 , \ctl_rf_c5_rf_prot3_reg/NET0131 , \ctl_rf_c5_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c5_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c5_rf_src_sel_reg/NET0131 , \ctl_rf_c5_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c5_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c5_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c5_rf_swidth_reg[0]/NET0131 , \ctl_rf_c5_rf_swidth_reg[1]/NET0131 , \ctl_rf_c5_rf_swidth_reg[2]/NET0131 , \ctl_rf_c5brbs_reg[16]/NET0131 , \ctl_rf_c5brbs_reg[17]/NET0131 , \ctl_rf_c5brbs_reg[18]/NET0131 , \ctl_rf_c5brbs_reg[19]/NET0131 , \ctl_rf_c5brbs_reg[20]/NET0131 , \ctl_rf_c5brbs_reg[21]/NET0131 , \ctl_rf_c5brbs_reg[22]/NET0131 , \ctl_rf_c5brbs_reg[23]/NET0131 , \ctl_rf_c5brbs_reg[24]/NET0131 , \ctl_rf_c5brbs_reg[25]/NET0131 , \ctl_rf_c5brbs_reg[26]/NET0131 , \ctl_rf_c5brbs_reg[27]/NET0131 , \ctl_rf_c5brbs_reg[28]/NET0131 , \ctl_rf_c5brbs_reg[29]/NET0131 , \ctl_rf_c5brbs_reg[30]/NET0131 , \ctl_rf_c5brbs_reg[31]/NET0131 , \ctl_rf_c5dmabs_reg[16]/NET0131 , \ctl_rf_c5dmabs_reg[17]/NET0131 , \ctl_rf_c5dmabs_reg[18]/NET0131 , \ctl_rf_c5dmabs_reg[19]/NET0131 , \ctl_rf_c5dmabs_reg[20]/NET0131 , \ctl_rf_c5dmabs_reg[21]/NET0131 , \ctl_rf_c5dmabs_reg[22]/NET0131 , \ctl_rf_c5dmabs_reg[23]/NET0131 , \ctl_rf_c5dmabs_reg[24]/NET0131 , \ctl_rf_c5dmabs_reg[25]/NET0131 , \ctl_rf_c5dmabs_reg[26]/NET0131 , \ctl_rf_c5dmabs_reg[27]/NET0131 , \ctl_rf_c5dmabs_reg[28]/NET0131 , \ctl_rf_c5dmabs_reg[29]/NET0131 , \ctl_rf_c5dmabs_reg[30]/NET0131 , \ctl_rf_c5dmabs_reg[31]/NET0131 , \ctl_rf_c6_rf_autold_reg/NET0131 , \ctl_rf_c6_rf_ch_en_reg/NET0131 , \ctl_rf_c6_rf_chabt_reg/NET0131 , \ctl_rf_c6_rf_chdad_reg[0]/NET0131 , \ctl_rf_c6_rf_chdad_reg[10]/NET0131 , \ctl_rf_c6_rf_chdad_reg[11]/P0002 , \ctl_rf_c6_rf_chdad_reg[12]/P0002 , \ctl_rf_c6_rf_chdad_reg[13]/NET0131 , \ctl_rf_c6_rf_chdad_reg[14]/P0002 , \ctl_rf_c6_rf_chdad_reg[15]/P0002 , \ctl_rf_c6_rf_chdad_reg[16]/NET0131 , \ctl_rf_c6_rf_chdad_reg[17]/NET0131 , \ctl_rf_c6_rf_chdad_reg[18]/NET0131 , \ctl_rf_c6_rf_chdad_reg[19]/NET0131 , \ctl_rf_c6_rf_chdad_reg[1]/NET0131 , \ctl_rf_c6_rf_chdad_reg[20]/P0002 , \ctl_rf_c6_rf_chdad_reg[21]/P0002 , \ctl_rf_c6_rf_chdad_reg[22]/P0002 , \ctl_rf_c6_rf_chdad_reg[23]/P0002 , \ctl_rf_c6_rf_chdad_reg[24]/P0002 , \ctl_rf_c6_rf_chdad_reg[25]/P0002 , \ctl_rf_c6_rf_chdad_reg[26]/P0002 , \ctl_rf_c6_rf_chdad_reg[27]/P0002 , \ctl_rf_c6_rf_chdad_reg[28]/P0002 , \ctl_rf_c6_rf_chdad_reg[29]/P0002 , \ctl_rf_c6_rf_chdad_reg[2]/NET0131 , \ctl_rf_c6_rf_chdad_reg[30]/P0002 , \ctl_rf_c6_rf_chdad_reg[31]/P0002 , \ctl_rf_c6_rf_chdad_reg[3]/P0002 , \ctl_rf_c6_rf_chdad_reg[4]/P0002 , \ctl_rf_c6_rf_chdad_reg[5]/P0002 , \ctl_rf_c6_rf_chdad_reg[6]/P0002 , \ctl_rf_c6_rf_chdad_reg[7]/P0002 , \ctl_rf_c6_rf_chdad_reg[8]/NET0131 , \ctl_rf_c6_rf_chdad_reg[9]/P0002 , \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c6_rf_chllp_on_reg/NET0131 , \ctl_rf_c6_rf_chllp_reg[0]/P0002 , \ctl_rf_c6_rf_chllp_reg[10]/NET0131 , \ctl_rf_c6_rf_chllp_reg[11]/NET0131 , \ctl_rf_c6_rf_chllp_reg[12]/NET0131 , \ctl_rf_c6_rf_chllp_reg[13]/NET0131 , \ctl_rf_c6_rf_chllp_reg[14]/NET0131 , \ctl_rf_c6_rf_chllp_reg[15]/NET0131 , \ctl_rf_c6_rf_chllp_reg[16]/NET0131 , \ctl_rf_c6_rf_chllp_reg[17]/NET0131 , \ctl_rf_c6_rf_chllp_reg[18]/NET0131 , \ctl_rf_c6_rf_chllp_reg[19]/NET0131 , \ctl_rf_c6_rf_chllp_reg[1]/P0002 , \ctl_rf_c6_rf_chllp_reg[20]/NET0131 , \ctl_rf_c6_rf_chllp_reg[21]/NET0131 , \ctl_rf_c6_rf_chllp_reg[22]/NET0131 , \ctl_rf_c6_rf_chllp_reg[23]/NET0131 , \ctl_rf_c6_rf_chllp_reg[24]/NET0131 , \ctl_rf_c6_rf_chllp_reg[25]/NET0131 , \ctl_rf_c6_rf_chllp_reg[26]/NET0131 , \ctl_rf_c6_rf_chllp_reg[27]/NET0131 , \ctl_rf_c6_rf_chllp_reg[28]/NET0131 , \ctl_rf_c6_rf_chllp_reg[29]/NET0131 , \ctl_rf_c6_rf_chllp_reg[2]/NET0131 , \ctl_rf_c6_rf_chllp_reg[30]/NET0131 , \ctl_rf_c6_rf_chllp_reg[31]/NET0131 , \ctl_rf_c6_rf_chllp_reg[3]/NET0131 , \ctl_rf_c6_rf_chllp_reg[4]/NET0131 , \ctl_rf_c6_rf_chllp_reg[5]/NET0131 , \ctl_rf_c6_rf_chllp_reg[6]/NET0131 , \ctl_rf_c6_rf_chllp_reg[7]/NET0131 , \ctl_rf_c6_rf_chllp_reg[8]/NET0131 , \ctl_rf_c6_rf_chllp_reg[9]/NET0131 , \ctl_rf_c6_rf_chllpen_reg/NET0131 , \ctl_rf_c6_rf_chpri_reg[0]/NET0131 , \ctl_rf_c6_rf_chpri_reg[1]/NET0131 , \ctl_rf_c6_rf_chsad_reg[0]/NET0131 , \ctl_rf_c6_rf_chsad_reg[10]/P0002 , \ctl_rf_c6_rf_chsad_reg[11]/NET0131 , \ctl_rf_c6_rf_chsad_reg[12]/NET0131 , \ctl_rf_c6_rf_chsad_reg[13]/P0002 , \ctl_rf_c6_rf_chsad_reg[14]/NET0131 , \ctl_rf_c6_rf_chsad_reg[15]/NET0131 , \ctl_rf_c6_rf_chsad_reg[16]/NET0131 , \ctl_rf_c6_rf_chsad_reg[17]/NET0131 , \ctl_rf_c6_rf_chsad_reg[18]/NET0131 , \ctl_rf_c6_rf_chsad_reg[19]/NET0131 , \ctl_rf_c6_rf_chsad_reg[1]/NET0131 , \ctl_rf_c6_rf_chsad_reg[20]/NET0131 , \ctl_rf_c6_rf_chsad_reg[21]/NET0131 , \ctl_rf_c6_rf_chsad_reg[22]/NET0131 , \ctl_rf_c6_rf_chsad_reg[23]/NET0131 , \ctl_rf_c6_rf_chsad_reg[24]/NET0131 , \ctl_rf_c6_rf_chsad_reg[25]/P0002 , \ctl_rf_c6_rf_chsad_reg[26]/P0002 , \ctl_rf_c6_rf_chsad_reg[27]/P0002 , \ctl_rf_c6_rf_chsad_reg[28]/P0002 , \ctl_rf_c6_rf_chsad_reg[29]/P0002 , \ctl_rf_c6_rf_chsad_reg[2]/NET0131 , \ctl_rf_c6_rf_chsad_reg[30]/P0002 , \ctl_rf_c6_rf_chsad_reg[31]/NET0131 , \ctl_rf_c6_rf_chsad_reg[3]/NET0131 , \ctl_rf_c6_rf_chsad_reg[4]/NET0131 , \ctl_rf_c6_rf_chsad_reg[5]/NET0131 , \ctl_rf_c6_rf_chsad_reg[6]/NET0131 , \ctl_rf_c6_rf_chsad_reg[7]/NET0131 , \ctl_rf_c6_rf_chsad_reg[8]/P0002 , \ctl_rf_c6_rf_chsad_reg[9]/NET0131 , \ctl_rf_c6_rf_chtsz_reg[0]/P0002 , \ctl_rf_c6_rf_chtsz_reg[10]/P0002 , \ctl_rf_c6_rf_chtsz_reg[11]/P0002 , \ctl_rf_c6_rf_chtsz_reg[1]/P0002 , \ctl_rf_c6_rf_chtsz_reg[2]/P0002 , \ctl_rf_c6_rf_chtsz_reg[3]/P0002 , \ctl_rf_c6_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c6_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c6_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c6_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c6_rf_chtsz_reg[8]/P0002 , \ctl_rf_c6_rf_chtsz_reg[9]/P0002 , \ctl_rf_c6_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c6_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c6_rf_dreqmode_reg/NET0131 , \ctl_rf_c6_rf_dst_sel_reg/NET0131 , \ctl_rf_c6_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c6_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c6_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c6_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c6_rf_int_err_msk_reg/NET0131 , \ctl_rf_c6_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c6_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c6_rf_mode_reg/NET0131 , \ctl_rf_c6_rf_prot1_reg/NET0131 , \ctl_rf_c6_rf_prot2_reg/NET0131 , \ctl_rf_c6_rf_prot3_reg/NET0131 , \ctl_rf_c6_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c6_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c6_rf_src_sel_reg/NET0131 , \ctl_rf_c6_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c6_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c6_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c6_rf_swidth_reg[0]/NET0131 , \ctl_rf_c6_rf_swidth_reg[1]/NET0131 , \ctl_rf_c6_rf_swidth_reg[2]/NET0131 , \ctl_rf_c6brbs_reg[16]/NET0131 , \ctl_rf_c6brbs_reg[17]/NET0131 , \ctl_rf_c6brbs_reg[18]/NET0131 , \ctl_rf_c6brbs_reg[19]/NET0131 , \ctl_rf_c6brbs_reg[20]/NET0131 , \ctl_rf_c6brbs_reg[21]/NET0131 , \ctl_rf_c6brbs_reg[22]/NET0131 , \ctl_rf_c6brbs_reg[23]/NET0131 , \ctl_rf_c6brbs_reg[24]/NET0131 , \ctl_rf_c6brbs_reg[25]/NET0131 , \ctl_rf_c6brbs_reg[26]/NET0131 , \ctl_rf_c6brbs_reg[27]/NET0131 , \ctl_rf_c6brbs_reg[28]/NET0131 , \ctl_rf_c6brbs_reg[29]/NET0131 , \ctl_rf_c6brbs_reg[30]/NET0131 , \ctl_rf_c6brbs_reg[31]/NET0131 , \ctl_rf_c6dmabs_reg[16]/NET0131 , \ctl_rf_c6dmabs_reg[17]/NET0131 , \ctl_rf_c6dmabs_reg[18]/NET0131 , \ctl_rf_c6dmabs_reg[19]/NET0131 , \ctl_rf_c6dmabs_reg[20]/NET0131 , \ctl_rf_c6dmabs_reg[21]/NET0131 , \ctl_rf_c6dmabs_reg[22]/NET0131 , \ctl_rf_c6dmabs_reg[23]/NET0131 , \ctl_rf_c6dmabs_reg[24]/NET0131 , \ctl_rf_c6dmabs_reg[25]/NET0131 , \ctl_rf_c6dmabs_reg[26]/NET0131 , \ctl_rf_c6dmabs_reg[27]/NET0131 , \ctl_rf_c6dmabs_reg[28]/NET0131 , \ctl_rf_c6dmabs_reg[29]/NET0131 , \ctl_rf_c6dmabs_reg[30]/NET0131 , \ctl_rf_c6dmabs_reg[31]/NET0131 , \ctl_rf_c7_rf_autold_reg/NET0131 , \ctl_rf_c7_rf_ch_en_reg/NET0131 , \ctl_rf_c7_rf_chabt_reg/NET0131 , \ctl_rf_c7_rf_chdad_reg[0]/NET0131 , \ctl_rf_c7_rf_chdad_reg[10]/P0002 , \ctl_rf_c7_rf_chdad_reg[11]/NET0131 , \ctl_rf_c7_rf_chdad_reg[12]/P0002 , \ctl_rf_c7_rf_chdad_reg[13]/NET0131 , \ctl_rf_c7_rf_chdad_reg[14]/NET0131 , \ctl_rf_c7_rf_chdad_reg[15]/NET0131 , \ctl_rf_c7_rf_chdad_reg[16]/NET0131 , \ctl_rf_c7_rf_chdad_reg[17]/NET0131 , \ctl_rf_c7_rf_chdad_reg[18]/NET0131 , \ctl_rf_c7_rf_chdad_reg[19]/NET0131 , \ctl_rf_c7_rf_chdad_reg[1]/NET0131 , \ctl_rf_c7_rf_chdad_reg[20]/P0002 , \ctl_rf_c7_rf_chdad_reg[21]/P0002 , \ctl_rf_c7_rf_chdad_reg[22]/P0002 , \ctl_rf_c7_rf_chdad_reg[23]/P0002 , \ctl_rf_c7_rf_chdad_reg[24]/P0002 , \ctl_rf_c7_rf_chdad_reg[25]/P0002 , \ctl_rf_c7_rf_chdad_reg[26]/P0002 , \ctl_rf_c7_rf_chdad_reg[27]/P0002 , \ctl_rf_c7_rf_chdad_reg[28]/P0002 , \ctl_rf_c7_rf_chdad_reg[29]/P0002 , \ctl_rf_c7_rf_chdad_reg[2]/NET0131 , \ctl_rf_c7_rf_chdad_reg[30]/P0002 , \ctl_rf_c7_rf_chdad_reg[31]/P0002 , \ctl_rf_c7_rf_chdad_reg[3]/P0002 , \ctl_rf_c7_rf_chdad_reg[4]/P0002 , \ctl_rf_c7_rf_chdad_reg[5]/P0002 , \ctl_rf_c7_rf_chdad_reg[6]/P0002 , \ctl_rf_c7_rf_chdad_reg[7]/P0002 , \ctl_rf_c7_rf_chdad_reg[8]/NET0131 , \ctl_rf_c7_rf_chdad_reg[9]/P0002 , \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131 , \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131 , \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131 , \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131 , \ctl_rf_c7_rf_chllp_on_reg/NET0131 , \ctl_rf_c7_rf_chllp_reg[0]/P0002 , \ctl_rf_c7_rf_chllp_reg[10]/NET0131 , \ctl_rf_c7_rf_chllp_reg[11]/NET0131 , \ctl_rf_c7_rf_chllp_reg[12]/NET0131 , \ctl_rf_c7_rf_chllp_reg[13]/NET0131 , \ctl_rf_c7_rf_chllp_reg[14]/NET0131 , \ctl_rf_c7_rf_chllp_reg[15]/NET0131 , \ctl_rf_c7_rf_chllp_reg[16]/NET0131 , \ctl_rf_c7_rf_chllp_reg[17]/NET0131 , \ctl_rf_c7_rf_chllp_reg[18]/NET0131 , \ctl_rf_c7_rf_chllp_reg[19]/NET0131 , \ctl_rf_c7_rf_chllp_reg[1]/P0002 , \ctl_rf_c7_rf_chllp_reg[20]/NET0131 , \ctl_rf_c7_rf_chllp_reg[21]/NET0131 , \ctl_rf_c7_rf_chllp_reg[22]/NET0131 , \ctl_rf_c7_rf_chllp_reg[23]/NET0131 , \ctl_rf_c7_rf_chllp_reg[24]/NET0131 , \ctl_rf_c7_rf_chllp_reg[25]/NET0131 , \ctl_rf_c7_rf_chllp_reg[26]/NET0131 , \ctl_rf_c7_rf_chllp_reg[27]/NET0131 , \ctl_rf_c7_rf_chllp_reg[28]/NET0131 , \ctl_rf_c7_rf_chllp_reg[29]/NET0131 , \ctl_rf_c7_rf_chllp_reg[2]/NET0131 , \ctl_rf_c7_rf_chllp_reg[30]/NET0131 , \ctl_rf_c7_rf_chllp_reg[31]/NET0131 , \ctl_rf_c7_rf_chllp_reg[3]/NET0131 , \ctl_rf_c7_rf_chllp_reg[4]/NET0131 , \ctl_rf_c7_rf_chllp_reg[5]/NET0131 , \ctl_rf_c7_rf_chllp_reg[6]/NET0131 , \ctl_rf_c7_rf_chllp_reg[7]/NET0131 , \ctl_rf_c7_rf_chllp_reg[8]/NET0131 , \ctl_rf_c7_rf_chllp_reg[9]/NET0131 , \ctl_rf_c7_rf_chllpen_reg/NET0131 , \ctl_rf_c7_rf_chpri_reg[0]/NET0131 , \ctl_rf_c7_rf_chpri_reg[1]/NET0131 , \ctl_rf_c7_rf_chsad_reg[0]/NET0131 , \ctl_rf_c7_rf_chsad_reg[10]/NET0131 , \ctl_rf_c7_rf_chsad_reg[11]/P0002 , \ctl_rf_c7_rf_chsad_reg[12]/NET0131 , \ctl_rf_c7_rf_chsad_reg[13]/P0002 , \ctl_rf_c7_rf_chsad_reg[14]/P0002 , \ctl_rf_c7_rf_chsad_reg[15]/P0002 , \ctl_rf_c7_rf_chsad_reg[16]/NET0131 , \ctl_rf_c7_rf_chsad_reg[17]/NET0131 , \ctl_rf_c7_rf_chsad_reg[18]/NET0131 , \ctl_rf_c7_rf_chsad_reg[19]/NET0131 , \ctl_rf_c7_rf_chsad_reg[1]/NET0131 , \ctl_rf_c7_rf_chsad_reg[20]/NET0131 , \ctl_rf_c7_rf_chsad_reg[21]/NET0131 , \ctl_rf_c7_rf_chsad_reg[22]/NET0131 , \ctl_rf_c7_rf_chsad_reg[23]/NET0131 , \ctl_rf_c7_rf_chsad_reg[24]/NET0131 , \ctl_rf_c7_rf_chsad_reg[25]/P0002 , \ctl_rf_c7_rf_chsad_reg[26]/P0002 , \ctl_rf_c7_rf_chsad_reg[27]/P0002 , \ctl_rf_c7_rf_chsad_reg[28]/P0002 , \ctl_rf_c7_rf_chsad_reg[29]/P0002 , \ctl_rf_c7_rf_chsad_reg[2]/NET0131 , \ctl_rf_c7_rf_chsad_reg[30]/P0002 , \ctl_rf_c7_rf_chsad_reg[31]/NET0131 , \ctl_rf_c7_rf_chsad_reg[3]/NET0131 , \ctl_rf_c7_rf_chsad_reg[4]/NET0131 , \ctl_rf_c7_rf_chsad_reg[5]/NET0131 , \ctl_rf_c7_rf_chsad_reg[6]/NET0131 , \ctl_rf_c7_rf_chsad_reg[7]/NET0131 , \ctl_rf_c7_rf_chsad_reg[8]/P0002 , \ctl_rf_c7_rf_chsad_reg[9]/NET0131 , \ctl_rf_c7_rf_chtsz_reg[0]/P0002 , \ctl_rf_c7_rf_chtsz_reg[10]/P0002 , \ctl_rf_c7_rf_chtsz_reg[11]/P0002 , \ctl_rf_c7_rf_chtsz_reg[1]/P0002 , \ctl_rf_c7_rf_chtsz_reg[2]/P0002 , \ctl_rf_c7_rf_chtsz_reg[3]/P0002 , \ctl_rf_c7_rf_chtsz_reg[4]/NET0131 , \ctl_rf_c7_rf_chtsz_reg[5]/NET0131 , \ctl_rf_c7_rf_chtsz_reg[6]/NET0131 , \ctl_rf_c7_rf_chtsz_reg[7]/NET0131 , \ctl_rf_c7_rf_chtsz_reg[8]/P0002 , \ctl_rf_c7_rf_chtsz_reg[9]/P0002 , \ctl_rf_c7_rf_dad_ctl0_reg/NET0131 , \ctl_rf_c7_rf_dad_ctl1_reg/NET0131 , \ctl_rf_c7_rf_dreqmode_reg/NET0131 , \ctl_rf_c7_rf_dst_sel_reg/NET0131 , \ctl_rf_c7_rf_dwidth_reg[0]/NET0131 , \ctl_rf_c7_rf_dwidth_reg[1]/NET0131 , \ctl_rf_c7_rf_dwidth_reg[2]/NET0131 , \ctl_rf_c7_rf_int_abt_msk_reg/NET0131 , \ctl_rf_c7_rf_int_err_msk_reg/NET0131 , \ctl_rf_c7_rf_int_tc1_msk_reg/NET0131 , \ctl_rf_c7_rf_int_tc_msk_reg/NET0131 , \ctl_rf_c7_rf_mode_reg/NET0131 , \ctl_rf_c7_rf_prot1_reg/NET0131 , \ctl_rf_c7_rf_prot2_reg/NET0131 , \ctl_rf_c7_rf_prot3_reg/NET0131 , \ctl_rf_c7_rf_sad_ctl0_reg/NET0131 , \ctl_rf_c7_rf_sad_ctl1_reg/NET0131 , \ctl_rf_c7_rf_src_sel_reg/NET0131 , \ctl_rf_c7_rf_src_sz_reg[0]/NET0131 , \ctl_rf_c7_rf_src_sz_reg[1]/NET0131 , \ctl_rf_c7_rf_src_sz_reg[2]/NET0131 , \ctl_rf_c7_rf_swidth_reg[0]/NET0131 , \ctl_rf_c7_rf_swidth_reg[1]/NET0131 , \ctl_rf_c7_rf_swidth_reg[2]/NET0131 , \ctl_rf_c7brbs_reg[16]/NET0131 , \ctl_rf_c7brbs_reg[17]/NET0131 , \ctl_rf_c7brbs_reg[18]/NET0131 , \ctl_rf_c7brbs_reg[19]/NET0131 , \ctl_rf_c7brbs_reg[20]/NET0131 , \ctl_rf_c7brbs_reg[21]/NET0131 , \ctl_rf_c7brbs_reg[22]/NET0131 , \ctl_rf_c7brbs_reg[23]/NET0131 , \ctl_rf_c7brbs_reg[24]/NET0131 , \ctl_rf_c7brbs_reg[25]/NET0131 , \ctl_rf_c7brbs_reg[26]/NET0131 , \ctl_rf_c7brbs_reg[27]/NET0131 , \ctl_rf_c7brbs_reg[28]/NET0131 , \ctl_rf_c7brbs_reg[29]/NET0131 , \ctl_rf_c7brbs_reg[30]/NET0131 , \ctl_rf_c7brbs_reg[31]/NET0131 , \ctl_rf_c7dmabs_reg[16]/NET0131 , \ctl_rf_c7dmabs_reg[17]/NET0131 , \ctl_rf_c7dmabs_reg[18]/NET0131 , \ctl_rf_c7dmabs_reg[19]/NET0131 , \ctl_rf_c7dmabs_reg[20]/NET0131 , \ctl_rf_c7dmabs_reg[21]/NET0131 , \ctl_rf_c7dmabs_reg[22]/NET0131 , \ctl_rf_c7dmabs_reg[23]/NET0131 , \ctl_rf_c7dmabs_reg[24]/NET0131 , \ctl_rf_c7dmabs_reg[25]/NET0131 , \ctl_rf_c7dmabs_reg[26]/NET0131 , \ctl_rf_c7dmabs_reg[27]/NET0131 , \ctl_rf_c7dmabs_reg[28]/NET0131 , \ctl_rf_c7dmabs_reg[29]/NET0131 , \ctl_rf_c7dmabs_reg[30]/NET0131 , \ctl_rf_c7dmabs_reg[31]/NET0131 , \ctl_rf_dmacen_reg/NET0131 , \ctl_rf_m0end_reg/NET0131 , \ctl_rf_m1end_reg/NET0131 , \ctl_rf_rf_sel_d1_reg/NET0131 , \ctl_rf_sync_reg[0]/NET0131 , \ctl_rf_sync_reg[1]/NET0131 , \ctl_rf_sync_reg[2]/NET0131 , \ctl_rf_sync_reg[3]/NET0131 , \ctl_rf_sync_reg[4]/NET0131 , \ctl_rf_sync_reg[5]/NET0131 , \ctl_rf_sync_reg[6]/NET0131 , \ctl_rf_sync_reg[7]/NET0131 , \ctl_rf_tc_reg[0]/NET0131 , \ctl_rf_tc_reg[1]/NET0131 , \ctl_rf_tc_reg[2]/NET0131 , \ctl_rf_tc_reg[3]/NET0131 , \ctl_rf_tc_reg[4]/NET0131 , \ctl_rf_tc_reg[5]/NET0131 , \ctl_rf_tc_reg[6]/NET0131 , \ctl_rf_tc_reg[7]/NET0131 , \de_bst_cnt_reg[0]/NET0131 , \de_bst_cnt_reg[2]/NET0131 , \de_bst_cnt_reg[3]/NET0131 , \de_bst_cnt_reg[4]/NET0131 , \de_bst_cnt_reg[5]/NET0131 , \de_bst_cnt_reg[6]/NET0131 , \de_bst_cnt_reg[7]/NET0131 , \de_bst_cnt_reg[8]/NET0131 , \de_de_st_reg[0]/NET0131 , \de_de_st_reg[1]/NET0131 , \de_de_st_reg[2]/NET0131 , \de_de_st_reg[5]/NET0131 , \de_de_st_reg[6]/NET0131 , \de_m0_arb_st_reg/NET0131 , \de_m0_is_llp_reg/NET0131 , \de_m1_arb_st_reg[0]/NET0131 , \de_m1_arb_st_reg[1]/NET0131 , \de_m1_is_llp_reg/NET0131 , \de_st_rd_msk_reg/NET0131 , \de_tsz_cnt_reg[0]/NET0131 , \de_tsz_cnt_reg[10]/NET0131 , \de_tsz_cnt_reg[11]/NET0131 , \de_tsz_cnt_reg[1]/NET0131 , \de_tsz_cnt_reg[2]/NET0131 , \de_tsz_cnt_reg[3]/NET0131 , \de_tsz_cnt_reg[4]/NET0131 , \de_tsz_cnt_reg[5]/NET0131 , \de_tsz_cnt_reg[6]/NET0131 , \de_tsz_cnt_reg[7]/NET0131 , \de_tsz_cnt_reg[8]/NET0131 , \de_tsz_cnt_reg[9]/NET0131 , \dma_ack[0]_pad , \dma_ack[1]_pad , \dma_ack[2]_pad , \dma_ack[3]_pad , \dma_ack[4]_pad , \dma_ack[5]_pad , \dma_ack[6]_pad , \dma_ack[7]_pad , \dma_tc[0]_pad , \dma_tc[1]_pad , \dma_tc[2]_pad , \dma_tc[3]_pad , \dma_tc[4]_pad , \dma_tc[5]_pad , \dma_tc[6]_pad , \dma_tc[7]_pad , \h0burst[0]_pad , \h0grant_pad , \h0readyin_pad , \h0req_pad , \h0resp[0]_pad , \h0resp[1]_pad , \h0write_pad , \h1burst[0]_pad , \h1prot[0]_pad , \h1rdt0_br[0]_pad , \h1rdt0_br[10]_pad , \h1rdt0_br[11]_pad , \h1rdt0_br[12]_pad , \h1rdt0_br[13]_pad , \h1rdt0_br[14]_pad , \h1rdt0_br[15]_pad , \h1rdt0_br[16]_pad , \h1rdt0_br[17]_pad , \h1rdt0_br[18]_pad , \h1rdt0_br[19]_pad , \h1rdt0_br[1]_pad , \h1rdt0_br[20]_pad , \h1rdt0_br[21]_pad , \h1rdt0_br[22]_pad , \h1rdt0_br[23]_pad , \h1rdt0_br[24]_pad , \h1rdt0_br[25]_pad , \h1rdt0_br[26]_pad , \h1rdt0_br[27]_pad , \h1rdt0_br[28]_pad , \h1rdt0_br[29]_pad , \h1rdt0_br[2]_pad , \h1rdt0_br[30]_pad , \h1rdt0_br[31]_pad , \h1rdt0_br[3]_pad , \h1rdt0_br[4]_pad , \h1rdt0_br[5]_pad , \h1rdt0_br[6]_pad , \h1rdt0_br[7]_pad , \h1rdt0_br[8]_pad , \h1rdt0_br[9]_pad , \h1rdt0_dma[0]_pad , \h1rdt0_dma[10]_pad , \h1rdt0_dma[11]_pad , \h1rdt0_dma[12]_pad , \h1rdt0_dma[13]_pad , \h1rdt0_dma[14]_pad , \h1rdt0_dma[15]_pad , \h1rdt0_dma[16]_pad , \h1rdt0_dma[17]_pad , \h1rdt0_dma[18]_pad , \h1rdt0_dma[19]_pad , \h1rdt0_dma[1]_pad , \h1rdt0_dma[20]_pad , \h1rdt0_dma[21]_pad , \h1rdt0_dma[22]_pad , \h1rdt0_dma[23]_pad , \h1rdt0_dma[24]_pad , \h1rdt0_dma[25]_pad , \h1rdt0_dma[26]_pad , \h1rdt0_dma[27]_pad , \h1rdt0_dma[28]_pad , \h1rdt0_dma[29]_pad , \h1rdt0_dma[2]_pad , \h1rdt0_dma[30]_pad , \h1rdt0_dma[31]_pad , \h1rdt0_dma[3]_pad , \h1rdt0_dma[4]_pad , \h1rdt0_dma[5]_pad , \h1rdt0_dma[6]_pad , \h1rdt0_dma[7]_pad , \h1rdt0_dma[8]_pad , \h1rdt0_dma[9]_pad , \h1rdt1_br[0]_pad , \h1rdt1_br[10]_pad , \h1rdt1_br[11]_pad , \h1rdt1_br[12]_pad , \h1rdt1_br[13]_pad , \h1rdt1_br[14]_pad , \h1rdt1_br[15]_pad , \h1rdt1_br[16]_pad , \h1rdt1_br[17]_pad , \h1rdt1_br[18]_pad , \h1rdt1_br[19]_pad , \h1rdt1_br[1]_pad , \h1rdt1_br[20]_pad , \h1rdt1_br[21]_pad , \h1rdt1_br[22]_pad , \h1rdt1_br[23]_pad , \h1rdt1_br[24]_pad , \h1rdt1_br[25]_pad , \h1rdt1_br[26]_pad , \h1rdt1_br[27]_pad , \h1rdt1_br[28]_pad , \h1rdt1_br[29]_pad , \h1rdt1_br[2]_pad , \h1rdt1_br[30]_pad , \h1rdt1_br[31]_pad , \h1rdt1_br[3]_pad , \h1rdt1_br[4]_pad , \h1rdt1_br[5]_pad , \h1rdt1_br[6]_pad , \h1rdt1_br[7]_pad , \h1rdt1_br[8]_pad , \h1rdt1_br[9]_pad , \h1rdt1_dma[0]_pad , \h1rdt1_dma[10]_pad , \h1rdt1_dma[11]_pad , \h1rdt1_dma[12]_pad , \h1rdt1_dma[13]_pad , \h1rdt1_dma[14]_pad , \h1rdt1_dma[15]_pad , \h1rdt1_dma[16]_pad , \h1rdt1_dma[17]_pad , \h1rdt1_dma[18]_pad , \h1rdt1_dma[19]_pad , \h1rdt1_dma[1]_pad , \h1rdt1_dma[20]_pad , \h1rdt1_dma[21]_pad , \h1rdt1_dma[22]_pad , \h1rdt1_dma[23]_pad , \h1rdt1_dma[24]_pad , \h1rdt1_dma[25]_pad , \h1rdt1_dma[26]_pad , \h1rdt1_dma[27]_pad , \h1rdt1_dma[28]_pad , \h1rdt1_dma[29]_pad , \h1rdt1_dma[2]_pad , \h1rdt1_dma[30]_pad , \h1rdt1_dma[31]_pad , \h1rdt1_dma[3]_pad , \h1rdt1_dma[4]_pad , \h1rdt1_dma[5]_pad , \h1rdt1_dma[6]_pad , \h1rdt1_dma[7]_pad , \h1rdt1_dma[8]_pad , \h1rdt1_dma[9]_pad , \h1rdt2_br[0]_pad , \h1rdt2_br[10]_pad , \h1rdt2_br[11]_pad , \h1rdt2_br[12]_pad , \h1rdt2_br[13]_pad , \h1rdt2_br[14]_pad , \h1rdt2_br[15]_pad , \h1rdt2_br[16]_pad , \h1rdt2_br[17]_pad , \h1rdt2_br[18]_pad , \h1rdt2_br[19]_pad , \h1rdt2_br[1]_pad , \h1rdt2_br[20]_pad , \h1rdt2_br[21]_pad , \h1rdt2_br[22]_pad , \h1rdt2_br[23]_pad , \h1rdt2_br[24]_pad , \h1rdt2_br[25]_pad , \h1rdt2_br[26]_pad , \h1rdt2_br[27]_pad , \h1rdt2_br[28]_pad , \h1rdt2_br[29]_pad , \h1rdt2_br[2]_pad , \h1rdt2_br[30]_pad , \h1rdt2_br[31]_pad , \h1rdt2_br[3]_pad , \h1rdt2_br[4]_pad , \h1rdt2_br[5]_pad , \h1rdt2_br[6]_pad , \h1rdt2_br[7]_pad , \h1rdt2_br[8]_pad , \h1rdt2_br[9]_pad , \h1rdt2_dma[0]_pad , \h1rdt2_dma[10]_pad , \h1rdt2_dma[11]_pad , \h1rdt2_dma[12]_pad , \h1rdt2_dma[13]_pad , \h1rdt2_dma[14]_pad , \h1rdt2_dma[15]_pad , \h1rdt2_dma[16]_pad , \h1rdt2_dma[17]_pad , \h1rdt2_dma[18]_pad , \h1rdt2_dma[19]_pad , \h1rdt2_dma[1]_pad , \h1rdt2_dma[20]_pad , \h1rdt2_dma[21]_pad , \h1rdt2_dma[22]_pad , \h1rdt2_dma[23]_pad , \h1rdt2_dma[24]_pad , \h1rdt2_dma[25]_pad , \h1rdt2_dma[26]_pad , \h1rdt2_dma[27]_pad , \h1rdt2_dma[28]_pad , \h1rdt2_dma[29]_pad , \h1rdt2_dma[2]_pad , \h1rdt2_dma[30]_pad , \h1rdt2_dma[31]_pad , \h1rdt2_dma[3]_pad , \h1rdt2_dma[4]_pad , \h1rdt2_dma[5]_pad , \h1rdt2_dma[6]_pad , \h1rdt2_dma[7]_pad , \h1rdt2_dma[8]_pad , \h1rdt2_dma[9]_pad , \h1rdt3_br[0]_pad , \h1rdt3_br[10]_pad , \h1rdt3_br[11]_pad , \h1rdt3_br[12]_pad , \h1rdt3_br[13]_pad , \h1rdt3_br[14]_pad , \h1rdt3_br[15]_pad , \h1rdt3_br[16]_pad , \h1rdt3_br[17]_pad , \h1rdt3_br[18]_pad , \h1rdt3_br[19]_pad , \h1rdt3_br[1]_pad , \h1rdt3_br[20]_pad , \h1rdt3_br[21]_pad , \h1rdt3_br[22]_pad , \h1rdt3_br[23]_pad , \h1rdt3_br[24]_pad , \h1rdt3_br[25]_pad , \h1rdt3_br[26]_pad , \h1rdt3_br[27]_pad , \h1rdt3_br[28]_pad , \h1rdt3_br[29]_pad , \h1rdt3_br[2]_pad , \h1rdt3_br[30]_pad , \h1rdt3_br[31]_pad , \h1rdt3_br[3]_pad , \h1rdt3_br[4]_pad , \h1rdt3_br[5]_pad , \h1rdt3_br[6]_pad , \h1rdt3_br[7]_pad , \h1rdt3_br[8]_pad , \h1rdt3_br[9]_pad , \h1rdt3_dma[0]_pad , \h1rdt3_dma[10]_pad , \h1rdt3_dma[11]_pad , \h1rdt3_dma[12]_pad , \h1rdt3_dma[13]_pad , \h1rdt3_dma[14]_pad , \h1rdt3_dma[15]_pad , \h1rdt3_dma[16]_pad , \h1rdt3_dma[17]_pad , \h1rdt3_dma[18]_pad , \h1rdt3_dma[19]_pad , \h1rdt3_dma[1]_pad , \h1rdt3_dma[20]_pad , \h1rdt3_dma[21]_pad , \h1rdt3_dma[22]_pad , \h1rdt3_dma[23]_pad , \h1rdt3_dma[24]_pad , \h1rdt3_dma[25]_pad , \h1rdt3_dma[26]_pad , \h1rdt3_dma[27]_pad , \h1rdt3_dma[28]_pad , \h1rdt3_dma[29]_pad , \h1rdt3_dma[2]_pad , \h1rdt3_dma[30]_pad , \h1rdt3_dma[31]_pad , \h1rdt3_dma[3]_pad , \h1rdt3_dma[4]_pad , \h1rdt3_dma[5]_pad , \h1rdt3_dma[6]_pad , \h1rdt3_dma[7]_pad , \h1rdt3_dma[8]_pad , \h1rdt3_dma[9]_pad , \h1rdt4_br[0]_pad , \h1rdt4_br[10]_pad , \h1rdt4_br[11]_pad , \h1rdt4_br[12]_pad , \h1rdt4_br[13]_pad , \h1rdt4_br[14]_pad , \h1rdt4_br[15]_pad , \h1rdt4_br[16]_pad , \h1rdt4_br[17]_pad , \h1rdt4_br[18]_pad , \h1rdt4_br[19]_pad , \h1rdt4_br[1]_pad , \h1rdt4_br[20]_pad , \h1rdt4_br[21]_pad , \h1rdt4_br[22]_pad , \h1rdt4_br[23]_pad , \h1rdt4_br[24]_pad , \h1rdt4_br[25]_pad , \h1rdt4_br[26]_pad , \h1rdt4_br[27]_pad , \h1rdt4_br[28]_pad , \h1rdt4_br[29]_pad , \h1rdt4_br[2]_pad , \h1rdt4_br[30]_pad , \h1rdt4_br[31]_pad , \h1rdt4_br[3]_pad , \h1rdt4_br[4]_pad , \h1rdt4_br[5]_pad , \h1rdt4_br[6]_pad , \h1rdt4_br[7]_pad , \h1rdt4_br[8]_pad , \h1rdt4_br[9]_pad , \h1rdt4_dma[0]_pad , \h1rdt4_dma[10]_pad , \h1rdt4_dma[11]_pad , \h1rdt4_dma[12]_pad , \h1rdt4_dma[13]_pad , \h1rdt4_dma[14]_pad , \h1rdt4_dma[15]_pad , \h1rdt4_dma[16]_pad , \h1rdt4_dma[17]_pad , \h1rdt4_dma[18]_pad , \h1rdt4_dma[19]_pad , \h1rdt4_dma[1]_pad , \h1rdt4_dma[20]_pad , \h1rdt4_dma[21]_pad , \h1rdt4_dma[22]_pad , \h1rdt4_dma[23]_pad , \h1rdt4_dma[24]_pad , \h1rdt4_dma[25]_pad , \h1rdt4_dma[26]_pad , \h1rdt4_dma[27]_pad , \h1rdt4_dma[28]_pad , \h1rdt4_dma[29]_pad , \h1rdt4_dma[2]_pad , \h1rdt4_dma[30]_pad , \h1rdt4_dma[31]_pad , \h1rdt4_dma[3]_pad , \h1rdt4_dma[4]_pad , \h1rdt4_dma[5]_pad , \h1rdt4_dma[6]_pad , \h1rdt4_dma[7]_pad , \h1rdt4_dma[8]_pad , \h1rdt4_dma[9]_pad , \h1rdt5_br[0]_pad , \h1rdt5_br[10]_pad , \h1rdt5_br[11]_pad , \h1rdt5_br[12]_pad , \h1rdt5_br[13]_pad , \h1rdt5_br[14]_pad , \h1rdt5_br[15]_pad , \h1rdt5_br[16]_pad , \h1rdt5_br[17]_pad , \h1rdt5_br[18]_pad , \h1rdt5_br[19]_pad , \h1rdt5_br[1]_pad , \h1rdt5_br[20]_pad , \h1rdt5_br[21]_pad , \h1rdt5_br[22]_pad , \h1rdt5_br[23]_pad , \h1rdt5_br[24]_pad , \h1rdt5_br[25]_pad , \h1rdt5_br[26]_pad , \h1rdt5_br[27]_pad , \h1rdt5_br[28]_pad , \h1rdt5_br[29]_pad , \h1rdt5_br[2]_pad , \h1rdt5_br[30]_pad , \h1rdt5_br[31]_pad , \h1rdt5_br[3]_pad , \h1rdt5_br[4]_pad , \h1rdt5_br[5]_pad , \h1rdt5_br[6]_pad , \h1rdt5_br[7]_pad , \h1rdt5_br[8]_pad , \h1rdt5_br[9]_pad , \h1rdt5_dma[0]_pad , \h1rdt5_dma[10]_pad , \h1rdt5_dma[11]_pad , \h1rdt5_dma[12]_pad , \h1rdt5_dma[13]_pad , \h1rdt5_dma[14]_pad , \h1rdt5_dma[15]_pad , \h1rdt5_dma[16]_pad , \h1rdt5_dma[17]_pad , \h1rdt5_dma[18]_pad , \h1rdt5_dma[19]_pad , \h1rdt5_dma[1]_pad , \h1rdt5_dma[20]_pad , \h1rdt5_dma[21]_pad , \h1rdt5_dma[22]_pad , \h1rdt5_dma[23]_pad , \h1rdt5_dma[24]_pad , \h1rdt5_dma[25]_pad , \h1rdt5_dma[26]_pad , \h1rdt5_dma[27]_pad , \h1rdt5_dma[28]_pad , \h1rdt5_dma[29]_pad , \h1rdt5_dma[2]_pad , \h1rdt5_dma[30]_pad , \h1rdt5_dma[31]_pad , \h1rdt5_dma[3]_pad , \h1rdt5_dma[4]_pad , \h1rdt5_dma[5]_pad , \h1rdt5_dma[6]_pad , \h1rdt5_dma[7]_pad , \h1rdt5_dma[8]_pad , \h1rdt5_dma[9]_pad , \h1rdt6_br[0]_pad , \h1rdt6_br[10]_pad , \h1rdt6_br[11]_pad , \h1rdt6_br[12]_pad , \h1rdt6_br[13]_pad , \h1rdt6_br[14]_pad , \h1rdt6_br[15]_pad , \h1rdt6_br[16]_pad , \h1rdt6_br[17]_pad , \h1rdt6_br[18]_pad , \h1rdt6_br[19]_pad , \h1rdt6_br[1]_pad , \h1rdt6_br[20]_pad , \h1rdt6_br[21]_pad , \h1rdt6_br[22]_pad , \h1rdt6_br[23]_pad , \h1rdt6_br[24]_pad , \h1rdt6_br[25]_pad , \h1rdt6_br[26]_pad , \h1rdt6_br[27]_pad , \h1rdt6_br[28]_pad , \h1rdt6_br[29]_pad , \h1rdt6_br[2]_pad , \h1rdt6_br[30]_pad , \h1rdt6_br[31]_pad , \h1rdt6_br[3]_pad , \h1rdt6_br[4]_pad , \h1rdt6_br[5]_pad , \h1rdt6_br[6]_pad , \h1rdt6_br[7]_pad , \h1rdt6_br[8]_pad , \h1rdt6_br[9]_pad , \h1rdt6_dma[0]_pad , \h1rdt6_dma[10]_pad , \h1rdt6_dma[11]_pad , \h1rdt6_dma[12]_pad , \h1rdt6_dma[13]_pad , \h1rdt6_dma[14]_pad , \h1rdt6_dma[15]_pad , \h1rdt6_dma[16]_pad , \h1rdt6_dma[17]_pad , \h1rdt6_dma[18]_pad , \h1rdt6_dma[19]_pad , \h1rdt6_dma[1]_pad , \h1rdt6_dma[20]_pad , \h1rdt6_dma[21]_pad , \h1rdt6_dma[22]_pad , \h1rdt6_dma[23]_pad , \h1rdt6_dma[24]_pad , \h1rdt6_dma[25]_pad , \h1rdt6_dma[26]_pad , \h1rdt6_dma[27]_pad , \h1rdt6_dma[28]_pad , \h1rdt6_dma[29]_pad , \h1rdt6_dma[2]_pad , \h1rdt6_dma[30]_pad , \h1rdt6_dma[31]_pad , \h1rdt6_dma[3]_pad , \h1rdt6_dma[4]_pad , \h1rdt6_dma[5]_pad , \h1rdt6_dma[6]_pad , \h1rdt6_dma[7]_pad , \h1rdt6_dma[8]_pad , \h1rdt6_dma[9]_pad , \h1rdt7_br[0]_pad , \h1rdt7_br[10]_pad , \h1rdt7_br[11]_pad , \h1rdt7_br[12]_pad , \h1rdt7_br[13]_pad , \h1rdt7_br[14]_pad , \h1rdt7_br[15]_pad , \h1rdt7_br[16]_pad , \h1rdt7_br[17]_pad , \h1rdt7_br[18]_pad , \h1rdt7_br[19]_pad , \h1rdt7_br[1]_pad , \h1rdt7_br[20]_pad , \h1rdt7_br[21]_pad , \h1rdt7_br[22]_pad , \h1rdt7_br[23]_pad , \h1rdt7_br[24]_pad , \h1rdt7_br[25]_pad , \h1rdt7_br[26]_pad , \h1rdt7_br[27]_pad , \h1rdt7_br[28]_pad , \h1rdt7_br[29]_pad , \h1rdt7_br[2]_pad , \h1rdt7_br[30]_pad , \h1rdt7_br[31]_pad , \h1rdt7_br[3]_pad , \h1rdt7_br[4]_pad , \h1rdt7_br[5]_pad , \h1rdt7_br[6]_pad , \h1rdt7_br[7]_pad , \h1rdt7_br[8]_pad , \h1rdt7_br[9]_pad , \h1rdt7_dma[0]_pad , \h1rdt7_dma[10]_pad , \h1rdt7_dma[11]_pad , \h1rdt7_dma[12]_pad , \h1rdt7_dma[13]_pad , \h1rdt7_dma[14]_pad , \h1rdt7_dma[15]_pad , \h1rdt7_dma[16]_pad , \h1rdt7_dma[17]_pad , \h1rdt7_dma[18]_pad , \h1rdt7_dma[19]_pad , \h1rdt7_dma[1]_pad , \h1rdt7_dma[20]_pad , \h1rdt7_dma[21]_pad , \h1rdt7_dma[22]_pad , \h1rdt7_dma[23]_pad , \h1rdt7_dma[24]_pad , \h1rdt7_dma[25]_pad , \h1rdt7_dma[26]_pad , \h1rdt7_dma[27]_pad , \h1rdt7_dma[28]_pad , \h1rdt7_dma[29]_pad , \h1rdt7_dma[2]_pad , \h1rdt7_dma[30]_pad , \h1rdt7_dma[31]_pad , \h1rdt7_dma[3]_pad , \h1rdt7_dma[4]_pad , \h1rdt7_dma[5]_pad , \h1rdt7_dma[6]_pad , \h1rdt7_dma[7]_pad , \h1rdt7_dma[8]_pad , \h1rdt7_dma[9]_pad , \h1rdy0_br_pad , \h1rdy0_dma_pad , \h1rdy1_br_pad , \h1rdy1_dma_pad , \h1rdy2_br_pad , \h1rdy2_dma_pad , \h1rdy3_br_pad , \h1rdy3_dma_pad , \h1rdy4_br_pad , \h1rdy4_dma_pad , \h1rdy5_br_pad , \h1rdy5_dma_pad , \h1rdy6_br_pad , \h1rdy6_dma_pad , \h1rdy7_br_pad , \h1rdy7_dma_pad , \h1rp0_br[0]_pad , \h1rp0_br[1]_pad , \h1rp0_dma[0]_pad , \h1rp0_dma[1]_pad , \h1rp1_br[0]_pad , \h1rp1_br[1]_pad , \h1rp1_dma[0]_pad , \h1rp1_dma[1]_pad , \h1rp2_br[0]_pad , \h1rp2_br[1]_pad , \h1rp2_dma[0]_pad , \h1rp2_dma[1]_pad , \h1rp3_br[0]_pad , \h1rp3_br[1]_pad , \h1rp3_dma[0]_pad , \h1rp3_dma[1]_pad , \h1rp4_br[0]_pad , \h1rp4_br[1]_pad , \h1rp4_dma[0]_pad , \h1rp4_dma[1]_pad , \h1rp5_br[0]_pad , \h1rp5_br[1]_pad , \h1rp5_dma[0]_pad , \h1rp5_dma[1]_pad , \h1rp6_br[0]_pad , \h1rp6_br[1]_pad , \h1rp6_dma[0]_pad , \h1rp6_dma[1]_pad , \h1rp7_br[0]_pad , \h1rp7_br[1]_pad , \h1rp7_dma[0]_pad , \h1rp7_dma[1]_pad , \h1size[0]_pad , \h1size[1]_pad , \h1size[2]_pad , \h1write_pad , \haddr[0]_pad , \haddr[1]_pad , \haddr[2]_pad , \haddr[3]_pad , \haddr[4]_pad , \haddr[5]_pad , \haddr[6]_pad , \haddr[7]_pad , \haddr[8]_pad , \hrdata_reg[0]_pad , \hrdata_reg[10]_pad , \hrdata_reg[11]_pad , \hrdata_reg[12]_pad , \hrdata_reg[13]_pad , \hrdata_reg[14]_pad , \hrdata_reg[15]_pad , \hrdata_reg[16]_pad , \hrdata_reg[17]_pad , \hrdata_reg[18]_pad , \hrdata_reg[19]_pad , \hrdata_reg[1]_pad , \hrdata_reg[20]_pad , \hrdata_reg[21]_pad , \hrdata_reg[22]_pad , \hrdata_reg[23]_pad , \hrdata_reg[24]_pad , \hrdata_reg[25]_pad , \hrdata_reg[26]_pad , \hrdata_reg[27]_pad , \hrdata_reg[28]_pad , \hrdata_reg[29]_pad , \hrdata_reg[2]_pad , \hrdata_reg[30]_pad , \hrdata_reg[31]_pad , \hrdata_reg[3]_pad , \hrdata_reg[4]_pad , \hrdata_reg[5]_pad , \hrdata_reg[6]_pad , \hrdata_reg[7]_pad , \hrdata_reg[8]_pad , \hrdata_reg[9]_pad , hreadyin_pad, hreadyout_br_pad, \hresp_br[0]_pad , \hresp_br[1]_pad , hsel_br_pad, hsel_reg_pad, \hsize[0]_pad , \hsize[1]_pad , \hsize[2]_pad , \htrans[0]_pad , \htrans[1]_pad , \hwdata[0]_pad , \hwdata[10]_pad , \hwdata[11]_pad , \hwdata[12]_pad , \hwdata[13]_pad , \hwdata[14]_pad , \hwdata[15]_pad , \hwdata[16]_pad , \hwdata[17]_pad , \hwdata[18]_pad , \hwdata[19]_pad , \hwdata[1]_pad , \hwdata[20]_pad , \hwdata[21]_pad , \hwdata[22]_pad , \hwdata[23]_pad , \hwdata[24]_pad , \hwdata[25]_pad , \hwdata[26]_pad , \hwdata[27]_pad , \hwdata[28]_pad , \hwdata[29]_pad , \hwdata[2]_pad , \hwdata[30]_pad , \hwdata[31]_pad , \hwdata[3]_pad , \hwdata[4]_pad , \hwdata[5]_pad , \hwdata[6]_pad , \hwdata[7]_pad , \hwdata[8]_pad , \hwdata[9]_pad , hwrite_pad, \m1_mux_hrdy_df_reg/NET0131 , \m1_mux_hrmxnof_reg/NET0131 , \m1_mux_hrp_df_reg[0]/NET0131 , \m1_mux_mux_no_reg[0]/NET0131 , \m1_mux_mux_no_reg[1]/NET0131 , \m1_mux_mux_no_reg[2]/NET0131 , \m1_mux_mux_no_reg[3]/NET0131 , \_al_n1 , \g16/_0_ , \g58487/_0_ , \g58489/_0_ , \g58491/_0_ , \g58493/_0_ , \g58495/_0_ , \g58497/_0_ , \g58499/_0_ , \g58500/_0_ , \g58501/_0_ , \g58502/_0_ , \g58504/_0_ , \g58505/_0_ , \g58507/_0_ , \g58508/_0_ , \g58509/_0_ , \g58510/_0_ , \g58556/_0_ , \g58557/_0_ , \g58558/_0_ , \g58559/_0_ , \g58560/_0_ , \g58561/_0_ , \g58562/_0_ , \g58563/_0_ , \g58566/_0_ , \g58567/_0_ , \g58568/_0_ , \g58569/_0_ , \g58570/_0_ , \g58571/_0_ , \g58572/_0_ , \g58573/_0_ , \g58574/_0_ , \g58575/_0_ , \g58576/_0_ , \g58577/_0_ , \g58578/_0_ , \g58579/_0_ , \g58580/_0_ , \g58581/_0_ , \g58584/_0_ , \g58585/_0_ , \g58586/_0_ , \g58587/_0_ , \g58588/_0_ , \g58589/_0_ , \g58590/_0_ , \g58591/_0_ , \g58592/_0_ , \g58593/_0_ , \g58594/_0_ , \g58595/_0_ , \g58596/_0_ , \g58597/_0_ , \g58598/_0_ , \g58599/_0_ , \g58600/_0_ , \g58601/_0_ , \g58602/_0_ , \g58603/_0_ , \g58604/_0_ , \g58605/_0_ , \g58606/_0_ , \g58607/_0_ , \g58608/_0_ , \g58609/_0_ , \g58610/_0_ , \g58611/_0_ , \g58612/_0_ , \g58613/_0_ , \g58614/_0_ , \g58615/_0_ , \g58616/_0_ , \g58617/_0_ , \g58618/_0_ , \g58619/_0_ , \g58620/_0_ , \g58621/_0_ , \g58622/_0_ , \g58623/_0_ , \g58624/_0_ , \g58625/_0_ , \g58626/_0_ , \g58627/_0_ , \g58723/_0_ , \g58734/_0_ , \g58737/_0_ , \g58741/_0_ , \g58749/_0_ , \g58754/_0_ , \g58762/_0_ , \g58763/_0_ , \g58764/_0_ , \g58765/_0_ , \g58766/_0_ , \g58767/_0_ , \g58768/_0_ , \g58769/_0_ , \g58770/_0_ , \g58771/_0_ , \g59788/_0_ , \g59832/_0_ , \g59873/_0_ , \g59874/_0_ , \g59893/_0_ , \g59894/_0_ , \g59895/_0_ , \g59896/_0_ , \g59923/_0_ , \g60031/_0_ , \g60032/_0_ , \g60033/_0_ , \g60036/_0_ , \g60037/_0_ , \g60038/_0_ , \g60165/_0_ , \g60186/_2__syn_2 , \g60187/_0_ , \g60188/_0_ , \g60258/_0_ , \g60259/_0_ , \g60260/_0_ , \g60261/_0_ , \g60263/_0_ , \g60264/_0_ , \g60265/_0_ , \g60266/_0_ , \g60267/_0_ , \g60303/_3_ , \g60360/_0_ , \g60361/_0_ , \g60401/_00_ , \g60428/_0_ , \g60429/_0_ , \g60448/_0_ , \g60449/_0_ , \g60974/_0_ , \g61072/_0_ , \g61073/_0_ , \g61074/_0_ , \g61075/_0_ , \g61076/_0_ , \g61077/_0_ , \g61078/_0_ , \g61079/_0_ , \g61486/_0_ , \g61502/_3_ , \g61879/_0_ , \g62077/_0_ , \g62078/_0_ , \g62079/_0_ , \g62080/_0_ , \g62081/_0_ , \g62082/_0_ , \g62083/_0_ , \g62084/_0_ , \g62085/_0_ , \g62086/_0_ , \g62087/_0_ , \g62088/_0_ , \g62089/_0_ , \g62090/_0_ , \g62091/_0_ , \g62629/_0_ , \g62630/_0_ , \g62631/_0_ , \g62632/_0_ , \g62633/_0_ , \g62634/_0_ , \g62635/_0_ , \g62637/_0_ , \g62638/_0_ , \g62639/_0_ , \g62641/_0_ , \g62643/_0_ , \g62645/_0_ , \g62646/_0_ , \g62647/_0_ , \g62648/_0_ , \g62649/_0_ , \g62650/_0_ , \g62651/_0_ , \g62652/_0_ , \g62655/_0_ , \g62656/_0_ , \g62657/_0_ , \g62658/_0_ , \g62659/_0_ , \g62660/_0_ , \g62661/_0_ , \g62662/_0_ , \g62663/_0_ , \g62664/_0_ , \g62665/_0_ , \g62667/_0_ , \g62668/_0_ , \g62669/_0_ , \g62670/_0_ , \g62671/_0_ , \g62672/_0_ , \g62673/_0_ , \g62674/_0_ , \g62675/_0_ , \g62676/_0_ , \g62677/_0_ , \g62678/_0_ , \g62679/_0_ , \g62680/_0_ , \g62681/_0_ , \g62682/_0_ , \g62683/_0_ , \g62684/_0_ , \g62685/_0_ , \g62686/_0_ , \g62687/_0_ , \g62688/_0_ , \g62689/_0_ , \g62690/_0_ , \g62691/_0_ , \g62692/_0_ , \g62693/_0_ , \g62694/_0_ , \g62695/_0_ , \g62696/_0_ , \g62697/_0_ , \g62698/_0_ , \g62699/_0_ , \g62700/_0_ , \g62701/_0_ , \g62702/_0_ , \g62703/_0_ , \g62704/_0_ , \g62705/_0_ , \g62706/_0_ , \g62707/_0_ , \g62708/_0_ , \g62709/_0_ , \g62710/_0_ , \g62711/_0_ , \g62712/_0_ , \g62713/_0_ , \g62714/_0_ , \g62715/_0_ , \g62716/_0_ , \g62721/_0_ , \g62722/_0_ , \g62723/_0_ , \g62725/_0_ , \g62726/_0_ , \g62727/_0_ , \g62728/_0_ , \g62729/_0_ , \g62730/_0_ , \g62731/_0_ , \g62732/_0_ , \g62733/_0_ , \g62734/_0_ , \g62735/_0_ , \g62736/_0_ , \g62737/_0_ , \g62738/_0_ , \g62739/_0_ , \g62740/_0_ , \g62741/_0_ , \g62742/_0_ , \g62743/_0_ , \g62744/_0_ , \g62745/_0_ , \g62746/_0_ , \g62747/_0_ , \g62748/_0_ , \g62749/_0_ , \g62750/_0_ , \g62751/_0_ , \g62752/_0_ , \g62753/_0_ , \g62754/_0_ , \g62755/_0_ , \g62756/_0_ , \g62757/_0_ , \g62758/_0_ , \g62759/_0_ , \g62760/_0_ , \g62761/_0_ , \g62762/_0_ , \g62763/_0_ , \g62764/_0_ , \g62765/_0_ , \g62766/_0_ , \g62767/_0_ , \g62768/_0_ , \g62769/_0_ , \g62770/_0_ , \g62771/_0_ , \g62772/_0_ , \g62773/_0_ , \g62774/_0_ , \g62775/_0_ , \g62776/_0_ , \g62777/_0_ , \g62778/_0_ , \g62779/_0_ , \g62780/_0_ , \g62781/_0_ , \g62783/_0_ , \g62784/_0_ , \g62785/_0_ , \g62786/_0_ , \g62787/_0_ , \g62788/_0_ , \g62789/_0_ , \g62790/_0_ , \g62791/_0_ , \g62792/_0_ , \g62793/_0_ , \g62794/_0_ , \g62795/_0_ , \g62797/_0_ , \g62798/_0_ , \g62799/_0_ , \g62800/_0_ , \g62801/_0_ , \g62802/_0_ , \g62803/_0_ , \g62804/_0_ , \g62805/_0_ , \g62806/_0_ , \g62807/_0_ , \g62808/_0_ , \g62809/_0_ , \g62810/_0_ , \g62811/_0_ , \g62812/_0_ , \g62813/_0_ , \g62814/_0_ , \g62815/_0_ , \g62816/_0_ , \g62817/_0_ , \g62818/_0_ , \g63108/_0_ , \g63117/_0_ , \g63125/_0_ , \g63126/_0_ , \g63127/_0_ , \g63128/_0_ , \g63129/_0_ , \g63130/_0_ , \g63131/_0_ , \g63132/_0_ , \g63133/_0_ , \g63134/_0_ , \g63135/_0_ , \g63136/_0_ , \g63137/_0_ , \g63138/_0_ , \g63139/_0_ , \g63140/_0_ , \g63141/_0_ , \g63142/_0_ , \g63143/_0_ , \g63144/_0_ , \g63145/_0_ , \g63146/_0_ , \g63147/_0_ , \g63148/_0_ , \g63149/_0_ , \g63150/_0_ , \g63151/_0_ , \g63152/_0_ , \g63153/_0_ , \g63154/_0_ , \g63155/_0_ , \g63156/_0_ , \g63157/_0_ , \g63159/_0_ , \g63160/_0_ , \g63161/_0_ , \g63162/_0_ , \g63163/_0_ , \g63164/_0_ , \g63165/_0_ , \g63166/_0_ , \g63167/_0_ , \g63168/_0_ , \g63169/_0_ , \g63170/_0_ , \g63171/_0_ , \g63172/_0_ , \g63173/_0_ , \g63174/_0_ , \g63175/_0_ , \g63176/_0_ , \g63177/_0_ , \g63178/_0_ , \g63179/_0_ , \g63180/_0_ , \g63181/_0_ , \g63182/_0_ , \g63183/_0_ , \g63184/_0_ , \g63185/_0_ , \g63186/_0_ , \g63187/_0_ , \g63188/_0_ , \g63189/_0_ , \g63190/_0_ , \g63191/_0_ , \g63192/_0_ , \g63193/_0_ , \g63194/_0_ , \g63195/_0_ , \g63196/_0_ , \g63197/_0_ , \g63198/_0_ , \g63199/_0_ , \g63200/_0_ , \g63201/_0_ , \g63202/_0_ , \g63203/_0_ , \g63204/_0_ , \g63205/_0_ , \g63206/_0_ , \g63207/_0_ , \g63208/_0_ , \g63209/_0_ , \g63210/_0_ , \g63211/_0_ , \g63212/_0_ , \g63213/_0_ , \g63214/_0_ , \g63215/_0_ , \g63216/_0_ , \g63217/_0_ , \g63218/_0_ , \g63219/_0_ , \g63220/_0_ , \g63221/_0_ , \g63222/_0_ , \g63223/_0_ , \g63224/_0_ , \g63225/_0_ , \g63226/_0_ , \g63228/_0_ , \g63229/_0_ , \g63231/_0_ , \g63232/_0_ , \g63233/_0_ , \g63234/_0_ , \g63235/_0_ , \g63236/_0_ , \g63237/_0_ , \g63238/_0_ , \g63239/_0_ , \g63240/_0_ , \g63241/_0_ , \g63242/_0_ , \g63244/_0_ , \g63246/_0_ , \g63247/_0_ , \g63248/_0_ , \g63249/_0_ , \g63250/_0_ , \g63251/_0_ , \g63252/_0_ , \g63253/_0_ , \g63254/_0_ , \g63255/_0_ , \g63256/_0_ , \g63257/_0_ , \g63258/_0_ , \g63259/_0_ , \g63260/_0_ , \g63261/_0_ , \g63262/_0_ , \g63263/_0_ , \g63264/_0_ , \g63265/_0_ , \g63266/_0_ , \g63267/_0_ , \g63268/_0_ , \g63269/_0_ , \g63270/_0_ , \g63272/_0_ , \g63291/_0_ , \g63292/_0_ , \g63293/_0_ , \g63294/_0_ , \g63295/_0_ , \g63298/_0_ , \g63299/_0_ , \g63300/_0_ , \g63301/_0_ , \g63302/_0_ , \g63303/_0_ , \g63304/_0_ , \g63305/_0_ , \g63306/_0_ , \g63307/_0_ , \g63308/_0_ , \g63309/_0_ , \g63310/_0_ , \g63311/_0_ , \g63312/_0_ , \g63313/_0_ , \g63314/_0_ , \g63315/_0_ , \g63316/_0_ , \g63317/_0_ , \g63318/_0_ , \g63320/_0_ , \g63322/_0_ , \g63323/_0_ , \g63324/_0_ , \g63325/_0_ , \g63326/_0_ , \g63327/_0_ , \g63328/_0_ , \g63329/_0_ , \g63330/_0_ , \g63331/_0_ , \g63332/_0_ , \g63333/_0_ , \g63334/_0_ , \g63335/_0_ , \g63336/_0_ , \g63337/_0_ , \g63338/_0_ , \g63339/_0_ , \g63340/_0_ , \g63341/_0_ , \g63342/_0_ , \g63343/_0_ , \g63344/_0_ , \g63345/_0_ , \g63346/_0_ , \g63347/_0_ , \g63348/_0_ , \g63349/_0_ , \g63350/_0_ , \g63351/_0_ , \g63352/_0_ , \g63353/_0_ , \g63354/_0_ , \g63355/_0_ , \g63356/_0_ , \g63357/_0_ , \g63358/_0_ , \g63359/_0_ , \g63360/_0_ , \g63361/_0_ , \g63362/_0_ , \g63363/_0_ , \g63364/_0_ , \g63365/_0_ , \g63366/_0_ , \g63367/_0_ , \g63368/_0_ , \g63369/_0_ , \g63370/_0_ , \g63371/_0_ , \g63372/_0_ , \g63373/_0_ , \g63374/_0_ , \g63375/_0_ , \g63376/_0_ , \g63377/_0_ , \g63378/_0_ , \g63379/_0_ , \g63380/_0_ , \g63383/_3_ , \g63386/_0_ , \g63387/_0_ , \g63388/_0_ , \g63389/_0_ , \g63390/_0_ , \g63391/_0_ , \g63392/_0_ , \g63419/_0_ , \g63421/_0_ , \g63422/_0_ , \g63423/_0_ , \g63424/_0_ , \g63425/_0_ , \g63536/_3_ , \g63625/_0_ , \g63628/_0_ , \g63871/_0_ , \g63874/_0_ , \g63889/_0_ , \g63933/_0_ , \g63945/_0_ , \g63959/_0_ , \g63962/_0_ , \g63974/_0_ , \g63977/_0_ , \g64035/_0_ , \g64435/_3_ , \g64939/_0_ , \g65149/_0_ , \g65632/_3_ , \g65633/_0_ , \g65634/_0_ , \g65635/_0_ , \g65636/_0_ , \g65638/_3_ , \g65640/_3_ , \g65999/_0_ , \g66912/_0_ , \g66914/_0_ , \g67555/_3_ , \g67564/_3_ , \g67567/_3_ , \g67735/_0_ , \g67736/_0_ , \g67737/_0_ , \g67738/_0_ , \g67758/_0_ , \g67760/_0_ , \g67761/_0_ , \g67763/_0_ , \g67766/_0_ , \g67810/_0_ , \g67816/_0_ , \g67902/_0_ , \g67927/_0_ , \g67936/_0_ , \g68067/_0_ , \g68068/_0_ , \g68069/_0_ , \g68070/_0_ , \g68071/_0_ , \g68072/_0_ , \g68073/_0_ , \g68074/_0_ , \g68075/_0_ , \g68076/_0_ , \g68077/_0_ , \g68078/_0_ , \g68079/_0_ , \g68080/_0_ , \g68081/_0_ , \g68082/_0_ , \g68083/_0_ , \g68084/_0_ , \g68085/_0_ , \g68086/_0_ , \g68087/_0_ , \g68088/_0_ , \g68089/_0_ , \g68090/_0_ , \g68091/_0_ , \g68096/_0_ , \g68160/_0_ , \g68218/_0_ , \g68219/_0_ , \g68220/_0_ , \g68221/_0_ , \g68222/_0_ , \g68226/_0_ , \g68247/_0_ , \g68252/_0_ , \g68632/_0_ , \g68633/_0_ , \g68635/_0_ , \g68640/_0_ , \g68642/_0_ , \g68643/_0_ , \g68644/_0_ , \g68645/_0_ , \g68649/_0_ , \g68668/_2_ , \g68670/_0_ , \g68681/_3_ , \g68689/_0_ , \g68690/_0_ , \g68691/_0_ , \g68692/_0_ , \g68693/_0_ , \g68694/_0_ , \g68695/_0_ , \g68737/_0_ , \g68742/_0_ , \g68745/_0_ , \g68750/_0_ , \g68759/_0_ , \g68761/_0_ , \g68774/_0_ , \g68775/_0_ , \g68776/_0_ , \g68777/_0_ , \g68778/_0_ , \g68780/_0_ , \g68781/_0_ , \g68782/_0_ , \g68783/_0_ , \g68784/_0_ , \g68785/_0_ , \g68786/_0_ , \g68787/_0_ , \g68790/_0_ , \g68791/_0_ , \g68793/_0_ , \g68794/_0_ , \g68795/_0_ , \g68796/_0_ , \g68797/_0_ , \g68804/_0_ , \g68805/_0_ , \g68807/_0_ , \g68809/_0_ , \g68864/_3_ , \g68865/_3_ , \g68866/_3_ , \g68867/_3_ , \g68868/_3_ , \g68869/_3_ , \g68870/_3_ , \g68871/_3_ , \g68872/_3_ , \g68873/_3_ , \g68874/_3_ , \g68875/_3_ , \g68876/_3_ , \g68877/_3_ , \g68878/_3_ , \g68879/_3_ , \g68880/_3_ , \g68881/_3_ , \g68882/_3_ , \g68883/_3_ , \g68884/_3_ , \g68885/_3_ , \g68886/_3_ , \g68887/_3_ , \g68888/_3_ , \g68889/_3_ , \g68890/_3_ , \g68891/_3_ , \g68892/_3_ , \g68893/_3_ , \g68894/_3_ , \g68895/_3_ , \g69037/_1__syn_2 , \g69077/_0_ , \g69081/_0_ , \g69084/_0_ , \g69085/_0_ , \g69086/_0_ , \g69088/_0_ , \g69094/_0_ , \g69095/_0_ , \g69097/_0_ , \g69114/_3_ , \g69116/_3_ , \g69118/_3_ , \g69120/_3_ , \g69122/_3_ , \g69124/_3_ , \g69126/_3_ , \g69128/_3_ , \g69581/_3_ , \g70303/_1__syn_2 , \g70304/_1__syn_2 , \g70305/_1__syn_2 , \g70306/_1__syn_2 , \g70353/_1__syn_2 , \g70359/_2_ , \g70364/_1__syn_2 , \g70375/_1__syn_2 , \g70380/_2_ , \g70383/_1__syn_2 , \g70394/_2_ , \g70395/_2_ , \g70396/_1__syn_2 , \g70398/_1__syn_2 , \g70407/_1_ , \g70416/_1__syn_2 , \g70418/_1__syn_2 , \g70419/_2_ , \g70424/_1_ , \g70465/_2_ , \g70511/_1_ , \g70512/_1_ , \g70513/_2_ , \g70514/_2_ , \g70516/_2_ , \g70518/_2_ , \g70519/_2_ , \g70520/_2_ , \g70530/_2_ , \g70534/_3_ , \g70536/_3_ , \g70540/_3_ , \g70541/_2_ , \g70545/_3_ , \g70546/_2_ , \g70547/_2_ , \g70550/_3_ , \g70551/_2_ , \g70552/_2_ , \g70558/_3_ , \g70559/_2_ , \g70560/_2_ , \g70562/_3_ , \g70564/_3_ , \g70567/_3_ , \g70568/_2_ , \g70571/_3_ , \g70577/_0_ , \g70578/_2_ , \g70585/_3_ , \g70586/_2_ , \g70587/_2_ , \g70588/_3_ , \g70602/_3_ , \g70841/_0_ , \g70842/_0_ , \g70843/_0_ , \g70844/_0_ , \g70845/_0_ , \g70846/_0_ , \g70847/_0_ , \g70848/_0_ , \g70849/_0_ , \g70850/_0_ , \g70851/_0_ , \g70852/_0_ , \g70853/_0_ , \g70854/_0_ , \g70855/_0_ , \g70856/_0_ , \g70857/_0_ , \g70858/_0_ , \g70859/_0_ , \g70860/_0_ , \g70861/_0_ , \g70862/_0_ , \g70863/_0_ , \g70864/_0_ , \g70865/_0_ , \g70866/_0_ , \g70867/_0_ , \g70868/_0_ , \g70869/_0_ , \g70870/_0_ , \g70871/_0_ , \g70872/_0_ , \g70944/_1__syn_2 , \g71042/_1__syn_2 , \g71064/_1__syn_2 , \g71065/_1__syn_2 , \g71076/_1__syn_2 , \g71077/_1__syn_2 , \g71202/_1__syn_2 , \g71204/_1__syn_2 , \g71236/_0_ , \g71237/_0_ , \g71241/_0_ , \g71242/_0_ , \g71245/_0_ , \g71246/_0_ , \g71306/_0_ , \g71308/_0_ , \g71309/_0_ , \g71310/_0_ , \g71355/_0_ , \g71416/_0_ , \g71417/_0_ , \g71420/_0_ , \g71432/_0_ , \g71434/_0_ , \g71435/_0_ , \g71436/_0_ , \g71446/_0_ , \g71449/_0_ , \g71451/_0_ , \g71452/_0_ , \g71485/_0_ , \g71494/_0_ , \g71499/_0_ , \g71500/_0_ , \g71501/_0_ , \g71502/_0_ , \g71503/_0_ , \g71504/_0_ , \g71505/_0_ , \g71506/_0_ , \g71815/_0_ , \g71823/_0_ , \g71832/_0_ , \g71833/_0__syn_2 , \g71837/_0_ , \g71838/_0_ , \g71846/_1__syn_2 , \g71847/_1__syn_2 , \g71849/_0_ , \g71854/_0_ , \g71858/_1__syn_2 , \g71859/_1__syn_2 , \g71863/_0_ , \g71867/_0_ , \g71869/_0_ , \g71872/_1_ , \g71873/_1__syn_2 , \g71874/_1__syn_2 , \g71875/_0_ , \g71877/_1__syn_2 , \g71881/_0_ , \g71906/_0_ , \g71907/_1__syn_2 , \g71910/_0_ , \g71911/_0_ , \g71912/_1__syn_2 , \g71913/_1__syn_2 , \g71914/_1__syn_2 , \g71918/_0_ , \g71921/_0_ , \g71922/_0_ , \g71929/_1__syn_2 , \g71931/_1__syn_2 , \g71938/_1__syn_2 , \g71942/_0_ , \g71946/_1__syn_2 , \g71947/_0_ , \g71951/_0_ , \g71958/_1__syn_2 , \g71965/_0_ , \g71970/_1__syn_2 , \g71972/_1__syn_2 , \g71973/_1__syn_2 , \g71986/_1__syn_2 , \g71987/_1__syn_2 , \g71990/_1__syn_2 , \g71991/_1__syn_2 , \g71992/_1__syn_2 , \g71994/_1__syn_2 , \g71997/_1__syn_2 , \g72001/_1__syn_2 , \g72013/_1__syn_2 , \g72021/_1__syn_2 , \g72030/_0_ , \g72031/_0__syn_2 , \g72036/_1__syn_2 , \g72038/_0_ , \g72042/_1__syn_2 , \g72047/_1__syn_2 , \g72048/_1__syn_2 , \g72049/_1__syn_2 , \g72056/_0_ , \g72064/_1__syn_2 , \g72073/_1__syn_2 , \g72075/_0_ , \g72078/_0_ , \g72081/_0_ , \g72091/_0_ , \g72096/_0_ , \g72100/_1__syn_2 , \g72113/_0_ , \g72118/_0_ , \g72121/_1__syn_2 , \g72122/_1__syn_2 , \g72125/_1__syn_2 , \g72128/_0_ , \g72140/_0_ , \g72144/_1__syn_2 , \g72154/_1__syn_2 , \g72159/_0_ , \g72164/_1__syn_2 , \g72165/_1__syn_2 , \g72167/_1__syn_2 , \g72170/_1__syn_2 , \g72172/_1__syn_2 , \g72173/_0_ , \g72177/_1__syn_2 , \g72189/_0_ , \g72194/_0_ , \g72196/_0_ , \g72198/_0_ , \g72206/_1__syn_2 , \g72209/_1__syn_2 , \g72210/_1__syn_2 , \g72211/_0_ , \g72215/_0_ , \g72227/_1__syn_2 , \g72229/_1__syn_2 , \g72230/_0_ , \g72239/_0_ , \g72250/_3_ , \g72251/_3_ , \g72252/_3_ , \g72253/_3_ , \g72254/_3_ , \g72255/_3_ , \g72256/_3_ , \g72257/_3_ , \g72259/_3_ , \g72260/_3_ , \g72261/_3_ , \g72262/_3_ , \g72263/_3_ , \g72264/_3_ , \g72265/_3_ , \g72266/_3_ , \g72267/_3_ , \g72273/_3_ , \g72275/_3_ , \g72282/_3_ , \g72285/_3_ , \g72293/_3_ , \g72304/_3_ , \g72305/_3_ , \g72306/_3_ , \g72307/_3_ , \g72309/_3_ , \g72310/_3_ , \g72324/_3_ , \g72325/_3_ , \g72326/_3_ , \g72327/_3_ , \g72711/_0_ , \g72763/_0_ , \g72966/_0_ , \g72967/_0_ , \g73018/_0_ , \g73058/_0_ , \g73062/_0_ , \g73067/_0_ , \g73068/_0_ , \g73207/_0_ , \g75007/_1__syn_2 , \g75568/_1_ , \g75792/_0_ , \g75836/_0_ , \g76027/_0_ , \g76034/_0_ , \g76108/_0_ , \g76130/_0_ , \g76266/_0_ , \g76315/_0_ , \g76569/_0_ , \g76714/_0_ , \g77122/_1__syn_2 , \g77709/_1_ , \g81909/_0_ , \g81922/_0_ , \g81926/_1__syn_2 , \g82197/_1_ , \g82272/_0_ , \g82291/_0_ , \g82716/_0_ , \g82718/_0_ , \g82738/_0_ , \g82769/_0_ , \g82775/_0_ , \g82779/_1__syn_2 , \g82804/_0_ , \g82810/_0_ , \g82817/_0_ , \g82823/_0_ , \g82835/_0_ , \g82841/_0_ , \g82847/_0_ , \g82853/_0_ , \g82859/_0_ , \g82862/_1__syn_2 , \g82956/_0_ , \g82959/_1_ , \g83020/_0_ , \g83025/_0_ , \g83078/_0_ , \g83083/_0_ , \g83121/_0_ , \g83135/_0_ , \g83205/_0_ , \g83240/_0_ , \g83509/_1__syn_2 , \g83769/_0_ , \h0lock_pad , \h1sel_br[7]_pad , \h1sel_dma[0]_pad , \h1sel_dma[4]_pad , \h1sel_dma[7]_pad );
	input \ahb_mst0_hsizeo_reg[0]/NET0131  ;
	input \ahb_mst0_hsizeo_reg[1]/NET0131  ;
	input \ahb_mst0_hsizeo_reg[2]/NET0131  ;
	input \ahb_mst0_m0_m1_diff_tx_reg/NET0131  ;
	input \ahb_mst0_mx_cmd_st_reg[0]/NET0131  ;
	input \ahb_mst0_mx_cmd_st_reg[1]/NET0131  ;
	input \ahb_mst0_mx_dtp_reg/NET0131  ;
	input \ahb_mst1_mx_cmd_st_reg[0]/NET0131  ;
	input \ahb_mst1_mx_cmd_st_reg[1]/NET0131  ;
	input \ahb_mst1_mx_dtp_reg/NET0131  ;
	input \ahb_slv_br_st_reg[0]/NET0131  ;
	input \ahb_slv_br_st_reg[1]/NET0131  ;
	input \ahb_slv_br_st_reg[2]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[2]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[3]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[4]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[5]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[6]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[7]/NET0131  ;
	input \ahb_slv_slv_ad_d1o_reg[8]/NET0131  ;
	input \ahb_slv_slv_br_req_reg/NET0131  ;
	input \ahb_slv_slv_pt_d1o_reg[0]/NET0131  ;
	input \ahb_slv_slv_pt_d1o_reg[1]/NET0131  ;
	input \ahb_slv_slv_pt_d1o_reg[2]/NET0131  ;
	input \ahb_slv_slv_pt_d1o_reg[3]/NET0131  ;
	input \ahb_slv_slv_sz_d1o_reg[0]/NET0131  ;
	input \ahb_slv_slv_sz_d1o_reg[1]/NET0131  ;
	input \ahb_slv_slv_sz_d1o_reg[2]/NET0131  ;
	input \ahb_slv_slv_wr_d1o_reg/NET0131  ;
	input \ch_sel_arb_ch_sel_reg[0]/P0000_reg_syn_2  ;
	input \ch_sel_arb_ch_sel_reg[1]/P0000_reg_syn_2  ;
	input \ch_sel_arb_ch_sel_reg[2]/P0000_reg_syn_2  ;
	input \ch_sel_arb_chcsr_reg_reg[10]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[11]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[12]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[13]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[15]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[16]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[17]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[18]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[19]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[1]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[20]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[2]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[3]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[4]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[5]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[6]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[8]/NET0131  ;
	input \ch_sel_arb_chcsr_reg_reg[9]/NET0131  ;
	input \ch_sel_arb_req_reg/NET0131  ;
	input \ch_sel_de_stup_d1_reg/NET0131  ;
	input \ch_sel_dma_reqd1_reg[0]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[1]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[2]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[3]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[4]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[5]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[6]/NET0131  ;
	input \ch_sel_dma_reqd1_reg[7]/NET0131  ;
	input \ch_sel_dma_reqd2_reg[0]/NET0131  ;
	input \ch_sel_dma_reqd2_reg[1]/P0001  ;
	input \ch_sel_dma_reqd2_reg[2]/P0001  ;
	input \ch_sel_dma_reqd2_reg[3]/P0001  ;
	input \ch_sel_dma_reqd2_reg[4]/NET0131  ;
	input \ch_sel_dma_reqd2_reg[5]/NET0131  ;
	input \ch_sel_dma_reqd2_reg[6]/NET0131  ;
	input \ch_sel_dma_reqd2_reg[7]/NET0131  ;
	input \ch_sel_dma_rrarb0_state_reg[0]/NET0131  ;
	input \ch_sel_dma_rrarb0_state_reg[1]/NET0131  ;
	input \ch_sel_dma_rrarb0_state_reg[2]/NET0131  ;
	input \ch_sel_dma_rrarb1_state_reg[0]/NET0131  ;
	input \ch_sel_dma_rrarb1_state_reg[1]/NET0131  ;
	input \ch_sel_dma_rrarb1_state_reg[2]/NET0131  ;
	input \ch_sel_dma_rrarb2_state_reg[0]/NET0131  ;
	input \ch_sel_dma_rrarb2_state_reg[1]/NET0131  ;
	input \ch_sel_dma_rrarb2_state_reg[2]/NET0131  ;
	input \ch_sel_dma_rrarb3_state_reg[0]/NET0131  ;
	input \ch_sel_dma_rrarb3_state_reg[1]/NET0131  ;
	input \ch_sel_dma_rrarb3_state_reg[2]/NET0131  ;
	input \ch_sel_fix_pri_sel_reg[0]/NET0131  ;
	input \ch_sel_fix_pri_sel_reg[1]/NET0131  ;
	input \ch_sel_vld_req_any_d1_reg/NET0131  ;
	input \ctl_rf_abt_reg[0]/NET0131  ;
	input \ctl_rf_abt_reg[1]/NET0131  ;
	input \ctl_rf_abt_reg[2]/NET0131  ;
	input \ctl_rf_abt_reg[3]/NET0131  ;
	input \ctl_rf_abt_reg[4]/NET0131  ;
	input \ctl_rf_abt_reg[5]/NET0131  ;
	input \ctl_rf_abt_reg[6]/NET0131  ;
	input \ctl_rf_abt_reg[7]/NET0131  ;
	input \ctl_rf_be_d1_reg[0]/P0001  ;
	input \ctl_rf_be_d1_reg[1]/P0001  ;
	input \ctl_rf_be_d1_reg[2]/P0001  ;
	input \ctl_rf_be_d1_reg[3]/P0001  ;
	input \ctl_rf_c0_rf_autold_reg/NET0131  ;
	input \ctl_rf_c0_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c0_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[10]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[11]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[12]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[13]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[14]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[15]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c0_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c0_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c0_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c0_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c0_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c0_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c0_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[10]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[11]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[12]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[13]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[14]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[15]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c0_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c0_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c0_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c0_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c0_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c0_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c0_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c0_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c0_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c0_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c0_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c0_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c0_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c0_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c0_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c0_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c0_rf_mode_reg/NET0131  ;
	input \ctl_rf_c0_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c0_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c0_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c0_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c0_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c0_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c0_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c0_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c0_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c0_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c0brbs_reg[16]/NET0131  ;
	input \ctl_rf_c0brbs_reg[17]/NET0131  ;
	input \ctl_rf_c0brbs_reg[18]/NET0131  ;
	input \ctl_rf_c0brbs_reg[19]/NET0131  ;
	input \ctl_rf_c0brbs_reg[20]/NET0131  ;
	input \ctl_rf_c0brbs_reg[21]/NET0131  ;
	input \ctl_rf_c0brbs_reg[22]/NET0131  ;
	input \ctl_rf_c0brbs_reg[23]/NET0131  ;
	input \ctl_rf_c0brbs_reg[24]/NET0131  ;
	input \ctl_rf_c0brbs_reg[25]/NET0131  ;
	input \ctl_rf_c0brbs_reg[26]/NET0131  ;
	input \ctl_rf_c0brbs_reg[27]/NET0131  ;
	input \ctl_rf_c0brbs_reg[28]/NET0131  ;
	input \ctl_rf_c0brbs_reg[29]/NET0131  ;
	input \ctl_rf_c0brbs_reg[30]/NET0131  ;
	input \ctl_rf_c0brbs_reg[31]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c0dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c1_rf_autold_reg/NET0131  ;
	input \ctl_rf_c1_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c1_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[10]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[11]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[12]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[13]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[14]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[15]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c1_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c1_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c1_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c1_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c1_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c1_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c1_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[10]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[11]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[12]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[13]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[14]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[15]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c1_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c1_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c1_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c1_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c1_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c1_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c1_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c1_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c1_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c1_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c1_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c1_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c1_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c1_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c1_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c1_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c1_rf_mode_reg/NET0131  ;
	input \ctl_rf_c1_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c1_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c1_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c1_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c1_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c1_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c1_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c1_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c1_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c1_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c1brbs_reg[16]/NET0131  ;
	input \ctl_rf_c1brbs_reg[17]/NET0131  ;
	input \ctl_rf_c1brbs_reg[18]/NET0131  ;
	input \ctl_rf_c1brbs_reg[19]/NET0131  ;
	input \ctl_rf_c1brbs_reg[20]/NET0131  ;
	input \ctl_rf_c1brbs_reg[21]/NET0131  ;
	input \ctl_rf_c1brbs_reg[22]/NET0131  ;
	input \ctl_rf_c1brbs_reg[23]/NET0131  ;
	input \ctl_rf_c1brbs_reg[24]/NET0131  ;
	input \ctl_rf_c1brbs_reg[25]/NET0131  ;
	input \ctl_rf_c1brbs_reg[26]/NET0131  ;
	input \ctl_rf_c1brbs_reg[27]/NET0131  ;
	input \ctl_rf_c1brbs_reg[28]/NET0131  ;
	input \ctl_rf_c1brbs_reg[29]/NET0131  ;
	input \ctl_rf_c1brbs_reg[30]/NET0131  ;
	input \ctl_rf_c1brbs_reg[31]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c1dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c2_rf_autold_reg/NET0131  ;
	input \ctl_rf_c2_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c2_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[10]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[11]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[12]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[13]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[14]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[15]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c2_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c2_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c2_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c2_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c2_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c2_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c2_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[10]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[11]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[12]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[13]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[14]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[15]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c2_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c2_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c2_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c2_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c2_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c2_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c2_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c2_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c2_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c2_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c2_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c2_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c2_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c2_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c2_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c2_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c2_rf_mode_reg/NET0131  ;
	input \ctl_rf_c2_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c2_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c2_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c2_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c2_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c2_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c2_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c2_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c2_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c2_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c2brbs_reg[16]/NET0131  ;
	input \ctl_rf_c2brbs_reg[17]/NET0131  ;
	input \ctl_rf_c2brbs_reg[18]/NET0131  ;
	input \ctl_rf_c2brbs_reg[19]/NET0131  ;
	input \ctl_rf_c2brbs_reg[20]/NET0131  ;
	input \ctl_rf_c2brbs_reg[21]/NET0131  ;
	input \ctl_rf_c2brbs_reg[22]/NET0131  ;
	input \ctl_rf_c2brbs_reg[23]/NET0131  ;
	input \ctl_rf_c2brbs_reg[24]/NET0131  ;
	input \ctl_rf_c2brbs_reg[25]/NET0131  ;
	input \ctl_rf_c2brbs_reg[26]/NET0131  ;
	input \ctl_rf_c2brbs_reg[27]/NET0131  ;
	input \ctl_rf_c2brbs_reg[28]/NET0131  ;
	input \ctl_rf_c2brbs_reg[29]/NET0131  ;
	input \ctl_rf_c2brbs_reg[30]/NET0131  ;
	input \ctl_rf_c2brbs_reg[31]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c2dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c3_rf_autold_reg/NET0131  ;
	input \ctl_rf_c3_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c3_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[10]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[11]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[12]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[13]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[14]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[15]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c3_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c3_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c3_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c3_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c3_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c3_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c3_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[10]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[11]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[12]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[13]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[14]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[15]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c3_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c3_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c3_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c3_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c3_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c3_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c3_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c3_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c3_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c3_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c3_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c3_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c3_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c3_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c3_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c3_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c3_rf_mode_reg/NET0131  ;
	input \ctl_rf_c3_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c3_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c3_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c3_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c3_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c3_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c3_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c3_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c3_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c3_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c3brbs_reg[16]/NET0131  ;
	input \ctl_rf_c3brbs_reg[17]/NET0131  ;
	input \ctl_rf_c3brbs_reg[18]/NET0131  ;
	input \ctl_rf_c3brbs_reg[19]/NET0131  ;
	input \ctl_rf_c3brbs_reg[20]/NET0131  ;
	input \ctl_rf_c3brbs_reg[21]/NET0131  ;
	input \ctl_rf_c3brbs_reg[22]/NET0131  ;
	input \ctl_rf_c3brbs_reg[23]/NET0131  ;
	input \ctl_rf_c3brbs_reg[24]/NET0131  ;
	input \ctl_rf_c3brbs_reg[25]/NET0131  ;
	input \ctl_rf_c3brbs_reg[26]/NET0131  ;
	input \ctl_rf_c3brbs_reg[27]/NET0131  ;
	input \ctl_rf_c3brbs_reg[28]/NET0131  ;
	input \ctl_rf_c3brbs_reg[29]/NET0131  ;
	input \ctl_rf_c3brbs_reg[30]/NET0131  ;
	input \ctl_rf_c3brbs_reg[31]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c3dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c4_rf_autold_reg/NET0131  ;
	input \ctl_rf_c4_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c4_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[10]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[11]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[12]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[13]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[14]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[15]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c4_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c4_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c4_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c4_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c4_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c4_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c4_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[10]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[11]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[12]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[13]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[14]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[15]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c4_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c4_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c4_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c4_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c4_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c4_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c4_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c4_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c4_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c4_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c4_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c4_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c4_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c4_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c4_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c4_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c4_rf_mode_reg/NET0131  ;
	input \ctl_rf_c4_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c4_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c4_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c4_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c4_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c4_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c4_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c4_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c4_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c4_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c4brbs_reg[16]/NET0131  ;
	input \ctl_rf_c4brbs_reg[17]/NET0131  ;
	input \ctl_rf_c4brbs_reg[18]/NET0131  ;
	input \ctl_rf_c4brbs_reg[19]/NET0131  ;
	input \ctl_rf_c4brbs_reg[20]/NET0131  ;
	input \ctl_rf_c4brbs_reg[21]/NET0131  ;
	input \ctl_rf_c4brbs_reg[22]/NET0131  ;
	input \ctl_rf_c4brbs_reg[23]/NET0131  ;
	input \ctl_rf_c4brbs_reg[24]/NET0131  ;
	input \ctl_rf_c4brbs_reg[25]/NET0131  ;
	input \ctl_rf_c4brbs_reg[26]/NET0131  ;
	input \ctl_rf_c4brbs_reg[27]/NET0131  ;
	input \ctl_rf_c4brbs_reg[28]/NET0131  ;
	input \ctl_rf_c4brbs_reg[29]/NET0131  ;
	input \ctl_rf_c4brbs_reg[30]/NET0131  ;
	input \ctl_rf_c4brbs_reg[31]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c4dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c5_rf_autold_reg/NET0131  ;
	input \ctl_rf_c5_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c5_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[10]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[11]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[12]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[13]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[14]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[15]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c5_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c5_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c5_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c5_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c5_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c5_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c5_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[10]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[11]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[12]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[13]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[14]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[15]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c5_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c5_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c5_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c5_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c5_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c5_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c5_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c5_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c5_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c5_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c5_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c5_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c5_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c5_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c5_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c5_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c5_rf_mode_reg/NET0131  ;
	input \ctl_rf_c5_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c5_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c5_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c5_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c5_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c5_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c5_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c5_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c5_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c5_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c5brbs_reg[16]/NET0131  ;
	input \ctl_rf_c5brbs_reg[17]/NET0131  ;
	input \ctl_rf_c5brbs_reg[18]/NET0131  ;
	input \ctl_rf_c5brbs_reg[19]/NET0131  ;
	input \ctl_rf_c5brbs_reg[20]/NET0131  ;
	input \ctl_rf_c5brbs_reg[21]/NET0131  ;
	input \ctl_rf_c5brbs_reg[22]/NET0131  ;
	input \ctl_rf_c5brbs_reg[23]/NET0131  ;
	input \ctl_rf_c5brbs_reg[24]/NET0131  ;
	input \ctl_rf_c5brbs_reg[25]/NET0131  ;
	input \ctl_rf_c5brbs_reg[26]/NET0131  ;
	input \ctl_rf_c5brbs_reg[27]/NET0131  ;
	input \ctl_rf_c5brbs_reg[28]/NET0131  ;
	input \ctl_rf_c5brbs_reg[29]/NET0131  ;
	input \ctl_rf_c5brbs_reg[30]/NET0131  ;
	input \ctl_rf_c5brbs_reg[31]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c5dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c6_rf_autold_reg/NET0131  ;
	input \ctl_rf_c6_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c6_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[10]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[11]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[12]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[13]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[14]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[15]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c6_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c6_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c6_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c6_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c6_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c6_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c6_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[10]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[11]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[12]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[13]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[14]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[15]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c6_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c6_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c6_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c6_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c6_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c6_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c6_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c6_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c6_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c6_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c6_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c6_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c6_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c6_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c6_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c6_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c6_rf_mode_reg/NET0131  ;
	input \ctl_rf_c6_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c6_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c6_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c6_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c6_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c6_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c6_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c6_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c6_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c6_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c6brbs_reg[16]/NET0131  ;
	input \ctl_rf_c6brbs_reg[17]/NET0131  ;
	input \ctl_rf_c6brbs_reg[18]/NET0131  ;
	input \ctl_rf_c6brbs_reg[19]/NET0131  ;
	input \ctl_rf_c6brbs_reg[20]/NET0131  ;
	input \ctl_rf_c6brbs_reg[21]/NET0131  ;
	input \ctl_rf_c6brbs_reg[22]/NET0131  ;
	input \ctl_rf_c6brbs_reg[23]/NET0131  ;
	input \ctl_rf_c6brbs_reg[24]/NET0131  ;
	input \ctl_rf_c6brbs_reg[25]/NET0131  ;
	input \ctl_rf_c6brbs_reg[26]/NET0131  ;
	input \ctl_rf_c6brbs_reg[27]/NET0131  ;
	input \ctl_rf_c6brbs_reg[28]/NET0131  ;
	input \ctl_rf_c6brbs_reg[29]/NET0131  ;
	input \ctl_rf_c6brbs_reg[30]/NET0131  ;
	input \ctl_rf_c6brbs_reg[31]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c6dmabs_reg[31]/NET0131  ;
	input \ctl_rf_c7_rf_autold_reg/NET0131  ;
	input \ctl_rf_c7_rf_ch_en_reg/NET0131  ;
	input \ctl_rf_c7_rf_chabt_reg/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[10]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[11]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[12]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[13]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[14]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[15]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[16]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[17]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[18]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[19]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[20]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[21]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[22]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[23]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[24]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[25]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[26]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[27]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[28]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[29]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[30]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[31]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[3]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[4]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[5]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[6]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[7]/P0002  ;
	input \ctl_rf_c7_rf_chdad_reg[8]/NET0131  ;
	input \ctl_rf_c7_rf_chdad_reg[9]/P0002  ;
	input \ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_on_reg/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[0]/P0002  ;
	input \ctl_rf_c7_rf_chllp_reg[10]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[11]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[12]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[13]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[14]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[15]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[16]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[17]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[18]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[19]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[1]/P0002  ;
	input \ctl_rf_c7_rf_chllp_reg[20]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[21]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[22]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[23]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[24]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[25]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[26]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[27]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[28]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[29]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[30]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[31]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[3]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[4]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[5]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[6]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[7]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[8]/NET0131  ;
	input \ctl_rf_c7_rf_chllp_reg[9]/NET0131  ;
	input \ctl_rf_c7_rf_chllpen_reg/NET0131  ;
	input \ctl_rf_c7_rf_chpri_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_chpri_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[10]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[11]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[12]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[13]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[14]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[15]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[16]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[17]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[18]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[19]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[20]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[21]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[22]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[23]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[24]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[25]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[26]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[27]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[28]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[29]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[30]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[31]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[3]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[4]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[5]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[6]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[7]/NET0131  ;
	input \ctl_rf_c7_rf_chsad_reg[8]/P0002  ;
	input \ctl_rf_c7_rf_chsad_reg[9]/NET0131  ;
	input \ctl_rf_c7_rf_chtsz_reg[0]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[10]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[11]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[1]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[2]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[3]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[4]/NET0131  ;
	input \ctl_rf_c7_rf_chtsz_reg[5]/NET0131  ;
	input \ctl_rf_c7_rf_chtsz_reg[6]/NET0131  ;
	input \ctl_rf_c7_rf_chtsz_reg[7]/NET0131  ;
	input \ctl_rf_c7_rf_chtsz_reg[8]/P0002  ;
	input \ctl_rf_c7_rf_chtsz_reg[9]/P0002  ;
	input \ctl_rf_c7_rf_dad_ctl0_reg/NET0131  ;
	input \ctl_rf_c7_rf_dad_ctl1_reg/NET0131  ;
	input \ctl_rf_c7_rf_dreqmode_reg/NET0131  ;
	input \ctl_rf_c7_rf_dst_sel_reg/NET0131  ;
	input \ctl_rf_c7_rf_dwidth_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_dwidth_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_dwidth_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_int_abt_msk_reg/NET0131  ;
	input \ctl_rf_c7_rf_int_err_msk_reg/NET0131  ;
	input \ctl_rf_c7_rf_int_tc1_msk_reg/NET0131  ;
	input \ctl_rf_c7_rf_int_tc_msk_reg/NET0131  ;
	input \ctl_rf_c7_rf_mode_reg/NET0131  ;
	input \ctl_rf_c7_rf_prot1_reg/NET0131  ;
	input \ctl_rf_c7_rf_prot2_reg/NET0131  ;
	input \ctl_rf_c7_rf_prot3_reg/NET0131  ;
	input \ctl_rf_c7_rf_sad_ctl0_reg/NET0131  ;
	input \ctl_rf_c7_rf_sad_ctl1_reg/NET0131  ;
	input \ctl_rf_c7_rf_src_sel_reg/NET0131  ;
	input \ctl_rf_c7_rf_src_sz_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_src_sz_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_src_sz_reg[2]/NET0131  ;
	input \ctl_rf_c7_rf_swidth_reg[0]/NET0131  ;
	input \ctl_rf_c7_rf_swidth_reg[1]/NET0131  ;
	input \ctl_rf_c7_rf_swidth_reg[2]/NET0131  ;
	input \ctl_rf_c7brbs_reg[16]/NET0131  ;
	input \ctl_rf_c7brbs_reg[17]/NET0131  ;
	input \ctl_rf_c7brbs_reg[18]/NET0131  ;
	input \ctl_rf_c7brbs_reg[19]/NET0131  ;
	input \ctl_rf_c7brbs_reg[20]/NET0131  ;
	input \ctl_rf_c7brbs_reg[21]/NET0131  ;
	input \ctl_rf_c7brbs_reg[22]/NET0131  ;
	input \ctl_rf_c7brbs_reg[23]/NET0131  ;
	input \ctl_rf_c7brbs_reg[24]/NET0131  ;
	input \ctl_rf_c7brbs_reg[25]/NET0131  ;
	input \ctl_rf_c7brbs_reg[26]/NET0131  ;
	input \ctl_rf_c7brbs_reg[27]/NET0131  ;
	input \ctl_rf_c7brbs_reg[28]/NET0131  ;
	input \ctl_rf_c7brbs_reg[29]/NET0131  ;
	input \ctl_rf_c7brbs_reg[30]/NET0131  ;
	input \ctl_rf_c7brbs_reg[31]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[16]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[17]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[18]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[19]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[20]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[21]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[22]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[23]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[24]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[25]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[26]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[27]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[28]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[29]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[30]/NET0131  ;
	input \ctl_rf_c7dmabs_reg[31]/NET0131  ;
	input \ctl_rf_dmacen_reg/NET0131  ;
	input \ctl_rf_m0end_reg/NET0131  ;
	input \ctl_rf_m1end_reg/NET0131  ;
	input \ctl_rf_rf_sel_d1_reg/NET0131  ;
	input \ctl_rf_sync_reg[0]/NET0131  ;
	input \ctl_rf_sync_reg[1]/NET0131  ;
	input \ctl_rf_sync_reg[2]/NET0131  ;
	input \ctl_rf_sync_reg[3]/NET0131  ;
	input \ctl_rf_sync_reg[4]/NET0131  ;
	input \ctl_rf_sync_reg[5]/NET0131  ;
	input \ctl_rf_sync_reg[6]/NET0131  ;
	input \ctl_rf_sync_reg[7]/NET0131  ;
	input \ctl_rf_tc_reg[0]/NET0131  ;
	input \ctl_rf_tc_reg[1]/NET0131  ;
	input \ctl_rf_tc_reg[2]/NET0131  ;
	input \ctl_rf_tc_reg[3]/NET0131  ;
	input \ctl_rf_tc_reg[4]/NET0131  ;
	input \ctl_rf_tc_reg[5]/NET0131  ;
	input \ctl_rf_tc_reg[6]/NET0131  ;
	input \ctl_rf_tc_reg[7]/NET0131  ;
	input \de_bst_cnt_reg[0]/NET0131  ;
	input \de_bst_cnt_reg[2]/NET0131  ;
	input \de_bst_cnt_reg[3]/NET0131  ;
	input \de_bst_cnt_reg[4]/NET0131  ;
	input \de_bst_cnt_reg[5]/NET0131  ;
	input \de_bst_cnt_reg[6]/NET0131  ;
	input \de_bst_cnt_reg[7]/NET0131  ;
	input \de_bst_cnt_reg[8]/NET0131  ;
	input \de_de_st_reg[0]/NET0131  ;
	input \de_de_st_reg[1]/NET0131  ;
	input \de_de_st_reg[2]/NET0131  ;
	input \de_de_st_reg[5]/NET0131  ;
	input \de_de_st_reg[6]/NET0131  ;
	input \de_m0_arb_st_reg/NET0131  ;
	input \de_m0_is_llp_reg/NET0131  ;
	input \de_m1_arb_st_reg[0]/NET0131  ;
	input \de_m1_arb_st_reg[1]/NET0131  ;
	input \de_m1_is_llp_reg/NET0131  ;
	input \de_st_rd_msk_reg/NET0131  ;
	input \de_tsz_cnt_reg[0]/NET0131  ;
	input \de_tsz_cnt_reg[10]/NET0131  ;
	input \de_tsz_cnt_reg[11]/NET0131  ;
	input \de_tsz_cnt_reg[1]/NET0131  ;
	input \de_tsz_cnt_reg[2]/NET0131  ;
	input \de_tsz_cnt_reg[3]/NET0131  ;
	input \de_tsz_cnt_reg[4]/NET0131  ;
	input \de_tsz_cnt_reg[5]/NET0131  ;
	input \de_tsz_cnt_reg[6]/NET0131  ;
	input \de_tsz_cnt_reg[7]/NET0131  ;
	input \de_tsz_cnt_reg[8]/NET0131  ;
	input \de_tsz_cnt_reg[9]/NET0131  ;
	input \dma_ack[0]_pad  ;
	input \dma_ack[1]_pad  ;
	input \dma_ack[2]_pad  ;
	input \dma_ack[3]_pad  ;
	input \dma_ack[4]_pad  ;
	input \dma_ack[5]_pad  ;
	input \dma_ack[6]_pad  ;
	input \dma_ack[7]_pad  ;
	input \dma_tc[0]_pad  ;
	input \dma_tc[1]_pad  ;
	input \dma_tc[2]_pad  ;
	input \dma_tc[3]_pad  ;
	input \dma_tc[4]_pad  ;
	input \dma_tc[5]_pad  ;
	input \dma_tc[6]_pad  ;
	input \dma_tc[7]_pad  ;
	input \h0burst[0]_pad  ;
	input \h0grant_pad  ;
	input \h0readyin_pad  ;
	input \h0req_pad  ;
	input \h0resp[0]_pad  ;
	input \h0resp[1]_pad  ;
	input \h0write_pad  ;
	input \h1burst[0]_pad  ;
	input \h1prot[0]_pad  ;
	input \h1rdt0_br[0]_pad  ;
	input \h1rdt0_br[10]_pad  ;
	input \h1rdt0_br[11]_pad  ;
	input \h1rdt0_br[12]_pad  ;
	input \h1rdt0_br[13]_pad  ;
	input \h1rdt0_br[14]_pad  ;
	input \h1rdt0_br[15]_pad  ;
	input \h1rdt0_br[16]_pad  ;
	input \h1rdt0_br[17]_pad  ;
	input \h1rdt0_br[18]_pad  ;
	input \h1rdt0_br[19]_pad  ;
	input \h1rdt0_br[1]_pad  ;
	input \h1rdt0_br[20]_pad  ;
	input \h1rdt0_br[21]_pad  ;
	input \h1rdt0_br[22]_pad  ;
	input \h1rdt0_br[23]_pad  ;
	input \h1rdt0_br[24]_pad  ;
	input \h1rdt0_br[25]_pad  ;
	input \h1rdt0_br[26]_pad  ;
	input \h1rdt0_br[27]_pad  ;
	input \h1rdt0_br[28]_pad  ;
	input \h1rdt0_br[29]_pad  ;
	input \h1rdt0_br[2]_pad  ;
	input \h1rdt0_br[30]_pad  ;
	input \h1rdt0_br[31]_pad  ;
	input \h1rdt0_br[3]_pad  ;
	input \h1rdt0_br[4]_pad  ;
	input \h1rdt0_br[5]_pad  ;
	input \h1rdt0_br[6]_pad  ;
	input \h1rdt0_br[7]_pad  ;
	input \h1rdt0_br[8]_pad  ;
	input \h1rdt0_br[9]_pad  ;
	input \h1rdt0_dma[0]_pad  ;
	input \h1rdt0_dma[10]_pad  ;
	input \h1rdt0_dma[11]_pad  ;
	input \h1rdt0_dma[12]_pad  ;
	input \h1rdt0_dma[13]_pad  ;
	input \h1rdt0_dma[14]_pad  ;
	input \h1rdt0_dma[15]_pad  ;
	input \h1rdt0_dma[16]_pad  ;
	input \h1rdt0_dma[17]_pad  ;
	input \h1rdt0_dma[18]_pad  ;
	input \h1rdt0_dma[19]_pad  ;
	input \h1rdt0_dma[1]_pad  ;
	input \h1rdt0_dma[20]_pad  ;
	input \h1rdt0_dma[21]_pad  ;
	input \h1rdt0_dma[22]_pad  ;
	input \h1rdt0_dma[23]_pad  ;
	input \h1rdt0_dma[24]_pad  ;
	input \h1rdt0_dma[25]_pad  ;
	input \h1rdt0_dma[26]_pad  ;
	input \h1rdt0_dma[27]_pad  ;
	input \h1rdt0_dma[28]_pad  ;
	input \h1rdt0_dma[29]_pad  ;
	input \h1rdt0_dma[2]_pad  ;
	input \h1rdt0_dma[30]_pad  ;
	input \h1rdt0_dma[31]_pad  ;
	input \h1rdt0_dma[3]_pad  ;
	input \h1rdt0_dma[4]_pad  ;
	input \h1rdt0_dma[5]_pad  ;
	input \h1rdt0_dma[6]_pad  ;
	input \h1rdt0_dma[7]_pad  ;
	input \h1rdt0_dma[8]_pad  ;
	input \h1rdt0_dma[9]_pad  ;
	input \h1rdt1_br[0]_pad  ;
	input \h1rdt1_br[10]_pad  ;
	input \h1rdt1_br[11]_pad  ;
	input \h1rdt1_br[12]_pad  ;
	input \h1rdt1_br[13]_pad  ;
	input \h1rdt1_br[14]_pad  ;
	input \h1rdt1_br[15]_pad  ;
	input \h1rdt1_br[16]_pad  ;
	input \h1rdt1_br[17]_pad  ;
	input \h1rdt1_br[18]_pad  ;
	input \h1rdt1_br[19]_pad  ;
	input \h1rdt1_br[1]_pad  ;
	input \h1rdt1_br[20]_pad  ;
	input \h1rdt1_br[21]_pad  ;
	input \h1rdt1_br[22]_pad  ;
	input \h1rdt1_br[23]_pad  ;
	input \h1rdt1_br[24]_pad  ;
	input \h1rdt1_br[25]_pad  ;
	input \h1rdt1_br[26]_pad  ;
	input \h1rdt1_br[27]_pad  ;
	input \h1rdt1_br[28]_pad  ;
	input \h1rdt1_br[29]_pad  ;
	input \h1rdt1_br[2]_pad  ;
	input \h1rdt1_br[30]_pad  ;
	input \h1rdt1_br[31]_pad  ;
	input \h1rdt1_br[3]_pad  ;
	input \h1rdt1_br[4]_pad  ;
	input \h1rdt1_br[5]_pad  ;
	input \h1rdt1_br[6]_pad  ;
	input \h1rdt1_br[7]_pad  ;
	input \h1rdt1_br[8]_pad  ;
	input \h1rdt1_br[9]_pad  ;
	input \h1rdt1_dma[0]_pad  ;
	input \h1rdt1_dma[10]_pad  ;
	input \h1rdt1_dma[11]_pad  ;
	input \h1rdt1_dma[12]_pad  ;
	input \h1rdt1_dma[13]_pad  ;
	input \h1rdt1_dma[14]_pad  ;
	input \h1rdt1_dma[15]_pad  ;
	input \h1rdt1_dma[16]_pad  ;
	input \h1rdt1_dma[17]_pad  ;
	input \h1rdt1_dma[18]_pad  ;
	input \h1rdt1_dma[19]_pad  ;
	input \h1rdt1_dma[1]_pad  ;
	input \h1rdt1_dma[20]_pad  ;
	input \h1rdt1_dma[21]_pad  ;
	input \h1rdt1_dma[22]_pad  ;
	input \h1rdt1_dma[23]_pad  ;
	input \h1rdt1_dma[24]_pad  ;
	input \h1rdt1_dma[25]_pad  ;
	input \h1rdt1_dma[26]_pad  ;
	input \h1rdt1_dma[27]_pad  ;
	input \h1rdt1_dma[28]_pad  ;
	input \h1rdt1_dma[29]_pad  ;
	input \h1rdt1_dma[2]_pad  ;
	input \h1rdt1_dma[30]_pad  ;
	input \h1rdt1_dma[31]_pad  ;
	input \h1rdt1_dma[3]_pad  ;
	input \h1rdt1_dma[4]_pad  ;
	input \h1rdt1_dma[5]_pad  ;
	input \h1rdt1_dma[6]_pad  ;
	input \h1rdt1_dma[7]_pad  ;
	input \h1rdt1_dma[8]_pad  ;
	input \h1rdt1_dma[9]_pad  ;
	input \h1rdt2_br[0]_pad  ;
	input \h1rdt2_br[10]_pad  ;
	input \h1rdt2_br[11]_pad  ;
	input \h1rdt2_br[12]_pad  ;
	input \h1rdt2_br[13]_pad  ;
	input \h1rdt2_br[14]_pad  ;
	input \h1rdt2_br[15]_pad  ;
	input \h1rdt2_br[16]_pad  ;
	input \h1rdt2_br[17]_pad  ;
	input \h1rdt2_br[18]_pad  ;
	input \h1rdt2_br[19]_pad  ;
	input \h1rdt2_br[1]_pad  ;
	input \h1rdt2_br[20]_pad  ;
	input \h1rdt2_br[21]_pad  ;
	input \h1rdt2_br[22]_pad  ;
	input \h1rdt2_br[23]_pad  ;
	input \h1rdt2_br[24]_pad  ;
	input \h1rdt2_br[25]_pad  ;
	input \h1rdt2_br[26]_pad  ;
	input \h1rdt2_br[27]_pad  ;
	input \h1rdt2_br[28]_pad  ;
	input \h1rdt2_br[29]_pad  ;
	input \h1rdt2_br[2]_pad  ;
	input \h1rdt2_br[30]_pad  ;
	input \h1rdt2_br[31]_pad  ;
	input \h1rdt2_br[3]_pad  ;
	input \h1rdt2_br[4]_pad  ;
	input \h1rdt2_br[5]_pad  ;
	input \h1rdt2_br[6]_pad  ;
	input \h1rdt2_br[7]_pad  ;
	input \h1rdt2_br[8]_pad  ;
	input \h1rdt2_br[9]_pad  ;
	input \h1rdt2_dma[0]_pad  ;
	input \h1rdt2_dma[10]_pad  ;
	input \h1rdt2_dma[11]_pad  ;
	input \h1rdt2_dma[12]_pad  ;
	input \h1rdt2_dma[13]_pad  ;
	input \h1rdt2_dma[14]_pad  ;
	input \h1rdt2_dma[15]_pad  ;
	input \h1rdt2_dma[16]_pad  ;
	input \h1rdt2_dma[17]_pad  ;
	input \h1rdt2_dma[18]_pad  ;
	input \h1rdt2_dma[19]_pad  ;
	input \h1rdt2_dma[1]_pad  ;
	input \h1rdt2_dma[20]_pad  ;
	input \h1rdt2_dma[21]_pad  ;
	input \h1rdt2_dma[22]_pad  ;
	input \h1rdt2_dma[23]_pad  ;
	input \h1rdt2_dma[24]_pad  ;
	input \h1rdt2_dma[25]_pad  ;
	input \h1rdt2_dma[26]_pad  ;
	input \h1rdt2_dma[27]_pad  ;
	input \h1rdt2_dma[28]_pad  ;
	input \h1rdt2_dma[29]_pad  ;
	input \h1rdt2_dma[2]_pad  ;
	input \h1rdt2_dma[30]_pad  ;
	input \h1rdt2_dma[31]_pad  ;
	input \h1rdt2_dma[3]_pad  ;
	input \h1rdt2_dma[4]_pad  ;
	input \h1rdt2_dma[5]_pad  ;
	input \h1rdt2_dma[6]_pad  ;
	input \h1rdt2_dma[7]_pad  ;
	input \h1rdt2_dma[8]_pad  ;
	input \h1rdt2_dma[9]_pad  ;
	input \h1rdt3_br[0]_pad  ;
	input \h1rdt3_br[10]_pad  ;
	input \h1rdt3_br[11]_pad  ;
	input \h1rdt3_br[12]_pad  ;
	input \h1rdt3_br[13]_pad  ;
	input \h1rdt3_br[14]_pad  ;
	input \h1rdt3_br[15]_pad  ;
	input \h1rdt3_br[16]_pad  ;
	input \h1rdt3_br[17]_pad  ;
	input \h1rdt3_br[18]_pad  ;
	input \h1rdt3_br[19]_pad  ;
	input \h1rdt3_br[1]_pad  ;
	input \h1rdt3_br[20]_pad  ;
	input \h1rdt3_br[21]_pad  ;
	input \h1rdt3_br[22]_pad  ;
	input \h1rdt3_br[23]_pad  ;
	input \h1rdt3_br[24]_pad  ;
	input \h1rdt3_br[25]_pad  ;
	input \h1rdt3_br[26]_pad  ;
	input \h1rdt3_br[27]_pad  ;
	input \h1rdt3_br[28]_pad  ;
	input \h1rdt3_br[29]_pad  ;
	input \h1rdt3_br[2]_pad  ;
	input \h1rdt3_br[30]_pad  ;
	input \h1rdt3_br[31]_pad  ;
	input \h1rdt3_br[3]_pad  ;
	input \h1rdt3_br[4]_pad  ;
	input \h1rdt3_br[5]_pad  ;
	input \h1rdt3_br[6]_pad  ;
	input \h1rdt3_br[7]_pad  ;
	input \h1rdt3_br[8]_pad  ;
	input \h1rdt3_br[9]_pad  ;
	input \h1rdt3_dma[0]_pad  ;
	input \h1rdt3_dma[10]_pad  ;
	input \h1rdt3_dma[11]_pad  ;
	input \h1rdt3_dma[12]_pad  ;
	input \h1rdt3_dma[13]_pad  ;
	input \h1rdt3_dma[14]_pad  ;
	input \h1rdt3_dma[15]_pad  ;
	input \h1rdt3_dma[16]_pad  ;
	input \h1rdt3_dma[17]_pad  ;
	input \h1rdt3_dma[18]_pad  ;
	input \h1rdt3_dma[19]_pad  ;
	input \h1rdt3_dma[1]_pad  ;
	input \h1rdt3_dma[20]_pad  ;
	input \h1rdt3_dma[21]_pad  ;
	input \h1rdt3_dma[22]_pad  ;
	input \h1rdt3_dma[23]_pad  ;
	input \h1rdt3_dma[24]_pad  ;
	input \h1rdt3_dma[25]_pad  ;
	input \h1rdt3_dma[26]_pad  ;
	input \h1rdt3_dma[27]_pad  ;
	input \h1rdt3_dma[28]_pad  ;
	input \h1rdt3_dma[29]_pad  ;
	input \h1rdt3_dma[2]_pad  ;
	input \h1rdt3_dma[30]_pad  ;
	input \h1rdt3_dma[31]_pad  ;
	input \h1rdt3_dma[3]_pad  ;
	input \h1rdt3_dma[4]_pad  ;
	input \h1rdt3_dma[5]_pad  ;
	input \h1rdt3_dma[6]_pad  ;
	input \h1rdt3_dma[7]_pad  ;
	input \h1rdt3_dma[8]_pad  ;
	input \h1rdt3_dma[9]_pad  ;
	input \h1rdt4_br[0]_pad  ;
	input \h1rdt4_br[10]_pad  ;
	input \h1rdt4_br[11]_pad  ;
	input \h1rdt4_br[12]_pad  ;
	input \h1rdt4_br[13]_pad  ;
	input \h1rdt4_br[14]_pad  ;
	input \h1rdt4_br[15]_pad  ;
	input \h1rdt4_br[16]_pad  ;
	input \h1rdt4_br[17]_pad  ;
	input \h1rdt4_br[18]_pad  ;
	input \h1rdt4_br[19]_pad  ;
	input \h1rdt4_br[1]_pad  ;
	input \h1rdt4_br[20]_pad  ;
	input \h1rdt4_br[21]_pad  ;
	input \h1rdt4_br[22]_pad  ;
	input \h1rdt4_br[23]_pad  ;
	input \h1rdt4_br[24]_pad  ;
	input \h1rdt4_br[25]_pad  ;
	input \h1rdt4_br[26]_pad  ;
	input \h1rdt4_br[27]_pad  ;
	input \h1rdt4_br[28]_pad  ;
	input \h1rdt4_br[29]_pad  ;
	input \h1rdt4_br[2]_pad  ;
	input \h1rdt4_br[30]_pad  ;
	input \h1rdt4_br[31]_pad  ;
	input \h1rdt4_br[3]_pad  ;
	input \h1rdt4_br[4]_pad  ;
	input \h1rdt4_br[5]_pad  ;
	input \h1rdt4_br[6]_pad  ;
	input \h1rdt4_br[7]_pad  ;
	input \h1rdt4_br[8]_pad  ;
	input \h1rdt4_br[9]_pad  ;
	input \h1rdt4_dma[0]_pad  ;
	input \h1rdt4_dma[10]_pad  ;
	input \h1rdt4_dma[11]_pad  ;
	input \h1rdt4_dma[12]_pad  ;
	input \h1rdt4_dma[13]_pad  ;
	input \h1rdt4_dma[14]_pad  ;
	input \h1rdt4_dma[15]_pad  ;
	input \h1rdt4_dma[16]_pad  ;
	input \h1rdt4_dma[17]_pad  ;
	input \h1rdt4_dma[18]_pad  ;
	input \h1rdt4_dma[19]_pad  ;
	input \h1rdt4_dma[1]_pad  ;
	input \h1rdt4_dma[20]_pad  ;
	input \h1rdt4_dma[21]_pad  ;
	input \h1rdt4_dma[22]_pad  ;
	input \h1rdt4_dma[23]_pad  ;
	input \h1rdt4_dma[24]_pad  ;
	input \h1rdt4_dma[25]_pad  ;
	input \h1rdt4_dma[26]_pad  ;
	input \h1rdt4_dma[27]_pad  ;
	input \h1rdt4_dma[28]_pad  ;
	input \h1rdt4_dma[29]_pad  ;
	input \h1rdt4_dma[2]_pad  ;
	input \h1rdt4_dma[30]_pad  ;
	input \h1rdt4_dma[31]_pad  ;
	input \h1rdt4_dma[3]_pad  ;
	input \h1rdt4_dma[4]_pad  ;
	input \h1rdt4_dma[5]_pad  ;
	input \h1rdt4_dma[6]_pad  ;
	input \h1rdt4_dma[7]_pad  ;
	input \h1rdt4_dma[8]_pad  ;
	input \h1rdt4_dma[9]_pad  ;
	input \h1rdt5_br[0]_pad  ;
	input \h1rdt5_br[10]_pad  ;
	input \h1rdt5_br[11]_pad  ;
	input \h1rdt5_br[12]_pad  ;
	input \h1rdt5_br[13]_pad  ;
	input \h1rdt5_br[14]_pad  ;
	input \h1rdt5_br[15]_pad  ;
	input \h1rdt5_br[16]_pad  ;
	input \h1rdt5_br[17]_pad  ;
	input \h1rdt5_br[18]_pad  ;
	input \h1rdt5_br[19]_pad  ;
	input \h1rdt5_br[1]_pad  ;
	input \h1rdt5_br[20]_pad  ;
	input \h1rdt5_br[21]_pad  ;
	input \h1rdt5_br[22]_pad  ;
	input \h1rdt5_br[23]_pad  ;
	input \h1rdt5_br[24]_pad  ;
	input \h1rdt5_br[25]_pad  ;
	input \h1rdt5_br[26]_pad  ;
	input \h1rdt5_br[27]_pad  ;
	input \h1rdt5_br[28]_pad  ;
	input \h1rdt5_br[29]_pad  ;
	input \h1rdt5_br[2]_pad  ;
	input \h1rdt5_br[30]_pad  ;
	input \h1rdt5_br[31]_pad  ;
	input \h1rdt5_br[3]_pad  ;
	input \h1rdt5_br[4]_pad  ;
	input \h1rdt5_br[5]_pad  ;
	input \h1rdt5_br[6]_pad  ;
	input \h1rdt5_br[7]_pad  ;
	input \h1rdt5_br[8]_pad  ;
	input \h1rdt5_br[9]_pad  ;
	input \h1rdt5_dma[0]_pad  ;
	input \h1rdt5_dma[10]_pad  ;
	input \h1rdt5_dma[11]_pad  ;
	input \h1rdt5_dma[12]_pad  ;
	input \h1rdt5_dma[13]_pad  ;
	input \h1rdt5_dma[14]_pad  ;
	input \h1rdt5_dma[15]_pad  ;
	input \h1rdt5_dma[16]_pad  ;
	input \h1rdt5_dma[17]_pad  ;
	input \h1rdt5_dma[18]_pad  ;
	input \h1rdt5_dma[19]_pad  ;
	input \h1rdt5_dma[1]_pad  ;
	input \h1rdt5_dma[20]_pad  ;
	input \h1rdt5_dma[21]_pad  ;
	input \h1rdt5_dma[22]_pad  ;
	input \h1rdt5_dma[23]_pad  ;
	input \h1rdt5_dma[24]_pad  ;
	input \h1rdt5_dma[25]_pad  ;
	input \h1rdt5_dma[26]_pad  ;
	input \h1rdt5_dma[27]_pad  ;
	input \h1rdt5_dma[28]_pad  ;
	input \h1rdt5_dma[29]_pad  ;
	input \h1rdt5_dma[2]_pad  ;
	input \h1rdt5_dma[30]_pad  ;
	input \h1rdt5_dma[31]_pad  ;
	input \h1rdt5_dma[3]_pad  ;
	input \h1rdt5_dma[4]_pad  ;
	input \h1rdt5_dma[5]_pad  ;
	input \h1rdt5_dma[6]_pad  ;
	input \h1rdt5_dma[7]_pad  ;
	input \h1rdt5_dma[8]_pad  ;
	input \h1rdt5_dma[9]_pad  ;
	input \h1rdt6_br[0]_pad  ;
	input \h1rdt6_br[10]_pad  ;
	input \h1rdt6_br[11]_pad  ;
	input \h1rdt6_br[12]_pad  ;
	input \h1rdt6_br[13]_pad  ;
	input \h1rdt6_br[14]_pad  ;
	input \h1rdt6_br[15]_pad  ;
	input \h1rdt6_br[16]_pad  ;
	input \h1rdt6_br[17]_pad  ;
	input \h1rdt6_br[18]_pad  ;
	input \h1rdt6_br[19]_pad  ;
	input \h1rdt6_br[1]_pad  ;
	input \h1rdt6_br[20]_pad  ;
	input \h1rdt6_br[21]_pad  ;
	input \h1rdt6_br[22]_pad  ;
	input \h1rdt6_br[23]_pad  ;
	input \h1rdt6_br[24]_pad  ;
	input \h1rdt6_br[25]_pad  ;
	input \h1rdt6_br[26]_pad  ;
	input \h1rdt6_br[27]_pad  ;
	input \h1rdt6_br[28]_pad  ;
	input \h1rdt6_br[29]_pad  ;
	input \h1rdt6_br[2]_pad  ;
	input \h1rdt6_br[30]_pad  ;
	input \h1rdt6_br[31]_pad  ;
	input \h1rdt6_br[3]_pad  ;
	input \h1rdt6_br[4]_pad  ;
	input \h1rdt6_br[5]_pad  ;
	input \h1rdt6_br[6]_pad  ;
	input \h1rdt6_br[7]_pad  ;
	input \h1rdt6_br[8]_pad  ;
	input \h1rdt6_br[9]_pad  ;
	input \h1rdt6_dma[0]_pad  ;
	input \h1rdt6_dma[10]_pad  ;
	input \h1rdt6_dma[11]_pad  ;
	input \h1rdt6_dma[12]_pad  ;
	input \h1rdt6_dma[13]_pad  ;
	input \h1rdt6_dma[14]_pad  ;
	input \h1rdt6_dma[15]_pad  ;
	input \h1rdt6_dma[16]_pad  ;
	input \h1rdt6_dma[17]_pad  ;
	input \h1rdt6_dma[18]_pad  ;
	input \h1rdt6_dma[19]_pad  ;
	input \h1rdt6_dma[1]_pad  ;
	input \h1rdt6_dma[20]_pad  ;
	input \h1rdt6_dma[21]_pad  ;
	input \h1rdt6_dma[22]_pad  ;
	input \h1rdt6_dma[23]_pad  ;
	input \h1rdt6_dma[24]_pad  ;
	input \h1rdt6_dma[25]_pad  ;
	input \h1rdt6_dma[26]_pad  ;
	input \h1rdt6_dma[27]_pad  ;
	input \h1rdt6_dma[28]_pad  ;
	input \h1rdt6_dma[29]_pad  ;
	input \h1rdt6_dma[2]_pad  ;
	input \h1rdt6_dma[30]_pad  ;
	input \h1rdt6_dma[31]_pad  ;
	input \h1rdt6_dma[3]_pad  ;
	input \h1rdt6_dma[4]_pad  ;
	input \h1rdt6_dma[5]_pad  ;
	input \h1rdt6_dma[6]_pad  ;
	input \h1rdt6_dma[7]_pad  ;
	input \h1rdt6_dma[8]_pad  ;
	input \h1rdt6_dma[9]_pad  ;
	input \h1rdt7_br[0]_pad  ;
	input \h1rdt7_br[10]_pad  ;
	input \h1rdt7_br[11]_pad  ;
	input \h1rdt7_br[12]_pad  ;
	input \h1rdt7_br[13]_pad  ;
	input \h1rdt7_br[14]_pad  ;
	input \h1rdt7_br[15]_pad  ;
	input \h1rdt7_br[16]_pad  ;
	input \h1rdt7_br[17]_pad  ;
	input \h1rdt7_br[18]_pad  ;
	input \h1rdt7_br[19]_pad  ;
	input \h1rdt7_br[1]_pad  ;
	input \h1rdt7_br[20]_pad  ;
	input \h1rdt7_br[21]_pad  ;
	input \h1rdt7_br[22]_pad  ;
	input \h1rdt7_br[23]_pad  ;
	input \h1rdt7_br[24]_pad  ;
	input \h1rdt7_br[25]_pad  ;
	input \h1rdt7_br[26]_pad  ;
	input \h1rdt7_br[27]_pad  ;
	input \h1rdt7_br[28]_pad  ;
	input \h1rdt7_br[29]_pad  ;
	input \h1rdt7_br[2]_pad  ;
	input \h1rdt7_br[30]_pad  ;
	input \h1rdt7_br[31]_pad  ;
	input \h1rdt7_br[3]_pad  ;
	input \h1rdt7_br[4]_pad  ;
	input \h1rdt7_br[5]_pad  ;
	input \h1rdt7_br[6]_pad  ;
	input \h1rdt7_br[7]_pad  ;
	input \h1rdt7_br[8]_pad  ;
	input \h1rdt7_br[9]_pad  ;
	input \h1rdt7_dma[0]_pad  ;
	input \h1rdt7_dma[10]_pad  ;
	input \h1rdt7_dma[11]_pad  ;
	input \h1rdt7_dma[12]_pad  ;
	input \h1rdt7_dma[13]_pad  ;
	input \h1rdt7_dma[14]_pad  ;
	input \h1rdt7_dma[15]_pad  ;
	input \h1rdt7_dma[16]_pad  ;
	input \h1rdt7_dma[17]_pad  ;
	input \h1rdt7_dma[18]_pad  ;
	input \h1rdt7_dma[19]_pad  ;
	input \h1rdt7_dma[1]_pad  ;
	input \h1rdt7_dma[20]_pad  ;
	input \h1rdt7_dma[21]_pad  ;
	input \h1rdt7_dma[22]_pad  ;
	input \h1rdt7_dma[23]_pad  ;
	input \h1rdt7_dma[24]_pad  ;
	input \h1rdt7_dma[25]_pad  ;
	input \h1rdt7_dma[26]_pad  ;
	input \h1rdt7_dma[27]_pad  ;
	input \h1rdt7_dma[28]_pad  ;
	input \h1rdt7_dma[29]_pad  ;
	input \h1rdt7_dma[2]_pad  ;
	input \h1rdt7_dma[30]_pad  ;
	input \h1rdt7_dma[31]_pad  ;
	input \h1rdt7_dma[3]_pad  ;
	input \h1rdt7_dma[4]_pad  ;
	input \h1rdt7_dma[5]_pad  ;
	input \h1rdt7_dma[6]_pad  ;
	input \h1rdt7_dma[7]_pad  ;
	input \h1rdt7_dma[8]_pad  ;
	input \h1rdt7_dma[9]_pad  ;
	input \h1rdy0_br_pad  ;
	input \h1rdy0_dma_pad  ;
	input \h1rdy1_br_pad  ;
	input \h1rdy1_dma_pad  ;
	input \h1rdy2_br_pad  ;
	input \h1rdy2_dma_pad  ;
	input \h1rdy3_br_pad  ;
	input \h1rdy3_dma_pad  ;
	input \h1rdy4_br_pad  ;
	input \h1rdy4_dma_pad  ;
	input \h1rdy5_br_pad  ;
	input \h1rdy5_dma_pad  ;
	input \h1rdy6_br_pad  ;
	input \h1rdy6_dma_pad  ;
	input \h1rdy7_br_pad  ;
	input \h1rdy7_dma_pad  ;
	input \h1rp0_br[0]_pad  ;
	input \h1rp0_br[1]_pad  ;
	input \h1rp0_dma[0]_pad  ;
	input \h1rp0_dma[1]_pad  ;
	input \h1rp1_br[0]_pad  ;
	input \h1rp1_br[1]_pad  ;
	input \h1rp1_dma[0]_pad  ;
	input \h1rp1_dma[1]_pad  ;
	input \h1rp2_br[0]_pad  ;
	input \h1rp2_br[1]_pad  ;
	input \h1rp2_dma[0]_pad  ;
	input \h1rp2_dma[1]_pad  ;
	input \h1rp3_br[0]_pad  ;
	input \h1rp3_br[1]_pad  ;
	input \h1rp3_dma[0]_pad  ;
	input \h1rp3_dma[1]_pad  ;
	input \h1rp4_br[0]_pad  ;
	input \h1rp4_br[1]_pad  ;
	input \h1rp4_dma[0]_pad  ;
	input \h1rp4_dma[1]_pad  ;
	input \h1rp5_br[0]_pad  ;
	input \h1rp5_br[1]_pad  ;
	input \h1rp5_dma[0]_pad  ;
	input \h1rp5_dma[1]_pad  ;
	input \h1rp6_br[0]_pad  ;
	input \h1rp6_br[1]_pad  ;
	input \h1rp6_dma[0]_pad  ;
	input \h1rp6_dma[1]_pad  ;
	input \h1rp7_br[0]_pad  ;
	input \h1rp7_br[1]_pad  ;
	input \h1rp7_dma[0]_pad  ;
	input \h1rp7_dma[1]_pad  ;
	input \h1size[0]_pad  ;
	input \h1size[1]_pad  ;
	input \h1size[2]_pad  ;
	input \h1write_pad  ;
	input \haddr[0]_pad  ;
	input \haddr[1]_pad  ;
	input \haddr[2]_pad  ;
	input \haddr[3]_pad  ;
	input \haddr[4]_pad  ;
	input \haddr[5]_pad  ;
	input \haddr[6]_pad  ;
	input \haddr[7]_pad  ;
	input \haddr[8]_pad  ;
	input \hrdata_reg[0]_pad  ;
	input \hrdata_reg[10]_pad  ;
	input \hrdata_reg[11]_pad  ;
	input \hrdata_reg[12]_pad  ;
	input \hrdata_reg[13]_pad  ;
	input \hrdata_reg[14]_pad  ;
	input \hrdata_reg[15]_pad  ;
	input \hrdata_reg[16]_pad  ;
	input \hrdata_reg[17]_pad  ;
	input \hrdata_reg[18]_pad  ;
	input \hrdata_reg[19]_pad  ;
	input \hrdata_reg[1]_pad  ;
	input \hrdata_reg[20]_pad  ;
	input \hrdata_reg[21]_pad  ;
	input \hrdata_reg[22]_pad  ;
	input \hrdata_reg[23]_pad  ;
	input \hrdata_reg[24]_pad  ;
	input \hrdata_reg[25]_pad  ;
	input \hrdata_reg[26]_pad  ;
	input \hrdata_reg[27]_pad  ;
	input \hrdata_reg[28]_pad  ;
	input \hrdata_reg[29]_pad  ;
	input \hrdata_reg[2]_pad  ;
	input \hrdata_reg[30]_pad  ;
	input \hrdata_reg[31]_pad  ;
	input \hrdata_reg[3]_pad  ;
	input \hrdata_reg[4]_pad  ;
	input \hrdata_reg[5]_pad  ;
	input \hrdata_reg[6]_pad  ;
	input \hrdata_reg[7]_pad  ;
	input \hrdata_reg[8]_pad  ;
	input \hrdata_reg[9]_pad  ;
	input hreadyin_pad ;
	input hreadyout_br_pad ;
	input \hresp_br[0]_pad  ;
	input \hresp_br[1]_pad  ;
	input hsel_br_pad ;
	input hsel_reg_pad ;
	input \hsize[0]_pad  ;
	input \hsize[1]_pad  ;
	input \hsize[2]_pad  ;
	input \htrans[0]_pad  ;
	input \htrans[1]_pad  ;
	input \hwdata[0]_pad  ;
	input \hwdata[10]_pad  ;
	input \hwdata[11]_pad  ;
	input \hwdata[12]_pad  ;
	input \hwdata[13]_pad  ;
	input \hwdata[14]_pad  ;
	input \hwdata[15]_pad  ;
	input \hwdata[16]_pad  ;
	input \hwdata[17]_pad  ;
	input \hwdata[18]_pad  ;
	input \hwdata[19]_pad  ;
	input \hwdata[1]_pad  ;
	input \hwdata[20]_pad  ;
	input \hwdata[21]_pad  ;
	input \hwdata[22]_pad  ;
	input \hwdata[23]_pad  ;
	input \hwdata[24]_pad  ;
	input \hwdata[25]_pad  ;
	input \hwdata[26]_pad  ;
	input \hwdata[27]_pad  ;
	input \hwdata[28]_pad  ;
	input \hwdata[29]_pad  ;
	input \hwdata[2]_pad  ;
	input \hwdata[30]_pad  ;
	input \hwdata[31]_pad  ;
	input \hwdata[3]_pad  ;
	input \hwdata[4]_pad  ;
	input \hwdata[5]_pad  ;
	input \hwdata[6]_pad  ;
	input \hwdata[7]_pad  ;
	input \hwdata[8]_pad  ;
	input \hwdata[9]_pad  ;
	input hwrite_pad ;
	input \m1_mux_hrdy_df_reg/NET0131  ;
	input \m1_mux_hrmxnof_reg/NET0131  ;
	input \m1_mux_hrp_df_reg[0]/NET0131  ;
	input \m1_mux_mux_no_reg[0]/NET0131  ;
	input \m1_mux_mux_no_reg[1]/NET0131  ;
	input \m1_mux_mux_no_reg[2]/NET0131  ;
	input \m1_mux_mux_no_reg[3]/NET0131  ;
	output \_al_n1  ;
	output \g16/_0_  ;
	output \g58487/_0_  ;
	output \g58489/_0_  ;
	output \g58491/_0_  ;
	output \g58493/_0_  ;
	output \g58495/_0_  ;
	output \g58497/_0_  ;
	output \g58499/_0_  ;
	output \g58500/_0_  ;
	output \g58501/_0_  ;
	output \g58502/_0_  ;
	output \g58504/_0_  ;
	output \g58505/_0_  ;
	output \g58507/_0_  ;
	output \g58508/_0_  ;
	output \g58509/_0_  ;
	output \g58510/_0_  ;
	output \g58556/_0_  ;
	output \g58557/_0_  ;
	output \g58558/_0_  ;
	output \g58559/_0_  ;
	output \g58560/_0_  ;
	output \g58561/_0_  ;
	output \g58562/_0_  ;
	output \g58563/_0_  ;
	output \g58566/_0_  ;
	output \g58567/_0_  ;
	output \g58568/_0_  ;
	output \g58569/_0_  ;
	output \g58570/_0_  ;
	output \g58571/_0_  ;
	output \g58572/_0_  ;
	output \g58573/_0_  ;
	output \g58574/_0_  ;
	output \g58575/_0_  ;
	output \g58576/_0_  ;
	output \g58577/_0_  ;
	output \g58578/_0_  ;
	output \g58579/_0_  ;
	output \g58580/_0_  ;
	output \g58581/_0_  ;
	output \g58584/_0_  ;
	output \g58585/_0_  ;
	output \g58586/_0_  ;
	output \g58587/_0_  ;
	output \g58588/_0_  ;
	output \g58589/_0_  ;
	output \g58590/_0_  ;
	output \g58591/_0_  ;
	output \g58592/_0_  ;
	output \g58593/_0_  ;
	output \g58594/_0_  ;
	output \g58595/_0_  ;
	output \g58596/_0_  ;
	output \g58597/_0_  ;
	output \g58598/_0_  ;
	output \g58599/_0_  ;
	output \g58600/_0_  ;
	output \g58601/_0_  ;
	output \g58602/_0_  ;
	output \g58603/_0_  ;
	output \g58604/_0_  ;
	output \g58605/_0_  ;
	output \g58606/_0_  ;
	output \g58607/_0_  ;
	output \g58608/_0_  ;
	output \g58609/_0_  ;
	output \g58610/_0_  ;
	output \g58611/_0_  ;
	output \g58612/_0_  ;
	output \g58613/_0_  ;
	output \g58614/_0_  ;
	output \g58615/_0_  ;
	output \g58616/_0_  ;
	output \g58617/_0_  ;
	output \g58618/_0_  ;
	output \g58619/_0_  ;
	output \g58620/_0_  ;
	output \g58621/_0_  ;
	output \g58622/_0_  ;
	output \g58623/_0_  ;
	output \g58624/_0_  ;
	output \g58625/_0_  ;
	output \g58626/_0_  ;
	output \g58627/_0_  ;
	output \g58723/_0_  ;
	output \g58734/_0_  ;
	output \g58737/_0_  ;
	output \g58741/_0_  ;
	output \g58749/_0_  ;
	output \g58754/_0_  ;
	output \g58762/_0_  ;
	output \g58763/_0_  ;
	output \g58764/_0_  ;
	output \g58765/_0_  ;
	output \g58766/_0_  ;
	output \g58767/_0_  ;
	output \g58768/_0_  ;
	output \g58769/_0_  ;
	output \g58770/_0_  ;
	output \g58771/_0_  ;
	output \g59788/_0_  ;
	output \g59832/_0_  ;
	output \g59873/_0_  ;
	output \g59874/_0_  ;
	output \g59893/_0_  ;
	output \g59894/_0_  ;
	output \g59895/_0_  ;
	output \g59896/_0_  ;
	output \g59923/_0_  ;
	output \g60031/_0_  ;
	output \g60032/_0_  ;
	output \g60033/_0_  ;
	output \g60036/_0_  ;
	output \g60037/_0_  ;
	output \g60038/_0_  ;
	output \g60165/_0_  ;
	output \g60186/_2__syn_2  ;
	output \g60187/_0_  ;
	output \g60188/_0_  ;
	output \g60258/_0_  ;
	output \g60259/_0_  ;
	output \g60260/_0_  ;
	output \g60261/_0_  ;
	output \g60263/_0_  ;
	output \g60264/_0_  ;
	output \g60265/_0_  ;
	output \g60266/_0_  ;
	output \g60267/_0_  ;
	output \g60303/_3_  ;
	output \g60360/_0_  ;
	output \g60361/_0_  ;
	output \g60401/_00_  ;
	output \g60428/_0_  ;
	output \g60429/_0_  ;
	output \g60448/_0_  ;
	output \g60449/_0_  ;
	output \g60974/_0_  ;
	output \g61072/_0_  ;
	output \g61073/_0_  ;
	output \g61074/_0_  ;
	output \g61075/_0_  ;
	output \g61076/_0_  ;
	output \g61077/_0_  ;
	output \g61078/_0_  ;
	output \g61079/_0_  ;
	output \g61486/_0_  ;
	output \g61502/_3_  ;
	output \g61879/_0_  ;
	output \g62077/_0_  ;
	output \g62078/_0_  ;
	output \g62079/_0_  ;
	output \g62080/_0_  ;
	output \g62081/_0_  ;
	output \g62082/_0_  ;
	output \g62083/_0_  ;
	output \g62084/_0_  ;
	output \g62085/_0_  ;
	output \g62086/_0_  ;
	output \g62087/_0_  ;
	output \g62088/_0_  ;
	output \g62089/_0_  ;
	output \g62090/_0_  ;
	output \g62091/_0_  ;
	output \g62629/_0_  ;
	output \g62630/_0_  ;
	output \g62631/_0_  ;
	output \g62632/_0_  ;
	output \g62633/_0_  ;
	output \g62634/_0_  ;
	output \g62635/_0_  ;
	output \g62637/_0_  ;
	output \g62638/_0_  ;
	output \g62639/_0_  ;
	output \g62641/_0_  ;
	output \g62643/_0_  ;
	output \g62645/_0_  ;
	output \g62646/_0_  ;
	output \g62647/_0_  ;
	output \g62648/_0_  ;
	output \g62649/_0_  ;
	output \g62650/_0_  ;
	output \g62651/_0_  ;
	output \g62652/_0_  ;
	output \g62655/_0_  ;
	output \g62656/_0_  ;
	output \g62657/_0_  ;
	output \g62658/_0_  ;
	output \g62659/_0_  ;
	output \g62660/_0_  ;
	output \g62661/_0_  ;
	output \g62662/_0_  ;
	output \g62663/_0_  ;
	output \g62664/_0_  ;
	output \g62665/_0_  ;
	output \g62667/_0_  ;
	output \g62668/_0_  ;
	output \g62669/_0_  ;
	output \g62670/_0_  ;
	output \g62671/_0_  ;
	output \g62672/_0_  ;
	output \g62673/_0_  ;
	output \g62674/_0_  ;
	output \g62675/_0_  ;
	output \g62676/_0_  ;
	output \g62677/_0_  ;
	output \g62678/_0_  ;
	output \g62679/_0_  ;
	output \g62680/_0_  ;
	output \g62681/_0_  ;
	output \g62682/_0_  ;
	output \g62683/_0_  ;
	output \g62684/_0_  ;
	output \g62685/_0_  ;
	output \g62686/_0_  ;
	output \g62687/_0_  ;
	output \g62688/_0_  ;
	output \g62689/_0_  ;
	output \g62690/_0_  ;
	output \g62691/_0_  ;
	output \g62692/_0_  ;
	output \g62693/_0_  ;
	output \g62694/_0_  ;
	output \g62695/_0_  ;
	output \g62696/_0_  ;
	output \g62697/_0_  ;
	output \g62698/_0_  ;
	output \g62699/_0_  ;
	output \g62700/_0_  ;
	output \g62701/_0_  ;
	output \g62702/_0_  ;
	output \g62703/_0_  ;
	output \g62704/_0_  ;
	output \g62705/_0_  ;
	output \g62706/_0_  ;
	output \g62707/_0_  ;
	output \g62708/_0_  ;
	output \g62709/_0_  ;
	output \g62710/_0_  ;
	output \g62711/_0_  ;
	output \g62712/_0_  ;
	output \g62713/_0_  ;
	output \g62714/_0_  ;
	output \g62715/_0_  ;
	output \g62716/_0_  ;
	output \g62721/_0_  ;
	output \g62722/_0_  ;
	output \g62723/_0_  ;
	output \g62725/_0_  ;
	output \g62726/_0_  ;
	output \g62727/_0_  ;
	output \g62728/_0_  ;
	output \g62729/_0_  ;
	output \g62730/_0_  ;
	output \g62731/_0_  ;
	output \g62732/_0_  ;
	output \g62733/_0_  ;
	output \g62734/_0_  ;
	output \g62735/_0_  ;
	output \g62736/_0_  ;
	output \g62737/_0_  ;
	output \g62738/_0_  ;
	output \g62739/_0_  ;
	output \g62740/_0_  ;
	output \g62741/_0_  ;
	output \g62742/_0_  ;
	output \g62743/_0_  ;
	output \g62744/_0_  ;
	output \g62745/_0_  ;
	output \g62746/_0_  ;
	output \g62747/_0_  ;
	output \g62748/_0_  ;
	output \g62749/_0_  ;
	output \g62750/_0_  ;
	output \g62751/_0_  ;
	output \g62752/_0_  ;
	output \g62753/_0_  ;
	output \g62754/_0_  ;
	output \g62755/_0_  ;
	output \g62756/_0_  ;
	output \g62757/_0_  ;
	output \g62758/_0_  ;
	output \g62759/_0_  ;
	output \g62760/_0_  ;
	output \g62761/_0_  ;
	output \g62762/_0_  ;
	output \g62763/_0_  ;
	output \g62764/_0_  ;
	output \g62765/_0_  ;
	output \g62766/_0_  ;
	output \g62767/_0_  ;
	output \g62768/_0_  ;
	output \g62769/_0_  ;
	output \g62770/_0_  ;
	output \g62771/_0_  ;
	output \g62772/_0_  ;
	output \g62773/_0_  ;
	output \g62774/_0_  ;
	output \g62775/_0_  ;
	output \g62776/_0_  ;
	output \g62777/_0_  ;
	output \g62778/_0_  ;
	output \g62779/_0_  ;
	output \g62780/_0_  ;
	output \g62781/_0_  ;
	output \g62783/_0_  ;
	output \g62784/_0_  ;
	output \g62785/_0_  ;
	output \g62786/_0_  ;
	output \g62787/_0_  ;
	output \g62788/_0_  ;
	output \g62789/_0_  ;
	output \g62790/_0_  ;
	output \g62791/_0_  ;
	output \g62792/_0_  ;
	output \g62793/_0_  ;
	output \g62794/_0_  ;
	output \g62795/_0_  ;
	output \g62797/_0_  ;
	output \g62798/_0_  ;
	output \g62799/_0_  ;
	output \g62800/_0_  ;
	output \g62801/_0_  ;
	output \g62802/_0_  ;
	output \g62803/_0_  ;
	output \g62804/_0_  ;
	output \g62805/_0_  ;
	output \g62806/_0_  ;
	output \g62807/_0_  ;
	output \g62808/_0_  ;
	output \g62809/_0_  ;
	output \g62810/_0_  ;
	output \g62811/_0_  ;
	output \g62812/_0_  ;
	output \g62813/_0_  ;
	output \g62814/_0_  ;
	output \g62815/_0_  ;
	output \g62816/_0_  ;
	output \g62817/_0_  ;
	output \g62818/_0_  ;
	output \g63108/_0_  ;
	output \g63117/_0_  ;
	output \g63125/_0_  ;
	output \g63126/_0_  ;
	output \g63127/_0_  ;
	output \g63128/_0_  ;
	output \g63129/_0_  ;
	output \g63130/_0_  ;
	output \g63131/_0_  ;
	output \g63132/_0_  ;
	output \g63133/_0_  ;
	output \g63134/_0_  ;
	output \g63135/_0_  ;
	output \g63136/_0_  ;
	output \g63137/_0_  ;
	output \g63138/_0_  ;
	output \g63139/_0_  ;
	output \g63140/_0_  ;
	output \g63141/_0_  ;
	output \g63142/_0_  ;
	output \g63143/_0_  ;
	output \g63144/_0_  ;
	output \g63145/_0_  ;
	output \g63146/_0_  ;
	output \g63147/_0_  ;
	output \g63148/_0_  ;
	output \g63149/_0_  ;
	output \g63150/_0_  ;
	output \g63151/_0_  ;
	output \g63152/_0_  ;
	output \g63153/_0_  ;
	output \g63154/_0_  ;
	output \g63155/_0_  ;
	output \g63156/_0_  ;
	output \g63157/_0_  ;
	output \g63159/_0_  ;
	output \g63160/_0_  ;
	output \g63161/_0_  ;
	output \g63162/_0_  ;
	output \g63163/_0_  ;
	output \g63164/_0_  ;
	output \g63165/_0_  ;
	output \g63166/_0_  ;
	output \g63167/_0_  ;
	output \g63168/_0_  ;
	output \g63169/_0_  ;
	output \g63170/_0_  ;
	output \g63171/_0_  ;
	output \g63172/_0_  ;
	output \g63173/_0_  ;
	output \g63174/_0_  ;
	output \g63175/_0_  ;
	output \g63176/_0_  ;
	output \g63177/_0_  ;
	output \g63178/_0_  ;
	output \g63179/_0_  ;
	output \g63180/_0_  ;
	output \g63181/_0_  ;
	output \g63182/_0_  ;
	output \g63183/_0_  ;
	output \g63184/_0_  ;
	output \g63185/_0_  ;
	output \g63186/_0_  ;
	output \g63187/_0_  ;
	output \g63188/_0_  ;
	output \g63189/_0_  ;
	output \g63190/_0_  ;
	output \g63191/_0_  ;
	output \g63192/_0_  ;
	output \g63193/_0_  ;
	output \g63194/_0_  ;
	output \g63195/_0_  ;
	output \g63196/_0_  ;
	output \g63197/_0_  ;
	output \g63198/_0_  ;
	output \g63199/_0_  ;
	output \g63200/_0_  ;
	output \g63201/_0_  ;
	output \g63202/_0_  ;
	output \g63203/_0_  ;
	output \g63204/_0_  ;
	output \g63205/_0_  ;
	output \g63206/_0_  ;
	output \g63207/_0_  ;
	output \g63208/_0_  ;
	output \g63209/_0_  ;
	output \g63210/_0_  ;
	output \g63211/_0_  ;
	output \g63212/_0_  ;
	output \g63213/_0_  ;
	output \g63214/_0_  ;
	output \g63215/_0_  ;
	output \g63216/_0_  ;
	output \g63217/_0_  ;
	output \g63218/_0_  ;
	output \g63219/_0_  ;
	output \g63220/_0_  ;
	output \g63221/_0_  ;
	output \g63222/_0_  ;
	output \g63223/_0_  ;
	output \g63224/_0_  ;
	output \g63225/_0_  ;
	output \g63226/_0_  ;
	output \g63228/_0_  ;
	output \g63229/_0_  ;
	output \g63231/_0_  ;
	output \g63232/_0_  ;
	output \g63233/_0_  ;
	output \g63234/_0_  ;
	output \g63235/_0_  ;
	output \g63236/_0_  ;
	output \g63237/_0_  ;
	output \g63238/_0_  ;
	output \g63239/_0_  ;
	output \g63240/_0_  ;
	output \g63241/_0_  ;
	output \g63242/_0_  ;
	output \g63244/_0_  ;
	output \g63246/_0_  ;
	output \g63247/_0_  ;
	output \g63248/_0_  ;
	output \g63249/_0_  ;
	output \g63250/_0_  ;
	output \g63251/_0_  ;
	output \g63252/_0_  ;
	output \g63253/_0_  ;
	output \g63254/_0_  ;
	output \g63255/_0_  ;
	output \g63256/_0_  ;
	output \g63257/_0_  ;
	output \g63258/_0_  ;
	output \g63259/_0_  ;
	output \g63260/_0_  ;
	output \g63261/_0_  ;
	output \g63262/_0_  ;
	output \g63263/_0_  ;
	output \g63264/_0_  ;
	output \g63265/_0_  ;
	output \g63266/_0_  ;
	output \g63267/_0_  ;
	output \g63268/_0_  ;
	output \g63269/_0_  ;
	output \g63270/_0_  ;
	output \g63272/_0_  ;
	output \g63291/_0_  ;
	output \g63292/_0_  ;
	output \g63293/_0_  ;
	output \g63294/_0_  ;
	output \g63295/_0_  ;
	output \g63298/_0_  ;
	output \g63299/_0_  ;
	output \g63300/_0_  ;
	output \g63301/_0_  ;
	output \g63302/_0_  ;
	output \g63303/_0_  ;
	output \g63304/_0_  ;
	output \g63305/_0_  ;
	output \g63306/_0_  ;
	output \g63307/_0_  ;
	output \g63308/_0_  ;
	output \g63309/_0_  ;
	output \g63310/_0_  ;
	output \g63311/_0_  ;
	output \g63312/_0_  ;
	output \g63313/_0_  ;
	output \g63314/_0_  ;
	output \g63315/_0_  ;
	output \g63316/_0_  ;
	output \g63317/_0_  ;
	output \g63318/_0_  ;
	output \g63320/_0_  ;
	output \g63322/_0_  ;
	output \g63323/_0_  ;
	output \g63324/_0_  ;
	output \g63325/_0_  ;
	output \g63326/_0_  ;
	output \g63327/_0_  ;
	output \g63328/_0_  ;
	output \g63329/_0_  ;
	output \g63330/_0_  ;
	output \g63331/_0_  ;
	output \g63332/_0_  ;
	output \g63333/_0_  ;
	output \g63334/_0_  ;
	output \g63335/_0_  ;
	output \g63336/_0_  ;
	output \g63337/_0_  ;
	output \g63338/_0_  ;
	output \g63339/_0_  ;
	output \g63340/_0_  ;
	output \g63341/_0_  ;
	output \g63342/_0_  ;
	output \g63343/_0_  ;
	output \g63344/_0_  ;
	output \g63345/_0_  ;
	output \g63346/_0_  ;
	output \g63347/_0_  ;
	output \g63348/_0_  ;
	output \g63349/_0_  ;
	output \g63350/_0_  ;
	output \g63351/_0_  ;
	output \g63352/_0_  ;
	output \g63353/_0_  ;
	output \g63354/_0_  ;
	output \g63355/_0_  ;
	output \g63356/_0_  ;
	output \g63357/_0_  ;
	output \g63358/_0_  ;
	output \g63359/_0_  ;
	output \g63360/_0_  ;
	output \g63361/_0_  ;
	output \g63362/_0_  ;
	output \g63363/_0_  ;
	output \g63364/_0_  ;
	output \g63365/_0_  ;
	output \g63366/_0_  ;
	output \g63367/_0_  ;
	output \g63368/_0_  ;
	output \g63369/_0_  ;
	output \g63370/_0_  ;
	output \g63371/_0_  ;
	output \g63372/_0_  ;
	output \g63373/_0_  ;
	output \g63374/_0_  ;
	output \g63375/_0_  ;
	output \g63376/_0_  ;
	output \g63377/_0_  ;
	output \g63378/_0_  ;
	output \g63379/_0_  ;
	output \g63380/_0_  ;
	output \g63383/_3_  ;
	output \g63386/_0_  ;
	output \g63387/_0_  ;
	output \g63388/_0_  ;
	output \g63389/_0_  ;
	output \g63390/_0_  ;
	output \g63391/_0_  ;
	output \g63392/_0_  ;
	output \g63419/_0_  ;
	output \g63421/_0_  ;
	output \g63422/_0_  ;
	output \g63423/_0_  ;
	output \g63424/_0_  ;
	output \g63425/_0_  ;
	output \g63536/_3_  ;
	output \g63625/_0_  ;
	output \g63628/_0_  ;
	output \g63871/_0_  ;
	output \g63874/_0_  ;
	output \g63889/_0_  ;
	output \g63933/_0_  ;
	output \g63945/_0_  ;
	output \g63959/_0_  ;
	output \g63962/_0_  ;
	output \g63974/_0_  ;
	output \g63977/_0_  ;
	output \g64035/_0_  ;
	output \g64435/_3_  ;
	output \g64939/_0_  ;
	output \g65149/_0_  ;
	output \g65632/_3_  ;
	output \g65633/_0_  ;
	output \g65634/_0_  ;
	output \g65635/_0_  ;
	output \g65636/_0_  ;
	output \g65638/_3_  ;
	output \g65640/_3_  ;
	output \g65999/_0_  ;
	output \g66912/_0_  ;
	output \g66914/_0_  ;
	output \g67555/_3_  ;
	output \g67564/_3_  ;
	output \g67567/_3_  ;
	output \g67735/_0_  ;
	output \g67736/_0_  ;
	output \g67737/_0_  ;
	output \g67738/_0_  ;
	output \g67758/_0_  ;
	output \g67760/_0_  ;
	output \g67761/_0_  ;
	output \g67763/_0_  ;
	output \g67766/_0_  ;
	output \g67810/_0_  ;
	output \g67816/_0_  ;
	output \g67902/_0_  ;
	output \g67927/_0_  ;
	output \g67936/_0_  ;
	output \g68067/_0_  ;
	output \g68068/_0_  ;
	output \g68069/_0_  ;
	output \g68070/_0_  ;
	output \g68071/_0_  ;
	output \g68072/_0_  ;
	output \g68073/_0_  ;
	output \g68074/_0_  ;
	output \g68075/_0_  ;
	output \g68076/_0_  ;
	output \g68077/_0_  ;
	output \g68078/_0_  ;
	output \g68079/_0_  ;
	output \g68080/_0_  ;
	output \g68081/_0_  ;
	output \g68082/_0_  ;
	output \g68083/_0_  ;
	output \g68084/_0_  ;
	output \g68085/_0_  ;
	output \g68086/_0_  ;
	output \g68087/_0_  ;
	output \g68088/_0_  ;
	output \g68089/_0_  ;
	output \g68090/_0_  ;
	output \g68091/_0_  ;
	output \g68096/_0_  ;
	output \g68160/_0_  ;
	output \g68218/_0_  ;
	output \g68219/_0_  ;
	output \g68220/_0_  ;
	output \g68221/_0_  ;
	output \g68222/_0_  ;
	output \g68226/_0_  ;
	output \g68247/_0_  ;
	output \g68252/_0_  ;
	output \g68632/_0_  ;
	output \g68633/_0_  ;
	output \g68635/_0_  ;
	output \g68640/_0_  ;
	output \g68642/_0_  ;
	output \g68643/_0_  ;
	output \g68644/_0_  ;
	output \g68645/_0_  ;
	output \g68649/_0_  ;
	output \g68668/_2_  ;
	output \g68670/_0_  ;
	output \g68681/_3_  ;
	output \g68689/_0_  ;
	output \g68690/_0_  ;
	output \g68691/_0_  ;
	output \g68692/_0_  ;
	output \g68693/_0_  ;
	output \g68694/_0_  ;
	output \g68695/_0_  ;
	output \g68737/_0_  ;
	output \g68742/_0_  ;
	output \g68745/_0_  ;
	output \g68750/_0_  ;
	output \g68759/_0_  ;
	output \g68761/_0_  ;
	output \g68774/_0_  ;
	output \g68775/_0_  ;
	output \g68776/_0_  ;
	output \g68777/_0_  ;
	output \g68778/_0_  ;
	output \g68780/_0_  ;
	output \g68781/_0_  ;
	output \g68782/_0_  ;
	output \g68783/_0_  ;
	output \g68784/_0_  ;
	output \g68785/_0_  ;
	output \g68786/_0_  ;
	output \g68787/_0_  ;
	output \g68790/_0_  ;
	output \g68791/_0_  ;
	output \g68793/_0_  ;
	output \g68794/_0_  ;
	output \g68795/_0_  ;
	output \g68796/_0_  ;
	output \g68797/_0_  ;
	output \g68804/_0_  ;
	output \g68805/_0_  ;
	output \g68807/_0_  ;
	output \g68809/_0_  ;
	output \g68864/_3_  ;
	output \g68865/_3_  ;
	output \g68866/_3_  ;
	output \g68867/_3_  ;
	output \g68868/_3_  ;
	output \g68869/_3_  ;
	output \g68870/_3_  ;
	output \g68871/_3_  ;
	output \g68872/_3_  ;
	output \g68873/_3_  ;
	output \g68874/_3_  ;
	output \g68875/_3_  ;
	output \g68876/_3_  ;
	output \g68877/_3_  ;
	output \g68878/_3_  ;
	output \g68879/_3_  ;
	output \g68880/_3_  ;
	output \g68881/_3_  ;
	output \g68882/_3_  ;
	output \g68883/_3_  ;
	output \g68884/_3_  ;
	output \g68885/_3_  ;
	output \g68886/_3_  ;
	output \g68887/_3_  ;
	output \g68888/_3_  ;
	output \g68889/_3_  ;
	output \g68890/_3_  ;
	output \g68891/_3_  ;
	output \g68892/_3_  ;
	output \g68893/_3_  ;
	output \g68894/_3_  ;
	output \g68895/_3_  ;
	output \g69037/_1__syn_2  ;
	output \g69077/_0_  ;
	output \g69081/_0_  ;
	output \g69084/_0_  ;
	output \g69085/_0_  ;
	output \g69086/_0_  ;
	output \g69088/_0_  ;
	output \g69094/_0_  ;
	output \g69095/_0_  ;
	output \g69097/_0_  ;
	output \g69114/_3_  ;
	output \g69116/_3_  ;
	output \g69118/_3_  ;
	output \g69120/_3_  ;
	output \g69122/_3_  ;
	output \g69124/_3_  ;
	output \g69126/_3_  ;
	output \g69128/_3_  ;
	output \g69581/_3_  ;
	output \g70303/_1__syn_2  ;
	output \g70304/_1__syn_2  ;
	output \g70305/_1__syn_2  ;
	output \g70306/_1__syn_2  ;
	output \g70353/_1__syn_2  ;
	output \g70359/_2_  ;
	output \g70364/_1__syn_2  ;
	output \g70375/_1__syn_2  ;
	output \g70380/_2_  ;
	output \g70383/_1__syn_2  ;
	output \g70394/_2_  ;
	output \g70395/_2_  ;
	output \g70396/_1__syn_2  ;
	output \g70398/_1__syn_2  ;
	output \g70407/_1_  ;
	output \g70416/_1__syn_2  ;
	output \g70418/_1__syn_2  ;
	output \g70419/_2_  ;
	output \g70424/_1_  ;
	output \g70465/_2_  ;
	output \g70511/_1_  ;
	output \g70512/_1_  ;
	output \g70513/_2_  ;
	output \g70514/_2_  ;
	output \g70516/_2_  ;
	output \g70518/_2_  ;
	output \g70519/_2_  ;
	output \g70520/_2_  ;
	output \g70530/_2_  ;
	output \g70534/_3_  ;
	output \g70536/_3_  ;
	output \g70540/_3_  ;
	output \g70541/_2_  ;
	output \g70545/_3_  ;
	output \g70546/_2_  ;
	output \g70547/_2_  ;
	output \g70550/_3_  ;
	output \g70551/_2_  ;
	output \g70552/_2_  ;
	output \g70558/_3_  ;
	output \g70559/_2_  ;
	output \g70560/_2_  ;
	output \g70562/_3_  ;
	output \g70564/_3_  ;
	output \g70567/_3_  ;
	output \g70568/_2_  ;
	output \g70571/_3_  ;
	output \g70577/_0_  ;
	output \g70578/_2_  ;
	output \g70585/_3_  ;
	output \g70586/_2_  ;
	output \g70587/_2_  ;
	output \g70588/_3_  ;
	output \g70602/_3_  ;
	output \g70841/_0_  ;
	output \g70842/_0_  ;
	output \g70843/_0_  ;
	output \g70844/_0_  ;
	output \g70845/_0_  ;
	output \g70846/_0_  ;
	output \g70847/_0_  ;
	output \g70848/_0_  ;
	output \g70849/_0_  ;
	output \g70850/_0_  ;
	output \g70851/_0_  ;
	output \g70852/_0_  ;
	output \g70853/_0_  ;
	output \g70854/_0_  ;
	output \g70855/_0_  ;
	output \g70856/_0_  ;
	output \g70857/_0_  ;
	output \g70858/_0_  ;
	output \g70859/_0_  ;
	output \g70860/_0_  ;
	output \g70861/_0_  ;
	output \g70862/_0_  ;
	output \g70863/_0_  ;
	output \g70864/_0_  ;
	output \g70865/_0_  ;
	output \g70866/_0_  ;
	output \g70867/_0_  ;
	output \g70868/_0_  ;
	output \g70869/_0_  ;
	output \g70870/_0_  ;
	output \g70871/_0_  ;
	output \g70872/_0_  ;
	output \g70944/_1__syn_2  ;
	output \g71042/_1__syn_2  ;
	output \g71064/_1__syn_2  ;
	output \g71065/_1__syn_2  ;
	output \g71076/_1__syn_2  ;
	output \g71077/_1__syn_2  ;
	output \g71202/_1__syn_2  ;
	output \g71204/_1__syn_2  ;
	output \g71236/_0_  ;
	output \g71237/_0_  ;
	output \g71241/_0_  ;
	output \g71242/_0_  ;
	output \g71245/_0_  ;
	output \g71246/_0_  ;
	output \g71306/_0_  ;
	output \g71308/_0_  ;
	output \g71309/_0_  ;
	output \g71310/_0_  ;
	output \g71355/_0_  ;
	output \g71416/_0_  ;
	output \g71417/_0_  ;
	output \g71420/_0_  ;
	output \g71432/_0_  ;
	output \g71434/_0_  ;
	output \g71435/_0_  ;
	output \g71436/_0_  ;
	output \g71446/_0_  ;
	output \g71449/_0_  ;
	output \g71451/_0_  ;
	output \g71452/_0_  ;
	output \g71485/_0_  ;
	output \g71494/_0_  ;
	output \g71499/_0_  ;
	output \g71500/_0_  ;
	output \g71501/_0_  ;
	output \g71502/_0_  ;
	output \g71503/_0_  ;
	output \g71504/_0_  ;
	output \g71505/_0_  ;
	output \g71506/_0_  ;
	output \g71815/_0_  ;
	output \g71823/_0_  ;
	output \g71832/_0_  ;
	output \g71833/_0__syn_2  ;
	output \g71837/_0_  ;
	output \g71838/_0_  ;
	output \g71846/_1__syn_2  ;
	output \g71847/_1__syn_2  ;
	output \g71849/_0_  ;
	output \g71854/_0_  ;
	output \g71858/_1__syn_2  ;
	output \g71859/_1__syn_2  ;
	output \g71863/_0_  ;
	output \g71867/_0_  ;
	output \g71869/_0_  ;
	output \g71872/_1_  ;
	output \g71873/_1__syn_2  ;
	output \g71874/_1__syn_2  ;
	output \g71875/_0_  ;
	output \g71877/_1__syn_2  ;
	output \g71881/_0_  ;
	output \g71906/_0_  ;
	output \g71907/_1__syn_2  ;
	output \g71910/_0_  ;
	output \g71911/_0_  ;
	output \g71912/_1__syn_2  ;
	output \g71913/_1__syn_2  ;
	output \g71914/_1__syn_2  ;
	output \g71918/_0_  ;
	output \g71921/_0_  ;
	output \g71922/_0_  ;
	output \g71929/_1__syn_2  ;
	output \g71931/_1__syn_2  ;
	output \g71938/_1__syn_2  ;
	output \g71942/_0_  ;
	output \g71946/_1__syn_2  ;
	output \g71947/_0_  ;
	output \g71951/_0_  ;
	output \g71958/_1__syn_2  ;
	output \g71965/_0_  ;
	output \g71970/_1__syn_2  ;
	output \g71972/_1__syn_2  ;
	output \g71973/_1__syn_2  ;
	output \g71986/_1__syn_2  ;
	output \g71987/_1__syn_2  ;
	output \g71990/_1__syn_2  ;
	output \g71991/_1__syn_2  ;
	output \g71992/_1__syn_2  ;
	output \g71994/_1__syn_2  ;
	output \g71997/_1__syn_2  ;
	output \g72001/_1__syn_2  ;
	output \g72013/_1__syn_2  ;
	output \g72021/_1__syn_2  ;
	output \g72030/_0_  ;
	output \g72031/_0__syn_2  ;
	output \g72036/_1__syn_2  ;
	output \g72038/_0_  ;
	output \g72042/_1__syn_2  ;
	output \g72047/_1__syn_2  ;
	output \g72048/_1__syn_2  ;
	output \g72049/_1__syn_2  ;
	output \g72056/_0_  ;
	output \g72064/_1__syn_2  ;
	output \g72073/_1__syn_2  ;
	output \g72075/_0_  ;
	output \g72078/_0_  ;
	output \g72081/_0_  ;
	output \g72091/_0_  ;
	output \g72096/_0_  ;
	output \g72100/_1__syn_2  ;
	output \g72113/_0_  ;
	output \g72118/_0_  ;
	output \g72121/_1__syn_2  ;
	output \g72122/_1__syn_2  ;
	output \g72125/_1__syn_2  ;
	output \g72128/_0_  ;
	output \g72140/_0_  ;
	output \g72144/_1__syn_2  ;
	output \g72154/_1__syn_2  ;
	output \g72159/_0_  ;
	output \g72164/_1__syn_2  ;
	output \g72165/_1__syn_2  ;
	output \g72167/_1__syn_2  ;
	output \g72170/_1__syn_2  ;
	output \g72172/_1__syn_2  ;
	output \g72173/_0_  ;
	output \g72177/_1__syn_2  ;
	output \g72189/_0_  ;
	output \g72194/_0_  ;
	output \g72196/_0_  ;
	output \g72198/_0_  ;
	output \g72206/_1__syn_2  ;
	output \g72209/_1__syn_2  ;
	output \g72210/_1__syn_2  ;
	output \g72211/_0_  ;
	output \g72215/_0_  ;
	output \g72227/_1__syn_2  ;
	output \g72229/_1__syn_2  ;
	output \g72230/_0_  ;
	output \g72239/_0_  ;
	output \g72250/_3_  ;
	output \g72251/_3_  ;
	output \g72252/_3_  ;
	output \g72253/_3_  ;
	output \g72254/_3_  ;
	output \g72255/_3_  ;
	output \g72256/_3_  ;
	output \g72257/_3_  ;
	output \g72259/_3_  ;
	output \g72260/_3_  ;
	output \g72261/_3_  ;
	output \g72262/_3_  ;
	output \g72263/_3_  ;
	output \g72264/_3_  ;
	output \g72265/_3_  ;
	output \g72266/_3_  ;
	output \g72267/_3_  ;
	output \g72273/_3_  ;
	output \g72275/_3_  ;
	output \g72282/_3_  ;
	output \g72285/_3_  ;
	output \g72293/_3_  ;
	output \g72304/_3_  ;
	output \g72305/_3_  ;
	output \g72306/_3_  ;
	output \g72307/_3_  ;
	output \g72309/_3_  ;
	output \g72310/_3_  ;
	output \g72324/_3_  ;
	output \g72325/_3_  ;
	output \g72326/_3_  ;
	output \g72327/_3_  ;
	output \g72711/_0_  ;
	output \g72763/_0_  ;
	output \g72966/_0_  ;
	output \g72967/_0_  ;
	output \g73018/_0_  ;
	output \g73058/_0_  ;
	output \g73062/_0_  ;
	output \g73067/_0_  ;
	output \g73068/_0_  ;
	output \g73207/_0_  ;
	output \g75007/_1__syn_2  ;
	output \g75568/_1_  ;
	output \g75792/_0_  ;
	output \g75836/_0_  ;
	output \g76027/_0_  ;
	output \g76034/_0_  ;
	output \g76108/_0_  ;
	output \g76130/_0_  ;
	output \g76266/_0_  ;
	output \g76315/_0_  ;
	output \g76569/_0_  ;
	output \g76714/_0_  ;
	output \g77122/_1__syn_2  ;
	output \g77709/_1_  ;
	output \g81909/_0_  ;
	output \g81922/_0_  ;
	output \g81926/_1__syn_2  ;
	output \g82197/_1_  ;
	output \g82272/_0_  ;
	output \g82291/_0_  ;
	output \g82716/_0_  ;
	output \g82718/_0_  ;
	output \g82738/_0_  ;
	output \g82769/_0_  ;
	output \g82775/_0_  ;
	output \g82779/_1__syn_2  ;
	output \g82804/_0_  ;
	output \g82810/_0_  ;
	output \g82817/_0_  ;
	output \g82823/_0_  ;
	output \g82835/_0_  ;
	output \g82841/_0_  ;
	output \g82847/_0_  ;
	output \g82853/_0_  ;
	output \g82859/_0_  ;
	output \g82862/_1__syn_2  ;
	output \g82956/_0_  ;
	output \g82959/_1_  ;
	output \g83020/_0_  ;
	output \g83025/_0_  ;
	output \g83078/_0_  ;
	output \g83083/_0_  ;
	output \g83121/_0_  ;
	output \g83135/_0_  ;
	output \g83205/_0_  ;
	output \g83240/_0_  ;
	output \g83509/_1__syn_2  ;
	output \g83769/_0_  ;
	output \h0lock_pad  ;
	output \h1sel_br[7]_pad  ;
	output \h1sel_dma[0]_pad  ;
	output \h1sel_dma[4]_pad  ;
	output \h1sel_dma[7]_pad  ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	LUT3 #(
		.INIT('h10)
	) name0 (
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w2229_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		_w2230_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w2231_
	);
	LUT4 #(
		.INIT('h2000)
	) name3 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w2232_
	);
	LUT4 #(
		.INIT('h8000)
	) name4 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2230_,
		_w2232_,
		_w2233_
	);
	LUT4 #(
		.INIT('h0200)
	) name5 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\ctl_rf_m0end_reg/NET0131 ,
		_w2234_
	);
	LUT4 #(
		.INIT('h0100)
	) name6 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\ctl_rf_m0end_reg/NET0131 ,
		_w2235_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name7 (
		\hwdata[31]_pad ,
		\hwdata[7]_pad ,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\hwdata[23]_pad ,
		_w2234_,
		_w2237_
	);
	LUT4 #(
		.INIT('heee2)
	) name9 (
		\ctl_rf_c1_rf_chsad_reg[7]/NET0131 ,
		_w2233_,
		_w2236_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		_w2239_
	);
	LUT4 #(
		.INIT('h8000)
	) name11 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2232_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name12 (
		\hwdata[17]_pad ,
		\hwdata[9]_pad ,
		_w2234_,
		_w2235_,
		_w2241_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\hwdata[1]_pad ,
		_w2234_,
		_w2242_
	);
	LUT4 #(
		.INIT('heee2)
	) name14 (
		\ctl_rf_c1_rf_chdad_reg[17]/NET0131 ,
		_w2240_,
		_w2241_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('h20)
	) name15 (
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w2244_
	);
	LUT4 #(
		.INIT('h8000)
	) name16 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2232_,
		_w2239_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name17 (
		\ctl_rf_c3_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2245_,
		_w2246_
	);
	LUT3 #(
		.INIT('h40)
	) name18 (
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w2248_
	);
	LUT4 #(
		.INIT('h0200)
	) name20 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w2249_
	);
	LUT4 #(
		.INIT('h8000)
	) name21 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2239_,
		_w2247_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name22 (
		\ctl_rf_c4_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h8000)
	) name23 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2232_,
		_w2239_,
		_w2247_,
		_w2252_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name24 (
		\ctl_rf_c5_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2252_,
		_w2253_
	);
	LUT3 #(
		.INIT('h80)
	) name25 (
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w2254_
	);
	LUT4 #(
		.INIT('h8000)
	) name26 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2239_,
		_w2249_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name27 (
		\ctl_rf_c6_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h8000)
	) name28 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2232_,
		_w2239_,
		_w2254_,
		_w2257_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name29 (
		\ctl_rf_c7_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h8000)
	) name30 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w2230_,
		_w2232_,
		_w2259_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name31 (
		\hwdata[31]_pad ,
		\hwdata[7]_pad ,
		_w2234_,
		_w2235_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\hwdata[15]_pad ,
		_w2234_,
		_w2261_
	);
	LUT4 #(
		.INIT('heee2)
	) name33 (
		\ctl_rf_c1_rf_chsad_reg[31]/NET0131 ,
		_w2259_,
		_w2260_,
		_w2261_,
		_w2262_
	);
	LUT4 #(
		.INIT('h8000)
	) name34 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2232_,
		_w2244_,
		_w2263_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name35 (
		\ctl_rf_c3_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2247_,
		_w2249_,
		_w2265_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name37 (
		\ctl_rf_c4_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h8000)
	) name38 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2249_,
		_w2254_,
		_w2267_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name39 (
		\ctl_rf_c6_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2267_,
		_w2268_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w2230_,
		_w2249_,
		_w2269_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name41 (
		\ctl_rf_c0_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h8000)
	) name42 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2239_,
		_w2244_,
		_w2249_,
		_w2271_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name43 (
		\ctl_rf_c2_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2271_,
		_w2272_
	);
	LUT4 #(
		.INIT('h8000)
	) name44 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2244_,
		_w2249_,
		_w2273_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name45 (
		\ctl_rf_c2_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2273_,
		_w2274_
	);
	LUT4 #(
		.INIT('h8000)
	) name46 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2232_,
		_w2247_,
		_w2275_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name47 (
		\ctl_rf_c5_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2275_,
		_w2276_
	);
	LUT4 #(
		.INIT('h8000)
	) name48 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2230_,
		_w2232_,
		_w2254_,
		_w2277_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name49 (
		\ctl_rf_c7_rf_chsad_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('h8000)
	) name50 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2239_,
		_w2249_,
		_w2279_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name51 (
		\ctl_rf_c0_rf_chdad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2279_,
		_w2280_
	);
	LUT4 #(
		.INIT('h8000)
	) name52 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2230_,
		_w2232_,
		_w2281_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name53 (
		\hwdata[13]_pad ,
		\hwdata[21]_pad ,
		_w2234_,
		_w2235_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\hwdata[5]_pad ,
		_w2234_,
		_w2283_
	);
	LUT4 #(
		.INIT('heee2)
	) name55 (
		\ctl_rf_c1_rf_chsad_reg[21]/NET0131 ,
		_w2281_,
		_w2282_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h8000)
	) name56 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2232_,
		_w2244_,
		_w2285_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name57 (
		\ctl_rf_c3_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2285_,
		_w2286_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2247_,
		_w2249_,
		_w2287_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name59 (
		\ctl_rf_c4_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2287_,
		_w2288_
	);
	LUT4 #(
		.INIT('h8000)
	) name60 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2232_,
		_w2247_,
		_w2289_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name61 (
		\ctl_rf_c5_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h8000)
	) name62 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2249_,
		_w2254_,
		_w2291_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name63 (
		\ctl_rf_c6_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h8000)
	) name64 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2232_,
		_w2254_,
		_w2293_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name65 (
		\ctl_rf_c7_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2293_,
		_w2294_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name66 (
		\hwdata[10]_pad ,
		\hwdata[18]_pad ,
		_w2234_,
		_w2235_,
		_w2295_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\hwdata[2]_pad ,
		_w2234_,
		_w2296_
	);
	LUT4 #(
		.INIT('heee2)
	) name68 (
		\ctl_rf_c1_rf_chdad_reg[18]/NET0131 ,
		_w2240_,
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name69 (
		\hwdata[11]_pad ,
		\hwdata[19]_pad ,
		_w2234_,
		_w2235_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\hwdata[3]_pad ,
		_w2234_,
		_w2299_
	);
	LUT4 #(
		.INIT('heee2)
	) name71 (
		\ctl_rf_c1_rf_chdad_reg[19]/NET0131 ,
		_w2240_,
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('heee2)
	) name72 (
		\ctl_rf_c3_rf_chdad_reg[18]/NET0131 ,
		_w2245_,
		_w2295_,
		_w2296_,
		_w2301_
	);
	LUT4 #(
		.INIT('heee2)
	) name73 (
		\ctl_rf_c3_rf_chdad_reg[19]/NET0131 ,
		_w2245_,
		_w2298_,
		_w2299_,
		_w2302_
	);
	LUT4 #(
		.INIT('heee2)
	) name74 (
		\ctl_rf_c3_rf_chsad_reg[18]/NET0131 ,
		_w2285_,
		_w2295_,
		_w2296_,
		_w2303_
	);
	LUT4 #(
		.INIT('heee2)
	) name75 (
		\ctl_rf_c3_rf_chsad_reg[19]/NET0131 ,
		_w2285_,
		_w2298_,
		_w2299_,
		_w2304_
	);
	LUT4 #(
		.INIT('heee2)
	) name76 (
		\ctl_rf_c4_rf_chdad_reg[19]/NET0131 ,
		_w2250_,
		_w2298_,
		_w2299_,
		_w2305_
	);
	LUT4 #(
		.INIT('heee2)
	) name77 (
		\ctl_rf_c4_rf_chdad_reg[18]/NET0131 ,
		_w2250_,
		_w2295_,
		_w2296_,
		_w2306_
	);
	LUT4 #(
		.INIT('heee2)
	) name78 (
		\ctl_rf_c4_rf_chsad_reg[18]/NET0131 ,
		_w2287_,
		_w2295_,
		_w2296_,
		_w2307_
	);
	LUT4 #(
		.INIT('heee2)
	) name79 (
		\ctl_rf_c4_rf_chsad_reg[19]/NET0131 ,
		_w2287_,
		_w2298_,
		_w2299_,
		_w2308_
	);
	LUT4 #(
		.INIT('heee2)
	) name80 (
		\ctl_rf_c5_rf_chdad_reg[18]/NET0131 ,
		_w2252_,
		_w2295_,
		_w2296_,
		_w2309_
	);
	LUT4 #(
		.INIT('heee2)
	) name81 (
		\ctl_rf_c5_rf_chdad_reg[19]/NET0131 ,
		_w2252_,
		_w2298_,
		_w2299_,
		_w2310_
	);
	LUT4 #(
		.INIT('heee2)
	) name82 (
		\ctl_rf_c5_rf_chsad_reg[18]/NET0131 ,
		_w2289_,
		_w2295_,
		_w2296_,
		_w2311_
	);
	LUT4 #(
		.INIT('heee2)
	) name83 (
		\ctl_rf_c5_rf_chsad_reg[19]/NET0131 ,
		_w2289_,
		_w2298_,
		_w2299_,
		_w2312_
	);
	LUT4 #(
		.INIT('heee2)
	) name84 (
		\ctl_rf_c6_rf_chdad_reg[18]/NET0131 ,
		_w2255_,
		_w2295_,
		_w2296_,
		_w2313_
	);
	LUT4 #(
		.INIT('heee2)
	) name85 (
		\ctl_rf_c6_rf_chdad_reg[19]/NET0131 ,
		_w2255_,
		_w2298_,
		_w2299_,
		_w2314_
	);
	LUT4 #(
		.INIT('heee2)
	) name86 (
		\ctl_rf_c6_rf_chsad_reg[18]/NET0131 ,
		_w2291_,
		_w2295_,
		_w2296_,
		_w2315_
	);
	LUT4 #(
		.INIT('heee2)
	) name87 (
		\ctl_rf_c6_rf_chsad_reg[19]/NET0131 ,
		_w2291_,
		_w2298_,
		_w2299_,
		_w2316_
	);
	LUT4 #(
		.INIT('heee2)
	) name88 (
		\ctl_rf_c7_rf_chsad_reg[18]/NET0131 ,
		_w2293_,
		_w2295_,
		_w2296_,
		_w2317_
	);
	LUT4 #(
		.INIT('heee2)
	) name89 (
		\ctl_rf_c7_rf_chsad_reg[19]/NET0131 ,
		_w2293_,
		_w2298_,
		_w2299_,
		_w2318_
	);
	LUT4 #(
		.INIT('h8000)
	) name90 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2230_,
		_w2249_,
		_w2319_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name91 (
		\ctl_rf_c0_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2319_,
		_w2320_
	);
	LUT4 #(
		.INIT('h8000)
	) name92 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2244_,
		_w2249_,
		_w2321_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name93 (
		\ctl_rf_c2_rf_chsad_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w2321_,
		_w2322_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name94 (
		\hwdata[14]_pad ,
		\hwdata[22]_pad ,
		_w2234_,
		_w2235_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\hwdata[6]_pad ,
		_w2234_,
		_w2324_
	);
	LUT4 #(
		.INIT('heee2)
	) name96 (
		\ctl_rf_c1_rf_chsad_reg[22]/NET0131 ,
		_w2281_,
		_w2323_,
		_w2324_,
		_w2325_
	);
	LUT4 #(
		.INIT('heee2)
	) name97 (
		\ctl_rf_c3_rf_chsad_reg[22]/NET0131 ,
		_w2285_,
		_w2323_,
		_w2324_,
		_w2326_
	);
	LUT4 #(
		.INIT('heee2)
	) name98 (
		\ctl_rf_c4_rf_chsad_reg[22]/NET0131 ,
		_w2287_,
		_w2323_,
		_w2324_,
		_w2327_
	);
	LUT4 #(
		.INIT('heee2)
	) name99 (
		\ctl_rf_c5_rf_chsad_reg[22]/NET0131 ,
		_w2289_,
		_w2323_,
		_w2324_,
		_w2328_
	);
	LUT4 #(
		.INIT('heee2)
	) name100 (
		\ctl_rf_c6_rf_chsad_reg[22]/NET0131 ,
		_w2291_,
		_w2323_,
		_w2324_,
		_w2329_
	);
	LUT4 #(
		.INIT('heee2)
	) name101 (
		\ctl_rf_c7_rf_chsad_reg[22]/NET0131 ,
		_w2293_,
		_w2323_,
		_w2324_,
		_w2330_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name102 (
		\hwdata[15]_pad ,
		\hwdata[23]_pad ,
		_w2234_,
		_w2235_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\hwdata[7]_pad ,
		_w2234_,
		_w2332_
	);
	LUT4 #(
		.INIT('heee2)
	) name104 (
		\ctl_rf_c1_rf_chsad_reg[23]/NET0131 ,
		_w2281_,
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT4 #(
		.INIT('heee2)
	) name105 (
		\ctl_rf_c3_rf_chsad_reg[23]/NET0131 ,
		_w2285_,
		_w2331_,
		_w2332_,
		_w2334_
	);
	LUT4 #(
		.INIT('heee2)
	) name106 (
		\ctl_rf_c4_rf_chsad_reg[23]/NET0131 ,
		_w2287_,
		_w2331_,
		_w2332_,
		_w2335_
	);
	LUT4 #(
		.INIT('heee2)
	) name107 (
		\ctl_rf_c5_rf_chsad_reg[23]/NET0131 ,
		_w2289_,
		_w2331_,
		_w2332_,
		_w2336_
	);
	LUT4 #(
		.INIT('heee2)
	) name108 (
		\ctl_rf_c6_rf_chsad_reg[23]/NET0131 ,
		_w2291_,
		_w2331_,
		_w2332_,
		_w2337_
	);
	LUT4 #(
		.INIT('heee2)
	) name109 (
		\ctl_rf_c7_rf_chsad_reg[23]/NET0131 ,
		_w2293_,
		_w2331_,
		_w2332_,
		_w2338_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name110 (
		\ctl_rf_c0_rf_chsad_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w2319_,
		_w2339_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name111 (
		\ctl_rf_c0_rf_chsad_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w2319_,
		_w2340_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name112 (
		\hwdata[12]_pad ,
		\hwdata[20]_pad ,
		_w2234_,
		_w2235_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\hwdata[4]_pad ,
		_w2234_,
		_w2342_
	);
	LUT4 #(
		.INIT('heee2)
	) name114 (
		\ctl_rf_c1_rf_chsad_reg[20]/NET0131 ,
		_w2281_,
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name115 (
		\hwdata[0]_pad ,
		\hwdata[24]_pad ,
		_w2234_,
		_w2235_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\hwdata[8]_pad ,
		_w2234_,
		_w2345_
	);
	LUT4 #(
		.INIT('heee2)
	) name117 (
		\ctl_rf_c1_rf_chsad_reg[24]/NET0131 ,
		_w2259_,
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT4 #(
		.INIT('heee2)
	) name118 (
		\ctl_rf_c2_rf_chdad_reg[18]/NET0131 ,
		_w2271_,
		_w2295_,
		_w2296_,
		_w2347_
	);
	LUT4 #(
		.INIT('heee2)
	) name119 (
		\ctl_rf_c2_rf_chdad_reg[19]/NET0131 ,
		_w2271_,
		_w2298_,
		_w2299_,
		_w2348_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name120 (
		\ctl_rf_c2_rf_chsad_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w2321_,
		_w2349_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name121 (
		\ctl_rf_c2_rf_chsad_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w2321_,
		_w2350_
	);
	LUT4 #(
		.INIT('heee2)
	) name122 (
		\ctl_rf_c3_rf_chsad_reg[20]/NET0131 ,
		_w2285_,
		_w2341_,
		_w2342_,
		_w2351_
	);
	LUT4 #(
		.INIT('heee2)
	) name123 (
		\ctl_rf_c3_rf_chsad_reg[24]/NET0131 ,
		_w2263_,
		_w2344_,
		_w2345_,
		_w2352_
	);
	LUT4 #(
		.INIT('heee2)
	) name124 (
		\ctl_rf_c4_rf_chsad_reg[20]/NET0131 ,
		_w2287_,
		_w2341_,
		_w2342_,
		_w2353_
	);
	LUT4 #(
		.INIT('heee2)
	) name125 (
		\ctl_rf_c4_rf_chsad_reg[24]/NET0131 ,
		_w2265_,
		_w2344_,
		_w2345_,
		_w2354_
	);
	LUT4 #(
		.INIT('heee2)
	) name126 (
		\ctl_rf_c6_rf_chsad_reg[20]/NET0131 ,
		_w2291_,
		_w2341_,
		_w2342_,
		_w2355_
	);
	LUT4 #(
		.INIT('heee2)
	) name127 (
		\ctl_rf_c6_rf_chsad_reg[24]/NET0131 ,
		_w2267_,
		_w2344_,
		_w2345_,
		_w2356_
	);
	LUT4 #(
		.INIT('heee2)
	) name128 (
		\ctl_rf_c0_rf_chdad_reg[18]/NET0131 ,
		_w2279_,
		_w2295_,
		_w2296_,
		_w2357_
	);
	LUT4 #(
		.INIT('heee2)
	) name129 (
		\ctl_rf_c0_rf_chdad_reg[19]/NET0131 ,
		_w2279_,
		_w2298_,
		_w2299_,
		_w2358_
	);
	LUT4 #(
		.INIT('heee2)
	) name130 (
		\ctl_rf_c0_rf_chsad_reg[20]/NET0131 ,
		_w2319_,
		_w2341_,
		_w2342_,
		_w2359_
	);
	LUT4 #(
		.INIT('heee2)
	) name131 (
		\ctl_rf_c0_rf_chsad_reg[22]/NET0131 ,
		_w2319_,
		_w2323_,
		_w2324_,
		_w2360_
	);
	LUT4 #(
		.INIT('heee2)
	) name132 (
		\ctl_rf_c0_rf_chsad_reg[23]/NET0131 ,
		_w2319_,
		_w2331_,
		_w2332_,
		_w2361_
	);
	LUT4 #(
		.INIT('heee2)
	) name133 (
		\ctl_rf_c0_rf_chsad_reg[24]/NET0131 ,
		_w2269_,
		_w2344_,
		_w2345_,
		_w2362_
	);
	LUT4 #(
		.INIT('heee2)
	) name134 (
		\ctl_rf_c2_rf_chsad_reg[20]/NET0131 ,
		_w2321_,
		_w2341_,
		_w2342_,
		_w2363_
	);
	LUT4 #(
		.INIT('heee2)
	) name135 (
		\ctl_rf_c2_rf_chsad_reg[22]/NET0131 ,
		_w2321_,
		_w2323_,
		_w2324_,
		_w2364_
	);
	LUT4 #(
		.INIT('heee2)
	) name136 (
		\ctl_rf_c2_rf_chsad_reg[23]/NET0131 ,
		_w2321_,
		_w2331_,
		_w2332_,
		_w2365_
	);
	LUT4 #(
		.INIT('heee2)
	) name137 (
		\ctl_rf_c2_rf_chsad_reg[24]/NET0131 ,
		_w2273_,
		_w2344_,
		_w2345_,
		_w2366_
	);
	LUT4 #(
		.INIT('heee2)
	) name138 (
		\ctl_rf_c5_rf_chsad_reg[20]/NET0131 ,
		_w2289_,
		_w2341_,
		_w2342_,
		_w2367_
	);
	LUT4 #(
		.INIT('heee2)
	) name139 (
		\ctl_rf_c5_rf_chsad_reg[24]/NET0131 ,
		_w2275_,
		_w2344_,
		_w2345_,
		_w2368_
	);
	LUT4 #(
		.INIT('heee2)
	) name140 (
		\ctl_rf_c7_rf_chsad_reg[20]/NET0131 ,
		_w2293_,
		_w2341_,
		_w2342_,
		_w2369_
	);
	LUT4 #(
		.INIT('heee2)
	) name141 (
		\ctl_rf_c7_rf_chsad_reg[24]/NET0131 ,
		_w2277_,
		_w2344_,
		_w2345_,
		_w2370_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name142 (
		\hwdata[16]_pad ,
		\hwdata[8]_pad ,
		_w2234_,
		_w2235_,
		_w2371_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\hwdata[0]_pad ,
		_w2234_,
		_w2372_
	);
	LUT4 #(
		.INIT('heee2)
	) name144 (
		\ctl_rf_c1_rf_chsad_reg[16]/NET0131 ,
		_w2281_,
		_w2371_,
		_w2372_,
		_w2373_
	);
	LUT4 #(
		.INIT('heee2)
	) name145 (
		\ctl_rf_c3_rf_chsad_reg[16]/NET0131 ,
		_w2285_,
		_w2371_,
		_w2372_,
		_w2374_
	);
	LUT4 #(
		.INIT('heee2)
	) name146 (
		\ctl_rf_c4_rf_chdad_reg[16]/NET0131 ,
		_w2250_,
		_w2371_,
		_w2372_,
		_w2375_
	);
	LUT4 #(
		.INIT('heee2)
	) name147 (
		\ctl_rf_c4_rf_chsad_reg[16]/NET0131 ,
		_w2287_,
		_w2371_,
		_w2372_,
		_w2376_
	);
	LUT4 #(
		.INIT('heee2)
	) name148 (
		\ctl_rf_c6_rf_chdad_reg[16]/NET0131 ,
		_w2255_,
		_w2371_,
		_w2372_,
		_w2377_
	);
	LUT4 #(
		.INIT('heee2)
	) name149 (
		\ctl_rf_c6_rf_chsad_reg[16]/NET0131 ,
		_w2291_,
		_w2371_,
		_w2372_,
		_w2378_
	);
	LUT4 #(
		.INIT('heee2)
	) name150 (
		\ctl_rf_c0_rf_chsad_reg[16]/NET0131 ,
		_w2319_,
		_w2371_,
		_w2372_,
		_w2379_
	);
	LUT4 #(
		.INIT('heee2)
	) name151 (
		\ctl_rf_c1_rf_chdad_reg[16]/NET0131 ,
		_w2240_,
		_w2371_,
		_w2372_,
		_w2380_
	);
	LUT4 #(
		.INIT('heee2)
	) name152 (
		\ctl_rf_c2_rf_chdad_reg[16]/NET0131 ,
		_w2271_,
		_w2371_,
		_w2372_,
		_w2381_
	);
	LUT4 #(
		.INIT('heee2)
	) name153 (
		\ctl_rf_c2_rf_chsad_reg[16]/NET0131 ,
		_w2321_,
		_w2371_,
		_w2372_,
		_w2382_
	);
	LUT4 #(
		.INIT('heee2)
	) name154 (
		\ctl_rf_c3_rf_chdad_reg[16]/NET0131 ,
		_w2245_,
		_w2371_,
		_w2372_,
		_w2383_
	);
	LUT4 #(
		.INIT('heee2)
	) name155 (
		\ctl_rf_c5_rf_chdad_reg[16]/NET0131 ,
		_w2252_,
		_w2371_,
		_w2372_,
		_w2384_
	);
	LUT4 #(
		.INIT('heee2)
	) name156 (
		\ctl_rf_c5_rf_chsad_reg[16]/NET0131 ,
		_w2289_,
		_w2371_,
		_w2372_,
		_w2385_
	);
	LUT4 #(
		.INIT('heee2)
	) name157 (
		\ctl_rf_c7_rf_chdad_reg[16]/NET0131 ,
		_w2257_,
		_w2371_,
		_w2372_,
		_w2386_
	);
	LUT4 #(
		.INIT('heee2)
	) name158 (
		\ctl_rf_c7_rf_chsad_reg[16]/NET0131 ,
		_w2293_,
		_w2371_,
		_w2372_,
		_w2387_
	);
	LUT4 #(
		.INIT('heee2)
	) name159 (
		\ctl_rf_c0_rf_chdad_reg[16]/NET0131 ,
		_w2279_,
		_w2371_,
		_w2372_,
		_w2388_
	);
	LUT4 #(
		.INIT('h0400)
	) name160 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2389_
	);
	LUT3 #(
		.INIT('h13)
	) name161 (
		\h1rdy2_br_pad ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h8000)
	) name162 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2391_
	);
	LUT4 #(
		.INIT('h4000)
	) name163 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2392_
	);
	LUT4 #(
		.INIT('h153f)
	) name164 (
		\h1rdy6_br_pad ,
		\h1rdy7_br_pad ,
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h0008)
	) name165 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2394_
	);
	LUT4 #(
		.INIT('h0002)
	) name166 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2395_
	);
	LUT4 #(
		.INIT('h153f)
	) name167 (
		\h1rdy1_dma_pad ,
		\h1rdy3_dma_pad ,
		_w2394_,
		_w2395_,
		_w2396_
	);
	LUT3 #(
		.INIT('h80)
	) name168 (
		_w2390_,
		_w2393_,
		_w2396_,
		_w2397_
	);
	LUT4 #(
		.INIT('h0800)
	) name169 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\h1rdy3_br_pad ,
		_w2398_,
		_w2399_
	);
	LUT4 #(
		.INIT('h0200)
	) name171 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2400_
	);
	LUT4 #(
		.INIT('h0020)
	) name172 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2401_
	);
	LUT4 #(
		.INIT('h135f)
	) name173 (
		\h1rdy1_br_pad ,
		\h1rdy5_dma_pad ,
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w2399_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h0080)
	) name175 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2404_
	);
	LUT4 #(
		.INIT('h1000)
	) name176 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2405_
	);
	LUT4 #(
		.INIT('h153f)
	) name177 (
		\h1rdy4_br_pad ,
		\h1rdy7_dma_pad ,
		_w2404_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('h0100)
	) name178 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2407_
	);
	LUT4 #(
		.INIT('h2000)
	) name179 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2408_
	);
	LUT4 #(
		.INIT('h135f)
	) name180 (
		\h1rdy0_br_pad ,
		\h1rdy5_br_pad ,
		_w2407_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h0004)
	) name181 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2410_
	);
	LUT4 #(
		.INIT('h0010)
	) name182 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2411_
	);
	LUT4 #(
		.INIT('h135f)
	) name183 (
		\h1rdy2_dma_pad ,
		\h1rdy4_dma_pad ,
		_w2410_,
		_w2411_,
		_w2412_
	);
	LUT4 #(
		.INIT('h0040)
	) name184 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2413_
	);
	LUT4 #(
		.INIT('h0001)
	) name185 (
		\m1_mux_mux_no_reg[0]/NET0131 ,
		\m1_mux_mux_no_reg[1]/NET0131 ,
		\m1_mux_mux_no_reg[2]/NET0131 ,
		\m1_mux_mux_no_reg[3]/NET0131 ,
		_w2414_
	);
	LUT4 #(
		.INIT('h153f)
	) name186 (
		\h1rdy0_dma_pad ,
		\h1rdy6_dma_pad ,
		_w2413_,
		_w2414_,
		_w2415_
	);
	LUT4 #(
		.INIT('h8000)
	) name187 (
		_w2406_,
		_w2409_,
		_w2412_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h80)
	) name188 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w2417_
	);
	LUT3 #(
		.INIT('h10)
	) name189 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		_w2418_
	);
	LUT4 #(
		.INIT('h0010)
	) name190 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2419_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\de_tsz_cnt_reg[10]/NET0131 ,
		\de_tsz_cnt_reg[11]/NET0131 ,
		_w2420_
	);
	LUT4 #(
		.INIT('h0001)
	) name192 (
		\de_tsz_cnt_reg[2]/NET0131 ,
		\de_tsz_cnt_reg[3]/NET0131 ,
		\de_tsz_cnt_reg[4]/NET0131 ,
		\de_tsz_cnt_reg[5]/NET0131 ,
		_w2421_
	);
	LUT4 #(
		.INIT('h0001)
	) name193 (
		\de_tsz_cnt_reg[6]/NET0131 ,
		\de_tsz_cnt_reg[7]/NET0131 ,
		\de_tsz_cnt_reg[8]/NET0131 ,
		\de_tsz_cnt_reg[9]/NET0131 ,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\de_tsz_cnt_reg[0]/NET0131 ,
		\de_tsz_cnt_reg[1]/NET0131 ,
		_w2423_
	);
	LUT4 #(
		.INIT('h8000)
	) name195 (
		_w2420_,
		_w2421_,
		_w2422_,
		_w2423_,
		_w2424_
	);
	LUT3 #(
		.INIT('ha8)
	) name196 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w2425_
	);
	LUT4 #(
		.INIT('h0001)
	) name197 (
		\de_bst_cnt_reg[5]/NET0131 ,
		\de_bst_cnt_reg[6]/NET0131 ,
		\de_bst_cnt_reg[7]/NET0131 ,
		\de_bst_cnt_reg[8]/NET0131 ,
		_w2426_
	);
	LUT4 #(
		.INIT('h0001)
	) name198 (
		\de_bst_cnt_reg[0]/NET0131 ,
		\de_bst_cnt_reg[2]/NET0131 ,
		\de_bst_cnt_reg[3]/NET0131 ,
		\de_bst_cnt_reg[4]/NET0131 ,
		_w2427_
	);
	LUT3 #(
		.INIT('h2a)
	) name199 (
		_w2425_,
		_w2426_,
		_w2427_,
		_w2428_
	);
	LUT4 #(
		.INIT('h135f)
	) name200 (
		\ahb_slv_slv_br_req_reg/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w2429_
	);
	LUT4 #(
		.INIT('h1055)
	) name201 (
		_w2419_,
		_w2424_,
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2431_
	);
	LUT3 #(
		.INIT('h01)
	) name203 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w2432_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w2431_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w2430_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		_w2417_,
		_w2434_,
		_w2435_
	);
	LUT4 #(
		.INIT('h0e00)
	) name207 (
		\ch_sel_arb_chcsr_reg_reg[3]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[4]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m1_arb_st_reg[0]/NET0131 ,
		_w2436_
	);
	LUT4 #(
		.INIT('h000e)
	) name208 (
		\ch_sel_arb_chcsr_reg_reg[5]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[6]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m1_arb_st_reg[0]/NET0131 ,
		_w2437_
	);
	LUT3 #(
		.INIT('h01)
	) name209 (
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2436_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('hba8a)
	) name210 (
		\h1burst[0]_pad ,
		_w2417_,
		_w2434_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		_w2440_
	);
	LUT3 #(
		.INIT('h40)
	) name212 (
		_w2417_,
		_w2434_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\m1_mux_hrmxnof_reg/NET0131 ,
		\m1_mux_hrp_df_reg[0]/NET0131 ,
		_w2442_
	);
	LUT3 #(
		.INIT('h13)
	) name214 (
		\h1rp0_br[0]_pad ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2407_,
		_w2443_
	);
	LUT4 #(
		.INIT('h153f)
	) name215 (
		\h1rp0_dma[0]_pad ,
		\h1rp4_dma[0]_pad ,
		_w2411_,
		_w2414_,
		_w2444_
	);
	LUT4 #(
		.INIT('h135f)
	) name216 (
		\h1rp2_br[0]_pad ,
		\h1rp2_dma[0]_pad ,
		_w2389_,
		_w2410_,
		_w2445_
	);
	LUT3 #(
		.INIT('h80)
	) name217 (
		_w2443_,
		_w2444_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\h1rp4_br[0]_pad ,
		_w2405_,
		_w2447_
	);
	LUT4 #(
		.INIT('h153f)
	) name219 (
		\h1rp1_br[0]_pad ,
		\h1rp3_br[0]_pad ,
		_w2398_,
		_w2400_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		_w2447_,
		_w2448_,
		_w2449_
	);
	LUT4 #(
		.INIT('h153f)
	) name221 (
		\h1rp1_dma[0]_pad ,
		\h1rp3_dma[0]_pad ,
		_w2394_,
		_w2395_,
		_w2450_
	);
	LUT4 #(
		.INIT('h153f)
	) name222 (
		\h1rp5_dma[0]_pad ,
		\h1rp6_br[0]_pad ,
		_w2392_,
		_w2401_,
		_w2451_
	);
	LUT4 #(
		.INIT('h153f)
	) name223 (
		\h1rp5_br[0]_pad ,
		\h1rp7_br[0]_pad ,
		_w2391_,
		_w2408_,
		_w2452_
	);
	LUT4 #(
		.INIT('h153f)
	) name224 (
		\h1rp6_dma[0]_pad ,
		\h1rp7_dma[0]_pad ,
		_w2404_,
		_w2413_,
		_w2453_
	);
	LUT4 #(
		.INIT('h8000)
	) name225 (
		_w2450_,
		_w2451_,
		_w2452_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('h1555)
	) name226 (
		_w2442_,
		_w2446_,
		_w2449_,
		_w2454_,
		_w2455_
	);
	LUT4 #(
		.INIT('h153f)
	) name227 (
		\h1rp0_dma[1]_pad ,
		\h1rp5_dma[1]_pad ,
		_w2401_,
		_w2414_,
		_w2456_
	);
	LUT4 #(
		.INIT('h135f)
	) name228 (
		\h1rp6_br[1]_pad ,
		\h1rp6_dma[1]_pad ,
		_w2392_,
		_w2413_,
		_w2457_
	);
	LUT4 #(
		.INIT('h153f)
	) name229 (
		\h1rp0_br[1]_pad ,
		\h1rp1_dma[1]_pad ,
		_w2395_,
		_w2407_,
		_w2458_
	);
	LUT4 #(
		.INIT('h153f)
	) name230 (
		\h1rp5_br[1]_pad ,
		\h1rp7_dma[1]_pad ,
		_w2404_,
		_w2408_,
		_w2459_
	);
	LUT4 #(
		.INIT('h8000)
	) name231 (
		_w2456_,
		_w2457_,
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT4 #(
		.INIT('h153f)
	) name232 (
		\h1rp1_br[1]_pad ,
		\h1rp7_br[1]_pad ,
		_w2391_,
		_w2400_,
		_w2461_
	);
	LUT4 #(
		.INIT('h135f)
	) name233 (
		\h1rp4_br[1]_pad ,
		\h1rp4_dma[1]_pad ,
		_w2405_,
		_w2411_,
		_w2462_
	);
	LUT4 #(
		.INIT('h153f)
	) name234 (
		\h1rp3_br[1]_pad ,
		\h1rp3_dma[1]_pad ,
		_w2394_,
		_w2398_,
		_w2463_
	);
	LUT4 #(
		.INIT('h135f)
	) name235 (
		\h1rp2_br[1]_pad ,
		\h1rp2_dma[1]_pad ,
		_w2389_,
		_w2410_,
		_w2464_
	);
	LUT4 #(
		.INIT('h8000)
	) name236 (
		_w2461_,
		_w2462_,
		_w2463_,
		_w2464_,
		_w2465_
	);
	LUT3 #(
		.INIT('h15)
	) name237 (
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2460_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\de_m1_arb_st_reg[0]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2467_
	);
	LUT3 #(
		.INIT('h02)
	) name239 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_m1_arb_st_reg[0]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2468_
	);
	LUT3 #(
		.INIT('h54)
	) name240 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[5]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[6]/NET0131 ,
		_w2469_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		\de_tsz_cnt_reg[0]/NET0131 ,
		\de_tsz_cnt_reg[1]/NET0131 ,
		_w2470_
	);
	LUT4 #(
		.INIT('h8000)
	) name242 (
		_w2420_,
		_w2421_,
		_w2422_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		\de_m1_arb_st_reg[0]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2472_
	);
	LUT4 #(
		.INIT('h4440)
	) name244 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[3]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[4]/NET0131 ,
		_w2473_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		_w2474_
	);
	LUT3 #(
		.INIT('h70)
	) name246 (
		_w2472_,
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT4 #(
		.INIT('h5700)
	) name247 (
		_w2468_,
		_w2469_,
		_w2471_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('hea00)
	) name248 (
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2460_,
		_w2465_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w2455_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('he)
	) name250 (
		_w2441_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst0_mx_dtp_reg/NET0131 ,
		_w2480_
	);
	LUT3 #(
		.INIT('h40)
	) name252 (
		\de_de_st_reg[5]/NET0131 ,
		\h0grant_pad ,
		\h0readyin_pad ,
		_w2481_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('h15)
	) name254 (
		\h0burst[0]_pad ,
		_w2480_,
		_w2481_,
		_w2483_
	);
	LUT3 #(
		.INIT('h54)
	) name255 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w2484_
	);
	LUT3 #(
		.INIT('h70)
	) name256 (
		_w2426_,
		_w2427_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w2486_
	);
	LUT3 #(
		.INIT('h07)
	) name258 (
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		\h0burst[0]_pad ,
		_w2487_
	);
	LUT4 #(
		.INIT('h1033)
	) name259 (
		_w2424_,
		_w2483_,
		_w2485_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('h0e00)
	) name260 (
		\ch_sel_arb_chcsr_reg_reg[3]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[4]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w2489_
	);
	LUT4 #(
		.INIT('h000e)
	) name261 (
		\ch_sel_arb_chcsr_reg_reg[5]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[6]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w2490_
	);
	LUT4 #(
		.INIT('h8880)
	) name262 (
		_w2480_,
		_w2481_,
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('hf400)
	) name263 (
		_w2424_,
		_w2485_,
		_w2486_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		_w2488_,
		_w2492_,
		_w2493_
	);
	LUT4 #(
		.INIT('h7770)
	) name265 (
		\ahb_mst0_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[5]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[6]/NET0131 ,
		_w2494_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w2495_
	);
	LUT3 #(
		.INIT('he0)
	) name267 (
		\ch_sel_arb_chcsr_reg_reg[3]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[4]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\ahb_mst0_mx_cmd_st_reg[0]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		_w2497_
	);
	LUT4 #(
		.INIT('h0008)
	) name269 (
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\h0grant_pad ,
		\h0resp[0]_pad ,
		\h0resp[1]_pad ,
		_w2498_
	);
	LUT3 #(
		.INIT('h70)
	) name270 (
		_w2496_,
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h1f00)
	) name271 (
		_w2471_,
		_w2494_,
		_w2495_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h40)
	) name272 (
		\ahb_mst0_mx_cmd_st_reg[0]/NET0131 ,
		_w2480_,
		_w2481_,
		_w2501_
	);
	LUT4 #(
		.INIT('hf400)
	) name273 (
		_w2424_,
		_w2485_,
		_w2486_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('he)
	) name274 (
		_w2500_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2504_
	);
	LUT3 #(
		.INIT('h20)
	) name276 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2505_
	);
	LUT4 #(
		.INIT('h0200)
	) name277 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_c4_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2506_
	);
	LUT4 #(
		.INIT('hf35f)
	) name278 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2507_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name279 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h7)
	) name281 (
		_w2507_,
		_w2508_,
		_w2510_
	);
	LUT3 #(
		.INIT('h80)
	) name282 (
		\de_de_st_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w2511_
	);
	LUT4 #(
		.INIT('h35ff)
	) name283 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2512_
	);
	LUT4 #(
		.INIT('hff35)
	) name284 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2513_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w2512_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h7)
	) name286 (
		_w2512_,
		_w2513_,
		_w2515_
	);
	LUT4 #(
		.INIT('h35ff)
	) name287 (
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2516_
	);
	LUT4 #(
		.INIT('hff35)
	) name288 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('h7)
	) name290 (
		_w2516_,
		_w2517_,
		_w2519_
	);
	LUT4 #(
		.INIT('h0888)
	) name291 (
		_w2512_,
		_w2513_,
		_w2516_,
		_w2517_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w2511_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('h00ca)
	) name293 (
		\ch_sel_dma_reqd1_reg[4]/NET0131 ,
		\ch_sel_dma_reqd2_reg[4]/NET0131 ,
		\ctl_rf_sync_reg[4]/NET0131 ,
		\dma_ack[4]_pad ,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		_w2505_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h4055)
	) name295 (
		_w2506_,
		_w2511_,
		_w2520_,
		_w2523_,
		_w2524_
	);
	LUT3 #(
		.INIT('h20)
	) name296 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2525_
	);
	LUT4 #(
		.INIT('h0200)
	) name297 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_c6_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2526_
	);
	LUT4 #(
		.INIT('h0777)
	) name298 (
		_w2512_,
		_w2513_,
		_w2516_,
		_w2517_,
		_w2527_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w2511_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h00ca)
	) name300 (
		\ch_sel_dma_reqd1_reg[6]/NET0131 ,
		\ch_sel_dma_reqd2_reg[6]/NET0131 ,
		\ctl_rf_sync_reg[6]/NET0131 ,
		\dma_ack[6]_pad ,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w2525_,
		_w2529_,
		_w2530_
	);
	LUT4 #(
		.INIT('h2033)
	) name302 (
		_w2511_,
		_w2526_,
		_w2527_,
		_w2530_,
		_w2531_
	);
	LUT3 #(
		.INIT('h20)
	) name303 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2532_
	);
	LUT4 #(
		.INIT('h0200)
	) name304 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\ctl_rf_c3_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2533_
	);
	LUT4 #(
		.INIT('h7000)
	) name305 (
		_w2512_,
		_w2513_,
		_w2516_,
		_w2517_,
		_w2534_
	);
	LUT3 #(
		.INIT('h2a)
	) name306 (
		\de_de_st_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w2535_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w2534_,
		_w2535_,
		_w2536_
	);
	LUT4 #(
		.INIT('h00ca)
	) name308 (
		\ch_sel_dma_reqd1_reg[3]/NET0131 ,
		\ch_sel_dma_reqd2_reg[3]/P0001 ,
		\ctl_rf_sync_reg[3]/NET0131 ,
		\dma_ack[3]_pad ,
		_w2537_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w2532_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('h4055)
	) name310 (
		_w2533_,
		_w2534_,
		_w2535_,
		_w2538_,
		_w2539_
	);
	LUT3 #(
		.INIT('h20)
	) name311 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2540_
	);
	LUT4 #(
		.INIT('h0200)
	) name312 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_c5_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2541_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w2520_,
		_w2535_,
		_w2542_
	);
	LUT4 #(
		.INIT('h00ca)
	) name314 (
		\ch_sel_dma_reqd1_reg[5]/NET0131 ,
		\ch_sel_dma_reqd2_reg[5]/NET0131 ,
		\ctl_rf_sync_reg[5]/NET0131 ,
		\dma_ack[5]_pad ,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w2540_,
		_w2543_,
		_w2544_
	);
	LUT4 #(
		.INIT('h080f)
	) name316 (
		_w2520_,
		_w2535_,
		_w2541_,
		_w2544_,
		_w2545_
	);
	LUT4 #(
		.INIT('h8000)
	) name317 (
		_w2524_,
		_w2531_,
		_w2539_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('h20)
	) name318 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2547_
	);
	LUT4 #(
		.INIT('h0200)
	) name319 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_c0_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2548_
	);
	LUT4 #(
		.INIT('h8000)
	) name320 (
		_w2512_,
		_w2513_,
		_w2516_,
		_w2517_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		_w2511_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h00ca)
	) name322 (
		\ch_sel_dma_reqd1_reg[0]/NET0131 ,
		\ch_sel_dma_reqd2_reg[0]/NET0131 ,
		\ctl_rf_sync_reg[0]/NET0131 ,
		\dma_ack[0]_pad ,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		_w2547_,
		_w2551_,
		_w2552_
	);
	LUT4 #(
		.INIT('h2033)
	) name324 (
		_w2511_,
		_w2548_,
		_w2549_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h20)
	) name325 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2554_
	);
	LUT4 #(
		.INIT('h0200)
	) name326 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_c2_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w2511_,
		_w2534_,
		_w2556_
	);
	LUT4 #(
		.INIT('h00ca)
	) name328 (
		\ch_sel_dma_reqd1_reg[2]/NET0131 ,
		\ch_sel_dma_reqd2_reg[2]/P0001 ,
		\ctl_rf_sync_reg[2]/NET0131 ,
		\dma_ack[2]_pad ,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		_w2554_,
		_w2557_,
		_w2558_
	);
	LUT4 #(
		.INIT('h080f)
	) name330 (
		_w2511_,
		_w2534_,
		_w2555_,
		_w2558_,
		_w2559_
	);
	LUT3 #(
		.INIT('h20)
	) name331 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2560_
	);
	LUT4 #(
		.INIT('h0200)
	) name332 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_c1_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w2535_,
		_w2549_,
		_w2562_
	);
	LUT4 #(
		.INIT('h00ca)
	) name334 (
		\ch_sel_dma_reqd1_reg[1]/NET0131 ,
		\ch_sel_dma_reqd2_reg[1]/P0001 ,
		\ctl_rf_sync_reg[1]/NET0131 ,
		\dma_ack[1]_pad ,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w2560_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h080f)
	) name336 (
		_w2535_,
		_w2549_,
		_w2561_,
		_w2564_,
		_w2565_
	);
	LUT3 #(
		.INIT('h20)
	) name337 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2566_
	);
	LUT4 #(
		.INIT('h0200)
	) name338 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\ctl_rf_c7_rf_mode_reg/NET0131 ,
		\ctl_rf_dmacen_reg/NET0131 ,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w2527_,
		_w2535_,
		_w2568_
	);
	LUT4 #(
		.INIT('h00ca)
	) name340 (
		\ch_sel_dma_reqd1_reg[7]/NET0131 ,
		\ch_sel_dma_reqd2_reg[7]/NET0131 ,
		\ctl_rf_sync_reg[7]/NET0131 ,
		\dma_ack[7]_pad ,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w2566_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('h080f)
	) name342 (
		_w2527_,
		_w2535_,
		_w2567_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('h8000)
	) name343 (
		_w2553_,
		_w2559_,
		_w2565_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h7)
	) name344 (
		_w2546_,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\ch_sel_vld_req_any_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2574_
	);
	LUT4 #(
		.INIT('h0001)
	) name346 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2575_
	);
	LUT4 #(
		.INIT('h0001)
	) name347 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2576_
	);
	LUT3 #(
		.INIT('h2a)
	) name348 (
		\de_de_st_reg[0]/NET0131 ,
		_w2575_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('h5111)
	) name349 (
		\ch_sel_de_stup_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2575_,
		_w2576_,
		_w2578_
	);
	LUT4 #(
		.INIT('h8f00)
	) name350 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		_w2504_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2581_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\ctl_rf_c0_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chpri_reg[1]/NET0131 ,
		_w2582_
	);
	LUT4 #(
		.INIT('h2030)
	) name354 (
		_w2553_,
		_w2565_,
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2584_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w2571_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w2583_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\ctl_rf_c3_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chpri_reg[1]/NET0131 ,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		_w2539_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		\ctl_rf_c2_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chpri_reg[1]/NET0131 ,
		_w2589_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w2559_,
		_w2589_,
		_w2590_
	);
	LUT4 #(
		.INIT('h8caf)
	) name362 (
		_w2553_,
		_w2559_,
		_w2582_,
		_w2589_,
		_w2591_
	);
	LUT4 #(
		.INIT('h0111)
	) name363 (
		_w2583_,
		_w2585_,
		_w2588_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\ctl_rf_c4_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chpri_reg[1]/NET0131 ,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w2524_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w2591_,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		_w2596_
	);
	LUT4 #(
		.INIT('h4044)
	) name368 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2504_,
		_w2531_,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('hd0)
	) name369 (
		_w2592_,
		_w2595_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2599_
	);
	LUT3 #(
		.INIT('h04)
	) name371 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2600_
	);
	LUT2 #(
		.INIT('h4)
	) name372 (
		_w2578_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w2574_,
		_w2600_,
		_w2602_
	);
	LUT4 #(
		.INIT('h080f)
	) name374 (
		_w2546_,
		_w2572_,
		_w2601_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2604_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w2545_,
		_w2604_,
		_w2605_
	);
	LUT4 #(
		.INIT('h8caf)
	) name377 (
		_w2539_,
		_w2545_,
		_w2587_,
		_w2604_,
		_w2606_
	);
	LUT3 #(
		.INIT('h10)
	) name378 (
		_w2583_,
		_w2585_,
		_w2606_,
		_w2607_
	);
	LUT4 #(
		.INIT('h4050)
	) name379 (
		_w2531_,
		_w2545_,
		_w2596_,
		_w2604_,
		_w2608_
	);
	LUT3 #(
		.INIT('h54)
	) name380 (
		_w2588_,
		_w2594_,
		_w2608_,
		_w2609_
	);
	LUT3 #(
		.INIT('h01)
	) name381 (
		_w2603_,
		_w2607_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h2300)
	) name382 (
		_w2524_,
		_w2545_,
		_w2593_,
		_w2604_,
		_w2611_
	);
	LUT3 #(
		.INIT('h32)
	) name383 (
		_w2588_,
		_w2590_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('h8acf)
	) name384 (
		_w2531_,
		_w2553_,
		_w2582_,
		_w2596_,
		_w2613_
	);
	LUT4 #(
		.INIT('h2030)
	) name385 (
		_w2531_,
		_w2571_,
		_w2584_,
		_w2596_,
		_w2614_
	);
	LUT4 #(
		.INIT('h8acf)
	) name386 (
		_w2524_,
		_w2559_,
		_w2589_,
		_w2593_,
		_w2615_
	);
	LUT3 #(
		.INIT('he0)
	) name387 (
		_w2613_,
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT3 #(
		.INIT('h02)
	) name388 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2617_
	);
	LUT4 #(
		.INIT('hfe00)
	) name389 (
		_w2579_,
		_w2612_,
		_w2616_,
		_w2617_,
		_w2618_
	);
	LUT4 #(
		.INIT('h0001)
	) name390 (
		_w2580_,
		_w2598_,
		_w2610_,
		_w2618_,
		_w2619_
	);
	LUT3 #(
		.INIT('hc8)
	) name391 (
		_w2588_,
		_w2591_,
		_w2611_,
		_w2620_
	);
	LUT3 #(
		.INIT('ha2)
	) name392 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2586_,
		_w2620_,
		_w2621_
	);
	LUT4 #(
		.INIT('h8acf)
	) name393 (
		_w2545_,
		_w2571_,
		_w2584_,
		_w2604_,
		_w2622_
	);
	LUT4 #(
		.INIT('h1500)
	) name394 (
		_w2583_,
		_w2588_,
		_w2591_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2608_,
		_w2624_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		_w2623_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2626_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w2578_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('h0400)
	) name399 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		\ch_sel_vld_req_any_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2628_
	);
	LUT4 #(
		.INIT('h080f)
	) name400 (
		_w2546_,
		_w2572_,
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT3 #(
		.INIT('h0e)
	) name401 (
		_w2621_,
		_w2625_,
		_w2629_,
		_w2630_
	);
	LUT3 #(
		.INIT('h08)
	) name402 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2631_
	);
	LUT4 #(
		.INIT('h4500)
	) name403 (
		_w2559_,
		_w2565_,
		_w2581_,
		_w2589_,
		_w2632_
	);
	LUT3 #(
		.INIT('h04)
	) name404 (
		_w2594_,
		_w2613_,
		_w2632_,
		_w2633_
	);
	LUT3 #(
		.INIT('h23)
	) name405 (
		_w2594_,
		_w2611_,
		_w2614_,
		_w2634_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name406 (
		_w2579_,
		_w2631_,
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2578_,
		_w2636_
	);
	LUT3 #(
		.INIT('h10)
	) name408 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_vld_req_any_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2637_
	);
	LUT4 #(
		.INIT('h080f)
	) name409 (
		_w2546_,
		_w2572_,
		_w2636_,
		_w2637_,
		_w2638_
	);
	LUT4 #(
		.INIT('h8acf)
	) name410 (
		_w2539_,
		_w2565_,
		_w2581_,
		_w2587_,
		_w2639_
	);
	LUT4 #(
		.INIT('hab00)
	) name411 (
		_w2594_,
		_w2605_,
		_w2614_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		_w2599_,
		_w2632_,
		_w2641_
	);
	LUT3 #(
		.INIT('h10)
	) name413 (
		_w2638_,
		_w2640_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w2583_,
		_w2591_,
		_w2643_
	);
	LUT4 #(
		.INIT('h1110)
	) name415 (
		_w2583_,
		_w2588_,
		_w2594_,
		_w2608_,
		_w2644_
	);
	LUT3 #(
		.INIT('h80)
	) name416 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2645_
	);
	LUT3 #(
		.INIT('h10)
	) name417 (
		_w2643_,
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('h01)
	) name418 (
		_w2635_,
		_w2642_,
		_w2646_,
		_w2647_
	);
	LUT3 #(
		.INIT('hdf)
	) name419 (
		_w2619_,
		_w2630_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		_w2578_,
		_w2649_
	);
	LUT3 #(
		.INIT('h10)
	) name421 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_vld_req_any_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2650_
	);
	LUT4 #(
		.INIT('h080f)
	) name422 (
		_w2546_,
		_w2572_,
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h4)
	) name423 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2652_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2653_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w2545_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2656_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w2571_,
		_w2656_,
		_w2657_
	);
	LUT4 #(
		.INIT('h2300)
	) name429 (
		_w2531_,
		_w2571_,
		_w2655_,
		_w2656_,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w2654_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2660_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		_w2565_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\ctl_rf_c3_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chpri_reg[1]/NET0131 ,
		_w2662_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		_w2539_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h8acf)
	) name435 (
		_w2539_,
		_w2565_,
		_w2660_,
		_w2662_,
		_w2664_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		\ctl_rf_c2_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chpri_reg[1]/NET0131 ,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w2559_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('h4500)
	) name438 (
		_w2559_,
		_w2565_,
		_w2660_,
		_w2665_,
		_w2667_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\ctl_rf_c0_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chpri_reg[1]/NET0131 ,
		_w2668_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w2553_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h8caf)
	) name441 (
		_w2531_,
		_w2553_,
		_w2655_,
		_w2668_,
		_w2670_
	);
	LUT3 #(
		.INIT('h10)
	) name442 (
		_w2664_,
		_w2667_,
		_w2670_,
		_w2671_
	);
	LUT4 #(
		.INIT('h4404)
	) name443 (
		_w2651_,
		_w2652_,
		_w2659_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2673_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		_w2578_,
		_w2673_,
		_w2674_
	);
	LUT4 #(
		.INIT('h8f00)
	) name446 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		\ctl_rf_c4_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chpri_reg[1]/NET0131 ,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w2524_,
		_w2676_,
		_w2677_
	);
	LUT4 #(
		.INIT('h2030)
	) name449 (
		_w2524_,
		_w2545_,
		_w2653_,
		_w2676_,
		_w2678_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w2663_,
		_w2678_,
		_w2679_
	);
	LUT3 #(
		.INIT('h32)
	) name451 (
		_w2663_,
		_w2666_,
		_w2678_,
		_w2680_
	);
	LUT4 #(
		.INIT('h8acf)
	) name452 (
		_w2524_,
		_w2559_,
		_w2665_,
		_w2676_,
		_w2681_
	);
	LUT3 #(
		.INIT('he0)
	) name453 (
		_w2658_,
		_w2670_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('h02)
	) name454 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2683_
	);
	LUT4 #(
		.INIT('hfe00)
	) name455 (
		_w2579_,
		_w2680_,
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('h08)
	) name456 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2685_
	);
	LUT3 #(
		.INIT('h0e)
	) name457 (
		_w2654_,
		_w2658_,
		_w2677_,
		_w2686_
	);
	LUT3 #(
		.INIT('h04)
	) name458 (
		_w2667_,
		_w2670_,
		_w2677_,
		_w2687_
	);
	LUT4 #(
		.INIT('hccc8)
	) name459 (
		_w2579_,
		_w2685_,
		_w2686_,
		_w2687_,
		_w2688_
	);
	LUT4 #(
		.INIT('h0001)
	) name460 (
		_w2672_,
		_w2675_,
		_w2684_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2690_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w2664_,
		_w2667_,
		_w2691_
	);
	LUT3 #(
		.INIT('he0)
	) name463 (
		_w2654_,
		_w2658_,
		_w2681_,
		_w2692_
	);
	LUT4 #(
		.INIT('h4440)
	) name464 (
		_w2651_,
		_w2690_,
		_w2691_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h00ea)
	) name465 (
		_w2658_,
		_w2661_,
		_w2670_,
		_w2677_,
		_w2694_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		_w2578_,
		_w2695_
	);
	LUT3 #(
		.INIT('h20)
	) name467 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_vld_req_any_d1_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2696_
	);
	LUT4 #(
		.INIT('h080f)
	) name468 (
		_w2546_,
		_w2572_,
		_w2695_,
		_w2696_,
		_w2697_
	);
	LUT4 #(
		.INIT('h00c4)
	) name469 (
		_w2679_,
		_w2690_,
		_w2694_,
		_w2697_,
		_w2698_
	);
	LUT3 #(
		.INIT('h80)
	) name470 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2699_
	);
	LUT4 #(
		.INIT('h4050)
	) name471 (
		_w2531_,
		_w2545_,
		_w2655_,
		_w2699_,
		_w2700_
	);
	LUT3 #(
		.INIT('h04)
	) name472 (
		_w2669_,
		_w2681_,
		_w2700_,
		_w2701_
	);
	LUT3 #(
		.INIT('h40)
	) name473 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		_w2702_
	);
	LUT4 #(
		.INIT('h8acf)
	) name474 (
		_w2531_,
		_w2553_,
		_w2668_,
		_w2702_,
		_w2703_
	);
	LUT3 #(
		.INIT('h10)
	) name475 (
		_w2664_,
		_w2667_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		_w2658_,
		_w2705_
	);
	LUT4 #(
		.INIT('haaa8)
	) name477 (
		_w2673_,
		_w2701_,
		_w2704_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h0301)
	) name478 (
		_w2664_,
		_w2667_,
		_w2669_,
		_w2678_,
		_w2707_
	);
	LUT4 #(
		.INIT('h0a08)
	) name479 (
		_w2652_,
		_w2657_,
		_w2697_,
		_w2707_,
		_w2708_
	);
	LUT4 #(
		.INIT('h0001)
	) name480 (
		_w2693_,
		_w2698_,
		_w2706_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h7)
	) name481 (
		_w2689_,
		_w2709_,
		_w2710_
	);
	LUT3 #(
		.INIT('h01)
	) name482 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2712_
	);
	LUT3 #(
		.INIT('h40)
	) name484 (
		_w2565_,
		_w2711_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		\ctl_rf_c3_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chpri_reg[1]/NET0131 ,
		_w2714_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w2539_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		\ctl_rf_c4_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chpri_reg[1]/NET0131 ,
		_w2716_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w2524_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('h4500)
	) name489 (
		_w2524_,
		_w2539_,
		_w2714_,
		_w2716_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		_w2531_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2721_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		_w2571_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h2300)
	) name494 (
		_w2531_,
		_w2571_,
		_w2719_,
		_w2721_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2724_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		_w2545_,
		_w2724_,
		_w2725_
	);
	LUT4 #(
		.INIT('h8caf)
	) name497 (
		_w2539_,
		_w2545_,
		_w2714_,
		_w2724_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		\ctl_rf_c2_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chpri_reg[1]/NET0131 ,
		_w2727_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		_w2559_,
		_w2727_,
		_w2728_
	);
	LUT3 #(
		.INIT('h8c)
	) name500 (
		_w2559_,
		_w2711_,
		_w2727_,
		_w2729_
	);
	LUT4 #(
		.INIT('h4500)
	) name501 (
		_w2718_,
		_w2723_,
		_w2726_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w2713_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		\ctl_rf_c0_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chpri_reg[1]/NET0131 ,
		_w2732_
	);
	LUT4 #(
		.INIT('h8acf)
	) name504 (
		_w2553_,
		_w2559_,
		_w2727_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h0301)
	) name505 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2718_,
		_w2726_,
		_w2733_,
		_w2734_
	);
	LUT4 #(
		.INIT('h8caf)
	) name506 (
		_w2524_,
		_w2531_,
		_w2716_,
		_w2719_,
		_w2735_
	);
	LUT4 #(
		.INIT('h2030)
	) name507 (
		_w2553_,
		_w2565_,
		_w2712_,
		_w2732_,
		_w2736_
	);
	LUT4 #(
		.INIT('hfac8)
	) name508 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2722_,
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		_w2738_
	);
	LUT3 #(
		.INIT('he0)
	) name510 (
		_w2734_,
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT3 #(
		.INIT('h51)
	) name511 (
		_w2579_,
		_w2731_,
		_w2739_,
		_w2740_
	);
	LUT3 #(
		.INIT('h02)
	) name512 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2741_
	);
	LUT4 #(
		.INIT('h4500)
	) name513 (
		_w2553_,
		_w2571_,
		_w2721_,
		_w2732_,
		_w2742_
	);
	LUT4 #(
		.INIT('hee0e)
	) name514 (
		_w2718_,
		_w2726_,
		_w2735_,
		_w2742_,
		_w2743_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name515 (
		_w2579_,
		_w2728_,
		_w2741_,
		_w2743_,
		_w2744_
	);
	LUT3 #(
		.INIT('h08)
	) name516 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w2723_,
		_w2725_,
		_w2746_
	);
	LUT3 #(
		.INIT('h54)
	) name518 (
		_w2717_,
		_w2723_,
		_w2725_,
		_w2747_
	);
	LUT3 #(
		.INIT('hc8)
	) name519 (
		_w2733_,
		_w2735_,
		_w2736_,
		_w2748_
	);
	LUT4 #(
		.INIT('hccc8)
	) name520 (
		_w2579_,
		_w2745_,
		_w2747_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('hccdf)
	) name521 (
		_w2715_,
		_w2720_,
		_w2733_,
		_w2736_,
		_w2750_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2751_
	);
	LUT3 #(
		.INIT('h10)
	) name523 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2752_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w2578_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w2574_,
		_w2752_,
		_w2754_
	);
	LUT4 #(
		.INIT('h080f)
	) name526 (
		_w2546_,
		_w2572_,
		_w2753_,
		_w2754_,
		_w2755_
	);
	LUT3 #(
		.INIT('h07)
	) name527 (
		_w2746_,
		_w2750_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2757_
	);
	LUT4 #(
		.INIT('h44c4)
	) name529 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		_w2720_,
		_w2726_,
		_w2736_,
		_w2758_
	);
	LUT3 #(
		.INIT('h01)
	) name530 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2759_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w2571_,
		_w2759_,
		_w2760_
	);
	LUT4 #(
		.INIT('h000b)
	) name532 (
		_w2718_,
		_w2733_,
		_w2736_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h7773)
	) name533 (
		_w2579_,
		_w2757_,
		_w2758_,
		_w2761_,
		_w2762_
	);
	LUT4 #(
		.INIT('h0100)
	) name534 (
		_w2744_,
		_w2749_,
		_w2756_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('hb)
	) name535 (
		_w2740_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		\ctl_rf_c3_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chpri_reg[1]/NET0131 ,
		_w2765_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		_w2539_,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2767_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		\ctl_rf_c0_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chpri_reg[1]/NET0131 ,
		_w2768_
	);
	LUT4 #(
		.INIT('h2030)
	) name540 (
		_w2553_,
		_w2565_,
		_w2767_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2771_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w2571_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h8caf)
	) name544 (
		_w2545_,
		_w2571_,
		_w2770_,
		_w2771_,
		_w2773_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\ctl_rf_c4_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chpri_reg[1]/NET0131 ,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w2524_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		_w2776_
	);
	LUT4 #(
		.INIT('h4500)
	) name548 (
		_w2531_,
		_w2545_,
		_w2770_,
		_w2776_,
		_w2777_
	);
	LUT4 #(
		.INIT('h000b)
	) name549 (
		_w2769_,
		_w2773_,
		_w2775_,
		_w2777_,
		_w2778_
	);
	LUT3 #(
		.INIT('h04)
	) name550 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2779_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		_w2578_,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w2574_,
		_w2779_,
		_w2781_
	);
	LUT4 #(
		.INIT('h080f)
	) name553 (
		_w2546_,
		_w2572_,
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2783_
	);
	LUT3 #(
		.INIT('ha8)
	) name555 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		_w2578_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h8f00)
	) name557 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h00f1)
	) name558 (
		_w2766_,
		_w2778_,
		_w2782_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name559 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2788_
	);
	LUT3 #(
		.INIT('h08)
	) name560 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2789_
	);
	LUT4 #(
		.INIT('h2030)
	) name561 (
		_w2524_,
		_w2545_,
		_w2770_,
		_w2774_,
		_w2790_
	);
	LUT4 #(
		.INIT('h8caf)
	) name562 (
		_w2524_,
		_w2531_,
		_w2774_,
		_w2776_,
		_w2791_
	);
	LUT3 #(
		.INIT('h13)
	) name563 (
		_w2772_,
		_w2790_,
		_w2791_,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		\ctl_rf_c2_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chpri_reg[1]/NET0131 ,
		_w2793_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w2559_,
		_w2793_,
		_w2794_
	);
	LUT4 #(
		.INIT('h8caf)
	) name566 (
		_w2553_,
		_w2559_,
		_w2768_,
		_w2793_,
		_w2795_
	);
	LUT3 #(
		.INIT('hc8)
	) name567 (
		_w2769_,
		_w2791_,
		_w2795_,
		_w2796_
	);
	LUT3 #(
		.INIT('ha2)
	) name568 (
		_w2789_,
		_w2792_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('h8caf)
	) name569 (
		_w2539_,
		_w2565_,
		_w2765_,
		_w2767_,
		_w2798_
	);
	LUT3 #(
		.INIT('h0e)
	) name570 (
		_w2769_,
		_w2795_,
		_w2798_,
		_w2799_
	);
	LUT3 #(
		.INIT('h10)
	) name571 (
		_w2775_,
		_w2777_,
		_w2795_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2801_
	);
	LUT3 #(
		.INIT('h80)
	) name573 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2802_
	);
	LUT3 #(
		.INIT('he0)
	) name574 (
		_w2799_,
		_w2800_,
		_w2802_,
		_w2803_
	);
	LUT3 #(
		.INIT('h02)
	) name575 (
		_w2787_,
		_w2797_,
		_w2803_,
		_w2804_
	);
	LUT3 #(
		.INIT('h01)
	) name576 (
		_w2769_,
		_w2772_,
		_w2795_,
		_w2805_
	);
	LUT3 #(
		.INIT('h10)
	) name577 (
		_w2772_,
		_w2790_,
		_w2798_,
		_w2806_
	);
	LUT3 #(
		.INIT('h40)
	) name578 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2807_
	);
	LUT2 #(
		.INIT('h4)
	) name579 (
		_w2578_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		_w2574_,
		_w2807_,
		_w2809_
	);
	LUT4 #(
		.INIT('h080f)
	) name581 (
		_w2546_,
		_w2572_,
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT3 #(
		.INIT('h01)
	) name582 (
		_w2805_,
		_w2806_,
		_w2810_,
		_w2811_
	);
	LUT3 #(
		.INIT('h45)
	) name583 (
		_w2772_,
		_w2775_,
		_w2795_,
		_w2812_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2813_
	);
	LUT3 #(
		.INIT('h20)
	) name585 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2814_
	);
	LUT3 #(
		.INIT('hb0)
	) name586 (
		_w2531_,
		_w2776_,
		_w2814_,
		_w2815_
	);
	LUT3 #(
		.INIT('hb0)
	) name587 (
		_w2799_,
		_w2812_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w2811_,
		_w2816_,
		_w2817_
	);
	LUT3 #(
		.INIT('h01)
	) name589 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2818_
	);
	LUT3 #(
		.INIT('h40)
	) name590 (
		_w2565_,
		_w2767_,
		_w2818_,
		_w2819_
	);
	LUT4 #(
		.INIT('h0105)
	) name591 (
		_w2766_,
		_w2772_,
		_w2790_,
		_w2791_,
		_w2820_
	);
	LUT3 #(
		.INIT('hb0)
	) name592 (
		_w2559_,
		_w2793_,
		_w2818_,
		_w2821_
	);
	LUT3 #(
		.INIT('h45)
	) name593 (
		_w2819_,
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('hcc04)
	) name594 (
		_w2769_,
		_w2773_,
		_w2795_,
		_w2798_,
		_w2823_
	);
	LUT3 #(
		.INIT('h10)
	) name595 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2824_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		_w2777_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w2823_,
		_w2825_,
		_w2826_
	);
	LUT3 #(
		.INIT('h51)
	) name598 (
		_w2579_,
		_w2822_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w2791_,
		_w2795_,
		_w2828_
	);
	LUT4 #(
		.INIT('h0054)
	) name600 (
		_w2579_,
		_w2794_,
		_w2820_,
		_w2828_,
		_w2829_
	);
	LUT3 #(
		.INIT('h02)
	) name601 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2830_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w2829_,
		_w2830_,
		_w2831_
	);
	LUT4 #(
		.INIT('hfff7)
	) name603 (
		_w2804_,
		_w2817_,
		_w2827_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		_w2834_
	);
	LUT3 #(
		.INIT('h07)
	) name606 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w2835_
	);
	LUT3 #(
		.INIT('h70)
	) name607 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w2836_
	);
	LUT4 #(
		.INIT('hc884)
	) name608 (
		\de_m1_is_llp_reg/NET0131 ,
		\h1size[2]_pad ,
		_w2425_,
		_w2834_,
		_w2837_
	);
	LUT4 #(
		.INIT('h0080)
	) name609 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[10]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w2838_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w2425_,
		_w2838_,
		_w2839_
	);
	LUT4 #(
		.INIT('h8880)
	) name611 (
		\ch_sel_arb_chcsr_reg_reg[13]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w2840_
	);
	LUT3 #(
		.INIT('h15)
	) name612 (
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w2835_,
		_w2840_,
		_w2841_
	);
	LUT4 #(
		.INIT('h5455)
	) name613 (
		_w2833_,
		_w2837_,
		_w2839_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('hba8a)
	) name614 (
		\h1size[2]_pad ,
		_w2417_,
		_w2434_,
		_w2842_,
		_w2843_
	);
	LUT3 #(
		.INIT('h40)
	) name615 (
		_w2539_,
		_w2587_,
		_w2599_,
		_w2844_
	);
	LUT4 #(
		.INIT('h8acf)
	) name616 (
		_w2553_,
		_w2565_,
		_w2581_,
		_w2582_,
		_w2845_
	);
	LUT4 #(
		.INIT('h8acf)
	) name617 (
		_w2531_,
		_w2571_,
		_w2584_,
		_w2596_,
		_w2846_
	);
	LUT4 #(
		.INIT('h8caf)
	) name618 (
		_w2524_,
		_w2545_,
		_w2593_,
		_w2604_,
		_w2847_
	);
	LUT4 #(
		.INIT('h8a00)
	) name619 (
		_w2599_,
		_w2845_,
		_w2846_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('haaa8)
	) name620 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2579_,
		_w2844_,
		_w2848_,
		_w2849_
	);
	LUT3 #(
		.INIT('h04)
	) name621 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2850_
	);
	LUT3 #(
		.INIT('h20)
	) name622 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2571_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h8caf)
	) name623 (
		_w2539_,
		_w2559_,
		_w2587_,
		_w2589_,
		_w2852_
	);
	LUT4 #(
		.INIT('h8088)
	) name624 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2845_,
		_w2847_,
		_w2852_,
		_w2853_
	);
	LUT3 #(
		.INIT('h45)
	) name625 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		_w2545_,
		_w2604_,
		_w2854_
	);
	LUT4 #(
		.INIT('h3b00)
	) name626 (
		_w2845_,
		_w2846_,
		_w2852_,
		_w2854_,
		_w2855_
	);
	LUT4 #(
		.INIT('h0203)
	) name627 (
		_w2638_,
		_w2851_,
		_w2853_,
		_w2855_,
		_w2856_
	);
	LUT4 #(
		.INIT('h8a00)
	) name628 (
		_w2631_,
		_w2845_,
		_w2846_,
		_w2847_,
		_w2857_
	);
	LUT3 #(
		.INIT('h04)
	) name629 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2858_
	);
	LUT3 #(
		.INIT('h45)
	) name630 (
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2565_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h4f00)
	) name631 (
		_w2846_,
		_w2847_,
		_w2852_,
		_w2859_,
		_w2860_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name632 (
		_w2504_,
		_w2845_,
		_w2846_,
		_w2852_,
		_w2861_
	);
	LUT4 #(
		.INIT('h2223)
	) name633 (
		_w2638_,
		_w2857_,
		_w2860_,
		_w2861_,
		_w2862_
	);
	LUT4 #(
		.INIT('hceff)
	) name634 (
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2849_,
		_w2856_,
		_w2862_,
		_w2863_
	);
	LUT4 #(
		.INIT('h8caf)
	) name635 (
		_w2539_,
		_w2559_,
		_w2765_,
		_w2793_,
		_w2864_
	);
	LUT4 #(
		.INIT('h8acf)
	) name636 (
		_w2524_,
		_w2545_,
		_w2770_,
		_w2774_,
		_w2865_
	);
	LUT4 #(
		.INIT('h8acf)
	) name637 (
		_w2531_,
		_w2571_,
		_w2771_,
		_w2776_,
		_w2866_
	);
	LUT3 #(
		.INIT('h10)
	) name638 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2867_
	);
	LUT3 #(
		.INIT('h8c)
	) name639 (
		_w2565_,
		_w2783_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h5d00)
	) name640 (
		_w2864_,
		_w2865_,
		_w2866_,
		_w2868_,
		_w2869_
	);
	LUT4 #(
		.INIT('h8acf)
	) name641 (
		_w2553_,
		_w2565_,
		_w2767_,
		_w2768_,
		_w2870_
	);
	LUT3 #(
		.INIT('h10)
	) name642 (
		\ch_sel_dma_rrarb2_state_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2871_
	);
	LUT3 #(
		.INIT('h8c)
	) name643 (
		_w2545_,
		_w2813_,
		_w2871_,
		_w2872_
	);
	LUT4 #(
		.INIT('h7300)
	) name644 (
		_w2864_,
		_w2866_,
		_w2870_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('h54)
	) name645 (
		_w2579_,
		_w2869_,
		_w2873_,
		_w2874_
	);
	LUT4 #(
		.INIT('h8808)
	) name646 (
		_w2788_,
		_w2865_,
		_w2866_,
		_w2870_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		_w2578_,
		_w2876_
	);
	LUT4 #(
		.INIT('h8f00)
	) name648 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2876_,
		_w2877_
	);
	LUT3 #(
		.INIT('h07)
	) name649 (
		\ch_sel_dma_rrarb2_state_reg[1]/NET0131 ,
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT3 #(
		.INIT('h40)
	) name650 (
		_w2539_,
		_w2765_,
		_w2779_,
		_w2879_
	);
	LUT4 #(
		.INIT('h8808)
	) name651 (
		_w2779_,
		_w2865_,
		_w2866_,
		_w2870_,
		_w2880_
	);
	LUT4 #(
		.INIT('ha200)
	) name652 (
		_w2801_,
		_w2864_,
		_w2865_,
		_w2870_,
		_w2881_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		_w2771_,
		_w2807_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w2571_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h0001)
	) name655 (
		_w2879_,
		_w2880_,
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT3 #(
		.INIT('hbf)
	) name656 (
		_w2874_,
		_w2878_,
		_w2884_,
		_w2885_
	);
	LUT3 #(
		.INIT('h40)
	) name657 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2887_
	);
	LUT3 #(
		.INIT('h40)
	) name659 (
		_w2571_,
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('h8acf)
	) name660 (
		_w2524_,
		_w2545_,
		_w2653_,
		_w2676_,
		_w2889_
	);
	LUT4 #(
		.INIT('h8caf)
	) name661 (
		_w2539_,
		_w2559_,
		_w2662_,
		_w2665_,
		_w2890_
	);
	LUT4 #(
		.INIT('h8acf)
	) name662 (
		_w2553_,
		_w2565_,
		_w2660_,
		_w2668_,
		_w2891_
	);
	LUT4 #(
		.INIT('h8a00)
	) name663 (
		_w2887_,
		_w2889_,
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('h8caf)
	) name664 (
		_w2531_,
		_w2571_,
		_w2655_,
		_w2656_,
		_w2893_
	);
	LUT4 #(
		.INIT('h8088)
	) name665 (
		_w2685_,
		_w2889_,
		_w2891_,
		_w2893_,
		_w2894_
	);
	LUT3 #(
		.INIT('hc8)
	) name666 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2895_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w2578_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h8f00)
	) name668 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h0001)
	) name669 (
		_w2888_,
		_w2892_,
		_w2894_,
		_w2897_,
		_w2898_
	);
	LUT3 #(
		.INIT('hc4)
	) name670 (
		_w2889_,
		_w2890_,
		_w2893_,
		_w2899_
	);
	LUT3 #(
		.INIT('h40)
	) name671 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2901_
	);
	LUT3 #(
		.INIT('hb0)
	) name673 (
		_w2565_,
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h2300)
	) name674 (
		_w2565_,
		_w2578_,
		_w2900_,
		_w2901_,
		_w2903_
	);
	LUT4 #(
		.INIT('h8c00)
	) name675 (
		_w2565_,
		_w2574_,
		_w2900_,
		_w2901_,
		_w2904_
	);
	LUT4 #(
		.INIT('h080f)
	) name676 (
		_w2546_,
		_w2572_,
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('h20aa)
	) name677 (
		_w2673_,
		_w2890_,
		_w2891_,
		_w2893_,
		_w2906_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name678 (
		_w2651_,
		_w2899_,
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT3 #(
		.INIT('h04)
	) name679 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2908_
	);
	LUT3 #(
		.INIT('h8a)
	) name680 (
		_w2889_,
		_w2891_,
		_w2893_,
		_w2909_
	);
	LUT3 #(
		.INIT('h23)
	) name681 (
		_w2539_,
		_w2578_,
		_w2662_,
		_w2910_
	);
	LUT3 #(
		.INIT('h8c)
	) name682 (
		_w2539_,
		_w2574_,
		_w2662_,
		_w2911_
	);
	LUT4 #(
		.INIT('h080f)
	) name683 (
		_w2546_,
		_w2572_,
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT3 #(
		.INIT('ha8)
	) name684 (
		_w2908_,
		_w2909_,
		_w2912_,
		_w2913_
	);
	LUT3 #(
		.INIT('h8c)
	) name685 (
		_w2545_,
		_w2652_,
		_w2653_,
		_w2914_
	);
	LUT4 #(
		.INIT('h4f00)
	) name686 (
		_w2890_,
		_w2891_,
		_w2893_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		_w2651_,
		_w2915_,
		_w2916_
	);
	LUT4 #(
		.INIT('hfff7)
	) name688 (
		_w2898_,
		_w2907_,
		_w2913_,
		_w2916_,
		_w2917_
	);
	LUT3 #(
		.INIT('h8a)
	) name689 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		_w2571_,
		_w2850_,
		_w2918_
	);
	LUT3 #(
		.INIT('h04)
	) name690 (
		\ch_sel_dma_rrarb1_state_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2919_
	);
	LUT2 #(
		.INIT('h4)
	) name691 (
		_w2545_,
		_w2919_,
		_w2920_
	);
	LUT3 #(
		.INIT('h31)
	) name692 (
		_w2846_,
		_w2918_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		_w2845_,
		_w2852_,
		_w2922_
	);
	LUT4 #(
		.INIT('haaa8)
	) name694 (
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2579_,
		_w2921_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		\ch_sel_dma_rrarb1_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb1_state_reg[2]/NET0131 ,
		_w2924_
	);
	LUT3 #(
		.INIT('hb0)
	) name696 (
		_w2565_,
		_w2858_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('h004f)
	) name697 (
		_w2539_,
		_w2587_,
		_w2600_,
		_w2631_,
		_w2926_
	);
	LUT3 #(
		.INIT('h70)
	) name698 (
		_w2852_,
		_w2925_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		_w2846_,
		_w2847_,
		_w2928_
	);
	LUT3 #(
		.INIT('h01)
	) name700 (
		_w2579_,
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('he)
	) name701 (
		_w2923_,
		_w2929_,
		_w2930_
	);
	LUT3 #(
		.INIT('hb0)
	) name702 (
		_w2539_,
		_w2765_,
		_w2779_,
		_w2931_
	);
	LUT4 #(
		.INIT('h0015)
	) name703 (
		_w2789_,
		_w2864_,
		_w2868_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		_w2865_,
		_w2866_,
		_w2933_
	);
	LUT3 #(
		.INIT('h01)
	) name705 (
		_w2579_,
		_w2932_,
		_w2933_,
		_w2934_
	);
	LUT3 #(
		.INIT('h80)
	) name706 (
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2795_,
		_w2798_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		\ch_sel_dma_rrarb2_state_reg[2]/NET0131 ,
		_w2578_,
		_w2936_
	);
	LUT4 #(
		.INIT('h8f00)
	) name708 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w2936_,
		_w2937_
	);
	LUT3 #(
		.INIT('h23)
	) name709 (
		_w2571_,
		_w2813_,
		_w2882_,
		_w2938_
	);
	LUT4 #(
		.INIT('h8caf)
	) name710 (
		_w2545_,
		_w2571_,
		_w2871_,
		_w2882_,
		_w2939_
	);
	LUT3 #(
		.INIT('h13)
	) name711 (
		_w2866_,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h01)
	) name712 (
		_w2935_,
		_w2937_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('hb)
	) name713 (
		_w2934_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('h8a)
	) name714 (
		\ch_sel_dma_rrarb3_state_reg[1]/NET0131 ,
		_w2571_,
		_w2886_,
		_w2943_
	);
	LUT3 #(
		.INIT('h40)
	) name715 (
		\ch_sel_dma_rrarb3_state_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2944_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		_w2545_,
		_w2944_,
		_w2945_
	);
	LUT3 #(
		.INIT('h31)
	) name717 (
		_w2893_,
		_w2943_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		_w2890_,
		_w2891_,
		_w2947_
	);
	LUT4 #(
		.INIT('haaa8)
	) name719 (
		\ch_sel_dma_rrarb3_state_reg[2]/NET0131 ,
		_w2579_,
		_w2946_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		_w2889_,
		_w2893_,
		_w2949_
	);
	LUT4 #(
		.INIT('h040f)
	) name721 (
		_w2539_,
		_w2662_,
		_w2685_,
		_w2908_,
		_w2950_
	);
	LUT3 #(
		.INIT('h70)
	) name722 (
		_w2890_,
		_w2902_,
		_w2950_,
		_w2951_
	);
	LUT3 #(
		.INIT('h01)
	) name723 (
		_w2579_,
		_w2949_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('he)
	) name724 (
		_w2948_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('h0073)
	) name725 (
		_w2565_,
		_w2711_,
		_w2712_,
		_w2741_,
		_w2954_
	);
	LUT4 #(
		.INIT('h8caf)
	) name726 (
		_w2539_,
		_w2559_,
		_w2714_,
		_w2727_,
		_w2955_
	);
	LUT4 #(
		.INIT('h8caf)
	) name727 (
		_w2524_,
		_w2545_,
		_w2716_,
		_w2724_,
		_w2956_
	);
	LUT4 #(
		.INIT('h8caf)
	) name728 (
		_w2531_,
		_w2571_,
		_w2719_,
		_w2721_,
		_w2957_
	);
	LUT4 #(
		.INIT('h1151)
	) name729 (
		_w2954_,
		_w2955_,
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h8acf)
	) name730 (
		_w2553_,
		_w2565_,
		_w2712_,
		_w2732_,
		_w2959_
	);
	LUT3 #(
		.INIT('h01)
	) name731 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		_w2960_
	);
	LUT2 #(
		.INIT('h4)
	) name732 (
		_w2545_,
		_w2960_,
		_w2961_
	);
	LUT3 #(
		.INIT('h8c)
	) name733 (
		_w2545_,
		_w2751_,
		_w2960_,
		_w2962_
	);
	LUT4 #(
		.INIT('h7300)
	) name734 (
		_w2955_,
		_w2957_,
		_w2959_,
		_w2962_,
		_w2963_
	);
	LUT3 #(
		.INIT('h54)
	) name735 (
		_w2579_,
		_w2958_,
		_w2963_,
		_w2964_
	);
	LUT3 #(
		.INIT('h04)
	) name736 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w2714_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w2539_,
		_w2966_,
		_w2967_
	);
	LUT3 #(
		.INIT('h01)
	) name739 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2969_
	);
	LUT3 #(
		.INIT('h40)
	) name741 (
		_w2571_,
		_w2968_,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w2967_,
		_w2970_,
		_w2971_
	);
	LUT3 #(
		.INIT('h01)
	) name743 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		_w2967_,
		_w2970_,
		_w2972_
	);
	LUT3 #(
		.INIT('h04)
	) name744 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2956_,
		_w2957_,
		_w2973_
	);
	LUT4 #(
		.INIT('hf200)
	) name745 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2955_,
		_w2956_,
		_w2959_,
		_w2974_
	);
	LUT4 #(
		.INIT('h0004)
	) name746 (
		_w2579_,
		_w2971_,
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT3 #(
		.INIT('hab)
	) name747 (
		_w2964_,
		_w2972_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('hcc40)
	) name748 (
		_w2424_,
		_w2482_,
		_w2485_,
		_w2486_,
		_w2977_
	);
	LUT3 #(
		.INIT('h8a)
	) name749 (
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		_w2571_,
		_w2968_,
		_w2978_
	);
	LUT3 #(
		.INIT('h0d)
	) name750 (
		_w2957_,
		_w2961_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		_w2955_,
		_w2959_,
		_w2980_
	);
	LUT4 #(
		.INIT('haaa8)
	) name752 (
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2579_,
		_w2979_,
		_w2980_,
		_w2981_
	);
	LUT3 #(
		.INIT('h04)
	) name753 (
		_w2559_,
		_w2727_,
		_w2965_,
		_w2982_
	);
	LUT3 #(
		.INIT('hf9)
	) name754 (
		\ch_sel_dma_rrarb0_state_reg[0]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[1]/NET0131 ,
		\ch_sel_dma_rrarb0_state_reg[2]/NET0131 ,
		_w2983_
	);
	LUT4 #(
		.INIT('h7300)
	) name755 (
		_w2565_,
		_w2711_,
		_w2712_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('h3332)
	) name756 (
		_w2715_,
		_w2745_,
		_w2982_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w2956_,
		_w2957_,
		_w2986_
	);
	LUT3 #(
		.INIT('h01)
	) name758 (
		_w2579_,
		_w2985_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('he)
	) name759 (
		_w2981_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		_w2989_
	);
	LUT3 #(
		.INIT('hf4)
	) name761 (
		_w2455_,
		_w2477_,
		_w2989_,
		_w2990_
	);
	LUT4 #(
		.INIT('h0100)
	) name762 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w2991_
	);
	LUT3 #(
		.INIT('h80)
	) name763 (
		_w2230_,
		_w2247_,
		_w2991_,
		_w2992_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name764 (
		\hwdata[15]_pad ,
		\hwdata[23]_pad ,
		_w2234_,
		_w2235_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\hwdata[31]_pad ,
		_w2234_,
		_w2994_
	);
	LUT4 #(
		.INIT('hbbb3)
	) name766 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2992_,
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name767 (
		\hwdata[0]_pad ,
		\hwdata[24]_pad ,
		_w2234_,
		_w2235_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\hwdata[16]_pad ,
		_w2234_,
		_w2997_
	);
	LUT2 #(
		.INIT('he)
	) name769 (
		_w2996_,
		_w2997_,
		_w2998_
	);
	LUT3 #(
		.INIT('ha8)
	) name770 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2996_,
		_w2997_,
		_w2999_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w2995_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('h2a)
	) name772 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3001_
	);
	LUT3 #(
		.INIT('h80)
	) name773 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3002_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name774 (
		_w2514_,
		_w2518_,
		_w3001_,
		_w3002_,
		_w3003_
	);
	LUT3 #(
		.INIT('h2a)
	) name775 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3004_
	);
	LUT3 #(
		.INIT('h80)
	) name776 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3005_
	);
	LUT4 #(
		.INIT('h67ef)
	) name777 (
		_w2514_,
		_w2518_,
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('h2a)
	) name778 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3007_
	);
	LUT3 #(
		.INIT('h80)
	) name779 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3008_
	);
	LUT4 #(
		.INIT('hcedf)
	) name780 (
		_w2514_,
		_w2518_,
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT3 #(
		.INIT('h80)
	) name781 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3010_
	);
	LUT3 #(
		.INIT('h2a)
	) name782 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3011_
	);
	LUT3 #(
		.INIT('h57)
	) name783 (
		_w2534_,
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('h8000)
	) name784 (
		_w3003_,
		_w3006_,
		_w3009_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h2)
	) name785 (
		_w2521_,
		_w3013_,
		_w3014_
	);
	LUT4 #(
		.INIT('h0001)
	) name786 (
		\ctl_rf_c2_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[30]/NET0131 ,
		_w3015_
	);
	LUT4 #(
		.INIT('h0001)
	) name787 (
		\ctl_rf_c2_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[27]/NET0131 ,
		_w3016_
	);
	LUT4 #(
		.INIT('h0001)
	) name788 (
		\ctl_rf_c2_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[9]/NET0131 ,
		_w3017_
	);
	LUT4 #(
		.INIT('h0001)
	) name789 (
		\ctl_rf_c2_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[5]/NET0131 ,
		_w3018_
	);
	LUT4 #(
		.INIT('h8000)
	) name790 (
		_w3015_,
		_w3016_,
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		\ctl_rf_c2_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[11]/NET0131 ,
		_w3020_
	);
	LUT4 #(
		.INIT('h0001)
	) name792 (
		\ctl_rf_c2_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[15]/NET0131 ,
		_w3021_
	);
	LUT4 #(
		.INIT('h0001)
	) name793 (
		\ctl_rf_c2_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[23]/NET0131 ,
		_w3022_
	);
	LUT4 #(
		.INIT('h0001)
	) name794 (
		\ctl_rf_c2_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c2_rf_chllp_reg[19]/NET0131 ,
		_w3023_
	);
	LUT4 #(
		.INIT('h8000)
	) name795 (
		_w3020_,
		_w3021_,
		_w3022_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h0888)
	) name796 (
		_w2509_,
		_w2534_,
		_w3019_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('h0001)
	) name797 (
		\ctl_rf_c4_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[30]/NET0131 ,
		_w3026_
	);
	LUT4 #(
		.INIT('h0001)
	) name798 (
		\ctl_rf_c4_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[27]/NET0131 ,
		_w3027_
	);
	LUT4 #(
		.INIT('h0001)
	) name799 (
		\ctl_rf_c4_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[9]/NET0131 ,
		_w3028_
	);
	LUT4 #(
		.INIT('h0001)
	) name800 (
		\ctl_rf_c4_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[5]/NET0131 ,
		_w3029_
	);
	LUT4 #(
		.INIT('h8000)
	) name801 (
		_w3026_,
		_w3027_,
		_w3028_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		\ctl_rf_c4_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[11]/NET0131 ,
		_w3031_
	);
	LUT4 #(
		.INIT('h0001)
	) name803 (
		\ctl_rf_c4_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[15]/NET0131 ,
		_w3032_
	);
	LUT4 #(
		.INIT('h0001)
	) name804 (
		\ctl_rf_c4_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[23]/NET0131 ,
		_w3033_
	);
	LUT4 #(
		.INIT('h0001)
	) name805 (
		\ctl_rf_c4_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[19]/NET0131 ,
		_w3034_
	);
	LUT4 #(
		.INIT('h8000)
	) name806 (
		_w3031_,
		_w3032_,
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('h0888)
	) name807 (
		_w2509_,
		_w2520_,
		_w3030_,
		_w3035_,
		_w3036_
	);
	LUT4 #(
		.INIT('h0001)
	) name808 (
		\ctl_rf_c1_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[30]/NET0131 ,
		_w3037_
	);
	LUT4 #(
		.INIT('h0001)
	) name809 (
		\ctl_rf_c1_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[27]/NET0131 ,
		_w3038_
	);
	LUT4 #(
		.INIT('h0001)
	) name810 (
		\ctl_rf_c1_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[9]/NET0131 ,
		_w3039_
	);
	LUT4 #(
		.INIT('h0001)
	) name811 (
		\ctl_rf_c1_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[5]/NET0131 ,
		_w3040_
	);
	LUT4 #(
		.INIT('h8000)
	) name812 (
		_w3037_,
		_w3038_,
		_w3039_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\ctl_rf_c1_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[11]/NET0131 ,
		_w3042_
	);
	LUT4 #(
		.INIT('h0001)
	) name814 (
		\ctl_rf_c1_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[15]/NET0131 ,
		_w3043_
	);
	LUT4 #(
		.INIT('h0001)
	) name815 (
		\ctl_rf_c1_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[23]/NET0131 ,
		_w3044_
	);
	LUT4 #(
		.INIT('h0001)
	) name816 (
		\ctl_rf_c1_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[19]/NET0131 ,
		_w3045_
	);
	LUT4 #(
		.INIT('h8000)
	) name817 (
		_w3042_,
		_w3043_,
		_w3044_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('h0444)
	) name818 (
		_w2509_,
		_w2549_,
		_w3041_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('h0001)
	) name819 (
		\ctl_rf_c3_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[30]/NET0131 ,
		_w3048_
	);
	LUT4 #(
		.INIT('h0001)
	) name820 (
		\ctl_rf_c3_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[27]/NET0131 ,
		_w3049_
	);
	LUT4 #(
		.INIT('h0001)
	) name821 (
		\ctl_rf_c3_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[9]/NET0131 ,
		_w3050_
	);
	LUT4 #(
		.INIT('h0001)
	) name822 (
		\ctl_rf_c3_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[5]/NET0131 ,
		_w3051_
	);
	LUT4 #(
		.INIT('h8000)
	) name823 (
		_w3048_,
		_w3049_,
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		\ctl_rf_c3_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[11]/NET0131 ,
		_w3053_
	);
	LUT4 #(
		.INIT('h0001)
	) name825 (
		\ctl_rf_c3_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[15]/NET0131 ,
		_w3054_
	);
	LUT4 #(
		.INIT('h0001)
	) name826 (
		\ctl_rf_c3_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[23]/NET0131 ,
		_w3055_
	);
	LUT4 #(
		.INIT('h0001)
	) name827 (
		\ctl_rf_c3_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[19]/NET0131 ,
		_w3056_
	);
	LUT4 #(
		.INIT('h8000)
	) name828 (
		_w3053_,
		_w3054_,
		_w3055_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h0444)
	) name829 (
		_w2509_,
		_w2534_,
		_w3052_,
		_w3057_,
		_w3058_
	);
	LUT4 #(
		.INIT('h0001)
	) name830 (
		_w3025_,
		_w3036_,
		_w3047_,
		_w3058_,
		_w3059_
	);
	LUT4 #(
		.INIT('h0001)
	) name831 (
		\ctl_rf_c7_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[30]/NET0131 ,
		_w3060_
	);
	LUT4 #(
		.INIT('h0001)
	) name832 (
		\ctl_rf_c7_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[27]/NET0131 ,
		_w3061_
	);
	LUT4 #(
		.INIT('h0001)
	) name833 (
		\ctl_rf_c7_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[9]/NET0131 ,
		_w3062_
	);
	LUT4 #(
		.INIT('h0001)
	) name834 (
		\ctl_rf_c7_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[5]/NET0131 ,
		_w3063_
	);
	LUT4 #(
		.INIT('h8000)
	) name835 (
		_w3060_,
		_w3061_,
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		\ctl_rf_c7_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[11]/NET0131 ,
		_w3065_
	);
	LUT4 #(
		.INIT('h0001)
	) name837 (
		\ctl_rf_c7_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[15]/NET0131 ,
		_w3066_
	);
	LUT4 #(
		.INIT('h0001)
	) name838 (
		\ctl_rf_c7_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[23]/NET0131 ,
		_w3067_
	);
	LUT4 #(
		.INIT('h0001)
	) name839 (
		\ctl_rf_c7_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[19]/NET0131 ,
		_w3068_
	);
	LUT4 #(
		.INIT('h8000)
	) name840 (
		_w3065_,
		_w3066_,
		_w3067_,
		_w3068_,
		_w3069_
	);
	LUT4 #(
		.INIT('h0444)
	) name841 (
		_w2509_,
		_w2527_,
		_w3064_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('h0001)
	) name842 (
		\ctl_rf_c5_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[30]/NET0131 ,
		_w3071_
	);
	LUT4 #(
		.INIT('h0001)
	) name843 (
		\ctl_rf_c5_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[27]/NET0131 ,
		_w3072_
	);
	LUT4 #(
		.INIT('h0001)
	) name844 (
		\ctl_rf_c5_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[9]/NET0131 ,
		_w3073_
	);
	LUT4 #(
		.INIT('h0001)
	) name845 (
		\ctl_rf_c5_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[5]/NET0131 ,
		_w3074_
	);
	LUT4 #(
		.INIT('h8000)
	) name846 (
		_w3071_,
		_w3072_,
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		\ctl_rf_c5_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[11]/NET0131 ,
		_w3076_
	);
	LUT4 #(
		.INIT('h0001)
	) name848 (
		\ctl_rf_c5_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[15]/NET0131 ,
		_w3077_
	);
	LUT4 #(
		.INIT('h0001)
	) name849 (
		\ctl_rf_c5_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[23]/NET0131 ,
		_w3078_
	);
	LUT4 #(
		.INIT('h0001)
	) name850 (
		\ctl_rf_c5_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[19]/NET0131 ,
		_w3079_
	);
	LUT4 #(
		.INIT('h8000)
	) name851 (
		_w3076_,
		_w3077_,
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0444)
	) name852 (
		_w2509_,
		_w2520_,
		_w3075_,
		_w3080_,
		_w3081_
	);
	LUT4 #(
		.INIT('h0001)
	) name853 (
		\ctl_rf_c0_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[30]/NET0131 ,
		_w3082_
	);
	LUT4 #(
		.INIT('h0001)
	) name854 (
		\ctl_rf_c0_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[27]/NET0131 ,
		_w3083_
	);
	LUT4 #(
		.INIT('h0001)
	) name855 (
		\ctl_rf_c0_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[9]/NET0131 ,
		_w3084_
	);
	LUT4 #(
		.INIT('h0001)
	) name856 (
		\ctl_rf_c0_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[5]/NET0131 ,
		_w3085_
	);
	LUT4 #(
		.INIT('h8000)
	) name857 (
		_w3082_,
		_w3083_,
		_w3084_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		\ctl_rf_c0_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[11]/NET0131 ,
		_w3087_
	);
	LUT4 #(
		.INIT('h0001)
	) name859 (
		\ctl_rf_c0_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[15]/NET0131 ,
		_w3088_
	);
	LUT4 #(
		.INIT('h0001)
	) name860 (
		\ctl_rf_c0_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[23]/NET0131 ,
		_w3089_
	);
	LUT4 #(
		.INIT('h0001)
	) name861 (
		\ctl_rf_c0_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c0_rf_chllp_reg[19]/NET0131 ,
		_w3090_
	);
	LUT4 #(
		.INIT('h8000)
	) name862 (
		_w3087_,
		_w3088_,
		_w3089_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h0888)
	) name863 (
		_w2509_,
		_w2549_,
		_w3086_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('h0001)
	) name864 (
		\ctl_rf_c6_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[30]/NET0131 ,
		_w3093_
	);
	LUT4 #(
		.INIT('h0001)
	) name865 (
		\ctl_rf_c6_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[27]/NET0131 ,
		_w3094_
	);
	LUT4 #(
		.INIT('h0001)
	) name866 (
		\ctl_rf_c6_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[9]/NET0131 ,
		_w3095_
	);
	LUT4 #(
		.INIT('h0001)
	) name867 (
		\ctl_rf_c6_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[5]/NET0131 ,
		_w3096_
	);
	LUT4 #(
		.INIT('h8000)
	) name868 (
		_w3093_,
		_w3094_,
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		\ctl_rf_c6_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[11]/NET0131 ,
		_w3098_
	);
	LUT4 #(
		.INIT('h0001)
	) name870 (
		\ctl_rf_c6_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[15]/NET0131 ,
		_w3099_
	);
	LUT4 #(
		.INIT('h0001)
	) name871 (
		\ctl_rf_c6_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[23]/NET0131 ,
		_w3100_
	);
	LUT4 #(
		.INIT('h0001)
	) name872 (
		\ctl_rf_c6_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[19]/NET0131 ,
		_w3101_
	);
	LUT4 #(
		.INIT('h8000)
	) name873 (
		_w3098_,
		_w3099_,
		_w3100_,
		_w3101_,
		_w3102_
	);
	LUT4 #(
		.INIT('h0888)
	) name874 (
		_w2509_,
		_w2527_,
		_w3097_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h0001)
	) name875 (
		_w3070_,
		_w3081_,
		_w3092_,
		_w3103_,
		_w3104_
	);
	LUT3 #(
		.INIT('h80)
	) name876 (
		_w2424_,
		_w2511_,
		_w2520_,
		_w3105_
	);
	LUT3 #(
		.INIT('h80)
	) name877 (
		_w3059_,
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h2)
	) name878 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2995_,
		_w3107_
	);
	LUT3 #(
		.INIT('h40)
	) name879 (
		\de_de_st_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3108_
	);
	LUT4 #(
		.INIT('ha222)
	) name880 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		_w2520_,
		_w3108_,
		_w3109_
	);
	LUT3 #(
		.INIT('hd0)
	) name881 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2995_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('habaa)
	) name882 (
		_w3000_,
		_w3014_,
		_w3106_,
		_w3110_,
		_w3111_
	);
	LUT4 #(
		.INIT('h1000)
	) name883 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w3112_
	);
	LUT3 #(
		.INIT('h80)
	) name884 (
		_w2230_,
		_w2247_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name885 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		_w2999_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		_w2542_,
		_w3013_,
		_w3116_
	);
	LUT3 #(
		.INIT('h80)
	) name888 (
		_w2424_,
		_w2520_,
		_w2535_,
		_w3117_
	);
	LUT3 #(
		.INIT('h80)
	) name889 (
		_w3059_,
		_w3104_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3114_,
		_w3119_
	);
	LUT3 #(
		.INIT('h15)
	) name891 (
		\de_de_st_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3120_
	);
	LUT4 #(
		.INIT('ha222)
	) name892 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		_w2520_,
		_w3120_,
		_w3121_
	);
	LUT3 #(
		.INIT('hd0)
	) name893 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3114_,
		_w3121_,
		_w3122_
	);
	LUT4 #(
		.INIT('habaa)
	) name894 (
		_w3115_,
		_w3116_,
		_w3118_,
		_w3122_,
		_w3123_
	);
	LUT3 #(
		.INIT('h80)
	) name895 (
		_w2230_,
		_w2254_,
		_w2991_,
		_w3124_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name896 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h2)
	) name897 (
		_w2999_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		_w2528_,
		_w3013_,
		_w3127_
	);
	LUT3 #(
		.INIT('h80)
	) name899 (
		_w2424_,
		_w2511_,
		_w2527_,
		_w3128_
	);
	LUT3 #(
		.INIT('h80)
	) name900 (
		_w3059_,
		_w3104_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h2)
	) name901 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3125_,
		_w3130_
	);
	LUT4 #(
		.INIT('ha222)
	) name902 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		_w2527_,
		_w3108_,
		_w3131_
	);
	LUT3 #(
		.INIT('hd0)
	) name903 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3125_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('habaa)
	) name904 (
		_w3126_,
		_w3127_,
		_w3129_,
		_w3132_,
		_w3133_
	);
	LUT3 #(
		.INIT('h80)
	) name905 (
		_w2230_,
		_w2254_,
		_w3112_,
		_w3134_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name906 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h2)
	) name907 (
		_w2999_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		_w2568_,
		_w3013_,
		_w3137_
	);
	LUT3 #(
		.INIT('h80)
	) name909 (
		_w2424_,
		_w2527_,
		_w2535_,
		_w3138_
	);
	LUT3 #(
		.INIT('h80)
	) name910 (
		_w3059_,
		_w3104_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3135_,
		_w3140_
	);
	LUT4 #(
		.INIT('ha222)
	) name912 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2527_,
		_w3120_,
		_w3141_
	);
	LUT3 #(
		.INIT('hd0)
	) name913 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3135_,
		_w3141_,
		_w3142_
	);
	LUT4 #(
		.INIT('habaa)
	) name914 (
		_w3136_,
		_w3137_,
		_w3139_,
		_w3142_,
		_w3143_
	);
	LUT3 #(
		.INIT('h80)
	) name915 (
		_w2229_,
		_w2230_,
		_w3112_,
		_w3144_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name916 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h2)
	) name917 (
		_w2999_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		_w2562_,
		_w3013_,
		_w3147_
	);
	LUT3 #(
		.INIT('h80)
	) name919 (
		_w2424_,
		_w2535_,
		_w2549_,
		_w3148_
	);
	LUT3 #(
		.INIT('h80)
	) name920 (
		_w3059_,
		_w3104_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3145_,
		_w3150_
	);
	LUT4 #(
		.INIT('ha222)
	) name922 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		_w2549_,
		_w3120_,
		_w3151_
	);
	LUT3 #(
		.INIT('hd0)
	) name923 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3145_,
		_w3151_,
		_w3152_
	);
	LUT4 #(
		.INIT('habaa)
	) name924 (
		_w3146_,
		_w3147_,
		_w3149_,
		_w3152_,
		_w3153_
	);
	LUT3 #(
		.INIT('h80)
	) name925 (
		_w2230_,
		_w2244_,
		_w2991_,
		_w3154_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name926 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h2)
	) name927 (
		_w2999_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w2556_,
		_w3013_,
		_w3157_
	);
	LUT3 #(
		.INIT('h80)
	) name929 (
		_w2424_,
		_w2511_,
		_w2534_,
		_w3158_
	);
	LUT3 #(
		.INIT('h80)
	) name930 (
		_w3059_,
		_w3104_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3155_,
		_w3160_
	);
	LUT4 #(
		.INIT('ha222)
	) name932 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		_w2534_,
		_w3108_,
		_w3161_
	);
	LUT3 #(
		.INIT('hd0)
	) name933 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3155_,
		_w3161_,
		_w3162_
	);
	LUT4 #(
		.INIT('habaa)
	) name934 (
		_w3156_,
		_w3157_,
		_w3159_,
		_w3162_,
		_w3163_
	);
	LUT3 #(
		.INIT('h80)
	) name935 (
		_w2230_,
		_w2244_,
		_w3112_,
		_w3164_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name936 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name937 (
		_w2999_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		_w2536_,
		_w3013_,
		_w3167_
	);
	LUT3 #(
		.INIT('h80)
	) name939 (
		_w2424_,
		_w2534_,
		_w2535_,
		_w3168_
	);
	LUT3 #(
		.INIT('h80)
	) name940 (
		_w3059_,
		_w3104_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3165_,
		_w3170_
	);
	LUT4 #(
		.INIT('ha222)
	) name942 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2534_,
		_w3120_,
		_w3171_
	);
	LUT3 #(
		.INIT('hd0)
	) name943 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3165_,
		_w3171_,
		_w3172_
	);
	LUT4 #(
		.INIT('habaa)
	) name944 (
		_w3166_,
		_w3167_,
		_w3169_,
		_w3172_,
		_w3173_
	);
	LUT3 #(
		.INIT('h80)
	) name945 (
		_w2229_,
		_w2230_,
		_w2991_,
		_w3174_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name946 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2993_,
		_w2994_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h2)
	) name947 (
		_w2999_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w2550_,
		_w3013_,
		_w3177_
	);
	LUT3 #(
		.INIT('h80)
	) name949 (
		_w2424_,
		_w2511_,
		_w2549_,
		_w3178_
	);
	LUT3 #(
		.INIT('h80)
	) name950 (
		_w3059_,
		_w3104_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3175_,
		_w3180_
	);
	LUT4 #(
		.INIT('ha222)
	) name952 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		_w2549_,
		_w3108_,
		_w3181_
	);
	LUT3 #(
		.INIT('hd0)
	) name953 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3175_,
		_w3181_,
		_w3182_
	);
	LUT4 #(
		.INIT('habaa)
	) name954 (
		_w3176_,
		_w3177_,
		_w3179_,
		_w3182_,
		_w3183_
	);
	LUT3 #(
		.INIT('h2a)
	) name955 (
		\ctl_rf_c1_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3184_
	);
	LUT3 #(
		.INIT('h80)
	) name956 (
		\ctl_rf_c2_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3185_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name957 (
		_w2514_,
		_w2518_,
		_w3184_,
		_w3185_,
		_w3186_
	);
	LUT3 #(
		.INIT('h2a)
	) name958 (
		\ctl_rf_c7_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3187_
	);
	LUT3 #(
		.INIT('h80)
	) name959 (
		\ctl_rf_c0_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3188_
	);
	LUT4 #(
		.INIT('h67ef)
	) name960 (
		_w2514_,
		_w2518_,
		_w3187_,
		_w3188_,
		_w3189_
	);
	LUT3 #(
		.INIT('h2a)
	) name961 (
		\ctl_rf_c3_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3190_
	);
	LUT3 #(
		.INIT('h80)
	) name962 (
		\ctl_rf_c6_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3191_
	);
	LUT4 #(
		.INIT('haebf)
	) name963 (
		_w2514_,
		_w2518_,
		_w3190_,
		_w3191_,
		_w3192_
	);
	LUT3 #(
		.INIT('h80)
	) name964 (
		\ctl_rf_c4_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3193_
	);
	LUT3 #(
		.INIT('h2a)
	) name965 (
		\ctl_rf_c5_rf_chtsz_reg[2]/P0002 ,
		_w2507_,
		_w2508_,
		_w3194_
	);
	LUT3 #(
		.INIT('h57)
	) name966 (
		_w2520_,
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h8000)
	) name967 (
		_w3186_,
		_w3189_,
		_w3192_,
		_w3195_,
		_w3196_
	);
	LUT4 #(
		.INIT('h7fff)
	) name968 (
		_w3186_,
		_w3189_,
		_w3192_,
		_w3195_,
		_w3197_
	);
	LUT3 #(
		.INIT('h2a)
	) name969 (
		\ctl_rf_c1_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3198_
	);
	LUT3 #(
		.INIT('h80)
	) name970 (
		\ctl_rf_c2_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3199_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name971 (
		_w2514_,
		_w2518_,
		_w3198_,
		_w3199_,
		_w3200_
	);
	LUT3 #(
		.INIT('h2a)
	) name972 (
		\ctl_rf_c7_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3201_
	);
	LUT3 #(
		.INIT('h80)
	) name973 (
		\ctl_rf_c0_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3202_
	);
	LUT4 #(
		.INIT('h67ef)
	) name974 (
		_w2514_,
		_w2518_,
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h2a)
	) name975 (
		\ctl_rf_c3_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3204_
	);
	LUT3 #(
		.INIT('h80)
	) name976 (
		\ctl_rf_c6_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3205_
	);
	LUT4 #(
		.INIT('haebf)
	) name977 (
		_w2514_,
		_w2518_,
		_w3204_,
		_w3205_,
		_w3206_
	);
	LUT3 #(
		.INIT('h80)
	) name978 (
		\ctl_rf_c4_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3207_
	);
	LUT3 #(
		.INIT('h2a)
	) name979 (
		\ctl_rf_c5_rf_chtsz_reg[4]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3208_
	);
	LUT3 #(
		.INIT('h57)
	) name980 (
		_w2520_,
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('h8000)
	) name981 (
		_w3200_,
		_w3203_,
		_w3206_,
		_w3209_,
		_w3210_
	);
	LUT4 #(
		.INIT('h7fff)
	) name982 (
		_w3200_,
		_w3203_,
		_w3206_,
		_w3209_,
		_w3211_
	);
	LUT3 #(
		.INIT('h2a)
	) name983 (
		\ctl_rf_c1_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3212_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		\ctl_rf_c2_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3213_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name985 (
		_w2514_,
		_w2518_,
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT3 #(
		.INIT('h2a)
	) name986 (
		\ctl_rf_c7_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3215_
	);
	LUT3 #(
		.INIT('h80)
	) name987 (
		\ctl_rf_c0_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3216_
	);
	LUT4 #(
		.INIT('h67ef)
	) name988 (
		_w2514_,
		_w2518_,
		_w3215_,
		_w3216_,
		_w3217_
	);
	LUT3 #(
		.INIT('h2a)
	) name989 (
		\ctl_rf_c3_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3218_
	);
	LUT3 #(
		.INIT('h80)
	) name990 (
		\ctl_rf_c6_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3219_
	);
	LUT4 #(
		.INIT('haebf)
	) name991 (
		_w2514_,
		_w2518_,
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT3 #(
		.INIT('h80)
	) name992 (
		\ctl_rf_c4_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3221_
	);
	LUT3 #(
		.INIT('h2a)
	) name993 (
		\ctl_rf_c5_rf_chtsz_reg[1]/P0002 ,
		_w2507_,
		_w2508_,
		_w3222_
	);
	LUT3 #(
		.INIT('h57)
	) name994 (
		_w2520_,
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT4 #(
		.INIT('h8000)
	) name995 (
		_w3214_,
		_w3217_,
		_w3220_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('h7fff)
	) name996 (
		_w3214_,
		_w3217_,
		_w3220_,
		_w3223_,
		_w3225_
	);
	LUT3 #(
		.INIT('h2a)
	) name997 (
		\ctl_rf_c1_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3226_
	);
	LUT3 #(
		.INIT('h80)
	) name998 (
		\ctl_rf_c2_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3227_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name999 (
		_w2514_,
		_w2518_,
		_w3226_,
		_w3227_,
		_w3228_
	);
	LUT3 #(
		.INIT('h2a)
	) name1000 (
		\ctl_rf_c7_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3229_
	);
	LUT3 #(
		.INIT('h80)
	) name1001 (
		\ctl_rf_c0_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3230_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1002 (
		_w2514_,
		_w2518_,
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT3 #(
		.INIT('h2a)
	) name1003 (
		\ctl_rf_c3_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3232_
	);
	LUT3 #(
		.INIT('h80)
	) name1004 (
		\ctl_rf_c6_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3233_
	);
	LUT4 #(
		.INIT('haebf)
	) name1005 (
		_w2514_,
		_w2518_,
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT3 #(
		.INIT('h80)
	) name1006 (
		\ctl_rf_c4_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3235_
	);
	LUT3 #(
		.INIT('h2a)
	) name1007 (
		\ctl_rf_c5_rf_chtsz_reg[11]/P0002 ,
		_w2507_,
		_w2508_,
		_w3236_
	);
	LUT3 #(
		.INIT('h57)
	) name1008 (
		_w2520_,
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('h8000)
	) name1009 (
		_w3228_,
		_w3231_,
		_w3234_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1010 (
		_w3228_,
		_w3231_,
		_w3234_,
		_w3237_,
		_w3239_
	);
	LUT4 #(
		.INIT('h8000)
	) name1011 (
		_w3196_,
		_w3210_,
		_w3224_,
		_w3238_,
		_w3240_
	);
	LUT3 #(
		.INIT('h2a)
	) name1012 (
		\ctl_rf_c1_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3241_
	);
	LUT3 #(
		.INIT('h80)
	) name1013 (
		\ctl_rf_c2_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3242_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1014 (
		_w2514_,
		_w2518_,
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT3 #(
		.INIT('h2a)
	) name1015 (
		\ctl_rf_c7_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3244_
	);
	LUT3 #(
		.INIT('h80)
	) name1016 (
		\ctl_rf_c0_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3245_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1017 (
		_w2514_,
		_w2518_,
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT3 #(
		.INIT('h2a)
	) name1018 (
		\ctl_rf_c3_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3247_
	);
	LUT3 #(
		.INIT('h80)
	) name1019 (
		\ctl_rf_c6_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3248_
	);
	LUT4 #(
		.INIT('haebf)
	) name1020 (
		_w2514_,
		_w2518_,
		_w3247_,
		_w3248_,
		_w3249_
	);
	LUT3 #(
		.INIT('h80)
	) name1021 (
		\ctl_rf_c4_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3250_
	);
	LUT3 #(
		.INIT('h2a)
	) name1022 (
		\ctl_rf_c5_rf_chtsz_reg[5]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3251_
	);
	LUT3 #(
		.INIT('h57)
	) name1023 (
		_w2520_,
		_w3250_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('h8000)
	) name1024 (
		_w3243_,
		_w3246_,
		_w3249_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1025 (
		_w3243_,
		_w3246_,
		_w3249_,
		_w3252_,
		_w3254_
	);
	LUT3 #(
		.INIT('h2a)
	) name1026 (
		\ctl_rf_c7_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3255_
	);
	LUT3 #(
		.INIT('h2a)
	) name1027 (
		\ctl_rf_c3_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3256_
	);
	LUT4 #(
		.INIT('habef)
	) name1028 (
		_w2514_,
		_w2518_,
		_w3255_,
		_w3256_,
		_w3257_
	);
	LUT3 #(
		.INIT('h2a)
	) name1029 (
		\ctl_rf_c1_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3258_
	);
	LUT3 #(
		.INIT('h80)
	) name1030 (
		\ctl_rf_c0_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3259_
	);
	LUT3 #(
		.INIT('h57)
	) name1031 (
		_w2549_,
		_w3258_,
		_w3259_,
		_w3260_
	);
	LUT3 #(
		.INIT('h80)
	) name1032 (
		\ctl_rf_c2_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3261_
	);
	LUT3 #(
		.INIT('h80)
	) name1033 (
		\ctl_rf_c6_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3262_
	);
	LUT4 #(
		.INIT('haebf)
	) name1034 (
		_w2514_,
		_w2518_,
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h80)
	) name1035 (
		\ctl_rf_c4_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3264_
	);
	LUT3 #(
		.INIT('h2a)
	) name1036 (
		\ctl_rf_c5_rf_chllpen_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w3265_
	);
	LUT3 #(
		.INIT('h57)
	) name1037 (
		_w2520_,
		_w3264_,
		_w3265_,
		_w3266_
	);
	LUT4 #(
		.INIT('h8000)
	) name1038 (
		_w3257_,
		_w3260_,
		_w3263_,
		_w3266_,
		_w3267_
	);
	LUT3 #(
		.INIT('h2a)
	) name1039 (
		\ctl_rf_c1_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3268_
	);
	LUT3 #(
		.INIT('h80)
	) name1040 (
		\ctl_rf_c2_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3269_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1041 (
		_w2514_,
		_w2518_,
		_w3268_,
		_w3269_,
		_w3270_
	);
	LUT3 #(
		.INIT('h2a)
	) name1042 (
		\ctl_rf_c7_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3271_
	);
	LUT3 #(
		.INIT('h80)
	) name1043 (
		\ctl_rf_c0_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3272_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1044 (
		_w2514_,
		_w2518_,
		_w3271_,
		_w3272_,
		_w3273_
	);
	LUT3 #(
		.INIT('h2a)
	) name1045 (
		\ctl_rf_c3_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3274_
	);
	LUT3 #(
		.INIT('h80)
	) name1046 (
		\ctl_rf_c6_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3275_
	);
	LUT4 #(
		.INIT('haebf)
	) name1047 (
		_w2514_,
		_w2518_,
		_w3274_,
		_w3275_,
		_w3276_
	);
	LUT3 #(
		.INIT('h80)
	) name1048 (
		\ctl_rf_c4_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3277_
	);
	LUT3 #(
		.INIT('h2a)
	) name1049 (
		\ctl_rf_c5_rf_chtsz_reg[3]/P0002 ,
		_w2507_,
		_w2508_,
		_w3278_
	);
	LUT3 #(
		.INIT('h57)
	) name1050 (
		_w2520_,
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT4 #(
		.INIT('h8000)
	) name1051 (
		_w3270_,
		_w3273_,
		_w3276_,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1052 (
		_w3270_,
		_w3273_,
		_w3276_,
		_w3279_,
		_w3281_
	);
	LUT3 #(
		.INIT('h2a)
	) name1053 (
		\ctl_rf_c1_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3282_
	);
	LUT3 #(
		.INIT('h80)
	) name1054 (
		\ctl_rf_c2_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3283_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1055 (
		_w2514_,
		_w2518_,
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT3 #(
		.INIT('h2a)
	) name1056 (
		\ctl_rf_c7_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3285_
	);
	LUT3 #(
		.INIT('h80)
	) name1057 (
		\ctl_rf_c0_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3286_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1058 (
		_w2514_,
		_w2518_,
		_w3285_,
		_w3286_,
		_w3287_
	);
	LUT3 #(
		.INIT('h2a)
	) name1059 (
		\ctl_rf_c3_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3288_
	);
	LUT3 #(
		.INIT('h80)
	) name1060 (
		\ctl_rf_c6_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3289_
	);
	LUT4 #(
		.INIT('haebf)
	) name1061 (
		_w2514_,
		_w2518_,
		_w3288_,
		_w3289_,
		_w3290_
	);
	LUT3 #(
		.INIT('h80)
	) name1062 (
		\ctl_rf_c4_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3291_
	);
	LUT3 #(
		.INIT('h2a)
	) name1063 (
		\ctl_rf_c5_rf_chtsz_reg[8]/P0002 ,
		_w2507_,
		_w2508_,
		_w3292_
	);
	LUT3 #(
		.INIT('h57)
	) name1064 (
		_w2520_,
		_w3291_,
		_w3292_,
		_w3293_
	);
	LUT4 #(
		.INIT('h8000)
	) name1065 (
		_w3284_,
		_w3287_,
		_w3290_,
		_w3293_,
		_w3294_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1066 (
		_w3284_,
		_w3287_,
		_w3290_,
		_w3293_,
		_w3295_
	);
	LUT4 #(
		.INIT('h8000)
	) name1067 (
		_w3253_,
		_w3267_,
		_w3280_,
		_w3294_,
		_w3296_
	);
	LUT3 #(
		.INIT('h2a)
	) name1068 (
		\ctl_rf_c1_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3297_
	);
	LUT3 #(
		.INIT('h80)
	) name1069 (
		\ctl_rf_c2_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3298_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1070 (
		_w2514_,
		_w2518_,
		_w3297_,
		_w3298_,
		_w3299_
	);
	LUT3 #(
		.INIT('h2a)
	) name1071 (
		\ctl_rf_c7_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3300_
	);
	LUT3 #(
		.INIT('h80)
	) name1072 (
		\ctl_rf_c0_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3301_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1073 (
		_w2514_,
		_w2518_,
		_w3300_,
		_w3301_,
		_w3302_
	);
	LUT3 #(
		.INIT('h2a)
	) name1074 (
		\ctl_rf_c3_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3303_
	);
	LUT3 #(
		.INIT('h80)
	) name1075 (
		\ctl_rf_c6_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3304_
	);
	LUT4 #(
		.INIT('haebf)
	) name1076 (
		_w2514_,
		_w2518_,
		_w3303_,
		_w3304_,
		_w3305_
	);
	LUT3 #(
		.INIT('h80)
	) name1077 (
		\ctl_rf_c4_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3306_
	);
	LUT3 #(
		.INIT('h2a)
	) name1078 (
		\ctl_rf_c5_rf_chtsz_reg[7]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3307_
	);
	LUT3 #(
		.INIT('h57)
	) name1079 (
		_w2520_,
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h8000)
	) name1080 (
		_w3299_,
		_w3302_,
		_w3305_,
		_w3308_,
		_w3309_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1081 (
		_w3299_,
		_w3302_,
		_w3305_,
		_w3308_,
		_w3310_
	);
	LUT3 #(
		.INIT('h2a)
	) name1082 (
		\ctl_rf_c1_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3311_
	);
	LUT3 #(
		.INIT('h80)
	) name1083 (
		\ctl_rf_c2_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3312_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1084 (
		_w2514_,
		_w2518_,
		_w3311_,
		_w3312_,
		_w3313_
	);
	LUT3 #(
		.INIT('h2a)
	) name1085 (
		\ctl_rf_c7_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3314_
	);
	LUT3 #(
		.INIT('h80)
	) name1086 (
		\ctl_rf_c0_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3315_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1087 (
		_w2514_,
		_w2518_,
		_w3314_,
		_w3315_,
		_w3316_
	);
	LUT3 #(
		.INIT('h2a)
	) name1088 (
		\ctl_rf_c3_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3317_
	);
	LUT3 #(
		.INIT('h80)
	) name1089 (
		\ctl_rf_c6_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3318_
	);
	LUT4 #(
		.INIT('haebf)
	) name1090 (
		_w2514_,
		_w2518_,
		_w3317_,
		_w3318_,
		_w3319_
	);
	LUT3 #(
		.INIT('h80)
	) name1091 (
		\ctl_rf_c4_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3320_
	);
	LUT3 #(
		.INIT('h2a)
	) name1092 (
		\ctl_rf_c5_rf_chtsz_reg[9]/P0002 ,
		_w2507_,
		_w2508_,
		_w3321_
	);
	LUT3 #(
		.INIT('h57)
	) name1093 (
		_w2520_,
		_w3320_,
		_w3321_,
		_w3322_
	);
	LUT4 #(
		.INIT('h8000)
	) name1094 (
		_w3313_,
		_w3316_,
		_w3319_,
		_w3322_,
		_w3323_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1095 (
		_w3313_,
		_w3316_,
		_w3319_,
		_w3322_,
		_w3324_
	);
	LUT3 #(
		.INIT('h2a)
	) name1096 (
		\ctl_rf_c1_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3325_
	);
	LUT3 #(
		.INIT('h80)
	) name1097 (
		\ctl_rf_c2_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3326_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1098 (
		_w2514_,
		_w2518_,
		_w3325_,
		_w3326_,
		_w3327_
	);
	LUT3 #(
		.INIT('h2a)
	) name1099 (
		\ctl_rf_c7_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3328_
	);
	LUT3 #(
		.INIT('h80)
	) name1100 (
		\ctl_rf_c0_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3329_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1101 (
		_w2514_,
		_w2518_,
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT3 #(
		.INIT('h2a)
	) name1102 (
		\ctl_rf_c3_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3331_
	);
	LUT3 #(
		.INIT('h80)
	) name1103 (
		\ctl_rf_c6_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3332_
	);
	LUT4 #(
		.INIT('haebf)
	) name1104 (
		_w2514_,
		_w2518_,
		_w3331_,
		_w3332_,
		_w3333_
	);
	LUT3 #(
		.INIT('h80)
	) name1105 (
		\ctl_rf_c4_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3334_
	);
	LUT3 #(
		.INIT('h2a)
	) name1106 (
		\ctl_rf_c5_rf_chtsz_reg[10]/P0002 ,
		_w2507_,
		_w2508_,
		_w3335_
	);
	LUT3 #(
		.INIT('h57)
	) name1107 (
		_w2520_,
		_w3334_,
		_w3335_,
		_w3336_
	);
	LUT4 #(
		.INIT('h8000)
	) name1108 (
		_w3327_,
		_w3330_,
		_w3333_,
		_w3336_,
		_w3337_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1109 (
		_w3327_,
		_w3330_,
		_w3333_,
		_w3336_,
		_w3338_
	);
	LUT3 #(
		.INIT('h2a)
	) name1110 (
		\ctl_rf_c1_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3339_
	);
	LUT3 #(
		.INIT('h80)
	) name1111 (
		\ctl_rf_c2_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3340_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1112 (
		_w2514_,
		_w2518_,
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT3 #(
		.INIT('h2a)
	) name1113 (
		\ctl_rf_c7_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3342_
	);
	LUT3 #(
		.INIT('h80)
	) name1114 (
		\ctl_rf_c0_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3343_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1115 (
		_w2514_,
		_w2518_,
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT3 #(
		.INIT('h2a)
	) name1116 (
		\ctl_rf_c3_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3345_
	);
	LUT3 #(
		.INIT('h80)
	) name1117 (
		\ctl_rf_c6_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3346_
	);
	LUT4 #(
		.INIT('haebf)
	) name1118 (
		_w2514_,
		_w2518_,
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT3 #(
		.INIT('h80)
	) name1119 (
		\ctl_rf_c4_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3348_
	);
	LUT3 #(
		.INIT('h2a)
	) name1120 (
		\ctl_rf_c5_rf_chtsz_reg[6]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3349_
	);
	LUT3 #(
		.INIT('h57)
	) name1121 (
		_w2520_,
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h8000)
	) name1122 (
		_w3341_,
		_w3344_,
		_w3347_,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1123 (
		_w3341_,
		_w3344_,
		_w3347_,
		_w3350_,
		_w3352_
	);
	LUT4 #(
		.INIT('h8000)
	) name1124 (
		_w3309_,
		_w3323_,
		_w3337_,
		_w3351_,
		_w3353_
	);
	LUT3 #(
		.INIT('h01)
	) name1125 (
		\de_de_st_reg[2]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		_w3354_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		\de_de_st_reg[0]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT3 #(
		.INIT('h2a)
	) name1128 (
		\ctl_rf_c1_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3357_
	);
	LUT3 #(
		.INIT('h80)
	) name1129 (
		\ctl_rf_c2_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3358_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name1130 (
		_w2514_,
		_w2518_,
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT3 #(
		.INIT('h2a)
	) name1131 (
		\ctl_rf_c7_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3360_
	);
	LUT3 #(
		.INIT('h80)
	) name1132 (
		\ctl_rf_c0_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3361_
	);
	LUT4 #(
		.INIT('h67ef)
	) name1133 (
		_w2514_,
		_w2518_,
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT3 #(
		.INIT('h2a)
	) name1134 (
		\ctl_rf_c3_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3363_
	);
	LUT3 #(
		.INIT('h80)
	) name1135 (
		\ctl_rf_c6_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3364_
	);
	LUT4 #(
		.INIT('haebf)
	) name1136 (
		_w2514_,
		_w2518_,
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('h80)
	) name1137 (
		\ctl_rf_c4_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3366_
	);
	LUT3 #(
		.INIT('h2a)
	) name1138 (
		\ctl_rf_c5_rf_chtsz_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w3367_
	);
	LUT3 #(
		.INIT('h57)
	) name1139 (
		_w2520_,
		_w3366_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('h8000)
	) name1140 (
		_w3359_,
		_w3362_,
		_w3365_,
		_w3368_,
		_w3369_
	);
	LUT4 #(
		.INIT('h7fff)
	) name1141 (
		_w3359_,
		_w3362_,
		_w3365_,
		_w3368_,
		_w3370_
	);
	LUT4 #(
		.INIT('ha222)
	) name1142 (
		\ch_sel_arb_req_reg/NET0131 ,
		\de_de_st_reg[0]/NET0131 ,
		_w2575_,
		_w2576_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name1143 (
		_w3369_,
		_w3371_,
		_w3372_
	);
	LUT3 #(
		.INIT('h80)
	) name1144 (
		_w3356_,
		_w3369_,
		_w3371_,
		_w3373_
	);
	LUT4 #(
		.INIT('h8000)
	) name1145 (
		_w3240_,
		_w3296_,
		_w3353_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h6)
	) name1146 (
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name1147 (
		\de_tsz_cnt_reg[0]/NET0131 ,
		\de_tsz_cnt_reg[1]/NET0131 ,
		_w3376_
	);
	LUT4 #(
		.INIT('h8000)
	) name1148 (
		_w2420_,
		_w2421_,
		_w2422_,
		_w3376_,
		_w3377_
	);
	LUT4 #(
		.INIT('h0002)
	) name1149 (
		\de_bst_cnt_reg[0]/NET0131 ,
		\de_bst_cnt_reg[2]/NET0131 ,
		\de_bst_cnt_reg[3]/NET0131 ,
		\de_bst_cnt_reg[4]/NET0131 ,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		_w2426_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		\de_de_st_reg[0]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w3380_
	);
	LUT2 #(
		.INIT('h8)
	) name1152 (
		_w3354_,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('hab00)
	) name1153 (
		_w3375_,
		_w3377_,
		_w3379_,
		_w3381_,
		_w3382_
	);
	LUT3 #(
		.INIT('h8a)
	) name1154 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w2468_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1156 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w3384_,
		_w3385_
	);
	LUT2 #(
		.INIT('h8)
	) name1157 (
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\h0readyin_pad ,
		_w3386_
	);
	LUT4 #(
		.INIT('h0200)
	) name1158 (
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		\h0readyin_pad ,
		_w3387_
	);
	LUT3 #(
		.INIT('h08)
	) name1159 (
		_w3354_,
		_w3380_,
		_w3387_,
		_w3388_
	);
	LUT3 #(
		.INIT('h45)
	) name1160 (
		_w3382_,
		_w3385_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('h8000)
	) name1161 (
		_w3240_,
		_w3296_,
		_w3353_,
		_w3372_,
		_w3390_
	);
	LUT3 #(
		.INIT('h80)
	) name1162 (
		\ch_sel_arb_req_reg/NET0131 ,
		_w3354_,
		_w3355_,
		_w3391_
	);
	LUT2 #(
		.INIT('h4)
	) name1163 (
		_w2577_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		_w3267_,
		_w3392_,
		_w3393_
	);
	LUT3 #(
		.INIT('h75)
	) name1165 (
		_w3389_,
		_w3390_,
		_w3393_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		\ahb_mst0_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		_w3395_
	);
	LUT4 #(
		.INIT('h008f)
	) name1167 (
		_w2496_,
		_w2497_,
		_w2498_,
		_w3395_,
		_w3396_
	);
	LUT4 #(
		.INIT('h000d)
	) name1168 (
		\ahb_mst0_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w3397_
	);
	LUT4 #(
		.INIT('h010f)
	) name1169 (
		_w2471_,
		_w2494_,
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('h5510)
	) name1170 (
		\h0req_pad ,
		_w2424_,
		_w2485_,
		_w2486_,
		_w3399_
	);
	LUT3 #(
		.INIT('h20)
	) name1171 (
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w3400_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\de_de_st_reg[5]/NET0131 ,
		\h0req_pad ,
		_w3401_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT3 #(
		.INIT('h70)
	) name1174 (
		_w2426_,
		_w2427_,
		_w3401_,
		_w3403_
	);
	LUT3 #(
		.INIT('h23)
	) name1175 (
		_w2424_,
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('hb)
	) name1176 (
		_w3399_,
		_w3404_,
		_w3405_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		\de_de_st_reg[0]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w3406_
	);
	LUT3 #(
		.INIT('h02)
	) name1178 (
		\de_de_st_reg[2]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		_w3407_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT4 #(
		.INIT('h5400)
	) name1180 (
		_w3375_,
		_w3377_,
		_w3379_,
		_w3381_,
		_w3409_
	);
	LUT4 #(
		.INIT('hfef0)
	) name1181 (
		_w3385_,
		_w3387_,
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h8000)
	) name1182 (
		_w2889_,
		_w2890_,
		_w2891_,
		_w2893_,
		_w3411_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w2579_,
		_w3411_,
		_w3412_
	);
	LUT4 #(
		.INIT('h8000)
	) name1184 (
		_w2845_,
		_w2846_,
		_w2847_,
		_w2852_,
		_w3413_
	);
	LUT4 #(
		.INIT('h8000)
	) name1185 (
		_w2795_,
		_w2798_,
		_w2865_,
		_w2866_,
		_w3414_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		\ch_sel_fix_pri_sel_reg[0]/NET0131 ,
		_w2578_,
		_w3415_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1187 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w3415_,
		_w3416_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1188 (
		_w2579_,
		_w3413_,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('hb)
	) name1189 (
		_w3412_,
		_w3417_,
		_w3418_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		\ch_sel_fix_pri_sel_reg[1]/NET0131 ,
		_w2578_,
		_w3419_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1191 (
		_w2546_,
		_w2572_,
		_w2574_,
		_w3419_,
		_w3420_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1192 (
		_w2579_,
		_w3411_,
		_w3414_,
		_w3420_,
		_w3421_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3422_
	);
	LUT3 #(
		.INIT('h2a)
	) name1194 (
		\hrdata_reg[16]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3423_
	);
	LUT4 #(
		.INIT('h0008)
	) name1195 (
		\ctl_rf_m0end_reg/NET0131 ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w3424_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3425_
	);
	LUT4 #(
		.INIT('h0100)
	) name1197 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3426_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3427_
	);
	LUT4 #(
		.INIT('hff35)
	) name1199 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3428_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1200 (
		\ctl_rf_c4_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3429_
	);
	LUT3 #(
		.INIT('h2a)
	) name1201 (
		_w3426_,
		_w3428_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3431_
	);
	LUT4 #(
		.INIT('h0010)
	) name1203 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3432_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1204 (
		\ctl_rf_c2_rf_chsad_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3433_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1205 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chdad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3434_
	);
	LUT3 #(
		.INIT('h2a)
	) name1206 (
		_w3432_,
		_w3433_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('h0400)
	) name1207 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3436_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1208 (
		\ctl_rf_c5_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3437_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1209 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3438_
	);
	LUT3 #(
		.INIT('h2a)
	) name1210 (
		_w3436_,
		_w3437_,
		_w3438_,
		_w3439_
	);
	LUT4 #(
		.INIT('h1000)
	) name1211 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3440_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1212 (
		\ctl_rf_c6_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3441_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1213 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3442_
	);
	LUT3 #(
		.INIT('h2a)
	) name1214 (
		_w3440_,
		_w3441_,
		_w3442_,
		_w3443_
	);
	LUT4 #(
		.INIT('h0001)
	) name1215 (
		_w3430_,
		_w3435_,
		_w3439_,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('h0001)
	) name1216 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3445_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1217 (
		\ctl_rf_c0_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3446_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1218 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3447_
	);
	LUT3 #(
		.INIT('h2a)
	) name1219 (
		_w3445_,
		_w3446_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h0004)
	) name1220 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3449_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1221 (
		\ctl_rf_c1_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3450_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1222 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3451_
	);
	LUT3 #(
		.INIT('h2a)
	) name1223 (
		_w3449_,
		_w3450_,
		_w3451_,
		_w3452_
	);
	LUT4 #(
		.INIT('h4000)
	) name1224 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3453_
	);
	LUT4 #(
		.INIT('hff35)
	) name1225 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3454_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1226 (
		\ctl_rf_c7_rf_chdad_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3455_
	);
	LUT3 #(
		.INIT('h2a)
	) name1227 (
		_w3453_,
		_w3454_,
		_w3455_,
		_w3456_
	);
	LUT4 #(
		.INIT('h0040)
	) name1228 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3457_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1229 (
		\ctl_rf_c3_rf_chsad_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3458_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1230 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chdad_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3459_
	);
	LUT3 #(
		.INIT('h2a)
	) name1231 (
		_w3457_,
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h0001)
	) name1232 (
		_w3448_,
		_w3452_,
		_w3456_,
		_w3460_,
		_w3461_
	);
	LUT4 #(
		.INIT('h0020)
	) name1233 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3462_
	);
	LUT4 #(
		.INIT('hff35)
	) name1234 (
		\ctl_rf_c2_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c2_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3463_
	);
	LUT4 #(
		.INIT('h8000)
	) name1235 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3464_
	);
	LUT4 #(
		.INIT('hff35)
	) name1236 (
		\ctl_rf_c7_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c7_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3465_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1237 (
		_w3462_,
		_w3463_,
		_w3464_,
		_w3465_,
		_w3466_
	);
	LUT4 #(
		.INIT('h0002)
	) name1238 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3467_
	);
	LUT4 #(
		.INIT('hff35)
	) name1239 (
		\ctl_rf_c0_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c0_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3468_
	);
	LUT4 #(
		.INIT('h0800)
	) name1240 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3469_
	);
	LUT4 #(
		.INIT('hff35)
	) name1241 (
		\ctl_rf_c5_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c5_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3470_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1242 (
		_w3467_,
		_w3468_,
		_w3469_,
		_w3470_,
		_w3471_
	);
	LUT4 #(
		.INIT('h0200)
	) name1243 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3472_
	);
	LUT4 #(
		.INIT('hff35)
	) name1244 (
		\ctl_rf_c4_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c4_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3473_
	);
	LUT4 #(
		.INIT('h0008)
	) name1245 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3474_
	);
	LUT4 #(
		.INIT('hff35)
	) name1246 (
		\ctl_rf_c1_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c1_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3475_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1247 (
		_w3472_,
		_w3473_,
		_w3474_,
		_w3475_,
		_w3476_
	);
	LUT4 #(
		.INIT('h0080)
	) name1248 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3477_
	);
	LUT4 #(
		.INIT('hff35)
	) name1249 (
		\ctl_rf_c3_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c3_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3478_
	);
	LUT4 #(
		.INIT('h2000)
	) name1250 (
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		_w3479_
	);
	LUT4 #(
		.INIT('hff35)
	) name1251 (
		\ctl_rf_c6_rf_chllp_reg[0]/P0002 ,
		\ctl_rf_c6_rf_chtsz_reg[0]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3480_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1252 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h8000)
	) name1253 (
		_w3466_,
		_w3471_,
		_w3476_,
		_w3481_,
		_w3482_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1254 (
		\haddr[8]_pad ,
		_w3444_,
		_w3461_,
		_w3482_,
		_w3483_
	);
	LUT3 #(
		.INIT('h01)
	) name1255 (
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w3484_
	);
	LUT4 #(
		.INIT('h0100)
	) name1256 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3485_
	);
	LUT4 #(
		.INIT('h4000)
	) name1257 (
		\de_de_st_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		_w2549_,
		_w3486_,
		_w3487_
	);
	LUT4 #(
		.INIT('h0020)
	) name1259 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3488_
	);
	LUT3 #(
		.INIT('h01)
	) name1260 (
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3489_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name1261 (
		\ctl_rf_c0_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[0]/NET0131 ,
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT4 #(
		.INIT('h0400)
	) name1262 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3491_
	);
	LUT4 #(
		.INIT('h0080)
	) name1263 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3492_
	);
	LUT4 #(
		.INIT('h153f)
	) name1264 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[0]/NET0131 ,
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT4 #(
		.INIT('h0200)
	) name1265 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3494_
	);
	LUT2 #(
		.INIT('h2)
	) name1266 (
		\ctl_rf_abt_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_int_abt_msk_reg/NET0131 ,
		_w3495_
	);
	LUT4 #(
		.INIT('h0001)
	) name1267 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3496_
	);
	LUT4 #(
		.INIT('h0777)
	) name1268 (
		\ctl_rf_dmacen_reg/NET0131 ,
		_w3494_,
		_w3495_,
		_w3496_,
		_w3497_
	);
	LUT3 #(
		.INIT('h80)
	) name1269 (
		_w3490_,
		_w3493_,
		_w3497_,
		_w3498_
	);
	LUT3 #(
		.INIT('h8a)
	) name1270 (
		_w3484_,
		_w3487_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h2a22)
	) name1271 (
		_w3424_,
		_w3484_,
		_w3487_,
		_w3498_,
		_w3500_
	);
	LUT3 #(
		.INIT('h8a)
	) name1272 (
		_w3422_,
		_w3483_,
		_w3500_,
		_w3501_
	);
	LUT4 #(
		.INIT('h8880)
	) name1273 (
		_w3422_,
		_w3424_,
		_w3483_,
		_w3499_,
		_w3502_
	);
	LUT4 #(
		.INIT('h0002)
	) name1274 (
		\ctl_rf_m0end_reg/NET0131 ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w3503_
	);
	LUT2 #(
		.INIT('h4)
	) name1275 (
		\haddr[8]_pad ,
		_w3503_,
		_w3504_
	);
	LUT3 #(
		.INIT('h04)
	) name1276 (
		\de_de_st_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3505_
	);
	LUT3 #(
		.INIT('h70)
	) name1277 (
		_w2507_,
		_w2508_,
		_w3505_,
		_w3506_
	);
	LUT3 #(
		.INIT('h20)
	) name1278 (
		\ctl_rf_c7_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3507_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1279 (
		\ctl_rf_c7_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c7_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3508_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1281 (
		_w2527_,
		_w3453_,
		_w3506_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('hff35)
	) name1282 (
		\ctl_rf_c6_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3511_
	);
	LUT4 #(
		.INIT('hff35)
	) name1283 (
		\ctl_rf_c3_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3512_
	);
	LUT4 #(
		.INIT('hf351)
	) name1284 (
		_w3477_,
		_w3479_,
		_w3511_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('hff35)
	) name1285 (
		\ctl_rf_c7_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3514_
	);
	LUT4 #(
		.INIT('hff35)
	) name1286 (
		\ctl_rf_c4_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3515_
	);
	LUT4 #(
		.INIT('hf531)
	) name1287 (
		_w3464_,
		_w3472_,
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT4 #(
		.INIT('hff35)
	) name1288 (
		\ctl_rf_c2_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3517_
	);
	LUT4 #(
		.INIT('hff35)
	) name1289 (
		\ctl_rf_c0_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3518_
	);
	LUT4 #(
		.INIT('hf531)
	) name1290 (
		_w3462_,
		_w3467_,
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('hff35)
	) name1291 (
		\ctl_rf_c1_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3520_
	);
	LUT4 #(
		.INIT('hff35)
	) name1292 (
		\ctl_rf_c5_rf_chllp_reg[8]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3521_
	);
	LUT4 #(
		.INIT('hf351)
	) name1293 (
		_w3469_,
		_w3474_,
		_w3520_,
		_w3521_,
		_w3522_
	);
	LUT4 #(
		.INIT('h8000)
	) name1294 (
		_w3513_,
		_w3516_,
		_w3519_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		_w3510_,
		_w3523_,
		_w3524_
	);
	LUT3 #(
		.INIT('h80)
	) name1296 (
		_w2507_,
		_w2508_,
		_w3505_,
		_w3525_
	);
	LUT3 #(
		.INIT('h20)
	) name1297 (
		\ctl_rf_c6_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3526_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1298 (
		\ctl_rf_c6_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c6_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3527_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1300 (
		_w2527_,
		_w3440_,
		_w3525_,
		_w3528_,
		_w3529_
	);
	LUT3 #(
		.INIT('h20)
	) name1301 (
		\ctl_rf_c1_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3530_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1302 (
		\ctl_rf_c1_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c1_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3531_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		_w3530_,
		_w3531_,
		_w3532_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1304 (
		_w2549_,
		_w3449_,
		_w3506_,
		_w3532_,
		_w3533_
	);
	LUT3 #(
		.INIT('h20)
	) name1305 (
		\ctl_rf_c5_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3534_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1306 (
		\ctl_rf_c5_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c5_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3535_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w3534_,
		_w3535_,
		_w3536_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1308 (
		_w2520_,
		_w3436_,
		_w3506_,
		_w3536_,
		_w3537_
	);
	LUT3 #(
		.INIT('h20)
	) name1309 (
		\ctl_rf_c2_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3538_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1310 (
		\ctl_rf_c2_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c2_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3539_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w3538_,
		_w3539_,
		_w3540_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1312 (
		_w2534_,
		_w3432_,
		_w3525_,
		_w3540_,
		_w3541_
	);
	LUT4 #(
		.INIT('h0001)
	) name1313 (
		_w3529_,
		_w3533_,
		_w3537_,
		_w3541_,
		_w3542_
	);
	LUT3 #(
		.INIT('h20)
	) name1314 (
		\ctl_rf_c0_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3543_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1315 (
		\ctl_rf_c0_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c0_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3544_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w3543_,
		_w3544_,
		_w3545_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1317 (
		_w2549_,
		_w3445_,
		_w3525_,
		_w3545_,
		_w3546_
	);
	LUT3 #(
		.INIT('h20)
	) name1318 (
		\ctl_rf_c3_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3547_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1319 (
		\ctl_rf_c3_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c3_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name1320 (
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1321 (
		_w2534_,
		_w3457_,
		_w3506_,
		_w3549_,
		_w3550_
	);
	LUT3 #(
		.INIT('h20)
	) name1322 (
		\ctl_rf_c4_rf_chsad_reg[8]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3551_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1323 (
		\ctl_rf_c4_rf_chdad_reg[8]/NET0131 ,
		\ctl_rf_c4_rf_dwidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3552_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w3551_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('h80cc)
	) name1325 (
		_w2520_,
		_w3426_,
		_w3525_,
		_w3553_,
		_w3554_
	);
	LUT4 #(
		.INIT('h0002)
	) name1326 (
		_w3503_,
		_w3546_,
		_w3550_,
		_w3554_,
		_w3555_
	);
	LUT4 #(
		.INIT('h1555)
	) name1327 (
		_w3504_,
		_w3524_,
		_w3542_,
		_w3555_,
		_w3556_
	);
	LUT4 #(
		.INIT('hff53)
	) name1328 (
		\ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3557_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1329 (
		\ctl_rf_c0_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c0_rf_chsad_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3558_
	);
	LUT4 #(
		.INIT('ha222)
	) name1330 (
		\haddr[8]_pad ,
		_w3445_,
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1331 (
		\ctl_rf_c2_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3560_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1332 (
		\ctl_rf_c2_rf_chsad_reg[16]/NET0131 ,
		\ctl_rf_c2_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3561_
	);
	LUT3 #(
		.INIT('h2a)
	) name1333 (
		_w3432_,
		_w3560_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1334 (
		\ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chsad_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3563_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1335 (
		\ctl_rf_c6_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c6_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3564_
	);
	LUT3 #(
		.INIT('h2a)
	) name1336 (
		_w3440_,
		_w3563_,
		_w3564_,
		_w3565_
	);
	LUT4 #(
		.INIT('hff53)
	) name1337 (
		\ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3566_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1338 (
		\ctl_rf_c1_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3567_
	);
	LUT3 #(
		.INIT('h2a)
	) name1339 (
		_w3449_,
		_w3566_,
		_w3567_,
		_w3568_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1340 (
		\ctl_rf_c7_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3569_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1341 (
		\ctl_rf_c7_rf_chsad_reg[16]/NET0131 ,
		\ctl_rf_c7_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3570_
	);
	LUT3 #(
		.INIT('h2a)
	) name1342 (
		_w3453_,
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT4 #(
		.INIT('h0001)
	) name1343 (
		_w3562_,
		_w3565_,
		_w3568_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		_w3559_,
		_w3572_,
		_w3573_
	);
	LUT4 #(
		.INIT('h135f)
	) name1345 (
		\ctl_rf_c1_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[16]/NET0131 ,
		_w3474_,
		_w3477_,
		_w3574_
	);
	LUT4 #(
		.INIT('h135f)
	) name1346 (
		\ctl_rf_c0_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[16]/NET0131 ,
		_w3467_,
		_w3472_,
		_w3575_
	);
	LUT4 #(
		.INIT('h135f)
	) name1347 (
		\ctl_rf_c5_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[16]/NET0131 ,
		_w3469_,
		_w3479_,
		_w3576_
	);
	LUT4 #(
		.INIT('h135f)
	) name1348 (
		\ctl_rf_c2_rf_chllp_reg[16]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[16]/NET0131 ,
		_w3462_,
		_w3464_,
		_w3577_
	);
	LUT4 #(
		.INIT('h8000)
	) name1349 (
		_w3574_,
		_w3575_,
		_w3576_,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1350 (
		\ctl_rf_c4_rf_chsad_reg[16]/NET0131 ,
		\ctl_rf_c4_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3579_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1351 (
		\ctl_rf_c4_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3580_
	);
	LUT3 #(
		.INIT('h2a)
	) name1352 (
		_w3426_,
		_w3579_,
		_w3580_,
		_w3581_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1353 (
		\ctl_rf_c5_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3582_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1354 (
		\ctl_rf_c5_rf_chsad_reg[16]/NET0131 ,
		\ctl_rf_c5_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3583_
	);
	LUT3 #(
		.INIT('h2a)
	) name1355 (
		_w3436_,
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1356 (
		\ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chsad_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3585_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1357 (
		\ctl_rf_c3_rf_chdad_reg[16]/NET0131 ,
		\ctl_rf_c3_rf_src_sz_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3586_
	);
	LUT3 #(
		.INIT('h2a)
	) name1358 (
		_w3457_,
		_w3585_,
		_w3586_,
		_w3587_
	);
	LUT3 #(
		.INIT('h01)
	) name1359 (
		_w3581_,
		_w3584_,
		_w3587_,
		_w3588_
	);
	LUT3 #(
		.INIT('hd0)
	) name1360 (
		_w3427_,
		_w3578_,
		_w3588_,
		_w3589_
	);
	LUT4 #(
		.INIT('h0200)
	) name1361 (
		\ctl_rf_c4dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3590_
	);
	LUT4 #(
		.INIT('h0800)
	) name1362 (
		\ctl_rf_c5dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3591_
	);
	LUT4 #(
		.INIT('h0002)
	) name1363 (
		\ctl_rf_c0dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3592_
	);
	LUT4 #(
		.INIT('h2000)
	) name1364 (
		\ctl_rf_c6dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3593_
	);
	LUT4 #(
		.INIT('h0001)
	) name1365 (
		_w3590_,
		_w3591_,
		_w3592_,
		_w3593_,
		_w3594_
	);
	LUT4 #(
		.INIT('h8000)
	) name1366 (
		\ctl_rf_c7dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3595_
	);
	LUT4 #(
		.INIT('h0020)
	) name1367 (
		\ctl_rf_c2dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3596_
	);
	LUT4 #(
		.INIT('h0008)
	) name1368 (
		\ctl_rf_c1dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3597_
	);
	LUT4 #(
		.INIT('h0080)
	) name1369 (
		\ctl_rf_c3dmabs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3598_
	);
	LUT4 #(
		.INIT('h0001)
	) name1370 (
		_w3595_,
		_w3596_,
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT3 #(
		.INIT('h2a)
	) name1371 (
		_w3431_,
		_w3594_,
		_w3599_,
		_w3600_
	);
	LUT4 #(
		.INIT('h0008)
	) name1372 (
		\ctl_rf_c1brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3601_
	);
	LUT4 #(
		.INIT('h0800)
	) name1373 (
		\ctl_rf_c5brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3602_
	);
	LUT4 #(
		.INIT('h0002)
	) name1374 (
		\ctl_rf_c0brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3603_
	);
	LUT4 #(
		.INIT('h8000)
	) name1375 (
		\ctl_rf_c7brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3604_
	);
	LUT4 #(
		.INIT('h0001)
	) name1376 (
		_w3601_,
		_w3602_,
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('h2000)
	) name1377 (
		\ctl_rf_c6brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3606_
	);
	LUT4 #(
		.INIT('h0020)
	) name1378 (
		\ctl_rf_c2brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3607_
	);
	LUT4 #(
		.INIT('h0200)
	) name1379 (
		\ctl_rf_c4brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3608_
	);
	LUT4 #(
		.INIT('h0080)
	) name1380 (
		\ctl_rf_c3brbs_reg[16]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3609_
	);
	LUT4 #(
		.INIT('h0001)
	) name1381 (
		_w3606_,
		_w3607_,
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT3 #(
		.INIT('h2a)
	) name1382 (
		_w3425_,
		_w3605_,
		_w3610_,
		_w3611_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1383 (
		\ctl_rf_abt_reg[0]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w3612_
	);
	LUT4 #(
		.INIT('h0008)
	) name1384 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3613_
	);
	LUT4 #(
		.INIT('h0040)
	) name1385 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		\haddr[5]_pad ,
		_w3614_
	);
	LUT4 #(
		.INIT('h0023)
	) name1386 (
		\ctl_rf_c0_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w3612_,
		_w3615_,
		_w3616_
	);
	LUT3 #(
		.INIT('h01)
	) name1388 (
		_w3600_,
		_w3611_,
		_w3616_,
		_w3617_
	);
	LUT4 #(
		.INIT('h5540)
	) name1389 (
		_w3503_,
		_w3573_,
		_w3589_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h3313)
	) name1390 (
		_w3501_,
		_w3502_,
		_w3556_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('hb)
	) name1391 (
		_w3423_,
		_w3619_,
		_w3620_
	);
	LUT3 #(
		.INIT('h2a)
	) name1392 (
		\hrdata_reg[8]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name1393 (
		_w3422_,
		_w3424_,
		_w3622_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\ctl_rf_c3_rf_chllp_reg[24]/NET0131 ,
		_w3477_,
		_w3623_
	);
	LUT4 #(
		.INIT('h135f)
	) name1395 (
		\ctl_rf_c2_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[24]/NET0131 ,
		_w3462_,
		_w3469_,
		_w3624_
	);
	LUT2 #(
		.INIT('h4)
	) name1396 (
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT4 #(
		.INIT('h135f)
	) name1397 (
		\ctl_rf_c0_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c1_rf_chllp_reg[24]/NET0131 ,
		_w3467_,
		_w3474_,
		_w3626_
	);
	LUT4 #(
		.INIT('h153f)
	) name1398 (
		\ctl_rf_c4_rf_chllp_reg[24]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[24]/NET0131 ,
		_w3464_,
		_w3472_,
		_w3627_
	);
	LUT4 #(
		.INIT('h135f)
	) name1399 (
		\ctl_rf_c1_rf_dreqmode_reg/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[24]/NET0131 ,
		_w3449_,
		_w3479_,
		_w3628_
	);
	LUT3 #(
		.INIT('h80)
	) name1400 (
		_w3626_,
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT3 #(
		.INIT('h2a)
	) name1401 (
		_w3427_,
		_w3625_,
		_w3629_,
		_w3630_
	);
	LUT3 #(
		.INIT('h80)
	) name1402 (
		\ctl_rf_c6_rf_chdad_reg[24]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3631_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1403 (
		\ctl_rf_c6_rf_chsad_reg[24]/NET0131 ,
		\ctl_rf_c6_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3632_
	);
	LUT3 #(
		.INIT('h8a)
	) name1404 (
		_w3440_,
		_w3631_,
		_w3632_,
		_w3633_
	);
	LUT3 #(
		.INIT('h80)
	) name1405 (
		\ctl_rf_c7_rf_chdad_reg[24]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3634_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1406 (
		\ctl_rf_c7_rf_chsad_reg[24]/NET0131 ,
		\ctl_rf_c7_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3635_
	);
	LUT3 #(
		.INIT('h8a)
	) name1407 (
		_w3453_,
		_w3634_,
		_w3635_,
		_w3636_
	);
	LUT3 #(
		.INIT('h02)
	) name1408 (
		\ctl_rf_c0_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3637_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1409 (
		\ctl_rf_c0_rf_chdad_reg[24]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3638_
	);
	LUT3 #(
		.INIT('h8a)
	) name1410 (
		_w3445_,
		_w3637_,
		_w3638_,
		_w3639_
	);
	LUT3 #(
		.INIT('h80)
	) name1411 (
		\ctl_rf_c5_rf_chdad_reg[24]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3640_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1412 (
		\ctl_rf_c5_rf_chsad_reg[24]/NET0131 ,
		\ctl_rf_c5_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3641_
	);
	LUT3 #(
		.INIT('h8a)
	) name1413 (
		_w3436_,
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT4 #(
		.INIT('h0001)
	) name1414 (
		_w3633_,
		_w3636_,
		_w3639_,
		_w3642_,
		_w3643_
	);
	LUT3 #(
		.INIT('h80)
	) name1415 (
		\ctl_rf_c3_rf_chdad_reg[24]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3644_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1416 (
		\ctl_rf_c3_rf_chsad_reg[24]/NET0131 ,
		\ctl_rf_c3_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3645_
	);
	LUT3 #(
		.INIT('h8a)
	) name1417 (
		_w3457_,
		_w3644_,
		_w3645_,
		_w3646_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1418 (
		\ctl_rf_c1_rf_chdad_reg[24]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3647_
	);
	LUT3 #(
		.INIT('ha2)
	) name1419 (
		\haddr[8]_pad ,
		_w3449_,
		_w3647_,
		_w3648_
	);
	LUT3 #(
		.INIT('h02)
	) name1420 (
		\ctl_rf_c4_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3649_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1421 (
		\ctl_rf_c4_rf_chdad_reg[24]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3650_
	);
	LUT3 #(
		.INIT('h8a)
	) name1422 (
		_w3426_,
		_w3649_,
		_w3650_,
		_w3651_
	);
	LUT3 #(
		.INIT('h02)
	) name1423 (
		\ctl_rf_c2_rf_dreqmode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3652_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1424 (
		\ctl_rf_c2_rf_chdad_reg[24]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3653_
	);
	LUT3 #(
		.INIT('h8a)
	) name1425 (
		_w3432_,
		_w3652_,
		_w3653_,
		_w3654_
	);
	LUT4 #(
		.INIT('h0004)
	) name1426 (
		_w3646_,
		_w3648_,
		_w3651_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h8)
	) name1427 (
		_w3643_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h0800)
	) name1428 (
		\ctl_rf_c5brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3657_
	);
	LUT4 #(
		.INIT('h2000)
	) name1429 (
		\ctl_rf_c6brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3658_
	);
	LUT4 #(
		.INIT('h0020)
	) name1430 (
		\ctl_rf_c2brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3659_
	);
	LUT4 #(
		.INIT('h0200)
	) name1431 (
		\ctl_rf_c4brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3660_
	);
	LUT4 #(
		.INIT('h0001)
	) name1432 (
		_w3657_,
		_w3658_,
		_w3659_,
		_w3660_,
		_w3661_
	);
	LUT4 #(
		.INIT('h0080)
	) name1433 (
		\ctl_rf_c3brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3662_
	);
	LUT4 #(
		.INIT('h0008)
	) name1434 (
		\ctl_rf_c1brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3663_
	);
	LUT4 #(
		.INIT('h0002)
	) name1435 (
		\ctl_rf_c0brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3664_
	);
	LUT4 #(
		.INIT('h8000)
	) name1436 (
		\ctl_rf_c7brbs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3665_
	);
	LUT4 #(
		.INIT('h0001)
	) name1437 (
		_w3662_,
		_w3663_,
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT3 #(
		.INIT('h2a)
	) name1438 (
		_w3425_,
		_w3661_,
		_w3666_,
		_w3667_
	);
	LUT4 #(
		.INIT('h0020)
	) name1439 (
		\ctl_rf_c2dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3668_
	);
	LUT4 #(
		.INIT('h2000)
	) name1440 (
		\ctl_rf_c6dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3669_
	);
	LUT4 #(
		.INIT('h0008)
	) name1441 (
		\ctl_rf_c1dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3670_
	);
	LUT4 #(
		.INIT('h0080)
	) name1442 (
		\ctl_rf_c3dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3671_
	);
	LUT4 #(
		.INIT('h0001)
	) name1443 (
		_w3668_,
		_w3669_,
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT4 #(
		.INIT('h0200)
	) name1444 (
		\ctl_rf_c4dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3673_
	);
	LUT4 #(
		.INIT('h0002)
	) name1445 (
		\ctl_rf_c0dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3674_
	);
	LUT4 #(
		.INIT('h0800)
	) name1446 (
		\ctl_rf_c5dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3675_
	);
	LUT4 #(
		.INIT('h8000)
	) name1447 (
		\ctl_rf_c7dmabs_reg[24]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3676_
	);
	LUT4 #(
		.INIT('h0001)
	) name1448 (
		_w3673_,
		_w3674_,
		_w3675_,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('h5111)
	) name1449 (
		\haddr[8]_pad ,
		_w3431_,
		_w3672_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h4)
	) name1450 (
		_w3667_,
		_w3678_,
		_w3679_
	);
	LUT3 #(
		.INIT('h8a)
	) name1451 (
		_w3422_,
		_w3667_,
		_w3678_,
		_w3680_
	);
	LUT4 #(
		.INIT('h1055)
	) name1452 (
		_w3622_,
		_w3630_,
		_w3656_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		\haddr[8]_pad ,
		_w3503_,
		_w3682_
	);
	LUT4 #(
		.INIT('h0001)
	) name1454 (
		_w3503_,
		_w3546_,
		_w3550_,
		_w3554_,
		_w3683_
	);
	LUT4 #(
		.INIT('h070f)
	) name1455 (
		_w3524_,
		_w3542_,
		_w3682_,
		_w3683_,
		_w3684_
	);
	LUT4 #(
		.INIT('haa80)
	) name1456 (
		_w3503_,
		_w3573_,
		_w3589_,
		_w3617_,
		_w3685_
	);
	LUT4 #(
		.INIT('hddcd)
	) name1457 (
		_w3424_,
		_w3681_,
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('hb)
	) name1458 (
		_w3621_,
		_w3686_,
		_w3687_
	);
	LUT3 #(
		.INIT('h2a)
	) name1459 (
		\hrdata_reg[24]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3688_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		\haddr[8]_pad ,
		_w3424_,
		_w3689_
	);
	LUT4 #(
		.INIT('h0002)
	) name1461 (
		_w3424_,
		_w3546_,
		_w3550_,
		_w3554_,
		_w3690_
	);
	LUT4 #(
		.INIT('h070f)
	) name1462 (
		_w3524_,
		_w3542_,
		_w3689_,
		_w3690_,
		_w3691_
	);
	LUT4 #(
		.INIT('h5510)
	) name1463 (
		_w3503_,
		_w3630_,
		_w3656_,
		_w3679_,
		_w3692_
	);
	LUT4 #(
		.INIT('h7500)
	) name1464 (
		_w3484_,
		_w3487_,
		_w3498_,
		_w3503_,
		_w3693_
	);
	LUT2 #(
		.INIT('h4)
	) name1465 (
		_w3483_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('h888a)
	) name1466 (
		_w3422_,
		_w3424_,
		_w3692_,
		_w3694_,
		_w3695_
	);
	LUT3 #(
		.INIT('hea)
	) name1467 (
		_w3688_,
		_w3691_,
		_w3695_,
		_w3696_
	);
	LUT3 #(
		.INIT('h20)
	) name1468 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3697_
	);
	LUT3 #(
		.INIT('h80)
	) name1469 (
		_w2507_,
		_w2508_,
		_w3697_,
		_w3698_
	);
	LUT3 #(
		.INIT('h80)
	) name1470 (
		_w2424_,
		_w2549_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		\de_de_st_reg[0]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3700_
	);
	LUT3 #(
		.INIT('h80)
	) name1472 (
		_w2507_,
		_w2508_,
		_w3700_,
		_w3701_
	);
	LUT3 #(
		.INIT('h2a)
	) name1473 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		_w2549_,
		_w3701_,
		_w3702_
	);
	LUT3 #(
		.INIT('h2a)
	) name1474 (
		\ctl_rf_c0_rf_chllpen_reg/NET0131 ,
		_w2549_,
		_w3698_,
		_w3703_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w3702_,
		_w3703_,
		_w3704_
	);
	LUT4 #(
		.INIT('hff70)
	) name1476 (
		_w3059_,
		_w3104_,
		_w3699_,
		_w3704_,
		_w3705_
	);
	LUT3 #(
		.INIT('h20)
	) name1477 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3706_
	);
	LUT3 #(
		.INIT('h70)
	) name1478 (
		_w2507_,
		_w2508_,
		_w3706_,
		_w3707_
	);
	LUT3 #(
		.INIT('h80)
	) name1479 (
		_w2424_,
		_w2549_,
		_w3707_,
		_w3708_
	);
	LUT3 #(
		.INIT('h70)
	) name1480 (
		_w2507_,
		_w2508_,
		_w3700_,
		_w3709_
	);
	LUT3 #(
		.INIT('h2a)
	) name1481 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		_w2549_,
		_w3709_,
		_w3710_
	);
	LUT3 #(
		.INIT('h2a)
	) name1482 (
		\ctl_rf_c1_rf_chllpen_reg/NET0131 ,
		_w2549_,
		_w3707_,
		_w3711_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT4 #(
		.INIT('hff70)
	) name1484 (
		_w3059_,
		_w3104_,
		_w3708_,
		_w3712_,
		_w3713_
	);
	LUT3 #(
		.INIT('h20)
	) name1485 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3714_
	);
	LUT3 #(
		.INIT('h80)
	) name1486 (
		_w2507_,
		_w2508_,
		_w3714_,
		_w3715_
	);
	LUT3 #(
		.INIT('h80)
	) name1487 (
		_w2424_,
		_w2534_,
		_w3715_,
		_w3716_
	);
	LUT3 #(
		.INIT('h2a)
	) name1488 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		_w2534_,
		_w3701_,
		_w3717_
	);
	LUT3 #(
		.INIT('h2a)
	) name1489 (
		\ctl_rf_c2_rf_chllpen_reg/NET0131 ,
		_w2534_,
		_w3715_,
		_w3718_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		_w3717_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('hff70)
	) name1491 (
		_w3059_,
		_w3104_,
		_w3716_,
		_w3719_,
		_w3720_
	);
	LUT3 #(
		.INIT('h20)
	) name1492 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3721_
	);
	LUT3 #(
		.INIT('h70)
	) name1493 (
		_w2507_,
		_w2508_,
		_w3721_,
		_w3722_
	);
	LUT3 #(
		.INIT('h80)
	) name1494 (
		_w2424_,
		_w2534_,
		_w3722_,
		_w3723_
	);
	LUT3 #(
		.INIT('h2a)
	) name1495 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2534_,
		_w3709_,
		_w3724_
	);
	LUT3 #(
		.INIT('h2a)
	) name1496 (
		\ctl_rf_c3_rf_chllpen_reg/NET0131 ,
		_w2534_,
		_w3722_,
		_w3725_
	);
	LUT2 #(
		.INIT('h4)
	) name1497 (
		_w3724_,
		_w3725_,
		_w3726_
	);
	LUT4 #(
		.INIT('hff70)
	) name1498 (
		_w3059_,
		_w3104_,
		_w3723_,
		_w3726_,
		_w3727_
	);
	LUT3 #(
		.INIT('h20)
	) name1499 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3728_
	);
	LUT3 #(
		.INIT('h80)
	) name1500 (
		_w2507_,
		_w2508_,
		_w3728_,
		_w3729_
	);
	LUT3 #(
		.INIT('h80)
	) name1501 (
		_w2424_,
		_w2520_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('h2a)
	) name1502 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		_w2520_,
		_w3701_,
		_w3731_
	);
	LUT3 #(
		.INIT('h2a)
	) name1503 (
		\ctl_rf_c4_rf_chllpen_reg/NET0131 ,
		_w2520_,
		_w3729_,
		_w3732_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w3731_,
		_w3732_,
		_w3733_
	);
	LUT4 #(
		.INIT('hff70)
	) name1505 (
		_w3059_,
		_w3104_,
		_w3730_,
		_w3733_,
		_w3734_
	);
	LUT3 #(
		.INIT('h20)
	) name1506 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3735_
	);
	LUT3 #(
		.INIT('h70)
	) name1507 (
		_w2507_,
		_w2508_,
		_w3735_,
		_w3736_
	);
	LUT3 #(
		.INIT('h80)
	) name1508 (
		_w2424_,
		_w2520_,
		_w3736_,
		_w3737_
	);
	LUT3 #(
		.INIT('h2a)
	) name1509 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		_w2520_,
		_w3709_,
		_w3738_
	);
	LUT3 #(
		.INIT('h2a)
	) name1510 (
		\ctl_rf_c5_rf_chllpen_reg/NET0131 ,
		_w2520_,
		_w3736_,
		_w3739_
	);
	LUT2 #(
		.INIT('h4)
	) name1511 (
		_w3738_,
		_w3739_,
		_w3740_
	);
	LUT4 #(
		.INIT('hff70)
	) name1512 (
		_w3059_,
		_w3104_,
		_w3737_,
		_w3740_,
		_w3741_
	);
	LUT3 #(
		.INIT('h20)
	) name1513 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3742_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		_w2507_,
		_w2508_,
		_w3742_,
		_w3743_
	);
	LUT3 #(
		.INIT('h80)
	) name1515 (
		_w2424_,
		_w2527_,
		_w3743_,
		_w3744_
	);
	LUT3 #(
		.INIT('h2a)
	) name1516 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		_w2527_,
		_w3701_,
		_w3745_
	);
	LUT3 #(
		.INIT('h2a)
	) name1517 (
		\ctl_rf_c6_rf_chllpen_reg/NET0131 ,
		_w2527_,
		_w3743_,
		_w3746_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT4 #(
		.INIT('hff70)
	) name1519 (
		_w3059_,
		_w3104_,
		_w3744_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('h20)
	) name1520 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3749_
	);
	LUT3 #(
		.INIT('h70)
	) name1521 (
		_w2507_,
		_w2508_,
		_w3749_,
		_w3750_
	);
	LUT3 #(
		.INIT('h80)
	) name1522 (
		_w2424_,
		_w2527_,
		_w3750_,
		_w3751_
	);
	LUT3 #(
		.INIT('h2a)
	) name1523 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2527_,
		_w3709_,
		_w3752_
	);
	LUT3 #(
		.INIT('h2a)
	) name1524 (
		\ctl_rf_c7_rf_chllpen_reg/NET0131 ,
		_w2527_,
		_w3750_,
		_w3753_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT4 #(
		.INIT('hff70)
	) name1526 (
		_w3059_,
		_w3104_,
		_w3751_,
		_w3754_,
		_w3755_
	);
	LUT3 #(
		.INIT('h10)
	) name1527 (
		\de_de_st_reg[2]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		_w3756_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		_w3406_,
		_w3756_,
		_w3757_
	);
	LUT3 #(
		.INIT('hf4)
	) name1529 (
		_w3267_,
		_w3392_,
		_w3757_,
		_w3758_
	);
	LUT3 #(
		.INIT('h15)
	) name1530 (
		\de_de_st_reg[0]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w3759_
	);
	LUT4 #(
		.INIT('h000e)
	) name1531 (
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		_w3760_
	);
	LUT4 #(
		.INIT('h0777)
	) name1532 (
		_w3406_,
		_w3756_,
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT4 #(
		.INIT('hdfd0)
	) name1533 (
		\ch_sel_arb_req_reg/NET0131 ,
		_w2577_,
		_w3356_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h2)
	) name1534 (
		\ch_sel_arb_req_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w3763_
	);
	LUT4 #(
		.INIT('hd500)
	) name1535 (
		\de_de_st_reg[0]/NET0131 ,
		_w2575_,
		_w2576_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		\ch_sel_arb_req_reg/NET0131 ,
		\ch_sel_de_stup_d1_reg/NET0131 ,
		_w3765_
	);
	LUT4 #(
		.INIT('hd500)
	) name1537 (
		\de_de_st_reg[0]/NET0131 ,
		_w2575_,
		_w2576_,
		_w3765_,
		_w3766_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1538 (
		_w2546_,
		_w2572_,
		_w3764_,
		_w3766_,
		_w3767_
	);
	LUT3 #(
		.INIT('h2a)
	) name1539 (
		\hrdata_reg[0]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3768_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1540 (
		_w3422_,
		_w3600_,
		_w3611_,
		_w3616_,
		_w3769_
	);
	LUT4 #(
		.INIT('h080f)
	) name1541 (
		_w3573_,
		_w3589_,
		_w3622_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		_w3768_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('haa20)
	) name1543 (
		_w3503_,
		_w3630_,
		_w3656_,
		_w3679_,
		_w3772_
	);
	LUT4 #(
		.INIT('h0075)
	) name1544 (
		_w3484_,
		_w3487_,
		_w3498_,
		_w3503_,
		_w3773_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w3483_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		_w3424_,
		_w3768_,
		_w3775_
	);
	LUT3 #(
		.INIT('he0)
	) name1547 (
		_w3772_,
		_w3774_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w3771_,
		_w3776_,
		_w3777_
	);
	LUT3 #(
		.INIT('h2a)
	) name1549 (
		\hrdata_reg[1]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3778_
	);
	LUT4 #(
		.INIT('hff53)
	) name1550 (
		\ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131 ,
		\ctl_rf_c0_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3779_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1551 (
		\ctl_rf_c0_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c0_rf_chsad_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3780_
	);
	LUT4 #(
		.INIT('ha222)
	) name1552 (
		\haddr[8]_pad ,
		_w3445_,
		_w3779_,
		_w3780_,
		_w3781_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1553 (
		\ctl_rf_c2_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3782_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1554 (
		\ctl_rf_c2_rf_chsad_reg[17]/NET0131 ,
		\ctl_rf_c2_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3783_
	);
	LUT3 #(
		.INIT('h2a)
	) name1555 (
		_w3432_,
		_w3782_,
		_w3783_,
		_w3784_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1556 (
		\ctl_rf_c4_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3785_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1557 (
		\ctl_rf_c4_rf_chsad_reg[17]/NET0131 ,
		\ctl_rf_c4_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3786_
	);
	LUT3 #(
		.INIT('h2a)
	) name1558 (
		_w3426_,
		_w3785_,
		_w3786_,
		_w3787_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1559 (
		\ctl_rf_c7_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3788_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1560 (
		\ctl_rf_c7_rf_chsad_reg[17]/NET0131 ,
		\ctl_rf_c7_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3789_
	);
	LUT3 #(
		.INIT('h2a)
	) name1561 (
		_w3453_,
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('hff53)
	) name1562 (
		\ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131 ,
		\ctl_rf_c1_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3791_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1563 (
		\ctl_rf_c1_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3792_
	);
	LUT3 #(
		.INIT('h2a)
	) name1564 (
		_w3449_,
		_w3791_,
		_w3792_,
		_w3793_
	);
	LUT4 #(
		.INIT('h0001)
	) name1565 (
		_w3784_,
		_w3787_,
		_w3790_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name1566 (
		_w3781_,
		_w3794_,
		_w3795_
	);
	LUT4 #(
		.INIT('h153f)
	) name1567 (
		\ctl_rf_c3_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[17]/NET0131 ,
		_w3469_,
		_w3477_,
		_w3796_
	);
	LUT4 #(
		.INIT('h135f)
	) name1568 (
		\ctl_rf_c0_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[17]/NET0131 ,
		_w3467_,
		_w3472_,
		_w3797_
	);
	LUT4 #(
		.INIT('h135f)
	) name1569 (
		\ctl_rf_c2_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[17]/NET0131 ,
		_w3462_,
		_w3479_,
		_w3798_
	);
	LUT4 #(
		.INIT('h153f)
	) name1570 (
		\ctl_rf_c1_rf_chllp_reg[17]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[17]/NET0131 ,
		_w3464_,
		_w3474_,
		_w3799_
	);
	LUT4 #(
		.INIT('h8000)
	) name1571 (
		_w3796_,
		_w3797_,
		_w3798_,
		_w3799_,
		_w3800_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1572 (
		\ctl_rf_c6_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c6_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3801_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1573 (
		\ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131 ,
		\ctl_rf_c6_rf_chsad_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3802_
	);
	LUT3 #(
		.INIT('h2a)
	) name1574 (
		_w3440_,
		_w3801_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1575 (
		\ctl_rf_c5_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3804_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1576 (
		\ctl_rf_c5_rf_chsad_reg[17]/NET0131 ,
		\ctl_rf_c5_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3805_
	);
	LUT3 #(
		.INIT('h2a)
	) name1577 (
		_w3436_,
		_w3804_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1578 (
		\ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131 ,
		\ctl_rf_c3_rf_chsad_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3807_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1579 (
		\ctl_rf_c3_rf_chdad_reg[17]/NET0131 ,
		\ctl_rf_c3_rf_src_sz_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3808_
	);
	LUT3 #(
		.INIT('h2a)
	) name1580 (
		_w3457_,
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT3 #(
		.INIT('h01)
	) name1581 (
		_w3803_,
		_w3806_,
		_w3809_,
		_w3810_
	);
	LUT3 #(
		.INIT('hd0)
	) name1582 (
		_w3427_,
		_w3800_,
		_w3810_,
		_w3811_
	);
	LUT4 #(
		.INIT('h0008)
	) name1583 (
		\ctl_rf_c1brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3812_
	);
	LUT4 #(
		.INIT('h0080)
	) name1584 (
		\ctl_rf_c3brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3813_
	);
	LUT4 #(
		.INIT('h0002)
	) name1585 (
		\ctl_rf_c0brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3814_
	);
	LUT4 #(
		.INIT('h8000)
	) name1586 (
		\ctl_rf_c7brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3815_
	);
	LUT4 #(
		.INIT('h0001)
	) name1587 (
		_w3812_,
		_w3813_,
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT4 #(
		.INIT('h2000)
	) name1588 (
		\ctl_rf_c6brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3817_
	);
	LUT4 #(
		.INIT('h0200)
	) name1589 (
		\ctl_rf_c4brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3818_
	);
	LUT4 #(
		.INIT('h0020)
	) name1590 (
		\ctl_rf_c2brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3819_
	);
	LUT4 #(
		.INIT('h0800)
	) name1591 (
		\ctl_rf_c5brbs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3820_
	);
	LUT4 #(
		.INIT('h0001)
	) name1592 (
		_w3817_,
		_w3818_,
		_w3819_,
		_w3820_,
		_w3821_
	);
	LUT3 #(
		.INIT('h2a)
	) name1593 (
		_w3425_,
		_w3816_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h0020)
	) name1594 (
		\ctl_rf_c2dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3823_
	);
	LUT4 #(
		.INIT('h0080)
	) name1595 (
		\ctl_rf_c3dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3824_
	);
	LUT4 #(
		.INIT('h0002)
	) name1596 (
		\ctl_rf_c0dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3825_
	);
	LUT4 #(
		.INIT('h2000)
	) name1597 (
		\ctl_rf_c6dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3826_
	);
	LUT4 #(
		.INIT('h0001)
	) name1598 (
		_w3823_,
		_w3824_,
		_w3825_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('h8000)
	) name1599 (
		\ctl_rf_c7dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3828_
	);
	LUT4 #(
		.INIT('h0200)
	) name1600 (
		\ctl_rf_c4dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3829_
	);
	LUT4 #(
		.INIT('h0008)
	) name1601 (
		\ctl_rf_c1dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3830_
	);
	LUT4 #(
		.INIT('h0800)
	) name1602 (
		\ctl_rf_c5dmabs_reg[17]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3831_
	);
	LUT4 #(
		.INIT('h0001)
	) name1603 (
		_w3828_,
		_w3829_,
		_w3830_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('h2a)
	) name1604 (
		_w3431_,
		_w3827_,
		_w3832_,
		_w3833_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1605 (
		\ctl_rf_abt_reg[1]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w3834_
	);
	LUT4 #(
		.INIT('h0023)
	) name1606 (
		\ctl_rf_c1_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT3 #(
		.INIT('h01)
	) name1608 (
		_w3822_,
		_w3833_,
		_w3836_,
		_w3837_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1609 (
		_w3422_,
		_w3822_,
		_w3833_,
		_w3836_,
		_w3838_
	);
	LUT4 #(
		.INIT('h4055)
	) name1610 (
		_w3622_,
		_w3795_,
		_w3811_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w3778_,
		_w3839_,
		_w3840_
	);
	LUT4 #(
		.INIT('h0800)
	) name1612 (
		\ctl_rf_c5dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3841_
	);
	LUT4 #(
		.INIT('h2000)
	) name1613 (
		\ctl_rf_c6dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3842_
	);
	LUT4 #(
		.INIT('h0020)
	) name1614 (
		\ctl_rf_c2dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3843_
	);
	LUT4 #(
		.INIT('h0200)
	) name1615 (
		\ctl_rf_c4dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3844_
	);
	LUT4 #(
		.INIT('h0001)
	) name1616 (
		_w3841_,
		_w3842_,
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT4 #(
		.INIT('h0080)
	) name1617 (
		\ctl_rf_c3dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3846_
	);
	LUT4 #(
		.INIT('h0008)
	) name1618 (
		\ctl_rf_c1dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3847_
	);
	LUT4 #(
		.INIT('h0002)
	) name1619 (
		\ctl_rf_c0dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3848_
	);
	LUT4 #(
		.INIT('h8000)
	) name1620 (
		\ctl_rf_c7dmabs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3849_
	);
	LUT4 #(
		.INIT('h0001)
	) name1621 (
		_w3846_,
		_w3847_,
		_w3848_,
		_w3849_,
		_w3850_
	);
	LUT3 #(
		.INIT('h2a)
	) name1622 (
		_w3431_,
		_w3845_,
		_w3850_,
		_w3851_
	);
	LUT4 #(
		.INIT('h0020)
	) name1623 (
		\ctl_rf_c2brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3852_
	);
	LUT4 #(
		.INIT('h2000)
	) name1624 (
		\ctl_rf_c6brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3853_
	);
	LUT4 #(
		.INIT('h0008)
	) name1625 (
		\ctl_rf_c1brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3854_
	);
	LUT4 #(
		.INIT('h0080)
	) name1626 (
		\ctl_rf_c3brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3855_
	);
	LUT4 #(
		.INIT('h0001)
	) name1627 (
		_w3852_,
		_w3853_,
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT4 #(
		.INIT('h0200)
	) name1628 (
		\ctl_rf_c4brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3857_
	);
	LUT4 #(
		.INIT('h0002)
	) name1629 (
		\ctl_rf_c0brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3858_
	);
	LUT4 #(
		.INIT('h0800)
	) name1630 (
		\ctl_rf_c5brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3859_
	);
	LUT4 #(
		.INIT('h8000)
	) name1631 (
		\ctl_rf_c7brbs_reg[25]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w3860_
	);
	LUT4 #(
		.INIT('h0001)
	) name1632 (
		_w3857_,
		_w3858_,
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT4 #(
		.INIT('h5111)
	) name1633 (
		\haddr[8]_pad ,
		_w3425_,
		_w3856_,
		_w3861_,
		_w3862_
	);
	LUT3 #(
		.INIT('h20)
	) name1634 (
		_w3503_,
		_w3851_,
		_w3862_,
		_w3863_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1635 (
		\ctl_rf_c4_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w3426_,
		_w3864_,
		_w3865_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1637 (
		\ctl_rf_c1_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3866_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1638 (
		\ctl_rf_c3_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3867_
	);
	LUT4 #(
		.INIT('hf531)
	) name1639 (
		_w3449_,
		_w3457_,
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h4)
	) name1640 (
		_w3865_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1641 (
		\ctl_rf_c7_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3870_
	);
	LUT3 #(
		.INIT('ha2)
	) name1642 (
		\haddr[8]_pad ,
		_w3453_,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1643 (
		\ctl_rf_c6_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3872_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1644 (
		\ctl_rf_c2_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3873_
	);
	LUT4 #(
		.INIT('hf351)
	) name1645 (
		_w3432_,
		_w3440_,
		_w3872_,
		_w3873_,
		_w3874_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1646 (
		\ctl_rf_c5_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3875_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1647 (
		\ctl_rf_c0_rf_chdad_reg[25]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[25]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3876_
	);
	LUT4 #(
		.INIT('hf531)
	) name1648 (
		_w3436_,
		_w3445_,
		_w3875_,
		_w3876_,
		_w3877_
	);
	LUT3 #(
		.INIT('h80)
	) name1649 (
		_w3871_,
		_w3874_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		_w3869_,
		_w3878_,
		_w3879_
	);
	LUT4 #(
		.INIT('h135f)
	) name1651 (
		\ctl_rf_c1_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[25]/NET0131 ,
		_w3474_,
		_w3477_,
		_w3880_
	);
	LUT4 #(
		.INIT('h135f)
	) name1652 (
		\ctl_rf_c0_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[25]/NET0131 ,
		_w3467_,
		_w3472_,
		_w3881_
	);
	LUT4 #(
		.INIT('h135f)
	) name1653 (
		\ctl_rf_c5_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[25]/NET0131 ,
		_w3469_,
		_w3479_,
		_w3882_
	);
	LUT4 #(
		.INIT('h135f)
	) name1654 (
		\ctl_rf_c2_rf_chllp_reg[25]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[25]/NET0131 ,
		_w3462_,
		_w3464_,
		_w3883_
	);
	LUT4 #(
		.INIT('h8000)
	) name1655 (
		_w3880_,
		_w3881_,
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT3 #(
		.INIT('hc4)
	) name1656 (
		_w3427_,
		_w3503_,
		_w3884_,
		_w3885_
	);
	LUT3 #(
		.INIT('h15)
	) name1657 (
		_w3863_,
		_w3879_,
		_w3885_,
		_w3886_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1658 (
		\ctl_rf_c7_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3887_
	);
	LUT4 #(
		.INIT('hff35)
	) name1659 (
		\ctl_rf_c7_rf_dst_sel_reg/NET0131 ,
		\ctl_rf_c7_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3888_
	);
	LUT3 #(
		.INIT('h2a)
	) name1660 (
		_w3453_,
		_w3887_,
		_w3888_,
		_w3889_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1661 (
		\ctl_rf_c3_rf_chsad_reg[1]/NET0131 ,
		\ctl_rf_c3_rf_dst_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3890_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1662 (
		\ctl_rf_c3_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c3_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3891_
	);
	LUT3 #(
		.INIT('h2a)
	) name1663 (
		_w3457_,
		_w3890_,
		_w3891_,
		_w3892_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1664 (
		\ctl_rf_c0_rf_chsad_reg[1]/NET0131 ,
		\ctl_rf_c0_rf_dst_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3893_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1665 (
		\ctl_rf_c0_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c0_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3894_
	);
	LUT3 #(
		.INIT('h2a)
	) name1666 (
		_w3445_,
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1667 (
		\ctl_rf_c1_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3896_
	);
	LUT4 #(
		.INIT('hff35)
	) name1668 (
		\ctl_rf_c1_rf_dst_sel_reg/NET0131 ,
		\ctl_rf_c1_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3897_
	);
	LUT3 #(
		.INIT('h2a)
	) name1669 (
		_w3449_,
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT4 #(
		.INIT('h0001)
	) name1670 (
		_w3889_,
		_w3892_,
		_w3895_,
		_w3898_,
		_w3899_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1671 (
		\ctl_rf_c5_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3900_
	);
	LUT4 #(
		.INIT('hff35)
	) name1672 (
		\ctl_rf_c5_rf_dst_sel_reg/NET0131 ,
		\ctl_rf_c5_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3901_
	);
	LUT3 #(
		.INIT('h2a)
	) name1673 (
		_w3436_,
		_w3900_,
		_w3901_,
		_w3902_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1674 (
		\ctl_rf_c6_rf_chsad_reg[1]/NET0131 ,
		\ctl_rf_c6_rf_dst_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3903_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1675 (
		\ctl_rf_c6_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c6_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3904_
	);
	LUT3 #(
		.INIT('h2a)
	) name1676 (
		_w3440_,
		_w3903_,
		_w3904_,
		_w3905_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1677 (
		\ctl_rf_c4_rf_chsad_reg[1]/NET0131 ,
		\ctl_rf_c4_rf_dst_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3906_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1678 (
		\ctl_rf_c4_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c4_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3907_
	);
	LUT3 #(
		.INIT('h2a)
	) name1679 (
		_w3426_,
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1680 (
		\ctl_rf_c2_rf_chdad_reg[1]/NET0131 ,
		\ctl_rf_c2_rf_chsad_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3909_
	);
	LUT4 #(
		.INIT('hff35)
	) name1681 (
		\ctl_rf_c2_rf_dst_sel_reg/NET0131 ,
		\ctl_rf_c2_rf_int_err_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3910_
	);
	LUT3 #(
		.INIT('h2a)
	) name1682 (
		_w3432_,
		_w3909_,
		_w3910_,
		_w3911_
	);
	LUT4 #(
		.INIT('h0001)
	) name1683 (
		_w3902_,
		_w3905_,
		_w3908_,
		_w3911_,
		_w3912_
	);
	LUT4 #(
		.INIT('hff35)
	) name1684 (
		\ctl_rf_c0_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c0_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3913_
	);
	LUT4 #(
		.INIT('hff35)
	) name1685 (
		\ctl_rf_c3_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c3_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3914_
	);
	LUT4 #(
		.INIT('hf531)
	) name1686 (
		_w3467_,
		_w3477_,
		_w3913_,
		_w3914_,
		_w3915_
	);
	LUT4 #(
		.INIT('hff35)
	) name1687 (
		\ctl_rf_c1_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c1_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3916_
	);
	LUT4 #(
		.INIT('hff35)
	) name1688 (
		\ctl_rf_c2_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c2_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3917_
	);
	LUT4 #(
		.INIT('hf351)
	) name1689 (
		_w3462_,
		_w3474_,
		_w3916_,
		_w3917_,
		_w3918_
	);
	LUT4 #(
		.INIT('hff35)
	) name1690 (
		\ctl_rf_c7_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c7_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3919_
	);
	LUT4 #(
		.INIT('hff35)
	) name1691 (
		\ctl_rf_c5_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c5_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3920_
	);
	LUT4 #(
		.INIT('hf531)
	) name1692 (
		_w3464_,
		_w3469_,
		_w3919_,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('hff35)
	) name1693 (
		\ctl_rf_c6_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c6_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3922_
	);
	LUT4 #(
		.INIT('hff35)
	) name1694 (
		\ctl_rf_c4_rf_chllp_reg[1]/P0002 ,
		\ctl_rf_c4_rf_chtsz_reg[1]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3923_
	);
	LUT4 #(
		.INIT('hf351)
	) name1695 (
		_w3472_,
		_w3479_,
		_w3922_,
		_w3923_,
		_w3924_
	);
	LUT4 #(
		.INIT('h8000)
	) name1696 (
		_w3915_,
		_w3918_,
		_w3921_,
		_w3924_,
		_w3925_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1697 (
		\haddr[8]_pad ,
		_w3899_,
		_w3912_,
		_w3925_,
		_w3926_
	);
	LUT4 #(
		.INIT('h1500)
	) name1698 (
		\de_de_st_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w3485_,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		_w2549_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h2)
	) name1700 (
		\ctl_rf_c1_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[4]_pad ,
		_w3929_
	);
	LUT3 #(
		.INIT('h02)
	) name1701 (
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[5]_pad ,
		_w3930_
	);
	LUT3 #(
		.INIT('h20)
	) name1702 (
		\ctl_rf_tc_reg[1]/NET0131 ,
		_w3929_,
		_w3930_,
		_w3931_
	);
	LUT4 #(
		.INIT('h135f)
	) name1703 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_m0end_reg/NET0131 ,
		_w3492_,
		_w3494_,
		_w3932_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1704 (
		\ctl_rf_abt_reg[1]/NET0131 ,
		\ctl_rf_c1_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c1_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[1]/NET0131 ,
		_w3933_
	);
	LUT4 #(
		.INIT('h7707)
	) name1705 (
		\ctl_rf_sync_reg[1]/NET0131 ,
		_w3491_,
		_w3496_,
		_w3933_,
		_w3934_
	);
	LUT3 #(
		.INIT('h40)
	) name1706 (
		_w3931_,
		_w3932_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('h1311)
	) name1707 (
		_w3484_,
		_w3503_,
		_w3928_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		_w3926_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w3424_,
		_w3778_,
		_w3938_
	);
	LUT3 #(
		.INIT('hd0)
	) name1710 (
		_w3886_,
		_w3937_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w3840_,
		_w3939_,
		_w3940_
	);
	LUT3 #(
		.INIT('h2a)
	) name1712 (
		\hrdata_reg[25]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3941_
	);
	LUT3 #(
		.INIT('h20)
	) name1713 (
		\ctl_rf_c2_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3942_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1714 (
		\ctl_rf_c2_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c2_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3943_
	);
	LUT3 #(
		.INIT('h8a)
	) name1715 (
		_w3432_,
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT3 #(
		.INIT('h20)
	) name1716 (
		\ctl_rf_c0_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3945_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1717 (
		\ctl_rf_c0_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c0_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3946_
	);
	LUT3 #(
		.INIT('h8a)
	) name1718 (
		_w3445_,
		_w3945_,
		_w3946_,
		_w3947_
	);
	LUT3 #(
		.INIT('h20)
	) name1719 (
		\ctl_rf_c3_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3948_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1720 (
		\ctl_rf_c3_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c3_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3949_
	);
	LUT3 #(
		.INIT('h8a)
	) name1721 (
		_w3457_,
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT3 #(
		.INIT('h20)
	) name1722 (
		\ctl_rf_c5_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3951_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1723 (
		\ctl_rf_c5_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c5_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3952_
	);
	LUT3 #(
		.INIT('h8a)
	) name1724 (
		_w3436_,
		_w3951_,
		_w3952_,
		_w3953_
	);
	LUT4 #(
		.INIT('h0001)
	) name1725 (
		_w3944_,
		_w3947_,
		_w3950_,
		_w3953_,
		_w3954_
	);
	LUT4 #(
		.INIT('hff35)
	) name1726 (
		\ctl_rf_c3_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3955_
	);
	LUT4 #(
		.INIT('hff35)
	) name1727 (
		\ctl_rf_c2_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3956_
	);
	LUT4 #(
		.INIT('hf351)
	) name1728 (
		_w3462_,
		_w3477_,
		_w3955_,
		_w3956_,
		_w3957_
	);
	LUT4 #(
		.INIT('hff35)
	) name1729 (
		\ctl_rf_c1_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3958_
	);
	LUT4 #(
		.INIT('hff35)
	) name1730 (
		\ctl_rf_c0_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3959_
	);
	LUT4 #(
		.INIT('hf351)
	) name1731 (
		_w3467_,
		_w3474_,
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT4 #(
		.INIT('hff35)
	) name1732 (
		\ctl_rf_c5_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3961_
	);
	LUT4 #(
		.INIT('hff35)
	) name1733 (
		\ctl_rf_c4_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3962_
	);
	LUT4 #(
		.INIT('hf531)
	) name1734 (
		_w3469_,
		_w3472_,
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('hff35)
	) name1735 (
		\ctl_rf_c6_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3964_
	);
	LUT4 #(
		.INIT('hff35)
	) name1736 (
		\ctl_rf_c7_rf_chllp_reg[9]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[9]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3965_
	);
	LUT4 #(
		.INIT('hf351)
	) name1737 (
		_w3464_,
		_w3479_,
		_w3964_,
		_w3965_,
		_w3966_
	);
	LUT4 #(
		.INIT('h8000)
	) name1738 (
		_w3957_,
		_w3960_,
		_w3963_,
		_w3966_,
		_w3967_
	);
	LUT3 #(
		.INIT('h20)
	) name1739 (
		\ctl_rf_c1_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3968_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1740 (
		\ctl_rf_c1_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c1_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3969_
	);
	LUT3 #(
		.INIT('h8a)
	) name1741 (
		_w3449_,
		_w3968_,
		_w3969_,
		_w3970_
	);
	LUT3 #(
		.INIT('h20)
	) name1742 (
		\ctl_rf_c4_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3971_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1743 (
		\ctl_rf_c4_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c4_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3972_
	);
	LUT3 #(
		.INIT('h8a)
	) name1744 (
		_w3426_,
		_w3971_,
		_w3972_,
		_w3973_
	);
	LUT3 #(
		.INIT('h20)
	) name1745 (
		\ctl_rf_c6_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3974_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1746 (
		\ctl_rf_c6_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c6_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3975_
	);
	LUT3 #(
		.INIT('h8a)
	) name1747 (
		_w3440_,
		_w3974_,
		_w3975_,
		_w3976_
	);
	LUT3 #(
		.INIT('h20)
	) name1748 (
		\ctl_rf_c7_rf_chsad_reg[9]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3977_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1749 (
		\ctl_rf_c7_rf_chdad_reg[9]/P0002 ,
		\ctl_rf_c7_rf_dwidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3978_
	);
	LUT3 #(
		.INIT('h8a)
	) name1750 (
		_w3453_,
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT4 #(
		.INIT('h0001)
	) name1751 (
		_w3970_,
		_w3973_,
		_w3976_,
		_w3979_,
		_w3980_
	);
	LUT4 #(
		.INIT('h8000)
	) name1752 (
		_w3424_,
		_w3954_,
		_w3967_,
		_w3980_,
		_w3981_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1753 (
		\hrdata_reg[25]_pad ,
		_w3422_,
		_w3689_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h10)
	) name1754 (
		_w3503_,
		_w3851_,
		_w3862_,
		_w3983_
	);
	LUT3 #(
		.INIT('h31)
	) name1755 (
		_w3427_,
		_w3503_,
		_w3884_,
		_w3984_
	);
	LUT3 #(
		.INIT('h13)
	) name1756 (
		_w3879_,
		_w3983_,
		_w3984_,
		_w3985_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1757 (
		_w3484_,
		_w3503_,
		_w3928_,
		_w3935_,
		_w3986_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		_w3926_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w3424_,
		_w3941_,
		_w3988_
	);
	LUT4 #(
		.INIT('h0455)
	) name1760 (
		_w3982_,
		_w3985_,
		_w3987_,
		_w3988_,
		_w3989_
	);
	LUT3 #(
		.INIT('h2a)
	) name1761 (
		\hrdata_reg[26]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w3990_
	);
	LUT3 #(
		.INIT('h20)
	) name1762 (
		\ctl_rf_c2_rf_chsad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3991_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1763 (
		\ctl_rf_c2_rf_chdad_reg[10]/P0002 ,
		\ctl_rf_c2_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3992_
	);
	LUT3 #(
		.INIT('h8a)
	) name1764 (
		_w3432_,
		_w3991_,
		_w3992_,
		_w3993_
	);
	LUT3 #(
		.INIT('h20)
	) name1765 (
		\ctl_rf_c0_rf_chsad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3994_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1766 (
		\ctl_rf_c0_rf_chdad_reg[10]/P0002 ,
		\ctl_rf_c0_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3995_
	);
	LUT3 #(
		.INIT('h8a)
	) name1767 (
		_w3445_,
		_w3994_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('h20)
	) name1768 (
		\ctl_rf_c5_rf_chsad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3997_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1769 (
		\ctl_rf_c5_rf_chdad_reg[10]/P0002 ,
		\ctl_rf_c5_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w3998_
	);
	LUT3 #(
		.INIT('h8a)
	) name1770 (
		_w3436_,
		_w3997_,
		_w3998_,
		_w3999_
	);
	LUT3 #(
		.INIT('h80)
	) name1771 (
		\ctl_rf_c3_rf_chdad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4000_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1772 (
		\ctl_rf_c3_rf_chsad_reg[10]/P0002 ,
		\ctl_rf_c3_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4001_
	);
	LUT3 #(
		.INIT('h8a)
	) name1773 (
		_w3457_,
		_w4000_,
		_w4001_,
		_w4002_
	);
	LUT4 #(
		.INIT('h0001)
	) name1774 (
		_w3993_,
		_w3996_,
		_w3999_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('hff35)
	) name1775 (
		\ctl_rf_c3_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4004_
	);
	LUT4 #(
		.INIT('hff35)
	) name1776 (
		\ctl_rf_c5_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4005_
	);
	LUT4 #(
		.INIT('hf351)
	) name1777 (
		_w3469_,
		_w3477_,
		_w4004_,
		_w4005_,
		_w4006_
	);
	LUT4 #(
		.INIT('hff35)
	) name1778 (
		\ctl_rf_c0_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4007_
	);
	LUT4 #(
		.INIT('hff35)
	) name1779 (
		\ctl_rf_c1_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4008_
	);
	LUT4 #(
		.INIT('hf531)
	) name1780 (
		_w3467_,
		_w3474_,
		_w4007_,
		_w4008_,
		_w4009_
	);
	LUT4 #(
		.INIT('hff35)
	) name1781 (
		\ctl_rf_c2_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4010_
	);
	LUT4 #(
		.INIT('hff35)
	) name1782 (
		\ctl_rf_c4_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4011_
	);
	LUT4 #(
		.INIT('hf531)
	) name1783 (
		_w3462_,
		_w3472_,
		_w4010_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('hff35)
	) name1784 (
		\ctl_rf_c6_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4013_
	);
	LUT4 #(
		.INIT('hff35)
	) name1785 (
		\ctl_rf_c7_rf_chllp_reg[10]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[10]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4014_
	);
	LUT4 #(
		.INIT('hf351)
	) name1786 (
		_w3464_,
		_w3479_,
		_w4013_,
		_w4014_,
		_w4015_
	);
	LUT4 #(
		.INIT('h8000)
	) name1787 (
		_w4006_,
		_w4009_,
		_w4012_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h80)
	) name1788 (
		\ctl_rf_c1_rf_chdad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4017_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1789 (
		\ctl_rf_c1_rf_chsad_reg[10]/P0002 ,
		\ctl_rf_c1_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4018_
	);
	LUT3 #(
		.INIT('h8a)
	) name1790 (
		_w3449_,
		_w4017_,
		_w4018_,
		_w4019_
	);
	LUT3 #(
		.INIT('h20)
	) name1791 (
		\ctl_rf_c4_rf_chsad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4020_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1792 (
		\ctl_rf_c4_rf_chdad_reg[10]/P0002 ,
		\ctl_rf_c4_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4021_
	);
	LUT3 #(
		.INIT('h8a)
	) name1793 (
		_w3426_,
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT3 #(
		.INIT('h20)
	) name1794 (
		\ctl_rf_c7_rf_chsad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4023_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1795 (
		\ctl_rf_c7_rf_chdad_reg[10]/P0002 ,
		\ctl_rf_c7_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4024_
	);
	LUT3 #(
		.INIT('h8a)
	) name1796 (
		_w3453_,
		_w4023_,
		_w4024_,
		_w4025_
	);
	LUT3 #(
		.INIT('h80)
	) name1797 (
		\ctl_rf_c6_rf_chdad_reg[10]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4026_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1798 (
		\ctl_rf_c6_rf_chsad_reg[10]/P0002 ,
		\ctl_rf_c6_rf_dwidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4027_
	);
	LUT3 #(
		.INIT('h8a)
	) name1799 (
		_w3440_,
		_w4026_,
		_w4027_,
		_w4028_
	);
	LUT4 #(
		.INIT('h0001)
	) name1800 (
		_w4019_,
		_w4022_,
		_w4025_,
		_w4028_,
		_w4029_
	);
	LUT4 #(
		.INIT('h8000)
	) name1801 (
		_w3424_,
		_w4003_,
		_w4016_,
		_w4029_,
		_w4030_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1802 (
		\hrdata_reg[26]_pad ,
		_w3422_,
		_w3689_,
		_w4030_,
		_w4031_
	);
	LUT4 #(
		.INIT('h0800)
	) name1803 (
		\ctl_rf_c5brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4032_
	);
	LUT4 #(
		.INIT('h2000)
	) name1804 (
		\ctl_rf_c6brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4033_
	);
	LUT4 #(
		.INIT('h0008)
	) name1805 (
		\ctl_rf_c1brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4034_
	);
	LUT4 #(
		.INIT('h0020)
	) name1806 (
		\ctl_rf_c2brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4035_
	);
	LUT4 #(
		.INIT('h0001)
	) name1807 (
		_w4032_,
		_w4033_,
		_w4034_,
		_w4035_,
		_w4036_
	);
	LUT4 #(
		.INIT('h0080)
	) name1808 (
		\ctl_rf_c3brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4037_
	);
	LUT4 #(
		.INIT('h0200)
	) name1809 (
		\ctl_rf_c4brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4038_
	);
	LUT4 #(
		.INIT('h0002)
	) name1810 (
		\ctl_rf_c0brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4039_
	);
	LUT4 #(
		.INIT('h8000)
	) name1811 (
		\ctl_rf_c7brbs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4040_
	);
	LUT4 #(
		.INIT('h0001)
	) name1812 (
		_w4037_,
		_w4038_,
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT3 #(
		.INIT('h2a)
	) name1813 (
		_w3425_,
		_w4036_,
		_w4041_,
		_w4042_
	);
	LUT4 #(
		.INIT('h0008)
	) name1814 (
		\ctl_rf_c1dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4043_
	);
	LUT4 #(
		.INIT('h2000)
	) name1815 (
		\ctl_rf_c6dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4044_
	);
	LUT4 #(
		.INIT('h0200)
	) name1816 (
		\ctl_rf_c4dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4045_
	);
	LUT4 #(
		.INIT('h0080)
	) name1817 (
		\ctl_rf_c3dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4046_
	);
	LUT4 #(
		.INIT('h0001)
	) name1818 (
		_w4043_,
		_w4044_,
		_w4045_,
		_w4046_,
		_w4047_
	);
	LUT4 #(
		.INIT('h0020)
	) name1819 (
		\ctl_rf_c2dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4048_
	);
	LUT4 #(
		.INIT('h0002)
	) name1820 (
		\ctl_rf_c0dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4049_
	);
	LUT4 #(
		.INIT('h0800)
	) name1821 (
		\ctl_rf_c5dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4050_
	);
	LUT4 #(
		.INIT('h8000)
	) name1822 (
		\ctl_rf_c7dmabs_reg[26]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4051_
	);
	LUT4 #(
		.INIT('h0001)
	) name1823 (
		_w4048_,
		_w4049_,
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT4 #(
		.INIT('h5111)
	) name1824 (
		\haddr[8]_pad ,
		_w3431_,
		_w4047_,
		_w4052_,
		_w4053_
	);
	LUT3 #(
		.INIT('h10)
	) name1825 (
		_w3503_,
		_w4042_,
		_w4053_,
		_w4054_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1826 (
		\ctl_rf_c3_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4055_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		_w3457_,
		_w4055_,
		_w4056_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1828 (
		\ctl_rf_c5_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4057_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1829 (
		\ctl_rf_c7_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4058_
	);
	LUT4 #(
		.INIT('hf531)
	) name1830 (
		_w3436_,
		_w3453_,
		_w4057_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h4)
	) name1831 (
		_w4056_,
		_w4059_,
		_w4060_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1832 (
		\ctl_rf_c2_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4061_
	);
	LUT3 #(
		.INIT('ha2)
	) name1833 (
		\haddr[8]_pad ,
		_w3432_,
		_w4061_,
		_w4062_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1834 (
		\ctl_rf_c0_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4063_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1835 (
		\ctl_rf_c6_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4064_
	);
	LUT4 #(
		.INIT('hf351)
	) name1836 (
		_w3440_,
		_w3445_,
		_w4063_,
		_w4064_,
		_w4065_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1837 (
		\ctl_rf_c1_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4066_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1838 (
		\ctl_rf_c4_rf_chdad_reg[26]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[26]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4067_
	);
	LUT4 #(
		.INIT('hf351)
	) name1839 (
		_w3426_,
		_w3449_,
		_w4066_,
		_w4067_,
		_w4068_
	);
	LUT3 #(
		.INIT('h80)
	) name1840 (
		_w4062_,
		_w4065_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name1841 (
		_w4060_,
		_w4069_,
		_w4070_
	);
	LUT4 #(
		.INIT('h135f)
	) name1842 (
		\ctl_rf_c0_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[26]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4071_
	);
	LUT4 #(
		.INIT('h135f)
	) name1843 (
		\ctl_rf_c1_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[26]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4072_
	);
	LUT4 #(
		.INIT('h135f)
	) name1844 (
		\ctl_rf_c5_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[26]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4073_
	);
	LUT4 #(
		.INIT('h135f)
	) name1845 (
		\ctl_rf_c2_rf_chllp_reg[26]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[26]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4074_
	);
	LUT4 #(
		.INIT('h8000)
	) name1846 (
		_w4071_,
		_w4072_,
		_w4073_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h31)
	) name1847 (
		_w3427_,
		_w3503_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('h15)
	) name1848 (
		_w4054_,
		_w4070_,
		_w4076_,
		_w4077_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1849 (
		\ctl_rf_c7_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4078_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1850 (
		\ctl_rf_c7_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4079_
	);
	LUT3 #(
		.INIT('h2a)
	) name1851 (
		_w3453_,
		_w4078_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1852 (
		\ctl_rf_c2_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4081_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1853 (
		\ctl_rf_c2_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4082_
	);
	LUT3 #(
		.INIT('h2a)
	) name1854 (
		_w3432_,
		_w4081_,
		_w4082_,
		_w4083_
	);
	LUT4 #(
		.INIT('hff53)
	) name1855 (
		\ctl_rf_c5_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c5_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4084_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1856 (
		\ctl_rf_c5_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4085_
	);
	LUT3 #(
		.INIT('h2a)
	) name1857 (
		_w3436_,
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1858 (
		\ctl_rf_c1_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4087_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1859 (
		\ctl_rf_c1_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4088_
	);
	LUT3 #(
		.INIT('h2a)
	) name1860 (
		_w3449_,
		_w4087_,
		_w4088_,
		_w4089_
	);
	LUT4 #(
		.INIT('h0001)
	) name1861 (
		_w4080_,
		_w4083_,
		_w4086_,
		_w4089_,
		_w4090_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1862 (
		\ctl_rf_c0_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4091_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1863 (
		\ctl_rf_c0_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4092_
	);
	LUT3 #(
		.INIT('h2a)
	) name1864 (
		_w3445_,
		_w4091_,
		_w4092_,
		_w4093_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1865 (
		\ctl_rf_c6_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4094_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1866 (
		\ctl_rf_c6_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4095_
	);
	LUT3 #(
		.INIT('h2a)
	) name1867 (
		_w3440_,
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT4 #(
		.INIT('hff53)
	) name1868 (
		\ctl_rf_c4_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c4_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4097_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1869 (
		\ctl_rf_c4_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c4_rf_chsad_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4098_
	);
	LUT3 #(
		.INIT('h2a)
	) name1870 (
		_w3426_,
		_w4097_,
		_w4098_,
		_w4099_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name1871 (
		\ctl_rf_c3_rf_chdad_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_int_abt_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4100_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1872 (
		\ctl_rf_c3_rf_chsad_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_src_sel_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4101_
	);
	LUT3 #(
		.INIT('h2a)
	) name1873 (
		_w3457_,
		_w4100_,
		_w4101_,
		_w4102_
	);
	LUT4 #(
		.INIT('h0001)
	) name1874 (
		_w4093_,
		_w4096_,
		_w4099_,
		_w4102_,
		_w4103_
	);
	LUT4 #(
		.INIT('hff35)
	) name1875 (
		\ctl_rf_c0_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4104_
	);
	LUT4 #(
		.INIT('hff35)
	) name1876 (
		\ctl_rf_c4_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4105_
	);
	LUT4 #(
		.INIT('hf531)
	) name1877 (
		_w3467_,
		_w3472_,
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('hff35)
	) name1878 (
		\ctl_rf_c1_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4107_
	);
	LUT4 #(
		.INIT('hff35)
	) name1879 (
		\ctl_rf_c2_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4108_
	);
	LUT4 #(
		.INIT('hf351)
	) name1880 (
		_w3462_,
		_w3474_,
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT4 #(
		.INIT('hff35)
	) name1881 (
		\ctl_rf_c7_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4110_
	);
	LUT4 #(
		.INIT('hff35)
	) name1882 (
		\ctl_rf_c5_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4111_
	);
	LUT4 #(
		.INIT('hf531)
	) name1883 (
		_w3464_,
		_w3469_,
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT4 #(
		.INIT('hff35)
	) name1884 (
		\ctl_rf_c3_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4113_
	);
	LUT4 #(
		.INIT('hff35)
	) name1885 (
		\ctl_rf_c6_rf_chllp_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[2]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4114_
	);
	LUT4 #(
		.INIT('hf531)
	) name1886 (
		_w3477_,
		_w3479_,
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT4 #(
		.INIT('h8000)
	) name1887 (
		_w4106_,
		_w4109_,
		_w4112_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1888 (
		\haddr[8]_pad ,
		_w4090_,
		_w4103_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h8)
	) name1889 (
		_w2534_,
		_w3486_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name1890 (
		\ctl_rf_c2_rf_int_tc1_msk_reg/NET0131 ,
		\haddr[4]_pad ,
		_w4119_
	);
	LUT3 #(
		.INIT('h08)
	) name1891 (
		\ctl_rf_tc_reg[2]/NET0131 ,
		_w3930_,
		_w4119_,
		_w4120_
	);
	LUT4 #(
		.INIT('h135f)
	) name1892 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_m1end_reg/NET0131 ,
		_w3492_,
		_w3494_,
		_w4121_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1893 (
		\ctl_rf_abt_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c2_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[2]/NET0131 ,
		_w4122_
	);
	LUT4 #(
		.INIT('h7707)
	) name1894 (
		\ctl_rf_sync_reg[2]/NET0131 ,
		_w3491_,
		_w3496_,
		_w4122_,
		_w4123_
	);
	LUT3 #(
		.INIT('h40)
	) name1895 (
		_w4120_,
		_w4121_,
		_w4123_,
		_w4124_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1896 (
		_w3484_,
		_w3503_,
		_w4118_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		_w4117_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w3424_,
		_w3990_,
		_w4127_
	);
	LUT4 #(
		.INIT('h0455)
	) name1899 (
		_w4031_,
		_w4077_,
		_w4126_,
		_w4127_,
		_w4128_
	);
	LUT3 #(
		.INIT('h2a)
	) name1900 (
		\hrdata_reg[27]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4129_
	);
	LUT3 #(
		.INIT('h20)
	) name1901 (
		\ctl_rf_c5_rf_chsad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4130_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1902 (
		\ctl_rf_c5_rf_chdad_reg[11]/P0002 ,
		\ctl_rf_c5_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4131_
	);
	LUT3 #(
		.INIT('h8a)
	) name1903 (
		_w3436_,
		_w4130_,
		_w4131_,
		_w4132_
	);
	LUT3 #(
		.INIT('h80)
	) name1904 (
		\ctl_rf_c0_rf_chdad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4133_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1905 (
		\ctl_rf_c0_rf_chsad_reg[11]/P0002 ,
		\ctl_rf_c0_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4134_
	);
	LUT3 #(
		.INIT('h8a)
	) name1906 (
		_w3445_,
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT3 #(
		.INIT('h80)
	) name1907 (
		\ctl_rf_c3_rf_chdad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4136_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1908 (
		\ctl_rf_c3_rf_chsad_reg[11]/P0002 ,
		\ctl_rf_c3_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4137_
	);
	LUT3 #(
		.INIT('h8a)
	) name1909 (
		_w3457_,
		_w4136_,
		_w4137_,
		_w4138_
	);
	LUT3 #(
		.INIT('h20)
	) name1910 (
		\ctl_rf_c2_rf_chsad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4139_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1911 (
		\ctl_rf_c2_rf_chdad_reg[11]/P0002 ,
		\ctl_rf_c2_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4140_
	);
	LUT3 #(
		.INIT('h8a)
	) name1912 (
		_w3432_,
		_w4139_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h0001)
	) name1913 (
		_w4132_,
		_w4135_,
		_w4138_,
		_w4141_,
		_w4142_
	);
	LUT4 #(
		.INIT('hff35)
	) name1914 (
		\ctl_rf_c3_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4143_
	);
	LUT4 #(
		.INIT('hff35)
	) name1915 (
		\ctl_rf_c2_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4144_
	);
	LUT4 #(
		.INIT('hf351)
	) name1916 (
		_w3462_,
		_w3477_,
		_w4143_,
		_w4144_,
		_w4145_
	);
	LUT4 #(
		.INIT('hff35)
	) name1917 (
		\ctl_rf_c1_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4146_
	);
	LUT4 #(
		.INIT('hff35)
	) name1918 (
		\ctl_rf_c0_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4147_
	);
	LUT4 #(
		.INIT('hf351)
	) name1919 (
		_w3467_,
		_w3474_,
		_w4146_,
		_w4147_,
		_w4148_
	);
	LUT4 #(
		.INIT('hff35)
	) name1920 (
		\ctl_rf_c5_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4149_
	);
	LUT4 #(
		.INIT('hff35)
	) name1921 (
		\ctl_rf_c4_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4150_
	);
	LUT4 #(
		.INIT('hf531)
	) name1922 (
		_w3469_,
		_w3472_,
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT4 #(
		.INIT('hff35)
	) name1923 (
		\ctl_rf_c6_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4152_
	);
	LUT4 #(
		.INIT('hff35)
	) name1924 (
		\ctl_rf_c7_rf_chllp_reg[11]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[11]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4153_
	);
	LUT4 #(
		.INIT('hf351)
	) name1925 (
		_w3464_,
		_w3479_,
		_w4152_,
		_w4153_,
		_w4154_
	);
	LUT4 #(
		.INIT('h8000)
	) name1926 (
		_w4145_,
		_w4148_,
		_w4151_,
		_w4154_,
		_w4155_
	);
	LUT3 #(
		.INIT('h20)
	) name1927 (
		\ctl_rf_c1_rf_chsad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4156_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1928 (
		\ctl_rf_c1_rf_chdad_reg[11]/P0002 ,
		\ctl_rf_c1_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4157_
	);
	LUT3 #(
		.INIT('h8a)
	) name1929 (
		_w3449_,
		_w4156_,
		_w4157_,
		_w4158_
	);
	LUT3 #(
		.INIT('h20)
	) name1930 (
		\ctl_rf_c4_rf_chsad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4159_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1931 (
		\ctl_rf_c4_rf_chdad_reg[11]/P0002 ,
		\ctl_rf_c4_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4160_
	);
	LUT3 #(
		.INIT('h8a)
	) name1932 (
		_w3426_,
		_w4159_,
		_w4160_,
		_w4161_
	);
	LUT3 #(
		.INIT('h20)
	) name1933 (
		\ctl_rf_c6_rf_chsad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4162_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1934 (
		\ctl_rf_c6_rf_chdad_reg[11]/P0002 ,
		\ctl_rf_c6_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4163_
	);
	LUT3 #(
		.INIT('h8a)
	) name1935 (
		_w3440_,
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT3 #(
		.INIT('h80)
	) name1936 (
		\ctl_rf_c7_rf_chdad_reg[11]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4165_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name1937 (
		\ctl_rf_c7_rf_chsad_reg[11]/P0002 ,
		\ctl_rf_c7_rf_swidth_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4166_
	);
	LUT3 #(
		.INIT('h8a)
	) name1938 (
		_w3453_,
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT4 #(
		.INIT('h0001)
	) name1939 (
		_w4158_,
		_w4161_,
		_w4164_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('h8000)
	) name1940 (
		_w3424_,
		_w4142_,
		_w4155_,
		_w4168_,
		_w4169_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1941 (
		\hrdata_reg[27]_pad ,
		_w3422_,
		_w3689_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h0800)
	) name1942 (
		\ctl_rf_c5dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4171_
	);
	LUT4 #(
		.INIT('h2000)
	) name1943 (
		\ctl_rf_c6dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4172_
	);
	LUT4 #(
		.INIT('h0008)
	) name1944 (
		\ctl_rf_c1dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4173_
	);
	LUT4 #(
		.INIT('h0020)
	) name1945 (
		\ctl_rf_c2dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4174_
	);
	LUT4 #(
		.INIT('h0001)
	) name1946 (
		_w4171_,
		_w4172_,
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT4 #(
		.INIT('h0080)
	) name1947 (
		\ctl_rf_c3dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4176_
	);
	LUT4 #(
		.INIT('h0200)
	) name1948 (
		\ctl_rf_c4dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4177_
	);
	LUT4 #(
		.INIT('h0002)
	) name1949 (
		\ctl_rf_c0dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4178_
	);
	LUT4 #(
		.INIT('h8000)
	) name1950 (
		\ctl_rf_c7dmabs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4179_
	);
	LUT4 #(
		.INIT('h0001)
	) name1951 (
		_w4176_,
		_w4177_,
		_w4178_,
		_w4179_,
		_w4180_
	);
	LUT3 #(
		.INIT('h2a)
	) name1952 (
		_w3431_,
		_w4175_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('h0008)
	) name1953 (
		\ctl_rf_c1brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4182_
	);
	LUT4 #(
		.INIT('h2000)
	) name1954 (
		\ctl_rf_c6brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4183_
	);
	LUT4 #(
		.INIT('h0200)
	) name1955 (
		\ctl_rf_c4brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4184_
	);
	LUT4 #(
		.INIT('h0080)
	) name1956 (
		\ctl_rf_c3brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4185_
	);
	LUT4 #(
		.INIT('h0001)
	) name1957 (
		_w4182_,
		_w4183_,
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('h0020)
	) name1958 (
		\ctl_rf_c2brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4187_
	);
	LUT4 #(
		.INIT('h0002)
	) name1959 (
		\ctl_rf_c0brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4188_
	);
	LUT4 #(
		.INIT('h0800)
	) name1960 (
		\ctl_rf_c5brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4189_
	);
	LUT4 #(
		.INIT('h8000)
	) name1961 (
		\ctl_rf_c7brbs_reg[27]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4190_
	);
	LUT4 #(
		.INIT('h0001)
	) name1962 (
		_w4187_,
		_w4188_,
		_w4189_,
		_w4190_,
		_w4191_
	);
	LUT4 #(
		.INIT('h5111)
	) name1963 (
		\haddr[8]_pad ,
		_w3425_,
		_w4186_,
		_w4191_,
		_w4192_
	);
	LUT3 #(
		.INIT('h10)
	) name1964 (
		_w3503_,
		_w4181_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1965 (
		\ctl_rf_c3_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		_w3457_,
		_w4194_,
		_w4195_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1967 (
		\ctl_rf_c5_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4196_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1968 (
		\ctl_rf_c6_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4197_
	);
	LUT4 #(
		.INIT('hf531)
	) name1969 (
		_w3436_,
		_w3440_,
		_w4196_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w4195_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1971 (
		\ctl_rf_c2_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4200_
	);
	LUT3 #(
		.INIT('ha2)
	) name1972 (
		\haddr[8]_pad ,
		_w3432_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1973 (
		\ctl_rf_c0_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4202_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1974 (
		\ctl_rf_c1_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4203_
	);
	LUT4 #(
		.INIT('hf531)
	) name1975 (
		_w3445_,
		_w3449_,
		_w4202_,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1976 (
		\ctl_rf_c4_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4205_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1977 (
		\ctl_rf_c7_rf_chdad_reg[27]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[27]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4206_
	);
	LUT4 #(
		.INIT('hf531)
	) name1978 (
		_w3426_,
		_w3453_,
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT3 #(
		.INIT('h80)
	) name1979 (
		_w4201_,
		_w4204_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w4199_,
		_w4208_,
		_w4209_
	);
	LUT4 #(
		.INIT('h135f)
	) name1981 (
		\ctl_rf_c0_rf_chllp_reg[27]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[27]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4210_
	);
	LUT4 #(
		.INIT('h135f)
	) name1982 (
		\ctl_rf_c1_rf_chllp_reg[27]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[27]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4211_
	);
	LUT4 #(
		.INIT('h135f)
	) name1983 (
		\ctl_rf_c5_rf_chllp_reg[27]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[27]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4212_
	);
	LUT4 #(
		.INIT('h135f)
	) name1984 (
		\ctl_rf_c2_rf_chllp_reg[27]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[27]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4213_
	);
	LUT4 #(
		.INIT('h8000)
	) name1985 (
		_w4210_,
		_w4211_,
		_w4212_,
		_w4213_,
		_w4214_
	);
	LUT3 #(
		.INIT('h31)
	) name1986 (
		_w3427_,
		_w3503_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h15)
	) name1987 (
		_w4193_,
		_w4209_,
		_w4215_,
		_w4216_
	);
	LUT3 #(
		.INIT('h20)
	) name1988 (
		\ctl_rf_c5_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4217_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1989 (
		\ctl_rf_c5_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c5_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4218_
	);
	LUT3 #(
		.INIT('h8a)
	) name1990 (
		_w3436_,
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT3 #(
		.INIT('h20)
	) name1991 (
		\ctl_rf_c3_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4220_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1992 (
		\ctl_rf_c3_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c3_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4221_
	);
	LUT3 #(
		.INIT('h8a)
	) name1993 (
		_w3457_,
		_w4220_,
		_w4221_,
		_w4222_
	);
	LUT3 #(
		.INIT('h20)
	) name1994 (
		\ctl_rf_c0_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4223_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1995 (
		\ctl_rf_c0_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c0_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4224_
	);
	LUT3 #(
		.INIT('h8a)
	) name1996 (
		_w3445_,
		_w4223_,
		_w4224_,
		_w4225_
	);
	LUT3 #(
		.INIT('h20)
	) name1997 (
		\ctl_rf_c2_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4226_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name1998 (
		\ctl_rf_c2_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c2_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4227_
	);
	LUT3 #(
		.INIT('h8a)
	) name1999 (
		_w3432_,
		_w4226_,
		_w4227_,
		_w4228_
	);
	LUT4 #(
		.INIT('h0001)
	) name2000 (
		_w4219_,
		_w4222_,
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT3 #(
		.INIT('h20)
	) name2001 (
		\ctl_rf_c7_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4230_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2002 (
		\ctl_rf_c7_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c7_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4231_
	);
	LUT3 #(
		.INIT('h8a)
	) name2003 (
		_w3453_,
		_w4230_,
		_w4231_,
		_w4232_
	);
	LUT3 #(
		.INIT('h20)
	) name2004 (
		\ctl_rf_c6_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4233_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2005 (
		\ctl_rf_c6_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c6_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4234_
	);
	LUT3 #(
		.INIT('h8a)
	) name2006 (
		_w3440_,
		_w4233_,
		_w4234_,
		_w4235_
	);
	LUT3 #(
		.INIT('h20)
	) name2007 (
		\ctl_rf_c1_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4236_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2008 (
		\ctl_rf_c1_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c1_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4237_
	);
	LUT3 #(
		.INIT('h8a)
	) name2009 (
		_w3449_,
		_w4236_,
		_w4237_,
		_w4238_
	);
	LUT3 #(
		.INIT('h20)
	) name2010 (
		\ctl_rf_c4_rf_chsad_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4239_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2011 (
		\ctl_rf_c4_rf_chdad_reg[3]/P0002 ,
		\ctl_rf_c4_rf_dad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4240_
	);
	LUT3 #(
		.INIT('h8a)
	) name2012 (
		_w3426_,
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT4 #(
		.INIT('h0001)
	) name2013 (
		_w4232_,
		_w4235_,
		_w4238_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('hff35)
	) name2014 (
		\ctl_rf_c2_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4243_
	);
	LUT4 #(
		.INIT('hff35)
	) name2015 (
		\ctl_rf_c7_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4244_
	);
	LUT4 #(
		.INIT('hf531)
	) name2016 (
		_w3462_,
		_w3464_,
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT4 #(
		.INIT('hff35)
	) name2017 (
		\ctl_rf_c4_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4246_
	);
	LUT4 #(
		.INIT('hff35)
	) name2018 (
		\ctl_rf_c3_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4247_
	);
	LUT4 #(
		.INIT('hf531)
	) name2019 (
		_w3472_,
		_w3477_,
		_w4246_,
		_w4247_,
		_w4248_
	);
	LUT4 #(
		.INIT('hff35)
	) name2020 (
		\ctl_rf_c6_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4249_
	);
	LUT4 #(
		.INIT('hff35)
	) name2021 (
		\ctl_rf_c5_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4250_
	);
	LUT4 #(
		.INIT('hf351)
	) name2022 (
		_w3469_,
		_w3479_,
		_w4249_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('hff35)
	) name2023 (
		\ctl_rf_c0_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4252_
	);
	LUT4 #(
		.INIT('hff35)
	) name2024 (
		\ctl_rf_c1_rf_chllp_reg[3]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[3]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4253_
	);
	LUT4 #(
		.INIT('hf531)
	) name2025 (
		_w3467_,
		_w3474_,
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h8000)
	) name2026 (
		_w4245_,
		_w4248_,
		_w4251_,
		_w4254_,
		_w4255_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2027 (
		\haddr[8]_pad ,
		_w4229_,
		_w4242_,
		_w4255_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		_w2534_,
		_w3927_,
		_w4257_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name2029 (
		\ctl_rf_c3_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[3]/NET0131 ,
		_w3488_,
		_w3489_,
		_w4258_
	);
	LUT2 #(
		.INIT('h2)
	) name2030 (
		\ctl_rf_abt_reg[3]/NET0131 ,
		\ctl_rf_c3_rf_int_abt_msk_reg/NET0131 ,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w3496_,
		_w4259_,
		_w4260_
	);
	LUT4 #(
		.INIT('h153f)
	) name2032 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[3]/NET0131 ,
		_w3491_,
		_w3492_,
		_w4261_
	);
	LUT3 #(
		.INIT('h20)
	) name2033 (
		_w4258_,
		_w4260_,
		_w4261_,
		_w4262_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2034 (
		_w3484_,
		_w3503_,
		_w4257_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h4)
	) name2035 (
		_w4256_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		_w3424_,
		_w4129_,
		_w4265_
	);
	LUT4 #(
		.INIT('h0455)
	) name2037 (
		_w4170_,
		_w4216_,
		_w4264_,
		_w4265_,
		_w4266_
	);
	LUT3 #(
		.INIT('h2a)
	) name2038 (
		\hrdata_reg[28]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4267_
	);
	LUT3 #(
		.INIT('h80)
	) name2039 (
		\ctl_rf_c0_rf_chdad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4268_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2040 (
		\ctl_rf_c0_rf_chsad_reg[12]/P0002 ,
		\ctl_rf_c0_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4269_
	);
	LUT3 #(
		.INIT('h8a)
	) name2041 (
		_w3445_,
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT3 #(
		.INIT('h20)
	) name2042 (
		\ctl_rf_c7_rf_chsad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4271_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2043 (
		\ctl_rf_c7_rf_chdad_reg[12]/P0002 ,
		\ctl_rf_c7_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4272_
	);
	LUT3 #(
		.INIT('h8a)
	) name2044 (
		_w3453_,
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT3 #(
		.INIT('h20)
	) name2045 (
		\ctl_rf_c6_rf_chsad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4274_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2046 (
		\ctl_rf_c6_rf_chdad_reg[12]/P0002 ,
		\ctl_rf_c6_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4275_
	);
	LUT3 #(
		.INIT('h8a)
	) name2047 (
		_w3440_,
		_w4274_,
		_w4275_,
		_w4276_
	);
	LUT3 #(
		.INIT('h80)
	) name2048 (
		\ctl_rf_c1_rf_chdad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4277_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2049 (
		\ctl_rf_c1_rf_chsad_reg[12]/P0002 ,
		\ctl_rf_c1_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4278_
	);
	LUT3 #(
		.INIT('h8a)
	) name2050 (
		_w3449_,
		_w4277_,
		_w4278_,
		_w4279_
	);
	LUT4 #(
		.INIT('h0001)
	) name2051 (
		_w4270_,
		_w4273_,
		_w4276_,
		_w4279_,
		_w4280_
	);
	LUT3 #(
		.INIT('h20)
	) name2052 (
		\ctl_rf_c5_rf_chsad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4281_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2053 (
		\ctl_rf_c5_rf_chdad_reg[12]/P0002 ,
		\ctl_rf_c5_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4282_
	);
	LUT3 #(
		.INIT('h8a)
	) name2054 (
		_w3436_,
		_w4281_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('h20)
	) name2055 (
		\ctl_rf_c2_rf_chsad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4284_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2056 (
		\ctl_rf_c2_rf_chdad_reg[12]/P0002 ,
		\ctl_rf_c2_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4285_
	);
	LUT3 #(
		.INIT('h8a)
	) name2057 (
		_w3432_,
		_w4284_,
		_w4285_,
		_w4286_
	);
	LUT3 #(
		.INIT('h20)
	) name2058 (
		\ctl_rf_c4_rf_chsad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4287_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2059 (
		\ctl_rf_c4_rf_chdad_reg[12]/P0002 ,
		\ctl_rf_c4_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4288_
	);
	LUT3 #(
		.INIT('h8a)
	) name2060 (
		_w3426_,
		_w4287_,
		_w4288_,
		_w4289_
	);
	LUT3 #(
		.INIT('h80)
	) name2061 (
		\ctl_rf_c3_rf_chdad_reg[12]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4290_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2062 (
		\ctl_rf_c3_rf_chsad_reg[12]/P0002 ,
		\ctl_rf_c3_rf_swidth_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4291_
	);
	LUT3 #(
		.INIT('h8a)
	) name2063 (
		_w3457_,
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT4 #(
		.INIT('h0001)
	) name2064 (
		_w4283_,
		_w4286_,
		_w4289_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		_w4280_,
		_w4293_,
		_w4294_
	);
	LUT4 #(
		.INIT('h135f)
	) name2066 (
		\ctl_rf_c5_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[12]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4295_
	);
	LUT4 #(
		.INIT('h135f)
	) name2067 (
		\ctl_rf_c1_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[12]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4296_
	);
	LUT4 #(
		.INIT('h153f)
	) name2068 (
		\ctl_rf_c0_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[12]/NET0131 ,
		_w3464_,
		_w3467_,
		_w4297_
	);
	LUT4 #(
		.INIT('h135f)
	) name2069 (
		\ctl_rf_c2_rf_chllp_reg[12]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[12]/NET0131 ,
		_w3462_,
		_w3472_,
		_w4298_
	);
	LUT4 #(
		.INIT('h8000)
	) name2070 (
		_w4295_,
		_w4296_,
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT3 #(
		.INIT('ha2)
	) name2071 (
		_w3424_,
		_w3427_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('h0222)
	) name2072 (
		_w3422_,
		_w3689_,
		_w4294_,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w4267_,
		_w4301_,
		_w4302_
	);
	LUT4 #(
		.INIT('h0800)
	) name2074 (
		\ctl_rf_c5dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4303_
	);
	LUT4 #(
		.INIT('h2000)
	) name2075 (
		\ctl_rf_c6dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4304_
	);
	LUT4 #(
		.INIT('h0008)
	) name2076 (
		\ctl_rf_c1dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4305_
	);
	LUT4 #(
		.INIT('h0020)
	) name2077 (
		\ctl_rf_c2dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4306_
	);
	LUT4 #(
		.INIT('h0001)
	) name2078 (
		_w4303_,
		_w4304_,
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT4 #(
		.INIT('h0080)
	) name2079 (
		\ctl_rf_c3dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4308_
	);
	LUT4 #(
		.INIT('h0200)
	) name2080 (
		\ctl_rf_c4dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4309_
	);
	LUT4 #(
		.INIT('h0002)
	) name2081 (
		\ctl_rf_c0dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4310_
	);
	LUT4 #(
		.INIT('h8000)
	) name2082 (
		\ctl_rf_c7dmabs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4311_
	);
	LUT4 #(
		.INIT('h0001)
	) name2083 (
		_w4308_,
		_w4309_,
		_w4310_,
		_w4311_,
		_w4312_
	);
	LUT3 #(
		.INIT('h2a)
	) name2084 (
		_w3431_,
		_w4307_,
		_w4312_,
		_w4313_
	);
	LUT4 #(
		.INIT('h0008)
	) name2085 (
		\ctl_rf_c1brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4314_
	);
	LUT4 #(
		.INIT('h2000)
	) name2086 (
		\ctl_rf_c6brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4315_
	);
	LUT4 #(
		.INIT('h0200)
	) name2087 (
		\ctl_rf_c4brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4316_
	);
	LUT4 #(
		.INIT('h0080)
	) name2088 (
		\ctl_rf_c3brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4317_
	);
	LUT4 #(
		.INIT('h0001)
	) name2089 (
		_w4314_,
		_w4315_,
		_w4316_,
		_w4317_,
		_w4318_
	);
	LUT4 #(
		.INIT('h0020)
	) name2090 (
		\ctl_rf_c2brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4319_
	);
	LUT4 #(
		.INIT('h0002)
	) name2091 (
		\ctl_rf_c0brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4320_
	);
	LUT4 #(
		.INIT('h0800)
	) name2092 (
		\ctl_rf_c5brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4321_
	);
	LUT4 #(
		.INIT('h8000)
	) name2093 (
		\ctl_rf_c7brbs_reg[28]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4322_
	);
	LUT4 #(
		.INIT('h0001)
	) name2094 (
		_w4319_,
		_w4320_,
		_w4321_,
		_w4322_,
		_w4323_
	);
	LUT4 #(
		.INIT('h5111)
	) name2095 (
		\haddr[8]_pad ,
		_w3425_,
		_w4318_,
		_w4323_,
		_w4324_
	);
	LUT3 #(
		.INIT('h10)
	) name2096 (
		_w3503_,
		_w4313_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2097 (
		\ctl_rf_c3_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4326_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		_w3457_,
		_w4326_,
		_w4327_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2099 (
		\ctl_rf_c5_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4328_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2100 (
		\ctl_rf_c6_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4329_
	);
	LUT4 #(
		.INIT('hf531)
	) name2101 (
		_w3436_,
		_w3440_,
		_w4328_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h4)
	) name2102 (
		_w4327_,
		_w4330_,
		_w4331_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2103 (
		\ctl_rf_c0_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4332_
	);
	LUT3 #(
		.INIT('ha2)
	) name2104 (
		\haddr[8]_pad ,
		_w3445_,
		_w4332_,
		_w4333_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2105 (
		\ctl_rf_c2_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4334_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2106 (
		\ctl_rf_c4_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4335_
	);
	LUT4 #(
		.INIT('hf351)
	) name2107 (
		_w3426_,
		_w3432_,
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2108 (
		\ctl_rf_c1_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4337_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2109 (
		\ctl_rf_c7_rf_chdad_reg[28]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[28]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4338_
	);
	LUT4 #(
		.INIT('hf531)
	) name2110 (
		_w3449_,
		_w3453_,
		_w4337_,
		_w4338_,
		_w4339_
	);
	LUT3 #(
		.INIT('h80)
	) name2111 (
		_w4333_,
		_w4336_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		_w4331_,
		_w4340_,
		_w4341_
	);
	LUT4 #(
		.INIT('h135f)
	) name2113 (
		\ctl_rf_c0_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[28]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4342_
	);
	LUT4 #(
		.INIT('h135f)
	) name2114 (
		\ctl_rf_c1_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[28]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4343_
	);
	LUT4 #(
		.INIT('h135f)
	) name2115 (
		\ctl_rf_c5_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[28]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4344_
	);
	LUT4 #(
		.INIT('h135f)
	) name2116 (
		\ctl_rf_c2_rf_chllp_reg[28]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[28]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4345_
	);
	LUT4 #(
		.INIT('h8000)
	) name2117 (
		_w4342_,
		_w4343_,
		_w4344_,
		_w4345_,
		_w4346_
	);
	LUT3 #(
		.INIT('h31)
	) name2118 (
		_w3427_,
		_w3503_,
		_w4346_,
		_w4347_
	);
	LUT3 #(
		.INIT('h15)
	) name2119 (
		_w4325_,
		_w4341_,
		_w4347_,
		_w4348_
	);
	LUT3 #(
		.INIT('h20)
	) name2120 (
		\ctl_rf_c4_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4349_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2121 (
		\ctl_rf_c4_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c4_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4350_
	);
	LUT3 #(
		.INIT('h8a)
	) name2122 (
		_w3426_,
		_w4349_,
		_w4350_,
		_w4351_
	);
	LUT3 #(
		.INIT('h20)
	) name2123 (
		\ctl_rf_c6_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4352_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2124 (
		\ctl_rf_c6_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c6_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4353_
	);
	LUT3 #(
		.INIT('h8a)
	) name2125 (
		_w3440_,
		_w4352_,
		_w4353_,
		_w4354_
	);
	LUT3 #(
		.INIT('h20)
	) name2126 (
		\ctl_rf_c7_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4355_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2127 (
		\ctl_rf_c7_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c7_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4356_
	);
	LUT3 #(
		.INIT('h8a)
	) name2128 (
		_w3453_,
		_w4355_,
		_w4356_,
		_w4357_
	);
	LUT3 #(
		.INIT('h20)
	) name2129 (
		\ctl_rf_c1_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4358_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2130 (
		\ctl_rf_c1_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c1_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4359_
	);
	LUT3 #(
		.INIT('h8a)
	) name2131 (
		_w3449_,
		_w4358_,
		_w4359_,
		_w4360_
	);
	LUT4 #(
		.INIT('h0001)
	) name2132 (
		_w4351_,
		_w4354_,
		_w4357_,
		_w4360_,
		_w4361_
	);
	LUT3 #(
		.INIT('h20)
	) name2133 (
		\ctl_rf_c0_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4362_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2134 (
		\ctl_rf_c0_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c0_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4363_
	);
	LUT3 #(
		.INIT('h8a)
	) name2135 (
		_w3445_,
		_w4362_,
		_w4363_,
		_w4364_
	);
	LUT3 #(
		.INIT('h20)
	) name2136 (
		\ctl_rf_c5_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4365_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2137 (
		\ctl_rf_c5_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c5_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4366_
	);
	LUT3 #(
		.INIT('h8a)
	) name2138 (
		_w3436_,
		_w4365_,
		_w4366_,
		_w4367_
	);
	LUT3 #(
		.INIT('h20)
	) name2139 (
		\ctl_rf_c3_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4368_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2140 (
		\ctl_rf_c3_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c3_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4369_
	);
	LUT3 #(
		.INIT('h8a)
	) name2141 (
		_w3457_,
		_w4368_,
		_w4369_,
		_w4370_
	);
	LUT3 #(
		.INIT('h20)
	) name2142 (
		\ctl_rf_c2_rf_chsad_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4371_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2143 (
		\ctl_rf_c2_rf_chdad_reg[4]/P0002 ,
		\ctl_rf_c2_rf_dad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4372_
	);
	LUT3 #(
		.INIT('h8a)
	) name2144 (
		_w3432_,
		_w4371_,
		_w4372_,
		_w4373_
	);
	LUT4 #(
		.INIT('h0001)
	) name2145 (
		_w4364_,
		_w4367_,
		_w4370_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('hff35)
	) name2146 (
		\ctl_rf_c7_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4375_
	);
	LUT4 #(
		.INIT('hff35)
	) name2147 (
		\ctl_rf_c2_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4376_
	);
	LUT4 #(
		.INIT('hf351)
	) name2148 (
		_w3462_,
		_w3464_,
		_w4375_,
		_w4376_,
		_w4377_
	);
	LUT4 #(
		.INIT('hff35)
	) name2149 (
		\ctl_rf_c1_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4378_
	);
	LUT4 #(
		.INIT('hff35)
	) name2150 (
		\ctl_rf_c0_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4379_
	);
	LUT4 #(
		.INIT('hf351)
	) name2151 (
		_w3467_,
		_w3474_,
		_w4378_,
		_w4379_,
		_w4380_
	);
	LUT4 #(
		.INIT('hff35)
	) name2152 (
		\ctl_rf_c5_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4381_
	);
	LUT4 #(
		.INIT('hff35)
	) name2153 (
		\ctl_rf_c6_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4382_
	);
	LUT4 #(
		.INIT('hf531)
	) name2154 (
		_w3469_,
		_w3479_,
		_w4381_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('hff35)
	) name2155 (
		\ctl_rf_c3_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4384_
	);
	LUT4 #(
		.INIT('hff35)
	) name2156 (
		\ctl_rf_c4_rf_chllp_reg[4]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[4]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4385_
	);
	LUT4 #(
		.INIT('hf351)
	) name2157 (
		_w3472_,
		_w3477_,
		_w4384_,
		_w4385_,
		_w4386_
	);
	LUT4 #(
		.INIT('h8000)
	) name2158 (
		_w4377_,
		_w4380_,
		_w4383_,
		_w4386_,
		_w4387_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2159 (
		\haddr[8]_pad ,
		_w4361_,
		_w4374_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		_w2520_,
		_w3486_,
		_w4389_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name2161 (
		\ctl_rf_c4_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[4]/NET0131 ,
		_w3488_,
		_w3489_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name2162 (
		\ctl_rf_abt_reg[4]/NET0131 ,
		\ctl_rf_c4_rf_int_abt_msk_reg/NET0131 ,
		_w4391_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		_w3496_,
		_w4391_,
		_w4392_
	);
	LUT4 #(
		.INIT('h153f)
	) name2164 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[4]/NET0131 ,
		_w3491_,
		_w3492_,
		_w4393_
	);
	LUT3 #(
		.INIT('h20)
	) name2165 (
		_w4390_,
		_w4392_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2166 (
		_w3484_,
		_w3503_,
		_w4389_,
		_w4394_,
		_w4395_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		_w4388_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w3424_,
		_w4267_,
		_w4397_
	);
	LUT3 #(
		.INIT('hd0)
	) name2169 (
		_w4348_,
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w4302_,
		_w4398_,
		_w4399_
	);
	LUT3 #(
		.INIT('h2a)
	) name2171 (
		\hrdata_reg[29]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4400_
	);
	LUT3 #(
		.INIT('h80)
	) name2172 (
		\ctl_rf_c7_rf_chdad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4401_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2173 (
		\ctl_rf_c7_rf_chsad_reg[13]/P0002 ,
		\ctl_rf_c7_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4402_
	);
	LUT3 #(
		.INIT('h8a)
	) name2174 (
		_w3453_,
		_w4401_,
		_w4402_,
		_w4403_
	);
	LUT3 #(
		.INIT('h20)
	) name2175 (
		\ctl_rf_c0_rf_chsad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4404_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2176 (
		\ctl_rf_c0_rf_chdad_reg[13]/P0002 ,
		\ctl_rf_c0_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4405_
	);
	LUT3 #(
		.INIT('h8a)
	) name2177 (
		_w3445_,
		_w4404_,
		_w4405_,
		_w4406_
	);
	LUT3 #(
		.INIT('h20)
	) name2178 (
		\ctl_rf_c3_rf_chsad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4407_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2179 (
		\ctl_rf_c3_rf_chdad_reg[13]/P0002 ,
		\ctl_rf_c3_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4408_
	);
	LUT3 #(
		.INIT('h8a)
	) name2180 (
		_w3457_,
		_w4407_,
		_w4408_,
		_w4409_
	);
	LUT3 #(
		.INIT('h80)
	) name2181 (
		\ctl_rf_c5_rf_chdad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4410_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2182 (
		\ctl_rf_c5_rf_chsad_reg[13]/P0002 ,
		\ctl_rf_c5_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4411_
	);
	LUT3 #(
		.INIT('h8a)
	) name2183 (
		_w3436_,
		_w4410_,
		_w4411_,
		_w4412_
	);
	LUT4 #(
		.INIT('h0001)
	) name2184 (
		_w4403_,
		_w4406_,
		_w4409_,
		_w4412_,
		_w4413_
	);
	LUT3 #(
		.INIT('h80)
	) name2185 (
		\ctl_rf_c6_rf_chdad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4414_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2186 (
		\ctl_rf_c6_rf_chsad_reg[13]/P0002 ,
		\ctl_rf_c6_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4415_
	);
	LUT3 #(
		.INIT('h8a)
	) name2187 (
		_w3440_,
		_w4414_,
		_w4415_,
		_w4416_
	);
	LUT3 #(
		.INIT('h20)
	) name2188 (
		\ctl_rf_c4_rf_chsad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4417_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2189 (
		\ctl_rf_c4_rf_chdad_reg[13]/P0002 ,
		\ctl_rf_c4_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4418_
	);
	LUT3 #(
		.INIT('h8a)
	) name2190 (
		_w3426_,
		_w4417_,
		_w4418_,
		_w4419_
	);
	LUT3 #(
		.INIT('h20)
	) name2191 (
		\ctl_rf_c2_rf_chsad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4420_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2192 (
		\ctl_rf_c2_rf_chdad_reg[13]/P0002 ,
		\ctl_rf_c2_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4421_
	);
	LUT3 #(
		.INIT('h8a)
	) name2193 (
		_w3432_,
		_w4420_,
		_w4421_,
		_w4422_
	);
	LUT3 #(
		.INIT('h80)
	) name2194 (
		\ctl_rf_c1_rf_chdad_reg[13]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4423_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2195 (
		\ctl_rf_c1_rf_chsad_reg[13]/P0002 ,
		\ctl_rf_c1_rf_swidth_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4424_
	);
	LUT3 #(
		.INIT('h8a)
	) name2196 (
		_w3449_,
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT4 #(
		.INIT('h0001)
	) name2197 (
		_w4416_,
		_w4419_,
		_w4422_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		_w4413_,
		_w4426_,
		_w4427_
	);
	LUT4 #(
		.INIT('h153f)
	) name2199 (
		\ctl_rf_c1_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[13]/NET0131 ,
		_w3472_,
		_w3474_,
		_w4428_
	);
	LUT4 #(
		.INIT('h135f)
	) name2200 (
		\ctl_rf_c2_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[13]/NET0131 ,
		_w3462_,
		_w3479_,
		_w4429_
	);
	LUT4 #(
		.INIT('h153f)
	) name2201 (
		\ctl_rf_c0_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[13]/NET0131 ,
		_w3464_,
		_w3467_,
		_w4430_
	);
	LUT4 #(
		.INIT('h153f)
	) name2202 (
		\ctl_rf_c3_rf_chllp_reg[13]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[13]/NET0131 ,
		_w3469_,
		_w3477_,
		_w4431_
	);
	LUT4 #(
		.INIT('h8000)
	) name2203 (
		_w4428_,
		_w4429_,
		_w4430_,
		_w4431_,
		_w4432_
	);
	LUT3 #(
		.INIT('ha2)
	) name2204 (
		_w3424_,
		_w3427_,
		_w4432_,
		_w4433_
	);
	LUT4 #(
		.INIT('h0222)
	) name2205 (
		_w3422_,
		_w3689_,
		_w4427_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w4400_,
		_w4434_,
		_w4435_
	);
	LUT4 #(
		.INIT('h0800)
	) name2207 (
		\ctl_rf_c5dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4436_
	);
	LUT4 #(
		.INIT('h2000)
	) name2208 (
		\ctl_rf_c6dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4437_
	);
	LUT4 #(
		.INIT('h0008)
	) name2209 (
		\ctl_rf_c1dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4438_
	);
	LUT4 #(
		.INIT('h0020)
	) name2210 (
		\ctl_rf_c2dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4439_
	);
	LUT4 #(
		.INIT('h0001)
	) name2211 (
		_w4436_,
		_w4437_,
		_w4438_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h0080)
	) name2212 (
		\ctl_rf_c3dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4441_
	);
	LUT4 #(
		.INIT('h0200)
	) name2213 (
		\ctl_rf_c4dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4442_
	);
	LUT4 #(
		.INIT('h0002)
	) name2214 (
		\ctl_rf_c0dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4443_
	);
	LUT4 #(
		.INIT('h8000)
	) name2215 (
		\ctl_rf_c7dmabs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4444_
	);
	LUT4 #(
		.INIT('h0001)
	) name2216 (
		_w4441_,
		_w4442_,
		_w4443_,
		_w4444_,
		_w4445_
	);
	LUT3 #(
		.INIT('h2a)
	) name2217 (
		_w3431_,
		_w4440_,
		_w4445_,
		_w4446_
	);
	LUT4 #(
		.INIT('h0008)
	) name2218 (
		\ctl_rf_c1brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4447_
	);
	LUT4 #(
		.INIT('h2000)
	) name2219 (
		\ctl_rf_c6brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4448_
	);
	LUT4 #(
		.INIT('h0200)
	) name2220 (
		\ctl_rf_c4brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4449_
	);
	LUT4 #(
		.INIT('h0080)
	) name2221 (
		\ctl_rf_c3brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4450_
	);
	LUT4 #(
		.INIT('h0001)
	) name2222 (
		_w4447_,
		_w4448_,
		_w4449_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h0020)
	) name2223 (
		\ctl_rf_c2brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4452_
	);
	LUT4 #(
		.INIT('h0002)
	) name2224 (
		\ctl_rf_c0brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4453_
	);
	LUT4 #(
		.INIT('h0800)
	) name2225 (
		\ctl_rf_c5brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4454_
	);
	LUT4 #(
		.INIT('h8000)
	) name2226 (
		\ctl_rf_c7brbs_reg[29]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4455_
	);
	LUT4 #(
		.INIT('h0001)
	) name2227 (
		_w4452_,
		_w4453_,
		_w4454_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('h5111)
	) name2228 (
		\haddr[8]_pad ,
		_w3425_,
		_w4451_,
		_w4456_,
		_w4457_
	);
	LUT3 #(
		.INIT('h10)
	) name2229 (
		_w3503_,
		_w4446_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2230 (
		\ctl_rf_c6_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4459_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		_w3440_,
		_w4459_,
		_w4460_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2232 (
		\ctl_rf_c7_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4461_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2233 (
		\ctl_rf_c3_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4462_
	);
	LUT4 #(
		.INIT('hf531)
	) name2234 (
		_w3453_,
		_w3457_,
		_w4461_,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h4)
	) name2235 (
		_w4460_,
		_w4463_,
		_w4464_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2236 (
		\ctl_rf_c1_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4465_
	);
	LUT3 #(
		.INIT('ha2)
	) name2237 (
		\haddr[8]_pad ,
		_w3449_,
		_w4465_,
		_w4466_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2238 (
		\ctl_rf_c4_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4467_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2239 (
		\ctl_rf_c2_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4468_
	);
	LUT4 #(
		.INIT('hf531)
	) name2240 (
		_w3426_,
		_w3432_,
		_w4467_,
		_w4468_,
		_w4469_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2241 (
		\ctl_rf_c0_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4470_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2242 (
		\ctl_rf_c5_rf_chdad_reg[29]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[29]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4471_
	);
	LUT4 #(
		.INIT('hf351)
	) name2243 (
		_w3436_,
		_w3445_,
		_w4470_,
		_w4471_,
		_w4472_
	);
	LUT3 #(
		.INIT('h80)
	) name2244 (
		_w4466_,
		_w4469_,
		_w4472_,
		_w4473_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		_w4464_,
		_w4473_,
		_w4474_
	);
	LUT4 #(
		.INIT('h135f)
	) name2246 (
		\ctl_rf_c1_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[29]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4475_
	);
	LUT4 #(
		.INIT('h135f)
	) name2247 (
		\ctl_rf_c0_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[29]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4476_
	);
	LUT4 #(
		.INIT('h135f)
	) name2248 (
		\ctl_rf_c5_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[29]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4477_
	);
	LUT4 #(
		.INIT('h135f)
	) name2249 (
		\ctl_rf_c2_rf_chllp_reg[29]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[29]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4478_
	);
	LUT4 #(
		.INIT('h8000)
	) name2250 (
		_w4475_,
		_w4476_,
		_w4477_,
		_w4478_,
		_w4479_
	);
	LUT3 #(
		.INIT('h31)
	) name2251 (
		_w3427_,
		_w3503_,
		_w4479_,
		_w4480_
	);
	LUT3 #(
		.INIT('h15)
	) name2252 (
		_w4458_,
		_w4474_,
		_w4480_,
		_w4481_
	);
	LUT3 #(
		.INIT('h20)
	) name2253 (
		\ctl_rf_c2_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4482_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2254 (
		\ctl_rf_c2_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c2_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4483_
	);
	LUT3 #(
		.INIT('h8a)
	) name2255 (
		_w3432_,
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT3 #(
		.INIT('h20)
	) name2256 (
		\ctl_rf_c3_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4485_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2257 (
		\ctl_rf_c3_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c3_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4486_
	);
	LUT3 #(
		.INIT('h8a)
	) name2258 (
		_w3457_,
		_w4485_,
		_w4486_,
		_w4487_
	);
	LUT3 #(
		.INIT('h20)
	) name2259 (
		\ctl_rf_c0_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4488_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2260 (
		\ctl_rf_c0_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c0_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4489_
	);
	LUT3 #(
		.INIT('h8a)
	) name2261 (
		_w3445_,
		_w4488_,
		_w4489_,
		_w4490_
	);
	LUT3 #(
		.INIT('h20)
	) name2262 (
		\ctl_rf_c5_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4491_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2263 (
		\ctl_rf_c5_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c5_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4492_
	);
	LUT3 #(
		.INIT('h8a)
	) name2264 (
		_w3436_,
		_w4491_,
		_w4492_,
		_w4493_
	);
	LUT4 #(
		.INIT('h0001)
	) name2265 (
		_w4484_,
		_w4487_,
		_w4490_,
		_w4493_,
		_w4494_
	);
	LUT3 #(
		.INIT('h20)
	) name2266 (
		\ctl_rf_c4_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4495_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2267 (
		\ctl_rf_c4_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c4_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4496_
	);
	LUT3 #(
		.INIT('h8a)
	) name2268 (
		_w3426_,
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT3 #(
		.INIT('h20)
	) name2269 (
		\ctl_rf_c6_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4498_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2270 (
		\ctl_rf_c6_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c6_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4499_
	);
	LUT3 #(
		.INIT('h8a)
	) name2271 (
		_w3440_,
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h20)
	) name2272 (
		\ctl_rf_c7_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4501_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2273 (
		\ctl_rf_c7_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c7_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4502_
	);
	LUT3 #(
		.INIT('h8a)
	) name2274 (
		_w3453_,
		_w4501_,
		_w4502_,
		_w4503_
	);
	LUT3 #(
		.INIT('h20)
	) name2275 (
		\ctl_rf_c1_rf_chsad_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4504_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2276 (
		\ctl_rf_c1_rf_chdad_reg[5]/P0002 ,
		\ctl_rf_c1_rf_sad_ctl0_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4505_
	);
	LUT3 #(
		.INIT('h8a)
	) name2277 (
		_w3449_,
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT4 #(
		.INIT('h0001)
	) name2278 (
		_w4497_,
		_w4500_,
		_w4503_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('hff35)
	) name2279 (
		\ctl_rf_c0_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4508_
	);
	LUT4 #(
		.INIT('hff35)
	) name2280 (
		\ctl_rf_c7_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4509_
	);
	LUT4 #(
		.INIT('hf351)
	) name2281 (
		_w3464_,
		_w3467_,
		_w4508_,
		_w4509_,
		_w4510_
	);
	LUT4 #(
		.INIT('hff35)
	) name2282 (
		\ctl_rf_c4_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4511_
	);
	LUT4 #(
		.INIT('hff35)
	) name2283 (
		\ctl_rf_c3_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4512_
	);
	LUT4 #(
		.INIT('hf531)
	) name2284 (
		_w3472_,
		_w3477_,
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT4 #(
		.INIT('hff35)
	) name2285 (
		\ctl_rf_c6_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4514_
	);
	LUT4 #(
		.INIT('hff35)
	) name2286 (
		\ctl_rf_c2_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4515_
	);
	LUT4 #(
		.INIT('hf351)
	) name2287 (
		_w3462_,
		_w3479_,
		_w4514_,
		_w4515_,
		_w4516_
	);
	LUT4 #(
		.INIT('hff35)
	) name2288 (
		\ctl_rf_c1_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4517_
	);
	LUT4 #(
		.INIT('hff35)
	) name2289 (
		\ctl_rf_c5_rf_chllp_reg[5]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[5]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4518_
	);
	LUT4 #(
		.INIT('hf351)
	) name2290 (
		_w3469_,
		_w3474_,
		_w4517_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('h8000)
	) name2291 (
		_w4510_,
		_w4513_,
		_w4516_,
		_w4519_,
		_w4520_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2292 (
		\haddr[8]_pad ,
		_w4494_,
		_w4507_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h8)
	) name2293 (
		_w2520_,
		_w3927_,
		_w4522_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name2294 (
		\ctl_rf_c5_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[5]/NET0131 ,
		_w3488_,
		_w3489_,
		_w4523_
	);
	LUT2 #(
		.INIT('h2)
	) name2295 (
		\ctl_rf_abt_reg[5]/NET0131 ,
		\ctl_rf_c5_rf_int_abt_msk_reg/NET0131 ,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		_w3496_,
		_w4524_,
		_w4525_
	);
	LUT4 #(
		.INIT('h153f)
	) name2297 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[5]/NET0131 ,
		_w3491_,
		_w3492_,
		_w4526_
	);
	LUT3 #(
		.INIT('h20)
	) name2298 (
		_w4523_,
		_w4525_,
		_w4526_,
		_w4527_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2299 (
		_w3484_,
		_w3503_,
		_w4522_,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name2300 (
		_w4521_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w3424_,
		_w4400_,
		_w4530_
	);
	LUT3 #(
		.INIT('hd0)
	) name2302 (
		_w4481_,
		_w4529_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w4435_,
		_w4531_,
		_w4532_
	);
	LUT3 #(
		.INIT('h2a)
	) name2304 (
		\hrdata_reg[2]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4533_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2305 (
		\ctl_rf_c0_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4534_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2306 (
		\ctl_rf_c0_rf_chsad_reg[18]/NET0131 ,
		\ctl_rf_c0_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4535_
	);
	LUT4 #(
		.INIT('ha222)
	) name2307 (
		\haddr[8]_pad ,
		_w3445_,
		_w4534_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('hf35f)
	) name2308 (
		\ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_chsad_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4537_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2309 (
		\ctl_rf_c2_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c2_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4538_
	);
	LUT3 #(
		.INIT('h2a)
	) name2310 (
		_w3432_,
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2311 (
		\ctl_rf_c6_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4540_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2312 (
		\ctl_rf_c6_rf_chsad_reg[18]/NET0131 ,
		\ctl_rf_c6_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4541_
	);
	LUT3 #(
		.INIT('h2a)
	) name2313 (
		_w3440_,
		_w4540_,
		_w4541_,
		_w4542_
	);
	LUT4 #(
		.INIT('hff53)
	) name2314 (
		\ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4543_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2315 (
		\ctl_rf_c1_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4544_
	);
	LUT3 #(
		.INIT('h2a)
	) name2316 (
		_w3449_,
		_w4543_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('hff53)
	) name2317 (
		\ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4546_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2318 (
		\ctl_rf_c7_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4547_
	);
	LUT3 #(
		.INIT('h2a)
	) name2319 (
		_w3453_,
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h0001)
	) name2320 (
		_w4539_,
		_w4542_,
		_w4545_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		_w4536_,
		_w4549_,
		_w4550_
	);
	LUT4 #(
		.INIT('h153f)
	) name2322 (
		\ctl_rf_c3_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[18]/NET0131 ,
		_w3469_,
		_w3477_,
		_w4551_
	);
	LUT4 #(
		.INIT('h135f)
	) name2323 (
		\ctl_rf_c0_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[18]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4552_
	);
	LUT4 #(
		.INIT('h135f)
	) name2324 (
		\ctl_rf_c2_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[18]/NET0131 ,
		_w3462_,
		_w3479_,
		_w4553_
	);
	LUT4 #(
		.INIT('h153f)
	) name2325 (
		\ctl_rf_c1_rf_chllp_reg[18]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[18]/NET0131 ,
		_w3464_,
		_w3474_,
		_w4554_
	);
	LUT4 #(
		.INIT('h8000)
	) name2326 (
		_w4551_,
		_w4552_,
		_w4553_,
		_w4554_,
		_w4555_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2327 (
		\ctl_rf_c4_rf_chsad_reg[18]/NET0131 ,
		\ctl_rf_c4_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4556_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2328 (
		\ctl_rf_c4_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4557_
	);
	LUT3 #(
		.INIT('h2a)
	) name2329 (
		_w3426_,
		_w4556_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('hff53)
	) name2330 (
		\ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4559_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2331 (
		\ctl_rf_c5_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4560_
	);
	LUT3 #(
		.INIT('h2a)
	) name2332 (
		_w3436_,
		_w4559_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2333 (
		\ctl_rf_c3_rf_chdad_reg[18]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4562_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2334 (
		\ctl_rf_c3_rf_chsad_reg[18]/NET0131 ,
		\ctl_rf_c3_rf_src_sz_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4563_
	);
	LUT3 #(
		.INIT('h2a)
	) name2335 (
		_w3457_,
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT3 #(
		.INIT('h01)
	) name2336 (
		_w4558_,
		_w4561_,
		_w4564_,
		_w4565_
	);
	LUT3 #(
		.INIT('hd0)
	) name2337 (
		_w3427_,
		_w4555_,
		_w4565_,
		_w4566_
	);
	LUT4 #(
		.INIT('h0008)
	) name2338 (
		\ctl_rf_c1brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4567_
	);
	LUT4 #(
		.INIT('h0080)
	) name2339 (
		\ctl_rf_c3brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4568_
	);
	LUT4 #(
		.INIT('h0002)
	) name2340 (
		\ctl_rf_c0brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4569_
	);
	LUT4 #(
		.INIT('h8000)
	) name2341 (
		\ctl_rf_c7brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4570_
	);
	LUT4 #(
		.INIT('h0001)
	) name2342 (
		_w4567_,
		_w4568_,
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT4 #(
		.INIT('h2000)
	) name2343 (
		\ctl_rf_c6brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4572_
	);
	LUT4 #(
		.INIT('h0200)
	) name2344 (
		\ctl_rf_c4brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4573_
	);
	LUT4 #(
		.INIT('h0020)
	) name2345 (
		\ctl_rf_c2brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4574_
	);
	LUT4 #(
		.INIT('h0800)
	) name2346 (
		\ctl_rf_c5brbs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4575_
	);
	LUT4 #(
		.INIT('h0001)
	) name2347 (
		_w4572_,
		_w4573_,
		_w4574_,
		_w4575_,
		_w4576_
	);
	LUT3 #(
		.INIT('h2a)
	) name2348 (
		_w3425_,
		_w4571_,
		_w4576_,
		_w4577_
	);
	LUT4 #(
		.INIT('h0020)
	) name2349 (
		\ctl_rf_c2dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4578_
	);
	LUT4 #(
		.INIT('h0080)
	) name2350 (
		\ctl_rf_c3dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4579_
	);
	LUT4 #(
		.INIT('h0002)
	) name2351 (
		\ctl_rf_c0dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4580_
	);
	LUT4 #(
		.INIT('h2000)
	) name2352 (
		\ctl_rf_c6dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4581_
	);
	LUT4 #(
		.INIT('h0001)
	) name2353 (
		_w4578_,
		_w4579_,
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT4 #(
		.INIT('h8000)
	) name2354 (
		\ctl_rf_c7dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4583_
	);
	LUT4 #(
		.INIT('h0200)
	) name2355 (
		\ctl_rf_c4dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4584_
	);
	LUT4 #(
		.INIT('h0008)
	) name2356 (
		\ctl_rf_c1dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4585_
	);
	LUT4 #(
		.INIT('h0800)
	) name2357 (
		\ctl_rf_c5dmabs_reg[18]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4586_
	);
	LUT4 #(
		.INIT('h0001)
	) name2358 (
		_w4583_,
		_w4584_,
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT3 #(
		.INIT('h2a)
	) name2359 (
		_w3431_,
		_w4582_,
		_w4587_,
		_w4588_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2360 (
		\ctl_rf_abt_reg[2]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w4589_
	);
	LUT4 #(
		.INIT('h0023)
	) name2361 (
		\ctl_rf_c2_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w4590_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w4589_,
		_w4590_,
		_w4591_
	);
	LUT3 #(
		.INIT('h01)
	) name2363 (
		_w4577_,
		_w4588_,
		_w4591_,
		_w4592_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2364 (
		_w3422_,
		_w4577_,
		_w4588_,
		_w4591_,
		_w4593_
	);
	LUT4 #(
		.INIT('h4055)
	) name2365 (
		_w3622_,
		_w4550_,
		_w4566_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w4533_,
		_w4594_,
		_w4595_
	);
	LUT3 #(
		.INIT('h20)
	) name2367 (
		_w3503_,
		_w4042_,
		_w4053_,
		_w4596_
	);
	LUT3 #(
		.INIT('hc4)
	) name2368 (
		_w3427_,
		_w3503_,
		_w4075_,
		_w4597_
	);
	LUT3 #(
		.INIT('h13)
	) name2369 (
		_w4070_,
		_w4596_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h1311)
	) name2370 (
		_w3484_,
		_w3503_,
		_w4118_,
		_w4124_,
		_w4599_
	);
	LUT2 #(
		.INIT('h4)
	) name2371 (
		_w4117_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h1)
	) name2372 (
		_w3424_,
		_w4533_,
		_w4601_
	);
	LUT3 #(
		.INIT('hd0)
	) name2373 (
		_w4598_,
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w4595_,
		_w4602_,
		_w4603_
	);
	LUT3 #(
		.INIT('h2a)
	) name2375 (
		\hrdata_reg[30]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4604_
	);
	LUT3 #(
		.INIT('h02)
	) name2376 (
		\ctl_rf_c0_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4605_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2377 (
		\ctl_rf_c0_rf_chdad_reg[14]/NET0131 ,
		\ctl_rf_c0_rf_chsad_reg[14]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4606_
	);
	LUT3 #(
		.INIT('h8a)
	) name2378 (
		_w3445_,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('h02)
	) name2379 (
		\ctl_rf_c7_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4608_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2380 (
		\ctl_rf_c7_rf_chdad_reg[14]/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[14]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4609_
	);
	LUT3 #(
		.INIT('h8a)
	) name2381 (
		_w3453_,
		_w4608_,
		_w4609_,
		_w4610_
	);
	LUT3 #(
		.INIT('h02)
	) name2382 (
		\ctl_rf_c6_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4611_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2383 (
		\ctl_rf_c6_rf_chdad_reg[14]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[14]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4612_
	);
	LUT3 #(
		.INIT('h8a)
	) name2384 (
		_w3440_,
		_w4611_,
		_w4612_,
		_w4613_
	);
	LUT3 #(
		.INIT('h02)
	) name2385 (
		\ctl_rf_c1_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4614_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2386 (
		\ctl_rf_c1_rf_chdad_reg[14]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[14]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4615_
	);
	LUT3 #(
		.INIT('h8a)
	) name2387 (
		_w3449_,
		_w4614_,
		_w4615_,
		_w4616_
	);
	LUT4 #(
		.INIT('h0001)
	) name2388 (
		_w4607_,
		_w4610_,
		_w4613_,
		_w4616_,
		_w4617_
	);
	LUT3 #(
		.INIT('h02)
	) name2389 (
		\ctl_rf_c3_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4618_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2390 (
		\ctl_rf_c3_rf_chdad_reg[14]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[14]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4619_
	);
	LUT3 #(
		.INIT('h8a)
	) name2391 (
		_w3457_,
		_w4618_,
		_w4619_,
		_w4620_
	);
	LUT3 #(
		.INIT('h02)
	) name2392 (
		\ctl_rf_c2_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4621_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2393 (
		\ctl_rf_c2_rf_chdad_reg[14]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[14]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4622_
	);
	LUT3 #(
		.INIT('h8a)
	) name2394 (
		_w3432_,
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT3 #(
		.INIT('h02)
	) name2395 (
		\ctl_rf_c4_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4624_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2396 (
		\ctl_rf_c4_rf_chdad_reg[14]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[14]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4625_
	);
	LUT3 #(
		.INIT('h8a)
	) name2397 (
		_w3426_,
		_w4624_,
		_w4625_,
		_w4626_
	);
	LUT3 #(
		.INIT('h02)
	) name2398 (
		\ctl_rf_c5_rf_autold_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4627_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2399 (
		\ctl_rf_c5_rf_chdad_reg[14]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[14]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4628_
	);
	LUT3 #(
		.INIT('h8a)
	) name2400 (
		_w3436_,
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT4 #(
		.INIT('h0001)
	) name2401 (
		_w4620_,
		_w4623_,
		_w4626_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		_w4617_,
		_w4630_,
		_w4631_
	);
	LUT4 #(
		.INIT('h135f)
	) name2403 (
		\ctl_rf_c5_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[14]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4632_
	);
	LUT4 #(
		.INIT('h135f)
	) name2404 (
		\ctl_rf_c1_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[14]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4633_
	);
	LUT4 #(
		.INIT('h153f)
	) name2405 (
		\ctl_rf_c0_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[14]/NET0131 ,
		_w3464_,
		_w3467_,
		_w4634_
	);
	LUT4 #(
		.INIT('h135f)
	) name2406 (
		\ctl_rf_c2_rf_chllp_reg[14]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[14]/NET0131 ,
		_w3462_,
		_w3472_,
		_w4635_
	);
	LUT4 #(
		.INIT('h8000)
	) name2407 (
		_w4632_,
		_w4633_,
		_w4634_,
		_w4635_,
		_w4636_
	);
	LUT3 #(
		.INIT('ha2)
	) name2408 (
		_w3424_,
		_w3427_,
		_w4636_,
		_w4637_
	);
	LUT4 #(
		.INIT('h0222)
	) name2409 (
		_w3422_,
		_w3689_,
		_w4631_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h1)
	) name2410 (
		_w4604_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h0800)
	) name2411 (
		\ctl_rf_c5dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4640_
	);
	LUT4 #(
		.INIT('h2000)
	) name2412 (
		\ctl_rf_c6dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4641_
	);
	LUT4 #(
		.INIT('h0008)
	) name2413 (
		\ctl_rf_c1dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4642_
	);
	LUT4 #(
		.INIT('h0020)
	) name2414 (
		\ctl_rf_c2dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4643_
	);
	LUT4 #(
		.INIT('h0001)
	) name2415 (
		_w4640_,
		_w4641_,
		_w4642_,
		_w4643_,
		_w4644_
	);
	LUT4 #(
		.INIT('h0080)
	) name2416 (
		\ctl_rf_c3dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4645_
	);
	LUT4 #(
		.INIT('h0200)
	) name2417 (
		\ctl_rf_c4dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4646_
	);
	LUT4 #(
		.INIT('h0002)
	) name2418 (
		\ctl_rf_c0dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4647_
	);
	LUT4 #(
		.INIT('h8000)
	) name2419 (
		\ctl_rf_c7dmabs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4648_
	);
	LUT4 #(
		.INIT('h0001)
	) name2420 (
		_w4645_,
		_w4646_,
		_w4647_,
		_w4648_,
		_w4649_
	);
	LUT3 #(
		.INIT('h2a)
	) name2421 (
		_w3431_,
		_w4644_,
		_w4649_,
		_w4650_
	);
	LUT4 #(
		.INIT('h0008)
	) name2422 (
		\ctl_rf_c1brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4651_
	);
	LUT4 #(
		.INIT('h8000)
	) name2423 (
		\ctl_rf_c7brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4652_
	);
	LUT4 #(
		.INIT('h0200)
	) name2424 (
		\ctl_rf_c4brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4653_
	);
	LUT4 #(
		.INIT('h0800)
	) name2425 (
		\ctl_rf_c5brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4654_
	);
	LUT4 #(
		.INIT('h0001)
	) name2426 (
		_w4651_,
		_w4652_,
		_w4653_,
		_w4654_,
		_w4655_
	);
	LUT4 #(
		.INIT('h0020)
	) name2427 (
		\ctl_rf_c2brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4656_
	);
	LUT4 #(
		.INIT('h0002)
	) name2428 (
		\ctl_rf_c0brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4657_
	);
	LUT4 #(
		.INIT('h0080)
	) name2429 (
		\ctl_rf_c3brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4658_
	);
	LUT4 #(
		.INIT('h2000)
	) name2430 (
		\ctl_rf_c6brbs_reg[30]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4659_
	);
	LUT4 #(
		.INIT('h0001)
	) name2431 (
		_w4656_,
		_w4657_,
		_w4658_,
		_w4659_,
		_w4660_
	);
	LUT4 #(
		.INIT('h5111)
	) name2432 (
		\haddr[8]_pad ,
		_w3425_,
		_w4655_,
		_w4660_,
		_w4661_
	);
	LUT3 #(
		.INIT('h10)
	) name2433 (
		_w3503_,
		_w4650_,
		_w4661_,
		_w4662_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2434 (
		\ctl_rf_c6_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c6_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4663_
	);
	LUT2 #(
		.INIT('h2)
	) name2435 (
		_w3440_,
		_w4663_,
		_w4664_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2436 (
		\ctl_rf_c7_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c7_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4665_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2437 (
		\ctl_rf_c3_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c3_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4666_
	);
	LUT4 #(
		.INIT('hf531)
	) name2438 (
		_w3453_,
		_w3457_,
		_w4665_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		_w4664_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2440 (
		\ctl_rf_c1_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c1_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4669_
	);
	LUT3 #(
		.INIT('ha2)
	) name2441 (
		\haddr[8]_pad ,
		_w3449_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2442 (
		\ctl_rf_c4_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c4_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4671_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2443 (
		\ctl_rf_c2_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c2_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4672_
	);
	LUT4 #(
		.INIT('hf531)
	) name2444 (
		_w3426_,
		_w3432_,
		_w4671_,
		_w4672_,
		_w4673_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2445 (
		\ctl_rf_c0_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c0_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4674_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2446 (
		\ctl_rf_c5_rf_chdad_reg[30]/P0002 ,
		\ctl_rf_c5_rf_chsad_reg[30]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4675_
	);
	LUT4 #(
		.INIT('hf351)
	) name2447 (
		_w3436_,
		_w3445_,
		_w4674_,
		_w4675_,
		_w4676_
	);
	LUT3 #(
		.INIT('h80)
	) name2448 (
		_w4670_,
		_w4673_,
		_w4676_,
		_w4677_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w4668_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h135f)
	) name2450 (
		\ctl_rf_c1_rf_chllp_reg[30]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[30]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4679_
	);
	LUT4 #(
		.INIT('h135f)
	) name2451 (
		\ctl_rf_c0_rf_chllp_reg[30]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[30]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4680_
	);
	LUT4 #(
		.INIT('h135f)
	) name2452 (
		\ctl_rf_c5_rf_chllp_reg[30]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[30]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4681_
	);
	LUT4 #(
		.INIT('h135f)
	) name2453 (
		\ctl_rf_c2_rf_chllp_reg[30]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[30]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4682_
	);
	LUT4 #(
		.INIT('h8000)
	) name2454 (
		_w4679_,
		_w4680_,
		_w4681_,
		_w4682_,
		_w4683_
	);
	LUT3 #(
		.INIT('h31)
	) name2455 (
		_w3427_,
		_w3503_,
		_w4683_,
		_w4684_
	);
	LUT3 #(
		.INIT('h15)
	) name2456 (
		_w4662_,
		_w4678_,
		_w4684_,
		_w4685_
	);
	LUT3 #(
		.INIT('h20)
	) name2457 (
		\ctl_rf_c5_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4686_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2458 (
		\ctl_rf_c5_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c5_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4687_
	);
	LUT3 #(
		.INIT('h8a)
	) name2459 (
		_w3436_,
		_w4686_,
		_w4687_,
		_w4688_
	);
	LUT3 #(
		.INIT('h20)
	) name2460 (
		\ctl_rf_c2_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4689_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2461 (
		\ctl_rf_c2_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c2_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4690_
	);
	LUT3 #(
		.INIT('h8a)
	) name2462 (
		_w3432_,
		_w4689_,
		_w4690_,
		_w4691_
	);
	LUT3 #(
		.INIT('h20)
	) name2463 (
		\ctl_rf_c0_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4692_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2464 (
		\ctl_rf_c0_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c0_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4693_
	);
	LUT3 #(
		.INIT('h8a)
	) name2465 (
		_w3445_,
		_w4692_,
		_w4693_,
		_w4694_
	);
	LUT3 #(
		.INIT('h20)
	) name2466 (
		\ctl_rf_c3_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4695_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2467 (
		\ctl_rf_c3_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c3_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4696_
	);
	LUT3 #(
		.INIT('h8a)
	) name2468 (
		_w3457_,
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT4 #(
		.INIT('h0001)
	) name2469 (
		_w4688_,
		_w4691_,
		_w4694_,
		_w4697_,
		_w4698_
	);
	LUT3 #(
		.INIT('h20)
	) name2470 (
		\ctl_rf_c7_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4699_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2471 (
		\ctl_rf_c7_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c7_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4700_
	);
	LUT3 #(
		.INIT('h8a)
	) name2472 (
		_w3453_,
		_w4699_,
		_w4700_,
		_w4701_
	);
	LUT3 #(
		.INIT('h20)
	) name2473 (
		\ctl_rf_c4_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4702_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2474 (
		\ctl_rf_c4_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c4_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4703_
	);
	LUT3 #(
		.INIT('h8a)
	) name2475 (
		_w3426_,
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT3 #(
		.INIT('h20)
	) name2476 (
		\ctl_rf_c1_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4705_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2477 (
		\ctl_rf_c1_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c1_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4706_
	);
	LUT3 #(
		.INIT('h8a)
	) name2478 (
		_w3449_,
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT3 #(
		.INIT('h20)
	) name2479 (
		\ctl_rf_c6_rf_chsad_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4708_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2480 (
		\ctl_rf_c6_rf_chdad_reg[6]/P0002 ,
		\ctl_rf_c6_rf_sad_ctl1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4709_
	);
	LUT3 #(
		.INIT('h8a)
	) name2481 (
		_w3440_,
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT4 #(
		.INIT('h0001)
	) name2482 (
		_w4701_,
		_w4704_,
		_w4707_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('hff35)
	) name2483 (
		\ctl_rf_c2_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4712_
	);
	LUT4 #(
		.INIT('hff35)
	) name2484 (
		\ctl_rf_c3_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4713_
	);
	LUT4 #(
		.INIT('hf531)
	) name2485 (
		_w3462_,
		_w3477_,
		_w4712_,
		_w4713_,
		_w4714_
	);
	LUT4 #(
		.INIT('hff35)
	) name2486 (
		\ctl_rf_c7_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4715_
	);
	LUT4 #(
		.INIT('hff35)
	) name2487 (
		\ctl_rf_c4_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4716_
	);
	LUT4 #(
		.INIT('hf531)
	) name2488 (
		_w3464_,
		_w3472_,
		_w4715_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('hff35)
	) name2489 (
		\ctl_rf_c6_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4718_
	);
	LUT4 #(
		.INIT('hff35)
	) name2490 (
		\ctl_rf_c5_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4719_
	);
	LUT4 #(
		.INIT('hf351)
	) name2491 (
		_w3469_,
		_w3479_,
		_w4718_,
		_w4719_,
		_w4720_
	);
	LUT4 #(
		.INIT('hff35)
	) name2492 (
		\ctl_rf_c0_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4721_
	);
	LUT4 #(
		.INIT('hff35)
	) name2493 (
		\ctl_rf_c1_rf_chllp_reg[6]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4722_
	);
	LUT4 #(
		.INIT('hf531)
	) name2494 (
		_w3467_,
		_w3474_,
		_w4721_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h8000)
	) name2495 (
		_w4714_,
		_w4717_,
		_w4720_,
		_w4723_,
		_w4724_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2496 (
		\haddr[8]_pad ,
		_w4698_,
		_w4711_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		_w2527_,
		_w3486_,
		_w4726_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name2498 (
		\ctl_rf_c6_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[6]/NET0131 ,
		_w3488_,
		_w3489_,
		_w4727_
	);
	LUT2 #(
		.INIT('h2)
	) name2499 (
		\ctl_rf_abt_reg[6]/NET0131 ,
		\ctl_rf_c6_rf_int_abt_msk_reg/NET0131 ,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		_w3496_,
		_w4728_,
		_w4729_
	);
	LUT4 #(
		.INIT('h153f)
	) name2501 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[6]/NET0131 ,
		_w3491_,
		_w3492_,
		_w4730_
	);
	LUT3 #(
		.INIT('h20)
	) name2502 (
		_w4727_,
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2503 (
		_w3484_,
		_w3503_,
		_w4726_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h4)
	) name2504 (
		_w4725_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w3424_,
		_w4604_,
		_w4734_
	);
	LUT3 #(
		.INIT('hd0)
	) name2506 (
		_w4685_,
		_w4733_,
		_w4734_,
		_w4735_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w4639_,
		_w4735_,
		_w4736_
	);
	LUT3 #(
		.INIT('h2a)
	) name2508 (
		\hrdata_reg[31]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4737_
	);
	LUT3 #(
		.INIT('h80)
	) name2509 (
		\ctl_rf_c0_rf_chdad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4738_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2510 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_c0_rf_chsad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4739_
	);
	LUT3 #(
		.INIT('h8a)
	) name2511 (
		_w3445_,
		_w4738_,
		_w4739_,
		_w4740_
	);
	LUT3 #(
		.INIT('h20)
	) name2512 (
		\ctl_rf_c6_rf_chsad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4741_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name2513 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_c6_rf_chdad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4742_
	);
	LUT3 #(
		.INIT('h8a)
	) name2514 (
		_w3440_,
		_w4741_,
		_w4742_,
		_w4743_
	);
	LUT3 #(
		.INIT('h80)
	) name2515 (
		\ctl_rf_c7_rf_chdad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4744_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2516 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4745_
	);
	LUT3 #(
		.INIT('h8a)
	) name2517 (
		_w3453_,
		_w4744_,
		_w4745_,
		_w4746_
	);
	LUT3 #(
		.INIT('h80)
	) name2518 (
		\ctl_rf_c1_rf_chdad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4747_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2519 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4748_
	);
	LUT3 #(
		.INIT('h8a)
	) name2520 (
		_w3449_,
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT4 #(
		.INIT('h0001)
	) name2521 (
		_w4740_,
		_w4743_,
		_w4746_,
		_w4749_,
		_w4750_
	);
	LUT3 #(
		.INIT('h80)
	) name2522 (
		\ctl_rf_c3_rf_chdad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4751_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2523 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\ctl_rf_c3_rf_chsad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4752_
	);
	LUT3 #(
		.INIT('h8a)
	) name2524 (
		_w3457_,
		_w4751_,
		_w4752_,
		_w4753_
	);
	LUT3 #(
		.INIT('h20)
	) name2525 (
		\ctl_rf_c2_rf_chsad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4754_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name2526 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_c2_rf_chdad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4755_
	);
	LUT3 #(
		.INIT('h8a)
	) name2527 (
		_w3432_,
		_w4754_,
		_w4755_,
		_w4756_
	);
	LUT3 #(
		.INIT('h20)
	) name2528 (
		\ctl_rf_c4_rf_chsad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4757_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name2529 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_c4_rf_chdad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4758_
	);
	LUT3 #(
		.INIT('h8a)
	) name2530 (
		_w3426_,
		_w4757_,
		_w4758_,
		_w4759_
	);
	LUT3 #(
		.INIT('h20)
	) name2531 (
		\ctl_rf_c5_rf_chsad_reg[15]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4760_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name2532 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_c5_rf_chdad_reg[15]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4761_
	);
	LUT3 #(
		.INIT('h8a)
	) name2533 (
		_w3436_,
		_w4760_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('h0001)
	) name2534 (
		_w4753_,
		_w4756_,
		_w4759_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		_w4750_,
		_w4763_,
		_w4764_
	);
	LUT4 #(
		.INIT('h135f)
	) name2536 (
		\ctl_rf_c5_rf_chllp_reg[15]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[15]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4765_
	);
	LUT4 #(
		.INIT('h135f)
	) name2537 (
		\ctl_rf_c0_rf_chllp_reg[15]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[15]/NET0131 ,
		_w3467_,
		_w3477_,
		_w4766_
	);
	LUT4 #(
		.INIT('h153f)
	) name2538 (
		\ctl_rf_c1_rf_chllp_reg[15]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[15]/NET0131 ,
		_w3464_,
		_w3474_,
		_w4767_
	);
	LUT4 #(
		.INIT('h135f)
	) name2539 (
		\ctl_rf_c2_rf_chllp_reg[15]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[15]/NET0131 ,
		_w3462_,
		_w3472_,
		_w4768_
	);
	LUT4 #(
		.INIT('h8000)
	) name2540 (
		_w4765_,
		_w4766_,
		_w4767_,
		_w4768_,
		_w4769_
	);
	LUT3 #(
		.INIT('ha2)
	) name2541 (
		_w3424_,
		_w3427_,
		_w4769_,
		_w4770_
	);
	LUT4 #(
		.INIT('h0222)
	) name2542 (
		_w3422_,
		_w3689_,
		_w4764_,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name2543 (
		_w4737_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2544 (
		\ctl_rf_c1_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c1_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4773_
	);
	LUT3 #(
		.INIT('h20)
	) name2545 (
		\ctl_rf_c1_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4774_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name2546 (
		\haddr[8]_pad ,
		_w3449_,
		_w4773_,
		_w4774_,
		_w4775_
	);
	LUT3 #(
		.INIT('h20)
	) name2547 (
		\ctl_rf_c7_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4776_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2548 (
		\ctl_rf_c7_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c7_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4777_
	);
	LUT3 #(
		.INIT('h8a)
	) name2549 (
		_w3453_,
		_w4776_,
		_w4777_,
		_w4778_
	);
	LUT3 #(
		.INIT('h80)
	) name2550 (
		\ctl_rf_c0_rf_chdad_reg[31]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4779_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2551 (
		\ctl_rf_c0_rf_chsad_reg[31]/NET0131 ,
		\ctl_rf_c0_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4780_
	);
	LUT3 #(
		.INIT('h8a)
	) name2552 (
		_w3445_,
		_w4779_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('h20)
	) name2553 (
		\ctl_rf_c5_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4782_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2554 (
		\ctl_rf_c5_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c5_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4783_
	);
	LUT3 #(
		.INIT('h8a)
	) name2555 (
		_w3436_,
		_w4782_,
		_w4783_,
		_w4784_
	);
	LUT3 #(
		.INIT('h20)
	) name2556 (
		\ctl_rf_c2_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4785_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2557 (
		\ctl_rf_c2_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c2_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4786_
	);
	LUT3 #(
		.INIT('h8a)
	) name2558 (
		_w3432_,
		_w4785_,
		_w4786_,
		_w4787_
	);
	LUT4 #(
		.INIT('h0001)
	) name2559 (
		_w4778_,
		_w4781_,
		_w4784_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w4775_,
		_w4788_,
		_w4789_
	);
	LUT4 #(
		.INIT('h135f)
	) name2561 (
		\ctl_rf_c0_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[31]/NET0131 ,
		_w3467_,
		_w3469_,
		_w4790_
	);
	LUT4 #(
		.INIT('h135f)
	) name2562 (
		\ctl_rf_c2_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[31]/NET0131 ,
		_w3462_,
		_w3479_,
		_w4791_
	);
	LUT4 #(
		.INIT('h135f)
	) name2563 (
		\ctl_rf_c1_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[31]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4792_
	);
	LUT4 #(
		.INIT('h153f)
	) name2564 (
		\ctl_rf_c4_rf_chllp_reg[31]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[31]/NET0131 ,
		_w3464_,
		_w3472_,
		_w4793_
	);
	LUT4 #(
		.INIT('h8000)
	) name2565 (
		_w4790_,
		_w4791_,
		_w4792_,
		_w4793_,
		_w4794_
	);
	LUT3 #(
		.INIT('h80)
	) name2566 (
		\ctl_rf_c3_rf_chdad_reg[31]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4795_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2567 (
		\ctl_rf_c3_rf_chsad_reg[31]/NET0131 ,
		\ctl_rf_c3_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4796_
	);
	LUT3 #(
		.INIT('h8a)
	) name2568 (
		_w3457_,
		_w4795_,
		_w4796_,
		_w4797_
	);
	LUT3 #(
		.INIT('h20)
	) name2569 (
		\ctl_rf_c4_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4798_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2570 (
		\ctl_rf_c4_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c4_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4799_
	);
	LUT3 #(
		.INIT('h8a)
	) name2571 (
		_w3426_,
		_w4798_,
		_w4799_,
		_w4800_
	);
	LUT3 #(
		.INIT('h20)
	) name2572 (
		\ctl_rf_c6_rf_chsad_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4801_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2573 (
		\ctl_rf_c6_rf_chdad_reg[31]/P0002 ,
		\ctl_rf_c6_rf_int_tc_msk_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4802_
	);
	LUT3 #(
		.INIT('h8a)
	) name2574 (
		_w3440_,
		_w4801_,
		_w4802_,
		_w4803_
	);
	LUT3 #(
		.INIT('h01)
	) name2575 (
		_w4797_,
		_w4800_,
		_w4803_,
		_w4804_
	);
	LUT3 #(
		.INIT('hd0)
	) name2576 (
		_w3427_,
		_w4794_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('h0800)
	) name2577 (
		\ctl_rf_c5brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4806_
	);
	LUT4 #(
		.INIT('h2000)
	) name2578 (
		\ctl_rf_c6brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4807_
	);
	LUT4 #(
		.INIT('h0008)
	) name2579 (
		\ctl_rf_c1brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4808_
	);
	LUT4 #(
		.INIT('h0020)
	) name2580 (
		\ctl_rf_c2brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4809_
	);
	LUT4 #(
		.INIT('h0001)
	) name2581 (
		_w4806_,
		_w4807_,
		_w4808_,
		_w4809_,
		_w4810_
	);
	LUT4 #(
		.INIT('h0080)
	) name2582 (
		\ctl_rf_c3brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4811_
	);
	LUT4 #(
		.INIT('h0200)
	) name2583 (
		\ctl_rf_c4brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4812_
	);
	LUT4 #(
		.INIT('h0002)
	) name2584 (
		\ctl_rf_c0brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4813_
	);
	LUT4 #(
		.INIT('h8000)
	) name2585 (
		\ctl_rf_c7brbs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4814_
	);
	LUT4 #(
		.INIT('h0001)
	) name2586 (
		_w4811_,
		_w4812_,
		_w4813_,
		_w4814_,
		_w4815_
	);
	LUT3 #(
		.INIT('h2a)
	) name2587 (
		_w3425_,
		_w4810_,
		_w4815_,
		_w4816_
	);
	LUT4 #(
		.INIT('h0008)
	) name2588 (
		\ctl_rf_c1dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4817_
	);
	LUT4 #(
		.INIT('h2000)
	) name2589 (
		\ctl_rf_c6dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4818_
	);
	LUT4 #(
		.INIT('h0200)
	) name2590 (
		\ctl_rf_c4dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4819_
	);
	LUT4 #(
		.INIT('h0080)
	) name2591 (
		\ctl_rf_c3dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4820_
	);
	LUT4 #(
		.INIT('h0001)
	) name2592 (
		_w4817_,
		_w4818_,
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT4 #(
		.INIT('h0020)
	) name2593 (
		\ctl_rf_c2dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4822_
	);
	LUT4 #(
		.INIT('h0002)
	) name2594 (
		\ctl_rf_c0dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4823_
	);
	LUT4 #(
		.INIT('h0800)
	) name2595 (
		\ctl_rf_c5dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4824_
	);
	LUT4 #(
		.INIT('h8000)
	) name2596 (
		\ctl_rf_c7dmabs_reg[31]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4825_
	);
	LUT4 #(
		.INIT('h0001)
	) name2597 (
		_w4822_,
		_w4823_,
		_w4824_,
		_w4825_,
		_w4826_
	);
	LUT4 #(
		.INIT('h5111)
	) name2598 (
		\haddr[8]_pad ,
		_w3431_,
		_w4821_,
		_w4826_,
		_w4827_
	);
	LUT2 #(
		.INIT('h4)
	) name2599 (
		_w4816_,
		_w4827_,
		_w4828_
	);
	LUT4 #(
		.INIT('h5540)
	) name2600 (
		_w3503_,
		_w4789_,
		_w4805_,
		_w4828_,
		_w4829_
	);
	LUT3 #(
		.INIT('h20)
	) name2601 (
		\ctl_rf_c4_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4830_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2602 (
		\ctl_rf_c4_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c4_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4831_
	);
	LUT3 #(
		.INIT('h8a)
	) name2603 (
		_w3426_,
		_w4830_,
		_w4831_,
		_w4832_
	);
	LUT3 #(
		.INIT('h20)
	) name2604 (
		\ctl_rf_c6_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4833_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2605 (
		\ctl_rf_c6_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c6_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4834_
	);
	LUT3 #(
		.INIT('h8a)
	) name2606 (
		_w3440_,
		_w4833_,
		_w4834_,
		_w4835_
	);
	LUT3 #(
		.INIT('h20)
	) name2607 (
		\ctl_rf_c7_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4836_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2608 (
		\ctl_rf_c7_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c7_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4837_
	);
	LUT3 #(
		.INIT('h8a)
	) name2609 (
		_w3453_,
		_w4836_,
		_w4837_,
		_w4838_
	);
	LUT3 #(
		.INIT('h20)
	) name2610 (
		\ctl_rf_c1_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4839_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2611 (
		\ctl_rf_c1_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c1_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4840_
	);
	LUT3 #(
		.INIT('h8a)
	) name2612 (
		_w3449_,
		_w4839_,
		_w4840_,
		_w4841_
	);
	LUT4 #(
		.INIT('h0001)
	) name2613 (
		_w4832_,
		_w4835_,
		_w4838_,
		_w4841_,
		_w4842_
	);
	LUT3 #(
		.INIT('h20)
	) name2614 (
		\ctl_rf_c0_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4843_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2615 (
		\ctl_rf_c0_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c0_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4844_
	);
	LUT3 #(
		.INIT('h8a)
	) name2616 (
		_w3445_,
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT3 #(
		.INIT('h20)
	) name2617 (
		\ctl_rf_c5_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4846_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2618 (
		\ctl_rf_c5_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c5_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4847_
	);
	LUT3 #(
		.INIT('h8a)
	) name2619 (
		_w3436_,
		_w4846_,
		_w4847_,
		_w4848_
	);
	LUT3 #(
		.INIT('h20)
	) name2620 (
		\ctl_rf_c3_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4849_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2621 (
		\ctl_rf_c3_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c3_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4850_
	);
	LUT3 #(
		.INIT('h8a)
	) name2622 (
		_w3457_,
		_w4849_,
		_w4850_,
		_w4851_
	);
	LUT3 #(
		.INIT('h20)
	) name2623 (
		\ctl_rf_c2_rf_chsad_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4852_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2624 (
		\ctl_rf_c2_rf_chdad_reg[7]/P0002 ,
		\ctl_rf_c2_rf_mode_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4853_
	);
	LUT3 #(
		.INIT('h8a)
	) name2625 (
		_w3432_,
		_w4852_,
		_w4853_,
		_w4854_
	);
	LUT4 #(
		.INIT('h0001)
	) name2626 (
		_w4845_,
		_w4848_,
		_w4851_,
		_w4854_,
		_w4855_
	);
	LUT4 #(
		.INIT('hff35)
	) name2627 (
		\ctl_rf_c3_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c3_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4856_
	);
	LUT4 #(
		.INIT('hff35)
	) name2628 (
		\ctl_rf_c0_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c0_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4857_
	);
	LUT4 #(
		.INIT('hf351)
	) name2629 (
		_w3467_,
		_w3477_,
		_w4856_,
		_w4857_,
		_w4858_
	);
	LUT4 #(
		.INIT('hff35)
	) name2630 (
		\ctl_rf_c5_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c5_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4859_
	);
	LUT4 #(
		.INIT('hff35)
	) name2631 (
		\ctl_rf_c1_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c1_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4860_
	);
	LUT4 #(
		.INIT('hf531)
	) name2632 (
		_w3469_,
		_w3474_,
		_w4859_,
		_w4860_,
		_w4861_
	);
	LUT4 #(
		.INIT('hff35)
	) name2633 (
		\ctl_rf_c2_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c2_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4862_
	);
	LUT4 #(
		.INIT('hff35)
	) name2634 (
		\ctl_rf_c7_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c7_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4863_
	);
	LUT4 #(
		.INIT('hf531)
	) name2635 (
		_w3462_,
		_w3464_,
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT4 #(
		.INIT('hff35)
	) name2636 (
		\ctl_rf_c4_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c4_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4865_
	);
	LUT4 #(
		.INIT('hff35)
	) name2637 (
		\ctl_rf_c6_rf_chllp_reg[7]/NET0131 ,
		\ctl_rf_c6_rf_chtsz_reg[7]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4866_
	);
	LUT4 #(
		.INIT('hf531)
	) name2638 (
		_w3472_,
		_w3479_,
		_w4865_,
		_w4866_,
		_w4867_
	);
	LUT4 #(
		.INIT('h8000)
	) name2639 (
		_w4858_,
		_w4861_,
		_w4864_,
		_w4867_,
		_w4868_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2640 (
		\haddr[8]_pad ,
		_w4842_,
		_w4855_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		_w2527_,
		_w3927_,
		_w4870_
	);
	LUT4 #(
		.INIT('h3b3f)
	) name2642 (
		\ctl_rf_c7_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[7]/NET0131 ,
		_w3488_,
		_w3489_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		\ctl_rf_abt_reg[7]/NET0131 ,
		\ctl_rf_c7_rf_int_abt_msk_reg/NET0131 ,
		_w4872_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		_w3496_,
		_w4872_,
		_w4873_
	);
	LUT4 #(
		.INIT('h153f)
	) name2645 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_sync_reg[7]/NET0131 ,
		_w3491_,
		_w3492_,
		_w4874_
	);
	LUT3 #(
		.INIT('h20)
	) name2646 (
		_w4871_,
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2647 (
		_w3484_,
		_w3503_,
		_w4870_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w4869_,
		_w4876_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w3424_,
		_w4737_,
		_w4878_
	);
	LUT3 #(
		.INIT('he0)
	) name2650 (
		_w4829_,
		_w4877_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h1)
	) name2651 (
		_w4772_,
		_w4879_,
		_w4880_
	);
	LUT3 #(
		.INIT('h2a)
	) name2652 (
		\hrdata_reg[3]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4881_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2653 (
		\ctl_rf_c0_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4882_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2654 (
		\ctl_rf_c0_rf_chsad_reg[19]/NET0131 ,
		\ctl_rf_c0_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4883_
	);
	LUT4 #(
		.INIT('ha222)
	) name2655 (
		\haddr[8]_pad ,
		_w3445_,
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('hf35f)
	) name2656 (
		\ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131 ,
		\ctl_rf_c2_rf_chsad_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4885_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2657 (
		\ctl_rf_c2_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c2_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4886_
	);
	LUT3 #(
		.INIT('h2a)
	) name2658 (
		_w3432_,
		_w4885_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2659 (
		\ctl_rf_c4_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4888_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2660 (
		\ctl_rf_c4_rf_chsad_reg[19]/NET0131 ,
		\ctl_rf_c4_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4889_
	);
	LUT3 #(
		.INIT('h2a)
	) name2661 (
		_w3426_,
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT4 #(
		.INIT('hff53)
	) name2662 (
		\ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131 ,
		\ctl_rf_c7_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4891_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2663 (
		\ctl_rf_c7_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c7_rf_chsad_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4892_
	);
	LUT3 #(
		.INIT('h2a)
	) name2664 (
		_w3453_,
		_w4891_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('hff53)
	) name2665 (
		\ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131 ,
		\ctl_rf_c1_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4894_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2666 (
		\ctl_rf_c1_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c1_rf_chsad_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4895_
	);
	LUT3 #(
		.INIT('h2a)
	) name2667 (
		_w3449_,
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT4 #(
		.INIT('h0001)
	) name2668 (
		_w4887_,
		_w4890_,
		_w4893_,
		_w4896_,
		_w4897_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		_w4884_,
		_w4897_,
		_w4898_
	);
	LUT4 #(
		.INIT('h135f)
	) name2670 (
		\ctl_rf_c1_rf_chllp_reg[19]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[19]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4899_
	);
	LUT4 #(
		.INIT('h135f)
	) name2671 (
		\ctl_rf_c0_rf_chllp_reg[19]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[19]/NET0131 ,
		_w3467_,
		_w3472_,
		_w4900_
	);
	LUT4 #(
		.INIT('h135f)
	) name2672 (
		\ctl_rf_c5_rf_chllp_reg[19]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[19]/NET0131 ,
		_w3469_,
		_w3479_,
		_w4901_
	);
	LUT4 #(
		.INIT('h135f)
	) name2673 (
		\ctl_rf_c2_rf_chllp_reg[19]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[19]/NET0131 ,
		_w3462_,
		_w3464_,
		_w4902_
	);
	LUT4 #(
		.INIT('h8000)
	) name2674 (
		_w4899_,
		_w4900_,
		_w4901_,
		_w4902_,
		_w4903_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2675 (
		\ctl_rf_c6_rf_chsad_reg[19]/NET0131 ,
		\ctl_rf_c6_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4904_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2676 (
		\ctl_rf_c6_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4905_
	);
	LUT3 #(
		.INIT('h2a)
	) name2677 (
		_w3440_,
		_w4904_,
		_w4905_,
		_w4906_
	);
	LUT4 #(
		.INIT('hff53)
	) name2678 (
		\ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131 ,
		\ctl_rf_c5_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4907_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2679 (
		\ctl_rf_c5_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4908_
	);
	LUT3 #(
		.INIT('h2a)
	) name2680 (
		_w3436_,
		_w4907_,
		_w4908_,
		_w4909_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name2681 (
		\ctl_rf_c3_rf_chdad_reg[19]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4910_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2682 (
		\ctl_rf_c3_rf_chsad_reg[19]/NET0131 ,
		\ctl_rf_c3_rf_prot1_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4911_
	);
	LUT3 #(
		.INIT('h2a)
	) name2683 (
		_w3457_,
		_w4910_,
		_w4911_,
		_w4912_
	);
	LUT3 #(
		.INIT('h01)
	) name2684 (
		_w4906_,
		_w4909_,
		_w4912_,
		_w4913_
	);
	LUT3 #(
		.INIT('hd0)
	) name2685 (
		_w3427_,
		_w4903_,
		_w4913_,
		_w4914_
	);
	LUT4 #(
		.INIT('h0008)
	) name2686 (
		\ctl_rf_c1dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4915_
	);
	LUT4 #(
		.INIT('h0080)
	) name2687 (
		\ctl_rf_c3dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4916_
	);
	LUT4 #(
		.INIT('h0002)
	) name2688 (
		\ctl_rf_c0dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4917_
	);
	LUT4 #(
		.INIT('h8000)
	) name2689 (
		\ctl_rf_c7dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4918_
	);
	LUT4 #(
		.INIT('h0001)
	) name2690 (
		_w4915_,
		_w4916_,
		_w4917_,
		_w4918_,
		_w4919_
	);
	LUT4 #(
		.INIT('h2000)
	) name2691 (
		\ctl_rf_c6dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4920_
	);
	LUT4 #(
		.INIT('h0200)
	) name2692 (
		\ctl_rf_c4dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4921_
	);
	LUT4 #(
		.INIT('h0020)
	) name2693 (
		\ctl_rf_c2dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4922_
	);
	LUT4 #(
		.INIT('h0800)
	) name2694 (
		\ctl_rf_c5dmabs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4923_
	);
	LUT4 #(
		.INIT('h0001)
	) name2695 (
		_w4920_,
		_w4921_,
		_w4922_,
		_w4923_,
		_w4924_
	);
	LUT3 #(
		.INIT('h2a)
	) name2696 (
		_w3431_,
		_w4919_,
		_w4924_,
		_w4925_
	);
	LUT4 #(
		.INIT('h0020)
	) name2697 (
		\ctl_rf_c2brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4926_
	);
	LUT4 #(
		.INIT('h0080)
	) name2698 (
		\ctl_rf_c3brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4927_
	);
	LUT4 #(
		.INIT('h0002)
	) name2699 (
		\ctl_rf_c0brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4928_
	);
	LUT4 #(
		.INIT('h2000)
	) name2700 (
		\ctl_rf_c6brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4929_
	);
	LUT4 #(
		.INIT('h0001)
	) name2701 (
		_w4926_,
		_w4927_,
		_w4928_,
		_w4929_,
		_w4930_
	);
	LUT4 #(
		.INIT('h8000)
	) name2702 (
		\ctl_rf_c7brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4931_
	);
	LUT4 #(
		.INIT('h0200)
	) name2703 (
		\ctl_rf_c4brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4932_
	);
	LUT4 #(
		.INIT('h0008)
	) name2704 (
		\ctl_rf_c1brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4933_
	);
	LUT4 #(
		.INIT('h0800)
	) name2705 (
		\ctl_rf_c5brbs_reg[19]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4934_
	);
	LUT4 #(
		.INIT('h0001)
	) name2706 (
		_w4931_,
		_w4932_,
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('h2a)
	) name2707 (
		_w3425_,
		_w4930_,
		_w4935_,
		_w4936_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2708 (
		\ctl_rf_abt_reg[3]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w4937_
	);
	LUT4 #(
		.INIT('h0023)
	) name2709 (
		\ctl_rf_c3_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w4938_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w4937_,
		_w4938_,
		_w4939_
	);
	LUT3 #(
		.INIT('h01)
	) name2711 (
		_w4925_,
		_w4936_,
		_w4939_,
		_w4940_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2712 (
		_w3422_,
		_w4925_,
		_w4936_,
		_w4939_,
		_w4941_
	);
	LUT4 #(
		.INIT('h4055)
	) name2713 (
		_w3622_,
		_w4898_,
		_w4914_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w4881_,
		_w4942_,
		_w4943_
	);
	LUT3 #(
		.INIT('h20)
	) name2715 (
		_w3503_,
		_w4181_,
		_w4192_,
		_w4944_
	);
	LUT3 #(
		.INIT('hc4)
	) name2716 (
		_w3427_,
		_w3503_,
		_w4214_,
		_w4945_
	);
	LUT3 #(
		.INIT('h13)
	) name2717 (
		_w4209_,
		_w4944_,
		_w4945_,
		_w4946_
	);
	LUT4 #(
		.INIT('h1311)
	) name2718 (
		_w3484_,
		_w3503_,
		_w4257_,
		_w4262_,
		_w4947_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w4256_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w3424_,
		_w4881_,
		_w4949_
	);
	LUT3 #(
		.INIT('hd0)
	) name2721 (
		_w4946_,
		_w4948_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w4943_,
		_w4950_,
		_w4951_
	);
	LUT3 #(
		.INIT('h2a)
	) name2723 (
		\hrdata_reg[4]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w4952_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2724 (
		\ctl_rf_c4_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c4_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4953_
	);
	LUT3 #(
		.INIT('h20)
	) name2725 (
		\ctl_rf_c4_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4954_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name2726 (
		\haddr[8]_pad ,
		_w3426_,
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT3 #(
		.INIT('h20)
	) name2727 (
		\ctl_rf_c6_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4956_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2728 (
		\ctl_rf_c6_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c6_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4957_
	);
	LUT3 #(
		.INIT('h8a)
	) name2729 (
		_w3440_,
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT3 #(
		.INIT('h80)
	) name2730 (
		\ctl_rf_c7_rf_chdad_reg[20]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4959_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2731 (
		\ctl_rf_c7_rf_chsad_reg[20]/NET0131 ,
		\ctl_rf_c7_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4960_
	);
	LUT3 #(
		.INIT('h8a)
	) name2732 (
		_w3453_,
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT3 #(
		.INIT('h20)
	) name2733 (
		\ctl_rf_c5_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4962_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2734 (
		\ctl_rf_c5_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c5_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4963_
	);
	LUT3 #(
		.INIT('h8a)
	) name2735 (
		_w3436_,
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT3 #(
		.INIT('h20)
	) name2736 (
		\ctl_rf_c2_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4965_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2737 (
		\ctl_rf_c2_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c2_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4966_
	);
	LUT3 #(
		.INIT('h8a)
	) name2738 (
		_w3432_,
		_w4965_,
		_w4966_,
		_w4967_
	);
	LUT4 #(
		.INIT('h0001)
	) name2739 (
		_w4958_,
		_w4961_,
		_w4964_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		_w4955_,
		_w4968_,
		_w4969_
	);
	LUT4 #(
		.INIT('h135f)
	) name2741 (
		\ctl_rf_c1_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[20]/NET0131 ,
		_w3474_,
		_w3477_,
		_w4970_
	);
	LUT4 #(
		.INIT('h135f)
	) name2742 (
		\ctl_rf_c0_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[20]/NET0131 ,
		_w3467_,
		_w3479_,
		_w4971_
	);
	LUT4 #(
		.INIT('h135f)
	) name2743 (
		\ctl_rf_c2_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[20]/NET0131 ,
		_w3462_,
		_w3472_,
		_w4972_
	);
	LUT4 #(
		.INIT('h153f)
	) name2744 (
		\ctl_rf_c5_rf_chllp_reg[20]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[20]/NET0131 ,
		_w3464_,
		_w3469_,
		_w4973_
	);
	LUT4 #(
		.INIT('h8000)
	) name2745 (
		_w4970_,
		_w4971_,
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT3 #(
		.INIT('h80)
	) name2746 (
		\ctl_rf_c0_rf_chdad_reg[20]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4975_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2747 (
		\ctl_rf_c0_rf_chsad_reg[20]/NET0131 ,
		\ctl_rf_c0_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4976_
	);
	LUT3 #(
		.INIT('h8a)
	) name2748 (
		_w3445_,
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT3 #(
		.INIT('h20)
	) name2749 (
		\ctl_rf_c3_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4978_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2750 (
		\ctl_rf_c3_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c3_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4979_
	);
	LUT3 #(
		.INIT('h8a)
	) name2751 (
		_w3457_,
		_w4978_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('h20)
	) name2752 (
		\ctl_rf_c1_rf_chsad_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4981_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2753 (
		\ctl_rf_c1_rf_chdad_reg[20]/P0002 ,
		\ctl_rf_c1_rf_prot2_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w4982_
	);
	LUT3 #(
		.INIT('h8a)
	) name2754 (
		_w3449_,
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('h01)
	) name2755 (
		_w4977_,
		_w4980_,
		_w4983_,
		_w4984_
	);
	LUT3 #(
		.INIT('hd0)
	) name2756 (
		_w3427_,
		_w4974_,
		_w4984_,
		_w4985_
	);
	LUT4 #(
		.INIT('h0008)
	) name2757 (
		\ctl_rf_c1dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4986_
	);
	LUT4 #(
		.INIT('h0080)
	) name2758 (
		\ctl_rf_c3dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4987_
	);
	LUT4 #(
		.INIT('h0002)
	) name2759 (
		\ctl_rf_c0dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4988_
	);
	LUT4 #(
		.INIT('h8000)
	) name2760 (
		\ctl_rf_c7dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4989_
	);
	LUT4 #(
		.INIT('h0001)
	) name2761 (
		_w4986_,
		_w4987_,
		_w4988_,
		_w4989_,
		_w4990_
	);
	LUT4 #(
		.INIT('h2000)
	) name2762 (
		\ctl_rf_c6dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4991_
	);
	LUT4 #(
		.INIT('h0200)
	) name2763 (
		\ctl_rf_c4dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4992_
	);
	LUT4 #(
		.INIT('h0020)
	) name2764 (
		\ctl_rf_c2dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4993_
	);
	LUT4 #(
		.INIT('h0800)
	) name2765 (
		\ctl_rf_c5dmabs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4994_
	);
	LUT4 #(
		.INIT('h0001)
	) name2766 (
		_w4991_,
		_w4992_,
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT3 #(
		.INIT('h2a)
	) name2767 (
		_w3431_,
		_w4990_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('h0020)
	) name2768 (
		\ctl_rf_c2brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4997_
	);
	LUT4 #(
		.INIT('h0080)
	) name2769 (
		\ctl_rf_c3brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4998_
	);
	LUT4 #(
		.INIT('h0002)
	) name2770 (
		\ctl_rf_c0brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w4999_
	);
	LUT4 #(
		.INIT('h2000)
	) name2771 (
		\ctl_rf_c6brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5000_
	);
	LUT4 #(
		.INIT('h0001)
	) name2772 (
		_w4997_,
		_w4998_,
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT4 #(
		.INIT('h8000)
	) name2773 (
		\ctl_rf_c7brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5002_
	);
	LUT4 #(
		.INIT('h0200)
	) name2774 (
		\ctl_rf_c4brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5003_
	);
	LUT4 #(
		.INIT('h0008)
	) name2775 (
		\ctl_rf_c1brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5004_
	);
	LUT4 #(
		.INIT('h0800)
	) name2776 (
		\ctl_rf_c5brbs_reg[20]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5005_
	);
	LUT4 #(
		.INIT('h0001)
	) name2777 (
		_w5002_,
		_w5003_,
		_w5004_,
		_w5005_,
		_w5006_
	);
	LUT3 #(
		.INIT('h2a)
	) name2778 (
		_w3425_,
		_w5001_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2779 (
		\ctl_rf_abt_reg[4]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w5008_
	);
	LUT4 #(
		.INIT('h0023)
	) name2780 (
		\ctl_rf_c4_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w5009_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2782 (
		_w3422_,
		_w4996_,
		_w5007_,
		_w5010_,
		_w5011_
	);
	LUT4 #(
		.INIT('h4055)
	) name2783 (
		_w3622_,
		_w4969_,
		_w4985_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h4)
	) name2784 (
		_w4952_,
		_w5012_,
		_w5013_
	);
	LUT3 #(
		.INIT('h20)
	) name2785 (
		_w3503_,
		_w4313_,
		_w4324_,
		_w5014_
	);
	LUT3 #(
		.INIT('hc4)
	) name2786 (
		_w3427_,
		_w3503_,
		_w4346_,
		_w5015_
	);
	LUT3 #(
		.INIT('h13)
	) name2787 (
		_w4341_,
		_w5014_,
		_w5015_,
		_w5016_
	);
	LUT4 #(
		.INIT('h1311)
	) name2788 (
		_w3484_,
		_w3503_,
		_w4389_,
		_w4394_,
		_w5017_
	);
	LUT2 #(
		.INIT('h4)
	) name2789 (
		_w4388_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w3424_,
		_w4952_,
		_w5019_
	);
	LUT3 #(
		.INIT('hd0)
	) name2791 (
		_w5016_,
		_w5018_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		_w5013_,
		_w5020_,
		_w5021_
	);
	LUT3 #(
		.INIT('h2a)
	) name2793 (
		\hrdata_reg[5]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5022_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2794 (
		\ctl_rf_c0_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c0_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5023_
	);
	LUT3 #(
		.INIT('h20)
	) name2795 (
		\ctl_rf_c0_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5024_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name2796 (
		\haddr[8]_pad ,
		_w3445_,
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('h20)
	) name2797 (
		\ctl_rf_c3_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5026_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2798 (
		\ctl_rf_c3_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c3_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5027_
	);
	LUT3 #(
		.INIT('h8a)
	) name2799 (
		_w3457_,
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT3 #(
		.INIT('h80)
	) name2800 (
		\ctl_rf_c5_rf_chdad_reg[21]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5029_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2801 (
		\ctl_rf_c5_rf_chsad_reg[21]/NET0131 ,
		\ctl_rf_c5_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5030_
	);
	LUT3 #(
		.INIT('h8a)
	) name2802 (
		_w3436_,
		_w5029_,
		_w5030_,
		_w5031_
	);
	LUT3 #(
		.INIT('h20)
	) name2803 (
		\ctl_rf_c1_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5032_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2804 (
		\ctl_rf_c1_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c1_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5033_
	);
	LUT3 #(
		.INIT('h8a)
	) name2805 (
		_w3449_,
		_w5032_,
		_w5033_,
		_w5034_
	);
	LUT3 #(
		.INIT('h20)
	) name2806 (
		\ctl_rf_c4_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5035_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2807 (
		\ctl_rf_c4_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c4_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5036_
	);
	LUT3 #(
		.INIT('h8a)
	) name2808 (
		_w3426_,
		_w5035_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('h0001)
	) name2809 (
		_w5028_,
		_w5031_,
		_w5034_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		_w5025_,
		_w5038_,
		_w5039_
	);
	LUT4 #(
		.INIT('h135f)
	) name2811 (
		\ctl_rf_c2_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[21]/NET0131 ,
		_w3462_,
		_w3472_,
		_w5040_
	);
	LUT4 #(
		.INIT('h135f)
	) name2812 (
		\ctl_rf_c1_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[21]/NET0131 ,
		_w3474_,
		_w3477_,
		_w5041_
	);
	LUT4 #(
		.INIT('h153f)
	) name2813 (
		\ctl_rf_c5_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[21]/NET0131 ,
		_w3464_,
		_w3469_,
		_w5042_
	);
	LUT4 #(
		.INIT('h135f)
	) name2814 (
		\ctl_rf_c0_rf_chllp_reg[21]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[21]/NET0131 ,
		_w3467_,
		_w3479_,
		_w5043_
	);
	LUT4 #(
		.INIT('h8000)
	) name2815 (
		_w5040_,
		_w5041_,
		_w5042_,
		_w5043_,
		_w5044_
	);
	LUT3 #(
		.INIT('h80)
	) name2816 (
		\ctl_rf_c7_rf_chdad_reg[21]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5045_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name2817 (
		\ctl_rf_c7_rf_chsad_reg[21]/NET0131 ,
		\ctl_rf_c7_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5046_
	);
	LUT3 #(
		.INIT('h8a)
	) name2818 (
		_w3453_,
		_w5045_,
		_w5046_,
		_w5047_
	);
	LUT3 #(
		.INIT('h20)
	) name2819 (
		\ctl_rf_c6_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5048_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2820 (
		\ctl_rf_c6_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c6_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5049_
	);
	LUT3 #(
		.INIT('h8a)
	) name2821 (
		_w3440_,
		_w5048_,
		_w5049_,
		_w5050_
	);
	LUT3 #(
		.INIT('h20)
	) name2822 (
		\ctl_rf_c2_rf_chsad_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5051_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2823 (
		\ctl_rf_c2_rf_chdad_reg[21]/P0002 ,
		\ctl_rf_c2_rf_prot3_reg/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5052_
	);
	LUT3 #(
		.INIT('h8a)
	) name2824 (
		_w3432_,
		_w5051_,
		_w5052_,
		_w5053_
	);
	LUT3 #(
		.INIT('h01)
	) name2825 (
		_w5047_,
		_w5050_,
		_w5053_,
		_w5054_
	);
	LUT3 #(
		.INIT('hd0)
	) name2826 (
		_w3427_,
		_w5044_,
		_w5054_,
		_w5055_
	);
	LUT4 #(
		.INIT('h0008)
	) name2827 (
		\ctl_rf_c1brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5056_
	);
	LUT4 #(
		.INIT('h0080)
	) name2828 (
		\ctl_rf_c3brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5057_
	);
	LUT4 #(
		.INIT('h0002)
	) name2829 (
		\ctl_rf_c0brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5058_
	);
	LUT4 #(
		.INIT('h8000)
	) name2830 (
		\ctl_rf_c7brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5059_
	);
	LUT4 #(
		.INIT('h0001)
	) name2831 (
		_w5056_,
		_w5057_,
		_w5058_,
		_w5059_,
		_w5060_
	);
	LUT4 #(
		.INIT('h2000)
	) name2832 (
		\ctl_rf_c6brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5061_
	);
	LUT4 #(
		.INIT('h0200)
	) name2833 (
		\ctl_rf_c4brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5062_
	);
	LUT4 #(
		.INIT('h0020)
	) name2834 (
		\ctl_rf_c2brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5063_
	);
	LUT4 #(
		.INIT('h0800)
	) name2835 (
		\ctl_rf_c5brbs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5064_
	);
	LUT4 #(
		.INIT('h0001)
	) name2836 (
		_w5061_,
		_w5062_,
		_w5063_,
		_w5064_,
		_w5065_
	);
	LUT3 #(
		.INIT('h2a)
	) name2837 (
		_w3425_,
		_w5060_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('h0020)
	) name2838 (
		\ctl_rf_c2dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5067_
	);
	LUT4 #(
		.INIT('h0080)
	) name2839 (
		\ctl_rf_c3dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5068_
	);
	LUT4 #(
		.INIT('h0002)
	) name2840 (
		\ctl_rf_c0dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5069_
	);
	LUT4 #(
		.INIT('h2000)
	) name2841 (
		\ctl_rf_c6dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5070_
	);
	LUT4 #(
		.INIT('h0001)
	) name2842 (
		_w5067_,
		_w5068_,
		_w5069_,
		_w5070_,
		_w5071_
	);
	LUT4 #(
		.INIT('h8000)
	) name2843 (
		\ctl_rf_c7dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5072_
	);
	LUT4 #(
		.INIT('h0200)
	) name2844 (
		\ctl_rf_c4dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5073_
	);
	LUT4 #(
		.INIT('h0008)
	) name2845 (
		\ctl_rf_c1dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5074_
	);
	LUT4 #(
		.INIT('h0800)
	) name2846 (
		\ctl_rf_c5dmabs_reg[21]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5075_
	);
	LUT4 #(
		.INIT('h0001)
	) name2847 (
		_w5072_,
		_w5073_,
		_w5074_,
		_w5075_,
		_w5076_
	);
	LUT3 #(
		.INIT('h2a)
	) name2848 (
		_w3431_,
		_w5071_,
		_w5076_,
		_w5077_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2849 (
		\ctl_rf_abt_reg[5]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w5078_
	);
	LUT4 #(
		.INIT('h0023)
	) name2850 (
		\ctl_rf_c5_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w5079_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w5078_,
		_w5079_,
		_w5080_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2852 (
		_w3422_,
		_w5066_,
		_w5077_,
		_w5080_,
		_w5081_
	);
	LUT4 #(
		.INIT('h4055)
	) name2853 (
		_w3622_,
		_w5039_,
		_w5055_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h4)
	) name2854 (
		_w5022_,
		_w5082_,
		_w5083_
	);
	LUT3 #(
		.INIT('h20)
	) name2855 (
		_w3503_,
		_w4446_,
		_w4457_,
		_w5084_
	);
	LUT3 #(
		.INIT('hc4)
	) name2856 (
		_w3427_,
		_w3503_,
		_w4479_,
		_w5085_
	);
	LUT3 #(
		.INIT('h13)
	) name2857 (
		_w4474_,
		_w5084_,
		_w5085_,
		_w5086_
	);
	LUT4 #(
		.INIT('h1311)
	) name2858 (
		_w3484_,
		_w3503_,
		_w4522_,
		_w4527_,
		_w5087_
	);
	LUT2 #(
		.INIT('h4)
	) name2859 (
		_w4521_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w3424_,
		_w5022_,
		_w5089_
	);
	LUT3 #(
		.INIT('hd0)
	) name2861 (
		_w5086_,
		_w5088_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name2862 (
		_w5083_,
		_w5090_,
		_w5091_
	);
	LUT3 #(
		.INIT('h2a)
	) name2863 (
		\hrdata_reg[6]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5092_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2864 (
		\ctl_rf_c7_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c7_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5093_
	);
	LUT3 #(
		.INIT('h20)
	) name2865 (
		\ctl_rf_c7_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5094_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name2866 (
		\haddr[8]_pad ,
		_w3453_,
		_w5093_,
		_w5094_,
		_w5095_
	);
	LUT3 #(
		.INIT('h20)
	) name2867 (
		\ctl_rf_c6_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5096_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2868 (
		\ctl_rf_c6_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c6_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5097_
	);
	LUT3 #(
		.INIT('h8a)
	) name2869 (
		_w3440_,
		_w5096_,
		_w5097_,
		_w5098_
	);
	LUT3 #(
		.INIT('h80)
	) name2870 (
		\ctl_rf_c4_rf_chdad_reg[22]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5099_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2871 (
		\ctl_rf_c4_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5100_
	);
	LUT3 #(
		.INIT('h8a)
	) name2872 (
		_w3426_,
		_w5099_,
		_w5100_,
		_w5101_
	);
	LUT3 #(
		.INIT('h20)
	) name2873 (
		\ctl_rf_c0_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5102_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2874 (
		\ctl_rf_c0_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c0_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5103_
	);
	LUT3 #(
		.INIT('h8a)
	) name2875 (
		_w3445_,
		_w5102_,
		_w5103_,
		_w5104_
	);
	LUT3 #(
		.INIT('h20)
	) name2876 (
		\ctl_rf_c3_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5105_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2877 (
		\ctl_rf_c3_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c3_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5106_
	);
	LUT3 #(
		.INIT('h8a)
	) name2878 (
		_w3457_,
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT4 #(
		.INIT('h0001)
	) name2879 (
		_w5098_,
		_w5101_,
		_w5104_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name2880 (
		_w5095_,
		_w5108_,
		_w5109_
	);
	LUT4 #(
		.INIT('h135f)
	) name2881 (
		\ctl_rf_c1_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[22]/NET0131 ,
		_w3474_,
		_w3477_,
		_w5110_
	);
	LUT4 #(
		.INIT('h135f)
	) name2882 (
		\ctl_rf_c0_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[22]/NET0131 ,
		_w3467_,
		_w3479_,
		_w5111_
	);
	LUT4 #(
		.INIT('h135f)
	) name2883 (
		\ctl_rf_c2_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c4_rf_chllp_reg[22]/NET0131 ,
		_w3462_,
		_w3472_,
		_w5112_
	);
	LUT4 #(
		.INIT('h153f)
	) name2884 (
		\ctl_rf_c5_rf_chllp_reg[22]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[22]/NET0131 ,
		_w3464_,
		_w3469_,
		_w5113_
	);
	LUT4 #(
		.INIT('h8000)
	) name2885 (
		_w5110_,
		_w5111_,
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT3 #(
		.INIT('h80)
	) name2886 (
		\ctl_rf_c5_rf_chdad_reg[22]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5115_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2887 (
		\ctl_rf_c5_rf_chpri_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5116_
	);
	LUT3 #(
		.INIT('h8a)
	) name2888 (
		_w3436_,
		_w5115_,
		_w5116_,
		_w5117_
	);
	LUT3 #(
		.INIT('h20)
	) name2889 (
		\ctl_rf_c2_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5118_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2890 (
		\ctl_rf_c2_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c2_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5119_
	);
	LUT3 #(
		.INIT('h8a)
	) name2891 (
		_w3432_,
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT3 #(
		.INIT('h20)
	) name2892 (
		\ctl_rf_c1_rf_chsad_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5121_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2893 (
		\ctl_rf_c1_rf_chdad_reg[22]/P0002 ,
		\ctl_rf_c1_rf_chpri_reg[0]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5122_
	);
	LUT3 #(
		.INIT('h8a)
	) name2894 (
		_w3449_,
		_w5121_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h01)
	) name2895 (
		_w5117_,
		_w5120_,
		_w5123_,
		_w5124_
	);
	LUT3 #(
		.INIT('hd0)
	) name2896 (
		_w3427_,
		_w5114_,
		_w5124_,
		_w5125_
	);
	LUT4 #(
		.INIT('h0008)
	) name2897 (
		\ctl_rf_c1brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5126_
	);
	LUT4 #(
		.INIT('h0080)
	) name2898 (
		\ctl_rf_c3brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5127_
	);
	LUT4 #(
		.INIT('h0002)
	) name2899 (
		\ctl_rf_c0brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5128_
	);
	LUT4 #(
		.INIT('h8000)
	) name2900 (
		\ctl_rf_c7brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5129_
	);
	LUT4 #(
		.INIT('h0001)
	) name2901 (
		_w5126_,
		_w5127_,
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT4 #(
		.INIT('h2000)
	) name2902 (
		\ctl_rf_c6brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5131_
	);
	LUT4 #(
		.INIT('h0200)
	) name2903 (
		\ctl_rf_c4brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5132_
	);
	LUT4 #(
		.INIT('h0020)
	) name2904 (
		\ctl_rf_c2brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5133_
	);
	LUT4 #(
		.INIT('h0800)
	) name2905 (
		\ctl_rf_c5brbs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5134_
	);
	LUT4 #(
		.INIT('h0001)
	) name2906 (
		_w5131_,
		_w5132_,
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT3 #(
		.INIT('h2a)
	) name2907 (
		_w3425_,
		_w5130_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('h0020)
	) name2908 (
		\ctl_rf_c2dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5137_
	);
	LUT4 #(
		.INIT('h0080)
	) name2909 (
		\ctl_rf_c3dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5138_
	);
	LUT4 #(
		.INIT('h0002)
	) name2910 (
		\ctl_rf_c0dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5139_
	);
	LUT4 #(
		.INIT('h2000)
	) name2911 (
		\ctl_rf_c6dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5140_
	);
	LUT4 #(
		.INIT('h0001)
	) name2912 (
		_w5137_,
		_w5138_,
		_w5139_,
		_w5140_,
		_w5141_
	);
	LUT4 #(
		.INIT('h8000)
	) name2913 (
		\ctl_rf_c7dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5142_
	);
	LUT4 #(
		.INIT('h0200)
	) name2914 (
		\ctl_rf_c4dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5143_
	);
	LUT4 #(
		.INIT('h0008)
	) name2915 (
		\ctl_rf_c1dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5144_
	);
	LUT4 #(
		.INIT('h0800)
	) name2916 (
		\ctl_rf_c5dmabs_reg[22]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5145_
	);
	LUT4 #(
		.INIT('h0001)
	) name2917 (
		_w5142_,
		_w5143_,
		_w5144_,
		_w5145_,
		_w5146_
	);
	LUT3 #(
		.INIT('h2a)
	) name2918 (
		_w3431_,
		_w5141_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2919 (
		\ctl_rf_abt_reg[6]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w5148_
	);
	LUT4 #(
		.INIT('h0023)
	) name2920 (
		\ctl_rf_c6_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name2921 (
		_w5148_,
		_w5149_,
		_w5150_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2922 (
		_w3422_,
		_w5136_,
		_w5147_,
		_w5150_,
		_w5151_
	);
	LUT4 #(
		.INIT('h4055)
	) name2923 (
		_w3622_,
		_w5109_,
		_w5125_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h4)
	) name2924 (
		_w5092_,
		_w5152_,
		_w5153_
	);
	LUT3 #(
		.INIT('h20)
	) name2925 (
		_w3503_,
		_w4650_,
		_w4661_,
		_w5154_
	);
	LUT3 #(
		.INIT('hc4)
	) name2926 (
		_w3427_,
		_w3503_,
		_w4683_,
		_w5155_
	);
	LUT3 #(
		.INIT('h13)
	) name2927 (
		_w4678_,
		_w5154_,
		_w5155_,
		_w5156_
	);
	LUT4 #(
		.INIT('h1311)
	) name2928 (
		_w3484_,
		_w3503_,
		_w4726_,
		_w4731_,
		_w5157_
	);
	LUT2 #(
		.INIT('h4)
	) name2929 (
		_w4725_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h1)
	) name2930 (
		_w3424_,
		_w5092_,
		_w5159_
	);
	LUT3 #(
		.INIT('hd0)
	) name2931 (
		_w5156_,
		_w5158_,
		_w5159_,
		_w5160_
	);
	LUT2 #(
		.INIT('h1)
	) name2932 (
		_w5153_,
		_w5160_,
		_w5161_
	);
	LUT3 #(
		.INIT('h2a)
	) name2933 (
		\hrdata_reg[7]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5162_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2934 (
		\ctl_rf_c4_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c4_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5163_
	);
	LUT3 #(
		.INIT('h20)
	) name2935 (
		\ctl_rf_c4_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5164_
	);
	LUT4 #(
		.INIT('hdd5d)
	) name2936 (
		\haddr[8]_pad ,
		_w3426_,
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT3 #(
		.INIT('h20)
	) name2937 (
		\ctl_rf_c1_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5166_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2938 (
		\ctl_rf_c1_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c1_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5167_
	);
	LUT3 #(
		.INIT('h8a)
	) name2939 (
		_w3449_,
		_w5166_,
		_w5167_,
		_w5168_
	);
	LUT3 #(
		.INIT('h80)
	) name2940 (
		\ctl_rf_c6_rf_chdad_reg[23]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5169_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2941 (
		\ctl_rf_c6_rf_chpri_reg[1]/NET0131 ,
		\ctl_rf_c6_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5170_
	);
	LUT3 #(
		.INIT('h8a)
	) name2942 (
		_w3440_,
		_w5169_,
		_w5170_,
		_w5171_
	);
	LUT3 #(
		.INIT('h20)
	) name2943 (
		\ctl_rf_c0_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5172_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2944 (
		\ctl_rf_c0_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c0_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5173_
	);
	LUT3 #(
		.INIT('h8a)
	) name2945 (
		_w3445_,
		_w5172_,
		_w5173_,
		_w5174_
	);
	LUT3 #(
		.INIT('h20)
	) name2946 (
		\ctl_rf_c2_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5175_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2947 (
		\ctl_rf_c2_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c2_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5176_
	);
	LUT3 #(
		.INIT('h8a)
	) name2948 (
		_w3432_,
		_w5175_,
		_w5176_,
		_w5177_
	);
	LUT4 #(
		.INIT('h0001)
	) name2949 (
		_w5168_,
		_w5171_,
		_w5174_,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h4)
	) name2950 (
		_w5165_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('h135f)
	) name2951 (
		\ctl_rf_c0_rf_chllp_reg[23]/NET0131 ,
		\ctl_rf_c5_rf_chllp_reg[23]/NET0131 ,
		_w3467_,
		_w3469_,
		_w5180_
	);
	LUT4 #(
		.INIT('h135f)
	) name2952 (
		\ctl_rf_c2_rf_chllp_reg[23]/NET0131 ,
		\ctl_rf_c6_rf_chllp_reg[23]/NET0131 ,
		_w3462_,
		_w3479_,
		_w5181_
	);
	LUT4 #(
		.INIT('h135f)
	) name2953 (
		\ctl_rf_c1_rf_chllp_reg[23]/NET0131 ,
		\ctl_rf_c3_rf_chllp_reg[23]/NET0131 ,
		_w3474_,
		_w3477_,
		_w5182_
	);
	LUT4 #(
		.INIT('h153f)
	) name2954 (
		\ctl_rf_c4_rf_chllp_reg[23]/NET0131 ,
		\ctl_rf_c7_rf_chllp_reg[23]/NET0131 ,
		_w3464_,
		_w3472_,
		_w5183_
	);
	LUT4 #(
		.INIT('h8000)
	) name2955 (
		_w5180_,
		_w5181_,
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('h80)
	) name2956 (
		\ctl_rf_c5_rf_chdad_reg[23]/P0002 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5185_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name2957 (
		\ctl_rf_c5_rf_chpri_reg[1]/NET0131 ,
		\ctl_rf_c5_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5186_
	);
	LUT3 #(
		.INIT('h8a)
	) name2958 (
		_w3436_,
		_w5185_,
		_w5186_,
		_w5187_
	);
	LUT3 #(
		.INIT('h20)
	) name2959 (
		\ctl_rf_c3_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5188_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2960 (
		\ctl_rf_c3_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c3_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5189_
	);
	LUT3 #(
		.INIT('h8a)
	) name2961 (
		_w3457_,
		_w5188_,
		_w5189_,
		_w5190_
	);
	LUT3 #(
		.INIT('h20)
	) name2962 (
		\ctl_rf_c7_rf_chsad_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5191_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name2963 (
		\ctl_rf_c7_rf_chdad_reg[23]/P0002 ,
		\ctl_rf_c7_rf_chpri_reg[1]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		_w5192_
	);
	LUT3 #(
		.INIT('h8a)
	) name2964 (
		_w3453_,
		_w5191_,
		_w5192_,
		_w5193_
	);
	LUT3 #(
		.INIT('h01)
	) name2965 (
		_w5187_,
		_w5190_,
		_w5193_,
		_w5194_
	);
	LUT3 #(
		.INIT('hd0)
	) name2966 (
		_w3427_,
		_w5184_,
		_w5194_,
		_w5195_
	);
	LUT4 #(
		.INIT('h0008)
	) name2967 (
		\ctl_rf_c1brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5196_
	);
	LUT4 #(
		.INIT('h0080)
	) name2968 (
		\ctl_rf_c3brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5197_
	);
	LUT4 #(
		.INIT('h0002)
	) name2969 (
		\ctl_rf_c0brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5198_
	);
	LUT4 #(
		.INIT('h8000)
	) name2970 (
		\ctl_rf_c7brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5199_
	);
	LUT4 #(
		.INIT('h0001)
	) name2971 (
		_w5196_,
		_w5197_,
		_w5198_,
		_w5199_,
		_w5200_
	);
	LUT4 #(
		.INIT('h2000)
	) name2972 (
		\ctl_rf_c6brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5201_
	);
	LUT4 #(
		.INIT('h0200)
	) name2973 (
		\ctl_rf_c4brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5202_
	);
	LUT4 #(
		.INIT('h0020)
	) name2974 (
		\ctl_rf_c2brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5203_
	);
	LUT4 #(
		.INIT('h0800)
	) name2975 (
		\ctl_rf_c5brbs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5204_
	);
	LUT4 #(
		.INIT('h0001)
	) name2976 (
		_w5201_,
		_w5202_,
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT3 #(
		.INIT('h2a)
	) name2977 (
		_w3425_,
		_w5200_,
		_w5205_,
		_w5206_
	);
	LUT4 #(
		.INIT('h0020)
	) name2978 (
		\ctl_rf_c2dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5207_
	);
	LUT4 #(
		.INIT('h0080)
	) name2979 (
		\ctl_rf_c3dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5208_
	);
	LUT4 #(
		.INIT('h0002)
	) name2980 (
		\ctl_rf_c0dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5209_
	);
	LUT4 #(
		.INIT('h2000)
	) name2981 (
		\ctl_rf_c6dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5210_
	);
	LUT4 #(
		.INIT('h0001)
	) name2982 (
		_w5207_,
		_w5208_,
		_w5209_,
		_w5210_,
		_w5211_
	);
	LUT4 #(
		.INIT('h8000)
	) name2983 (
		\ctl_rf_c7dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5212_
	);
	LUT4 #(
		.INIT('h0200)
	) name2984 (
		\ctl_rf_c4dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5213_
	);
	LUT4 #(
		.INIT('h0008)
	) name2985 (
		\ctl_rf_c1dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5214_
	);
	LUT4 #(
		.INIT('h0800)
	) name2986 (
		\ctl_rf_c5dmabs_reg[23]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[3]_pad ,
		\haddr[4]_pad ,
		_w5215_
	);
	LUT4 #(
		.INIT('h0001)
	) name2987 (
		_w5212_,
		_w5213_,
		_w5214_,
		_w5215_,
		_w5216_
	);
	LUT3 #(
		.INIT('h2a)
	) name2988 (
		_w3431_,
		_w5211_,
		_w5216_,
		_w5217_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2989 (
		\ctl_rf_abt_reg[7]/NET0131 ,
		\haddr[6]_pad ,
		\haddr[7]_pad ,
		\haddr[8]_pad ,
		_w5218_
	);
	LUT4 #(
		.INIT('h0023)
	) name2990 (
		\ctl_rf_c7_rf_int_abt_msk_reg/NET0131 ,
		\haddr[8]_pad ,
		_w3613_,
		_w3614_,
		_w5219_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		_w5218_,
		_w5219_,
		_w5220_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2992 (
		_w3422_,
		_w5206_,
		_w5217_,
		_w5220_,
		_w5221_
	);
	LUT4 #(
		.INIT('h4055)
	) name2993 (
		_w3622_,
		_w5179_,
		_w5195_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name2994 (
		_w5162_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('haa80)
	) name2995 (
		_w3503_,
		_w4789_,
		_w4805_,
		_w4828_,
		_w5224_
	);
	LUT4 #(
		.INIT('h1311)
	) name2996 (
		_w3484_,
		_w3503_,
		_w4870_,
		_w4875_,
		_w5225_
	);
	LUT2 #(
		.INIT('h4)
	) name2997 (
		_w4869_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name2998 (
		_w3424_,
		_w5162_,
		_w5227_
	);
	LUT3 #(
		.INIT('he0)
	) name2999 (
		_w5224_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h1)
	) name3000 (
		_w5223_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		_w5230_
	);
	LUT4 #(
		.INIT('h8000)
	) name3002 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w5231_
	);
	LUT4 #(
		.INIT('h8000)
	) name3003 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w5230_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3004 (
		\hwdata[29]_pad ,
		\hwdata[5]_pad ,
		_w2234_,
		_w2235_,
		_w5233_
	);
	LUT2 #(
		.INIT('h8)
	) name3005 (
		\hwdata[21]_pad ,
		_w2234_,
		_w5234_
	);
	LUT4 #(
		.INIT('heee2)
	) name3006 (
		\ctl_rf_c1_rf_chtsz_reg[5]/NET0131 ,
		_w5232_,
		_w5233_,
		_w5234_,
		_w5235_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3007 (
		\hwdata[30]_pad ,
		\hwdata[6]_pad ,
		_w2234_,
		_w2235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\hwdata[22]_pad ,
		_w2234_,
		_w5237_
	);
	LUT4 #(
		.INIT('heee2)
	) name3009 (
		\ctl_rf_c1_rf_chtsz_reg[6]/NET0131 ,
		_w5232_,
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3010 (
		\ctl_rf_c1_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5232_,
		_w5239_
	);
	LUT4 #(
		.INIT('h8000)
	) name3011 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2232_,
		_w2244_,
		_w5240_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3012 (
		\ctl_rf_c3_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5240_,
		_w5241_
	);
	LUT4 #(
		.INIT('h8000)
	) name3013 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2244_,
		_w5230_,
		_w5231_,
		_w5242_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3014 (
		\ctl_rf_c3_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5242_,
		_w5243_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3015 (
		\ctl_rf_c3_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5242_,
		_w5244_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3016 (
		\ctl_rf_c3_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5242_,
		_w5245_
	);
	LUT4 #(
		.INIT('h8000)
	) name3017 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2247_,
		_w2249_,
		_w5246_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3018 (
		\ctl_rf_c4_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5246_,
		_w5247_
	);
	LUT4 #(
		.INIT('h2000)
	) name3019 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w5248_
	);
	LUT4 #(
		.INIT('h8000)
	) name3020 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2247_,
		_w5230_,
		_w5248_,
		_w5249_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3021 (
		\ctl_rf_c4_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5249_,
		_w5250_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3022 (
		\ctl_rf_c4_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5249_,
		_w5251_
	);
	LUT4 #(
		.INIT('h8000)
	) name3023 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2232_,
		_w2247_,
		_w5252_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3024 (
		\ctl_rf_c5_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5252_,
		_w5253_
	);
	LUT4 #(
		.INIT('h8000)
	) name3025 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2247_,
		_w5230_,
		_w5231_,
		_w5254_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3026 (
		\ctl_rf_c5_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5254_,
		_w5255_
	);
	LUT4 #(
		.INIT('h8000)
	) name3027 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2249_,
		_w2254_,
		_w5256_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3028 (
		\ctl_rf_c6_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5256_,
		_w5257_
	);
	LUT4 #(
		.INIT('h2000)
	) name3029 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		_w5258_
	);
	LUT4 #(
		.INIT('h8000)
	) name3030 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2248_,
		_w2254_,
		_w5258_,
		_w5259_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3031 (
		\ctl_rf_c6_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5259_,
		_w5260_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3032 (
		\ctl_rf_c6_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5259_,
		_w5261_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3033 (
		\ctl_rf_c6_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5259_,
		_w5262_
	);
	LUT4 #(
		.INIT('h8000)
	) name3034 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2232_,
		_w2254_,
		_w5263_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3035 (
		\ctl_rf_c7_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5263_,
		_w5264_
	);
	LUT4 #(
		.INIT('h8000)
	) name3036 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2231_,
		_w2254_,
		_w5258_,
		_w5265_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3037 (
		\ctl_rf_c7_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5265_,
		_w5266_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3038 (
		\ctl_rf_c7_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5265_,
		_w5267_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3039 (
		\ctl_rf_c7_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5265_,
		_w5268_
	);
	LUT4 #(
		.INIT('h8000)
	) name3040 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2230_,
		_w2249_,
		_w5269_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3041 (
		\ctl_rf_c0_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5269_,
		_w5270_
	);
	LUT4 #(
		.INIT('h8000)
	) name3042 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w5230_,
		_w5248_,
		_w5271_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3043 (
		\ctl_rf_c0_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5271_,
		_w5272_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3044 (
		\ctl_rf_c0_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5271_,
		_w5273_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3045 (
		\ctl_rf_c0_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5271_,
		_w5274_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3046 (
		\hwdata[28]_pad ,
		\hwdata[4]_pad ,
		_w2234_,
		_w2235_,
		_w5275_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		\hwdata[20]_pad ,
		_w2234_,
		_w5276_
	);
	LUT4 #(
		.INIT('heee2)
	) name3048 (
		\ctl_rf_c1_rf_chtsz_reg[4]/NET0131 ,
		_w5232_,
		_w5275_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('h8000)
	) name3049 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2230_,
		_w2244_,
		_w2249_,
		_w5278_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3050 (
		\ctl_rf_c2_rf_chsad_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5278_,
		_w5279_
	);
	LUT4 #(
		.INIT('h8000)
	) name3051 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2244_,
		_w5230_,
		_w5248_,
		_w5280_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3052 (
		\ctl_rf_c2_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5280_,
		_w5281_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3053 (
		\ctl_rf_c2_rf_chtsz_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5280_,
		_w5282_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3054 (
		\ctl_rf_c2_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5280_,
		_w5283_
	);
	LUT4 #(
		.INIT('heee2)
	) name3055 (
		\ctl_rf_c3_rf_chtsz_reg[4]/NET0131 ,
		_w5242_,
		_w5275_,
		_w5276_,
		_w5284_
	);
	LUT4 #(
		.INIT('heee2)
	) name3056 (
		\ctl_rf_c4_rf_chtsz_reg[4]/NET0131 ,
		_w5249_,
		_w5275_,
		_w5276_,
		_w5285_
	);
	LUT4 #(
		.INIT('heee2)
	) name3057 (
		\ctl_rf_c6_rf_chtsz_reg[4]/NET0131 ,
		_w5259_,
		_w5275_,
		_w5276_,
		_w5286_
	);
	LUT4 #(
		.INIT('heee2)
	) name3058 (
		\ctl_rf_c7_rf_chtsz_reg[4]/NET0131 ,
		_w5265_,
		_w5275_,
		_w5276_,
		_w5287_
	);
	LUT4 #(
		.INIT('h8000)
	) name3059 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w2232_,
		_w2239_,
		_w5288_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3060 (
		\hwdata[10]_pad ,
		\hwdata[18]_pad ,
		_w2234_,
		_w2235_,
		_w5289_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		\hwdata[26]_pad ,
		_w2234_,
		_w5290_
	);
	LUT4 #(
		.INIT('heee2)
	) name3062 (
		\ctl_rf_c1_rf_chdad_reg[10]/NET0131 ,
		_w5288_,
		_w5289_,
		_w5290_,
		_w5291_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3063 (
		\hwdata[12]_pad ,
		\hwdata[20]_pad ,
		_w2234_,
		_w2235_,
		_w5292_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		\hwdata[28]_pad ,
		_w2234_,
		_w5293_
	);
	LUT4 #(
		.INIT('heee2)
	) name3065 (
		\ctl_rf_c1_rf_chdad_reg[12]/NET0131 ,
		_w5288_,
		_w5292_,
		_w5293_,
		_w5294_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3066 (
		\ctl_rf_c1_rf_chdad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5288_,
		_w5295_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3067 (
		\hwdata[16]_pad ,
		\hwdata[8]_pad ,
		_w2234_,
		_w2235_,
		_w5296_
	);
	LUT2 #(
		.INIT('h8)
	) name3068 (
		\hwdata[24]_pad ,
		_w2234_,
		_w5297_
	);
	LUT4 #(
		.INIT('heee2)
	) name3069 (
		\ctl_rf_c1_rf_chdad_reg[8]/NET0131 ,
		_w5288_,
		_w5296_,
		_w5297_,
		_w5298_
	);
	LUT4 #(
		.INIT('h8000)
	) name3070 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w2230_,
		_w2232_,
		_w5299_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3071 (
		\hwdata[11]_pad ,
		\hwdata[19]_pad ,
		_w2234_,
		_w2235_,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name3072 (
		\hwdata[27]_pad ,
		_w2234_,
		_w5301_
	);
	LUT4 #(
		.INIT('heee2)
	) name3073 (
		\ctl_rf_c1_rf_chsad_reg[11]/NET0131 ,
		_w5299_,
		_w5300_,
		_w5301_,
		_w5302_
	);
	LUT4 #(
		.INIT('heee2)
	) name3074 (
		\ctl_rf_c1_rf_chsad_reg[5]/NET0131 ,
		_w2233_,
		_w5233_,
		_w5234_,
		_w5303_
	);
	LUT4 #(
		.INIT('heee2)
	) name3075 (
		\ctl_rf_c1_rf_chsad_reg[6]/NET0131 ,
		_w2233_,
		_w5236_,
		_w5237_,
		_w5304_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3076 (
		\hwdata[17]_pad ,
		\hwdata[9]_pad ,
		_w2234_,
		_w2235_,
		_w5305_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		\hwdata[25]_pad ,
		_w2234_,
		_w5306_
	);
	LUT4 #(
		.INIT('heee2)
	) name3078 (
		\ctl_rf_c1_rf_chsad_reg[9]/NET0131 ,
		_w5299_,
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('h8000)
	) name3079 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2232_,
		_w2239_,
		_w2244_,
		_w5308_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3080 (
		\ctl_rf_c3_rf_chdad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5308_,
		_w5309_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3081 (
		\ctl_rf_c3_rf_chdad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5308_,
		_w5310_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3082 (
		\ctl_rf_c3_rf_chdad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5308_,
		_w5311_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3083 (
		\ctl_rf_c3_rf_chdad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5308_,
		_w5312_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3084 (
		\ctl_rf_c3_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5308_,
		_w5313_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3085 (
		\ctl_rf_c3_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5240_,
		_w5314_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3086 (
		\ctl_rf_c3_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5240_,
		_w5315_
	);
	LUT4 #(
		.INIT('h8000)
	) name3087 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2232_,
		_w2244_,
		_w5316_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3088 (
		\ctl_rf_c3_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5316_,
		_w5317_
	);
	LUT4 #(
		.INIT('h8000)
	) name3089 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2239_,
		_w2247_,
		_w2249_,
		_w5318_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3090 (
		\ctl_rf_c4_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h8000)
	) name3091 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2247_,
		_w2249_,
		_w5320_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3092 (
		\ctl_rf_c4_rf_chsad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5320_,
		_w5321_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3093 (
		\ctl_rf_c4_rf_chsad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5320_,
		_w5322_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3094 (
		\ctl_rf_c4_rf_chsad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5320_,
		_w5323_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3095 (
		\ctl_rf_c4_rf_chsad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5320_,
		_w5324_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3096 (
		\ctl_rf_c4_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5246_,
		_w5325_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3097 (
		\ctl_rf_c4_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5246_,
		_w5326_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3098 (
		\ctl_rf_c4_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5320_,
		_w5327_
	);
	LUT4 #(
		.INIT('h8000)
	) name3099 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2232_,
		_w2239_,
		_w2247_,
		_w5328_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3100 (
		\ctl_rf_c5_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5328_,
		_w5329_
	);
	LUT4 #(
		.INIT('h8000)
	) name3101 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2232_,
		_w2247_,
		_w5330_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3102 (
		\ctl_rf_c5_rf_chsad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3103 (
		\ctl_rf_c5_rf_chsad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5330_,
		_w5332_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3104 (
		\ctl_rf_c5_rf_chsad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5330_,
		_w5333_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3105 (
		\ctl_rf_c5_rf_chsad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5330_,
		_w5334_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3106 (
		\ctl_rf_c5_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5252_,
		_w5335_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3107 (
		\ctl_rf_c5_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5252_,
		_w5336_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3108 (
		\ctl_rf_c5_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5330_,
		_w5337_
	);
	LUT4 #(
		.INIT('h8000)
	) name3109 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2239_,
		_w2249_,
		_w2254_,
		_w5338_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3110 (
		\ctl_rf_c6_rf_chdad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5338_,
		_w5339_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3111 (
		\ctl_rf_c6_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5338_,
		_w5340_
	);
	LUT4 #(
		.INIT('h8000)
	) name3112 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2249_,
		_w2254_,
		_w5341_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3113 (
		\ctl_rf_c6_rf_chsad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5341_,
		_w5342_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3114 (
		\ctl_rf_c6_rf_chsad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5341_,
		_w5343_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3115 (
		\ctl_rf_c6_rf_chsad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5341_,
		_w5344_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3116 (
		\ctl_rf_c6_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5256_,
		_w5345_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3117 (
		\ctl_rf_c6_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5256_,
		_w5346_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3118 (
		\ctl_rf_c6_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5341_,
		_w5347_
	);
	LUT4 #(
		.INIT('h8000)
	) name3119 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2232_,
		_w2239_,
		_w2254_,
		_w5348_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3120 (
		\ctl_rf_c7_rf_chdad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3121 (
		\ctl_rf_c7_rf_chdad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5348_,
		_w5350_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3122 (
		\ctl_rf_c7_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5348_,
		_w5351_
	);
	LUT4 #(
		.INIT('h8000)
	) name3123 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2232_,
		_w2254_,
		_w5352_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3124 (
		\ctl_rf_c7_rf_chsad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5352_,
		_w5353_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3125 (
		\ctl_rf_c7_rf_chsad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5352_,
		_w5354_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3126 (
		\ctl_rf_c7_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5263_,
		_w5355_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3127 (
		\ctl_rf_c7_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5263_,
		_w5356_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3128 (
		\ctl_rf_c7_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5352_,
		_w5357_
	);
	LUT4 #(
		.INIT('heee2)
	) name3129 (
		\ctl_rf_c1_rf_chsad_reg[0]/NET0131 ,
		_w2233_,
		_w2996_,
		_w2997_,
		_w5358_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3130 (
		\hwdata[1]_pad ,
		\hwdata[25]_pad ,
		_w2234_,
		_w2235_,
		_w5359_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		\hwdata[17]_pad ,
		_w2234_,
		_w5360_
	);
	LUT4 #(
		.INIT('heee2)
	) name3132 (
		\ctl_rf_c1_rf_chsad_reg[1]/NET0131 ,
		_w2233_,
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3133 (
		\hwdata[26]_pad ,
		\hwdata[2]_pad ,
		_w2234_,
		_w2235_,
		_w5362_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		\hwdata[18]_pad ,
		_w2234_,
		_w5363_
	);
	LUT4 #(
		.INIT('heee2)
	) name3135 (
		\ctl_rf_c1_rf_chsad_reg[2]/NET0131 ,
		_w2233_,
		_w5362_,
		_w5363_,
		_w5364_
	);
	LUT4 #(
		.INIT('heee2)
	) name3136 (
		\ctl_rf_c1_rf_chsad_reg[4]/NET0131 ,
		_w2233_,
		_w5275_,
		_w5276_,
		_w5365_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3137 (
		\ctl_rf_c3_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5240_,
		_w5366_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3138 (
		\hwdata[13]_pad ,
		\hwdata[21]_pad ,
		_w2234_,
		_w2235_,
		_w5367_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		\hwdata[29]_pad ,
		_w2234_,
		_w5368_
	);
	LUT4 #(
		.INIT('heee2)
	) name3140 (
		\ctl_rf_c3_rf_chsad_reg[13]/NET0131 ,
		_w5316_,
		_w5367_,
		_w5368_,
		_w5369_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3141 (
		\hwdata[14]_pad ,
		\hwdata[22]_pad ,
		_w2234_,
		_w2235_,
		_w5370_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		\hwdata[30]_pad ,
		_w2234_,
		_w5371_
	);
	LUT4 #(
		.INIT('heee2)
	) name3143 (
		\ctl_rf_c3_rf_chsad_reg[14]/NET0131 ,
		_w5316_,
		_w5370_,
		_w5371_,
		_w5372_
	);
	LUT4 #(
		.INIT('heee2)
	) name3144 (
		\ctl_rf_c3_rf_chsad_reg[1]/NET0131 ,
		_w5240_,
		_w5359_,
		_w5360_,
		_w5373_
	);
	LUT4 #(
		.INIT('heee2)
	) name3145 (
		\ctl_rf_c3_rf_chsad_reg[2]/NET0131 ,
		_w5240_,
		_w5362_,
		_w5363_,
		_w5374_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3146 (
		\hwdata[27]_pad ,
		\hwdata[3]_pad ,
		_w2234_,
		_w2235_,
		_w5375_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		\hwdata[19]_pad ,
		_w2234_,
		_w5376_
	);
	LUT4 #(
		.INIT('heee2)
	) name3148 (
		\ctl_rf_c3_rf_chsad_reg[3]/NET0131 ,
		_w5240_,
		_w5375_,
		_w5376_,
		_w5377_
	);
	LUT4 #(
		.INIT('heee2)
	) name3149 (
		\ctl_rf_c3_rf_chsad_reg[4]/NET0131 ,
		_w5240_,
		_w5275_,
		_w5276_,
		_w5378_
	);
	LUT4 #(
		.INIT('h8000)
	) name3150 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2247_,
		_w2249_,
		_w5379_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3151 (
		\ctl_rf_c4_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5379_,
		_w5380_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3152 (
		\ctl_rf_c4_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5379_,
		_w5381_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3153 (
		\ctl_rf_c4_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5379_,
		_w5382_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3154 (
		\ctl_rf_c4_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5246_,
		_w5383_
	);
	LUT4 #(
		.INIT('heee2)
	) name3155 (
		\ctl_rf_c4_rf_chsad_reg[13]/NET0131 ,
		_w5320_,
		_w5367_,
		_w5368_,
		_w5384_
	);
	LUT4 #(
		.INIT('heee2)
	) name3156 (
		\ctl_rf_c4_rf_chsad_reg[14]/NET0131 ,
		_w5320_,
		_w5370_,
		_w5371_,
		_w5385_
	);
	LUT4 #(
		.INIT('heee2)
	) name3157 (
		\ctl_rf_c4_rf_chsad_reg[1]/NET0131 ,
		_w5246_,
		_w5359_,
		_w5360_,
		_w5386_
	);
	LUT4 #(
		.INIT('heee2)
	) name3158 (
		\ctl_rf_c4_rf_chsad_reg[2]/NET0131 ,
		_w5246_,
		_w5362_,
		_w5363_,
		_w5387_
	);
	LUT4 #(
		.INIT('heee2)
	) name3159 (
		\ctl_rf_c4_rf_chsad_reg[3]/NET0131 ,
		_w5246_,
		_w5375_,
		_w5376_,
		_w5388_
	);
	LUT4 #(
		.INIT('heee2)
	) name3160 (
		\ctl_rf_c4_rf_chsad_reg[4]/NET0131 ,
		_w5246_,
		_w5275_,
		_w5276_,
		_w5389_
	);
	LUT4 #(
		.INIT('h8000)
	) name3161 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2249_,
		_w2254_,
		_w5390_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3162 (
		\ctl_rf_c6_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5390_,
		_w5391_
	);
	LUT4 #(
		.INIT('heee2)
	) name3163 (
		\ctl_rf_c6_rf_chdad_reg[13]/NET0131 ,
		_w5338_,
		_w5367_,
		_w5368_,
		_w5392_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3164 (
		\ctl_rf_c6_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5390_,
		_w5393_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3165 (
		\ctl_rf_c6_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5390_,
		_w5394_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3166 (
		\ctl_rf_c6_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5256_,
		_w5395_
	);
	LUT4 #(
		.INIT('heee2)
	) name3167 (
		\ctl_rf_c6_rf_chsad_reg[14]/NET0131 ,
		_w5341_,
		_w5370_,
		_w5371_,
		_w5396_
	);
	LUT4 #(
		.INIT('heee2)
	) name3168 (
		\ctl_rf_c6_rf_chsad_reg[1]/NET0131 ,
		_w5256_,
		_w5359_,
		_w5360_,
		_w5397_
	);
	LUT4 #(
		.INIT('heee2)
	) name3169 (
		\ctl_rf_c6_rf_chsad_reg[2]/NET0131 ,
		_w5256_,
		_w5362_,
		_w5363_,
		_w5398_
	);
	LUT4 #(
		.INIT('heee2)
	) name3170 (
		\ctl_rf_c6_rf_chsad_reg[3]/NET0131 ,
		_w5256_,
		_w5375_,
		_w5376_,
		_w5399_
	);
	LUT4 #(
		.INIT('heee2)
	) name3171 (
		\ctl_rf_c6_rf_chsad_reg[4]/NET0131 ,
		_w5256_,
		_w5275_,
		_w5276_,
		_w5400_
	);
	LUT4 #(
		.INIT('h8000)
	) name3172 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2239_,
		_w2249_,
		_w5401_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3173 (
		\ctl_rf_c0_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5401_,
		_w5402_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3174 (
		\ctl_rf_c0_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5401_,
		_w5403_
	);
	LUT4 #(
		.INIT('h8000)
	) name3175 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w2239_,
		_w2249_,
		_w5404_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3176 (
		\ctl_rf_c0_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3177 (
		\ctl_rf_c0_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5269_,
		_w5406_
	);
	LUT4 #(
		.INIT('h8000)
	) name3178 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w2230_,
		_w2249_,
		_w5407_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3179 (
		\ctl_rf_c0_rf_chsad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5407_,
		_w5408_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3180 (
		\ctl_rf_c0_rf_chsad_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5407_,
		_w5409_
	);
	LUT4 #(
		.INIT('heee2)
	) name3181 (
		\ctl_rf_c0_rf_chsad_reg[1]/NET0131 ,
		_w5269_,
		_w5359_,
		_w5360_,
		_w5410_
	);
	LUT4 #(
		.INIT('heee2)
	) name3182 (
		\ctl_rf_c0_rf_chsad_reg[2]/NET0131 ,
		_w5269_,
		_w5362_,
		_w5363_,
		_w5411_
	);
	LUT4 #(
		.INIT('heee2)
	) name3183 (
		\ctl_rf_c0_rf_chsad_reg[3]/NET0131 ,
		_w5269_,
		_w5375_,
		_w5376_,
		_w5412_
	);
	LUT4 #(
		.INIT('heee2)
	) name3184 (
		\ctl_rf_c0_rf_chsad_reg[4]/NET0131 ,
		_w5269_,
		_w5275_,
		_w5276_,
		_w5413_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3185 (
		\ctl_rf_c0_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5269_,
		_w5414_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3186 (
		\ctl_rf_c0_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5269_,
		_w5415_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3187 (
		\ctl_rf_c0_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5407_,
		_w5416_
	);
	LUT4 #(
		.INIT('heee2)
	) name3188 (
		\ctl_rf_c0_rf_chtsz_reg[4]/NET0131 ,
		_w5271_,
		_w5275_,
		_w5276_,
		_w5417_
	);
	LUT4 #(
		.INIT('h8000)
	) name3189 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2232_,
		_w2239_,
		_w5418_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3190 (
		\ctl_rf_c1_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5418_,
		_w5419_
	);
	LUT4 #(
		.INIT('heee2)
	) name3191 (
		\ctl_rf_c1_rf_chdad_reg[13]/NET0131 ,
		_w5288_,
		_w5367_,
		_w5368_,
		_w5420_
	);
	LUT4 #(
		.INIT('heee2)
	) name3192 (
		\ctl_rf_c1_rf_chdad_reg[14]/NET0131 ,
		_w5288_,
		_w5370_,
		_w5371_,
		_w5421_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3193 (
		\ctl_rf_c1_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5418_,
		_w5422_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3194 (
		\ctl_rf_c1_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5418_,
		_w5423_
	);
	LUT4 #(
		.INIT('h8000)
	) name3195 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2244_,
		_w2249_,
		_w5424_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3196 (
		\ctl_rf_c2_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5424_,
		_w5425_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3197 (
		\ctl_rf_c2_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5424_,
		_w5426_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3198 (
		\ctl_rf_c2_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5424_,
		_w5427_
	);
	LUT4 #(
		.INIT('h8000)
	) name3199 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2239_,
		_w2244_,
		_w2249_,
		_w5428_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3200 (
		\ctl_rf_c2_rf_chdad_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5428_,
		_w5429_
	);
	LUT4 #(
		.INIT('h8000)
	) name3201 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2230_,
		_w2244_,
		_w2249_,
		_w5430_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3202 (
		\ctl_rf_c2_rf_chsad_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5430_,
		_w5431_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3203 (
		\ctl_rf_c2_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5278_,
		_w5432_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3204 (
		\ctl_rf_c2_rf_chsad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5430_,
		_w5433_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3205 (
		\ctl_rf_c2_rf_chsad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5430_,
		_w5434_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3206 (
		\ctl_rf_c2_rf_chsad_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5430_,
		_w5435_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3207 (
		\ctl_rf_c2_rf_chsad_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5430_,
		_w5436_
	);
	LUT4 #(
		.INIT('heee2)
	) name3208 (
		\ctl_rf_c2_rf_chsad_reg[1]/NET0131 ,
		_w5278_,
		_w5359_,
		_w5360_,
		_w5437_
	);
	LUT4 #(
		.INIT('heee2)
	) name3209 (
		\ctl_rf_c2_rf_chsad_reg[2]/NET0131 ,
		_w5278_,
		_w5362_,
		_w5363_,
		_w5438_
	);
	LUT4 #(
		.INIT('heee2)
	) name3210 (
		\ctl_rf_c2_rf_chsad_reg[3]/NET0131 ,
		_w5278_,
		_w5375_,
		_w5376_,
		_w5439_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3211 (
		\ctl_rf_c2_rf_chsad_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5278_,
		_w5440_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3212 (
		\ctl_rf_c2_rf_chsad_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5278_,
		_w5441_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3213 (
		\ctl_rf_c2_rf_chsad_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5278_,
		_w5442_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3214 (
		\ctl_rf_c2_rf_chsad_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5430_,
		_w5443_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3215 (
		\ctl_rf_c2_rf_chtsz_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5280_,
		_w5444_
	);
	LUT4 #(
		.INIT('h8000)
	) name3216 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2232_,
		_w2239_,
		_w2244_,
		_w5445_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3217 (
		\ctl_rf_c3_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5445_,
		_w5446_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3218 (
		\ctl_rf_c3_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5445_,
		_w5447_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3219 (
		\ctl_rf_c3_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5445_,
		_w5448_
	);
	LUT4 #(
		.INIT('h8000)
	) name3220 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2232_,
		_w2239_,
		_w2247_,
		_w5449_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3221 (
		\ctl_rf_c5_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('heee2)
	) name3222 (
		\ctl_rf_c5_rf_chdad_reg[13]/NET0131 ,
		_w5328_,
		_w5367_,
		_w5368_,
		_w5451_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3223 (
		\ctl_rf_c5_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5449_,
		_w5452_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3224 (
		\ctl_rf_c5_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5252_,
		_w5453_
	);
	LUT4 #(
		.INIT('heee2)
	) name3225 (
		\ctl_rf_c5_rf_chsad_reg[14]/NET0131 ,
		_w5330_,
		_w5370_,
		_w5371_,
		_w5454_
	);
	LUT4 #(
		.INIT('heee2)
	) name3226 (
		\ctl_rf_c5_rf_chsad_reg[1]/NET0131 ,
		_w5252_,
		_w5359_,
		_w5360_,
		_w5455_
	);
	LUT4 #(
		.INIT('heee2)
	) name3227 (
		\ctl_rf_c5_rf_chsad_reg[2]/NET0131 ,
		_w5252_,
		_w5362_,
		_w5363_,
		_w5456_
	);
	LUT4 #(
		.INIT('heee2)
	) name3228 (
		\ctl_rf_c5_rf_chsad_reg[3]/NET0131 ,
		_w5252_,
		_w5375_,
		_w5376_,
		_w5457_
	);
	LUT4 #(
		.INIT('heee2)
	) name3229 (
		\ctl_rf_c5_rf_chsad_reg[4]/NET0131 ,
		_w5252_,
		_w5275_,
		_w5276_,
		_w5458_
	);
	LUT4 #(
		.INIT('h8000)
	) name3230 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2232_,
		_w2239_,
		_w2254_,
		_w5459_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3231 (
		\ctl_rf_c7_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5459_,
		_w5460_
	);
	LUT4 #(
		.INIT('heee2)
	) name3232 (
		\ctl_rf_c7_rf_chdad_reg[13]/NET0131 ,
		_w5348_,
		_w5367_,
		_w5368_,
		_w5461_
	);
	LUT4 #(
		.INIT('heee2)
	) name3233 (
		\ctl_rf_c7_rf_chdad_reg[14]/NET0131 ,
		_w5348_,
		_w5370_,
		_w5371_,
		_w5462_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3234 (
		\ctl_rf_c7_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5459_,
		_w5463_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3235 (
		\ctl_rf_c7_rf_chdad_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5459_,
		_w5464_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3236 (
		\ctl_rf_c7_rf_chsad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5263_,
		_w5465_
	);
	LUT4 #(
		.INIT('heee2)
	) name3237 (
		\ctl_rf_c7_rf_chsad_reg[1]/NET0131 ,
		_w5263_,
		_w5359_,
		_w5360_,
		_w5466_
	);
	LUT4 #(
		.INIT('heee2)
	) name3238 (
		\ctl_rf_c7_rf_chsad_reg[2]/NET0131 ,
		_w5263_,
		_w5362_,
		_w5363_,
		_w5467_
	);
	LUT4 #(
		.INIT('heee2)
	) name3239 (
		\ctl_rf_c7_rf_chsad_reg[3]/NET0131 ,
		_w5263_,
		_w5375_,
		_w5376_,
		_w5468_
	);
	LUT4 #(
		.INIT('heee2)
	) name3240 (
		\ctl_rf_c7_rf_chsad_reg[4]/NET0131 ,
		_w5263_,
		_w5275_,
		_w5276_,
		_w5469_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3241 (
		\ctl_rf_c0_rf_chdad_reg[0]/NET0131 ,
		_w2996_,
		_w2997_,
		_w5401_,
		_w5470_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3242 (
		\ctl_rf_c0_rf_chdad_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5404_,
		_w5471_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3243 (
		\ctl_rf_c0_rf_chdad_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5404_,
		_w5472_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3244 (
		\ctl_rf_c0_rf_chdad_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5404_,
		_w5473_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3245 (
		\ctl_rf_c0_rf_chdad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5404_,
		_w5474_
	);
	LUT3 #(
		.INIT('h40)
	) name3246 (
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		\m1_mux_hrp_df_reg[0]/NET0131 ,
		_w5475_
	);
	LUT4 #(
		.INIT('h8000)
	) name3247 (
		\m1_mux_hrp_df_reg[0]/NET0131 ,
		_w2390_,
		_w2393_,
		_w2396_,
		_w5476_
	);
	LUT4 #(
		.INIT('h070f)
	) name3248 (
		_w2403_,
		_w2416_,
		_w5475_,
		_w5476_,
		_w5477_
	);
	LUT3 #(
		.INIT('h8c)
	) name3249 (
		\ctl_rf_c4dmabs_reg[16]/NET0131 ,
		\ctl_rf_c4dmabs_reg[17]/NET0131 ,
		\ctl_rf_c4dmabs_reg[22]/NET0131 ,
		_w5478_
	);
	LUT4 #(
		.INIT('h000b)
	) name3250 (
		\ctl_rf_c4dmabs_reg[16]/NET0131 ,
		\ctl_rf_c4dmabs_reg[20]/NET0131 ,
		\ctl_rf_c4dmabs_reg[21]/NET0131 ,
		\ctl_rf_c4dmabs_reg[22]/NET0131 ,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		\ctl_rf_c4dmabs_reg[18]/NET0131 ,
		\ctl_rf_c4dmabs_reg[19]/NET0131 ,
		_w5480_
	);
	LUT4 #(
		.INIT('hab00)
	) name3252 (
		\ctl_rf_c4dmabs_reg[23]/NET0131 ,
		_w5478_,
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT4 #(
		.INIT('h0001)
	) name3253 (
		\ctl_rf_c4dmabs_reg[28]/NET0131 ,
		\ctl_rf_c4dmabs_reg[29]/NET0131 ,
		\ctl_rf_c4dmabs_reg[30]/NET0131 ,
		\ctl_rf_c4dmabs_reg[31]/NET0131 ,
		_w5482_
	);
	LUT4 #(
		.INIT('h0001)
	) name3254 (
		\ctl_rf_c4dmabs_reg[24]/NET0131 ,
		\ctl_rf_c4dmabs_reg[25]/NET0131 ,
		\ctl_rf_c4dmabs_reg[26]/NET0131 ,
		\ctl_rf_c4dmabs_reg[27]/NET0131 ,
		_w5483_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		_w5482_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h4)
	) name3256 (
		_w5481_,
		_w5484_,
		_w5485_
	);
	LUT3 #(
		.INIT('h8c)
	) name3257 (
		\ctl_rf_c6dmabs_reg[16]/NET0131 ,
		\ctl_rf_c6dmabs_reg[17]/NET0131 ,
		\ctl_rf_c6dmabs_reg[22]/NET0131 ,
		_w5486_
	);
	LUT4 #(
		.INIT('h000b)
	) name3258 (
		\ctl_rf_c6dmabs_reg[16]/NET0131 ,
		\ctl_rf_c6dmabs_reg[20]/NET0131 ,
		\ctl_rf_c6dmabs_reg[21]/NET0131 ,
		\ctl_rf_c6dmabs_reg[22]/NET0131 ,
		_w5487_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		\ctl_rf_c6dmabs_reg[18]/NET0131 ,
		\ctl_rf_c6dmabs_reg[19]/NET0131 ,
		_w5488_
	);
	LUT4 #(
		.INIT('hab00)
	) name3260 (
		\ctl_rf_c6dmabs_reg[23]/NET0131 ,
		_w5486_,
		_w5487_,
		_w5488_,
		_w5489_
	);
	LUT4 #(
		.INIT('h0001)
	) name3261 (
		\ctl_rf_c6dmabs_reg[28]/NET0131 ,
		\ctl_rf_c6dmabs_reg[29]/NET0131 ,
		\ctl_rf_c6dmabs_reg[30]/NET0131 ,
		\ctl_rf_c6dmabs_reg[31]/NET0131 ,
		_w5490_
	);
	LUT4 #(
		.INIT('h0001)
	) name3262 (
		\ctl_rf_c6dmabs_reg[24]/NET0131 ,
		\ctl_rf_c6dmabs_reg[25]/NET0131 ,
		\ctl_rf_c6dmabs_reg[26]/NET0131 ,
		\ctl_rf_c6dmabs_reg[27]/NET0131 ,
		_w5491_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		_w5490_,
		_w5491_,
		_w5492_
	);
	LUT2 #(
		.INIT('h4)
	) name3264 (
		_w5489_,
		_w5492_,
		_w5493_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3265 (
		_w5481_,
		_w5484_,
		_w5489_,
		_w5492_,
		_w5494_
	);
	LUT3 #(
		.INIT('h8c)
	) name3266 (
		\ctl_rf_c3dmabs_reg[16]/NET0131 ,
		\ctl_rf_c3dmabs_reg[17]/NET0131 ,
		\ctl_rf_c3dmabs_reg[22]/NET0131 ,
		_w5495_
	);
	LUT4 #(
		.INIT('h000b)
	) name3267 (
		\ctl_rf_c3dmabs_reg[16]/NET0131 ,
		\ctl_rf_c3dmabs_reg[20]/NET0131 ,
		\ctl_rf_c3dmabs_reg[21]/NET0131 ,
		\ctl_rf_c3dmabs_reg[22]/NET0131 ,
		_w5496_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		\ctl_rf_c3dmabs_reg[18]/NET0131 ,
		\ctl_rf_c3dmabs_reg[19]/NET0131 ,
		_w5497_
	);
	LUT4 #(
		.INIT('hab00)
	) name3269 (
		\ctl_rf_c3dmabs_reg[23]/NET0131 ,
		_w5495_,
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT4 #(
		.INIT('h0001)
	) name3270 (
		\ctl_rf_c3dmabs_reg[28]/NET0131 ,
		\ctl_rf_c3dmabs_reg[29]/NET0131 ,
		\ctl_rf_c3dmabs_reg[30]/NET0131 ,
		\ctl_rf_c3dmabs_reg[31]/NET0131 ,
		_w5499_
	);
	LUT4 #(
		.INIT('h0001)
	) name3271 (
		\ctl_rf_c3dmabs_reg[24]/NET0131 ,
		\ctl_rf_c3dmabs_reg[25]/NET0131 ,
		\ctl_rf_c3dmabs_reg[26]/NET0131 ,
		\ctl_rf_c3dmabs_reg[27]/NET0131 ,
		_w5500_
	);
	LUT2 #(
		.INIT('h8)
	) name3272 (
		_w5499_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h4)
	) name3273 (
		_w5498_,
		_w5501_,
		_w5502_
	);
	LUT3 #(
		.INIT('h8c)
	) name3274 (
		\ctl_rf_c5dmabs_reg[16]/NET0131 ,
		\ctl_rf_c5dmabs_reg[17]/NET0131 ,
		\ctl_rf_c5dmabs_reg[22]/NET0131 ,
		_w5503_
	);
	LUT4 #(
		.INIT('h000b)
	) name3275 (
		\ctl_rf_c5dmabs_reg[16]/NET0131 ,
		\ctl_rf_c5dmabs_reg[20]/NET0131 ,
		\ctl_rf_c5dmabs_reg[21]/NET0131 ,
		\ctl_rf_c5dmabs_reg[22]/NET0131 ,
		_w5504_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		\ctl_rf_c5dmabs_reg[18]/NET0131 ,
		\ctl_rf_c5dmabs_reg[19]/NET0131 ,
		_w5505_
	);
	LUT4 #(
		.INIT('hab00)
	) name3277 (
		\ctl_rf_c5dmabs_reg[23]/NET0131 ,
		_w5503_,
		_w5504_,
		_w5505_,
		_w5506_
	);
	LUT4 #(
		.INIT('h0001)
	) name3278 (
		\ctl_rf_c5dmabs_reg[28]/NET0131 ,
		\ctl_rf_c5dmabs_reg[29]/NET0131 ,
		\ctl_rf_c5dmabs_reg[30]/NET0131 ,
		\ctl_rf_c5dmabs_reg[31]/NET0131 ,
		_w5507_
	);
	LUT4 #(
		.INIT('h0001)
	) name3279 (
		\ctl_rf_c5dmabs_reg[24]/NET0131 ,
		\ctl_rf_c5dmabs_reg[25]/NET0131 ,
		\ctl_rf_c5dmabs_reg[26]/NET0131 ,
		\ctl_rf_c5dmabs_reg[27]/NET0131 ,
		_w5508_
	);
	LUT2 #(
		.INIT('h8)
	) name3280 (
		_w5507_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h4)
	) name3281 (
		_w5506_,
		_w5509_,
		_w5510_
	);
	LUT3 #(
		.INIT('h8c)
	) name3282 (
		\ctl_rf_c7dmabs_reg[16]/NET0131 ,
		\ctl_rf_c7dmabs_reg[17]/NET0131 ,
		\ctl_rf_c7dmabs_reg[22]/NET0131 ,
		_w5511_
	);
	LUT4 #(
		.INIT('h000b)
	) name3283 (
		\ctl_rf_c7dmabs_reg[16]/NET0131 ,
		\ctl_rf_c7dmabs_reg[20]/NET0131 ,
		\ctl_rf_c7dmabs_reg[21]/NET0131 ,
		\ctl_rf_c7dmabs_reg[22]/NET0131 ,
		_w5512_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		\ctl_rf_c7dmabs_reg[18]/NET0131 ,
		\ctl_rf_c7dmabs_reg[19]/NET0131 ,
		_w5513_
	);
	LUT4 #(
		.INIT('hab00)
	) name3285 (
		\ctl_rf_c7dmabs_reg[23]/NET0131 ,
		_w5511_,
		_w5512_,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h0001)
	) name3286 (
		\ctl_rf_c7dmabs_reg[28]/NET0131 ,
		\ctl_rf_c7dmabs_reg[29]/NET0131 ,
		\ctl_rf_c7dmabs_reg[30]/NET0131 ,
		\ctl_rf_c7dmabs_reg[31]/NET0131 ,
		_w5515_
	);
	LUT4 #(
		.INIT('h0001)
	) name3287 (
		\ctl_rf_c7dmabs_reg[24]/NET0131 ,
		\ctl_rf_c7dmabs_reg[25]/NET0131 ,
		\ctl_rf_c7dmabs_reg[26]/NET0131 ,
		\ctl_rf_c7dmabs_reg[27]/NET0131 ,
		_w5516_
	);
	LUT2 #(
		.INIT('h8)
	) name3288 (
		_w5515_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h4)
	) name3289 (
		_w5514_,
		_w5517_,
		_w5518_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3290 (
		_w5506_,
		_w5509_,
		_w5514_,
		_w5517_,
		_w5519_
	);
	LUT3 #(
		.INIT('h8c)
	) name3291 (
		\ctl_rf_c2dmabs_reg[16]/NET0131 ,
		\ctl_rf_c2dmabs_reg[17]/NET0131 ,
		\ctl_rf_c2dmabs_reg[22]/NET0131 ,
		_w5520_
	);
	LUT4 #(
		.INIT('h000b)
	) name3292 (
		\ctl_rf_c2dmabs_reg[16]/NET0131 ,
		\ctl_rf_c2dmabs_reg[20]/NET0131 ,
		\ctl_rf_c2dmabs_reg[21]/NET0131 ,
		\ctl_rf_c2dmabs_reg[22]/NET0131 ,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		\ctl_rf_c2dmabs_reg[18]/NET0131 ,
		\ctl_rf_c2dmabs_reg[19]/NET0131 ,
		_w5522_
	);
	LUT4 #(
		.INIT('hab00)
	) name3294 (
		\ctl_rf_c2dmabs_reg[23]/NET0131 ,
		_w5520_,
		_w5521_,
		_w5522_,
		_w5523_
	);
	LUT4 #(
		.INIT('h0001)
	) name3295 (
		\ctl_rf_c2dmabs_reg[28]/NET0131 ,
		\ctl_rf_c2dmabs_reg[29]/NET0131 ,
		\ctl_rf_c2dmabs_reg[30]/NET0131 ,
		\ctl_rf_c2dmabs_reg[31]/NET0131 ,
		_w5524_
	);
	LUT4 #(
		.INIT('h0001)
	) name3296 (
		\ctl_rf_c2dmabs_reg[24]/NET0131 ,
		\ctl_rf_c2dmabs_reg[25]/NET0131 ,
		\ctl_rf_c2dmabs_reg[26]/NET0131 ,
		\ctl_rf_c2dmabs_reg[27]/NET0131 ,
		_w5525_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		_w5524_,
		_w5525_,
		_w5526_
	);
	LUT2 #(
		.INIT('h4)
	) name3298 (
		_w5523_,
		_w5526_,
		_w5527_
	);
	LUT3 #(
		.INIT('h8c)
	) name3299 (
		\ctl_rf_c1dmabs_reg[16]/NET0131 ,
		\ctl_rf_c1dmabs_reg[17]/NET0131 ,
		\ctl_rf_c1dmabs_reg[22]/NET0131 ,
		_w5528_
	);
	LUT4 #(
		.INIT('h000b)
	) name3300 (
		\ctl_rf_c1dmabs_reg[16]/NET0131 ,
		\ctl_rf_c1dmabs_reg[20]/NET0131 ,
		\ctl_rf_c1dmabs_reg[21]/NET0131 ,
		\ctl_rf_c1dmabs_reg[22]/NET0131 ,
		_w5529_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		\ctl_rf_c1dmabs_reg[18]/NET0131 ,
		\ctl_rf_c1dmabs_reg[19]/NET0131 ,
		_w5530_
	);
	LUT4 #(
		.INIT('hab00)
	) name3302 (
		\ctl_rf_c1dmabs_reg[23]/NET0131 ,
		_w5528_,
		_w5529_,
		_w5530_,
		_w5531_
	);
	LUT4 #(
		.INIT('h0001)
	) name3303 (
		\ctl_rf_c1dmabs_reg[28]/NET0131 ,
		\ctl_rf_c1dmabs_reg[29]/NET0131 ,
		\ctl_rf_c1dmabs_reg[30]/NET0131 ,
		\ctl_rf_c1dmabs_reg[31]/NET0131 ,
		_w5532_
	);
	LUT4 #(
		.INIT('h0001)
	) name3304 (
		\ctl_rf_c1dmabs_reg[24]/NET0131 ,
		\ctl_rf_c1dmabs_reg[25]/NET0131 ,
		\ctl_rf_c1dmabs_reg[26]/NET0131 ,
		\ctl_rf_c1dmabs_reg[27]/NET0131 ,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name3305 (
		_w5532_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h4)
	) name3306 (
		_w5531_,
		_w5534_,
		_w5535_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3307 (
		_w5523_,
		_w5526_,
		_w5531_,
		_w5534_,
		_w5536_
	);
	LUT4 #(
		.INIT('h2000)
	) name3308 (
		_w5494_,
		_w5502_,
		_w5519_,
		_w5536_,
		_w5537_
	);
	LUT3 #(
		.INIT('h8c)
	) name3309 (
		\ctl_rf_c0dmabs_reg[16]/NET0131 ,
		\ctl_rf_c0dmabs_reg[17]/NET0131 ,
		\ctl_rf_c0dmabs_reg[22]/NET0131 ,
		_w5538_
	);
	LUT4 #(
		.INIT('h000b)
	) name3310 (
		\ctl_rf_c0dmabs_reg[16]/NET0131 ,
		\ctl_rf_c0dmabs_reg[20]/NET0131 ,
		\ctl_rf_c0dmabs_reg[21]/NET0131 ,
		\ctl_rf_c0dmabs_reg[22]/NET0131 ,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		\ctl_rf_c0dmabs_reg[18]/NET0131 ,
		\ctl_rf_c0dmabs_reg[19]/NET0131 ,
		_w5540_
	);
	LUT4 #(
		.INIT('hab00)
	) name3312 (
		\ctl_rf_c0dmabs_reg[23]/NET0131 ,
		_w5538_,
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('h0001)
	) name3313 (
		\ctl_rf_c0dmabs_reg[28]/NET0131 ,
		\ctl_rf_c0dmabs_reg[29]/NET0131 ,
		\ctl_rf_c0dmabs_reg[30]/NET0131 ,
		\ctl_rf_c0dmabs_reg[31]/NET0131 ,
		_w5542_
	);
	LUT4 #(
		.INIT('h0001)
	) name3314 (
		\ctl_rf_c0dmabs_reg[24]/NET0131 ,
		\ctl_rf_c0dmabs_reg[25]/NET0131 ,
		\ctl_rf_c0dmabs_reg[26]/NET0131 ,
		\ctl_rf_c0dmabs_reg[27]/NET0131 ,
		_w5543_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		_w5542_,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		_w5541_,
		_w5544_,
		_w5545_
	);
	LUT3 #(
		.INIT('h8c)
	) name3317 (
		\ctl_rf_c0brbs_reg[16]/NET0131 ,
		\ctl_rf_c0brbs_reg[17]/NET0131 ,
		\ctl_rf_c0brbs_reg[22]/NET0131 ,
		_w5546_
	);
	LUT4 #(
		.INIT('h000b)
	) name3318 (
		\ctl_rf_c0brbs_reg[16]/NET0131 ,
		\ctl_rf_c0brbs_reg[20]/NET0131 ,
		\ctl_rf_c0brbs_reg[21]/NET0131 ,
		\ctl_rf_c0brbs_reg[22]/NET0131 ,
		_w5547_
	);
	LUT2 #(
		.INIT('h1)
	) name3319 (
		\ctl_rf_c0brbs_reg[18]/NET0131 ,
		\ctl_rf_c0brbs_reg[19]/NET0131 ,
		_w5548_
	);
	LUT4 #(
		.INIT('hab00)
	) name3320 (
		\ctl_rf_c0brbs_reg[23]/NET0131 ,
		_w5546_,
		_w5547_,
		_w5548_,
		_w5549_
	);
	LUT4 #(
		.INIT('h0001)
	) name3321 (
		\ctl_rf_c0brbs_reg[28]/NET0131 ,
		\ctl_rf_c0brbs_reg[29]/NET0131 ,
		\ctl_rf_c0brbs_reg[30]/NET0131 ,
		\ctl_rf_c0brbs_reg[31]/NET0131 ,
		_w5550_
	);
	LUT4 #(
		.INIT('h0001)
	) name3322 (
		\ctl_rf_c0brbs_reg[24]/NET0131 ,
		\ctl_rf_c0brbs_reg[25]/NET0131 ,
		\ctl_rf_c0brbs_reg[26]/NET0131 ,
		\ctl_rf_c0brbs_reg[27]/NET0131 ,
		_w5551_
	);
	LUT2 #(
		.INIT('h8)
	) name3323 (
		_w5550_,
		_w5551_,
		_w5552_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		_w5549_,
		_w5552_,
		_w5553_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3325 (
		_w5541_,
		_w5544_,
		_w5549_,
		_w5552_,
		_w5554_
	);
	LUT3 #(
		.INIT('h8c)
	) name3326 (
		\ctl_rf_c1brbs_reg[16]/NET0131 ,
		\ctl_rf_c1brbs_reg[17]/NET0131 ,
		\ctl_rf_c1brbs_reg[22]/NET0131 ,
		_w5555_
	);
	LUT4 #(
		.INIT('h000b)
	) name3327 (
		\ctl_rf_c1brbs_reg[16]/NET0131 ,
		\ctl_rf_c1brbs_reg[20]/NET0131 ,
		\ctl_rf_c1brbs_reg[21]/NET0131 ,
		\ctl_rf_c1brbs_reg[22]/NET0131 ,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		\ctl_rf_c1brbs_reg[18]/NET0131 ,
		\ctl_rf_c1brbs_reg[19]/NET0131 ,
		_w5557_
	);
	LUT4 #(
		.INIT('hab00)
	) name3329 (
		\ctl_rf_c1brbs_reg[23]/NET0131 ,
		_w5555_,
		_w5556_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('h0001)
	) name3330 (
		\ctl_rf_c1brbs_reg[28]/NET0131 ,
		\ctl_rf_c1brbs_reg[29]/NET0131 ,
		\ctl_rf_c1brbs_reg[30]/NET0131 ,
		\ctl_rf_c1brbs_reg[31]/NET0131 ,
		_w5559_
	);
	LUT4 #(
		.INIT('h0001)
	) name3331 (
		\ctl_rf_c1brbs_reg[24]/NET0131 ,
		\ctl_rf_c1brbs_reg[25]/NET0131 ,
		\ctl_rf_c1brbs_reg[26]/NET0131 ,
		\ctl_rf_c1brbs_reg[27]/NET0131 ,
		_w5560_
	);
	LUT2 #(
		.INIT('h8)
	) name3332 (
		_w5559_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h4)
	) name3333 (
		_w5558_,
		_w5561_,
		_w5562_
	);
	LUT3 #(
		.INIT('h8c)
	) name3334 (
		\ctl_rf_c2brbs_reg[16]/NET0131 ,
		\ctl_rf_c2brbs_reg[17]/NET0131 ,
		\ctl_rf_c2brbs_reg[22]/NET0131 ,
		_w5563_
	);
	LUT4 #(
		.INIT('h000b)
	) name3335 (
		\ctl_rf_c2brbs_reg[16]/NET0131 ,
		\ctl_rf_c2brbs_reg[20]/NET0131 ,
		\ctl_rf_c2brbs_reg[21]/NET0131 ,
		\ctl_rf_c2brbs_reg[22]/NET0131 ,
		_w5564_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		\ctl_rf_c2brbs_reg[18]/NET0131 ,
		\ctl_rf_c2brbs_reg[19]/NET0131 ,
		_w5565_
	);
	LUT4 #(
		.INIT('hab00)
	) name3337 (
		\ctl_rf_c2brbs_reg[23]/NET0131 ,
		_w5563_,
		_w5564_,
		_w5565_,
		_w5566_
	);
	LUT4 #(
		.INIT('h0001)
	) name3338 (
		\ctl_rf_c2brbs_reg[28]/NET0131 ,
		\ctl_rf_c2brbs_reg[29]/NET0131 ,
		\ctl_rf_c2brbs_reg[30]/NET0131 ,
		\ctl_rf_c2brbs_reg[31]/NET0131 ,
		_w5567_
	);
	LUT4 #(
		.INIT('h0001)
	) name3339 (
		\ctl_rf_c2brbs_reg[24]/NET0131 ,
		\ctl_rf_c2brbs_reg[25]/NET0131 ,
		\ctl_rf_c2brbs_reg[26]/NET0131 ,
		\ctl_rf_c2brbs_reg[27]/NET0131 ,
		_w5568_
	);
	LUT2 #(
		.INIT('h8)
	) name3340 (
		_w5567_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('h4)
	) name3341 (
		_w5566_,
		_w5569_,
		_w5570_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3342 (
		_w5558_,
		_w5561_,
		_w5566_,
		_w5569_,
		_w5571_
	);
	LUT2 #(
		.INIT('h8)
	) name3343 (
		_w5554_,
		_w5571_,
		_w5572_
	);
	LUT4 #(
		.INIT('h007f)
	) name3344 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w2431_,
		_w5573_
	);
	LUT3 #(
		.INIT('h8c)
	) name3345 (
		\ctl_rf_c6brbs_reg[16]/NET0131 ,
		\ctl_rf_c6brbs_reg[17]/NET0131 ,
		\ctl_rf_c6brbs_reg[22]/NET0131 ,
		_w5574_
	);
	LUT4 #(
		.INIT('h000b)
	) name3346 (
		\ctl_rf_c6brbs_reg[16]/NET0131 ,
		\ctl_rf_c6brbs_reg[20]/NET0131 ,
		\ctl_rf_c6brbs_reg[21]/NET0131 ,
		\ctl_rf_c6brbs_reg[22]/NET0131 ,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		\ctl_rf_c6brbs_reg[18]/NET0131 ,
		\ctl_rf_c6brbs_reg[19]/NET0131 ,
		_w5576_
	);
	LUT4 #(
		.INIT('hab00)
	) name3348 (
		\ctl_rf_c6brbs_reg[23]/NET0131 ,
		_w5574_,
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT4 #(
		.INIT('h0001)
	) name3349 (
		\ctl_rf_c6brbs_reg[28]/NET0131 ,
		\ctl_rf_c6brbs_reg[29]/NET0131 ,
		\ctl_rf_c6brbs_reg[30]/NET0131 ,
		\ctl_rf_c6brbs_reg[31]/NET0131 ,
		_w5578_
	);
	LUT4 #(
		.INIT('h0001)
	) name3350 (
		\ctl_rf_c6brbs_reg[24]/NET0131 ,
		\ctl_rf_c6brbs_reg[25]/NET0131 ,
		\ctl_rf_c6brbs_reg[26]/NET0131 ,
		\ctl_rf_c6brbs_reg[27]/NET0131 ,
		_w5579_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w5578_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		_w5577_,
		_w5580_,
		_w5581_
	);
	LUT3 #(
		.INIT('h8c)
	) name3353 (
		\ctl_rf_c7brbs_reg[16]/NET0131 ,
		\ctl_rf_c7brbs_reg[17]/NET0131 ,
		\ctl_rf_c7brbs_reg[22]/NET0131 ,
		_w5582_
	);
	LUT4 #(
		.INIT('h000b)
	) name3354 (
		\ctl_rf_c7brbs_reg[16]/NET0131 ,
		\ctl_rf_c7brbs_reg[20]/NET0131 ,
		\ctl_rf_c7brbs_reg[21]/NET0131 ,
		\ctl_rf_c7brbs_reg[22]/NET0131 ,
		_w5583_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		\ctl_rf_c7brbs_reg[18]/NET0131 ,
		\ctl_rf_c7brbs_reg[19]/NET0131 ,
		_w5584_
	);
	LUT4 #(
		.INIT('hab00)
	) name3356 (
		\ctl_rf_c7brbs_reg[23]/NET0131 ,
		_w5582_,
		_w5583_,
		_w5584_,
		_w5585_
	);
	LUT4 #(
		.INIT('h0001)
	) name3357 (
		\ctl_rf_c7brbs_reg[28]/NET0131 ,
		\ctl_rf_c7brbs_reg[29]/NET0131 ,
		\ctl_rf_c7brbs_reg[30]/NET0131 ,
		\ctl_rf_c7brbs_reg[31]/NET0131 ,
		_w5586_
	);
	LUT4 #(
		.INIT('h0001)
	) name3358 (
		\ctl_rf_c7brbs_reg[24]/NET0131 ,
		\ctl_rf_c7brbs_reg[25]/NET0131 ,
		\ctl_rf_c7brbs_reg[26]/NET0131 ,
		\ctl_rf_c7brbs_reg[27]/NET0131 ,
		_w5587_
	);
	LUT2 #(
		.INIT('h8)
	) name3359 (
		_w5586_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name3360 (
		_w5585_,
		_w5588_,
		_w5589_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3361 (
		_w5577_,
		_w5580_,
		_w5585_,
		_w5588_,
		_w5590_
	);
	LUT3 #(
		.INIT('h8c)
	) name3362 (
		\ctl_rf_c5brbs_reg[16]/NET0131 ,
		\ctl_rf_c5brbs_reg[17]/NET0131 ,
		\ctl_rf_c5brbs_reg[22]/NET0131 ,
		_w5591_
	);
	LUT4 #(
		.INIT('h000b)
	) name3363 (
		\ctl_rf_c5brbs_reg[16]/NET0131 ,
		\ctl_rf_c5brbs_reg[20]/NET0131 ,
		\ctl_rf_c5brbs_reg[21]/NET0131 ,
		\ctl_rf_c5brbs_reg[22]/NET0131 ,
		_w5592_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		\ctl_rf_c5brbs_reg[18]/NET0131 ,
		\ctl_rf_c5brbs_reg[19]/NET0131 ,
		_w5593_
	);
	LUT4 #(
		.INIT('hab00)
	) name3365 (
		\ctl_rf_c5brbs_reg[23]/NET0131 ,
		_w5591_,
		_w5592_,
		_w5593_,
		_w5594_
	);
	LUT4 #(
		.INIT('h0001)
	) name3366 (
		\ctl_rf_c5brbs_reg[28]/NET0131 ,
		\ctl_rf_c5brbs_reg[29]/NET0131 ,
		\ctl_rf_c5brbs_reg[30]/NET0131 ,
		\ctl_rf_c5brbs_reg[31]/NET0131 ,
		_w5595_
	);
	LUT4 #(
		.INIT('h0001)
	) name3367 (
		\ctl_rf_c5brbs_reg[24]/NET0131 ,
		\ctl_rf_c5brbs_reg[25]/NET0131 ,
		\ctl_rf_c5brbs_reg[26]/NET0131 ,
		\ctl_rf_c5brbs_reg[27]/NET0131 ,
		_w5596_
	);
	LUT2 #(
		.INIT('h8)
	) name3368 (
		_w5595_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h4)
	) name3369 (
		_w5594_,
		_w5597_,
		_w5598_
	);
	LUT3 #(
		.INIT('h8c)
	) name3370 (
		\ctl_rf_c3brbs_reg[16]/NET0131 ,
		\ctl_rf_c3brbs_reg[17]/NET0131 ,
		\ctl_rf_c3brbs_reg[22]/NET0131 ,
		_w5599_
	);
	LUT4 #(
		.INIT('h000b)
	) name3371 (
		\ctl_rf_c3brbs_reg[16]/NET0131 ,
		\ctl_rf_c3brbs_reg[20]/NET0131 ,
		\ctl_rf_c3brbs_reg[21]/NET0131 ,
		\ctl_rf_c3brbs_reg[22]/NET0131 ,
		_w5600_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		\ctl_rf_c3brbs_reg[18]/NET0131 ,
		\ctl_rf_c3brbs_reg[19]/NET0131 ,
		_w5601_
	);
	LUT4 #(
		.INIT('hab00)
	) name3373 (
		\ctl_rf_c3brbs_reg[23]/NET0131 ,
		_w5599_,
		_w5600_,
		_w5601_,
		_w5602_
	);
	LUT4 #(
		.INIT('h0001)
	) name3374 (
		\ctl_rf_c3brbs_reg[28]/NET0131 ,
		\ctl_rf_c3brbs_reg[29]/NET0131 ,
		\ctl_rf_c3brbs_reg[30]/NET0131 ,
		\ctl_rf_c3brbs_reg[31]/NET0131 ,
		_w5603_
	);
	LUT4 #(
		.INIT('h0001)
	) name3375 (
		\ctl_rf_c3brbs_reg[24]/NET0131 ,
		\ctl_rf_c3brbs_reg[25]/NET0131 ,
		\ctl_rf_c3brbs_reg[26]/NET0131 ,
		\ctl_rf_c3brbs_reg[27]/NET0131 ,
		_w5604_
	);
	LUT2 #(
		.INIT('h8)
	) name3376 (
		_w5603_,
		_w5604_,
		_w5605_
	);
	LUT2 #(
		.INIT('h4)
	) name3377 (
		_w5602_,
		_w5605_,
		_w5606_
	);
	LUT3 #(
		.INIT('h8c)
	) name3378 (
		\ctl_rf_c4brbs_reg[16]/NET0131 ,
		\ctl_rf_c4brbs_reg[17]/NET0131 ,
		\ctl_rf_c4brbs_reg[22]/NET0131 ,
		_w5607_
	);
	LUT4 #(
		.INIT('h000b)
	) name3379 (
		\ctl_rf_c4brbs_reg[16]/NET0131 ,
		\ctl_rf_c4brbs_reg[20]/NET0131 ,
		\ctl_rf_c4brbs_reg[21]/NET0131 ,
		\ctl_rf_c4brbs_reg[22]/NET0131 ,
		_w5608_
	);
	LUT2 #(
		.INIT('h1)
	) name3380 (
		\ctl_rf_c4brbs_reg[18]/NET0131 ,
		\ctl_rf_c4brbs_reg[19]/NET0131 ,
		_w5609_
	);
	LUT4 #(
		.INIT('hab00)
	) name3381 (
		\ctl_rf_c4brbs_reg[23]/NET0131 ,
		_w5607_,
		_w5608_,
		_w5609_,
		_w5610_
	);
	LUT4 #(
		.INIT('h0001)
	) name3382 (
		\ctl_rf_c4brbs_reg[28]/NET0131 ,
		\ctl_rf_c4brbs_reg[29]/NET0131 ,
		\ctl_rf_c4brbs_reg[30]/NET0131 ,
		\ctl_rf_c4brbs_reg[31]/NET0131 ,
		_w5611_
	);
	LUT4 #(
		.INIT('h0001)
	) name3383 (
		\ctl_rf_c4brbs_reg[24]/NET0131 ,
		\ctl_rf_c4brbs_reg[25]/NET0131 ,
		\ctl_rf_c4brbs_reg[26]/NET0131 ,
		\ctl_rf_c4brbs_reg[27]/NET0131 ,
		_w5612_
	);
	LUT2 #(
		.INIT('h8)
	) name3384 (
		_w5611_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h4)
	) name3385 (
		_w5610_,
		_w5613_,
		_w5614_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3386 (
		_w5602_,
		_w5605_,
		_w5610_,
		_w5613_,
		_w5615_
	);
	LUT3 #(
		.INIT('h20)
	) name3387 (
		_w5590_,
		_w5598_,
		_w5615_,
		_w5616_
	);
	LUT4 #(
		.INIT('h8000)
	) name3388 (
		_w5537_,
		_w5572_,
		_w5573_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('hb)
	) name3389 (
		_w2440_,
		_w5617_,
		_w5618_
	);
	LUT3 #(
		.INIT('h73)
	) name3390 (
		_w2440_,
		_w5477_,
		_w5617_,
		_w5619_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		_w5537_,
		_w5554_,
		_w5620_
	);
	LUT4 #(
		.INIT('h4044)
	) name3392 (
		_w5602_,
		_w5605_,
		_w5610_,
		_w5613_,
		_w5621_
	);
	LUT4 #(
		.INIT('h0800)
	) name3393 (
		_w5571_,
		_w5590_,
		_w5598_,
		_w5621_,
		_w5622_
	);
	LUT3 #(
		.INIT('heb)
	) name3394 (
		_w5581_,
		_w5589_,
		_w5598_,
		_w5623_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		_w5571_,
		_w5615_,
		_w5624_
	);
	LUT4 #(
		.INIT('h4044)
	) name3396 (
		_w5558_,
		_w5561_,
		_w5566_,
		_w5569_,
		_w5625_
	);
	LUT4 #(
		.INIT('h2000)
	) name3397 (
		_w5590_,
		_w5598_,
		_w5615_,
		_w5625_,
		_w5626_
	);
	LUT4 #(
		.INIT('h0045)
	) name3398 (
		_w5622_,
		_w5623_,
		_w5624_,
		_w5626_,
		_w5627_
	);
	LUT3 #(
		.INIT('h80)
	) name3399 (
		_w5494_,
		_w5502_,
		_w5519_,
		_w5628_
	);
	LUT4 #(
		.INIT('h4b44)
	) name3400 (
		_w5506_,
		_w5509_,
		_w5514_,
		_w5517_,
		_w5629_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name3401 (
		_w5494_,
		_w5502_,
		_w5535_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name3402 (
		_w5628_,
		_w5630_,
		_w5631_
	);
	LUT4 #(
		.INIT('h0020)
	) name3403 (
		_w5494_,
		_w5502_,
		_w5519_,
		_w5527_,
		_w5632_
	);
	LUT4 #(
		.INIT('h0302)
	) name3404 (
		_w5536_,
		_w5537_,
		_w5545_,
		_w5632_,
		_w5633_
	);
	LUT4 #(
		.INIT('h2f22)
	) name3405 (
		_w5620_,
		_w5627_,
		_w5631_,
		_w5633_,
		_w5634_
	);
	LUT4 #(
		.INIT('h4000)
	) name3406 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w5635_
	);
	LUT4 #(
		.INIT('h8000)
	) name3407 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w5230_,
		_w5635_,
		_w5636_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3408 (
		\ctl_rf_c1_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5636_,
		_w5637_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3409 (
		\ctl_rf_c1_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5636_,
		_w5638_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3410 (
		\ctl_rf_c1_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5636_,
		_w5639_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3411 (
		\ctl_rf_c1_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5636_,
		_w5640_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3412 (
		\ctl_rf_c1_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5636_,
		_w5641_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3413 (
		\ctl_rf_c1_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5636_,
		_w5642_
	);
	LUT4 #(
		.INIT('h8000)
	) name3414 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w5230_,
		_w5635_,
		_w5643_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3415 (
		\ctl_rf_c1_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5643_,
		_w5644_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3416 (
		\ctl_rf_c1_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5643_,
		_w5645_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3417 (
		\ctl_rf_c1_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5643_,
		_w5646_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3418 (
		\ctl_rf_c1_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5643_,
		_w5647_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3419 (
		\ctl_rf_c1_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5643_,
		_w5648_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3420 (
		\ctl_rf_c1_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5643_,
		_w5649_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3421 (
		\ctl_rf_c1_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5643_,
		_w5650_
	);
	LUT4 #(
		.INIT('h8000)
	) name3422 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w5230_,
		_w5635_,
		_w5651_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name3423 (
		\hwdata[1]_pad ,
		\hwdata[25]_pad ,
		_w2234_,
		_w2235_,
		_w5652_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		\hwdata[9]_pad ,
		_w2234_,
		_w5653_
	);
	LUT4 #(
		.INIT('heee2)
	) name3425 (
		\ctl_rf_c1_rf_chllp_reg[25]/NET0131 ,
		_w5651_,
		_w5652_,
		_w5653_,
		_w5654_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3426 (
		\hwdata[26]_pad ,
		\hwdata[2]_pad ,
		_w2234_,
		_w2235_,
		_w5655_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		\hwdata[10]_pad ,
		_w2234_,
		_w5656_
	);
	LUT4 #(
		.INIT('heee2)
	) name3428 (
		\ctl_rf_c1_rf_chllp_reg[26]/NET0131 ,
		_w5651_,
		_w5655_,
		_w5656_,
		_w5657_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3429 (
		\hwdata[27]_pad ,
		\hwdata[3]_pad ,
		_w2234_,
		_w2235_,
		_w5658_
	);
	LUT2 #(
		.INIT('h8)
	) name3430 (
		\hwdata[11]_pad ,
		_w2234_,
		_w5659_
	);
	LUT4 #(
		.INIT('heee2)
	) name3431 (
		\ctl_rf_c1_rf_chllp_reg[27]/NET0131 ,
		_w5651_,
		_w5658_,
		_w5659_,
		_w5660_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3432 (
		\hwdata[28]_pad ,
		\hwdata[4]_pad ,
		_w2234_,
		_w2235_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name3433 (
		\hwdata[12]_pad ,
		_w2234_,
		_w5662_
	);
	LUT4 #(
		.INIT('heee2)
	) name3434 (
		\ctl_rf_c1_rf_chllp_reg[28]/NET0131 ,
		_w5651_,
		_w5661_,
		_w5662_,
		_w5663_
	);
	LUT4 #(
		.INIT('h8000)
	) name3435 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w5230_,
		_w5635_,
		_w5664_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3436 (
		\ctl_rf_c1_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5664_,
		_w5665_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3437 (
		\ctl_rf_c1_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5664_,
		_w5666_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3438 (
		\ctl_rf_c1_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5664_,
		_w5667_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3439 (
		\ctl_rf_c1_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5664_,
		_w5668_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3440 (
		\ctl_rf_c1_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5636_,
		_w5669_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3441 (
		\ctl_rf_c1_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5636_,
		_w5670_
	);
	LUT4 #(
		.INIT('h8000)
	) name3442 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2244_,
		_w5230_,
		_w5635_,
		_w5671_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3443 (
		\ctl_rf_c3_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5671_,
		_w5672_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3444 (
		\ctl_rf_c3_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5671_,
		_w5673_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3445 (
		\ctl_rf_c3_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5671_,
		_w5674_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3446 (
		\ctl_rf_c3_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5671_,
		_w5675_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3447 (
		\ctl_rf_c3_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5671_,
		_w5676_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3448 (
		\ctl_rf_c3_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5671_,
		_w5677_
	);
	LUT4 #(
		.INIT('h8000)
	) name3449 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2244_,
		_w5230_,
		_w5635_,
		_w5678_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3450 (
		\ctl_rf_c3_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5678_,
		_w5679_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3451 (
		\ctl_rf_c3_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5678_,
		_w5680_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3452 (
		\ctl_rf_c3_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5678_,
		_w5681_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3453 (
		\ctl_rf_c3_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5678_,
		_w5682_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3454 (
		\ctl_rf_c3_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5678_,
		_w5683_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3455 (
		\ctl_rf_c3_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5678_,
		_w5684_
	);
	LUT4 #(
		.INIT('h8000)
	) name3456 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2244_,
		_w5230_,
		_w5635_,
		_w5685_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3457 (
		\ctl_rf_c3_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5685_,
		_w5686_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3458 (
		\ctl_rf_c3_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5685_,
		_w5687_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3459 (
		\ctl_rf_c3_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5685_,
		_w5688_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3460 (
		\ctl_rf_c3_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5685_,
		_w5689_
	);
	LUT4 #(
		.INIT('h8000)
	) name3461 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2244_,
		_w5230_,
		_w5635_,
		_w5690_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3462 (
		\ctl_rf_c3_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5690_,
		_w5691_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3463 (
		\ctl_rf_c3_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5690_,
		_w5692_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3464 (
		\ctl_rf_c3_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5690_,
		_w5693_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3465 (
		\ctl_rf_c3_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5690_,
		_w5694_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3466 (
		\ctl_rf_c3_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5671_,
		_w5695_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3467 (
		\ctl_rf_c3_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5671_,
		_w5696_
	);
	LUT4 #(
		.INIT('h1000)
	) name3468 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w5697_
	);
	LUT4 #(
		.INIT('h8000)
	) name3469 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2247_,
		_w5230_,
		_w5697_,
		_w5698_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3470 (
		\ctl_rf_c4_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3471 (
		\ctl_rf_c4_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5698_,
		_w5700_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3472 (
		\ctl_rf_c4_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5698_,
		_w5701_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3473 (
		\ctl_rf_c4_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5698_,
		_w5702_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3474 (
		\ctl_rf_c4_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5698_,
		_w5703_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3475 (
		\ctl_rf_c4_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5698_,
		_w5704_
	);
	LUT4 #(
		.INIT('h8000)
	) name3476 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2247_,
		_w5230_,
		_w5697_,
		_w5705_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3477 (
		\ctl_rf_c4_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5705_,
		_w5706_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3478 (
		\ctl_rf_c4_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5705_,
		_w5707_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3479 (
		\ctl_rf_c4_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5705_,
		_w5708_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3480 (
		\ctl_rf_c4_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5705_,
		_w5709_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3481 (
		\ctl_rf_c4_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5705_,
		_w5710_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3482 (
		\ctl_rf_c4_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5705_,
		_w5711_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3483 (
		\ctl_rf_c4_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5705_,
		_w5712_
	);
	LUT4 #(
		.INIT('h8000)
	) name3484 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2247_,
		_w5230_,
		_w5697_,
		_w5713_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3485 (
		\ctl_rf_c4_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5713_,
		_w5714_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3486 (
		\ctl_rf_c4_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5713_,
		_w5715_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3487 (
		\ctl_rf_c4_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5713_,
		_w5716_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3488 (
		\ctl_rf_c4_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5713_,
		_w5717_
	);
	LUT4 #(
		.INIT('h8000)
	) name3489 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2247_,
		_w5230_,
		_w5697_,
		_w5718_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3490 (
		\ctl_rf_c4_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5718_,
		_w5719_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3491 (
		\ctl_rf_c4_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5718_,
		_w5720_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3492 (
		\ctl_rf_c4_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5718_,
		_w5721_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3493 (
		\ctl_rf_c4_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5718_,
		_w5722_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3494 (
		\ctl_rf_c4_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5698_,
		_w5723_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3495 (
		\ctl_rf_c4_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5698_,
		_w5724_
	);
	LUT4 #(
		.INIT('h8000)
	) name3496 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2247_,
		_w5230_,
		_w5635_,
		_w5725_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3497 (
		\ctl_rf_c5_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5725_,
		_w5726_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3498 (
		\ctl_rf_c5_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5725_,
		_w5727_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3499 (
		\ctl_rf_c5_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5725_,
		_w5728_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3500 (
		\ctl_rf_c5_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5725_,
		_w5729_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3501 (
		\ctl_rf_c5_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5725_,
		_w5730_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3502 (
		\ctl_rf_c5_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5725_,
		_w5731_
	);
	LUT4 #(
		.INIT('h8000)
	) name3503 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2247_,
		_w5230_,
		_w5635_,
		_w5732_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3504 (
		\ctl_rf_c5_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5732_,
		_w5733_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3505 (
		\ctl_rf_c5_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5732_,
		_w5734_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3506 (
		\ctl_rf_c5_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5732_,
		_w5735_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3507 (
		\ctl_rf_c5_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5732_,
		_w5736_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3508 (
		\ctl_rf_c5_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5732_,
		_w5737_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3509 (
		\ctl_rf_c5_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5732_,
		_w5738_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3510 (
		\ctl_rf_c5_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5732_,
		_w5739_
	);
	LUT4 #(
		.INIT('h8000)
	) name3511 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2247_,
		_w5230_,
		_w5635_,
		_w5740_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3512 (
		\ctl_rf_c5_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5740_,
		_w5741_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3513 (
		\ctl_rf_c5_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5740_,
		_w5742_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3514 (
		\ctl_rf_c5_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5740_,
		_w5743_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3515 (
		\ctl_rf_c5_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5740_,
		_w5744_
	);
	LUT4 #(
		.INIT('h8000)
	) name3516 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2247_,
		_w5230_,
		_w5635_,
		_w5745_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3517 (
		\ctl_rf_c5_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5745_,
		_w5746_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3518 (
		\ctl_rf_c5_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5745_,
		_w5747_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3519 (
		\ctl_rf_c5_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5745_,
		_w5748_
	);
	LUT3 #(
		.INIT('h2a)
	) name3520 (
		\hrdata_reg[17]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5749_
	);
	LUT4 #(
		.INIT('h8000)
	) name3521 (
		_w3503_,
		_w3954_,
		_w3967_,
		_w3980_,
		_w5750_
	);
	LUT3 #(
		.INIT('h54)
	) name3522 (
		_w3424_,
		_w3504_,
		_w5750_,
		_w5751_
	);
	LUT4 #(
		.INIT('hfff5)
	) name3523 (
		\ctl_rf_m0end_reg/NET0131 ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w5752_
	);
	LUT4 #(
		.INIT('hf800)
	) name3524 (
		_w3795_,
		_w3811_,
		_w3837_,
		_w5752_,
		_w5753_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3525 (
		_w3424_,
		_w3484_,
		_w3928_,
		_w3935_,
		_w5754_
	);
	LUT3 #(
		.INIT('h8a)
	) name3526 (
		_w3422_,
		_w3926_,
		_w5754_,
		_w5755_
	);
	LUT4 #(
		.INIT('habaa)
	) name3527 (
		_w5749_,
		_w5751_,
		_w5753_,
		_w5755_,
		_w5756_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3528 (
		\ctl_rf_c5_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5745_,
		_w5757_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3529 (
		\ctl_rf_c5_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5725_,
		_w5758_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3530 (
		\ctl_rf_c5_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5725_,
		_w5759_
	);
	LUT3 #(
		.INIT('h2a)
	) name3531 (
		\hrdata_reg[18]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5760_
	);
	LUT4 #(
		.INIT('h8000)
	) name3532 (
		_w3503_,
		_w4003_,
		_w4016_,
		_w4029_,
		_w5761_
	);
	LUT3 #(
		.INIT('h54)
	) name3533 (
		_w3424_,
		_w3504_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('hf800)
	) name3534 (
		_w4550_,
		_w4566_,
		_w4592_,
		_w5752_,
		_w5763_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3535 (
		_w3424_,
		_w3484_,
		_w4118_,
		_w4124_,
		_w5764_
	);
	LUT3 #(
		.INIT('h8a)
	) name3536 (
		_w3422_,
		_w4117_,
		_w5764_,
		_w5765_
	);
	LUT4 #(
		.INIT('habaa)
	) name3537 (
		_w5760_,
		_w5762_,
		_w5763_,
		_w5765_,
		_w5766_
	);
	LUT4 #(
		.INIT('h1000)
	) name3538 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		_w5767_
	);
	LUT4 #(
		.INIT('h8000)
	) name3539 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2248_,
		_w2254_,
		_w5767_,
		_w5768_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3540 (
		\ctl_rf_c6_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5768_,
		_w5769_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3541 (
		\ctl_rf_c6_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5768_,
		_w5770_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3542 (
		\ctl_rf_c6_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5768_,
		_w5771_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3543 (
		\ctl_rf_c6_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5768_,
		_w5772_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3544 (
		\ctl_rf_c6_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5768_,
		_w5773_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3545 (
		\ctl_rf_c6_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5768_,
		_w5774_
	);
	LUT4 #(
		.INIT('h8000)
	) name3546 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2248_,
		_w2254_,
		_w5767_,
		_w5775_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3547 (
		\ctl_rf_c6_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3548 (
		\ctl_rf_c6_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5775_,
		_w5777_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3549 (
		\ctl_rf_c6_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5775_,
		_w5778_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3550 (
		\ctl_rf_c6_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5775_,
		_w5779_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3551 (
		\ctl_rf_c6_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5775_,
		_w5780_
	);
	LUT4 #(
		.INIT('h8000)
	) name3552 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2248_,
		_w2254_,
		_w5767_,
		_w5781_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3553 (
		\ctl_rf_c6_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3554 (
		\ctl_rf_c6_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5781_,
		_w5783_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3555 (
		\ctl_rf_c6_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5781_,
		_w5784_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3556 (
		\ctl_rf_c6_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5781_,
		_w5785_
	);
	LUT4 #(
		.INIT('h8000)
	) name3557 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2248_,
		_w2254_,
		_w5767_,
		_w5786_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3558 (
		\ctl_rf_c6_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5786_,
		_w5787_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3559 (
		\ctl_rf_c6_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5786_,
		_w5788_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3560 (
		\ctl_rf_c6_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5786_,
		_w5789_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3561 (
		\ctl_rf_c6_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5786_,
		_w5790_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3562 (
		\ctl_rf_c6_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5768_,
		_w5791_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3563 (
		\ctl_rf_c6_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5768_,
		_w5792_
	);
	LUT3 #(
		.INIT('h2a)
	) name3564 (
		\hrdata_reg[19]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5793_
	);
	LUT4 #(
		.INIT('h8000)
	) name3565 (
		_w3503_,
		_w4142_,
		_w4155_,
		_w4168_,
		_w5794_
	);
	LUT3 #(
		.INIT('h54)
	) name3566 (
		_w3424_,
		_w3504_,
		_w5794_,
		_w5795_
	);
	LUT4 #(
		.INIT('hf800)
	) name3567 (
		_w4898_,
		_w4914_,
		_w4940_,
		_w5752_,
		_w5796_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3568 (
		_w3424_,
		_w3484_,
		_w4257_,
		_w4262_,
		_w5797_
	);
	LUT3 #(
		.INIT('h8a)
	) name3569 (
		_w3422_,
		_w4256_,
		_w5797_,
		_w5798_
	);
	LUT4 #(
		.INIT('habaa)
	) name3570 (
		_w5793_,
		_w5795_,
		_w5796_,
		_w5798_,
		_w5799_
	);
	LUT3 #(
		.INIT('h2a)
	) name3571 (
		\hrdata_reg[20]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5800_
	);
	LUT4 #(
		.INIT('h5554)
	) name3572 (
		_w3503_,
		_w4996_,
		_w5007_,
		_w5010_,
		_w5801_
	);
	LUT3 #(
		.INIT('h70)
	) name3573 (
		_w4969_,
		_w4985_,
		_w5801_,
		_w5802_
	);
	LUT4 #(
		.INIT('hc040)
	) name3574 (
		_w3427_,
		_w4280_,
		_w4293_,
		_w4299_,
		_w5803_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		\haddr[8]_pad ,
		_w3503_,
		_w5804_
	);
	LUT3 #(
		.INIT('h45)
	) name3576 (
		_w3424_,
		_w5803_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3577 (
		_w3424_,
		_w3484_,
		_w4389_,
		_w4394_,
		_w5806_
	);
	LUT3 #(
		.INIT('h8a)
	) name3578 (
		_w3422_,
		_w4388_,
		_w5806_,
		_w5807_
	);
	LUT4 #(
		.INIT('hefaa)
	) name3579 (
		_w5800_,
		_w5802_,
		_w5805_,
		_w5807_,
		_w5808_
	);
	LUT3 #(
		.INIT('h2a)
	) name3580 (
		\hrdata_reg[21]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5809_
	);
	LUT4 #(
		.INIT('h5554)
	) name3581 (
		_w3503_,
		_w5066_,
		_w5077_,
		_w5080_,
		_w5810_
	);
	LUT3 #(
		.INIT('h70)
	) name3582 (
		_w5039_,
		_w5055_,
		_w5810_,
		_w5811_
	);
	LUT4 #(
		.INIT('hc040)
	) name3583 (
		_w3427_,
		_w4413_,
		_w4426_,
		_w4432_,
		_w5812_
	);
	LUT3 #(
		.INIT('h51)
	) name3584 (
		_w3424_,
		_w5804_,
		_w5812_,
		_w5813_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3585 (
		_w3424_,
		_w3484_,
		_w4522_,
		_w4527_,
		_w5814_
	);
	LUT3 #(
		.INIT('h8a)
	) name3586 (
		_w3422_,
		_w4521_,
		_w5814_,
		_w5815_
	);
	LUT4 #(
		.INIT('hefaa)
	) name3587 (
		_w5809_,
		_w5811_,
		_w5813_,
		_w5815_,
		_w5816_
	);
	LUT4 #(
		.INIT('h8000)
	) name3588 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2231_,
		_w2254_,
		_w5767_,
		_w5817_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3589 (
		\ctl_rf_c7_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5817_,
		_w5818_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3590 (
		\ctl_rf_c7_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5817_,
		_w5819_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3591 (
		\ctl_rf_c7_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5817_,
		_w5820_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3592 (
		\ctl_rf_c7_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5817_,
		_w5821_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3593 (
		\ctl_rf_c7_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5817_,
		_w5822_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3594 (
		\ctl_rf_c7_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5817_,
		_w5823_
	);
	LUT4 #(
		.INIT('h8000)
	) name3595 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2231_,
		_w2254_,
		_w5767_,
		_w5824_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3596 (
		\ctl_rf_c7_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5824_,
		_w5825_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3597 (
		\ctl_rf_c7_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5824_,
		_w5826_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3598 (
		\ctl_rf_c7_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5824_,
		_w5827_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3599 (
		\ctl_rf_c7_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5824_,
		_w5828_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3600 (
		\ctl_rf_c7_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5824_,
		_w5829_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3601 (
		\ctl_rf_c7_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5824_,
		_w5830_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3602 (
		\ctl_rf_c7_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5824_,
		_w5831_
	);
	LUT4 #(
		.INIT('h8000)
	) name3603 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2231_,
		_w2254_,
		_w5767_,
		_w5832_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3604 (
		\ctl_rf_c7_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5832_,
		_w5833_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3605 (
		\ctl_rf_c7_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5832_,
		_w5834_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3606 (
		\ctl_rf_c7_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5832_,
		_w5835_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3607 (
		\ctl_rf_c7_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5832_,
		_w5836_
	);
	LUT4 #(
		.INIT('h8000)
	) name3608 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2231_,
		_w2254_,
		_w5767_,
		_w5837_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3609 (
		\ctl_rf_c7_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5837_,
		_w5838_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3610 (
		\ctl_rf_c7_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5837_,
		_w5839_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3611 (
		\ctl_rf_c7_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5837_,
		_w5840_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3612 (
		\ctl_rf_c7_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5837_,
		_w5841_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3613 (
		\ctl_rf_c7_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5817_,
		_w5842_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3614 (
		\ctl_rf_c7_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5817_,
		_w5843_
	);
	LUT3 #(
		.INIT('h2a)
	) name3615 (
		\hrdata_reg[22]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5844_
	);
	LUT4 #(
		.INIT('h5554)
	) name3616 (
		_w3503_,
		_w5136_,
		_w5147_,
		_w5150_,
		_w5845_
	);
	LUT3 #(
		.INIT('h70)
	) name3617 (
		_w5109_,
		_w5125_,
		_w5845_,
		_w5846_
	);
	LUT4 #(
		.INIT('hc040)
	) name3618 (
		_w3427_,
		_w4617_,
		_w4630_,
		_w4636_,
		_w5847_
	);
	LUT3 #(
		.INIT('h51)
	) name3619 (
		_w3424_,
		_w5804_,
		_w5847_,
		_w5848_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3620 (
		_w3424_,
		_w3484_,
		_w4726_,
		_w4731_,
		_w5849_
	);
	LUT3 #(
		.INIT('h8a)
	) name3621 (
		_w3422_,
		_w4725_,
		_w5849_,
		_w5850_
	);
	LUT4 #(
		.INIT('hefaa)
	) name3622 (
		_w5844_,
		_w5846_,
		_w5848_,
		_w5850_,
		_w5851_
	);
	LUT3 #(
		.INIT('h2a)
	) name3623 (
		\hrdata_reg[23]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w5852_
	);
	LUT4 #(
		.INIT('h5554)
	) name3624 (
		_w3503_,
		_w5206_,
		_w5217_,
		_w5220_,
		_w5853_
	);
	LUT3 #(
		.INIT('h70)
	) name3625 (
		_w5179_,
		_w5195_,
		_w5853_,
		_w5854_
	);
	LUT4 #(
		.INIT('hc040)
	) name3626 (
		_w3427_,
		_w4750_,
		_w4763_,
		_w4769_,
		_w5855_
	);
	LUT3 #(
		.INIT('h51)
	) name3627 (
		_w3424_,
		_w5804_,
		_w5855_,
		_w5856_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3628 (
		_w3424_,
		_w3484_,
		_w4870_,
		_w4875_,
		_w5857_
	);
	LUT3 #(
		.INIT('h8a)
	) name3629 (
		_w3422_,
		_w4869_,
		_w5857_,
		_w5858_
	);
	LUT4 #(
		.INIT('hefaa)
	) name3630 (
		_w5852_,
		_w5854_,
		_w5856_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('he)
	) name3631 (
		_w2431_,
		_w5617_,
		_w5860_
	);
	LUT4 #(
		.INIT('h8000)
	) name3632 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w5230_,
		_w5697_,
		_w5861_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3633 (
		\ctl_rf_c0_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5861_,
		_w5862_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3634 (
		\ctl_rf_c0_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5861_,
		_w5863_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3635 (
		\ctl_rf_c0_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5861_,
		_w5864_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3636 (
		\ctl_rf_c0_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5861_,
		_w5865_
	);
	LUT4 #(
		.INIT('h8000)
	) name3637 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w5230_,
		_w5697_,
		_w5866_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3638 (
		\ctl_rf_c0_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h8000)
	) name3639 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w5230_,
		_w5697_,
		_w5868_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3640 (
		\ctl_rf_c0_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5868_,
		_w5869_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3641 (
		\ctl_rf_c0_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5868_,
		_w5870_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3642 (
		\ctl_rf_c0_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5868_,
		_w5871_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3643 (
		\ctl_rf_c0_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5861_,
		_w5872_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3644 (
		\ctl_rf_c0_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5861_,
		_w5873_
	);
	LUT4 #(
		.INIT('h8000)
	) name3645 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2244_,
		_w5230_,
		_w5697_,
		_w5874_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3646 (
		\ctl_rf_c2_rf_chllp_reg[10]/NET0131 ,
		_w5289_,
		_w5290_,
		_w5874_,
		_w5875_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3647 (
		\ctl_rf_c2_rf_chllp_reg[11]/NET0131 ,
		_w5300_,
		_w5301_,
		_w5874_,
		_w5876_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3648 (
		\ctl_rf_c2_rf_chllp_reg[12]/NET0131 ,
		_w5292_,
		_w5293_,
		_w5874_,
		_w5877_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3649 (
		\ctl_rf_c2_rf_chllp_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5874_,
		_w5878_
	);
	LUT4 #(
		.INIT('h8000)
	) name3650 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2244_,
		_w5230_,
		_w5697_,
		_w5879_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3651 (
		\ctl_rf_c2_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3652 (
		\ctl_rf_c2_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5879_,
		_w5881_
	);
	LUT4 #(
		.INIT('h8000)
	) name3653 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2244_,
		_w5230_,
		_w5697_,
		_w5882_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3654 (
		\ctl_rf_c2_rf_chllp_reg[28]/NET0131 ,
		_w5661_,
		_w5662_,
		_w5882_,
		_w5883_
	);
	LUT4 #(
		.INIT('h8000)
	) name3655 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2244_,
		_w5230_,
		_w5697_,
		_w5884_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3656 (
		\ctl_rf_c2_rf_chllp_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5884_,
		_w5885_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3657 (
		\ctl_rf_c2_rf_chllp_reg[6]/NET0131 ,
		_w5236_,
		_w5237_,
		_w5884_,
		_w5886_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3658 (
		\ctl_rf_c2_rf_chllp_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5884_,
		_w5887_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3659 (
		\ctl_rf_c2_rf_chllp_reg[8]/NET0131 ,
		_w5296_,
		_w5297_,
		_w5874_,
		_w5888_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3660 (
		\ctl_rf_c2_rf_chllp_reg[9]/NET0131 ,
		_w5305_,
		_w5306_,
		_w5874_,
		_w5889_
	);
	LUT4 #(
		.INIT('h0400)
	) name3661 (
		_w5577_,
		_w5580_,
		_w5585_,
		_w5588_,
		_w5890_
	);
	LUT4 #(
		.INIT('h0600)
	) name3662 (
		_w5581_,
		_w5589_,
		_w5598_,
		_w5615_,
		_w5891_
	);
	LUT4 #(
		.INIT('h5155)
	) name3663 (
		_w5570_,
		_w5590_,
		_w5598_,
		_w5621_,
		_w5892_
	);
	LUT2 #(
		.INIT('h4)
	) name3664 (
		_w5891_,
		_w5892_,
		_w5893_
	);
	LUT4 #(
		.INIT('h0400)
	) name3665 (
		_w5562_,
		_w5590_,
		_w5598_,
		_w5615_,
		_w5894_
	);
	LUT4 #(
		.INIT('h8880)
	) name3666 (
		_w5537_,
		_w5554_,
		_w5571_,
		_w5894_,
		_w5895_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3667 (
		_w5481_,
		_w5484_,
		_w5506_,
		_w5509_,
		_w5896_
	);
	LUT4 #(
		.INIT('h0400)
	) name3668 (
		_w5489_,
		_w5492_,
		_w5514_,
		_w5517_,
		_w5897_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3669 (
		_w5489_,
		_w5492_,
		_w5514_,
		_w5517_,
		_w5898_
	);
	LUT4 #(
		.INIT('h1200)
	) name3670 (
		_w5493_,
		_w5502_,
		_w5518_,
		_w5896_,
		_w5899_
	);
	LUT4 #(
		.INIT('h007f)
	) name3671 (
		_w5494_,
		_w5502_,
		_w5519_,
		_w5527_,
		_w5900_
	);
	LUT2 #(
		.INIT('h4)
	) name3672 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT4 #(
		.INIT('h0020)
	) name3673 (
		_w5494_,
		_w5502_,
		_w5519_,
		_w5535_,
		_w5902_
	);
	LUT4 #(
		.INIT('h0302)
	) name3674 (
		_w5536_,
		_w5537_,
		_w5545_,
		_w5902_,
		_w5903_
	);
	LUT4 #(
		.INIT('h4f44)
	) name3675 (
		_w5893_,
		_w5895_,
		_w5901_,
		_w5903_,
		_w5904_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3676 (
		\ctl_rf_c0_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5861_,
		_w5905_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3677 (
		\ctl_rf_c0_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5861_,
		_w5906_
	);
	LUT4 #(
		.INIT('h8000)
	) name3678 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w5230_,
		_w5697_,
		_w5907_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3679 (
		\ctl_rf_c0_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5907_,
		_w5908_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3680 (
		\ctl_rf_c0_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5907_,
		_w5909_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3681 (
		\ctl_rf_c0_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5866_,
		_w5910_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3682 (
		\ctl_rf_c0_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5866_,
		_w5911_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3683 (
		\ctl_rf_c0_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5866_,
		_w5912_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3684 (
		\ctl_rf_c0_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5868_,
		_w5913_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3685 (
		\ctl_rf_c1_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5643_,
		_w5914_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3686 (
		\ctl_rf_c1_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5651_,
		_w5915_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3687 (
		\hwdata[29]_pad ,
		\hwdata[5]_pad ,
		_w2234_,
		_w2235_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name3688 (
		\hwdata[13]_pad ,
		_w2234_,
		_w5917_
	);
	LUT4 #(
		.INIT('heee2)
	) name3689 (
		\ctl_rf_c1_rf_chllp_reg[29]/NET0131 ,
		_w5651_,
		_w5916_,
		_w5917_,
		_w5918_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3690 (
		\ctl_rf_c1_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5664_,
		_w5919_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name3691 (
		\hwdata[30]_pad ,
		\hwdata[6]_pad ,
		_w2234_,
		_w2235_,
		_w5920_
	);
	LUT2 #(
		.INIT('h8)
	) name3692 (
		\hwdata[14]_pad ,
		_w2234_,
		_w5921_
	);
	LUT4 #(
		.INIT('heee2)
	) name3693 (
		\ctl_rf_c1_rf_chllp_reg[30]/NET0131 ,
		_w5651_,
		_w5920_,
		_w5921_,
		_w5922_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3694 (
		\ctl_rf_c1_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5651_,
		_w5923_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3695 (
		\ctl_rf_c1_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5664_,
		_w5924_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3696 (
		\ctl_rf_c2_rf_chllp_reg[13]/NET0131 ,
		_w5367_,
		_w5368_,
		_w5874_,
		_w5925_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3697 (
		\ctl_rf_c2_rf_chllp_reg[14]/NET0131 ,
		_w5370_,
		_w5371_,
		_w5874_,
		_w5926_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3698 (
		\ctl_rf_c2_rf_chllp_reg[16]/NET0131 ,
		_w2371_,
		_w2372_,
		_w5879_,
		_w5927_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3699 (
		\ctl_rf_c2_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5879_,
		_w5928_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3700 (
		\ctl_rf_c2_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5879_,
		_w5929_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3701 (
		\ctl_rf_c2_rf_chllp_reg[19]/NET0131 ,
		_w2298_,
		_w2299_,
		_w5879_,
		_w5930_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3702 (
		\ctl_rf_c2_rf_chllp_reg[25]/NET0131 ,
		_w5652_,
		_w5653_,
		_w5882_,
		_w5931_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3703 (
		\ctl_rf_c2_rf_chllp_reg[26]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5882_,
		_w5932_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3704 (
		\ctl_rf_c2_rf_chllp_reg[27]/NET0131 ,
		_w5658_,
		_w5659_,
		_w5882_,
		_w5933_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3705 (
		\ctl_rf_c2_rf_chllp_reg[4]/NET0131 ,
		_w5275_,
		_w5276_,
		_w5884_,
		_w5934_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3706 (
		\ctl_rf_c3_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5678_,
		_w5935_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3707 (
		\ctl_rf_c3_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5685_,
		_w5936_
	);
	LUT4 #(
		.INIT('heee2)
	) name3708 (
		\ctl_rf_c3_rf_chllp_reg[29]/NET0131 ,
		_w5685_,
		_w5916_,
		_w5917_,
		_w5937_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3709 (
		\ctl_rf_c3_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5690_,
		_w5938_
	);
	LUT4 #(
		.INIT('heee2)
	) name3710 (
		\ctl_rf_c3_rf_chllp_reg[30]/NET0131 ,
		_w5685_,
		_w5920_,
		_w5921_,
		_w5939_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3711 (
		\ctl_rf_c3_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5685_,
		_w5940_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3712 (
		\ctl_rf_c3_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5690_,
		_w5941_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3713 (
		\ctl_rf_c4_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5705_,
		_w5942_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3714 (
		\ctl_rf_c4_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5713_,
		_w5943_
	);
	LUT4 #(
		.INIT('heee2)
	) name3715 (
		\ctl_rf_c4_rf_chllp_reg[29]/NET0131 ,
		_w5713_,
		_w5916_,
		_w5917_,
		_w5944_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3716 (
		\ctl_rf_c4_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5718_,
		_w5945_
	);
	LUT4 #(
		.INIT('heee2)
	) name3717 (
		\ctl_rf_c4_rf_chllp_reg[30]/NET0131 ,
		_w5713_,
		_w5920_,
		_w5921_,
		_w5946_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3718 (
		\ctl_rf_c4_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5713_,
		_w5947_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3719 (
		\ctl_rf_c4_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5718_,
		_w5948_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3720 (
		\ctl_rf_c5_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5732_,
		_w5949_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3721 (
		\ctl_rf_c5_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5740_,
		_w5950_
	);
	LUT4 #(
		.INIT('heee2)
	) name3722 (
		\ctl_rf_c5_rf_chllp_reg[29]/NET0131 ,
		_w5740_,
		_w5916_,
		_w5917_,
		_w5951_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3723 (
		\ctl_rf_c5_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5745_,
		_w5952_
	);
	LUT4 #(
		.INIT('heee2)
	) name3724 (
		\ctl_rf_c5_rf_chllp_reg[30]/NET0131 ,
		_w5740_,
		_w5920_,
		_w5921_,
		_w5953_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3725 (
		\ctl_rf_c5_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5740_,
		_w5954_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3726 (
		\ctl_rf_c5_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5745_,
		_w5955_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3727 (
		\ctl_rf_c6_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5775_,
		_w5956_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3728 (
		\ctl_rf_c6_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5781_,
		_w5957_
	);
	LUT4 #(
		.INIT('heee2)
	) name3729 (
		\ctl_rf_c6_rf_chllp_reg[29]/NET0131 ,
		_w5781_,
		_w5916_,
		_w5917_,
		_w5958_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3730 (
		\ctl_rf_c6_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5786_,
		_w5959_
	);
	LUT4 #(
		.INIT('heee2)
	) name3731 (
		\ctl_rf_c6_rf_chllp_reg[30]/NET0131 ,
		_w5781_,
		_w5920_,
		_w5921_,
		_w5960_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3732 (
		\ctl_rf_c6_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5781_,
		_w5961_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3733 (
		\ctl_rf_c6_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5786_,
		_w5962_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3734 (
		\ctl_rf_c7_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5824_,
		_w5963_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3735 (
		\ctl_rf_c7_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5832_,
		_w5964_
	);
	LUT4 #(
		.INIT('heee2)
	) name3736 (
		\ctl_rf_c7_rf_chllp_reg[29]/NET0131 ,
		_w5832_,
		_w5916_,
		_w5917_,
		_w5965_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3737 (
		\ctl_rf_c7_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5837_,
		_w5966_
	);
	LUT4 #(
		.INIT('heee2)
	) name3738 (
		\ctl_rf_c7_rf_chllp_reg[30]/NET0131 ,
		_w5832_,
		_w5920_,
		_w5921_,
		_w5967_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3739 (
		\ctl_rf_c7_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5832_,
		_w5968_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3740 (
		\ctl_rf_c7_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5837_,
		_w5969_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3741 (
		\ctl_rf_c0_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5907_,
		_w5970_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3742 (
		\ctl_rf_c2_rf_chllp_reg[23]/NET0131 ,
		_w2331_,
		_w2332_,
		_w5879_,
		_w5971_
	);
	LUT2 #(
		.INIT('h8)
	) name3743 (
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w5972_
	);
	LUT3 #(
		.INIT('h80)
	) name3744 (
		\ch_sel_arb_chcsr_reg_reg[17]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w5973_
	);
	LUT2 #(
		.INIT('h8)
	) name3745 (
		\ch_sel_arb_chcsr_reg_reg[15]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[16]/NET0131 ,
		_w5974_
	);
	LUT3 #(
		.INIT('h2a)
	) name3746 (
		\de_bst_cnt_reg[8]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w5975_
	);
	LUT3 #(
		.INIT('hf8)
	) name3747 (
		_w5973_,
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3748 (
		\ctl_rf_c0_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5907_,
		_w5977_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3749 (
		\ctl_rf_c0_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5866_,
		_w5978_
	);
	LUT4 #(
		.INIT('heee2)
	) name3750 (
		\ctl_rf_c0_rf_chllp_reg[29]/NET0131 ,
		_w5866_,
		_w5916_,
		_w5917_,
		_w5979_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3751 (
		\ctl_rf_c0_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5868_,
		_w5980_
	);
	LUT4 #(
		.INIT('heee2)
	) name3752 (
		\ctl_rf_c0_rf_chllp_reg[30]/NET0131 ,
		_w5866_,
		_w5920_,
		_w5921_,
		_w5981_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3753 (
		\ctl_rf_c0_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5866_,
		_w5982_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3754 (
		\ctl_rf_c0_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5868_,
		_w5983_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3755 (
		\ctl_rf_c2_rf_chllp_reg[20]/NET0131 ,
		_w2341_,
		_w2342_,
		_w5879_,
		_w5984_
	);
	LUT4 #(
		.INIT('heee2)
	) name3756 (
		\ctl_rf_c2_rf_chllp_reg[29]/NET0131 ,
		_w5882_,
		_w5916_,
		_w5917_,
		_w5985_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3757 (
		\ctl_rf_c2_rf_chllp_reg[2]/NET0131 ,
		_w5362_,
		_w5363_,
		_w5884_,
		_w5986_
	);
	LUT4 #(
		.INIT('heee2)
	) name3758 (
		\ctl_rf_c2_rf_chllp_reg[30]/NET0131 ,
		_w5882_,
		_w5920_,
		_w5921_,
		_w5987_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3759 (
		\ctl_rf_c2_rf_chllp_reg[31]/NET0131 ,
		_w2260_,
		_w2261_,
		_w5882_,
		_w5988_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name3760 (
		\ctl_rf_c2_rf_chllp_reg[3]/NET0131 ,
		_w5375_,
		_w5376_,
		_w5884_,
		_w5989_
	);
	LUT4 #(
		.INIT('hc884)
	) name3761 (
		\de_m1_is_llp_reg/NET0131 ,
		\h1size[1]_pad ,
		_w2425_,
		_w2834_,
		_w5990_
	);
	LUT4 #(
		.INIT('h8880)
	) name3762 (
		\ch_sel_arb_chcsr_reg_reg[12]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w5991_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		_w2835_,
		_w5991_,
		_w5992_
	);
	LUT4 #(
		.INIT('h0080)
	) name3764 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[9]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w5993_
	);
	LUT3 #(
		.INIT('hab)
	) name3765 (
		_w2425_,
		_w2836_,
		_w5993_,
		_w5994_
	);
	LUT4 #(
		.INIT('h5455)
	) name3766 (
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w5990_,
		_w5992_,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h8)
	) name3767 (
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w5996_
	);
	LUT2 #(
		.INIT('he)
	) name3768 (
		_w5995_,
		_w5996_,
		_w5997_
	);
	LUT4 #(
		.INIT('hff10)
	) name3769 (
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w5998_
	);
	LUT4 #(
		.INIT('h0706)
	) name3770 (
		_w5590_,
		_w5598_,
		_w5614_,
		_w5890_,
		_w5999_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3771 (
		_w5594_,
		_w5597_,
		_w5602_,
		_w5605_,
		_w6000_
	);
	LUT3 #(
		.INIT('h13)
	) name3772 (
		_w5590_,
		_w5615_,
		_w6000_,
		_w6001_
	);
	LUT4 #(
		.INIT('h0008)
	) name3773 (
		_w5537_,
		_w5572_,
		_w5999_,
		_w6001_,
		_w6002_
	);
	LUT4 #(
		.INIT('h99fe)
	) name3774 (
		_w5485_,
		_w5510_,
		_w5897_,
		_w5898_,
		_w6003_
	);
	LUT3 #(
		.INIT('h04)
	) name3775 (
		_w5502_,
		_w5536_,
		_w5545_,
		_w6004_
	);
	LUT3 #(
		.INIT('h10)
	) name3776 (
		_w5537_,
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('he)
	) name3777 (
		_w6002_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h2)
	) name3778 (
		\de_de_st_reg[5]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6007_
	);
	LUT3 #(
		.INIT('h8a)
	) name3779 (
		\de_m1_arb_st_reg[0]/NET0131 ,
		_w2418_,
		_w6007_,
		_w6008_
	);
	LUT3 #(
		.INIT('h40)
	) name3780 (
		_w2418_,
		_w2467_,
		_w3400_,
		_w6009_
	);
	LUT2 #(
		.INIT('he)
	) name3781 (
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT3 #(
		.INIT('h2a)
	) name3782 (
		\hrdata_reg[10]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6011_
	);
	LUT4 #(
		.INIT('h4000)
	) name3783 (
		_w3503_,
		_w4003_,
		_w4016_,
		_w4029_,
		_w6012_
	);
	LUT3 #(
		.INIT('h54)
	) name3784 (
		_w3424_,
		_w3682_,
		_w6012_,
		_w6013_
	);
	LUT4 #(
		.INIT('hf800)
	) name3785 (
		_w4550_,
		_w4566_,
		_w4592_,
		_w3503_,
		_w6014_
	);
	LUT3 #(
		.INIT('h20)
	) name3786 (
		_w3424_,
		_w4042_,
		_w4053_,
		_w6015_
	);
	LUT3 #(
		.INIT('ha2)
	) name3787 (
		_w3424_,
		_w3427_,
		_w4075_,
		_w6016_
	);
	LUT4 #(
		.INIT('h020a)
	) name3788 (
		_w3422_,
		_w4070_,
		_w6015_,
		_w6016_,
		_w6017_
	);
	LUT4 #(
		.INIT('habaa)
	) name3789 (
		_w6011_,
		_w6013_,
		_w6014_,
		_w6017_,
		_w6018_
	);
	LUT3 #(
		.INIT('h2a)
	) name3790 (
		\hrdata_reg[11]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6019_
	);
	LUT4 #(
		.INIT('h4000)
	) name3791 (
		_w3503_,
		_w4142_,
		_w4155_,
		_w4168_,
		_w6020_
	);
	LUT3 #(
		.INIT('h54)
	) name3792 (
		_w3424_,
		_w3682_,
		_w6020_,
		_w6021_
	);
	LUT4 #(
		.INIT('hf800)
	) name3793 (
		_w4898_,
		_w4914_,
		_w4940_,
		_w3503_,
		_w6022_
	);
	LUT3 #(
		.INIT('h20)
	) name3794 (
		_w3424_,
		_w4181_,
		_w4192_,
		_w6023_
	);
	LUT3 #(
		.INIT('ha2)
	) name3795 (
		_w3424_,
		_w3427_,
		_w4214_,
		_w6024_
	);
	LUT4 #(
		.INIT('h020a)
	) name3796 (
		_w3422_,
		_w4209_,
		_w6023_,
		_w6024_,
		_w6025_
	);
	LUT4 #(
		.INIT('habaa)
	) name3797 (
		_w6019_,
		_w6021_,
		_w6022_,
		_w6025_,
		_w6026_
	);
	LUT3 #(
		.INIT('h2a)
	) name3798 (
		\hrdata_reg[12]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6027_
	);
	LUT3 #(
		.INIT('h20)
	) name3799 (
		_w3424_,
		_w4313_,
		_w4324_,
		_w6028_
	);
	LUT3 #(
		.INIT('ha2)
	) name3800 (
		_w3424_,
		_w3427_,
		_w4346_,
		_w6029_
	);
	LUT4 #(
		.INIT('h020a)
	) name3801 (
		_w3422_,
		_w4341_,
		_w6028_,
		_w6029_,
		_w6030_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3802 (
		_w3503_,
		_w4996_,
		_w5007_,
		_w5010_,
		_w6031_
	);
	LUT4 #(
		.INIT('h4055)
	) name3803 (
		_w3424_,
		_w4969_,
		_w4985_,
		_w6031_,
		_w6032_
	);
	LUT2 #(
		.INIT('h2)
	) name3804 (
		\haddr[8]_pad ,
		_w3503_,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		_w5803_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('heeae)
	) name3806 (
		_w6027_,
		_w6030_,
		_w6032_,
		_w6034_,
		_w6035_
	);
	LUT3 #(
		.INIT('h2a)
	) name3807 (
		\hrdata_reg[13]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6036_
	);
	LUT3 #(
		.INIT('h20)
	) name3808 (
		_w3424_,
		_w4446_,
		_w4457_,
		_w6037_
	);
	LUT3 #(
		.INIT('ha2)
	) name3809 (
		_w3424_,
		_w3427_,
		_w4479_,
		_w6038_
	);
	LUT4 #(
		.INIT('h020a)
	) name3810 (
		_w3422_,
		_w4474_,
		_w6037_,
		_w6038_,
		_w6039_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3811 (
		_w3503_,
		_w5066_,
		_w5077_,
		_w5080_,
		_w6040_
	);
	LUT4 #(
		.INIT('h4055)
	) name3812 (
		_w3424_,
		_w5039_,
		_w5055_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h4)
	) name3813 (
		_w5812_,
		_w6033_,
		_w6042_
	);
	LUT4 #(
		.INIT('heeae)
	) name3814 (
		_w6036_,
		_w6039_,
		_w6041_,
		_w6042_,
		_w6043_
	);
	LUT3 #(
		.INIT('h2a)
	) name3815 (
		\hrdata_reg[14]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6044_
	);
	LUT3 #(
		.INIT('h20)
	) name3816 (
		_w3424_,
		_w4650_,
		_w4661_,
		_w6045_
	);
	LUT3 #(
		.INIT('ha2)
	) name3817 (
		_w3424_,
		_w3427_,
		_w4683_,
		_w6046_
	);
	LUT4 #(
		.INIT('h020a)
	) name3818 (
		_w3422_,
		_w4678_,
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3819 (
		_w3503_,
		_w5136_,
		_w5147_,
		_w5150_,
		_w6048_
	);
	LUT4 #(
		.INIT('h4055)
	) name3820 (
		_w3424_,
		_w5109_,
		_w5125_,
		_w6048_,
		_w6049_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w5847_,
		_w6033_,
		_w6050_
	);
	LUT4 #(
		.INIT('heeae)
	) name3822 (
		_w6044_,
		_w6047_,
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT3 #(
		.INIT('h2a)
	) name3823 (
		\hrdata_reg[15]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6052_
	);
	LUT3 #(
		.INIT('h8a)
	) name3824 (
		_w3422_,
		_w4816_,
		_w4827_,
		_w6053_
	);
	LUT4 #(
		.INIT('h4055)
	) name3825 (
		_w3622_,
		_w4789_,
		_w4805_,
		_w6053_,
		_w6054_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3826 (
		_w3503_,
		_w5206_,
		_w5217_,
		_w5220_,
		_w6055_
	);
	LUT4 #(
		.INIT('h4055)
	) name3827 (
		_w3424_,
		_w5179_,
		_w5195_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h4)
	) name3828 (
		_w5855_,
		_w6033_,
		_w6057_
	);
	LUT4 #(
		.INIT('hbbab)
	) name3829 (
		_w6052_,
		_w6054_,
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('h2a)
	) name3830 (
		\hrdata_reg[9]_pad ,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w6059_
	);
	LUT4 #(
		.INIT('h4000)
	) name3831 (
		_w3503_,
		_w3954_,
		_w3967_,
		_w3980_,
		_w6060_
	);
	LUT3 #(
		.INIT('h54)
	) name3832 (
		_w3424_,
		_w3682_,
		_w6060_,
		_w6061_
	);
	LUT4 #(
		.INIT('hf800)
	) name3833 (
		_w3795_,
		_w3811_,
		_w3837_,
		_w3503_,
		_w6062_
	);
	LUT3 #(
		.INIT('h20)
	) name3834 (
		_w3424_,
		_w3851_,
		_w3862_,
		_w6063_
	);
	LUT3 #(
		.INIT('ha2)
	) name3835 (
		_w3424_,
		_w3427_,
		_w3884_,
		_w6064_
	);
	LUT4 #(
		.INIT('h020a)
	) name3836 (
		_w3422_,
		_w3879_,
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT4 #(
		.INIT('habaa)
	) name3837 (
		_w6059_,
		_w6061_,
		_w6062_,
		_w6065_,
		_w6066_
	);
	LUT4 #(
		.INIT('hc884)
	) name3838 (
		\de_m1_is_llp_reg/NET0131 ,
		\h1size[0]_pad ,
		_w2425_,
		_w2834_,
		_w6067_
	);
	LUT4 #(
		.INIT('h0080)
	) name3839 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[8]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w6068_
	);
	LUT4 #(
		.INIT('h8880)
	) name3840 (
		\ch_sel_arb_chcsr_reg_reg[11]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w6069_
	);
	LUT4 #(
		.INIT('h23af)
	) name3841 (
		_w2425_,
		_w2835_,
		_w6068_,
		_w6069_,
		_w6070_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name3842 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6067_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		_w6072_
	);
	LUT3 #(
		.INIT('h0d)
	) name3844 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w6073_
	);
	LUT4 #(
		.INIT('ha882)
	) name3845 (
		\ahb_mst0_hsizeo_reg[1]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w2484_,
		_w6072_,
		_w6074_
	);
	LUT4 #(
		.INIT('h0020)
	) name3846 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[9]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w6075_
	);
	LUT2 #(
		.INIT('h4)
	) name3847 (
		_w2484_,
		_w6075_,
		_w6076_
	);
	LUT4 #(
		.INIT('h2220)
	) name3848 (
		\ch_sel_arb_chcsr_reg_reg[12]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w6077_
	);
	LUT4 #(
		.INIT('hf8fd)
	) name3849 (
		\de_m0_is_llp_reg/NET0131 ,
		_w2484_,
		_w6072_,
		_w6077_,
		_w6078_
	);
	LUT3 #(
		.INIT('hef)
	) name3850 (
		_w6074_,
		_w6076_,
		_w6078_,
		_w6079_
	);
	LUT3 #(
		.INIT('h20)
	) name3851 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6080_
	);
	LUT4 #(
		.INIT('h8000)
	) name3852 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		_w2390_,
		_w2393_,
		_w2396_,
		_w6081_
	);
	LUT4 #(
		.INIT('h070f)
	) name3853 (
		_w2403_,
		_w2416_,
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT4 #(
		.INIT('h0800)
	) name3854 (
		hreadyin_pad,
		hsel_br_pad,
		\htrans[0]_pad ,
		\htrans[1]_pad ,
		_w6083_
	);
	LUT4 #(
		.INIT('h1001)
	) name3855 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		hreadyout_br_pad,
		\hresp_br[0]_pad ,
		\hresp_br[1]_pad ,
		_w6084_
	);
	LUT4 #(
		.INIT('h8000)
	) name3856 (
		hreadyout_br_pad,
		hsel_br_pad,
		\htrans[0]_pad ,
		\htrans[1]_pad ,
		_w6085_
	);
	LUT4 #(
		.INIT('h0001)
	) name3857 (
		\ahb_slv_br_st_reg[1]/NET0131 ,
		_w6083_,
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h8)
	) name3858 (
		_w6082_,
		_w6086_,
		_w6087_
	);
	LUT3 #(
		.INIT('h40)
	) name3859 (
		\ch_sel_arb_chcsr_reg_reg[17]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6088_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		\ch_sel_arb_chcsr_reg_reg[15]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[16]/NET0131 ,
		_w6089_
	);
	LUT3 #(
		.INIT('h2a)
	) name3861 (
		\de_bst_cnt_reg[0]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6090_
	);
	LUT3 #(
		.INIT('hf8)
	) name3862 (
		_w6088_,
		_w6089_,
		_w6090_,
		_w6091_
	);
	LUT3 #(
		.INIT('h2a)
	) name3863 (
		\de_bst_cnt_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name3864 (
		\ch_sel_arb_chcsr_reg_reg[15]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[16]/NET0131 ,
		_w6093_
	);
	LUT3 #(
		.INIT('hec)
	) name3865 (
		_w6088_,
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT3 #(
		.INIT('h2a)
	) name3866 (
		\de_bst_cnt_reg[3]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6095_
	);
	LUT2 #(
		.INIT('h4)
	) name3867 (
		\ch_sel_arb_chcsr_reg_reg[15]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[16]/NET0131 ,
		_w6096_
	);
	LUT3 #(
		.INIT('hec)
	) name3868 (
		_w6088_,
		_w6095_,
		_w6096_,
		_w6097_
	);
	LUT3 #(
		.INIT('h2a)
	) name3869 (
		\de_bst_cnt_reg[4]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6098_
	);
	LUT3 #(
		.INIT('hf8)
	) name3870 (
		_w5974_,
		_w6088_,
		_w6098_,
		_w6099_
	);
	LUT3 #(
		.INIT('h2a)
	) name3871 (
		\de_bst_cnt_reg[5]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6100_
	);
	LUT3 #(
		.INIT('hf8)
	) name3872 (
		_w5973_,
		_w6089_,
		_w6100_,
		_w6101_
	);
	LUT3 #(
		.INIT('h2a)
	) name3873 (
		\de_bst_cnt_reg[7]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6102_
	);
	LUT3 #(
		.INIT('hf8)
	) name3874 (
		_w5973_,
		_w6096_,
		_w6102_,
		_w6103_
	);
	LUT3 #(
		.INIT('h2a)
	) name3875 (
		\de_bst_cnt_reg[6]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w6104_
	);
	LUT3 #(
		.INIT('hf8)
	) name3876 (
		_w5973_,
		_w6093_,
		_w6104_,
		_w6105_
	);
	LUT4 #(
		.INIT('ha882)
	) name3877 (
		\ahb_mst0_hsizeo_reg[0]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w2484_,
		_w6072_,
		_w6106_
	);
	LUT4 #(
		.INIT('h0020)
	) name3878 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[8]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w6107_
	);
	LUT4 #(
		.INIT('h2220)
	) name3879 (
		\ch_sel_arb_chcsr_reg_reg[11]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w6108_
	);
	LUT4 #(
		.INIT('h23af)
	) name3880 (
		_w2484_,
		_w6073_,
		_w6107_,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('hb)
	) name3881 (
		_w6106_,
		_w6109_,
		_w6110_
	);
	LUT4 #(
		.INIT('ha882)
	) name3882 (
		\ahb_mst0_hsizeo_reg[2]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w2484_,
		_w6072_,
		_w6111_
	);
	LUT4 #(
		.INIT('h2220)
	) name3883 (
		\ch_sel_arb_chcsr_reg_reg[13]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[2]/NET0131 ,
		_w6112_
	);
	LUT4 #(
		.INIT('h0008)
	) name3884 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[10]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w6113_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name3885 (
		_w2484_,
		_w6073_,
		_w6112_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('hb)
	) name3886 (
		_w6111_,
		_w6114_,
		_w6115_
	);
	LUT2 #(
		.INIT('h8)
	) name3887 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w6116_
	);
	LUT3 #(
		.INIT('h13)
	) name3888 (
		\de_de_st_reg[6]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w6117_
	);
	LUT3 #(
		.INIT('h45)
	) name3889 (
		_w2431_,
		_w6116_,
		_w6117_,
		_w6118_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3890 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6120_
	);
	LUT4 #(
		.INIT('h0008)
	) name3892 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6121_
	);
	LUT3 #(
		.INIT('h54)
	) name3893 (
		_w2431_,
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3894 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w6122_,
		_w6123_
	);
	LUT3 #(
		.INIT('hf2)
	) name3895 (
		\h1write_pad ,
		_w6119_,
		_w6123_,
		_w6124_
	);
	LUT3 #(
		.INIT('hac)
	) name3896 (
		\ahb_slv_slv_pt_d1o_reg[2]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[19]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6125_
	);
	LUT3 #(
		.INIT('hac)
	) name3897 (
		\ahb_slv_slv_pt_d1o_reg[3]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[20]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6126_
	);
	LUT3 #(
		.INIT('hac)
	) name3898 (
		\ahb_slv_slv_pt_d1o_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[18]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6127_
	);
	LUT2 #(
		.INIT('he)
	) name3899 (
		_w2993_,
		_w2994_,
		_w6128_
	);
	LUT4 #(
		.INIT('h8000)
	) name3900 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2230_,
		_w3112_,
		_w6129_
	);
	LUT3 #(
		.INIT('he0)
	) name3901 (
		_w2993_,
		_w2994_,
		_w6129_,
		_w6130_
	);
	LUT4 #(
		.INIT('h0080)
	) name3902 (
		_w2549_,
		_w3001_,
		_w3700_,
		_w6129_,
		_w6131_
	);
	LUT2 #(
		.INIT('he)
	) name3903 (
		_w6130_,
		_w6131_,
		_w6132_
	);
	LUT4 #(
		.INIT('h8000)
	) name3904 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2244_,
		_w2991_,
		_w6133_
	);
	LUT3 #(
		.INIT('he0)
	) name3905 (
		_w2993_,
		_w2994_,
		_w6133_,
		_w6134_
	);
	LUT4 #(
		.INIT('h0080)
	) name3906 (
		_w2534_,
		_w3010_,
		_w3700_,
		_w6133_,
		_w6135_
	);
	LUT2 #(
		.INIT('he)
	) name3907 (
		_w6134_,
		_w6135_,
		_w6136_
	);
	LUT4 #(
		.INIT('h8000)
	) name3908 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2244_,
		_w3112_,
		_w6137_
	);
	LUT3 #(
		.INIT('he0)
	) name3909 (
		_w2993_,
		_w2994_,
		_w6137_,
		_w6138_
	);
	LUT4 #(
		.INIT('h0080)
	) name3910 (
		_w2534_,
		_w3011_,
		_w3700_,
		_w6137_,
		_w6139_
	);
	LUT2 #(
		.INIT('he)
	) name3911 (
		_w6138_,
		_w6139_,
		_w6140_
	);
	LUT4 #(
		.INIT('h8000)
	) name3912 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2229_,
		_w2230_,
		_w2991_,
		_w6141_
	);
	LUT3 #(
		.INIT('he0)
	) name3913 (
		_w2993_,
		_w2994_,
		_w6141_,
		_w6142_
	);
	LUT4 #(
		.INIT('h0080)
	) name3914 (
		_w2549_,
		_w3005_,
		_w3700_,
		_w6141_,
		_w6143_
	);
	LUT2 #(
		.INIT('he)
	) name3915 (
		_w6142_,
		_w6143_,
		_w6144_
	);
	LUT4 #(
		.INIT('h8000)
	) name3916 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2247_,
		_w2991_,
		_w6145_
	);
	LUT3 #(
		.INIT('he0)
	) name3917 (
		_w2993_,
		_w2994_,
		_w6145_,
		_w6146_
	);
	LUT4 #(
		.INIT('h0080)
	) name3918 (
		_w2520_,
		_w3002_,
		_w3700_,
		_w6145_,
		_w6147_
	);
	LUT2 #(
		.INIT('he)
	) name3919 (
		_w6146_,
		_w6147_,
		_w6148_
	);
	LUT4 #(
		.INIT('h8000)
	) name3920 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2247_,
		_w3112_,
		_w6149_
	);
	LUT3 #(
		.INIT('he0)
	) name3921 (
		_w2993_,
		_w2994_,
		_w6149_,
		_w6150_
	);
	LUT4 #(
		.INIT('h0080)
	) name3922 (
		_w2520_,
		_w3007_,
		_w3700_,
		_w6149_,
		_w6151_
	);
	LUT2 #(
		.INIT('he)
	) name3923 (
		_w6150_,
		_w6151_,
		_w6152_
	);
	LUT4 #(
		.INIT('h8000)
	) name3924 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2254_,
		_w2991_,
		_w6153_
	);
	LUT3 #(
		.INIT('he0)
	) name3925 (
		_w2993_,
		_w2994_,
		_w6153_,
		_w6154_
	);
	LUT4 #(
		.INIT('h0080)
	) name3926 (
		_w2527_,
		_w3008_,
		_w3700_,
		_w6153_,
		_w6155_
	);
	LUT2 #(
		.INIT('he)
	) name3927 (
		_w6154_,
		_w6155_,
		_w6156_
	);
	LUT4 #(
		.INIT('h8000)
	) name3928 (
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w2230_,
		_w2254_,
		_w3112_,
		_w6157_
	);
	LUT3 #(
		.INIT('he0)
	) name3929 (
		_w2993_,
		_w2994_,
		_w6157_,
		_w6158_
	);
	LUT4 #(
		.INIT('h0080)
	) name3930 (
		_w2527_,
		_w3004_,
		_w3700_,
		_w6157_,
		_w6159_
	);
	LUT2 #(
		.INIT('he)
	) name3931 (
		_w6158_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h4)
	) name3932 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		_w6161_
	);
	LUT2 #(
		.INIT('h1)
	) name3933 (
		_w6083_,
		_w6161_,
		_w6162_
	);
	LUT4 #(
		.INIT('h00ea)
	) name3934 (
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2460_,
		_w2465_,
		_w6083_,
		_w6163_
	);
	LUT3 #(
		.INIT('h13)
	) name3935 (
		_w2455_,
		_w6162_,
		_w6163_,
		_w6164_
	);
	LUT3 #(
		.INIT('h23)
	) name3936 (
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m1_is_llp_reg/NET0131 ,
		_w6165_
	);
	LUT3 #(
		.INIT('h80)
	) name3937 (
		\ctl_rf_c2_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6166_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w2534_,
		_w6166_,
		_w6167_
	);
	LUT3 #(
		.INIT('h80)
	) name3939 (
		\ctl_rf_c0_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6168_
	);
	LUT3 #(
		.INIT('h2a)
	) name3940 (
		\ctl_rf_c5_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6169_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name3941 (
		_w2514_,
		_w2518_,
		_w6168_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		_w6167_,
		_w6170_,
		_w6171_
	);
	LUT3 #(
		.INIT('h80)
	) name3943 (
		\ctl_rf_c6_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6172_
	);
	LUT3 #(
		.INIT('h2a)
	) name3944 (
		\de_de_st_reg[6]/NET0131 ,
		_w2527_,
		_w6172_,
		_w6173_
	);
	LUT3 #(
		.INIT('h80)
	) name3945 (
		\ctl_rf_c4_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6174_
	);
	LUT3 #(
		.INIT('h2a)
	) name3946 (
		\ctl_rf_c3_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6175_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name3947 (
		_w2514_,
		_w2518_,
		_w6174_,
		_w6175_,
		_w6176_
	);
	LUT3 #(
		.INIT('h2a)
	) name3948 (
		\ctl_rf_c1_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6177_
	);
	LUT3 #(
		.INIT('h2a)
	) name3949 (
		\ctl_rf_c7_rf_chllp_reg[0]/P0002 ,
		_w2507_,
		_w2508_,
		_w6178_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name3950 (
		_w2514_,
		_w2518_,
		_w6177_,
		_w6178_,
		_w6179_
	);
	LUT3 #(
		.INIT('h80)
	) name3951 (
		_w6173_,
		_w6176_,
		_w6179_,
		_w6180_
	);
	LUT3 #(
		.INIT('h15)
	) name3952 (
		_w6165_,
		_w6171_,
		_w6180_,
		_w6181_
	);
	LUT3 #(
		.INIT('h10)
	) name3953 (
		\ahb_slv_br_st_reg[0]/NET0131 ,
		\ahb_slv_br_st_reg[1]/NET0131 ,
		\ahb_slv_br_st_reg[2]/NET0131 ,
		_w6182_
	);
	LUT3 #(
		.INIT('h04)
	) name3954 (
		\ahb_slv_br_st_reg[0]/NET0131 ,
		\ahb_slv_br_st_reg[1]/NET0131 ,
		\ahb_slv_br_st_reg[2]/NET0131 ,
		_w6183_
	);
	LUT3 #(
		.INIT('h02)
	) name3955 (
		\ahb_slv_br_st_reg[0]/NET0131 ,
		\ahb_slv_br_st_reg[1]/NET0131 ,
		\ahb_slv_br_st_reg[2]/NET0131 ,
		_w6184_
	);
	LUT3 #(
		.INIT('h13)
	) name3956 (
		_w6083_,
		_w6183_,
		_w6184_,
		_w6185_
	);
	LUT4 #(
		.INIT('he9eb)
	) name3957 (
		\ahb_slv_br_st_reg[0]/NET0131 ,
		\ahb_slv_br_st_reg[1]/NET0131 ,
		\ahb_slv_br_st_reg[2]/NET0131 ,
		_w6083_,
		_w6186_
	);
	LUT4 #(
		.INIT('hea00)
	) name3958 (
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w2460_,
		_w2465_,
		_w6185_,
		_w6187_
	);
	LUT3 #(
		.INIT('hec)
	) name3959 (
		_w2455_,
		_w6186_,
		_w6187_,
		_w6188_
	);
	LUT3 #(
		.INIT('h10)
	) name3960 (
		\de_de_st_reg[5]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w6189_
	);
	LUT3 #(
		.INIT('hf8)
	) name3961 (
		_w6171_,
		_w6180_,
		_w6189_,
		_w6190_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		_w6083_,
		_w6184_,
		_w6191_
	);
	LUT3 #(
		.INIT('h40)
	) name3963 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_slv_slv_br_req_reg/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		_w6192_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		_w6192_,
		_w3383_,
		_w6193_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3965 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w6193_,
		_w6194_
	);
	LUT3 #(
		.INIT('h23)
	) name3966 (
		_w6191_,
		_w6185_,
		_w6194_,
		_w6195_
	);
	LUT3 #(
		.INIT('hd0)
	) name3967 (
		_w2455_,
		_w2466_,
		_w6182_,
		_w6196_
	);
	LUT2 #(
		.INIT('h8)
	) name3968 (
		_w6183_,
		_w6194_,
		_w6197_
	);
	LUT2 #(
		.INIT('he)
	) name3969 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h8)
	) name3970 (
		\ctl_rf_c0_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6199_
	);
	LUT3 #(
		.INIT('h80)
	) name3971 (
		_w2507_,
		_w2508_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h8)
	) name3972 (
		_w2549_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h1)
	) name3973 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6202_
	);
	LUT2 #(
		.INIT('h8)
	) name3974 (
		\ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6203_
	);
	LUT3 #(
		.INIT('he0)
	) name3975 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h8)
	) name3976 (
		_w6201_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h2)
	) name3977 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		_w6206_
	);
	LUT3 #(
		.INIT('he0)
	) name3978 (
		_w2996_,
		_w2997_,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name3979 (
		_w3175_,
		_w6207_,
		_w6208_
	);
	LUT3 #(
		.INIT('h06)
	) name3980 (
		\ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6205_,
		_w6208_,
		_w6209_
	);
	LUT4 #(
		.INIT('h1333)
	) name3981 (
		\ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6201_,
		_w6204_,
		_w6210_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		\ctl_rf_c0_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6211_
	);
	LUT3 #(
		.INIT('h80)
	) name3983 (
		_w6201_,
		_w6204_,
		_w6211_,
		_w6212_
	);
	LUT3 #(
		.INIT('h01)
	) name3984 (
		_w6208_,
		_w6210_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		\ctl_rf_c1_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6214_
	);
	LUT3 #(
		.INIT('h70)
	) name3986 (
		_w2507_,
		_w2508_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		_w2549_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6217_
	);
	LUT2 #(
		.INIT('h8)
	) name3989 (
		\ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6218_
	);
	LUT3 #(
		.INIT('he0)
	) name3990 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		_w6216_,
		_w6219_,
		_w6220_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		_w6221_
	);
	LUT3 #(
		.INIT('he0)
	) name3993 (
		_w2996_,
		_w2997_,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h4)
	) name3994 (
		_w3145_,
		_w6222_,
		_w6223_
	);
	LUT3 #(
		.INIT('h06)
	) name3995 (
		\ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6220_,
		_w6223_,
		_w6224_
	);
	LUT4 #(
		.INIT('h1333)
	) name3996 (
		\ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6216_,
		_w6219_,
		_w6225_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		\ctl_rf_c1_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c1_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6226_
	);
	LUT3 #(
		.INIT('h80)
	) name3998 (
		_w6216_,
		_w6219_,
		_w6226_,
		_w6227_
	);
	LUT3 #(
		.INIT('h01)
	) name3999 (
		_w6223_,
		_w6225_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h8)
	) name4000 (
		\ctl_rf_c2_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6229_
	);
	LUT3 #(
		.INIT('h80)
	) name4001 (
		_w2507_,
		_w2508_,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		_w2534_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6232_
	);
	LUT2 #(
		.INIT('h8)
	) name4004 (
		\ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6233_
	);
	LUT3 #(
		.INIT('he0)
	) name4005 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		_w6231_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h2)
	) name4007 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		_w6236_
	);
	LUT3 #(
		.INIT('he0)
	) name4008 (
		_w2996_,
		_w2997_,
		_w6236_,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name4009 (
		_w3155_,
		_w6237_,
		_w6238_
	);
	LUT3 #(
		.INIT('h06)
	) name4010 (
		\ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6235_,
		_w6238_,
		_w6239_
	);
	LUT4 #(
		.INIT('h1333)
	) name4011 (
		\ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6231_,
		_w6234_,
		_w6240_
	);
	LUT2 #(
		.INIT('h8)
	) name4012 (
		\ctl_rf_c2_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6241_
	);
	LUT3 #(
		.INIT('h80)
	) name4013 (
		_w6231_,
		_w6234_,
		_w6241_,
		_w6242_
	);
	LUT3 #(
		.INIT('h01)
	) name4014 (
		_w6238_,
		_w6240_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h8)
	) name4015 (
		\ctl_rf_c3_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6244_
	);
	LUT3 #(
		.INIT('h70)
	) name4016 (
		_w2507_,
		_w2508_,
		_w6244_,
		_w6245_
	);
	LUT2 #(
		.INIT('h8)
	) name4017 (
		_w2534_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h1)
	) name4018 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6247_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		\ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6248_
	);
	LUT3 #(
		.INIT('he0)
	) name4020 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h8)
	) name4021 (
		_w6246_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h2)
	) name4022 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		_w6251_
	);
	LUT3 #(
		.INIT('he0)
	) name4023 (
		_w2996_,
		_w2997_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h4)
	) name4024 (
		_w3165_,
		_w6252_,
		_w6253_
	);
	LUT3 #(
		.INIT('h06)
	) name4025 (
		\ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6250_,
		_w6253_,
		_w6254_
	);
	LUT4 #(
		.INIT('h1333)
	) name4026 (
		\ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6246_,
		_w6249_,
		_w6255_
	);
	LUT2 #(
		.INIT('h8)
	) name4027 (
		\ctl_rf_c3_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6256_
	);
	LUT3 #(
		.INIT('h80)
	) name4028 (
		_w6246_,
		_w6249_,
		_w6256_,
		_w6257_
	);
	LUT3 #(
		.INIT('h01)
	) name4029 (
		_w6253_,
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h8)
	) name4030 (
		\ctl_rf_c4_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6259_
	);
	LUT3 #(
		.INIT('h80)
	) name4031 (
		_w2507_,
		_w2508_,
		_w6259_,
		_w6260_
	);
	LUT2 #(
		.INIT('h8)
	) name4032 (
		_w2520_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h1)
	) name4033 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6262_
	);
	LUT2 #(
		.INIT('h8)
	) name4034 (
		\ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6263_
	);
	LUT3 #(
		.INIT('he0)
	) name4035 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6263_,
		_w6264_
	);
	LUT2 #(
		.INIT('h8)
	) name4036 (
		_w6261_,
		_w6264_,
		_w6265_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		_w6266_
	);
	LUT3 #(
		.INIT('he0)
	) name4038 (
		_w2996_,
		_w2997_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h4)
	) name4039 (
		_w2995_,
		_w6267_,
		_w6268_
	);
	LUT3 #(
		.INIT('h06)
	) name4040 (
		\ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6265_,
		_w6268_,
		_w6269_
	);
	LUT4 #(
		.INIT('h1333)
	) name4041 (
		\ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6261_,
		_w6264_,
		_w6270_
	);
	LUT2 #(
		.INIT('h8)
	) name4042 (
		\ctl_rf_c4_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6271_
	);
	LUT3 #(
		.INIT('h80)
	) name4043 (
		_w6261_,
		_w6264_,
		_w6271_,
		_w6272_
	);
	LUT3 #(
		.INIT('h01)
	) name4044 (
		_w6268_,
		_w6270_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h8)
	) name4045 (
		\ctl_rf_c5_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6274_
	);
	LUT3 #(
		.INIT('h70)
	) name4046 (
		_w2507_,
		_w2508_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h8)
	) name4047 (
		_w2520_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6277_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		\ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6278_
	);
	LUT3 #(
		.INIT('he0)
	) name4050 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h8)
	) name4051 (
		_w6276_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h2)
	) name4052 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		_w6281_
	);
	LUT3 #(
		.INIT('he0)
	) name4053 (
		_w2996_,
		_w2997_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h4)
	) name4054 (
		_w3114_,
		_w6282_,
		_w6283_
	);
	LUT3 #(
		.INIT('h06)
	) name4055 (
		\ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6280_,
		_w6283_,
		_w6284_
	);
	LUT4 #(
		.INIT('h1333)
	) name4056 (
		\ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6276_,
		_w6279_,
		_w6285_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		\ctl_rf_c5_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6286_
	);
	LUT3 #(
		.INIT('h80)
	) name4058 (
		_w6276_,
		_w6279_,
		_w6286_,
		_w6287_
	);
	LUT3 #(
		.INIT('h01)
	) name4059 (
		_w6283_,
		_w6285_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h8)
	) name4060 (
		\ctl_rf_c6_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6289_
	);
	LUT3 #(
		.INIT('h80)
	) name4061 (
		_w2507_,
		_w2508_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h8)
	) name4062 (
		_w2527_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6292_
	);
	LUT2 #(
		.INIT('h8)
	) name4064 (
		\ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6293_
	);
	LUT3 #(
		.INIT('he0)
	) name4065 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h8)
	) name4066 (
		_w6291_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h2)
	) name4067 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		_w6296_
	);
	LUT3 #(
		.INIT('he0)
	) name4068 (
		_w2996_,
		_w2997_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h4)
	) name4069 (
		_w3125_,
		_w6297_,
		_w6298_
	);
	LUT3 #(
		.INIT('h06)
	) name4070 (
		\ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6295_,
		_w6298_,
		_w6299_
	);
	LUT4 #(
		.INIT('h1333)
	) name4071 (
		\ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6291_,
		_w6294_,
		_w6300_
	);
	LUT2 #(
		.INIT('h8)
	) name4072 (
		\ctl_rf_c6_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6301_
	);
	LUT3 #(
		.INIT('h80)
	) name4073 (
		_w6291_,
		_w6294_,
		_w6301_,
		_w6302_
	);
	LUT3 #(
		.INIT('h01)
	) name4074 (
		_w6298_,
		_w6300_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\ctl_rf_c7_rf_chllp_on_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		_w6304_
	);
	LUT3 #(
		.INIT('h70)
	) name4076 (
		_w2507_,
		_w2508_,
		_w6304_,
		_w6305_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		_w2527_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6307_
	);
	LUT2 #(
		.INIT('h8)
	) name4079 (
		\ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6308_
	);
	LUT3 #(
		.INIT('he0)
	) name4080 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		_w2424_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		_w6306_,
		_w6309_,
		_w6310_
	);
	LUT2 #(
		.INIT('h2)
	) name4082 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		_w6311_
	);
	LUT3 #(
		.INIT('he0)
	) name4083 (
		_w2996_,
		_w2997_,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h4)
	) name4084 (
		_w3135_,
		_w6312_,
		_w6313_
	);
	LUT3 #(
		.INIT('h06)
	) name4085 (
		\ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131 ,
		_w6310_,
		_w6313_,
		_w6314_
	);
	LUT4 #(
		.INIT('h1333)
	) name4086 (
		\ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6306_,
		_w6309_,
		_w6315_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		\ctl_rf_c7_rf_chllp_cnt_reg[2]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[3]/NET0131 ,
		_w6316_
	);
	LUT3 #(
		.INIT('h80)
	) name4088 (
		_w6306_,
		_w6309_,
		_w6316_,
		_w6317_
	);
	LUT3 #(
		.INIT('h01)
	) name4089 (
		_w6313_,
		_w6315_,
		_w6317_,
		_w6318_
	);
	LUT3 #(
		.INIT('ha2)
	) name4090 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		\m1_mux_hrp_df_reg[0]/NET0131 ,
		_w6319_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4091 (
		_w2446_,
		_w2449_,
		_w2454_,
		_w6319_,
		_w6320_
	);
	LUT3 #(
		.INIT('h10)
	) name4092 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		hreadyout_br_pad,
		\hresp_br[0]_pad ,
		_w6321_
	);
	LUT3 #(
		.INIT('h54)
	) name4093 (
		_w6085_,
		_w6320_,
		_w6321_,
		_w6322_
	);
	LUT3 #(
		.INIT('ha6)
	) name4094 (
		\ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6201_,
		_w6202_,
		_w6323_
	);
	LUT2 #(
		.INIT('h4)
	) name4095 (
		_w6208_,
		_w6323_,
		_w6324_
	);
	LUT3 #(
		.INIT('ha6)
	) name4096 (
		\ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6216_,
		_w6217_,
		_w6325_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		_w6223_,
		_w6325_,
		_w6326_
	);
	LUT3 #(
		.INIT('ha6)
	) name4098 (
		\ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6276_,
		_w6277_,
		_w6327_
	);
	LUT2 #(
		.INIT('h4)
	) name4099 (
		_w6283_,
		_w6327_,
		_w6328_
	);
	LUT3 #(
		.INIT('ha6)
	) name4100 (
		\ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6231_,
		_w6232_,
		_w6329_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		_w6238_,
		_w6329_,
		_w6330_
	);
	LUT3 #(
		.INIT('ha6)
	) name4102 (
		\ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6246_,
		_w6247_,
		_w6331_
	);
	LUT2 #(
		.INIT('h4)
	) name4103 (
		_w6253_,
		_w6331_,
		_w6332_
	);
	LUT3 #(
		.INIT('ha6)
	) name4104 (
		\ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6261_,
		_w6262_,
		_w6333_
	);
	LUT2 #(
		.INIT('h4)
	) name4105 (
		_w6268_,
		_w6333_,
		_w6334_
	);
	LUT3 #(
		.INIT('ha6)
	) name4106 (
		\ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6291_,
		_w6292_,
		_w6335_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w6298_,
		_w6335_,
		_w6336_
	);
	LUT3 #(
		.INIT('ha6)
	) name4108 (
		\ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131 ,
		_w6306_,
		_w6307_,
		_w6337_
	);
	LUT2 #(
		.INIT('h4)
	) name4109 (
		_w6313_,
		_w6337_,
		_w6338_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4110 (
		\ctl_rf_c0_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c0_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6201_,
		_w6202_,
		_w6339_
	);
	LUT2 #(
		.INIT('h4)
	) name4111 (
		_w6208_,
		_w6339_,
		_w6340_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4112 (
		\ctl_rf_c1_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c1_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6216_,
		_w6217_,
		_w6341_
	);
	LUT2 #(
		.INIT('h4)
	) name4113 (
		_w6223_,
		_w6341_,
		_w6342_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4114 (
		\ctl_rf_c2_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c2_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6231_,
		_w6232_,
		_w6343_
	);
	LUT2 #(
		.INIT('h4)
	) name4115 (
		_w6238_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4116 (
		\ctl_rf_c3_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c3_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6246_,
		_w6247_,
		_w6345_
	);
	LUT2 #(
		.INIT('h4)
	) name4117 (
		_w6253_,
		_w6345_,
		_w6346_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4118 (
		\ctl_rf_c4_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c4_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6261_,
		_w6262_,
		_w6347_
	);
	LUT2 #(
		.INIT('h4)
	) name4119 (
		_w6268_,
		_w6347_,
		_w6348_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4120 (
		\ctl_rf_c5_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c5_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6276_,
		_w6277_,
		_w6349_
	);
	LUT2 #(
		.INIT('h4)
	) name4121 (
		_w6283_,
		_w6349_,
		_w6350_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4122 (
		\ctl_rf_c6_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c6_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6291_,
		_w6292_,
		_w6351_
	);
	LUT2 #(
		.INIT('h4)
	) name4123 (
		_w6298_,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4124 (
		\ctl_rf_c7_rf_chllp_cnt_reg[0]/NET0131 ,
		\ctl_rf_c7_rf_chllp_cnt_reg[1]/NET0131 ,
		_w6306_,
		_w6307_,
		_w6353_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w6313_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h2)
	) name4126 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6355_
	);
	LUT3 #(
		.INIT('h10)
	) name4127 (
		\ahb_slv_br_st_reg[2]/NET0131 ,
		hreadyout_br_pad,
		\hresp_br[1]_pad ,
		_w6356_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		_w6085_,
		_w6356_,
		_w6357_
	);
	LUT4 #(
		.INIT('h70ff)
	) name4129 (
		_w2460_,
		_w2465_,
		_w6355_,
		_w6357_,
		_w6358_
	);
	LUT2 #(
		.INIT('h2)
	) name4130 (
		_w5537_,
		_w5545_,
		_w6359_
	);
	LUT4 #(
		.INIT('h0100)
	) name4131 (
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w6360_
	);
	LUT3 #(
		.INIT('h10)
	) name4132 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w6361_
	);
	LUT3 #(
		.INIT('h40)
	) name4133 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w6362_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4134 (
		\ctl_rf_abt_reg[0]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6363_
	);
	LUT3 #(
		.INIT('h2a)
	) name4135 (
		\ctl_rf_abt_reg[0]/NET0131 ,
		\hwdata[0]_pad ,
		_w2234_,
		_w6364_
	);
	LUT3 #(
		.INIT('h23)
	) name4136 (
		_w2371_,
		_w6363_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('hb)
	) name4137 (
		_w3702_,
		_w6365_,
		_w6366_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4138 (
		\ctl_rf_abt_reg[2]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6367_
	);
	LUT3 #(
		.INIT('h2a)
	) name4139 (
		\ctl_rf_abt_reg[2]/NET0131 ,
		\hwdata[2]_pad ,
		_w2234_,
		_w6368_
	);
	LUT3 #(
		.INIT('h23)
	) name4140 (
		_w2295_,
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('hb)
	) name4141 (
		_w3717_,
		_w6369_,
		_w6370_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4142 (
		\ctl_rf_abt_reg[1]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6371_
	);
	LUT3 #(
		.INIT('h2a)
	) name4143 (
		\ctl_rf_abt_reg[1]/NET0131 ,
		\hwdata[1]_pad ,
		_w2234_,
		_w6372_
	);
	LUT3 #(
		.INIT('h23)
	) name4144 (
		_w2241_,
		_w6371_,
		_w6372_,
		_w6373_
	);
	LUT2 #(
		.INIT('hb)
	) name4145 (
		_w3710_,
		_w6373_,
		_w6374_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4146 (
		\ctl_rf_abt_reg[3]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6375_
	);
	LUT3 #(
		.INIT('h2a)
	) name4147 (
		\ctl_rf_abt_reg[3]/NET0131 ,
		\hwdata[3]_pad ,
		_w2234_,
		_w6376_
	);
	LUT3 #(
		.INIT('h23)
	) name4148 (
		_w2298_,
		_w6375_,
		_w6376_,
		_w6377_
	);
	LUT2 #(
		.INIT('hb)
	) name4149 (
		_w3724_,
		_w6377_,
		_w6378_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4150 (
		\ctl_rf_abt_reg[4]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6379_
	);
	LUT3 #(
		.INIT('h2a)
	) name4151 (
		\ctl_rf_abt_reg[4]/NET0131 ,
		\hwdata[4]_pad ,
		_w2234_,
		_w6380_
	);
	LUT3 #(
		.INIT('h23)
	) name4152 (
		_w2341_,
		_w6379_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('hb)
	) name4153 (
		_w3731_,
		_w6381_,
		_w6382_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4154 (
		\ctl_rf_abt_reg[5]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6383_
	);
	LUT3 #(
		.INIT('h2a)
	) name4155 (
		\ctl_rf_abt_reg[5]/NET0131 ,
		\hwdata[5]_pad ,
		_w2234_,
		_w6384_
	);
	LUT3 #(
		.INIT('h23)
	) name4156 (
		_w2282_,
		_w6383_,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('hb)
	) name4157 (
		_w3738_,
		_w6385_,
		_w6386_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4158 (
		\ctl_rf_abt_reg[6]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6387_
	);
	LUT3 #(
		.INIT('h2a)
	) name4159 (
		\ctl_rf_abt_reg[6]/NET0131 ,
		\hwdata[6]_pad ,
		_w2234_,
		_w6388_
	);
	LUT3 #(
		.INIT('h23)
	) name4160 (
		_w2323_,
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT2 #(
		.INIT('hb)
	) name4161 (
		_w3745_,
		_w6389_,
		_w6390_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4162 (
		\ctl_rf_abt_reg[7]/NET0131 ,
		_w6360_,
		_w6361_,
		_w6362_,
		_w6391_
	);
	LUT3 #(
		.INIT('h2a)
	) name4163 (
		\ctl_rf_abt_reg[7]/NET0131 ,
		\hwdata[7]_pad ,
		_w2234_,
		_w6392_
	);
	LUT3 #(
		.INIT('h23)
	) name4164 (
		_w2331_,
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('hb)
	) name4165 (
		_w3752_,
		_w6393_,
		_w6394_
	);
	LUT3 #(
		.INIT('h20)
	) name4166 (
		\h1prot[0]_pad ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6395_
	);
	LUT4 #(
		.INIT('h8000)
	) name4167 (
		\h1prot[0]_pad ,
		_w2390_,
		_w2393_,
		_w2396_,
		_w6396_
	);
	LUT4 #(
		.INIT('h070f)
	) name4168 (
		_w2403_,
		_w2416_,
		_w6395_,
		_w6396_,
		_w6397_
	);
	LUT4 #(
		.INIT('h8088)
	) name4169 (
		\ahb_slv_slv_pt_d1o_reg[0]/NET0131 ,
		\de_m1_arb_st_reg[1]/NET0131 ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6398_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4170 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w6398_,
		_w6399_
	);
	LUT2 #(
		.INIT('hd)
	) name4171 (
		_w6397_,
		_w6399_,
		_w6400_
	);
	LUT4 #(
		.INIT('he0ee)
	) name4172 (
		\ahb_mst1_mx_cmd_st_reg[0]/NET0131 ,
		\ahb_mst1_mx_cmd_st_reg[1]/NET0131 ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6401_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4173 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w6401_,
		_w6402_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4174 (
		_w2397_,
		_w2403_,
		_w2416_,
		_w3383_,
		_w6403_
	);
	LUT3 #(
		.INIT('h20)
	) name4175 (
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		\m1_mux_hrdy_df_reg/NET0131 ,
		\m1_mux_hrmxnof_reg/NET0131 ,
		_w6404_
	);
	LUT4 #(
		.INIT('h8000)
	) name4176 (
		\ahb_mst1_mx_dtp_reg/NET0131 ,
		_w2390_,
		_w2393_,
		_w2396_,
		_w6405_
	);
	LUT4 #(
		.INIT('h070f)
	) name4177 (
		_w2403_,
		_w2416_,
		_w6404_,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('hb)
	) name4178 (
		_w6403_,
		_w6406_,
		_w6407_
	);
	LUT2 #(
		.INIT('h4)
	) name4179 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w6408_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4180 (
		\ctl_rf_tc_reg[7]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6409_
	);
	LUT3 #(
		.INIT('h2a)
	) name4181 (
		\ctl_rf_tc_reg[7]/NET0131 ,
		\hwdata[23]_pad ,
		_w2234_,
		_w6410_
	);
	LUT3 #(
		.INIT('h23)
	) name4182 (
		_w2236_,
		_w6409_,
		_w6410_,
		_w6411_
	);
	LUT3 #(
		.INIT('h15)
	) name4183 (
		\ctl_rf_c7_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6412_
	);
	LUT4 #(
		.INIT('h8000)
	) name4184 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2527_,
		_w6412_,
		_w6413_
	);
	LUT2 #(
		.INIT('hd)
	) name4185 (
		_w6411_,
		_w6413_,
		_w6414_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4186 (
		\ctl_rf_tc_reg[3]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6415_
	);
	LUT3 #(
		.INIT('h2a)
	) name4187 (
		\ctl_rf_tc_reg[3]/NET0131 ,
		\hwdata[19]_pad ,
		_w2234_,
		_w6416_
	);
	LUT3 #(
		.INIT('h23)
	) name4188 (
		_w5375_,
		_w6415_,
		_w6416_,
		_w6417_
	);
	LUT3 #(
		.INIT('h15)
	) name4189 (
		\ctl_rf_c3_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6418_
	);
	LUT4 #(
		.INIT('h8000)
	) name4190 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2534_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('hd)
	) name4191 (
		_w6417_,
		_w6419_,
		_w6420_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4192 (
		\ctl_rf_tc_reg[0]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6421_
	);
	LUT3 #(
		.INIT('h2a)
	) name4193 (
		\ctl_rf_tc_reg[0]/NET0131 ,
		\hwdata[16]_pad ,
		_w2234_,
		_w6422_
	);
	LUT3 #(
		.INIT('h23)
	) name4194 (
		_w2996_,
		_w6421_,
		_w6422_,
		_w6423_
	);
	LUT3 #(
		.INIT('h40)
	) name4195 (
		\ctl_rf_c0_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6424_
	);
	LUT4 #(
		.INIT('h8000)
	) name4196 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2549_,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('hd)
	) name4197 (
		_w6423_,
		_w6425_,
		_w6426_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4198 (
		\ctl_rf_tc_reg[1]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6427_
	);
	LUT3 #(
		.INIT('h2a)
	) name4199 (
		\ctl_rf_tc_reg[1]/NET0131 ,
		\hwdata[17]_pad ,
		_w2234_,
		_w6428_
	);
	LUT3 #(
		.INIT('h23)
	) name4200 (
		_w5359_,
		_w6427_,
		_w6428_,
		_w6429_
	);
	LUT3 #(
		.INIT('h15)
	) name4201 (
		\ctl_rf_c1_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6430_
	);
	LUT4 #(
		.INIT('h8000)
	) name4202 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2549_,
		_w6430_,
		_w6431_
	);
	LUT2 #(
		.INIT('hd)
	) name4203 (
		_w6429_,
		_w6431_,
		_w6432_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4204 (
		\ctl_rf_tc_reg[4]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6433_
	);
	LUT3 #(
		.INIT('h2a)
	) name4205 (
		\ctl_rf_tc_reg[4]/NET0131 ,
		\hwdata[20]_pad ,
		_w2234_,
		_w6434_
	);
	LUT3 #(
		.INIT('h23)
	) name4206 (
		_w5275_,
		_w6433_,
		_w6434_,
		_w6435_
	);
	LUT3 #(
		.INIT('h40)
	) name4207 (
		\ctl_rf_c4_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6436_
	);
	LUT4 #(
		.INIT('h8000)
	) name4208 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2520_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('hd)
	) name4209 (
		_w6435_,
		_w6437_,
		_w6438_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4210 (
		\ctl_rf_tc_reg[2]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6439_
	);
	LUT3 #(
		.INIT('h2a)
	) name4211 (
		\ctl_rf_tc_reg[2]/NET0131 ,
		\hwdata[18]_pad ,
		_w2234_,
		_w6440_
	);
	LUT3 #(
		.INIT('h23)
	) name4212 (
		_w5362_,
		_w6439_,
		_w6440_,
		_w6441_
	);
	LUT3 #(
		.INIT('h40)
	) name4213 (
		\ctl_rf_c2_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6442_
	);
	LUT4 #(
		.INIT('h8000)
	) name4214 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2534_,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('hd)
	) name4215 (
		_w6441_,
		_w6443_,
		_w6444_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4216 (
		\ctl_rf_tc_reg[6]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6445_
	);
	LUT3 #(
		.INIT('h2a)
	) name4217 (
		\ctl_rf_tc_reg[6]/NET0131 ,
		\hwdata[22]_pad ,
		_w2234_,
		_w6446_
	);
	LUT3 #(
		.INIT('h23)
	) name4218 (
		_w5236_,
		_w6445_,
		_w6446_,
		_w6447_
	);
	LUT3 #(
		.INIT('h40)
	) name4219 (
		\ctl_rf_c6_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6448_
	);
	LUT4 #(
		.INIT('h8000)
	) name4220 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2527_,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('hd)
	) name4221 (
		_w6447_,
		_w6449_,
		_w6450_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4222 (
		\ctl_rf_tc_reg[5]/NET0131 ,
		_w2249_,
		_w6360_,
		_w6408_,
		_w6451_
	);
	LUT3 #(
		.INIT('h2a)
	) name4223 (
		\ctl_rf_tc_reg[5]/NET0131 ,
		\hwdata[21]_pad ,
		_w2234_,
		_w6452_
	);
	LUT3 #(
		.INIT('h23)
	) name4224 (
		_w5233_,
		_w6451_,
		_w6452_,
		_w6453_
	);
	LUT3 #(
		.INIT('h15)
	) name4225 (
		\ctl_rf_c5_rf_int_tc_msk_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6454_
	);
	LUT4 #(
		.INIT('h8000)
	) name4226 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w2520_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('hd)
	) name4227 (
		_w6453_,
		_w6455_,
		_w6456_
	);
	LUT3 #(
		.INIT('h80)
	) name4228 (
		\ctl_rf_c2_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6457_
	);
	LUT3 #(
		.INIT('h2a)
	) name4229 (
		\ctl_rf_c1_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6458_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4230 (
		_w2514_,
		_w2518_,
		_w6457_,
		_w6458_,
		_w6459_
	);
	LUT3 #(
		.INIT('h2a)
	) name4231 (
		\ctl_rf_c7_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6460_
	);
	LUT3 #(
		.INIT('h80)
	) name4232 (
		\ctl_rf_c0_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6461_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4233 (
		_w2514_,
		_w2518_,
		_w6460_,
		_w6461_,
		_w6462_
	);
	LUT3 #(
		.INIT('h2a)
	) name4234 (
		\ctl_rf_c3_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6463_
	);
	LUT3 #(
		.INIT('h80)
	) name4235 (
		\ctl_rf_c6_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6464_
	);
	LUT4 #(
		.INIT('haebf)
	) name4236 (
		_w2514_,
		_w2518_,
		_w6463_,
		_w6464_,
		_w6465_
	);
	LUT3 #(
		.INIT('h2a)
	) name4237 (
		\ctl_rf_c5_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6466_
	);
	LUT3 #(
		.INIT('h80)
	) name4238 (
		\ctl_rf_c4_rf_dwidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6467_
	);
	LUT3 #(
		.INIT('h57)
	) name4239 (
		_w2520_,
		_w6466_,
		_w6467_,
		_w6468_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4240 (
		_w6459_,
		_w6462_,
		_w6465_,
		_w6468_,
		_w6469_
	);
	LUT3 #(
		.INIT('h80)
	) name4241 (
		\ctl_rf_c2_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6470_
	);
	LUT3 #(
		.INIT('h2a)
	) name4242 (
		\ctl_rf_c1_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6471_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4243 (
		_w2514_,
		_w2518_,
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT3 #(
		.INIT('h2a)
	) name4244 (
		\ctl_rf_c7_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6473_
	);
	LUT3 #(
		.INIT('h80)
	) name4245 (
		\ctl_rf_c0_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6474_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4246 (
		_w2514_,
		_w2518_,
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT3 #(
		.INIT('h2a)
	) name4247 (
		\ctl_rf_c3_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6476_
	);
	LUT3 #(
		.INIT('h80)
	) name4248 (
		\ctl_rf_c6_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6477_
	);
	LUT4 #(
		.INIT('haebf)
	) name4249 (
		_w2514_,
		_w2518_,
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT3 #(
		.INIT('h2a)
	) name4250 (
		\ctl_rf_c5_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6479_
	);
	LUT3 #(
		.INIT('h80)
	) name4251 (
		\ctl_rf_c4_rf_dst_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6480_
	);
	LUT3 #(
		.INIT('h57)
	) name4252 (
		_w2520_,
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4253 (
		_w6472_,
		_w6475_,
		_w6478_,
		_w6481_,
		_w6482_
	);
	LUT3 #(
		.INIT('h80)
	) name4254 (
		\ctl_rf_c2_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6483_
	);
	LUT3 #(
		.INIT('h2a)
	) name4255 (
		\ctl_rf_c1_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6484_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4256 (
		_w2514_,
		_w2518_,
		_w6483_,
		_w6484_,
		_w6485_
	);
	LUT3 #(
		.INIT('h2a)
	) name4257 (
		\ctl_rf_c7_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6486_
	);
	LUT3 #(
		.INIT('h80)
	) name4258 (
		\ctl_rf_c0_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6487_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4259 (
		_w2514_,
		_w2518_,
		_w6486_,
		_w6487_,
		_w6488_
	);
	LUT3 #(
		.INIT('h2a)
	) name4260 (
		\ctl_rf_c3_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6489_
	);
	LUT3 #(
		.INIT('h80)
	) name4261 (
		\ctl_rf_c6_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6490_
	);
	LUT4 #(
		.INIT('haebf)
	) name4262 (
		_w2514_,
		_w2518_,
		_w6489_,
		_w6490_,
		_w6491_
	);
	LUT3 #(
		.INIT('h2a)
	) name4263 (
		\ctl_rf_c5_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6492_
	);
	LUT3 #(
		.INIT('h80)
	) name4264 (
		\ctl_rf_c4_rf_swidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6493_
	);
	LUT3 #(
		.INIT('h57)
	) name4265 (
		_w2520_,
		_w6492_,
		_w6493_,
		_w6494_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4266 (
		_w6485_,
		_w6488_,
		_w6491_,
		_w6494_,
		_w6495_
	);
	LUT3 #(
		.INIT('h80)
	) name4267 (
		\ctl_rf_c2_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6496_
	);
	LUT3 #(
		.INIT('h2a)
	) name4268 (
		\ctl_rf_c1_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6497_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4269 (
		_w2514_,
		_w2518_,
		_w6496_,
		_w6497_,
		_w6498_
	);
	LUT3 #(
		.INIT('h2a)
	) name4270 (
		\ctl_rf_c7_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6499_
	);
	LUT3 #(
		.INIT('h80)
	) name4271 (
		\ctl_rf_c0_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6500_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4272 (
		_w2514_,
		_w2518_,
		_w6499_,
		_w6500_,
		_w6501_
	);
	LUT3 #(
		.INIT('h2a)
	) name4273 (
		\ctl_rf_c3_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6502_
	);
	LUT3 #(
		.INIT('h80)
	) name4274 (
		\ctl_rf_c6_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6503_
	);
	LUT4 #(
		.INIT('haebf)
	) name4275 (
		_w2514_,
		_w2518_,
		_w6502_,
		_w6503_,
		_w6504_
	);
	LUT3 #(
		.INIT('h2a)
	) name4276 (
		\ctl_rf_c5_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6505_
	);
	LUT3 #(
		.INIT('h80)
	) name4277 (
		\ctl_rf_c4_rf_dwidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6506_
	);
	LUT3 #(
		.INIT('h57)
	) name4278 (
		_w2520_,
		_w6505_,
		_w6506_,
		_w6507_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4279 (
		_w6498_,
		_w6501_,
		_w6504_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('h80)
	) name4280 (
		\ctl_rf_c2_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6509_
	);
	LUT3 #(
		.INIT('h2a)
	) name4281 (
		\ctl_rf_c1_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6510_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4282 (
		_w2514_,
		_w2518_,
		_w6509_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('h2a)
	) name4283 (
		\ctl_rf_c7_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6512_
	);
	LUT3 #(
		.INIT('h80)
	) name4284 (
		\ctl_rf_c0_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6513_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4285 (
		_w2514_,
		_w2518_,
		_w6512_,
		_w6513_,
		_w6514_
	);
	LUT3 #(
		.INIT('h2a)
	) name4286 (
		\ctl_rf_c3_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6515_
	);
	LUT3 #(
		.INIT('h80)
	) name4287 (
		\ctl_rf_c6_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6516_
	);
	LUT4 #(
		.INIT('haebf)
	) name4288 (
		_w2514_,
		_w2518_,
		_w6515_,
		_w6516_,
		_w6517_
	);
	LUT3 #(
		.INIT('h2a)
	) name4289 (
		\ctl_rf_c5_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6518_
	);
	LUT3 #(
		.INIT('h80)
	) name4290 (
		\ctl_rf_c4_rf_prot1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6519_
	);
	LUT3 #(
		.INIT('h57)
	) name4291 (
		_w2520_,
		_w6518_,
		_w6519_,
		_w6520_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4292 (
		_w6511_,
		_w6514_,
		_w6517_,
		_w6520_,
		_w6521_
	);
	LUT3 #(
		.INIT('h80)
	) name4293 (
		\ctl_rf_c2_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6522_
	);
	LUT3 #(
		.INIT('h2a)
	) name4294 (
		\ctl_rf_c1_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6523_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4295 (
		_w2514_,
		_w2518_,
		_w6522_,
		_w6523_,
		_w6524_
	);
	LUT3 #(
		.INIT('h2a)
	) name4296 (
		\ctl_rf_c7_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6525_
	);
	LUT3 #(
		.INIT('h80)
	) name4297 (
		\ctl_rf_c0_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6526_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4298 (
		_w2514_,
		_w2518_,
		_w6525_,
		_w6526_,
		_w6527_
	);
	LUT3 #(
		.INIT('h2a)
	) name4299 (
		\ctl_rf_c3_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6528_
	);
	LUT3 #(
		.INIT('h80)
	) name4300 (
		\ctl_rf_c6_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6529_
	);
	LUT4 #(
		.INIT('haebf)
	) name4301 (
		_w2514_,
		_w2518_,
		_w6528_,
		_w6529_,
		_w6530_
	);
	LUT3 #(
		.INIT('h2a)
	) name4302 (
		\ctl_rf_c5_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6531_
	);
	LUT3 #(
		.INIT('h80)
	) name4303 (
		\ctl_rf_c4_rf_sad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6532_
	);
	LUT3 #(
		.INIT('h57)
	) name4304 (
		_w2520_,
		_w6531_,
		_w6532_,
		_w6533_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4305 (
		_w6524_,
		_w6527_,
		_w6530_,
		_w6533_,
		_w6534_
	);
	LUT3 #(
		.INIT('h80)
	) name4306 (
		\ctl_rf_c2_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6535_
	);
	LUT3 #(
		.INIT('h2a)
	) name4307 (
		\ctl_rf_c1_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6536_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4308 (
		_w2514_,
		_w2518_,
		_w6535_,
		_w6536_,
		_w6537_
	);
	LUT3 #(
		.INIT('h2a)
	) name4309 (
		\ctl_rf_c7_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6538_
	);
	LUT3 #(
		.INIT('h80)
	) name4310 (
		\ctl_rf_c0_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6539_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4311 (
		_w2514_,
		_w2518_,
		_w6538_,
		_w6539_,
		_w6540_
	);
	LUT3 #(
		.INIT('h2a)
	) name4312 (
		\ctl_rf_c3_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6541_
	);
	LUT3 #(
		.INIT('h80)
	) name4313 (
		\ctl_rf_c6_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6542_
	);
	LUT4 #(
		.INIT('haebf)
	) name4314 (
		_w2514_,
		_w2518_,
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT3 #(
		.INIT('h2a)
	) name4315 (
		\ctl_rf_c5_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6544_
	);
	LUT3 #(
		.INIT('h80)
	) name4316 (
		\ctl_rf_c4_rf_swidth_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6545_
	);
	LUT3 #(
		.INIT('h57)
	) name4317 (
		_w2520_,
		_w6544_,
		_w6545_,
		_w6546_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4318 (
		_w6537_,
		_w6540_,
		_w6543_,
		_w6546_,
		_w6547_
	);
	LUT3 #(
		.INIT('h80)
	) name4319 (
		\ctl_rf_c2_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6548_
	);
	LUT3 #(
		.INIT('h2a)
	) name4320 (
		\ctl_rf_c1_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6549_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4321 (
		_w2514_,
		_w2518_,
		_w6548_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h2a)
	) name4322 (
		\ctl_rf_c7_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6551_
	);
	LUT3 #(
		.INIT('h80)
	) name4323 (
		\ctl_rf_c0_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6552_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4324 (
		_w2514_,
		_w2518_,
		_w6551_,
		_w6552_,
		_w6553_
	);
	LUT3 #(
		.INIT('h2a)
	) name4325 (
		\ctl_rf_c3_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6554_
	);
	LUT3 #(
		.INIT('h80)
	) name4326 (
		\ctl_rf_c6_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6555_
	);
	LUT4 #(
		.INIT('haebf)
	) name4327 (
		_w2514_,
		_w2518_,
		_w6554_,
		_w6555_,
		_w6556_
	);
	LUT3 #(
		.INIT('h2a)
	) name4328 (
		\ctl_rf_c5_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6557_
	);
	LUT3 #(
		.INIT('h80)
	) name4329 (
		\ctl_rf_c4_rf_swidth_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6558_
	);
	LUT3 #(
		.INIT('h57)
	) name4330 (
		_w2520_,
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4331 (
		_w6550_,
		_w6553_,
		_w6556_,
		_w6559_,
		_w6560_
	);
	LUT3 #(
		.INIT('h80)
	) name4332 (
		\ctl_rf_c2_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6561_
	);
	LUT3 #(
		.INIT('h2a)
	) name4333 (
		\ctl_rf_c1_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6562_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4334 (
		_w2514_,
		_w2518_,
		_w6561_,
		_w6562_,
		_w6563_
	);
	LUT3 #(
		.INIT('h2a)
	) name4335 (
		\ctl_rf_c7_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6564_
	);
	LUT3 #(
		.INIT('h80)
	) name4336 (
		\ctl_rf_c0_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6565_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4337 (
		_w2514_,
		_w2518_,
		_w6564_,
		_w6565_,
		_w6566_
	);
	LUT3 #(
		.INIT('h2a)
	) name4338 (
		\ctl_rf_c3_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6567_
	);
	LUT3 #(
		.INIT('h80)
	) name4339 (
		\ctl_rf_c6_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6568_
	);
	LUT4 #(
		.INIT('haebf)
	) name4340 (
		_w2514_,
		_w2518_,
		_w6567_,
		_w6568_,
		_w6569_
	);
	LUT3 #(
		.INIT('h2a)
	) name4341 (
		\ctl_rf_c5_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6570_
	);
	LUT3 #(
		.INIT('h80)
	) name4342 (
		\ctl_rf_c4_rf_src_sz_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6571_
	);
	LUT3 #(
		.INIT('h57)
	) name4343 (
		_w2520_,
		_w6570_,
		_w6571_,
		_w6572_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4344 (
		_w6563_,
		_w6566_,
		_w6569_,
		_w6572_,
		_w6573_
	);
	LUT3 #(
		.INIT('h80)
	) name4345 (
		\ctl_rf_c2_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6574_
	);
	LUT3 #(
		.INIT('h2a)
	) name4346 (
		\ctl_rf_c1_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6575_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4347 (
		_w2514_,
		_w2518_,
		_w6574_,
		_w6575_,
		_w6576_
	);
	LUT3 #(
		.INIT('h2a)
	) name4348 (
		\ctl_rf_c7_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6577_
	);
	LUT3 #(
		.INIT('h80)
	) name4349 (
		\ctl_rf_c0_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6578_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4350 (
		_w2514_,
		_w2518_,
		_w6577_,
		_w6578_,
		_w6579_
	);
	LUT3 #(
		.INIT('h2a)
	) name4351 (
		\ctl_rf_c3_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6580_
	);
	LUT3 #(
		.INIT('h80)
	) name4352 (
		\ctl_rf_c6_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6581_
	);
	LUT4 #(
		.INIT('haebf)
	) name4353 (
		_w2514_,
		_w2518_,
		_w6580_,
		_w6581_,
		_w6582_
	);
	LUT3 #(
		.INIT('h2a)
	) name4354 (
		\ctl_rf_c5_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6583_
	);
	LUT3 #(
		.INIT('h80)
	) name4355 (
		\ctl_rf_c4_rf_src_sel_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6584_
	);
	LUT3 #(
		.INIT('h57)
	) name4356 (
		_w2520_,
		_w6583_,
		_w6584_,
		_w6585_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4357 (
		_w6576_,
		_w6579_,
		_w6582_,
		_w6585_,
		_w6586_
	);
	LUT3 #(
		.INIT('h80)
	) name4358 (
		\ctl_rf_c2_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6587_
	);
	LUT3 #(
		.INIT('h2a)
	) name4359 (
		\ctl_rf_c1_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6588_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4360 (
		_w2514_,
		_w2518_,
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT3 #(
		.INIT('h2a)
	) name4361 (
		\ctl_rf_c7_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6590_
	);
	LUT3 #(
		.INIT('h80)
	) name4362 (
		\ctl_rf_c0_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6591_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4363 (
		_w2514_,
		_w2518_,
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('h2a)
	) name4364 (
		\ctl_rf_c3_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6593_
	);
	LUT3 #(
		.INIT('h80)
	) name4365 (
		\ctl_rf_c6_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6594_
	);
	LUT4 #(
		.INIT('haebf)
	) name4366 (
		_w2514_,
		_w2518_,
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT3 #(
		.INIT('h2a)
	) name4367 (
		\ctl_rf_c5_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6596_
	);
	LUT3 #(
		.INIT('h80)
	) name4368 (
		\ctl_rf_c4_rf_dad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6597_
	);
	LUT3 #(
		.INIT('h57)
	) name4369 (
		_w2520_,
		_w6596_,
		_w6597_,
		_w6598_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4370 (
		_w6589_,
		_w6592_,
		_w6595_,
		_w6598_,
		_w6599_
	);
	LUT3 #(
		.INIT('h80)
	) name4371 (
		\ctl_rf_c2_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6600_
	);
	LUT3 #(
		.INIT('h2a)
	) name4372 (
		\ctl_rf_c1_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6601_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4373 (
		_w2514_,
		_w2518_,
		_w6600_,
		_w6601_,
		_w6602_
	);
	LUT3 #(
		.INIT('h2a)
	) name4374 (
		\ctl_rf_c7_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6603_
	);
	LUT3 #(
		.INIT('h80)
	) name4375 (
		\ctl_rf_c0_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6604_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4376 (
		_w2514_,
		_w2518_,
		_w6603_,
		_w6604_,
		_w6605_
	);
	LUT3 #(
		.INIT('h2a)
	) name4377 (
		\ctl_rf_c3_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6606_
	);
	LUT3 #(
		.INIT('h80)
	) name4378 (
		\ctl_rf_c6_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6607_
	);
	LUT4 #(
		.INIT('haebf)
	) name4379 (
		_w2514_,
		_w2518_,
		_w6606_,
		_w6607_,
		_w6608_
	);
	LUT3 #(
		.INIT('h2a)
	) name4380 (
		\ctl_rf_c5_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6609_
	);
	LUT3 #(
		.INIT('h80)
	) name4381 (
		\ctl_rf_c4_rf_dad_ctl1_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6610_
	);
	LUT3 #(
		.INIT('h57)
	) name4382 (
		_w2520_,
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4383 (
		_w6602_,
		_w6605_,
		_w6608_,
		_w6611_,
		_w6612_
	);
	LUT3 #(
		.INIT('h80)
	) name4384 (
		\ctl_rf_c2_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6613_
	);
	LUT3 #(
		.INIT('h2a)
	) name4385 (
		\ctl_rf_c1_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6614_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4386 (
		_w2514_,
		_w2518_,
		_w6613_,
		_w6614_,
		_w6615_
	);
	LUT3 #(
		.INIT('h2a)
	) name4387 (
		\ctl_rf_c7_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6616_
	);
	LUT3 #(
		.INIT('h80)
	) name4388 (
		\ctl_rf_c0_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6617_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4389 (
		_w2514_,
		_w2518_,
		_w6616_,
		_w6617_,
		_w6618_
	);
	LUT3 #(
		.INIT('h2a)
	) name4390 (
		\ctl_rf_c3_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6619_
	);
	LUT3 #(
		.INIT('h80)
	) name4391 (
		\ctl_rf_c6_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6620_
	);
	LUT4 #(
		.INIT('haebf)
	) name4392 (
		_w2514_,
		_w2518_,
		_w6619_,
		_w6620_,
		_w6621_
	);
	LUT3 #(
		.INIT('h2a)
	) name4393 (
		\ctl_rf_c5_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6622_
	);
	LUT3 #(
		.INIT('h80)
	) name4394 (
		\ctl_rf_c4_rf_sad_ctl0_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6623_
	);
	LUT3 #(
		.INIT('h57)
	) name4395 (
		_w2520_,
		_w6622_,
		_w6623_,
		_w6624_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4396 (
		_w6615_,
		_w6618_,
		_w6621_,
		_w6624_,
		_w6625_
	);
	LUT3 #(
		.INIT('h80)
	) name4397 (
		\ctl_rf_c2_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6626_
	);
	LUT3 #(
		.INIT('h2a)
	) name4398 (
		\ctl_rf_c1_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6627_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4399 (
		_w2514_,
		_w2518_,
		_w6626_,
		_w6627_,
		_w6628_
	);
	LUT3 #(
		.INIT('h2a)
	) name4400 (
		\ctl_rf_c7_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6629_
	);
	LUT3 #(
		.INIT('h80)
	) name4401 (
		\ctl_rf_c0_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6630_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4402 (
		_w2514_,
		_w2518_,
		_w6629_,
		_w6630_,
		_w6631_
	);
	LUT3 #(
		.INIT('h2a)
	) name4403 (
		\ctl_rf_c3_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6632_
	);
	LUT3 #(
		.INIT('h80)
	) name4404 (
		\ctl_rf_c6_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6633_
	);
	LUT4 #(
		.INIT('haebf)
	) name4405 (
		_w2514_,
		_w2518_,
		_w6632_,
		_w6633_,
		_w6634_
	);
	LUT3 #(
		.INIT('h2a)
	) name4406 (
		\ctl_rf_c5_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6635_
	);
	LUT3 #(
		.INIT('h80)
	) name4407 (
		\ctl_rf_c4_rf_dwidth_reg[0]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6636_
	);
	LUT3 #(
		.INIT('h57)
	) name4408 (
		_w2520_,
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4409 (
		_w6628_,
		_w6631_,
		_w6634_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h80)
	) name4410 (
		\ctl_rf_c2_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6639_
	);
	LUT3 #(
		.INIT('h2a)
	) name4411 (
		\ctl_rf_c1_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6640_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4412 (
		_w2514_,
		_w2518_,
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT3 #(
		.INIT('h2a)
	) name4413 (
		\ctl_rf_c7_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6642_
	);
	LUT3 #(
		.INIT('h80)
	) name4414 (
		\ctl_rf_c0_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6643_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4415 (
		_w2514_,
		_w2518_,
		_w6642_,
		_w6643_,
		_w6644_
	);
	LUT3 #(
		.INIT('h2a)
	) name4416 (
		\ctl_rf_c3_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6645_
	);
	LUT3 #(
		.INIT('h80)
	) name4417 (
		\ctl_rf_c6_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6646_
	);
	LUT4 #(
		.INIT('haebf)
	) name4418 (
		_w2514_,
		_w2518_,
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT3 #(
		.INIT('h2a)
	) name4419 (
		\ctl_rf_c5_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6648_
	);
	LUT3 #(
		.INIT('h80)
	) name4420 (
		\ctl_rf_c4_rf_prot2_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6649_
	);
	LUT3 #(
		.INIT('h57)
	) name4421 (
		_w2520_,
		_w6648_,
		_w6649_,
		_w6650_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4422 (
		_w6641_,
		_w6644_,
		_w6647_,
		_w6650_,
		_w6651_
	);
	LUT3 #(
		.INIT('h80)
	) name4423 (
		\ctl_rf_c2_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6652_
	);
	LUT3 #(
		.INIT('h2a)
	) name4424 (
		\ctl_rf_c1_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6653_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4425 (
		_w2514_,
		_w2518_,
		_w6652_,
		_w6653_,
		_w6654_
	);
	LUT3 #(
		.INIT('h2a)
	) name4426 (
		\ctl_rf_c7_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6655_
	);
	LUT3 #(
		.INIT('h80)
	) name4427 (
		\ctl_rf_c0_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6656_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4428 (
		_w2514_,
		_w2518_,
		_w6655_,
		_w6656_,
		_w6657_
	);
	LUT3 #(
		.INIT('h2a)
	) name4429 (
		\ctl_rf_c3_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6658_
	);
	LUT3 #(
		.INIT('h80)
	) name4430 (
		\ctl_rf_c6_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6659_
	);
	LUT4 #(
		.INIT('haebf)
	) name4431 (
		_w2514_,
		_w2518_,
		_w6658_,
		_w6659_,
		_w6660_
	);
	LUT3 #(
		.INIT('h2a)
	) name4432 (
		\ctl_rf_c5_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6661_
	);
	LUT3 #(
		.INIT('h80)
	) name4433 (
		\ctl_rf_c4_rf_src_sz_reg[1]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6662_
	);
	LUT3 #(
		.INIT('h57)
	) name4434 (
		_w2520_,
		_w6661_,
		_w6662_,
		_w6663_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4435 (
		_w6654_,
		_w6657_,
		_w6660_,
		_w6663_,
		_w6664_
	);
	LUT3 #(
		.INIT('h80)
	) name4436 (
		\ctl_rf_c2_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6665_
	);
	LUT3 #(
		.INIT('h2a)
	) name4437 (
		\ctl_rf_c1_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6666_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4438 (
		_w2514_,
		_w2518_,
		_w6665_,
		_w6666_,
		_w6667_
	);
	LUT3 #(
		.INIT('h2a)
	) name4439 (
		\ctl_rf_c7_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6668_
	);
	LUT3 #(
		.INIT('h80)
	) name4440 (
		\ctl_rf_c0_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6669_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4441 (
		_w2514_,
		_w2518_,
		_w6668_,
		_w6669_,
		_w6670_
	);
	LUT3 #(
		.INIT('h2a)
	) name4442 (
		\ctl_rf_c3_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6671_
	);
	LUT3 #(
		.INIT('h80)
	) name4443 (
		\ctl_rf_c6_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6672_
	);
	LUT4 #(
		.INIT('haebf)
	) name4444 (
		_w2514_,
		_w2518_,
		_w6671_,
		_w6672_,
		_w6673_
	);
	LUT3 #(
		.INIT('h2a)
	) name4445 (
		\ctl_rf_c5_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6674_
	);
	LUT3 #(
		.INIT('h80)
	) name4446 (
		\ctl_rf_c4_rf_prot3_reg/NET0131 ,
		_w2507_,
		_w2508_,
		_w6675_
	);
	LUT3 #(
		.INIT('h57)
	) name4447 (
		_w2520_,
		_w6674_,
		_w6675_,
		_w6676_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4448 (
		_w6667_,
		_w6670_,
		_w6673_,
		_w6676_,
		_w6677_
	);
	LUT3 #(
		.INIT('h80)
	) name4449 (
		\ctl_rf_c2_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6678_
	);
	LUT3 #(
		.INIT('h2a)
	) name4450 (
		\ctl_rf_c1_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6679_
	);
	LUT4 #(
		.INIT('h37bf)
	) name4451 (
		_w2514_,
		_w2518_,
		_w6678_,
		_w6679_,
		_w6680_
	);
	LUT3 #(
		.INIT('h2a)
	) name4452 (
		\ctl_rf_c7_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6681_
	);
	LUT3 #(
		.INIT('h80)
	) name4453 (
		\ctl_rf_c0_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6682_
	);
	LUT4 #(
		.INIT('h67ef)
	) name4454 (
		_w2514_,
		_w2518_,
		_w6681_,
		_w6682_,
		_w6683_
	);
	LUT3 #(
		.INIT('h2a)
	) name4455 (
		\ctl_rf_c3_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6684_
	);
	LUT3 #(
		.INIT('h80)
	) name4456 (
		\ctl_rf_c6_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6685_
	);
	LUT4 #(
		.INIT('haebf)
	) name4457 (
		_w2514_,
		_w2518_,
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('h2a)
	) name4458 (
		\ctl_rf_c5_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6687_
	);
	LUT3 #(
		.INIT('h80)
	) name4459 (
		\ctl_rf_c4_rf_src_sz_reg[2]/NET0131 ,
		_w2507_,
		_w2508_,
		_w6688_
	);
	LUT3 #(
		.INIT('h57)
	) name4460 (
		_w2520_,
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4461 (
		_w6680_,
		_w6683_,
		_w6686_,
		_w6689_,
		_w6690_
	);
	LUT4 #(
		.INIT('h153f)
	) name4462 (
		\h1rdt0_dma[13]_pad ,
		\h1rdt1_br[13]_pad ,
		_w2400_,
		_w2414_,
		_w6691_
	);
	LUT4 #(
		.INIT('h153f)
	) name4463 (
		\h1rdt2_dma[13]_pad ,
		\h1rdt4_br[13]_pad ,
		_w2405_,
		_w2410_,
		_w6692_
	);
	LUT4 #(
		.INIT('h153f)
	) name4464 (
		\h1rdt5_dma[13]_pad ,
		\h1rdt7_br[13]_pad ,
		_w2391_,
		_w2401_,
		_w6693_
	);
	LUT4 #(
		.INIT('h153f)
	) name4465 (
		\h1rdt1_dma[13]_pad ,
		\h1rdt6_br[13]_pad ,
		_w2392_,
		_w2395_,
		_w6694_
	);
	LUT4 #(
		.INIT('h8000)
	) name4466 (
		_w6691_,
		_w6692_,
		_w6693_,
		_w6694_,
		_w6695_
	);
	LUT4 #(
		.INIT('h153f)
	) name4467 (
		\h1rdt4_dma[13]_pad ,
		\h1rdt5_br[13]_pad ,
		_w2408_,
		_w2411_,
		_w6696_
	);
	LUT4 #(
		.INIT('h135f)
	) name4468 (
		\h1rdt3_dma[13]_pad ,
		\h1rdt6_dma[13]_pad ,
		_w2394_,
		_w2413_,
		_w6697_
	);
	LUT4 #(
		.INIT('h153f)
	) name4469 (
		\h1rdt0_br[13]_pad ,
		\h1rdt3_br[13]_pad ,
		_w2398_,
		_w2407_,
		_w6698_
	);
	LUT4 #(
		.INIT('h135f)
	) name4470 (
		\h1rdt2_br[13]_pad ,
		\h1rdt7_dma[13]_pad ,
		_w2389_,
		_w2404_,
		_w6699_
	);
	LUT4 #(
		.INIT('h8000)
	) name4471 (
		_w6696_,
		_w6697_,
		_w6698_,
		_w6699_,
		_w6700_
	);
	LUT3 #(
		.INIT('h02)
	) name4472 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		_w6701_
	);
	LUT2 #(
		.INIT('h9)
	) name4473 (
		\ctl_rf_m0end_reg/NET0131 ,
		\ctl_rf_m1end_reg/NET0131 ,
		_w6702_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		_w6701_,
		_w6702_,
		_w6703_
	);
	LUT3 #(
		.INIT('h01)
	) name4475 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		_w6704_
	);
	LUT3 #(
		.INIT('hcd)
	) name4476 (
		_w6701_,
		_w6702_,
		_w6704_,
		_w6705_
	);
	LUT3 #(
		.INIT('h70)
	) name4477 (
		_w6695_,
		_w6700_,
		_w6705_,
		_w6706_
	);
	LUT4 #(
		.INIT('h135f)
	) name4478 (
		\h1rdt1_br[21]_pad ,
		\h1rdt6_dma[21]_pad ,
		_w2400_,
		_w2413_,
		_w6707_
	);
	LUT4 #(
		.INIT('h153f)
	) name4479 (
		\h1rdt5_br[21]_pad ,
		\h1rdt5_dma[21]_pad ,
		_w2401_,
		_w2408_,
		_w6708_
	);
	LUT4 #(
		.INIT('h153f)
	) name4480 (
		\h1rdt0_br[21]_pad ,
		\h1rdt3_br[21]_pad ,
		_w2398_,
		_w2407_,
		_w6709_
	);
	LUT4 #(
		.INIT('h135f)
	) name4481 (
		\h1rdt2_br[21]_pad ,
		\h1rdt3_dma[21]_pad ,
		_w2389_,
		_w2394_,
		_w6710_
	);
	LUT4 #(
		.INIT('h8000)
	) name4482 (
		_w6707_,
		_w6708_,
		_w6709_,
		_w6710_,
		_w6711_
	);
	LUT4 #(
		.INIT('h135f)
	) name4483 (
		\h1rdt1_dma[21]_pad ,
		\h1rdt2_dma[21]_pad ,
		_w2395_,
		_w2410_,
		_w6712_
	);
	LUT4 #(
		.INIT('h153f)
	) name4484 (
		\h1rdt4_br[21]_pad ,
		\h1rdt6_br[21]_pad ,
		_w2392_,
		_w2405_,
		_w6713_
	);
	LUT4 #(
		.INIT('h153f)
	) name4485 (
		\h1rdt4_dma[21]_pad ,
		\h1rdt7_br[21]_pad ,
		_w2391_,
		_w2411_,
		_w6714_
	);
	LUT4 #(
		.INIT('h153f)
	) name4486 (
		\h1rdt0_dma[21]_pad ,
		\h1rdt7_dma[21]_pad ,
		_w2404_,
		_w2414_,
		_w6715_
	);
	LUT4 #(
		.INIT('h8000)
	) name4487 (
		_w6712_,
		_w6713_,
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT3 #(
		.INIT('h10)
	) name4488 (
		_w6701_,
		_w6702_,
		_w6704_,
		_w6717_
	);
	LUT3 #(
		.INIT('h70)
	) name4489 (
		_w6711_,
		_w6716_,
		_w6717_,
		_w6718_
	);
	LUT4 #(
		.INIT('h153f)
	) name4490 (
		\h1rdt1_br[29]_pad ,
		\h1rdt2_br[29]_pad ,
		_w2389_,
		_w2400_,
		_w6719_
	);
	LUT4 #(
		.INIT('h153f)
	) name4491 (
		\h1rdt4_dma[29]_pad ,
		\h1rdt6_br[29]_pad ,
		_w2392_,
		_w2411_,
		_w6720_
	);
	LUT4 #(
		.INIT('h153f)
	) name4492 (
		\h1rdt1_dma[29]_pad ,
		\h1rdt7_br[29]_pad ,
		_w2391_,
		_w2395_,
		_w6721_
	);
	LUT4 #(
		.INIT('h153f)
	) name4493 (
		\h1rdt0_dma[29]_pad ,
		\h1rdt4_br[29]_pad ,
		_w2405_,
		_w2414_,
		_w6722_
	);
	LUT4 #(
		.INIT('h8000)
	) name4494 (
		_w6719_,
		_w6720_,
		_w6721_,
		_w6722_,
		_w6723_
	);
	LUT4 #(
		.INIT('h135f)
	) name4495 (
		\h1rdt3_dma[29]_pad ,
		\h1rdt7_dma[29]_pad ,
		_w2394_,
		_w2404_,
		_w6724_
	);
	LUT4 #(
		.INIT('h153f)
	) name4496 (
		\h1rdt2_dma[29]_pad ,
		\h1rdt5_dma[29]_pad ,
		_w2401_,
		_w2410_,
		_w6725_
	);
	LUT4 #(
		.INIT('h135f)
	) name4497 (
		\h1rdt3_br[29]_pad ,
		\h1rdt6_dma[29]_pad ,
		_w2398_,
		_w2413_,
		_w6726_
	);
	LUT4 #(
		.INIT('h135f)
	) name4498 (
		\h1rdt0_br[29]_pad ,
		\h1rdt5_br[29]_pad ,
		_w2407_,
		_w2408_,
		_w6727_
	);
	LUT4 #(
		.INIT('h8000)
	) name4499 (
		_w6724_,
		_w6725_,
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT3 #(
		.INIT('h2a)
	) name4500 (
		_w6703_,
		_w6723_,
		_w6728_,
		_w6729_
	);
	LUT3 #(
		.INIT('hfe)
	) name4501 (
		_w6706_,
		_w6718_,
		_w6729_,
		_w6730_
	);
	LUT4 #(
		.INIT('h153f)
	) name4502 (
		\h1rdt0_br[14]_pad ,
		\h1rdt2_br[14]_pad ,
		_w2389_,
		_w2407_,
		_w6731_
	);
	LUT4 #(
		.INIT('h153f)
	) name4503 (
		\h1rdt4_dma[14]_pad ,
		\h1rdt6_br[14]_pad ,
		_w2392_,
		_w2411_,
		_w6732_
	);
	LUT4 #(
		.INIT('h153f)
	) name4504 (
		\h1rdt1_br[14]_pad ,
		\h1rdt7_br[14]_pad ,
		_w2391_,
		_w2400_,
		_w6733_
	);
	LUT4 #(
		.INIT('h153f)
	) name4505 (
		\h1rdt0_dma[14]_pad ,
		\h1rdt7_dma[14]_pad ,
		_w2404_,
		_w2414_,
		_w6734_
	);
	LUT4 #(
		.INIT('h8000)
	) name4506 (
		_w6731_,
		_w6732_,
		_w6733_,
		_w6734_,
		_w6735_
	);
	LUT4 #(
		.INIT('h135f)
	) name4507 (
		\h1rdt4_br[14]_pad ,
		\h1rdt5_br[14]_pad ,
		_w2405_,
		_w2408_,
		_w6736_
	);
	LUT4 #(
		.INIT('h135f)
	) name4508 (
		\h1rdt1_dma[14]_pad ,
		\h1rdt2_dma[14]_pad ,
		_w2395_,
		_w2410_,
		_w6737_
	);
	LUT4 #(
		.INIT('h153f)
	) name4509 (
		\h1rdt3_br[14]_pad ,
		\h1rdt3_dma[14]_pad ,
		_w2394_,
		_w2398_,
		_w6738_
	);
	LUT4 #(
		.INIT('h135f)
	) name4510 (
		\h1rdt5_dma[14]_pad ,
		\h1rdt6_dma[14]_pad ,
		_w2401_,
		_w2413_,
		_w6739_
	);
	LUT4 #(
		.INIT('h8000)
	) name4511 (
		_w6736_,
		_w6737_,
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT3 #(
		.INIT('h2a)
	) name4512 (
		_w6705_,
		_w6735_,
		_w6740_,
		_w6741_
	);
	LUT4 #(
		.INIT('h135f)
	) name4513 (
		\h1rdt1_dma[22]_pad ,
		\h1rdt5_br[22]_pad ,
		_w2395_,
		_w2408_,
		_w6742_
	);
	LUT4 #(
		.INIT('h153f)
	) name4514 (
		\h1rdt4_dma[22]_pad ,
		\h1rdt7_dma[22]_pad ,
		_w2404_,
		_w2411_,
		_w6743_
	);
	LUT4 #(
		.INIT('h153f)
	) name4515 (
		\h1rdt3_br[22]_pad ,
		\h1rdt3_dma[22]_pad ,
		_w2394_,
		_w2398_,
		_w6744_
	);
	LUT4 #(
		.INIT('h153f)
	) name4516 (
		\h1rdt0_dma[22]_pad ,
		\h1rdt6_dma[22]_pad ,
		_w2413_,
		_w2414_,
		_w6745_
	);
	LUT4 #(
		.INIT('h8000)
	) name4517 (
		_w6742_,
		_w6743_,
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT4 #(
		.INIT('h153f)
	) name4518 (
		\h1rdt0_br[22]_pad ,
		\h1rdt6_br[22]_pad ,
		_w2392_,
		_w2407_,
		_w6747_
	);
	LUT4 #(
		.INIT('h153f)
	) name4519 (
		\h1rdt4_br[22]_pad ,
		\h1rdt5_dma[22]_pad ,
		_w2401_,
		_w2405_,
		_w6748_
	);
	LUT4 #(
		.INIT('h135f)
	) name4520 (
		\h1rdt2_br[22]_pad ,
		\h1rdt7_br[22]_pad ,
		_w2389_,
		_w2391_,
		_w6749_
	);
	LUT4 #(
		.INIT('h135f)
	) name4521 (
		\h1rdt1_br[22]_pad ,
		\h1rdt2_dma[22]_pad ,
		_w2400_,
		_w2410_,
		_w6750_
	);
	LUT4 #(
		.INIT('h8000)
	) name4522 (
		_w6747_,
		_w6748_,
		_w6749_,
		_w6750_,
		_w6751_
	);
	LUT3 #(
		.INIT('h2a)
	) name4523 (
		_w6717_,
		_w6746_,
		_w6751_,
		_w6752_
	);
	LUT4 #(
		.INIT('h153f)
	) name4524 (
		\h1rdt0_br[30]_pad ,
		\h1rdt5_dma[30]_pad ,
		_w2401_,
		_w2407_,
		_w6753_
	);
	LUT4 #(
		.INIT('h153f)
	) name4525 (
		\h1rdt0_dma[30]_pad ,
		\h1rdt6_br[30]_pad ,
		_w2392_,
		_w2414_,
		_w6754_
	);
	LUT4 #(
		.INIT('h153f)
	) name4526 (
		\h1rdt5_br[30]_pad ,
		\h1rdt7_br[30]_pad ,
		_w2391_,
		_w2408_,
		_w6755_
	);
	LUT4 #(
		.INIT('h135f)
	) name4527 (
		\h1rdt4_br[30]_pad ,
		\h1rdt4_dma[30]_pad ,
		_w2405_,
		_w2411_,
		_w6756_
	);
	LUT4 #(
		.INIT('h8000)
	) name4528 (
		_w6753_,
		_w6754_,
		_w6755_,
		_w6756_,
		_w6757_
	);
	LUT4 #(
		.INIT('h153f)
	) name4529 (
		\h1rdt6_dma[30]_pad ,
		\h1rdt7_dma[30]_pad ,
		_w2404_,
		_w2413_,
		_w6758_
	);
	LUT4 #(
		.INIT('h153f)
	) name4530 (
		\h1rdt1_br[30]_pad ,
		\h1rdt2_br[30]_pad ,
		_w2389_,
		_w2400_,
		_w6759_
	);
	LUT4 #(
		.INIT('h153f)
	) name4531 (
		\h1rdt2_dma[30]_pad ,
		\h1rdt3_br[30]_pad ,
		_w2398_,
		_w2410_,
		_w6760_
	);
	LUT4 #(
		.INIT('h153f)
	) name4532 (
		\h1rdt1_dma[30]_pad ,
		\h1rdt3_dma[30]_pad ,
		_w2394_,
		_w2395_,
		_w6761_
	);
	LUT4 #(
		.INIT('h8000)
	) name4533 (
		_w6758_,
		_w6759_,
		_w6760_,
		_w6761_,
		_w6762_
	);
	LUT3 #(
		.INIT('h2a)
	) name4534 (
		_w6703_,
		_w6757_,
		_w6762_,
		_w6763_
	);
	LUT3 #(
		.INIT('hfe)
	) name4535 (
		_w6741_,
		_w6752_,
		_w6763_,
		_w6764_
	);
	LUT4 #(
		.INIT('h153f)
	) name4536 (
		\h1rdt4_br[15]_pad ,
		\h1rdt6_br[15]_pad ,
		_w2392_,
		_w2405_,
		_w6765_
	);
	LUT4 #(
		.INIT('h153f)
	) name4537 (
		\h1rdt1_dma[15]_pad ,
		\h1rdt2_br[15]_pad ,
		_w2389_,
		_w2395_,
		_w6766_
	);
	LUT4 #(
		.INIT('h153f)
	) name4538 (
		\h1rdt0_dma[15]_pad ,
		\h1rdt7_br[15]_pad ,
		_w2391_,
		_w2414_,
		_w6767_
	);
	LUT4 #(
		.INIT('h135f)
	) name4539 (
		\h1rdt1_br[15]_pad ,
		\h1rdt2_dma[15]_pad ,
		_w2400_,
		_w2410_,
		_w6768_
	);
	LUT4 #(
		.INIT('h8000)
	) name4540 (
		_w6765_,
		_w6766_,
		_w6767_,
		_w6768_,
		_w6769_
	);
	LUT4 #(
		.INIT('h135f)
	) name4541 (
		\h1rdt5_br[15]_pad ,
		\h1rdt6_dma[15]_pad ,
		_w2408_,
		_w2413_,
		_w6770_
	);
	LUT4 #(
		.INIT('h153f)
	) name4542 (
		\h1rdt4_dma[15]_pad ,
		\h1rdt7_dma[15]_pad ,
		_w2404_,
		_w2411_,
		_w6771_
	);
	LUT4 #(
		.INIT('h135f)
	) name4543 (
		\h1rdt3_br[15]_pad ,
		\h1rdt5_dma[15]_pad ,
		_w2398_,
		_w2401_,
		_w6772_
	);
	LUT4 #(
		.INIT('h153f)
	) name4544 (
		\h1rdt0_br[15]_pad ,
		\h1rdt3_dma[15]_pad ,
		_w2394_,
		_w2407_,
		_w6773_
	);
	LUT4 #(
		.INIT('h8000)
	) name4545 (
		_w6770_,
		_w6771_,
		_w6772_,
		_w6773_,
		_w6774_
	);
	LUT3 #(
		.INIT('h2a)
	) name4546 (
		_w6705_,
		_w6769_,
		_w6774_,
		_w6775_
	);
	LUT4 #(
		.INIT('h135f)
	) name4547 (
		\h1rdt3_dma[23]_pad ,
		\h1rdt5_dma[23]_pad ,
		_w2394_,
		_w2401_,
		_w6776_
	);
	LUT4 #(
		.INIT('h153f)
	) name4548 (
		\h1rdt0_dma[23]_pad ,
		\h1rdt5_br[23]_pad ,
		_w2408_,
		_w2414_,
		_w6777_
	);
	LUT4 #(
		.INIT('h135f)
	) name4549 (
		\h1rdt3_br[23]_pad ,
		\h1rdt4_br[23]_pad ,
		_w2398_,
		_w2405_,
		_w6778_
	);
	LUT4 #(
		.INIT('h135f)
	) name4550 (
		\h1rdt1_dma[23]_pad ,
		\h1rdt4_dma[23]_pad ,
		_w2395_,
		_w2411_,
		_w6779_
	);
	LUT4 #(
		.INIT('h8000)
	) name4551 (
		_w6776_,
		_w6777_,
		_w6778_,
		_w6779_,
		_w6780_
	);
	LUT4 #(
		.INIT('h135f)
	) name4552 (
		\h1rdt0_br[23]_pad ,
		\h1rdt6_dma[23]_pad ,
		_w2407_,
		_w2413_,
		_w6781_
	);
	LUT4 #(
		.INIT('h153f)
	) name4553 (
		\h1rdt2_dma[23]_pad ,
		\h1rdt7_dma[23]_pad ,
		_w2404_,
		_w2410_,
		_w6782_
	);
	LUT4 #(
		.INIT('h153f)
	) name4554 (
		\h1rdt1_br[23]_pad ,
		\h1rdt7_br[23]_pad ,
		_w2391_,
		_w2400_,
		_w6783_
	);
	LUT4 #(
		.INIT('h135f)
	) name4555 (
		\h1rdt2_br[23]_pad ,
		\h1rdt6_br[23]_pad ,
		_w2389_,
		_w2392_,
		_w6784_
	);
	LUT4 #(
		.INIT('h8000)
	) name4556 (
		_w6781_,
		_w6782_,
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT3 #(
		.INIT('h2a)
	) name4557 (
		_w6717_,
		_w6780_,
		_w6785_,
		_w6786_
	);
	LUT4 #(
		.INIT('h153f)
	) name4558 (
		\h1rdt0_br[31]_pad ,
		\h1rdt5_dma[31]_pad ,
		_w2401_,
		_w2407_,
		_w6787_
	);
	LUT4 #(
		.INIT('h153f)
	) name4559 (
		\h1rdt1_br[31]_pad ,
		\h1rdt6_br[31]_pad ,
		_w2392_,
		_w2400_,
		_w6788_
	);
	LUT4 #(
		.INIT('h135f)
	) name4560 (
		\h1rdt7_br[31]_pad ,
		\h1rdt7_dma[31]_pad ,
		_w2391_,
		_w2404_,
		_w6789_
	);
	LUT4 #(
		.INIT('h135f)
	) name4561 (
		\h1rdt2_br[31]_pad ,
		\h1rdt4_br[31]_pad ,
		_w2389_,
		_w2405_,
		_w6790_
	);
	LUT4 #(
		.INIT('h8000)
	) name4562 (
		_w6787_,
		_w6788_,
		_w6789_,
		_w6790_,
		_w6791_
	);
	LUT4 #(
		.INIT('h153f)
	) name4563 (
		\h1rdt0_dma[31]_pad ,
		\h1rdt4_dma[31]_pad ,
		_w2411_,
		_w2414_,
		_w6792_
	);
	LUT4 #(
		.INIT('h135f)
	) name4564 (
		\h1rdt5_br[31]_pad ,
		\h1rdt6_dma[31]_pad ,
		_w2408_,
		_w2413_,
		_w6793_
	);
	LUT4 #(
		.INIT('h153f)
	) name4565 (
		\h1rdt2_dma[31]_pad ,
		\h1rdt3_br[31]_pad ,
		_w2398_,
		_w2410_,
		_w6794_
	);
	LUT4 #(
		.INIT('h153f)
	) name4566 (
		\h1rdt1_dma[31]_pad ,
		\h1rdt3_dma[31]_pad ,
		_w2394_,
		_w2395_,
		_w6795_
	);
	LUT4 #(
		.INIT('h8000)
	) name4567 (
		_w6792_,
		_w6793_,
		_w6794_,
		_w6795_,
		_w6796_
	);
	LUT3 #(
		.INIT('h2a)
	) name4568 (
		_w6703_,
		_w6791_,
		_w6796_,
		_w6797_
	);
	LUT3 #(
		.INIT('hfe)
	) name4569 (
		_w6775_,
		_w6786_,
		_w6797_,
		_w6798_
	);
	LUT4 #(
		.INIT('h135f)
	) name4570 (
		\h1rdt2_br[16]_pad ,
		\h1rdt6_dma[16]_pad ,
		_w2389_,
		_w2413_,
		_w6799_
	);
	LUT4 #(
		.INIT('h153f)
	) name4571 (
		\h1rdt0_dma[16]_pad ,
		\h1rdt5_br[16]_pad ,
		_w2408_,
		_w2414_,
		_w6800_
	);
	LUT4 #(
		.INIT('h153f)
	) name4572 (
		\h1rdt3_br[16]_pad ,
		\h1rdt6_br[16]_pad ,
		_w2392_,
		_w2398_,
		_w6801_
	);
	LUT4 #(
		.INIT('h135f)
	) name4573 (
		\h1rdt1_br[16]_pad ,
		\h1rdt4_dma[16]_pad ,
		_w2400_,
		_w2411_,
		_w6802_
	);
	LUT4 #(
		.INIT('h8000)
	) name4574 (
		_w6799_,
		_w6800_,
		_w6801_,
		_w6802_,
		_w6803_
	);
	LUT4 #(
		.INIT('h135f)
	) name4575 (
		\h1rdt3_dma[16]_pad ,
		\h1rdt5_dma[16]_pad ,
		_w2394_,
		_w2401_,
		_w6804_
	);
	LUT4 #(
		.INIT('h135f)
	) name4576 (
		\h1rdt1_dma[16]_pad ,
		\h1rdt2_dma[16]_pad ,
		_w2395_,
		_w2410_,
		_w6805_
	);
	LUT4 #(
		.INIT('h153f)
	) name4577 (
		\h1rdt4_br[16]_pad ,
		\h1rdt7_br[16]_pad ,
		_w2391_,
		_w2405_,
		_w6806_
	);
	LUT4 #(
		.INIT('h153f)
	) name4578 (
		\h1rdt0_br[16]_pad ,
		\h1rdt7_dma[16]_pad ,
		_w2404_,
		_w2407_,
		_w6807_
	);
	LUT4 #(
		.INIT('h8000)
	) name4579 (
		_w6804_,
		_w6805_,
		_w6806_,
		_w6807_,
		_w6808_
	);
	LUT3 #(
		.INIT('h2a)
	) name4580 (
		_w6705_,
		_w6803_,
		_w6808_,
		_w6809_
	);
	LUT4 #(
		.INIT('h135f)
	) name4581 (
		\h1rdt1_br[8]_pad ,
		\h1rdt5_br[8]_pad ,
		_w2400_,
		_w2408_,
		_w6810_
	);
	LUT4 #(
		.INIT('h153f)
	) name4582 (
		\h1rdt0_dma[8]_pad ,
		\h1rdt6_dma[8]_pad ,
		_w2413_,
		_w2414_,
		_w6811_
	);
	LUT4 #(
		.INIT('h153f)
	) name4583 (
		\h1rdt0_br[8]_pad ,
		\h1rdt3_br[8]_pad ,
		_w2398_,
		_w2407_,
		_w6812_
	);
	LUT4 #(
		.INIT('h153f)
	) name4584 (
		\h1rdt4_dma[8]_pad ,
		\h1rdt7_dma[8]_pad ,
		_w2404_,
		_w2411_,
		_w6813_
	);
	LUT4 #(
		.INIT('h8000)
	) name4585 (
		_w6810_,
		_w6811_,
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT4 #(
		.INIT('h135f)
	) name4586 (
		\h1rdt1_dma[8]_pad ,
		\h1rdt2_dma[8]_pad ,
		_w2395_,
		_w2410_,
		_w6815_
	);
	LUT4 #(
		.INIT('h135f)
	) name4587 (
		\h1rdt3_dma[8]_pad ,
		\h1rdt5_dma[8]_pad ,
		_w2394_,
		_w2401_,
		_w6816_
	);
	LUT4 #(
		.INIT('h153f)
	) name4588 (
		\h1rdt6_br[8]_pad ,
		\h1rdt7_br[8]_pad ,
		_w2391_,
		_w2392_,
		_w6817_
	);
	LUT4 #(
		.INIT('h135f)
	) name4589 (
		\h1rdt2_br[8]_pad ,
		\h1rdt4_br[8]_pad ,
		_w2389_,
		_w2405_,
		_w6818_
	);
	LUT4 #(
		.INIT('h8000)
	) name4590 (
		_w6815_,
		_w6816_,
		_w6817_,
		_w6818_,
		_w6819_
	);
	LUT3 #(
		.INIT('h2a)
	) name4591 (
		_w6717_,
		_w6814_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('h153f)
	) name4592 (
		\h1rdt0_br[0]_pad ,
		\h1rdt5_dma[0]_pad ,
		_w2401_,
		_w2407_,
		_w6821_
	);
	LUT4 #(
		.INIT('h153f)
	) name4593 (
		\h1rdt0_dma[0]_pad ,
		\h1rdt4_br[0]_pad ,
		_w2405_,
		_w2414_,
		_w6822_
	);
	LUT4 #(
		.INIT('h135f)
	) name4594 (
		\h1rdt2_br[0]_pad ,
		\h1rdt7_br[0]_pad ,
		_w2389_,
		_w2391_,
		_w6823_
	);
	LUT4 #(
		.INIT('h153f)
	) name4595 (
		\h1rdt4_dma[0]_pad ,
		\h1rdt6_br[0]_pad ,
		_w2392_,
		_w2411_,
		_w6824_
	);
	LUT4 #(
		.INIT('h8000)
	) name4596 (
		_w6821_,
		_w6822_,
		_w6823_,
		_w6824_,
		_w6825_
	);
	LUT4 #(
		.INIT('h153f)
	) name4597 (
		\h1rdt6_dma[0]_pad ,
		\h1rdt7_dma[0]_pad ,
		_w2404_,
		_w2413_,
		_w6826_
	);
	LUT4 #(
		.INIT('h135f)
	) name4598 (
		\h1rdt1_br[0]_pad ,
		\h1rdt5_br[0]_pad ,
		_w2400_,
		_w2408_,
		_w6827_
	);
	LUT4 #(
		.INIT('h153f)
	) name4599 (
		\h1rdt2_dma[0]_pad ,
		\h1rdt3_br[0]_pad ,
		_w2398_,
		_w2410_,
		_w6828_
	);
	LUT4 #(
		.INIT('h153f)
	) name4600 (
		\h1rdt1_dma[0]_pad ,
		\h1rdt3_dma[0]_pad ,
		_w2394_,
		_w2395_,
		_w6829_
	);
	LUT4 #(
		.INIT('h8000)
	) name4601 (
		_w6826_,
		_w6827_,
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT3 #(
		.INIT('h2a)
	) name4602 (
		_w6703_,
		_w6825_,
		_w6830_,
		_w6831_
	);
	LUT3 #(
		.INIT('hfe)
	) name4603 (
		_w6809_,
		_w6820_,
		_w6831_,
		_w6832_
	);
	LUT4 #(
		.INIT('h135f)
	) name4604 (
		\h1rdt2_br[17]_pad ,
		\h1rdt6_dma[17]_pad ,
		_w2389_,
		_w2413_,
		_w6833_
	);
	LUT4 #(
		.INIT('h153f)
	) name4605 (
		\h1rdt5_br[17]_pad ,
		\h1rdt5_dma[17]_pad ,
		_w2401_,
		_w2408_,
		_w6834_
	);
	LUT4 #(
		.INIT('h153f)
	) name4606 (
		\h1rdt2_dma[17]_pad ,
		\h1rdt3_br[17]_pad ,
		_w2398_,
		_w2410_,
		_w6835_
	);
	LUT4 #(
		.INIT('h135f)
	) name4607 (
		\h1rdt3_dma[17]_pad ,
		\h1rdt7_dma[17]_pad ,
		_w2394_,
		_w2404_,
		_w6836_
	);
	LUT4 #(
		.INIT('h8000)
	) name4608 (
		_w6833_,
		_w6834_,
		_w6835_,
		_w6836_,
		_w6837_
	);
	LUT4 #(
		.INIT('h153f)
	) name4609 (
		\h1rdt4_br[17]_pad ,
		\h1rdt6_br[17]_pad ,
		_w2392_,
		_w2405_,
		_w6838_
	);
	LUT4 #(
		.INIT('h153f)
	) name4610 (
		\h1rdt0_br[17]_pad ,
		\h1rdt1_dma[17]_pad ,
		_w2395_,
		_w2407_,
		_w6839_
	);
	LUT4 #(
		.INIT('h153f)
	) name4611 (
		\h1rdt4_dma[17]_pad ,
		\h1rdt7_br[17]_pad ,
		_w2391_,
		_w2411_,
		_w6840_
	);
	LUT4 #(
		.INIT('h153f)
	) name4612 (
		\h1rdt0_dma[17]_pad ,
		\h1rdt1_br[17]_pad ,
		_w2400_,
		_w2414_,
		_w6841_
	);
	LUT4 #(
		.INIT('h8000)
	) name4613 (
		_w6838_,
		_w6839_,
		_w6840_,
		_w6841_,
		_w6842_
	);
	LUT3 #(
		.INIT('h2a)
	) name4614 (
		_w6705_,
		_w6837_,
		_w6842_,
		_w6843_
	);
	LUT4 #(
		.INIT('h135f)
	) name4615 (
		\h1rdt1_dma[9]_pad ,
		\h1rdt2_dma[9]_pad ,
		_w2395_,
		_w2410_,
		_w6844_
	);
	LUT4 #(
		.INIT('h135f)
	) name4616 (
		\h1rdt3_dma[9]_pad ,
		\h1rdt4_dma[9]_pad ,
		_w2394_,
		_w2411_,
		_w6845_
	);
	LUT4 #(
		.INIT('h153f)
	) name4617 (
		\h1rdt5_br[9]_pad ,
		\h1rdt7_br[9]_pad ,
		_w2391_,
		_w2408_,
		_w6846_
	);
	LUT4 #(
		.INIT('h153f)
	) name4618 (
		\h1rdt0_dma[9]_pad ,
		\h1rdt5_dma[9]_pad ,
		_w2401_,
		_w2414_,
		_w6847_
	);
	LUT4 #(
		.INIT('h8000)
	) name4619 (
		_w6844_,
		_w6845_,
		_w6846_,
		_w6847_,
		_w6848_
	);
	LUT4 #(
		.INIT('h153f)
	) name4620 (
		\h1rdt6_dma[9]_pad ,
		\h1rdt7_dma[9]_pad ,
		_w2404_,
		_w2413_,
		_w6849_
	);
	LUT4 #(
		.INIT('h153f)
	) name4621 (
		\h1rdt1_br[9]_pad ,
		\h1rdt2_br[9]_pad ,
		_w2389_,
		_w2400_,
		_w6850_
	);
	LUT4 #(
		.INIT('h153f)
	) name4622 (
		\h1rdt0_br[9]_pad ,
		\h1rdt3_br[9]_pad ,
		_w2398_,
		_w2407_,
		_w6851_
	);
	LUT4 #(
		.INIT('h153f)
	) name4623 (
		\h1rdt4_br[9]_pad ,
		\h1rdt6_br[9]_pad ,
		_w2392_,
		_w2405_,
		_w6852_
	);
	LUT4 #(
		.INIT('h8000)
	) name4624 (
		_w6849_,
		_w6850_,
		_w6851_,
		_w6852_,
		_w6853_
	);
	LUT3 #(
		.INIT('h2a)
	) name4625 (
		_w6717_,
		_w6848_,
		_w6853_,
		_w6854_
	);
	LUT4 #(
		.INIT('h135f)
	) name4626 (
		\h1rdt1_dma[1]_pad ,
		\h1rdt2_dma[1]_pad ,
		_w2395_,
		_w2410_,
		_w6855_
	);
	LUT4 #(
		.INIT('h135f)
	) name4627 (
		\h1rdt3_dma[1]_pad ,
		\h1rdt6_dma[1]_pad ,
		_w2394_,
		_w2413_,
		_w6856_
	);
	LUT4 #(
		.INIT('h153f)
	) name4628 (
		\h1rdt0_dma[1]_pad ,
		\h1rdt7_br[1]_pad ,
		_w2391_,
		_w2414_,
		_w6857_
	);
	LUT4 #(
		.INIT('h135f)
	) name4629 (
		\h1rdt5_dma[1]_pad ,
		\h1rdt7_dma[1]_pad ,
		_w2401_,
		_w2404_,
		_w6858_
	);
	LUT4 #(
		.INIT('h8000)
	) name4630 (
		_w6855_,
		_w6856_,
		_w6857_,
		_w6858_,
		_w6859_
	);
	LUT4 #(
		.INIT('h153f)
	) name4631 (
		\h1rdt1_br[1]_pad ,
		\h1rdt2_br[1]_pad ,
		_w2389_,
		_w2400_,
		_w6860_
	);
	LUT4 #(
		.INIT('h153f)
	) name4632 (
		\h1rdt4_dma[1]_pad ,
		\h1rdt5_br[1]_pad ,
		_w2408_,
		_w2411_,
		_w6861_
	);
	LUT4 #(
		.INIT('h153f)
	) name4633 (
		\h1rdt0_br[1]_pad ,
		\h1rdt3_br[1]_pad ,
		_w2398_,
		_w2407_,
		_w6862_
	);
	LUT4 #(
		.INIT('h153f)
	) name4634 (
		\h1rdt4_br[1]_pad ,
		\h1rdt6_br[1]_pad ,
		_w2392_,
		_w2405_,
		_w6863_
	);
	LUT4 #(
		.INIT('h8000)
	) name4635 (
		_w6860_,
		_w6861_,
		_w6862_,
		_w6863_,
		_w6864_
	);
	LUT3 #(
		.INIT('h2a)
	) name4636 (
		_w6703_,
		_w6859_,
		_w6864_,
		_w6865_
	);
	LUT3 #(
		.INIT('hfe)
	) name4637 (
		_w6843_,
		_w6854_,
		_w6865_,
		_w6866_
	);
	LUT4 #(
		.INIT('h135f)
	) name4638 (
		\h1rdt1_br[18]_pad ,
		\h1rdt7_dma[18]_pad ,
		_w2400_,
		_w2404_,
		_w6867_
	);
	LUT4 #(
		.INIT('h153f)
	) name4639 (
		\h1rdt0_dma[18]_pad ,
		\h1rdt5_br[18]_pad ,
		_w2408_,
		_w2414_,
		_w6868_
	);
	LUT4 #(
		.INIT('h153f)
	) name4640 (
		\h1rdt3_br[18]_pad ,
		\h1rdt6_br[18]_pad ,
		_w2392_,
		_w2398_,
		_w6869_
	);
	LUT4 #(
		.INIT('h135f)
	) name4641 (
		\h1rdt4_dma[18]_pad ,
		\h1rdt6_dma[18]_pad ,
		_w2411_,
		_w2413_,
		_w6870_
	);
	LUT4 #(
		.INIT('h8000)
	) name4642 (
		_w6867_,
		_w6868_,
		_w6869_,
		_w6870_,
		_w6871_
	);
	LUT4 #(
		.INIT('h135f)
	) name4643 (
		\h1rdt3_dma[18]_pad ,
		\h1rdt5_dma[18]_pad ,
		_w2394_,
		_w2401_,
		_w6872_
	);
	LUT4 #(
		.INIT('h135f)
	) name4644 (
		\h1rdt1_dma[18]_pad ,
		\h1rdt2_dma[18]_pad ,
		_w2395_,
		_w2410_,
		_w6873_
	);
	LUT4 #(
		.INIT('h153f)
	) name4645 (
		\h1rdt4_br[18]_pad ,
		\h1rdt7_br[18]_pad ,
		_w2391_,
		_w2405_,
		_w6874_
	);
	LUT4 #(
		.INIT('h153f)
	) name4646 (
		\h1rdt0_br[18]_pad ,
		\h1rdt2_br[18]_pad ,
		_w2389_,
		_w2407_,
		_w6875_
	);
	LUT4 #(
		.INIT('h8000)
	) name4647 (
		_w6872_,
		_w6873_,
		_w6874_,
		_w6875_,
		_w6876_
	);
	LUT3 #(
		.INIT('h2a)
	) name4648 (
		_w6705_,
		_w6871_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('h153f)
	) name4649 (
		\h1rdt0_dma[10]_pad ,
		\h1rdt2_dma[10]_pad ,
		_w2410_,
		_w2414_,
		_w6878_
	);
	LUT4 #(
		.INIT('h153f)
	) name4650 (
		\h1rdt1_dma[10]_pad ,
		\h1rdt3_dma[10]_pad ,
		_w2394_,
		_w2395_,
		_w6879_
	);
	LUT4 #(
		.INIT('h153f)
	) name4651 (
		\h1rdt3_br[10]_pad ,
		\h1rdt6_br[10]_pad ,
		_w2392_,
		_w2398_,
		_w6880_
	);
	LUT4 #(
		.INIT('h153f)
	) name4652 (
		\h1rdt4_br[10]_pad ,
		\h1rdt5_dma[10]_pad ,
		_w2401_,
		_w2405_,
		_w6881_
	);
	LUT4 #(
		.INIT('h8000)
	) name4653 (
		_w6878_,
		_w6879_,
		_w6880_,
		_w6881_,
		_w6882_
	);
	LUT4 #(
		.INIT('h153f)
	) name4654 (
		\h1rdt6_dma[10]_pad ,
		\h1rdt7_dma[10]_pad ,
		_w2404_,
		_w2413_,
		_w6883_
	);
	LUT4 #(
		.INIT('h135f)
	) name4655 (
		\h1rdt0_br[10]_pad ,
		\h1rdt5_br[10]_pad ,
		_w2407_,
		_w2408_,
		_w6884_
	);
	LUT4 #(
		.INIT('h135f)
	) name4656 (
		\h1rdt2_br[10]_pad ,
		\h1rdt7_br[10]_pad ,
		_w2389_,
		_w2391_,
		_w6885_
	);
	LUT4 #(
		.INIT('h135f)
	) name4657 (
		\h1rdt1_br[10]_pad ,
		\h1rdt4_dma[10]_pad ,
		_w2400_,
		_w2411_,
		_w6886_
	);
	LUT4 #(
		.INIT('h8000)
	) name4658 (
		_w6883_,
		_w6884_,
		_w6885_,
		_w6886_,
		_w6887_
	);
	LUT3 #(
		.INIT('h2a)
	) name4659 (
		_w6717_,
		_w6882_,
		_w6887_,
		_w6888_
	);
	LUT4 #(
		.INIT('h135f)
	) name4660 (
		\h1rdt3_dma[2]_pad ,
		\h1rdt5_dma[2]_pad ,
		_w2394_,
		_w2401_,
		_w6889_
	);
	LUT4 #(
		.INIT('h153f)
	) name4661 (
		\h1rdt2_dma[2]_pad ,
		\h1rdt6_br[2]_pad ,
		_w2392_,
		_w2410_,
		_w6890_
	);
	LUT4 #(
		.INIT('h135f)
	) name4662 (
		\h1rdt2_br[2]_pad ,
		\h1rdt7_br[2]_pad ,
		_w2389_,
		_w2391_,
		_w6891_
	);
	LUT4 #(
		.INIT('h135f)
	) name4663 (
		\h1rdt4_br[2]_pad ,
		\h1rdt6_dma[2]_pad ,
		_w2405_,
		_w2413_,
		_w6892_
	);
	LUT4 #(
		.INIT('h8000)
	) name4664 (
		_w6889_,
		_w6890_,
		_w6891_,
		_w6892_,
		_w6893_
	);
	LUT4 #(
		.INIT('h153f)
	) name4665 (
		\h1rdt0_dma[2]_pad ,
		\h1rdt1_dma[2]_pad ,
		_w2395_,
		_w2414_,
		_w6894_
	);
	LUT4 #(
		.INIT('h153f)
	) name4666 (
		\h1rdt4_dma[2]_pad ,
		\h1rdt7_dma[2]_pad ,
		_w2404_,
		_w2411_,
		_w6895_
	);
	LUT4 #(
		.INIT('h135f)
	) name4667 (
		\h1rdt3_br[2]_pad ,
		\h1rdt5_br[2]_pad ,
		_w2398_,
		_w2408_,
		_w6896_
	);
	LUT4 #(
		.INIT('h153f)
	) name4668 (
		\h1rdt0_br[2]_pad ,
		\h1rdt1_br[2]_pad ,
		_w2400_,
		_w2407_,
		_w6897_
	);
	LUT4 #(
		.INIT('h8000)
	) name4669 (
		_w6894_,
		_w6895_,
		_w6896_,
		_w6897_,
		_w6898_
	);
	LUT3 #(
		.INIT('h2a)
	) name4670 (
		_w6703_,
		_w6893_,
		_w6898_,
		_w6899_
	);
	LUT3 #(
		.INIT('hfe)
	) name4671 (
		_w6877_,
		_w6888_,
		_w6899_,
		_w6900_
	);
	LUT4 #(
		.INIT('h135f)
	) name4672 (
		\h1rdt2_br[19]_pad ,
		\h1rdt7_dma[19]_pad ,
		_w2389_,
		_w2404_,
		_w6901_
	);
	LUT4 #(
		.INIT('h135f)
	) name4673 (
		\h1rdt3_dma[19]_pad ,
		\h1rdt5_br[19]_pad ,
		_w2394_,
		_w2408_,
		_w6902_
	);
	LUT4 #(
		.INIT('h153f)
	) name4674 (
		\h1rdt6_br[19]_pad ,
		\h1rdt7_br[19]_pad ,
		_w2391_,
		_w2392_,
		_w6903_
	);
	LUT4 #(
		.INIT('h135f)
	) name4675 (
		\h1rdt0_br[19]_pad ,
		\h1rdt6_dma[19]_pad ,
		_w2407_,
		_w2413_,
		_w6904_
	);
	LUT4 #(
		.INIT('h8000)
	) name4676 (
		_w6901_,
		_w6902_,
		_w6903_,
		_w6904_,
		_w6905_
	);
	LUT4 #(
		.INIT('h153f)
	) name4677 (
		\h1rdt0_dma[19]_pad ,
		\h1rdt5_dma[19]_pad ,
		_w2401_,
		_w2414_,
		_w6906_
	);
	LUT4 #(
		.INIT('h135f)
	) name4678 (
		\h1rdt1_dma[19]_pad ,
		\h1rdt2_dma[19]_pad ,
		_w2395_,
		_w2410_,
		_w6907_
	);
	LUT4 #(
		.INIT('h135f)
	) name4679 (
		\h1rdt3_br[19]_pad ,
		\h1rdt4_br[19]_pad ,
		_w2398_,
		_w2405_,
		_w6908_
	);
	LUT4 #(
		.INIT('h135f)
	) name4680 (
		\h1rdt1_br[19]_pad ,
		\h1rdt4_dma[19]_pad ,
		_w2400_,
		_w2411_,
		_w6909_
	);
	LUT4 #(
		.INIT('h8000)
	) name4681 (
		_w6906_,
		_w6907_,
		_w6908_,
		_w6909_,
		_w6910_
	);
	LUT3 #(
		.INIT('h2a)
	) name4682 (
		_w6705_,
		_w6905_,
		_w6910_,
		_w6911_
	);
	LUT4 #(
		.INIT('h153f)
	) name4683 (
		\h1rdt0_br[11]_pad ,
		\h1rdt3_dma[11]_pad ,
		_w2394_,
		_w2407_,
		_w6912_
	);
	LUT4 #(
		.INIT('h135f)
	) name4684 (
		\h1rdt6_br[11]_pad ,
		\h1rdt6_dma[11]_pad ,
		_w2392_,
		_w2413_,
		_w6913_
	);
	LUT4 #(
		.INIT('h153f)
	) name4685 (
		\h1rdt0_dma[11]_pad ,
		\h1rdt7_br[11]_pad ,
		_w2391_,
		_w2414_,
		_w6914_
	);
	LUT4 #(
		.INIT('h153f)
	) name4686 (
		\h1rdt4_br[11]_pad ,
		\h1rdt7_dma[11]_pad ,
		_w2404_,
		_w2405_,
		_w6915_
	);
	LUT4 #(
		.INIT('h8000)
	) name4687 (
		_w6912_,
		_w6913_,
		_w6914_,
		_w6915_,
		_w6916_
	);
	LUT4 #(
		.INIT('h153f)
	) name4688 (
		\h1rdt1_br[11]_pad ,
		\h1rdt2_br[11]_pad ,
		_w2389_,
		_w2400_,
		_w6917_
	);
	LUT4 #(
		.INIT('h153f)
	) name4689 (
		\h1rdt4_dma[11]_pad ,
		\h1rdt5_br[11]_pad ,
		_w2408_,
		_w2411_,
		_w6918_
	);
	LUT4 #(
		.INIT('h153f)
	) name4690 (
		\h1rdt2_dma[11]_pad ,
		\h1rdt3_br[11]_pad ,
		_w2398_,
		_w2410_,
		_w6919_
	);
	LUT4 #(
		.INIT('h135f)
	) name4691 (
		\h1rdt1_dma[11]_pad ,
		\h1rdt5_dma[11]_pad ,
		_w2395_,
		_w2401_,
		_w6920_
	);
	LUT4 #(
		.INIT('h8000)
	) name4692 (
		_w6917_,
		_w6918_,
		_w6919_,
		_w6920_,
		_w6921_
	);
	LUT3 #(
		.INIT('h2a)
	) name4693 (
		_w6717_,
		_w6916_,
		_w6921_,
		_w6922_
	);
	LUT4 #(
		.INIT('h135f)
	) name4694 (
		\h1rdt3_dma[3]_pad ,
		\h1rdt5_dma[3]_pad ,
		_w2394_,
		_w2401_,
		_w6923_
	);
	LUT4 #(
		.INIT('h135f)
	) name4695 (
		\h1rdt5_br[3]_pad ,
		\h1rdt6_dma[3]_pad ,
		_w2408_,
		_w2413_,
		_w6924_
	);
	LUT4 #(
		.INIT('h153f)
	) name4696 (
		\h1rdt3_br[3]_pad ,
		\h1rdt6_br[3]_pad ,
		_w2392_,
		_w2398_,
		_w6925_
	);
	LUT4 #(
		.INIT('h153f)
	) name4697 (
		\h1rdt4_dma[3]_pad ,
		\h1rdt7_dma[3]_pad ,
		_w2404_,
		_w2411_,
		_w6926_
	);
	LUT4 #(
		.INIT('h8000)
	) name4698 (
		_w6923_,
		_w6924_,
		_w6925_,
		_w6926_,
		_w6927_
	);
	LUT4 #(
		.INIT('h153f)
	) name4699 (
		\h1rdt1_br[3]_pad ,
		\h1rdt2_br[3]_pad ,
		_w2389_,
		_w2400_,
		_w6928_
	);
	LUT4 #(
		.INIT('h153f)
	) name4700 (
		\h1rdt0_dma[3]_pad ,
		\h1rdt4_br[3]_pad ,
		_w2405_,
		_w2414_,
		_w6929_
	);
	LUT4 #(
		.INIT('h153f)
	) name4701 (
		\h1rdt0_br[3]_pad ,
		\h1rdt7_br[3]_pad ,
		_w2391_,
		_w2407_,
		_w6930_
	);
	LUT4 #(
		.INIT('h135f)
	) name4702 (
		\h1rdt1_dma[3]_pad ,
		\h1rdt2_dma[3]_pad ,
		_w2395_,
		_w2410_,
		_w6931_
	);
	LUT4 #(
		.INIT('h8000)
	) name4703 (
		_w6928_,
		_w6929_,
		_w6930_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('h2a)
	) name4704 (
		_w6703_,
		_w6927_,
		_w6932_,
		_w6933_
	);
	LUT3 #(
		.INIT('hfe)
	) name4705 (
		_w6911_,
		_w6922_,
		_w6933_,
		_w6934_
	);
	LUT4 #(
		.INIT('h153f)
	) name4706 (
		\h1rdt0_br[25]_pad ,
		\h1rdt4_br[25]_pad ,
		_w2405_,
		_w2407_,
		_w6935_
	);
	LUT4 #(
		.INIT('h135f)
	) name4707 (
		\h1rdt2_dma[25]_pad ,
		\h1rdt4_dma[25]_pad ,
		_w2410_,
		_w2411_,
		_w6936_
	);
	LUT4 #(
		.INIT('h153f)
	) name4708 (
		\h1rdt5_br[25]_pad ,
		\h1rdt7_br[25]_pad ,
		_w2391_,
		_w2408_,
		_w6937_
	);
	LUT4 #(
		.INIT('h153f)
	) name4709 (
		\h1rdt1_dma[25]_pad ,
		\h1rdt6_br[25]_pad ,
		_w2392_,
		_w2395_,
		_w6938_
	);
	LUT4 #(
		.INIT('h8000)
	) name4710 (
		_w6935_,
		_w6936_,
		_w6937_,
		_w6938_,
		_w6939_
	);
	LUT4 #(
		.INIT('h135f)
	) name4711 (
		\h1rdt2_br[25]_pad ,
		\h1rdt7_dma[25]_pad ,
		_w2389_,
		_w2404_,
		_w6940_
	);
	LUT4 #(
		.INIT('h135f)
	) name4712 (
		\h1rdt1_br[25]_pad ,
		\h1rdt6_dma[25]_pad ,
		_w2400_,
		_w2413_,
		_w6941_
	);
	LUT4 #(
		.INIT('h153f)
	) name4713 (
		\h1rdt0_dma[25]_pad ,
		\h1rdt3_br[25]_pad ,
		_w2398_,
		_w2414_,
		_w6942_
	);
	LUT4 #(
		.INIT('h135f)
	) name4714 (
		\h1rdt3_dma[25]_pad ,
		\h1rdt5_dma[25]_pad ,
		_w2394_,
		_w2401_,
		_w6943_
	);
	LUT4 #(
		.INIT('h8000)
	) name4715 (
		_w6940_,
		_w6941_,
		_w6942_,
		_w6943_,
		_w6944_
	);
	LUT3 #(
		.INIT('h2a)
	) name4716 (
		_w6717_,
		_w6939_,
		_w6944_,
		_w6945_
	);
	LUT3 #(
		.INIT('h2a)
	) name4717 (
		_w6705_,
		_w6859_,
		_w6864_,
		_w6946_
	);
	LUT3 #(
		.INIT('h2a)
	) name4718 (
		_w6703_,
		_w6837_,
		_w6842_,
		_w6947_
	);
	LUT3 #(
		.INIT('hfe)
	) name4719 (
		_w6945_,
		_w6946_,
		_w6947_,
		_w6948_
	);
	LUT4 #(
		.INIT('h135f)
	) name4720 (
		\h1rdt3_dma[20]_pad ,
		\h1rdt5_dma[20]_pad ,
		_w2394_,
		_w2401_,
		_w6949_
	);
	LUT4 #(
		.INIT('h135f)
	) name4721 (
		\h1rdt4_br[20]_pad ,
		\h1rdt4_dma[20]_pad ,
		_w2405_,
		_w2411_,
		_w6950_
	);
	LUT4 #(
		.INIT('h135f)
	) name4722 (
		\h1rdt1_dma[20]_pad ,
		\h1rdt3_br[20]_pad ,
		_w2395_,
		_w2398_,
		_w6951_
	);
	LUT4 #(
		.INIT('h153f)
	) name4723 (
		\h1rdt5_br[20]_pad ,
		\h1rdt6_br[20]_pad ,
		_w2392_,
		_w2408_,
		_w6952_
	);
	LUT4 #(
		.INIT('h8000)
	) name4724 (
		_w6949_,
		_w6950_,
		_w6951_,
		_w6952_,
		_w6953_
	);
	LUT4 #(
		.INIT('h153f)
	) name4725 (
		\h1rdt0_br[20]_pad ,
		\h1rdt2_br[20]_pad ,
		_w2389_,
		_w2407_,
		_w6954_
	);
	LUT4 #(
		.INIT('h135f)
	) name4726 (
		\h1rdt1_br[20]_pad ,
		\h1rdt2_dma[20]_pad ,
		_w2400_,
		_w2410_,
		_w6955_
	);
	LUT4 #(
		.INIT('h153f)
	) name4727 (
		\h1rdt0_dma[20]_pad ,
		\h1rdt7_br[20]_pad ,
		_w2391_,
		_w2414_,
		_w6956_
	);
	LUT4 #(
		.INIT('h153f)
	) name4728 (
		\h1rdt6_dma[20]_pad ,
		\h1rdt7_dma[20]_pad ,
		_w2404_,
		_w2413_,
		_w6957_
	);
	LUT4 #(
		.INIT('h8000)
	) name4729 (
		_w6954_,
		_w6955_,
		_w6956_,
		_w6957_,
		_w6958_
	);
	LUT3 #(
		.INIT('h2a)
	) name4730 (
		_w6705_,
		_w6953_,
		_w6958_,
		_w6959_
	);
	LUT4 #(
		.INIT('h153f)
	) name4731 (
		\h1rdt0_dma[12]_pad ,
		\h1rdt4_br[12]_pad ,
		_w2405_,
		_w2414_,
		_w6960_
	);
	LUT4 #(
		.INIT('h135f)
	) name4732 (
		\h1rdt2_dma[12]_pad ,
		\h1rdt4_dma[12]_pad ,
		_w2410_,
		_w2411_,
		_w6961_
	);
	LUT4 #(
		.INIT('h153f)
	) name4733 (
		\h1rdt3_br[12]_pad ,
		\h1rdt3_dma[12]_pad ,
		_w2394_,
		_w2398_,
		_w6962_
	);
	LUT4 #(
		.INIT('h135f)
	) name4734 (
		\h1rdt6_br[12]_pad ,
		\h1rdt6_dma[12]_pad ,
		_w2392_,
		_w2413_,
		_w6963_
	);
	LUT4 #(
		.INIT('h8000)
	) name4735 (
		_w6960_,
		_w6961_,
		_w6962_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('h153f)
	) name4736 (
		\h1rdt1_dma[12]_pad ,
		\h1rdt2_br[12]_pad ,
		_w2389_,
		_w2395_,
		_w6965_
	);
	LUT4 #(
		.INIT('h135f)
	) name4737 (
		\h1rdt1_br[12]_pad ,
		\h1rdt5_dma[12]_pad ,
		_w2400_,
		_w2401_,
		_w6966_
	);
	LUT4 #(
		.INIT('h153f)
	) name4738 (
		\h1rdt0_br[12]_pad ,
		\h1rdt7_br[12]_pad ,
		_w2391_,
		_w2407_,
		_w6967_
	);
	LUT4 #(
		.INIT('h153f)
	) name4739 (
		\h1rdt5_br[12]_pad ,
		\h1rdt7_dma[12]_pad ,
		_w2404_,
		_w2408_,
		_w6968_
	);
	LUT4 #(
		.INIT('h8000)
	) name4740 (
		_w6965_,
		_w6966_,
		_w6967_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h2a)
	) name4741 (
		_w6717_,
		_w6964_,
		_w6969_,
		_w6970_
	);
	LUT4 #(
		.INIT('h135f)
	) name4742 (
		\h1rdt5_br[4]_pad ,
		\h1rdt6_dma[4]_pad ,
		_w2408_,
		_w2413_,
		_w6971_
	);
	LUT4 #(
		.INIT('h135f)
	) name4743 (
		\h1rdt1_br[4]_pad ,
		\h1rdt5_dma[4]_pad ,
		_w2400_,
		_w2401_,
		_w6972_
	);
	LUT4 #(
		.INIT('h153f)
	) name4744 (
		\h1rdt0_br[4]_pad ,
		\h1rdt3_br[4]_pad ,
		_w2398_,
		_w2407_,
		_w6973_
	);
	LUT4 #(
		.INIT('h135f)
	) name4745 (
		\h1rdt2_br[4]_pad ,
		\h1rdt3_dma[4]_pad ,
		_w2389_,
		_w2394_,
		_w6974_
	);
	LUT4 #(
		.INIT('h8000)
	) name4746 (
		_w6971_,
		_w6972_,
		_w6973_,
		_w6974_,
		_w6975_
	);
	LUT4 #(
		.INIT('h135f)
	) name4747 (
		\h1rdt1_dma[4]_pad ,
		\h1rdt2_dma[4]_pad ,
		_w2395_,
		_w2410_,
		_w6976_
	);
	LUT4 #(
		.INIT('h153f)
	) name4748 (
		\h1rdt4_br[4]_pad ,
		\h1rdt6_br[4]_pad ,
		_w2392_,
		_w2405_,
		_w6977_
	);
	LUT4 #(
		.INIT('h153f)
	) name4749 (
		\h1rdt4_dma[4]_pad ,
		\h1rdt7_br[4]_pad ,
		_w2391_,
		_w2411_,
		_w6978_
	);
	LUT4 #(
		.INIT('h153f)
	) name4750 (
		\h1rdt0_dma[4]_pad ,
		\h1rdt7_dma[4]_pad ,
		_w2404_,
		_w2414_,
		_w6979_
	);
	LUT4 #(
		.INIT('h8000)
	) name4751 (
		_w6976_,
		_w6977_,
		_w6978_,
		_w6979_,
		_w6980_
	);
	LUT3 #(
		.INIT('h2a)
	) name4752 (
		_w6703_,
		_w6975_,
		_w6980_,
		_w6981_
	);
	LUT3 #(
		.INIT('hfe)
	) name4753 (
		_w6959_,
		_w6970_,
		_w6981_,
		_w6982_
	);
	LUT3 #(
		.INIT('h70)
	) name4754 (
		_w6695_,
		_w6700_,
		_w6717_,
		_w6983_
	);
	LUT3 #(
		.INIT('h2a)
	) name4755 (
		_w6705_,
		_w6711_,
		_w6716_,
		_w6984_
	);
	LUT4 #(
		.INIT('h135f)
	) name4756 (
		\h1rdt2_br[5]_pad ,
		\h1rdt6_dma[5]_pad ,
		_w2389_,
		_w2413_,
		_w6985_
	);
	LUT4 #(
		.INIT('h153f)
	) name4757 (
		\h1rdt5_br[5]_pad ,
		\h1rdt5_dma[5]_pad ,
		_w2401_,
		_w2408_,
		_w6986_
	);
	LUT4 #(
		.INIT('h153f)
	) name4758 (
		\h1rdt0_br[5]_pad ,
		\h1rdt3_br[5]_pad ,
		_w2398_,
		_w2407_,
		_w6987_
	);
	LUT4 #(
		.INIT('h153f)
	) name4759 (
		\h1rdt1_br[5]_pad ,
		\h1rdt3_dma[5]_pad ,
		_w2394_,
		_w2400_,
		_w6988_
	);
	LUT4 #(
		.INIT('h8000)
	) name4760 (
		_w6985_,
		_w6986_,
		_w6987_,
		_w6988_,
		_w6989_
	);
	LUT4 #(
		.INIT('h135f)
	) name4761 (
		\h1rdt1_dma[5]_pad ,
		\h1rdt2_dma[5]_pad ,
		_w2395_,
		_w2410_,
		_w6990_
	);
	LUT4 #(
		.INIT('h153f)
	) name4762 (
		\h1rdt4_br[5]_pad ,
		\h1rdt6_br[5]_pad ,
		_w2392_,
		_w2405_,
		_w6991_
	);
	LUT4 #(
		.INIT('h153f)
	) name4763 (
		\h1rdt4_dma[5]_pad ,
		\h1rdt7_br[5]_pad ,
		_w2391_,
		_w2411_,
		_w6992_
	);
	LUT4 #(
		.INIT('h153f)
	) name4764 (
		\h1rdt0_dma[5]_pad ,
		\h1rdt7_dma[5]_pad ,
		_w2404_,
		_w2414_,
		_w6993_
	);
	LUT4 #(
		.INIT('h8000)
	) name4765 (
		_w6990_,
		_w6991_,
		_w6992_,
		_w6993_,
		_w6994_
	);
	LUT3 #(
		.INIT('h2a)
	) name4766 (
		_w6703_,
		_w6989_,
		_w6994_,
		_w6995_
	);
	LUT3 #(
		.INIT('hfe)
	) name4767 (
		_w6983_,
		_w6984_,
		_w6995_,
		_w6996_
	);
	LUT3 #(
		.INIT('h2a)
	) name4768 (
		_w6717_,
		_w6735_,
		_w6740_,
		_w6997_
	);
	LUT3 #(
		.INIT('h2a)
	) name4769 (
		_w6705_,
		_w6746_,
		_w6751_,
		_w6998_
	);
	LUT4 #(
		.INIT('h135f)
	) name4770 (
		\h1rdt6_br[6]_pad ,
		\h1rdt6_dma[6]_pad ,
		_w2392_,
		_w2413_,
		_w6999_
	);
	LUT4 #(
		.INIT('h153f)
	) name4771 (
		\h1rdt0_br[6]_pad ,
		\h1rdt1_br[6]_pad ,
		_w2400_,
		_w2407_,
		_w7000_
	);
	LUT4 #(
		.INIT('h153f)
	) name4772 (
		\h1rdt5_br[6]_pad ,
		\h1rdt7_br[6]_pad ,
		_w2391_,
		_w2408_,
		_w7001_
	);
	LUT4 #(
		.INIT('h153f)
	) name4773 (
		\h1rdt0_dma[6]_pad ,
		\h1rdt2_br[6]_pad ,
		_w2389_,
		_w2414_,
		_w7002_
	);
	LUT4 #(
		.INIT('h8000)
	) name4774 (
		_w6999_,
		_w7000_,
		_w7001_,
		_w7002_,
		_w7003_
	);
	LUT4 #(
		.INIT('h135f)
	) name4775 (
		\h1rdt4_br[6]_pad ,
		\h1rdt4_dma[6]_pad ,
		_w2405_,
		_w2411_,
		_w7004_
	);
	LUT4 #(
		.INIT('h135f)
	) name4776 (
		\h1rdt1_dma[6]_pad ,
		\h1rdt2_dma[6]_pad ,
		_w2395_,
		_w2410_,
		_w7005_
	);
	LUT4 #(
		.INIT('h135f)
	) name4777 (
		\h1rdt3_br[6]_pad ,
		\h1rdt5_dma[6]_pad ,
		_w2398_,
		_w2401_,
		_w7006_
	);
	LUT4 #(
		.INIT('h135f)
	) name4778 (
		\h1rdt3_dma[6]_pad ,
		\h1rdt7_dma[6]_pad ,
		_w2394_,
		_w2404_,
		_w7007_
	);
	LUT4 #(
		.INIT('h8000)
	) name4779 (
		_w7004_,
		_w7005_,
		_w7006_,
		_w7007_,
		_w7008_
	);
	LUT3 #(
		.INIT('h2a)
	) name4780 (
		_w6703_,
		_w7003_,
		_w7008_,
		_w7009_
	);
	LUT3 #(
		.INIT('hfe)
	) name4781 (
		_w6997_,
		_w6998_,
		_w7009_,
		_w7010_
	);
	LUT3 #(
		.INIT('h2a)
	) name4782 (
		_w6717_,
		_w6769_,
		_w6774_,
		_w7011_
	);
	LUT3 #(
		.INIT('h2a)
	) name4783 (
		_w6705_,
		_w6780_,
		_w6785_,
		_w7012_
	);
	LUT4 #(
		.INIT('h153f)
	) name4784 (
		\h1rdt1_dma[7]_pad ,
		\h1rdt3_dma[7]_pad ,
		_w2394_,
		_w2395_,
		_w7013_
	);
	LUT4 #(
		.INIT('h135f)
	) name4785 (
		\h1rdt0_br[7]_pad ,
		\h1rdt0_dma[7]_pad ,
		_w2407_,
		_w2414_,
		_w7014_
	);
	LUT4 #(
		.INIT('h135f)
	) name4786 (
		\h1rdt2_br[7]_pad ,
		\h1rdt7_br[7]_pad ,
		_w2389_,
		_w2391_,
		_w7015_
	);
	LUT4 #(
		.INIT('h153f)
	) name4787 (
		\h1rdt4_dma[7]_pad ,
		\h1rdt5_dma[7]_pad ,
		_w2401_,
		_w2411_,
		_w7016_
	);
	LUT4 #(
		.INIT('h8000)
	) name4788 (
		_w7013_,
		_w7014_,
		_w7015_,
		_w7016_,
		_w7017_
	);
	LUT4 #(
		.INIT('h153f)
	) name4789 (
		\h1rdt5_br[7]_pad ,
		\h1rdt6_br[7]_pad ,
		_w2392_,
		_w2408_,
		_w7018_
	);
	LUT4 #(
		.INIT('h135f)
	) name4790 (
		\h1rdt1_br[7]_pad ,
		\h1rdt4_br[7]_pad ,
		_w2400_,
		_w2405_,
		_w7019_
	);
	LUT4 #(
		.INIT('h135f)
	) name4791 (
		\h1rdt3_br[7]_pad ,
		\h1rdt6_dma[7]_pad ,
		_w2398_,
		_w2413_,
		_w7020_
	);
	LUT4 #(
		.INIT('h153f)
	) name4792 (
		\h1rdt2_dma[7]_pad ,
		\h1rdt7_dma[7]_pad ,
		_w2404_,
		_w2410_,
		_w7021_
	);
	LUT4 #(
		.INIT('h8000)
	) name4793 (
		_w7018_,
		_w7019_,
		_w7020_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h2a)
	) name4794 (
		_w6703_,
		_w7017_,
		_w7022_,
		_w7023_
	);
	LUT3 #(
		.INIT('hfe)
	) name4795 (
		_w7011_,
		_w7012_,
		_w7023_,
		_w7024_
	);
	LUT4 #(
		.INIT('h153f)
	) name4796 (
		\h1rdt0_br[24]_pad ,
		\h1rdt4_br[24]_pad ,
		_w2405_,
		_w2407_,
		_w7025_
	);
	LUT4 #(
		.INIT('h135f)
	) name4797 (
		\h1rdt2_br[24]_pad ,
		\h1rdt5_br[24]_pad ,
		_w2389_,
		_w2408_,
		_w7026_
	);
	LUT4 #(
		.INIT('h153f)
	) name4798 (
		\h1rdt6_dma[24]_pad ,
		\h1rdt7_br[24]_pad ,
		_w2391_,
		_w2413_,
		_w7027_
	);
	LUT4 #(
		.INIT('h153f)
	) name4799 (
		\h1rdt0_dma[24]_pad ,
		\h1rdt1_br[24]_pad ,
		_w2400_,
		_w2414_,
		_w7028_
	);
	LUT4 #(
		.INIT('h8000)
	) name4800 (
		_w7025_,
		_w7026_,
		_w7027_,
		_w7028_,
		_w7029_
	);
	LUT4 #(
		.INIT('h153f)
	) name4801 (
		\h1rdt4_dma[24]_pad ,
		\h1rdt7_dma[24]_pad ,
		_w2404_,
		_w2411_,
		_w7030_
	);
	LUT4 #(
		.INIT('h135f)
	) name4802 (
		\h1rdt3_dma[24]_pad ,
		\h1rdt5_dma[24]_pad ,
		_w2394_,
		_w2401_,
		_w7031_
	);
	LUT4 #(
		.INIT('h153f)
	) name4803 (
		\h1rdt2_dma[24]_pad ,
		\h1rdt3_br[24]_pad ,
		_w2398_,
		_w2410_,
		_w7032_
	);
	LUT4 #(
		.INIT('h153f)
	) name4804 (
		\h1rdt1_dma[24]_pad ,
		\h1rdt6_br[24]_pad ,
		_w2392_,
		_w2395_,
		_w7033_
	);
	LUT4 #(
		.INIT('h8000)
	) name4805 (
		_w7030_,
		_w7031_,
		_w7032_,
		_w7033_,
		_w7034_
	);
	LUT3 #(
		.INIT('h2a)
	) name4806 (
		_w6705_,
		_w7029_,
		_w7034_,
		_w7035_
	);
	LUT3 #(
		.INIT('h2a)
	) name4807 (
		_w6717_,
		_w6825_,
		_w6830_,
		_w7036_
	);
	LUT3 #(
		.INIT('h2a)
	) name4808 (
		_w6703_,
		_w6814_,
		_w6819_,
		_w7037_
	);
	LUT3 #(
		.INIT('hfe)
	) name4809 (
		_w7035_,
		_w7036_,
		_w7037_,
		_w7038_
	);
	LUT3 #(
		.INIT('h2a)
	) name4810 (
		_w6705_,
		_w6939_,
		_w6944_,
		_w7039_
	);
	LUT3 #(
		.INIT('h2a)
	) name4811 (
		_w6717_,
		_w6859_,
		_w6864_,
		_w7040_
	);
	LUT3 #(
		.INIT('h2a)
	) name4812 (
		_w6703_,
		_w6848_,
		_w6853_,
		_w7041_
	);
	LUT3 #(
		.INIT('hfe)
	) name4813 (
		_w7039_,
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h135f)
	) name4814 (
		\h1rdt0_br[26]_pad ,
		\h1rdt4_dma[26]_pad ,
		_w2407_,
		_w2411_,
		_w7043_
	);
	LUT4 #(
		.INIT('h153f)
	) name4815 (
		\h1rdt2_dma[26]_pad ,
		\h1rdt6_br[26]_pad ,
		_w2392_,
		_w2410_,
		_w7044_
	);
	LUT4 #(
		.INIT('h153f)
	) name4816 (
		\h1rdt1_br[26]_pad ,
		\h1rdt3_br[26]_pad ,
		_w2398_,
		_w2400_,
		_w7045_
	);
	LUT4 #(
		.INIT('h153f)
	) name4817 (
		\h1rdt0_dma[26]_pad ,
		\h1rdt5_br[26]_pad ,
		_w2408_,
		_w2414_,
		_w7046_
	);
	LUT4 #(
		.INIT('h8000)
	) name4818 (
		_w7043_,
		_w7044_,
		_w7045_,
		_w7046_,
		_w7047_
	);
	LUT4 #(
		.INIT('h135f)
	) name4819 (
		\h1rdt1_dma[26]_pad ,
		\h1rdt5_dma[26]_pad ,
		_w2395_,
		_w2401_,
		_w7048_
	);
	LUT4 #(
		.INIT('h135f)
	) name4820 (
		\h1rdt2_br[26]_pad ,
		\h1rdt3_dma[26]_pad ,
		_w2389_,
		_w2394_,
		_w7049_
	);
	LUT4 #(
		.INIT('h135f)
	) name4821 (
		\h1rdt7_br[26]_pad ,
		\h1rdt7_dma[26]_pad ,
		_w2391_,
		_w2404_,
		_w7050_
	);
	LUT4 #(
		.INIT('h135f)
	) name4822 (
		\h1rdt4_br[26]_pad ,
		\h1rdt6_dma[26]_pad ,
		_w2405_,
		_w2413_,
		_w7051_
	);
	LUT4 #(
		.INIT('h8000)
	) name4823 (
		_w7048_,
		_w7049_,
		_w7050_,
		_w7051_,
		_w7052_
	);
	LUT3 #(
		.INIT('h2a)
	) name4824 (
		_w6705_,
		_w7047_,
		_w7052_,
		_w7053_
	);
	LUT3 #(
		.INIT('h2a)
	) name4825 (
		_w6717_,
		_w6893_,
		_w6898_,
		_w7054_
	);
	LUT3 #(
		.INIT('h2a)
	) name4826 (
		_w6703_,
		_w6882_,
		_w6887_,
		_w7055_
	);
	LUT3 #(
		.INIT('hfe)
	) name4827 (
		_w7053_,
		_w7054_,
		_w7055_,
		_w7056_
	);
	LUT4 #(
		.INIT('h135f)
	) name4828 (
		\h1rdt2_br[27]_pad ,
		\h1rdt6_dma[27]_pad ,
		_w2389_,
		_w2413_,
		_w7057_
	);
	LUT4 #(
		.INIT('h153f)
	) name4829 (
		\h1rdt1_dma[27]_pad ,
		\h1rdt3_dma[27]_pad ,
		_w2394_,
		_w2395_,
		_w7058_
	);
	LUT4 #(
		.INIT('h153f)
	) name4830 (
		\h1rdt0_br[27]_pad ,
		\h1rdt7_br[27]_pad ,
		_w2391_,
		_w2407_,
		_w7059_
	);
	LUT4 #(
		.INIT('h153f)
	) name4831 (
		\h1rdt2_dma[27]_pad ,
		\h1rdt5_dma[27]_pad ,
		_w2401_,
		_w2410_,
		_w7060_
	);
	LUT4 #(
		.INIT('h8000)
	) name4832 (
		_w7057_,
		_w7058_,
		_w7059_,
		_w7060_,
		_w7061_
	);
	LUT4 #(
		.INIT('h153f)
	) name4833 (
		\h1rdt4_br[27]_pad ,
		\h1rdt6_br[27]_pad ,
		_w2392_,
		_w2405_,
		_w7062_
	);
	LUT4 #(
		.INIT('h153f)
	) name4834 (
		\h1rdt0_dma[27]_pad ,
		\h1rdt5_br[27]_pad ,
		_w2408_,
		_w2414_,
		_w7063_
	);
	LUT4 #(
		.INIT('h153f)
	) name4835 (
		\h1rdt1_br[27]_pad ,
		\h1rdt3_br[27]_pad ,
		_w2398_,
		_w2400_,
		_w7064_
	);
	LUT4 #(
		.INIT('h153f)
	) name4836 (
		\h1rdt4_dma[27]_pad ,
		\h1rdt7_dma[27]_pad ,
		_w2404_,
		_w2411_,
		_w7065_
	);
	LUT4 #(
		.INIT('h8000)
	) name4837 (
		_w7062_,
		_w7063_,
		_w7064_,
		_w7065_,
		_w7066_
	);
	LUT3 #(
		.INIT('h2a)
	) name4838 (
		_w6705_,
		_w7061_,
		_w7066_,
		_w7067_
	);
	LUT3 #(
		.INIT('h2a)
	) name4839 (
		_w6717_,
		_w6927_,
		_w6932_,
		_w7068_
	);
	LUT3 #(
		.INIT('h2a)
	) name4840 (
		_w6703_,
		_w6916_,
		_w6921_,
		_w7069_
	);
	LUT3 #(
		.INIT('hfe)
	) name4841 (
		_w7067_,
		_w7068_,
		_w7069_,
		_w7070_
	);
	LUT4 #(
		.INIT('h135f)
	) name4842 (
		\h1rdt2_br[28]_pad ,
		\h1rdt6_dma[28]_pad ,
		_w2389_,
		_w2413_,
		_w7071_
	);
	LUT4 #(
		.INIT('h135f)
	) name4843 (
		\h1rdt3_dma[28]_pad ,
		\h1rdt5_br[28]_pad ,
		_w2394_,
		_w2408_,
		_w7072_
	);
	LUT4 #(
		.INIT('h153f)
	) name4844 (
		\h1rdt0_br[28]_pad ,
		\h1rdt3_br[28]_pad ,
		_w2398_,
		_w2407_,
		_w7073_
	);
	LUT4 #(
		.INIT('h135f)
	) name4845 (
		\h1rdt1_br[28]_pad ,
		\h1rdt5_dma[28]_pad ,
		_w2400_,
		_w2401_,
		_w7074_
	);
	LUT4 #(
		.INIT('h8000)
	) name4846 (
		_w7071_,
		_w7072_,
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('h135f)
	) name4847 (
		\h1rdt1_dma[28]_pad ,
		\h1rdt2_dma[28]_pad ,
		_w2395_,
		_w2410_,
		_w7076_
	);
	LUT4 #(
		.INIT('h153f)
	) name4848 (
		\h1rdt4_br[28]_pad ,
		\h1rdt6_br[28]_pad ,
		_w2392_,
		_w2405_,
		_w7077_
	);
	LUT4 #(
		.INIT('h153f)
	) name4849 (
		\h1rdt4_dma[28]_pad ,
		\h1rdt7_br[28]_pad ,
		_w2391_,
		_w2411_,
		_w7078_
	);
	LUT4 #(
		.INIT('h153f)
	) name4850 (
		\h1rdt0_dma[28]_pad ,
		\h1rdt7_dma[28]_pad ,
		_w2404_,
		_w2414_,
		_w7079_
	);
	LUT4 #(
		.INIT('h8000)
	) name4851 (
		_w7076_,
		_w7077_,
		_w7078_,
		_w7079_,
		_w7080_
	);
	LUT3 #(
		.INIT('h2a)
	) name4852 (
		_w6705_,
		_w7075_,
		_w7080_,
		_w7081_
	);
	LUT3 #(
		.INIT('h2a)
	) name4853 (
		_w6717_,
		_w6975_,
		_w6980_,
		_w7082_
	);
	LUT3 #(
		.INIT('h2a)
	) name4854 (
		_w6703_,
		_w6964_,
		_w6969_,
		_w7083_
	);
	LUT3 #(
		.INIT('hfe)
	) name4855 (
		_w7081_,
		_w7082_,
		_w7083_,
		_w7084_
	);
	LUT3 #(
		.INIT('h2a)
	) name4856 (
		_w6717_,
		_w6989_,
		_w6994_,
		_w7085_
	);
	LUT3 #(
		.INIT('h2a)
	) name4857 (
		_w6705_,
		_w6723_,
		_w6728_,
		_w7086_
	);
	LUT3 #(
		.INIT('h70)
	) name4858 (
		_w6695_,
		_w6700_,
		_w6703_,
		_w7087_
	);
	LUT3 #(
		.INIT('hfe)
	) name4859 (
		_w7085_,
		_w7086_,
		_w7087_,
		_w7088_
	);
	LUT3 #(
		.INIT('h2a)
	) name4860 (
		_w6717_,
		_w7047_,
		_w7052_,
		_w7089_
	);
	LUT3 #(
		.INIT('h2a)
	) name4861 (
		_w6705_,
		_w6893_,
		_w6898_,
		_w7090_
	);
	LUT3 #(
		.INIT('h2a)
	) name4862 (
		_w6703_,
		_w6871_,
		_w6876_,
		_w7091_
	);
	LUT3 #(
		.INIT('hfe)
	) name4863 (
		_w7089_,
		_w7090_,
		_w7091_,
		_w7092_
	);
	LUT3 #(
		.INIT('h2a)
	) name4864 (
		_w6717_,
		_w7003_,
		_w7008_,
		_w7093_
	);
	LUT3 #(
		.INIT('h2a)
	) name4865 (
		_w6705_,
		_w6757_,
		_w6762_,
		_w7094_
	);
	LUT3 #(
		.INIT('h2a)
	) name4866 (
		_w6703_,
		_w6735_,
		_w6740_,
		_w7095_
	);
	LUT3 #(
		.INIT('hfe)
	) name4867 (
		_w7093_,
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT3 #(
		.INIT('h2a)
	) name4868 (
		_w6717_,
		_w7017_,
		_w7022_,
		_w7097_
	);
	LUT3 #(
		.INIT('h2a)
	) name4869 (
		_w6705_,
		_w6791_,
		_w6796_,
		_w7098_
	);
	LUT3 #(
		.INIT('h2a)
	) name4870 (
		_w6703_,
		_w6769_,
		_w6774_,
		_w7099_
	);
	LUT3 #(
		.INIT('hfe)
	) name4871 (
		_w7097_,
		_w7098_,
		_w7099_,
		_w7100_
	);
	LUT3 #(
		.INIT('h2a)
	) name4872 (
		_w6717_,
		_w7061_,
		_w7066_,
		_w7101_
	);
	LUT3 #(
		.INIT('h2a)
	) name4873 (
		_w6705_,
		_w6927_,
		_w6932_,
		_w7102_
	);
	LUT3 #(
		.INIT('h2a)
	) name4874 (
		_w6703_,
		_w6905_,
		_w6910_,
		_w7103_
	);
	LUT3 #(
		.INIT('hfe)
	) name4875 (
		_w7101_,
		_w7102_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('h2a)
	) name4876 (
		_w6717_,
		_w7075_,
		_w7080_,
		_w7105_
	);
	LUT3 #(
		.INIT('h2a)
	) name4877 (
		_w6705_,
		_w6975_,
		_w6980_,
		_w7106_
	);
	LUT3 #(
		.INIT('h2a)
	) name4878 (
		_w6703_,
		_w6953_,
		_w6958_,
		_w7107_
	);
	LUT3 #(
		.INIT('hfe)
	) name4879 (
		_w7105_,
		_w7106_,
		_w7107_,
		_w7108_
	);
	LUT3 #(
		.INIT('h2a)
	) name4880 (
		_w6705_,
		_w6989_,
		_w6994_,
		_w7109_
	);
	LUT3 #(
		.INIT('h2a)
	) name4881 (
		_w6717_,
		_w6723_,
		_w6728_,
		_w7110_
	);
	LUT3 #(
		.INIT('h2a)
	) name4882 (
		_w6703_,
		_w6711_,
		_w6716_,
		_w7111_
	);
	LUT3 #(
		.INIT('hfe)
	) name4883 (
		_w7109_,
		_w7110_,
		_w7111_,
		_w7112_
	);
	LUT3 #(
		.INIT('h2a)
	) name4884 (
		_w6705_,
		_w7003_,
		_w7008_,
		_w7113_
	);
	LUT3 #(
		.INIT('h2a)
	) name4885 (
		_w6717_,
		_w6757_,
		_w6762_,
		_w7114_
	);
	LUT3 #(
		.INIT('h2a)
	) name4886 (
		_w6703_,
		_w6746_,
		_w6751_,
		_w7115_
	);
	LUT3 #(
		.INIT('hfe)
	) name4887 (
		_w7113_,
		_w7114_,
		_w7115_,
		_w7116_
	);
	LUT3 #(
		.INIT('h2a)
	) name4888 (
		_w6705_,
		_w7017_,
		_w7022_,
		_w7117_
	);
	LUT3 #(
		.INIT('h2a)
	) name4889 (
		_w6717_,
		_w6791_,
		_w6796_,
		_w7118_
	);
	LUT3 #(
		.INIT('h2a)
	) name4890 (
		_w6703_,
		_w6780_,
		_w6785_,
		_w7119_
	);
	LUT3 #(
		.INIT('hfe)
	) name4891 (
		_w7117_,
		_w7118_,
		_w7119_,
		_w7120_
	);
	LUT3 #(
		.INIT('h2a)
	) name4892 (
		_w6717_,
		_w6803_,
		_w6808_,
		_w7121_
	);
	LUT3 #(
		.INIT('h2a)
	) name4893 (
		_w6705_,
		_w6814_,
		_w6819_,
		_w7122_
	);
	LUT3 #(
		.INIT('h2a)
	) name4894 (
		_w6703_,
		_w7029_,
		_w7034_,
		_w7123_
	);
	LUT3 #(
		.INIT('hfe)
	) name4895 (
		_w7121_,
		_w7122_,
		_w7123_,
		_w7124_
	);
	LUT3 #(
		.INIT('h2a)
	) name4896 (
		_w6717_,
		_w6837_,
		_w6842_,
		_w7125_
	);
	LUT3 #(
		.INIT('h2a)
	) name4897 (
		_w6705_,
		_w6848_,
		_w6853_,
		_w7126_
	);
	LUT3 #(
		.INIT('h2a)
	) name4898 (
		_w6703_,
		_w6939_,
		_w6944_,
		_w7127_
	);
	LUT3 #(
		.INIT('hfe)
	) name4899 (
		_w7125_,
		_w7126_,
		_w7127_,
		_w7128_
	);
	LUT3 #(
		.INIT('h2a)
	) name4900 (
		_w6717_,
		_w7029_,
		_w7034_,
		_w7129_
	);
	LUT3 #(
		.INIT('h2a)
	) name4901 (
		_w6705_,
		_w6825_,
		_w6830_,
		_w7130_
	);
	LUT3 #(
		.INIT('h2a)
	) name4902 (
		_w6703_,
		_w6803_,
		_w6808_,
		_w7131_
	);
	LUT3 #(
		.INIT('hfe)
	) name4903 (
		_w7129_,
		_w7130_,
		_w7131_,
		_w7132_
	);
	LUT3 #(
		.INIT('h2a)
	) name4904 (
		_w6717_,
		_w6871_,
		_w6876_,
		_w7133_
	);
	LUT3 #(
		.INIT('h2a)
	) name4905 (
		_w6705_,
		_w6882_,
		_w6887_,
		_w7134_
	);
	LUT3 #(
		.INIT('h2a)
	) name4906 (
		_w6703_,
		_w7047_,
		_w7052_,
		_w7135_
	);
	LUT3 #(
		.INIT('hfe)
	) name4907 (
		_w7133_,
		_w7134_,
		_w7135_,
		_w7136_
	);
	LUT3 #(
		.INIT('h2a)
	) name4908 (
		_w6717_,
		_w6905_,
		_w6910_,
		_w7137_
	);
	LUT3 #(
		.INIT('h2a)
	) name4909 (
		_w6705_,
		_w6916_,
		_w6921_,
		_w7138_
	);
	LUT3 #(
		.INIT('h2a)
	) name4910 (
		_w6703_,
		_w7061_,
		_w7066_,
		_w7139_
	);
	LUT3 #(
		.INIT('hfe)
	) name4911 (
		_w7137_,
		_w7138_,
		_w7139_,
		_w7140_
	);
	LUT3 #(
		.INIT('h2a)
	) name4912 (
		_w6717_,
		_w6953_,
		_w6958_,
		_w7141_
	);
	LUT3 #(
		.INIT('h2a)
	) name4913 (
		_w6705_,
		_w6964_,
		_w6969_,
		_w7142_
	);
	LUT3 #(
		.INIT('h2a)
	) name4914 (
		_w6703_,
		_w7075_,
		_w7080_,
		_w7143_
	);
	LUT3 #(
		.INIT('hfe)
	) name4915 (
		_w7141_,
		_w7142_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('hca00)
	) name4916 (
		\ch_sel_dma_reqd1_reg[4]/NET0131 ,
		\ch_sel_dma_reqd2_reg[4]/NET0131 ,
		\ctl_rf_sync_reg[4]/NET0131 ,
		\dma_ack[4]_pad ,
		_w7145_
	);
	LUT2 #(
		.INIT('h4)
	) name4917 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_c4_rf_mode_reg/NET0131 ,
		_w7146_
	);
	LUT4 #(
		.INIT('h0040)
	) name4918 (
		\ctl_rf_c4_rf_chabt_reg/NET0131 ,
		\ctl_rf_c4_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[4]_pad ,
		_w7147_
	);
	LUT3 #(
		.INIT('h80)
	) name4919 (
		_w2507_,
		_w2508_,
		_w7147_,
		_w7148_
	);
	LUT3 #(
		.INIT('hec)
	) name4920 (
		_w2520_,
		_w7145_,
		_w7148_,
		_w7149_
	);
	LUT4 #(
		.INIT('hca00)
	) name4921 (
		\ch_sel_dma_reqd1_reg[1]/NET0131 ,
		\ch_sel_dma_reqd2_reg[1]/P0001 ,
		\ctl_rf_sync_reg[1]/NET0131 ,
		\dma_ack[1]_pad ,
		_w7150_
	);
	LUT2 #(
		.INIT('h4)
	) name4922 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_c1_rf_mode_reg/NET0131 ,
		_w7151_
	);
	LUT4 #(
		.INIT('h0040)
	) name4923 (
		\ctl_rf_c1_rf_chabt_reg/NET0131 ,
		\ctl_rf_c1_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[1]_pad ,
		_w7152_
	);
	LUT3 #(
		.INIT('h70)
	) name4924 (
		_w2507_,
		_w2508_,
		_w7152_,
		_w7153_
	);
	LUT3 #(
		.INIT('hec)
	) name4925 (
		_w2549_,
		_w7150_,
		_w7153_,
		_w7154_
	);
	LUT4 #(
		.INIT('h4155)
	) name4926 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w7155_
	);
	LUT3 #(
		.INIT('h15)
	) name4927 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		_w2426_,
		_w2427_,
		_w7156_
	);
	LUT4 #(
		.INIT('h0405)
	) name4928 (
		\de_de_st_reg[5]/NET0131 ,
		_w2424_,
		_w7155_,
		_w7156_,
		_w7157_
	);
	LUT4 #(
		.INIT('hca00)
	) name4929 (
		\ch_sel_dma_reqd1_reg[7]/NET0131 ,
		\ch_sel_dma_reqd2_reg[7]/NET0131 ,
		\ctl_rf_sync_reg[7]/NET0131 ,
		\dma_ack[7]_pad ,
		_w7158_
	);
	LUT2 #(
		.INIT('h4)
	) name4930 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\ctl_rf_c7_rf_mode_reg/NET0131 ,
		_w7159_
	);
	LUT4 #(
		.INIT('h0040)
	) name4931 (
		\ctl_rf_c7_rf_chabt_reg/NET0131 ,
		\ctl_rf_c7_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[7]_pad ,
		_w7160_
	);
	LUT3 #(
		.INIT('h70)
	) name4932 (
		_w2507_,
		_w2508_,
		_w7160_,
		_w7161_
	);
	LUT3 #(
		.INIT('hec)
	) name4933 (
		_w2527_,
		_w7158_,
		_w7161_,
		_w7162_
	);
	LUT4 #(
		.INIT('hca00)
	) name4934 (
		\ch_sel_dma_reqd1_reg[2]/NET0131 ,
		\ch_sel_dma_reqd2_reg[2]/P0001 ,
		\ctl_rf_sync_reg[2]/NET0131 ,
		\dma_ack[2]_pad ,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name4935 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_c2_rf_mode_reg/NET0131 ,
		_w7164_
	);
	LUT4 #(
		.INIT('h0040)
	) name4936 (
		\ctl_rf_c2_rf_chabt_reg/NET0131 ,
		\ctl_rf_c2_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[2]_pad ,
		_w7165_
	);
	LUT3 #(
		.INIT('h80)
	) name4937 (
		_w2507_,
		_w2508_,
		_w7165_,
		_w7166_
	);
	LUT3 #(
		.INIT('hec)
	) name4938 (
		_w2534_,
		_w7163_,
		_w7166_,
		_w7167_
	);
	LUT4 #(
		.INIT('hca00)
	) name4939 (
		\ch_sel_dma_reqd1_reg[3]/NET0131 ,
		\ch_sel_dma_reqd2_reg[3]/P0001 ,
		\ctl_rf_sync_reg[3]/NET0131 ,
		\dma_ack[3]_pad ,
		_w7168_
	);
	LUT2 #(
		.INIT('h4)
	) name4940 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\ctl_rf_c3_rf_mode_reg/NET0131 ,
		_w7169_
	);
	LUT4 #(
		.INIT('h0040)
	) name4941 (
		\ctl_rf_c3_rf_chabt_reg/NET0131 ,
		\ctl_rf_c3_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[3]_pad ,
		_w7170_
	);
	LUT3 #(
		.INIT('h70)
	) name4942 (
		_w2507_,
		_w2508_,
		_w7170_,
		_w7171_
	);
	LUT3 #(
		.INIT('hec)
	) name4943 (
		_w2534_,
		_w7168_,
		_w7171_,
		_w7172_
	);
	LUT4 #(
		.INIT('hca00)
	) name4944 (
		\ch_sel_dma_reqd1_reg[5]/NET0131 ,
		\ch_sel_dma_reqd2_reg[5]/NET0131 ,
		\ctl_rf_sync_reg[5]/NET0131 ,
		\dma_ack[5]_pad ,
		_w7173_
	);
	LUT2 #(
		.INIT('h4)
	) name4945 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_c5_rf_mode_reg/NET0131 ,
		_w7174_
	);
	LUT4 #(
		.INIT('h0040)
	) name4946 (
		\ctl_rf_c5_rf_chabt_reg/NET0131 ,
		\ctl_rf_c5_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[5]_pad ,
		_w7175_
	);
	LUT3 #(
		.INIT('h70)
	) name4947 (
		_w2507_,
		_w2508_,
		_w7175_,
		_w7176_
	);
	LUT3 #(
		.INIT('hec)
	) name4948 (
		_w2520_,
		_w7173_,
		_w7176_,
		_w7177_
	);
	LUT4 #(
		.INIT('hca00)
	) name4949 (
		\ch_sel_dma_reqd1_reg[6]/NET0131 ,
		\ch_sel_dma_reqd2_reg[6]/NET0131 ,
		\ctl_rf_sync_reg[6]/NET0131 ,
		\dma_ack[6]_pad ,
		_w7178_
	);
	LUT2 #(
		.INIT('h4)
	) name4950 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_c6_rf_mode_reg/NET0131 ,
		_w7179_
	);
	LUT4 #(
		.INIT('h0040)
	) name4951 (
		\ctl_rf_c6_rf_chabt_reg/NET0131 ,
		\ctl_rf_c6_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[6]_pad ,
		_w7180_
	);
	LUT3 #(
		.INIT('h80)
	) name4952 (
		_w2507_,
		_w2508_,
		_w7180_,
		_w7181_
	);
	LUT3 #(
		.INIT('hec)
	) name4953 (
		_w2527_,
		_w7178_,
		_w7181_,
		_w7182_
	);
	LUT4 #(
		.INIT('hca00)
	) name4954 (
		\ch_sel_dma_reqd1_reg[0]/NET0131 ,
		\ch_sel_dma_reqd2_reg[0]/NET0131 ,
		\ctl_rf_sync_reg[0]/NET0131 ,
		\dma_ack[0]_pad ,
		_w7183_
	);
	LUT2 #(
		.INIT('h4)
	) name4955 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_c0_rf_mode_reg/NET0131 ,
		_w7184_
	);
	LUT4 #(
		.INIT('h0040)
	) name4956 (
		\ctl_rf_c0_rf_chabt_reg/NET0131 ,
		\ctl_rf_c0_rf_mode_reg/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\dma_ack[0]_pad ,
		_w7185_
	);
	LUT3 #(
		.INIT('h80)
	) name4957 (
		_w2507_,
		_w2508_,
		_w7185_,
		_w7186_
	);
	LUT3 #(
		.INIT('hec)
	) name4958 (
		_w2549_,
		_w7183_,
		_w7186_,
		_w7187_
	);
	LUT4 #(
		.INIT('hca00)
	) name4959 (
		\ch_sel_dma_reqd1_reg[2]/NET0131 ,
		\ch_sel_dma_reqd2_reg[2]/P0001 ,
		\ctl_rf_sync_reg[2]/NET0131 ,
		\dma_tc[2]_pad ,
		_w7188_
	);
	LUT3 #(
		.INIT('h80)
	) name4960 (
		_w2507_,
		_w2508_,
		_w7164_,
		_w7189_
	);
	LUT2 #(
		.INIT('h2)
	) name4961 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[2]_pad ,
		_w7190_
	);
	LUT4 #(
		.INIT('h8000)
	) name4962 (
		_w2424_,
		_w2534_,
		_w7189_,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('he)
	) name4963 (
		_w7188_,
		_w7191_,
		_w7192_
	);
	LUT4 #(
		.INIT('hca00)
	) name4964 (
		\ch_sel_dma_reqd1_reg[7]/NET0131 ,
		\ch_sel_dma_reqd2_reg[7]/NET0131 ,
		\ctl_rf_sync_reg[7]/NET0131 ,
		\dma_tc[7]_pad ,
		_w7193_
	);
	LUT3 #(
		.INIT('h70)
	) name4965 (
		_w2507_,
		_w2508_,
		_w7159_,
		_w7194_
	);
	LUT2 #(
		.INIT('h2)
	) name4966 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[7]_pad ,
		_w7195_
	);
	LUT4 #(
		.INIT('h8000)
	) name4967 (
		_w2424_,
		_w2527_,
		_w7194_,
		_w7195_,
		_w7196_
	);
	LUT2 #(
		.INIT('he)
	) name4968 (
		_w7193_,
		_w7196_,
		_w7197_
	);
	LUT4 #(
		.INIT('hca00)
	) name4969 (
		\ch_sel_dma_reqd1_reg[3]/NET0131 ,
		\ch_sel_dma_reqd2_reg[3]/P0001 ,
		\ctl_rf_sync_reg[3]/NET0131 ,
		\dma_tc[3]_pad ,
		_w7198_
	);
	LUT3 #(
		.INIT('h70)
	) name4970 (
		_w2507_,
		_w2508_,
		_w7169_,
		_w7199_
	);
	LUT2 #(
		.INIT('h2)
	) name4971 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[3]_pad ,
		_w7200_
	);
	LUT4 #(
		.INIT('h8000)
	) name4972 (
		_w2424_,
		_w2534_,
		_w7199_,
		_w7200_,
		_w7201_
	);
	LUT2 #(
		.INIT('he)
	) name4973 (
		_w7198_,
		_w7201_,
		_w7202_
	);
	LUT4 #(
		.INIT('hca00)
	) name4974 (
		\ch_sel_dma_reqd1_reg[5]/NET0131 ,
		\ch_sel_dma_reqd2_reg[5]/NET0131 ,
		\ctl_rf_sync_reg[5]/NET0131 ,
		\dma_tc[5]_pad ,
		_w7203_
	);
	LUT3 #(
		.INIT('h70)
	) name4975 (
		_w2507_,
		_w2508_,
		_w7174_,
		_w7204_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[5]_pad ,
		_w7205_
	);
	LUT4 #(
		.INIT('h8000)
	) name4977 (
		_w2424_,
		_w2520_,
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('he)
	) name4978 (
		_w7203_,
		_w7206_,
		_w7207_
	);
	LUT4 #(
		.INIT('hca00)
	) name4979 (
		\ch_sel_dma_reqd1_reg[0]/NET0131 ,
		\ch_sel_dma_reqd2_reg[0]/NET0131 ,
		\ctl_rf_sync_reg[0]/NET0131 ,
		\dma_tc[0]_pad ,
		_w7208_
	);
	LUT3 #(
		.INIT('h80)
	) name4980 (
		_w2507_,
		_w2508_,
		_w7184_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name4981 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[0]_pad ,
		_w7210_
	);
	LUT4 #(
		.INIT('h8000)
	) name4982 (
		_w2424_,
		_w2549_,
		_w7209_,
		_w7210_,
		_w7211_
	);
	LUT2 #(
		.INIT('he)
	) name4983 (
		_w7208_,
		_w7211_,
		_w7212_
	);
	LUT4 #(
		.INIT('hca00)
	) name4984 (
		\ch_sel_dma_reqd1_reg[1]/NET0131 ,
		\ch_sel_dma_reqd2_reg[1]/P0001 ,
		\ctl_rf_sync_reg[1]/NET0131 ,
		\dma_tc[1]_pad ,
		_w7213_
	);
	LUT3 #(
		.INIT('h70)
	) name4985 (
		_w2507_,
		_w2508_,
		_w7151_,
		_w7214_
	);
	LUT2 #(
		.INIT('h2)
	) name4986 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[1]_pad ,
		_w7215_
	);
	LUT4 #(
		.INIT('h8000)
	) name4987 (
		_w2424_,
		_w2549_,
		_w7214_,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('he)
	) name4988 (
		_w7213_,
		_w7216_,
		_w7217_
	);
	LUT4 #(
		.INIT('hca00)
	) name4989 (
		\ch_sel_dma_reqd1_reg[4]/NET0131 ,
		\ch_sel_dma_reqd2_reg[4]/NET0131 ,
		\ctl_rf_sync_reg[4]/NET0131 ,
		\dma_tc[4]_pad ,
		_w7218_
	);
	LUT3 #(
		.INIT('h80)
	) name4990 (
		_w2507_,
		_w2508_,
		_w7146_,
		_w7219_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[4]_pad ,
		_w7220_
	);
	LUT4 #(
		.INIT('h8000)
	) name4992 (
		_w2424_,
		_w2520_,
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT2 #(
		.INIT('he)
	) name4993 (
		_w7218_,
		_w7221_,
		_w7222_
	);
	LUT4 #(
		.INIT('hca00)
	) name4994 (
		\ch_sel_dma_reqd1_reg[6]/NET0131 ,
		\ch_sel_dma_reqd2_reg[6]/NET0131 ,
		\ctl_rf_sync_reg[6]/NET0131 ,
		\dma_tc[6]_pad ,
		_w7223_
	);
	LUT3 #(
		.INIT('h80)
	) name4995 (
		_w2507_,
		_w2508_,
		_w7179_,
		_w7224_
	);
	LUT2 #(
		.INIT('h2)
	) name4996 (
		\de_de_st_reg[5]/NET0131 ,
		\dma_tc[6]_pad ,
		_w7225_
	);
	LUT4 #(
		.INIT('h8000)
	) name4997 (
		_w2424_,
		_w2527_,
		_w7224_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('he)
	) name4998 (
		_w7223_,
		_w7226_,
		_w7227_
	);
	LUT4 #(
		.INIT('h8000)
	) name4999 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2247_,
		_w2991_,
		_w7228_
	);
	LUT4 #(
		.INIT('h8000)
	) name5000 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2247_,
		_w3112_,
		_w7229_
	);
	LUT4 #(
		.INIT('h8000)
	) name5001 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2254_,
		_w3112_,
		_w7230_
	);
	LUT4 #(
		.INIT('h8000)
	) name5002 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2254_,
		_w2991_,
		_w7231_
	);
	LUT3 #(
		.INIT('h10)
	) name5003 (
		_w2993_,
		_w2994_,
		_w6141_,
		_w7232_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3135_,
		_w7233_
	);
	LUT4 #(
		.INIT('h8000)
	) name5005 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2239_,
		_w2991_,
		_w7234_
	);
	LUT4 #(
		.INIT('h8000)
	) name5006 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2229_,
		_w2239_,
		_w3112_,
		_w7235_
	);
	LUT2 #(
		.INIT('h2)
	) name5007 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3114_,
		_w7236_
	);
	LUT3 #(
		.INIT('h10)
	) name5008 (
		_w2993_,
		_w2994_,
		_w6133_,
		_w7237_
	);
	LUT2 #(
		.INIT('h2)
	) name5009 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3114_,
		_w7238_
	);
	LUT3 #(
		.INIT('h10)
	) name5010 (
		_w2993_,
		_w2994_,
		_w6137_,
		_w7239_
	);
	LUT3 #(
		.INIT('h10)
	) name5011 (
		_w2993_,
		_w2994_,
		_w6129_,
		_w7240_
	);
	LUT3 #(
		.INIT('h10)
	) name5012 (
		_w2993_,
		_w2994_,
		_w6149_,
		_w7241_
	);
	LUT4 #(
		.INIT('h8000)
	) name5013 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2244_,
		_w3112_,
		_w7242_
	);
	LUT4 #(
		.INIT('h8000)
	) name5014 (
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w2239_,
		_w2244_,
		_w2991_,
		_w7243_
	);
	LUT3 #(
		.INIT('h10)
	) name5015 (
		_w2993_,
		_w2994_,
		_w6157_,
		_w7244_
	);
	LUT2 #(
		.INIT('h2)
	) name5016 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3135_,
		_w7245_
	);
	LUT3 #(
		.INIT('h10)
	) name5017 (
		_w2993_,
		_w2994_,
		_w6145_,
		_w7246_
	);
	LUT3 #(
		.INIT('h10)
	) name5018 (
		_w2993_,
		_w2994_,
		_w6153_,
		_w7247_
	);
	LUT2 #(
		.INIT('h2)
	) name5019 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2995_,
		_w7248_
	);
	LUT2 #(
		.INIT('h2)
	) name5020 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2995_,
		_w7249_
	);
	LUT2 #(
		.INIT('h2)
	) name5021 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3125_,
		_w7250_
	);
	LUT2 #(
		.INIT('h2)
	) name5022 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3125_,
		_w7251_
	);
	LUT2 #(
		.INIT('h2)
	) name5023 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3155_,
		_w7252_
	);
	LUT2 #(
		.INIT('h2)
	) name5024 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3175_,
		_w7253_
	);
	LUT2 #(
		.INIT('h2)
	) name5025 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3145_,
		_w7254_
	);
	LUT2 #(
		.INIT('h2)
	) name5026 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3155_,
		_w7255_
	);
	LUT2 #(
		.INIT('h2)
	) name5027 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3165_,
		_w7256_
	);
	LUT2 #(
		.INIT('h2)
	) name5028 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3165_,
		_w7257_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5029 (
		\ctl_rf_c0_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_c6_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[0]/NET0131 ,
		\ctl_rf_tc_reg[6]/NET0131 ,
		_w7258_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5030 (
		\ctl_rf_c3_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_c7_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[3]/NET0131 ,
		\ctl_rf_tc_reg[7]/NET0131 ,
		_w7259_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5031 (
		\ctl_rf_c1_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_c2_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[1]/NET0131 ,
		\ctl_rf_tc_reg[2]/NET0131 ,
		_w7260_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5032 (
		\ctl_rf_c4_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_c5_rf_int_tc1_msk_reg/NET0131 ,
		\ctl_rf_tc_reg[4]/NET0131 ,
		\ctl_rf_tc_reg[5]/NET0131 ,
		_w7261_
	);
	LUT4 #(
		.INIT('h8000)
	) name5033 (
		_w7258_,
		_w7259_,
		_w7260_,
		_w7261_,
		_w7262_
	);
	LUT4 #(
		.INIT('h7fff)
	) name5034 (
		_w7258_,
		_w7259_,
		_w7260_,
		_w7261_,
		_w7263_
	);
	LUT4 #(
		.INIT('hf531)
	) name5035 (
		\ctl_rf_abt_reg[4]/NET0131 ,
		\ctl_rf_abt_reg[5]/NET0131 ,
		\ctl_rf_c4_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c5_rf_int_abt_msk_reg/NET0131 ,
		_w7264_
	);
	LUT4 #(
		.INIT('hf531)
	) name5036 (
		\ctl_rf_abt_reg[6]/NET0131 ,
		\ctl_rf_abt_reg[7]/NET0131 ,
		\ctl_rf_c6_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c7_rf_int_abt_msk_reg/NET0131 ,
		_w7265_
	);
	LUT4 #(
		.INIT('hf531)
	) name5037 (
		\ctl_rf_abt_reg[0]/NET0131 ,
		\ctl_rf_abt_reg[1]/NET0131 ,
		\ctl_rf_c0_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c1_rf_int_abt_msk_reg/NET0131 ,
		_w7266_
	);
	LUT4 #(
		.INIT('hf531)
	) name5038 (
		\ctl_rf_abt_reg[2]/NET0131 ,
		\ctl_rf_abt_reg[3]/NET0131 ,
		\ctl_rf_c2_rf_int_abt_msk_reg/NET0131 ,
		\ctl_rf_c3_rf_int_abt_msk_reg/NET0131 ,
		_w7267_
	);
	LUT4 #(
		.INIT('h8000)
	) name5039 (
		_w7264_,
		_w7265_,
		_w7266_,
		_w7267_,
		_w7268_
	);
	LUT2 #(
		.INIT('h7)
	) name5040 (
		_w7262_,
		_w7268_,
		_w7269_
	);
	LUT2 #(
		.INIT('h2)
	) name5041 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w3145_,
		_w7270_
	);
	LUT2 #(
		.INIT('h2)
	) name5042 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w3175_,
		_w7271_
	);
	LUT4 #(
		.INIT('h8000)
	) name5043 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ctl_rf_be_d1_reg[0]/P0001 ,
		_w3112_,
		_w6360_,
		_w7272_
	);
	LUT3 #(
		.INIT('h80)
	) name5044 (
		_w2232_,
		_w6360_,
		_w6408_,
		_w7273_
	);
	LUT4 #(
		.INIT('h0200)
	) name5045 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[20]_pad ,
		_w7274_
	);
	LUT3 #(
		.INIT('h02)
	) name5046 (
		_w6701_,
		_w6702_,
		_w7274_,
		_w7275_
	);
	LUT3 #(
		.INIT('h8a)
	) name5047 (
		\hwdata[4]_pad ,
		_w6702_,
		_w6704_,
		_w7276_
	);
	LUT4 #(
		.INIT('h0100)
	) name5048 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[28]_pad ,
		_w7277_
	);
	LUT3 #(
		.INIT('hab)
	) name5049 (
		_w6702_,
		_w7274_,
		_w7277_,
		_w7278_
	);
	LUT4 #(
		.INIT('h1011)
	) name5050 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7275_,
		_w7276_,
		_w7278_,
		_w7279_
	);
	LUT4 #(
		.INIT('h0200)
	) name5051 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[16]_pad ,
		_w7280_
	);
	LUT3 #(
		.INIT('h02)
	) name5052 (
		_w6701_,
		_w6702_,
		_w7280_,
		_w7281_
	);
	LUT3 #(
		.INIT('h8a)
	) name5053 (
		\hwdata[0]_pad ,
		_w6702_,
		_w6704_,
		_w7282_
	);
	LUT4 #(
		.INIT('h0100)
	) name5054 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[24]_pad ,
		_w7283_
	);
	LUT3 #(
		.INIT('hab)
	) name5055 (
		_w6702_,
		_w7280_,
		_w7283_,
		_w7284_
	);
	LUT4 #(
		.INIT('h1011)
	) name5056 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7281_,
		_w7282_,
		_w7284_,
		_w7285_
	);
	LUT4 #(
		.INIT('h0200)
	) name5057 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[3]_pad ,
		_w7286_
	);
	LUT3 #(
		.INIT('h02)
	) name5058 (
		_w6701_,
		_w6702_,
		_w7286_,
		_w7287_
	);
	LUT3 #(
		.INIT('h8a)
	) name5059 (
		\hwdata[19]_pad ,
		_w6702_,
		_w6704_,
		_w7288_
	);
	LUT4 #(
		.INIT('h0100)
	) name5060 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[11]_pad ,
		_w7289_
	);
	LUT3 #(
		.INIT('hab)
	) name5061 (
		_w6702_,
		_w7286_,
		_w7289_,
		_w7290_
	);
	LUT4 #(
		.INIT('h1011)
	) name5062 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7287_,
		_w7288_,
		_w7290_,
		_w7291_
	);
	LUT4 #(
		.INIT('h0200)
	) name5063 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[7]_pad ,
		_w7292_
	);
	LUT3 #(
		.INIT('h02)
	) name5064 (
		_w6701_,
		_w6702_,
		_w7292_,
		_w7293_
	);
	LUT3 #(
		.INIT('h8a)
	) name5065 (
		\hwdata[23]_pad ,
		_w6702_,
		_w6704_,
		_w7294_
	);
	LUT4 #(
		.INIT('h0100)
	) name5066 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[15]_pad ,
		_w7295_
	);
	LUT3 #(
		.INIT('hab)
	) name5067 (
		_w6702_,
		_w7292_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('h1011)
	) name5068 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7293_,
		_w7294_,
		_w7296_,
		_w7297_
	);
	LUT4 #(
		.INIT('h0200)
	) name5069 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[26]_pad ,
		_w7298_
	);
	LUT3 #(
		.INIT('h02)
	) name5070 (
		_w6701_,
		_w6702_,
		_w7298_,
		_w7299_
	);
	LUT3 #(
		.INIT('h8a)
	) name5071 (
		\hwdata[10]_pad ,
		_w6702_,
		_w6704_,
		_w7300_
	);
	LUT4 #(
		.INIT('h0100)
	) name5072 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[18]_pad ,
		_w7301_
	);
	LUT3 #(
		.INIT('hab)
	) name5073 (
		_w6702_,
		_w7298_,
		_w7301_,
		_w7302_
	);
	LUT4 #(
		.INIT('h1011)
	) name5074 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7299_,
		_w7300_,
		_w7302_,
		_w7303_
	);
	LUT4 #(
		.INIT('h0200)
	) name5075 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[27]_pad ,
		_w7304_
	);
	LUT3 #(
		.INIT('h02)
	) name5076 (
		_w6701_,
		_w6702_,
		_w7304_,
		_w7305_
	);
	LUT3 #(
		.INIT('h8a)
	) name5077 (
		\hwdata[11]_pad ,
		_w6702_,
		_w6704_,
		_w7306_
	);
	LUT4 #(
		.INIT('h0100)
	) name5078 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[19]_pad ,
		_w7307_
	);
	LUT3 #(
		.INIT('hab)
	) name5079 (
		_w6702_,
		_w7304_,
		_w7307_,
		_w7308_
	);
	LUT4 #(
		.INIT('h1011)
	) name5080 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7305_,
		_w7306_,
		_w7308_,
		_w7309_
	);
	LUT4 #(
		.INIT('h0200)
	) name5081 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[28]_pad ,
		_w7310_
	);
	LUT3 #(
		.INIT('h02)
	) name5082 (
		_w6701_,
		_w6702_,
		_w7310_,
		_w7311_
	);
	LUT3 #(
		.INIT('h8a)
	) name5083 (
		\hwdata[12]_pad ,
		_w6702_,
		_w6704_,
		_w7312_
	);
	LUT4 #(
		.INIT('h0100)
	) name5084 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[20]_pad ,
		_w7313_
	);
	LUT3 #(
		.INIT('hab)
	) name5085 (
		_w6702_,
		_w7310_,
		_w7313_,
		_w7314_
	);
	LUT4 #(
		.INIT('h1011)
	) name5086 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7311_,
		_w7312_,
		_w7314_,
		_w7315_
	);
	LUT4 #(
		.INIT('h0200)
	) name5087 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[29]_pad ,
		_w7316_
	);
	LUT3 #(
		.INIT('h02)
	) name5088 (
		_w6701_,
		_w6702_,
		_w7316_,
		_w7317_
	);
	LUT3 #(
		.INIT('h8a)
	) name5089 (
		\hwdata[13]_pad ,
		_w6702_,
		_w6704_,
		_w7318_
	);
	LUT4 #(
		.INIT('h0100)
	) name5090 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[21]_pad ,
		_w7319_
	);
	LUT3 #(
		.INIT('hab)
	) name5091 (
		_w6702_,
		_w7316_,
		_w7319_,
		_w7320_
	);
	LUT4 #(
		.INIT('h1011)
	) name5092 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7317_,
		_w7318_,
		_w7320_,
		_w7321_
	);
	LUT4 #(
		.INIT('h0200)
	) name5093 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[30]_pad ,
		_w7322_
	);
	LUT3 #(
		.INIT('h02)
	) name5094 (
		_w6701_,
		_w6702_,
		_w7322_,
		_w7323_
	);
	LUT3 #(
		.INIT('h8a)
	) name5095 (
		\hwdata[14]_pad ,
		_w6702_,
		_w6704_,
		_w7324_
	);
	LUT4 #(
		.INIT('h0100)
	) name5096 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[22]_pad ,
		_w7325_
	);
	LUT3 #(
		.INIT('hab)
	) name5097 (
		_w6702_,
		_w7322_,
		_w7325_,
		_w7326_
	);
	LUT4 #(
		.INIT('h1011)
	) name5098 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7323_,
		_w7324_,
		_w7326_,
		_w7327_
	);
	LUT4 #(
		.INIT('h0200)
	) name5099 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[10]_pad ,
		_w7328_
	);
	LUT3 #(
		.INIT('h02)
	) name5100 (
		_w6701_,
		_w6702_,
		_w7328_,
		_w7329_
	);
	LUT3 #(
		.INIT('h8a)
	) name5101 (
		\hwdata[26]_pad ,
		_w6702_,
		_w6704_,
		_w7330_
	);
	LUT4 #(
		.INIT('h0100)
	) name5102 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[2]_pad ,
		_w7331_
	);
	LUT3 #(
		.INIT('hab)
	) name5103 (
		_w6702_,
		_w7328_,
		_w7331_,
		_w7332_
	);
	LUT4 #(
		.INIT('h1011)
	) name5104 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7329_,
		_w7330_,
		_w7332_,
		_w7333_
	);
	LUT4 #(
		.INIT('h0200)
	) name5105 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[31]_pad ,
		_w7334_
	);
	LUT3 #(
		.INIT('h02)
	) name5106 (
		_w6701_,
		_w6702_,
		_w7334_,
		_w7335_
	);
	LUT3 #(
		.INIT('h8a)
	) name5107 (
		\hwdata[15]_pad ,
		_w6702_,
		_w6704_,
		_w7336_
	);
	LUT4 #(
		.INIT('h0100)
	) name5108 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[23]_pad ,
		_w7337_
	);
	LUT3 #(
		.INIT('hab)
	) name5109 (
		_w6702_,
		_w7334_,
		_w7337_,
		_w7338_
	);
	LUT4 #(
		.INIT('h1011)
	) name5110 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7335_,
		_w7336_,
		_w7338_,
		_w7339_
	);
	LUT4 #(
		.INIT('h0200)
	) name5111 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[0]_pad ,
		_w7340_
	);
	LUT3 #(
		.INIT('h02)
	) name5112 (
		_w6701_,
		_w6702_,
		_w7340_,
		_w7341_
	);
	LUT3 #(
		.INIT('h8a)
	) name5113 (
		\hwdata[16]_pad ,
		_w6702_,
		_w6704_,
		_w7342_
	);
	LUT4 #(
		.INIT('h0100)
	) name5114 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[8]_pad ,
		_w7343_
	);
	LUT3 #(
		.INIT('hab)
	) name5115 (
		_w6702_,
		_w7340_,
		_w7343_,
		_w7344_
	);
	LUT4 #(
		.INIT('h1011)
	) name5116 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7341_,
		_w7342_,
		_w7344_,
		_w7345_
	);
	LUT4 #(
		.INIT('h0200)
	) name5117 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[1]_pad ,
		_w7346_
	);
	LUT3 #(
		.INIT('h02)
	) name5118 (
		_w6701_,
		_w6702_,
		_w7346_,
		_w7347_
	);
	LUT3 #(
		.INIT('h8a)
	) name5119 (
		\hwdata[17]_pad ,
		_w6702_,
		_w6704_,
		_w7348_
	);
	LUT4 #(
		.INIT('h0100)
	) name5120 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[9]_pad ,
		_w7349_
	);
	LUT3 #(
		.INIT('hab)
	) name5121 (
		_w6702_,
		_w7346_,
		_w7349_,
		_w7350_
	);
	LUT4 #(
		.INIT('h1011)
	) name5122 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7347_,
		_w7348_,
		_w7350_,
		_w7351_
	);
	LUT4 #(
		.INIT('h0200)
	) name5123 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[2]_pad ,
		_w7352_
	);
	LUT3 #(
		.INIT('h02)
	) name5124 (
		_w6701_,
		_w6702_,
		_w7352_,
		_w7353_
	);
	LUT3 #(
		.INIT('h8a)
	) name5125 (
		\hwdata[18]_pad ,
		_w6702_,
		_w6704_,
		_w7354_
	);
	LUT4 #(
		.INIT('h0100)
	) name5126 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[10]_pad ,
		_w7355_
	);
	LUT3 #(
		.INIT('hab)
	) name5127 (
		_w6702_,
		_w7352_,
		_w7355_,
		_w7356_
	);
	LUT4 #(
		.INIT('h1011)
	) name5128 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7353_,
		_w7354_,
		_w7356_,
		_w7357_
	);
	LUT4 #(
		.INIT('h0200)
	) name5129 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[17]_pad ,
		_w7358_
	);
	LUT3 #(
		.INIT('h02)
	) name5130 (
		_w6701_,
		_w6702_,
		_w7358_,
		_w7359_
	);
	LUT3 #(
		.INIT('h8a)
	) name5131 (
		\hwdata[1]_pad ,
		_w6702_,
		_w6704_,
		_w7360_
	);
	LUT4 #(
		.INIT('h0100)
	) name5132 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[25]_pad ,
		_w7361_
	);
	LUT3 #(
		.INIT('hab)
	) name5133 (
		_w6702_,
		_w7358_,
		_w7361_,
		_w7362_
	);
	LUT4 #(
		.INIT('h1011)
	) name5134 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7359_,
		_w7360_,
		_w7362_,
		_w7363_
	);
	LUT4 #(
		.INIT('h0200)
	) name5135 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[4]_pad ,
		_w7364_
	);
	LUT3 #(
		.INIT('h02)
	) name5136 (
		_w6701_,
		_w6702_,
		_w7364_,
		_w7365_
	);
	LUT3 #(
		.INIT('h8a)
	) name5137 (
		\hwdata[20]_pad ,
		_w6702_,
		_w6704_,
		_w7366_
	);
	LUT4 #(
		.INIT('h0100)
	) name5138 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[12]_pad ,
		_w7367_
	);
	LUT3 #(
		.INIT('hab)
	) name5139 (
		_w6702_,
		_w7364_,
		_w7367_,
		_w7368_
	);
	LUT4 #(
		.INIT('h1011)
	) name5140 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7365_,
		_w7366_,
		_w7368_,
		_w7369_
	);
	LUT4 #(
		.INIT('h0200)
	) name5141 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[5]_pad ,
		_w7370_
	);
	LUT3 #(
		.INIT('h02)
	) name5142 (
		_w6701_,
		_w6702_,
		_w7370_,
		_w7371_
	);
	LUT3 #(
		.INIT('h8a)
	) name5143 (
		\hwdata[21]_pad ,
		_w6702_,
		_w6704_,
		_w7372_
	);
	LUT4 #(
		.INIT('h0100)
	) name5144 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[13]_pad ,
		_w7373_
	);
	LUT3 #(
		.INIT('hab)
	) name5145 (
		_w6702_,
		_w7370_,
		_w7373_,
		_w7374_
	);
	LUT4 #(
		.INIT('h1011)
	) name5146 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7371_,
		_w7372_,
		_w7374_,
		_w7375_
	);
	LUT4 #(
		.INIT('h0200)
	) name5147 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[6]_pad ,
		_w7376_
	);
	LUT3 #(
		.INIT('h02)
	) name5148 (
		_w6701_,
		_w6702_,
		_w7376_,
		_w7377_
	);
	LUT3 #(
		.INIT('h8a)
	) name5149 (
		\hwdata[22]_pad ,
		_w6702_,
		_w6704_,
		_w7378_
	);
	LUT4 #(
		.INIT('h0100)
	) name5150 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[14]_pad ,
		_w7379_
	);
	LUT3 #(
		.INIT('hab)
	) name5151 (
		_w6702_,
		_w7376_,
		_w7379_,
		_w7380_
	);
	LUT4 #(
		.INIT('h1011)
	) name5152 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7377_,
		_w7378_,
		_w7380_,
		_w7381_
	);
	LUT4 #(
		.INIT('h0200)
	) name5153 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[8]_pad ,
		_w7382_
	);
	LUT3 #(
		.INIT('h02)
	) name5154 (
		_w6701_,
		_w6702_,
		_w7382_,
		_w7383_
	);
	LUT3 #(
		.INIT('h8a)
	) name5155 (
		\hwdata[24]_pad ,
		_w6702_,
		_w6704_,
		_w7384_
	);
	LUT4 #(
		.INIT('h0100)
	) name5156 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[0]_pad ,
		_w7385_
	);
	LUT3 #(
		.INIT('hab)
	) name5157 (
		_w6702_,
		_w7382_,
		_w7385_,
		_w7386_
	);
	LUT4 #(
		.INIT('h1011)
	) name5158 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7383_,
		_w7384_,
		_w7386_,
		_w7387_
	);
	LUT4 #(
		.INIT('h0200)
	) name5159 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[11]_pad ,
		_w7388_
	);
	LUT3 #(
		.INIT('h02)
	) name5160 (
		_w6701_,
		_w6702_,
		_w7388_,
		_w7389_
	);
	LUT3 #(
		.INIT('h8a)
	) name5161 (
		\hwdata[27]_pad ,
		_w6702_,
		_w6704_,
		_w7390_
	);
	LUT4 #(
		.INIT('h0100)
	) name5162 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[3]_pad ,
		_w7391_
	);
	LUT3 #(
		.INIT('hab)
	) name5163 (
		_w6702_,
		_w7388_,
		_w7391_,
		_w7392_
	);
	LUT4 #(
		.INIT('h1011)
	) name5164 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7389_,
		_w7390_,
		_w7392_,
		_w7393_
	);
	LUT4 #(
		.INIT('h0200)
	) name5165 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[12]_pad ,
		_w7394_
	);
	LUT3 #(
		.INIT('h02)
	) name5166 (
		_w6701_,
		_w6702_,
		_w7394_,
		_w7395_
	);
	LUT3 #(
		.INIT('h8a)
	) name5167 (
		\hwdata[28]_pad ,
		_w6702_,
		_w6704_,
		_w7396_
	);
	LUT4 #(
		.INIT('h0100)
	) name5168 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[4]_pad ,
		_w7397_
	);
	LUT3 #(
		.INIT('hab)
	) name5169 (
		_w6702_,
		_w7394_,
		_w7397_,
		_w7398_
	);
	LUT4 #(
		.INIT('h1011)
	) name5170 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7395_,
		_w7396_,
		_w7398_,
		_w7399_
	);
	LUT4 #(
		.INIT('h0200)
	) name5171 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[18]_pad ,
		_w7400_
	);
	LUT3 #(
		.INIT('h02)
	) name5172 (
		_w6701_,
		_w6702_,
		_w7400_,
		_w7401_
	);
	LUT3 #(
		.INIT('h8a)
	) name5173 (
		\hwdata[2]_pad ,
		_w6702_,
		_w6704_,
		_w7402_
	);
	LUT4 #(
		.INIT('h0100)
	) name5174 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[26]_pad ,
		_w7403_
	);
	LUT3 #(
		.INIT('hab)
	) name5175 (
		_w6702_,
		_w7400_,
		_w7403_,
		_w7404_
	);
	LUT4 #(
		.INIT('h1011)
	) name5176 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7401_,
		_w7402_,
		_w7404_,
		_w7405_
	);
	LUT4 #(
		.INIT('h0200)
	) name5177 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[14]_pad ,
		_w7406_
	);
	LUT3 #(
		.INIT('h02)
	) name5178 (
		_w6701_,
		_w6702_,
		_w7406_,
		_w7407_
	);
	LUT3 #(
		.INIT('h8a)
	) name5179 (
		\hwdata[30]_pad ,
		_w6702_,
		_w6704_,
		_w7408_
	);
	LUT4 #(
		.INIT('h0100)
	) name5180 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[6]_pad ,
		_w7409_
	);
	LUT3 #(
		.INIT('hab)
	) name5181 (
		_w6702_,
		_w7406_,
		_w7409_,
		_w7410_
	);
	LUT4 #(
		.INIT('h1011)
	) name5182 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7407_,
		_w7408_,
		_w7410_,
		_w7411_
	);
	LUT4 #(
		.INIT('h0200)
	) name5183 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[15]_pad ,
		_w7412_
	);
	LUT3 #(
		.INIT('h02)
	) name5184 (
		_w6701_,
		_w6702_,
		_w7412_,
		_w7413_
	);
	LUT3 #(
		.INIT('h8a)
	) name5185 (
		\hwdata[31]_pad ,
		_w6702_,
		_w6704_,
		_w7414_
	);
	LUT4 #(
		.INIT('h0100)
	) name5186 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[7]_pad ,
		_w7415_
	);
	LUT3 #(
		.INIT('hab)
	) name5187 (
		_w6702_,
		_w7412_,
		_w7415_,
		_w7416_
	);
	LUT4 #(
		.INIT('h1011)
	) name5188 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7413_,
		_w7414_,
		_w7416_,
		_w7417_
	);
	LUT4 #(
		.INIT('h0200)
	) name5189 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[21]_pad ,
		_w7418_
	);
	LUT3 #(
		.INIT('h02)
	) name5190 (
		_w6701_,
		_w6702_,
		_w7418_,
		_w7419_
	);
	LUT3 #(
		.INIT('h8a)
	) name5191 (
		\hwdata[5]_pad ,
		_w6702_,
		_w6704_,
		_w7420_
	);
	LUT4 #(
		.INIT('h0100)
	) name5192 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[29]_pad ,
		_w7421_
	);
	LUT3 #(
		.INIT('hab)
	) name5193 (
		_w6702_,
		_w7418_,
		_w7421_,
		_w7422_
	);
	LUT4 #(
		.INIT('h1011)
	) name5194 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7419_,
		_w7420_,
		_w7422_,
		_w7423_
	);
	LUT4 #(
		.INIT('h0200)
	) name5195 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[22]_pad ,
		_w7424_
	);
	LUT3 #(
		.INIT('h02)
	) name5196 (
		_w6701_,
		_w6702_,
		_w7424_,
		_w7425_
	);
	LUT3 #(
		.INIT('h8a)
	) name5197 (
		\hwdata[6]_pad ,
		_w6702_,
		_w6704_,
		_w7426_
	);
	LUT4 #(
		.INIT('h0100)
	) name5198 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[30]_pad ,
		_w7427_
	);
	LUT3 #(
		.INIT('hab)
	) name5199 (
		_w6702_,
		_w7424_,
		_w7427_,
		_w7428_
	);
	LUT4 #(
		.INIT('h1011)
	) name5200 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7425_,
		_w7426_,
		_w7428_,
		_w7429_
	);
	LUT4 #(
		.INIT('h0200)
	) name5201 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[23]_pad ,
		_w7430_
	);
	LUT3 #(
		.INIT('h02)
	) name5202 (
		_w6701_,
		_w6702_,
		_w7430_,
		_w7431_
	);
	LUT3 #(
		.INIT('h8a)
	) name5203 (
		\hwdata[7]_pad ,
		_w6702_,
		_w6704_,
		_w7432_
	);
	LUT4 #(
		.INIT('h0100)
	) name5204 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[31]_pad ,
		_w7433_
	);
	LUT3 #(
		.INIT('hab)
	) name5205 (
		_w6702_,
		_w7430_,
		_w7433_,
		_w7434_
	);
	LUT4 #(
		.INIT('h1011)
	) name5206 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7431_,
		_w7432_,
		_w7434_,
		_w7435_
	);
	LUT4 #(
		.INIT('h0200)
	) name5207 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[24]_pad ,
		_w7436_
	);
	LUT3 #(
		.INIT('h02)
	) name5208 (
		_w6701_,
		_w6702_,
		_w7436_,
		_w7437_
	);
	LUT3 #(
		.INIT('h8a)
	) name5209 (
		\hwdata[8]_pad ,
		_w6702_,
		_w6704_,
		_w7438_
	);
	LUT4 #(
		.INIT('h0100)
	) name5210 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[16]_pad ,
		_w7439_
	);
	LUT3 #(
		.INIT('hab)
	) name5211 (
		_w6702_,
		_w7436_,
		_w7439_,
		_w7440_
	);
	LUT4 #(
		.INIT('h1011)
	) name5212 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7437_,
		_w7438_,
		_w7440_,
		_w7441_
	);
	LUT4 #(
		.INIT('h0200)
	) name5213 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[25]_pad ,
		_w7442_
	);
	LUT3 #(
		.INIT('h02)
	) name5214 (
		_w6701_,
		_w6702_,
		_w7442_,
		_w7443_
	);
	LUT3 #(
		.INIT('h8a)
	) name5215 (
		\hwdata[9]_pad ,
		_w6702_,
		_w6704_,
		_w7444_
	);
	LUT4 #(
		.INIT('h0100)
	) name5216 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[17]_pad ,
		_w7445_
	);
	LUT3 #(
		.INIT('hab)
	) name5217 (
		_w6702_,
		_w7442_,
		_w7445_,
		_w7446_
	);
	LUT4 #(
		.INIT('h1011)
	) name5218 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7443_,
		_w7444_,
		_w7446_,
		_w7447_
	);
	LUT4 #(
		.INIT('h0200)
	) name5219 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[9]_pad ,
		_w7448_
	);
	LUT3 #(
		.INIT('h02)
	) name5220 (
		_w6701_,
		_w6702_,
		_w7448_,
		_w7449_
	);
	LUT3 #(
		.INIT('h8a)
	) name5221 (
		\hwdata[25]_pad ,
		_w6702_,
		_w6704_,
		_w7450_
	);
	LUT4 #(
		.INIT('h0100)
	) name5222 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[1]_pad ,
		_w7451_
	);
	LUT3 #(
		.INIT('hab)
	) name5223 (
		_w6702_,
		_w7448_,
		_w7451_,
		_w7452_
	);
	LUT4 #(
		.INIT('h1011)
	) name5224 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7449_,
		_w7450_,
		_w7452_,
		_w7453_
	);
	LUT4 #(
		.INIT('h0200)
	) name5225 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[13]_pad ,
		_w7454_
	);
	LUT3 #(
		.INIT('h02)
	) name5226 (
		_w6701_,
		_w6702_,
		_w7454_,
		_w7455_
	);
	LUT3 #(
		.INIT('h8a)
	) name5227 (
		\hwdata[29]_pad ,
		_w6702_,
		_w6704_,
		_w7456_
	);
	LUT4 #(
		.INIT('h0100)
	) name5228 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[5]_pad ,
		_w7457_
	);
	LUT3 #(
		.INIT('hab)
	) name5229 (
		_w6702_,
		_w7454_,
		_w7457_,
		_w7458_
	);
	LUT4 #(
		.INIT('h1011)
	) name5230 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7455_,
		_w7456_,
		_w7458_,
		_w7459_
	);
	LUT4 #(
		.INIT('h0200)
	) name5231 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[19]_pad ,
		_w7460_
	);
	LUT3 #(
		.INIT('h02)
	) name5232 (
		_w6701_,
		_w6702_,
		_w7460_,
		_w7461_
	);
	LUT3 #(
		.INIT('h8a)
	) name5233 (
		\hwdata[3]_pad ,
		_w6702_,
		_w6704_,
		_w7462_
	);
	LUT4 #(
		.INIT('h0100)
	) name5234 (
		\ahb_slv_slv_sz_d1o_reg[0]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[1]/NET0131 ,
		\ahb_slv_slv_sz_d1o_reg[2]/NET0131 ,
		\hwdata[27]_pad ,
		_w7463_
	);
	LUT3 #(
		.INIT('hab)
	) name5235 (
		_w6702_,
		_w7460_,
		_w7463_,
		_w7464_
	);
	LUT4 #(
		.INIT('h1011)
	) name5236 (
		\de_m0_arb_st_reg/NET0131 ,
		_w7461_,
		_w7462_,
		_w7464_,
		_w7465_
	);
	LUT3 #(
		.INIT('h10)
	) name5237 (
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\ctl_rf_rf_sel_d1_reg/NET0131 ,
		_w7466_
	);
	LUT4 #(
		.INIT('h1000)
	) name5238 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w7467_
	);
	LUT3 #(
		.INIT('h10)
	) name5239 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w7468_
	);
	LUT3 #(
		.INIT('h80)
	) name5240 (
		_w7466_,
		_w7467_,
		_w7468_,
		_w7469_
	);
	LUT4 #(
		.INIT('h2000)
	) name5241 (
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w7470_
	);
	LUT3 #(
		.INIT('h20)
	) name5242 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w7471_
	);
	LUT3 #(
		.INIT('h80)
	) name5243 (
		_w7466_,
		_w7470_,
		_w7471_,
		_w7472_
	);
	LUT4 #(
		.INIT('h1000)
	) name5244 (
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w7473_
	);
	LUT3 #(
		.INIT('h80)
	) name5245 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w7474_
	);
	LUT3 #(
		.INIT('h80)
	) name5246 (
		_w7466_,
		_w7473_,
		_w7474_,
		_w7475_
	);
	LUT3 #(
		.INIT('h80)
	) name5247 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7476_
	);
	LUT3 #(
		.INIT('h80)
	) name5248 (
		_w7466_,
		_w7473_,
		_w7476_,
		_w7477_
	);
	LUT4 #(
		.INIT('h0400)
	) name5249 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w7478_
	);
	LUT3 #(
		.INIT('h80)
	) name5250 (
		_w6362_,
		_w7466_,
		_w7478_,
		_w7479_
	);
	LUT3 #(
		.INIT('h40)
	) name5251 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7480_
	);
	LUT3 #(
		.INIT('h80)
	) name5252 (
		_w7466_,
		_w7478_,
		_w7480_,
		_w7481_
	);
	LUT3 #(
		.INIT('h10)
	) name5253 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7482_
	);
	LUT3 #(
		.INIT('h80)
	) name5254 (
		_w7466_,
		_w7467_,
		_w7482_,
		_w7483_
	);
	LUT3 #(
		.INIT('h20)
	) name5255 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7484_
	);
	LUT3 #(
		.INIT('h80)
	) name5256 (
		_w7466_,
		_w7470_,
		_w7484_,
		_w7485_
	);
	LUT4 #(
		.INIT('h1011)
	) name5257 (
		_w2472_,
		_w7281_,
		_w7282_,
		_w7284_,
		_w7486_
	);
	LUT4 #(
		.INIT('h1011)
	) name5258 (
		_w2472_,
		_w7455_,
		_w7456_,
		_w7458_,
		_w7487_
	);
	LUT4 #(
		.INIT('h1011)
	) name5259 (
		_w2472_,
		_w7401_,
		_w7402_,
		_w7404_,
		_w7488_
	);
	LUT4 #(
		.INIT('h1011)
	) name5260 (
		_w2472_,
		_w7413_,
		_w7414_,
		_w7416_,
		_w7489_
	);
	LUT4 #(
		.INIT('h1011)
	) name5261 (
		_w2472_,
		_w7347_,
		_w7348_,
		_w7350_,
		_w7490_
	);
	LUT4 #(
		.INIT('h1011)
	) name5262 (
		_w2472_,
		_w7449_,
		_w7450_,
		_w7452_,
		_w7491_
	);
	LUT4 #(
		.INIT('h1011)
	) name5263 (
		_w2472_,
		_w7461_,
		_w7462_,
		_w7464_,
		_w7492_
	);
	LUT4 #(
		.INIT('h1011)
	) name5264 (
		_w2472_,
		_w7335_,
		_w7336_,
		_w7338_,
		_w7493_
	);
	LUT4 #(
		.INIT('h1011)
	) name5265 (
		_w2472_,
		_w7407_,
		_w7408_,
		_w7410_,
		_w7494_
	);
	LUT4 #(
		.INIT('h1011)
	) name5266 (
		_w2472_,
		_w7395_,
		_w7396_,
		_w7398_,
		_w7495_
	);
	LUT4 #(
		.INIT('h1011)
	) name5267 (
		_w2472_,
		_w7419_,
		_w7420_,
		_w7422_,
		_w7496_
	);
	LUT4 #(
		.INIT('h1011)
	) name5268 (
		_w2472_,
		_w7317_,
		_w7318_,
		_w7320_,
		_w7497_
	);
	LUT4 #(
		.INIT('h1011)
	) name5269 (
		_w2472_,
		_w7431_,
		_w7432_,
		_w7434_,
		_w7498_
	);
	LUT4 #(
		.INIT('h1011)
	) name5270 (
		_w2472_,
		_w7425_,
		_w7426_,
		_w7428_,
		_w7499_
	);
	LUT4 #(
		.INIT('h1011)
	) name5271 (
		_w2472_,
		_w7437_,
		_w7438_,
		_w7440_,
		_w7500_
	);
	LUT4 #(
		.INIT('h1011)
	) name5272 (
		_w2472_,
		_w7299_,
		_w7300_,
		_w7302_,
		_w7501_
	);
	LUT4 #(
		.INIT('h1011)
	) name5273 (
		_w2472_,
		_w7341_,
		_w7342_,
		_w7344_,
		_w7502_
	);
	LUT4 #(
		.INIT('h1011)
	) name5274 (
		_w2472_,
		_w7389_,
		_w7390_,
		_w7392_,
		_w7503_
	);
	LUT4 #(
		.INIT('h1011)
	) name5275 (
		_w2472_,
		_w7287_,
		_w7288_,
		_w7290_,
		_w7504_
	);
	LUT4 #(
		.INIT('h1011)
	) name5276 (
		_w2472_,
		_w7311_,
		_w7312_,
		_w7314_,
		_w7505_
	);
	LUT4 #(
		.INIT('h1011)
	) name5277 (
		_w2472_,
		_w7353_,
		_w7354_,
		_w7356_,
		_w7506_
	);
	LUT4 #(
		.INIT('h1011)
	) name5278 (
		_w2472_,
		_w7293_,
		_w7294_,
		_w7296_,
		_w7507_
	);
	LUT4 #(
		.INIT('h1011)
	) name5279 (
		_w2472_,
		_w7371_,
		_w7372_,
		_w7374_,
		_w7508_
	);
	LUT4 #(
		.INIT('h1011)
	) name5280 (
		_w2472_,
		_w7329_,
		_w7330_,
		_w7332_,
		_w7509_
	);
	LUT4 #(
		.INIT('h1011)
	) name5281 (
		_w2472_,
		_w7305_,
		_w7306_,
		_w7308_,
		_w7510_
	);
	LUT4 #(
		.INIT('h1011)
	) name5282 (
		_w2472_,
		_w7323_,
		_w7324_,
		_w7326_,
		_w7511_
	);
	LUT4 #(
		.INIT('h1011)
	) name5283 (
		_w2472_,
		_w7359_,
		_w7360_,
		_w7362_,
		_w7512_
	);
	LUT4 #(
		.INIT('h1011)
	) name5284 (
		_w2472_,
		_w7365_,
		_w7366_,
		_w7368_,
		_w7513_
	);
	LUT4 #(
		.INIT('h1011)
	) name5285 (
		_w2472_,
		_w7377_,
		_w7378_,
		_w7380_,
		_w7514_
	);
	LUT4 #(
		.INIT('h1011)
	) name5286 (
		_w2472_,
		_w7383_,
		_w7384_,
		_w7386_,
		_w7515_
	);
	LUT4 #(
		.INIT('h1011)
	) name5287 (
		_w2472_,
		_w7275_,
		_w7276_,
		_w7278_,
		_w7516_
	);
	LUT4 #(
		.INIT('h1011)
	) name5288 (
		_w2472_,
		_w7443_,
		_w7444_,
		_w7446_,
		_w7517_
	);
	LUT4 #(
		.INIT('h8000)
	) name5289 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w2239_,
		_w2249_,
		_w7518_
	);
	LUT3 #(
		.INIT('h80)
	) name5290 (
		_w6362_,
		_w7466_,
		_w7467_,
		_w7519_
	);
	LUT4 #(
		.INIT('h8000)
	) name5291 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w5230_,
		_w5248_,
		_w7520_
	);
	LUT3 #(
		.INIT('h80)
	) name5292 (
		_w7466_,
		_w7468_,
		_w7478_,
		_w7521_
	);
	LUT3 #(
		.INIT('h80)
	) name5293 (
		_w7466_,
		_w7478_,
		_w7482_,
		_w7522_
	);
	LUT4 #(
		.INIT('h8000)
	) name5294 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2229_,
		_w2232_,
		_w2239_,
		_w7523_
	);
	LUT3 #(
		.INIT('h80)
	) name5295 (
		_w7466_,
		_w7473_,
		_w7484_,
		_w7524_
	);
	LUT4 #(
		.INIT('h0800)
	) name5296 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\ahb_slv_slv_wr_d1o_reg/NET0131 ,
		_w7525_
	);
	LUT3 #(
		.INIT('h80)
	) name5297 (
		_w7466_,
		_w7480_,
		_w7525_,
		_w7526_
	);
	LUT4 #(
		.INIT('h8000)
	) name5298 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2239_,
		_w2244_,
		_w2249_,
		_w7527_
	);
	LUT3 #(
		.INIT('h80)
	) name5299 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7528_
	);
	LUT3 #(
		.INIT('h80)
	) name5300 (
		_w7466_,
		_w7478_,
		_w7528_,
		_w7529_
	);
	LUT3 #(
		.INIT('h80)
	) name5301 (
		_w7466_,
		_w7525_,
		_w7528_,
		_w7530_
	);
	LUT4 #(
		.INIT('h8000)
	) name5302 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2244_,
		_w5230_,
		_w5248_,
		_w7531_
	);
	LUT3 #(
		.INIT('h20)
	) name5303 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w7532_
	);
	LUT3 #(
		.INIT('h80)
	) name5304 (
		_w7466_,
		_w7467_,
		_w7532_,
		_w7533_
	);
	LUT3 #(
		.INIT('h20)
	) name5305 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w7534_
	);
	LUT3 #(
		.INIT('h80)
	) name5306 (
		_w7466_,
		_w7467_,
		_w7534_,
		_w7535_
	);
	LUT3 #(
		.INIT('h80)
	) name5307 (
		_w7466_,
		_w7478_,
		_w7532_,
		_w7536_
	);
	LUT4 #(
		.INIT('h8000)
	) name5308 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2232_,
		_w2239_,
		_w2244_,
		_w7537_
	);
	LUT3 #(
		.INIT('h80)
	) name5309 (
		_w7466_,
		_w7525_,
		_w7532_,
		_w7538_
	);
	LUT3 #(
		.INIT('h80)
	) name5310 (
		_w7466_,
		_w7525_,
		_w7534_,
		_w7539_
	);
	LUT4 #(
		.INIT('h8000)
	) name5311 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2247_,
		_w5230_,
		_w5248_,
		_w7540_
	);
	LUT4 #(
		.INIT('h8000)
	) name5312 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2232_,
		_w2239_,
		_w2247_,
		_w7541_
	);
	LUT3 #(
		.INIT('h80)
	) name5313 (
		_w7466_,
		_w7478_,
		_w7534_,
		_w7542_
	);
	LUT4 #(
		.INIT('h8000)
	) name5314 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2247_,
		_w5230_,
		_w5231_,
		_w7543_
	);
	LUT3 #(
		.INIT('h80)
	) name5315 (
		_w7466_,
		_w7471_,
		_w7473_,
		_w7544_
	);
	LUT3 #(
		.INIT('h80)
	) name5316 (
		_w6362_,
		_w7466_,
		_w7525_,
		_w7545_
	);
	LUT4 #(
		.INIT('h8000)
	) name5317 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2248_,
		_w2254_,
		_w5258_,
		_w7546_
	);
	LUT3 #(
		.INIT('h80)
	) name5318 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\ctl_rf_be_d1_reg[2]/P0001 ,
		_w7547_
	);
	LUT3 #(
		.INIT('h80)
	) name5319 (
		_w7466_,
		_w7467_,
		_w7547_,
		_w7548_
	);
	LUT3 #(
		.INIT('h80)
	) name5320 (
		_w7466_,
		_w7467_,
		_w7528_,
		_w7549_
	);
	LUT3 #(
		.INIT('h80)
	) name5321 (
		_w7466_,
		_w7478_,
		_w7547_,
		_w7550_
	);
	LUT4 #(
		.INIT('h8000)
	) name5322 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2232_,
		_w2239_,
		_w2254_,
		_w7551_
	);
	LUT4 #(
		.INIT('h8000)
	) name5323 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2231_,
		_w2254_,
		_w5258_,
		_w7552_
	);
	LUT3 #(
		.INIT('h80)
	) name5324 (
		_w7466_,
		_w7467_,
		_w7480_,
		_w7553_
	);
	LUT3 #(
		.INIT('h80)
	) name5325 (
		_w7466_,
		_w7468_,
		_w7525_,
		_w7554_
	);
	LUT3 #(
		.INIT('h80)
	) name5326 (
		_w7466_,
		_w7525_,
		_w7547_,
		_w7555_
	);
	LUT3 #(
		.INIT('h80)
	) name5327 (
		_w7466_,
		_w7470_,
		_w7476_,
		_w7556_
	);
	LUT3 #(
		.INIT('h80)
	) name5328 (
		_w7466_,
		_w7470_,
		_w7474_,
		_w7557_
	);
	LUT3 #(
		.INIT('h80)
	) name5329 (
		_w7466_,
		_w7482_,
		_w7525_,
		_w7558_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5330 (
		\ctl_rf_c0_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c0_rf_chllp_on_reg/NET0131 ,
		_w3086_,
		_w3091_,
		_w7559_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5331 (
		\ctl_rf_c1_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c1_rf_chllp_on_reg/NET0131 ,
		_w3041_,
		_w3046_,
		_w7560_
	);
	LUT4 #(
		.INIT('h8000)
	) name5332 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2229_,
		_w5230_,
		_w5231_,
		_w7561_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5333 (
		\ctl_rf_c2_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c2_rf_chllp_on_reg/NET0131 ,
		_w3019_,
		_w3024_,
		_w7562_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5334 (
		\ctl_rf_c3_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c3_rf_chllp_on_reg/NET0131 ,
		_w3052_,
		_w3057_,
		_w7563_
	);
	LUT4 #(
		.INIT('h8000)
	) name5335 (
		\ctl_rf_be_d1_reg[1]/P0001 ,
		_w2244_,
		_w5230_,
		_w5231_,
		_w7564_
	);
	LUT4 #(
		.INIT('h8000)
	) name5336 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2239_,
		_w2247_,
		_w2249_,
		_w7565_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5337 (
		\ctl_rf_c4_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c4_rf_chllp_on_reg/NET0131 ,
		_w3030_,
		_w3035_,
		_w7566_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5338 (
		\ctl_rf_c5_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c5_rf_chllp_on_reg/NET0131 ,
		_w3075_,
		_w3080_,
		_w7567_
	);
	LUT4 #(
		.INIT('h8000)
	) name5339 (
		\ctl_rf_be_d1_reg[3]/P0001 ,
		_w2239_,
		_w2249_,
		_w2254_,
		_w7568_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5340 (
		\ctl_rf_c6_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c6_rf_chllp_on_reg/NET0131 ,
		_w3097_,
		_w3102_,
		_w7569_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5341 (
		\ctl_rf_c7_rf_ch_en_reg/NET0131 ,
		\ctl_rf_c7_rf_chllp_on_reg/NET0131 ,
		_w3064_,
		_w3069_,
		_w7570_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name5342 (
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[6]/NET0131 ,
		\de_m0_is_llp_reg/NET0131 ,
		_w7571_
	);
	LUT4 #(
		.INIT('h2000)
	) name5343 (
		\ahb_mst0_m0_m1_diff_tx_reg/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\h0readyin_pad ,
		_w7572_
	);
	LUT4 #(
		.INIT('hffc4)
	) name5344 (
		\h0readyin_pad ,
		\h0write_pad ,
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT2 #(
		.INIT('he)
	) name5345 (
		_w5359_,
		_w5360_,
		_w7574_
	);
	LUT2 #(
		.INIT('he)
	) name5346 (
		_w2344_,
		_w2345_,
		_w7575_
	);
	LUT2 #(
		.INIT('he)
	) name5347 (
		_w5652_,
		_w5653_,
		_w7576_
	);
	LUT2 #(
		.INIT('he)
	) name5348 (
		_w5655_,
		_w5656_,
		_w7577_
	);
	LUT2 #(
		.INIT('he)
	) name5349 (
		_w5658_,
		_w5659_,
		_w7578_
	);
	LUT2 #(
		.INIT('he)
	) name5350 (
		_w5661_,
		_w5662_,
		_w7579_
	);
	LUT2 #(
		.INIT('he)
	) name5351 (
		_w5916_,
		_w5917_,
		_w7580_
	);
	LUT2 #(
		.INIT('he)
	) name5352 (
		_w5362_,
		_w5363_,
		_w7581_
	);
	LUT2 #(
		.INIT('he)
	) name5353 (
		_w5920_,
		_w5921_,
		_w7582_
	);
	LUT2 #(
		.INIT('he)
	) name5354 (
		_w2260_,
		_w2261_,
		_w7583_
	);
	LUT2 #(
		.INIT('he)
	) name5355 (
		_w5375_,
		_w5376_,
		_w7584_
	);
	LUT2 #(
		.INIT('he)
	) name5356 (
		_w5275_,
		_w5276_,
		_w7585_
	);
	LUT2 #(
		.INIT('he)
	) name5357 (
		_w5233_,
		_w5234_,
		_w7586_
	);
	LUT2 #(
		.INIT('he)
	) name5358 (
		_w5236_,
		_w5237_,
		_w7587_
	);
	LUT2 #(
		.INIT('he)
	) name5359 (
		_w2236_,
		_w2237_,
		_w7588_
	);
	LUT2 #(
		.INIT('he)
	) name5360 (
		_w5296_,
		_w5297_,
		_w7589_
	);
	LUT2 #(
		.INIT('he)
	) name5361 (
		_w5305_,
		_w5306_,
		_w7590_
	);
	LUT2 #(
		.INIT('he)
	) name5362 (
		_w2371_,
		_w2372_,
		_w7591_
	);
	LUT2 #(
		.INIT('he)
	) name5363 (
		_w5292_,
		_w5293_,
		_w7592_
	);
	LUT2 #(
		.INIT('he)
	) name5364 (
		_w2241_,
		_w2242_,
		_w7593_
	);
	LUT2 #(
		.INIT('he)
	) name5365 (
		_w2295_,
		_w2296_,
		_w7594_
	);
	LUT2 #(
		.INIT('he)
	) name5366 (
		_w2298_,
		_w2299_,
		_w7595_
	);
	LUT2 #(
		.INIT('he)
	) name5367 (
		_w2341_,
		_w2342_,
		_w7596_
	);
	LUT2 #(
		.INIT('he)
	) name5368 (
		_w2282_,
		_w2283_,
		_w7597_
	);
	LUT2 #(
		.INIT('he)
	) name5369 (
		_w2323_,
		_w2324_,
		_w7598_
	);
	LUT2 #(
		.INIT('he)
	) name5370 (
		_w2331_,
		_w2332_,
		_w7599_
	);
	LUT2 #(
		.INIT('he)
	) name5371 (
		_w5370_,
		_w5371_,
		_w7600_
	);
	LUT2 #(
		.INIT('he)
	) name5372 (
		_w5289_,
		_w5290_,
		_w7601_
	);
	LUT2 #(
		.INIT('he)
	) name5373 (
		_w5300_,
		_w5301_,
		_w7602_
	);
	LUT2 #(
		.INIT('he)
	) name5374 (
		_w5367_,
		_w5368_,
		_w7603_
	);
	LUT2 #(
		.INIT('h6)
	) name5375 (
		\ahb_slv_slv_ad_d1o_reg[4]/NET0131 ,
		\haddr[4]_pad ,
		_w7604_
	);
	LUT2 #(
		.INIT('h6)
	) name5376 (
		\ahb_slv_slv_ad_d1o_reg[8]/NET0131 ,
		\haddr[8]_pad ,
		_w7605_
	);
	LUT3 #(
		.INIT('h80)
	) name5377 (
		hreadyin_pad,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w7606_
	);
	LUT3 #(
		.INIT('h10)
	) name5378 (
		_w7604_,
		_w7605_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h2)
	) name5379 (
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\haddr[7]_pad ,
		_w7608_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5380 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\haddr[3]_pad ,
		\haddr[5]_pad ,
		_w7609_
	);
	LUT2 #(
		.INIT('h4)
	) name5381 (
		_w7608_,
		_w7609_,
		_w7610_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5382 (
		\ahb_slv_slv_ad_d1o_reg[5]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[7]/NET0131 ,
		\haddr[5]_pad ,
		\haddr[7]_pad ,
		_w7611_
	);
	LUT4 #(
		.INIT('hf531)
	) name5383 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\haddr[2]_pad ,
		\haddr[6]_pad ,
		_w7612_
	);
	LUT3 #(
		.INIT('hb0)
	) name5384 (
		\ahb_slv_slv_ad_d1o_reg[2]/NET0131 ,
		\haddr[2]_pad ,
		hwrite_pad,
		_w7613_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name5385 (
		\ahb_slv_slv_ad_d1o_reg[3]/NET0131 ,
		\ahb_slv_slv_ad_d1o_reg[6]/NET0131 ,
		\haddr[3]_pad ,
		\haddr[6]_pad ,
		_w7614_
	);
	LUT4 #(
		.INIT('h8000)
	) name5386 (
		_w7611_,
		_w7612_,
		_w7613_,
		_w7614_,
		_w7615_
	);
	LUT3 #(
		.INIT('h7f)
	) name5387 (
		_w7607_,
		_w7610_,
		_w7615_,
		_w7616_
	);
	LUT2 #(
		.INIT('h4)
	) name5388 (
		\de_de_st_reg[5]/NET0131 ,
		\de_m0_arb_st_reg/NET0131 ,
		_w7617_
	);
	LUT3 #(
		.INIT('h40)
	) name5389 (
		\ch_sel_arb_chcsr_reg_reg[1]/NET0131 ,
		\ch_sel_arb_chcsr_reg_reg[2]/NET0131 ,
		\de_de_st_reg[1]/NET0131 ,
		_w7618_
	);
	LUT2 #(
		.INIT('he)
	) name5390 (
		_w7617_,
		_w7618_,
		_w7619_
	);
	LUT4 #(
		.INIT('hffcb)
	) name5391 (
		\haddr[1]_pad ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w7620_
	);
	LUT3 #(
		.INIT('h01)
	) name5392 (
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name5393 (
		\haddr[0]_pad ,
		\haddr[1]_pad ,
		_w7622_
	);
	LUT3 #(
		.INIT('hd5)
	) name5394 (
		_w7620_,
		_w7621_,
		_w7622_,
		_w7623_
	);
	LUT2 #(
		.INIT('h2)
	) name5395 (
		\haddr[0]_pad ,
		\haddr[1]_pad ,
		_w7624_
	);
	LUT3 #(
		.INIT('hd5)
	) name5396 (
		_w7620_,
		_w7621_,
		_w7624_,
		_w7625_
	);
	LUT4 #(
		.INIT('h0002)
	) name5397 (
		\haddr[1]_pad ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w7626_
	);
	LUT4 #(
		.INIT('hffc7)
	) name5398 (
		\haddr[1]_pad ,
		\hsize[0]_pad ,
		\hsize[1]_pad ,
		\hsize[2]_pad ,
		_w7627_
	);
	LUT3 #(
		.INIT('h4f)
	) name5399 (
		\haddr[0]_pad ,
		_w7626_,
		_w7627_,
		_w7628_
	);
	LUT3 #(
		.INIT('h8f)
	) name5400 (
		\haddr[0]_pad ,
		_w7626_,
		_w7627_,
		_w7629_
	);
	LUT4 #(
		.INIT('ha800)
	) name5401 (
		hreadyin_pad,
		hsel_br_pad,
		hsel_reg_pad,
		\htrans[1]_pad ,
		_w7630_
	);
	LUT2 #(
		.INIT('h8)
	) name5402 (
		\ch_sel_dma_reqd1_reg[5]/NET0131 ,
		\ctl_rf_sync_reg[5]/NET0131 ,
		_w7631_
	);
	LUT2 #(
		.INIT('h8)
	) name5403 (
		\ch_sel_dma_reqd1_reg[7]/NET0131 ,
		\ctl_rf_sync_reg[7]/NET0131 ,
		_w7632_
	);
	LUT2 #(
		.INIT('h8)
	) name5404 (
		\ch_sel_dma_reqd1_reg[1]/NET0131 ,
		\ctl_rf_sync_reg[1]/NET0131 ,
		_w7633_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		\ch_sel_dma_reqd1_reg[0]/NET0131 ,
		\ctl_rf_sync_reg[0]/NET0131 ,
		_w7634_
	);
	LUT2 #(
		.INIT('h8)
	) name5406 (
		\ch_sel_dma_reqd1_reg[4]/NET0131 ,
		\ctl_rf_sync_reg[4]/NET0131 ,
		_w7635_
	);
	LUT2 #(
		.INIT('h8)
	) name5407 (
		\ch_sel_dma_reqd1_reg[3]/NET0131 ,
		\ctl_rf_sync_reg[3]/NET0131 ,
		_w7636_
	);
	LUT2 #(
		.INIT('h8)
	) name5408 (
		\ch_sel_dma_reqd1_reg[6]/NET0131 ,
		\ctl_rf_sync_reg[6]/NET0131 ,
		_w7637_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\ch_sel_dma_reqd1_reg[2]/NET0131 ,
		\ctl_rf_sync_reg[2]/NET0131 ,
		_w7638_
	);
	LUT3 #(
		.INIT('hac)
	) name5410 (
		\ahb_mst0_mx_cmd_st_reg[1]/NET0131 ,
		\ahb_mst0_mx_dtp_reg/NET0131 ,
		\h0readyin_pad ,
		_w7639_
	);
	LUT3 #(
		.INIT('h5c)
	) name5411 (
		\de_de_st_reg[1]/NET0131 ,
		\de_de_st_reg[5]/NET0131 ,
		\de_st_rd_msk_reg/NET0131 ,
		_w7640_
	);
	LUT4 #(
		.INIT('heee2)
	) name5412 (
		\ctl_rf_c7_rf_chdad_reg[18]/NET0131 ,
		_w2257_,
		_w2295_,
		_w2296_,
		_w7641_
	);
	LUT4 #(
		.INIT('heee2)
	) name5413 (
		\ctl_rf_c7_rf_chdad_reg[19]/NET0131 ,
		_w2257_,
		_w2298_,
		_w2299_,
		_w7642_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5414 (
		\ctl_rf_c2_rf_chllp_reg[24]/NET0131 ,
		_w2344_,
		_w2345_,
		_w5882_,
		_w7643_
	);
	LUT4 #(
		.INIT('heee2)
	) name5415 (
		\ctl_rf_c1_rf_chsad_reg[18]/NET0131 ,
		_w2281_,
		_w2295_,
		_w2296_,
		_w7644_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5416 (
		\ctl_rf_c5_rf_chdad_reg[1]/NET0131 ,
		_w5359_,
		_w5360_,
		_w5449_,
		_w7645_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5417 (
		\ctl_rf_c5_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5254_,
		_w7646_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5418 (
		\ctl_rf_c5_rf_chtsz_reg[5]/NET0131 ,
		_w5233_,
		_w5234_,
		_w5254_,
		_w7647_
	);
	LUT4 #(
		.INIT('heee2)
	) name5419 (
		\ctl_rf_c5_rf_chtsz_reg[4]/NET0131 ,
		_w5254_,
		_w5275_,
		_w5276_,
		_w7648_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5420 (
		\ctl_rf_c6_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2291_,
		_w7649_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5421 (
		\ctl_rf_c7_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2293_,
		_w7650_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5422 (
		\ctl_rf_c3_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2285_,
		_w7651_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5423 (
		\ctl_rf_c4_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2287_,
		_w7652_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5424 (
		\ctl_rf_c5_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2289_,
		_w7653_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5425 (
		\ctl_rf_c1_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2281_,
		_w7654_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5426 (
		\ctl_rf_c0_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2319_,
		_w7655_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5427 (
		\ctl_rf_c2_rf_chsad_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w2321_,
		_w7656_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5428 (
		\ctl_rf_c4_rf_chtsz_reg[7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5249_,
		_w7657_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5429 (
		\ctl_rf_c2_rf_chsad_reg[15]/NET0131 ,
		_w2993_,
		_w2994_,
		_w5430_,
		_w7658_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5430 (
		\ctl_rf_c6_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5775_,
		_w7659_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5431 (
		\ctl_rf_c0_rf_chllp_reg[18]/NET0131 ,
		_w2295_,
		_w2296_,
		_w5907_,
		_w7660_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5432 (
		\ctl_rf_c6_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5775_,
		_w7661_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5433 (
		\ctl_rf_c0_rf_chllp_reg[22]/NET0131 ,
		_w2323_,
		_w2324_,
		_w5907_,
		_w7662_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5434 (
		\ctl_rf_c0_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5907_,
		_w7663_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5435 (
		\ctl_rf_c0_rf_chllp_reg[17]/NET0131 ,
		_w2241_,
		_w2242_,
		_w5907_,
		_w7664_
	);
	LUT4 #(
		.INIT('heee2)
	) name5436 (
		\ctl_rf_c1_rf_chsad_reg[19]/NET0131 ,
		_w2281_,
		_w2298_,
		_w2299_,
		_w7665_
	);
	LUT4 #(
		.INIT('heee2)
	) name5437 (
		\ctl_rf_c1_rf_chsad_reg[3]/NET0131 ,
		_w2233_,
		_w5375_,
		_w5376_,
		_w7666_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name5438 (
		\ctl_rf_c3_rf_chllp_reg[21]/NET0131 ,
		_w2282_,
		_w2283_,
		_w5678_,
		_w7667_
	);
	assign \_al_n1  = 1'b1;
	assign \g16/_0_  = _w2238_ ;
	assign \g58487/_0_  = _w2243_ ;
	assign \g58489/_0_  = _w2246_ ;
	assign \g58491/_0_  = _w2251_ ;
	assign \g58493/_0_  = _w2253_ ;
	assign \g58495/_0_  = _w2256_ ;
	assign \g58497/_0_  = _w2258_ ;
	assign \g58499/_0_  = _w2262_ ;
	assign \g58500/_0_  = _w2264_ ;
	assign \g58501/_0_  = _w2266_ ;
	assign \g58502/_0_  = _w2268_ ;
	assign \g58504/_0_  = _w2270_ ;
	assign \g58505/_0_  = _w2272_ ;
	assign \g58507/_0_  = _w2274_ ;
	assign \g58508/_0_  = _w2276_ ;
	assign \g58509/_0_  = _w2278_ ;
	assign \g58510/_0_  = _w2280_ ;
	assign \g58556/_0_  = _w2284_ ;
	assign \g58557/_0_  = _w2286_ ;
	assign \g58558/_0_  = _w2288_ ;
	assign \g58559/_0_  = _w2290_ ;
	assign \g58560/_0_  = _w2292_ ;
	assign \g58561/_0_  = _w2294_ ;
	assign \g58562/_0_  = _w2297_ ;
	assign \g58563/_0_  = _w2300_ ;
	assign \g58566/_0_  = _w2301_ ;
	assign \g58567/_0_  = _w2302_ ;
	assign \g58568/_0_  = _w2303_ ;
	assign \g58569/_0_  = _w2304_ ;
	assign \g58570/_0_  = _w2305_ ;
	assign \g58571/_0_  = _w2306_ ;
	assign \g58572/_0_  = _w2307_ ;
	assign \g58573/_0_  = _w2308_ ;
	assign \g58574/_0_  = _w2309_ ;
	assign \g58575/_0_  = _w2310_ ;
	assign \g58576/_0_  = _w2311_ ;
	assign \g58577/_0_  = _w2312_ ;
	assign \g58578/_0_  = _w2313_ ;
	assign \g58579/_0_  = _w2314_ ;
	assign \g58580/_0_  = _w2315_ ;
	assign \g58581/_0_  = _w2316_ ;
	assign \g58584/_0_  = _w2317_ ;
	assign \g58585/_0_  = _w2318_ ;
	assign \g58586/_0_  = _w2320_ ;
	assign \g58587/_0_  = _w2322_ ;
	assign \g58588/_0_  = _w2325_ ;
	assign \g58589/_0_  = _w2326_ ;
	assign \g58590/_0_  = _w2327_ ;
	assign \g58591/_0_  = _w2328_ ;
	assign \g58592/_0_  = _w2329_ ;
	assign \g58593/_0_  = _w2330_ ;
	assign \g58594/_0_  = _w2333_ ;
	assign \g58595/_0_  = _w2334_ ;
	assign \g58596/_0_  = _w2335_ ;
	assign \g58597/_0_  = _w2336_ ;
	assign \g58598/_0_  = _w2337_ ;
	assign \g58599/_0_  = _w2338_ ;
	assign \g58600/_0_  = _w2339_ ;
	assign \g58601/_0_  = _w2340_ ;
	assign \g58602/_0_  = _w2343_ ;
	assign \g58603/_0_  = _w2346_ ;
	assign \g58604/_0_  = _w2347_ ;
	assign \g58605/_0_  = _w2348_ ;
	assign \g58606/_0_  = _w2349_ ;
	assign \g58607/_0_  = _w2350_ ;
	assign \g58608/_0_  = _w2351_ ;
	assign \g58609/_0_  = _w2352_ ;
	assign \g58610/_0_  = _w2353_ ;
	assign \g58611/_0_  = _w2354_ ;
	assign \g58612/_0_  = _w2355_ ;
	assign \g58613/_0_  = _w2356_ ;
	assign \g58614/_0_  = _w2357_ ;
	assign \g58615/_0_  = _w2358_ ;
	assign \g58616/_0_  = _w2359_ ;
	assign \g58617/_0_  = _w2360_ ;
	assign \g58618/_0_  = _w2361_ ;
	assign \g58619/_0_  = _w2362_ ;
	assign \g58620/_0_  = _w2363_ ;
	assign \g58621/_0_  = _w2364_ ;
	assign \g58622/_0_  = _w2365_ ;
	assign \g58623/_0_  = _w2366_ ;
	assign \g58624/_0_  = _w2367_ ;
	assign \g58625/_0_  = _w2368_ ;
	assign \g58626/_0_  = _w2369_ ;
	assign \g58627/_0_  = _w2370_ ;
	assign \g58723/_0_  = _w2373_ ;
	assign \g58734/_0_  = _w2374_ ;
	assign \g58737/_0_  = _w2375_ ;
	assign \g58741/_0_  = _w2376_ ;
	assign \g58749/_0_  = _w2377_ ;
	assign \g58754/_0_  = _w2378_ ;
	assign \g58762/_0_  = _w2379_ ;
	assign \g58763/_0_  = _w2380_ ;
	assign \g58764/_0_  = _w2381_ ;
	assign \g58765/_0_  = _w2382_ ;
	assign \g58766/_0_  = _w2383_ ;
	assign \g58767/_0_  = _w2384_ ;
	assign \g58768/_0_  = _w2385_ ;
	assign \g58769/_0_  = _w2386_ ;
	assign \g58770/_0_  = _w2387_ ;
	assign \g58771/_0_  = _w2388_ ;
	assign \g59788/_0_  = _w2439_ ;
	assign \g59832/_0_  = _w2479_ ;
	assign \g59873/_0_  = _w2493_ ;
	assign \g59874/_0_  = _w2503_ ;
	assign \g59893/_0_  = _w2648_ ;
	assign \g59894/_0_  = _w2710_ ;
	assign \g59895/_0_  = _w2764_ ;
	assign \g59896/_0_  = _w2832_ ;
	assign \g59923/_0_  = _w2843_ ;
	assign \g60031/_0_  = _w2863_ ;
	assign \g60032/_0_  = _w2885_ ;
	assign \g60033/_0_  = _w2917_ ;
	assign \g60036/_0_  = _w2930_ ;
	assign \g60037/_0_  = _w2942_ ;
	assign \g60038/_0_  = _w2953_ ;
	assign \g60165/_0_  = _w2976_ ;
	assign \g60186/_2__syn_2  = _w2977_ ;
	assign \g60187/_0_  = _w2988_ ;
	assign \g60188/_0_  = _w2990_ ;
	assign \g60258/_0_  = _w3111_ ;
	assign \g60259/_0_  = _w3123_ ;
	assign \g60260/_0_  = _w3133_ ;
	assign \g60261/_0_  = _w3143_ ;
	assign \g60263/_0_  = _w3153_ ;
	assign \g60264/_0_  = _w3163_ ;
	assign \g60265/_0_  = _w3173_ ;
	assign \g60266/_0_  = _w3183_ ;
	assign \g60267/_0_  = _w3374_ ;
	assign \g60303/_3_  = _w3394_ ;
	assign \g60360/_0_  = _w3398_ ;
	assign \g60361/_0_  = _w3405_ ;
	assign \g60401/_00_  = _w3410_ ;
	assign \g60428/_0_  = _w3418_ ;
	assign \g60429/_0_  = _w3421_ ;
	assign \g60448/_0_  = _w3620_ ;
	assign \g60449/_0_  = _w3687_ ;
	assign \g60974/_0_  = _w3696_ ;
	assign \g61072/_0_  = _w3705_ ;
	assign \g61073/_0_  = _w3713_ ;
	assign \g61074/_0_  = _w3720_ ;
	assign \g61075/_0_  = _w3727_ ;
	assign \g61076/_0_  = _w3734_ ;
	assign \g61077/_0_  = _w3741_ ;
	assign \g61078/_0_  = _w3748_ ;
	assign \g61079/_0_  = _w3755_ ;
	assign \g61486/_0_  = _w3758_ ;
	assign \g61502/_3_  = _w3762_ ;
	assign \g61879/_0_  = _w3767_ ;
	assign \g62077/_0_  = _w3777_ ;
	assign \g62078/_0_  = _w3940_ ;
	assign \g62079/_0_  = _w3989_ ;
	assign \g62080/_0_  = _w4128_ ;
	assign \g62081/_0_  = _w4266_ ;
	assign \g62082/_0_  = _w4399_ ;
	assign \g62083/_0_  = _w4532_ ;
	assign \g62084/_0_  = _w4603_ ;
	assign \g62085/_0_  = _w4736_ ;
	assign \g62086/_0_  = _w4880_ ;
	assign \g62087/_0_  = _w4951_ ;
	assign \g62088/_0_  = _w5021_ ;
	assign \g62089/_0_  = _w5091_ ;
	assign \g62090/_0_  = _w5161_ ;
	assign \g62091/_0_  = _w5229_ ;
	assign \g62629/_0_  = _w5235_ ;
	assign \g62630/_0_  = _w5238_ ;
	assign \g62631/_0_  = _w5239_ ;
	assign \g62632/_0_  = _w5241_ ;
	assign \g62633/_0_  = _w5243_ ;
	assign \g62634/_0_  = _w5244_ ;
	assign \g62635/_0_  = _w5245_ ;
	assign \g62637/_0_  = _w5247_ ;
	assign \g62638/_0_  = _w5250_ ;
	assign \g62639/_0_  = _w5251_ ;
	assign \g62641/_0_  = _w5253_ ;
	assign \g62643/_0_  = _w5255_ ;
	assign \g62645/_0_  = _w5257_ ;
	assign \g62646/_0_  = _w5260_ ;
	assign \g62647/_0_  = _w5261_ ;
	assign \g62648/_0_  = _w5262_ ;
	assign \g62649/_0_  = _w5264_ ;
	assign \g62650/_0_  = _w5266_ ;
	assign \g62651/_0_  = _w5267_ ;
	assign \g62652/_0_  = _w5268_ ;
	assign \g62655/_0_  = _w5270_ ;
	assign \g62656/_0_  = _w5272_ ;
	assign \g62657/_0_  = _w5273_ ;
	assign \g62658/_0_  = _w5274_ ;
	assign \g62659/_0_  = _w5277_ ;
	assign \g62660/_0_  = _w5279_ ;
	assign \g62661/_0_  = _w5281_ ;
	assign \g62662/_0_  = _w5282_ ;
	assign \g62663/_0_  = _w5283_ ;
	assign \g62664/_0_  = _w5284_ ;
	assign \g62665/_0_  = _w5285_ ;
	assign \g62667/_0_  = _w5286_ ;
	assign \g62668/_0_  = _w5287_ ;
	assign \g62669/_0_  = _w5291_ ;
	assign \g62670/_0_  = _w5294_ ;
	assign \g62671/_0_  = _w5295_ ;
	assign \g62672/_0_  = _w5298_ ;
	assign \g62673/_0_  = _w5302_ ;
	assign \g62674/_0_  = _w5303_ ;
	assign \g62675/_0_  = _w5304_ ;
	assign \g62676/_0_  = _w5307_ ;
	assign \g62677/_0_  = _w5309_ ;
	assign \g62678/_0_  = _w5310_ ;
	assign \g62679/_0_  = _w5311_ ;
	assign \g62680/_0_  = _w5312_ ;
	assign \g62681/_0_  = _w5313_ ;
	assign \g62682/_0_  = _w5314_ ;
	assign \g62683/_0_  = _w5315_ ;
	assign \g62684/_0_  = _w5317_ ;
	assign \g62685/_0_  = _w5319_ ;
	assign \g62686/_0_  = _w5321_ ;
	assign \g62687/_0_  = _w5322_ ;
	assign \g62688/_0_  = _w5323_ ;
	assign \g62689/_0_  = _w5324_ ;
	assign \g62690/_0_  = _w5325_ ;
	assign \g62691/_0_  = _w5326_ ;
	assign \g62692/_0_  = _w5327_ ;
	assign \g62693/_0_  = _w5329_ ;
	assign \g62694/_0_  = _w5331_ ;
	assign \g62695/_0_  = _w5332_ ;
	assign \g62696/_0_  = _w5333_ ;
	assign \g62697/_0_  = _w5334_ ;
	assign \g62698/_0_  = _w5335_ ;
	assign \g62699/_0_  = _w5336_ ;
	assign \g62700/_0_  = _w5337_ ;
	assign \g62701/_0_  = _w5339_ ;
	assign \g62702/_0_  = _w5340_ ;
	assign \g62703/_0_  = _w5342_ ;
	assign \g62704/_0_  = _w5343_ ;
	assign \g62705/_0_  = _w5344_ ;
	assign \g62706/_0_  = _w5345_ ;
	assign \g62707/_0_  = _w5346_ ;
	assign \g62708/_0_  = _w5347_ ;
	assign \g62709/_0_  = _w5349_ ;
	assign \g62710/_0_  = _w5350_ ;
	assign \g62711/_0_  = _w5351_ ;
	assign \g62712/_0_  = _w5353_ ;
	assign \g62713/_0_  = _w5354_ ;
	assign \g62714/_0_  = _w5355_ ;
	assign \g62715/_0_  = _w5356_ ;
	assign \g62716/_0_  = _w5357_ ;
	assign \g62721/_0_  = _w5358_ ;
	assign \g62722/_0_  = _w5361_ ;
	assign \g62723/_0_  = _w5364_ ;
	assign \g62725/_0_  = _w5365_ ;
	assign \g62726/_0_  = _w5366_ ;
	assign \g62727/_0_  = _w5369_ ;
	assign \g62728/_0_  = _w5372_ ;
	assign \g62729/_0_  = _w5373_ ;
	assign \g62730/_0_  = _w5374_ ;
	assign \g62731/_0_  = _w5377_ ;
	assign \g62732/_0_  = _w5378_ ;
	assign \g62733/_0_  = _w5380_ ;
	assign \g62734/_0_  = _w5381_ ;
	assign \g62735/_0_  = _w5382_ ;
	assign \g62736/_0_  = _w5383_ ;
	assign \g62737/_0_  = _w5384_ ;
	assign \g62738/_0_  = _w5385_ ;
	assign \g62739/_0_  = _w5386_ ;
	assign \g62740/_0_  = _w5387_ ;
	assign \g62741/_0_  = _w5388_ ;
	assign \g62742/_0_  = _w5389_ ;
	assign \g62743/_0_  = _w5391_ ;
	assign \g62744/_0_  = _w5392_ ;
	assign \g62745/_0_  = _w5393_ ;
	assign \g62746/_0_  = _w5394_ ;
	assign \g62747/_0_  = _w5395_ ;
	assign \g62748/_0_  = _w5396_ ;
	assign \g62749/_0_  = _w5397_ ;
	assign \g62750/_0_  = _w5398_ ;
	assign \g62751/_0_  = _w5399_ ;
	assign \g62752/_0_  = _w5400_ ;
	assign \g62753/_0_  = _w5402_ ;
	assign \g62754/_0_  = _w5403_ ;
	assign \g62755/_0_  = _w5405_ ;
	assign \g62756/_0_  = _w5406_ ;
	assign \g62757/_0_  = _w5408_ ;
	assign \g62758/_0_  = _w5409_ ;
	assign \g62759/_0_  = _w5410_ ;
	assign \g62760/_0_  = _w5411_ ;
	assign \g62761/_0_  = _w5412_ ;
	assign \g62762/_0_  = _w5413_ ;
	assign \g62763/_0_  = _w5414_ ;
	assign \g62764/_0_  = _w5415_ ;
	assign \g62765/_0_  = _w5416_ ;
	assign \g62766/_0_  = _w5417_ ;
	assign \g62767/_0_  = _w5419_ ;
	assign \g62768/_0_  = _w5420_ ;
	assign \g62769/_0_  = _w5421_ ;
	assign \g62770/_0_  = _w5422_ ;
	assign \g62771/_0_  = _w5423_ ;
	assign \g62772/_0_  = _w5425_ ;
	assign \g62773/_0_  = _w5426_ ;
	assign \g62774/_0_  = _w5427_ ;
	assign \g62775/_0_  = _w5429_ ;
	assign \g62776/_0_  = _w5431_ ;
	assign \g62777/_0_  = _w5432_ ;
	assign \g62778/_0_  = _w5433_ ;
	assign \g62779/_0_  = _w5434_ ;
	assign \g62780/_0_  = _w5435_ ;
	assign \g62781/_0_  = _w5436_ ;
	assign \g62783/_0_  = _w5437_ ;
	assign \g62784/_0_  = _w5438_ ;
	assign \g62785/_0_  = _w5439_ ;
	assign \g62786/_0_  = _w5440_ ;
	assign \g62787/_0_  = _w5441_ ;
	assign \g62788/_0_  = _w5442_ ;
	assign \g62789/_0_  = _w5443_ ;
	assign \g62790/_0_  = _w5444_ ;
	assign \g62791/_0_  = _w5446_ ;
	assign \g62792/_0_  = _w5447_ ;
	assign \g62793/_0_  = _w5448_ ;
	assign \g62794/_0_  = _w5450_ ;
	assign \g62795/_0_  = _w5451_ ;
	assign \g62797/_0_  = _w5452_ ;
	assign \g62798/_0_  = _w5453_ ;
	assign \g62799/_0_  = _w5454_ ;
	assign \g62800/_0_  = _w5455_ ;
	assign \g62801/_0_  = _w5456_ ;
	assign \g62802/_0_  = _w5457_ ;
	assign \g62803/_0_  = _w5458_ ;
	assign \g62804/_0_  = _w5460_ ;
	assign \g62805/_0_  = _w5461_ ;
	assign \g62806/_0_  = _w5462_ ;
	assign \g62807/_0_  = _w5463_ ;
	assign \g62808/_0_  = _w5464_ ;
	assign \g62809/_0_  = _w5465_ ;
	assign \g62810/_0_  = _w5466_ ;
	assign \g62811/_0_  = _w5467_ ;
	assign \g62812/_0_  = _w5468_ ;
	assign \g62813/_0_  = _w5469_ ;
	assign \g62814/_0_  = _w5470_ ;
	assign \g62815/_0_  = _w5471_ ;
	assign \g62816/_0_  = _w5472_ ;
	assign \g62817/_0_  = _w5473_ ;
	assign \g62818/_0_  = _w5474_ ;
	assign \g63108/_0_  = _w5619_ ;
	assign \g63117/_0_  = _w5634_ ;
	assign \g63125/_0_  = _w5637_ ;
	assign \g63126/_0_  = _w5638_ ;
	assign \g63127/_0_  = _w5639_ ;
	assign \g63128/_0_  = _w5640_ ;
	assign \g63129/_0_  = _w5641_ ;
	assign \g63130/_0_  = _w5642_ ;
	assign \g63131/_0_  = _w5644_ ;
	assign \g63132/_0_  = _w5645_ ;
	assign \g63133/_0_  = _w5646_ ;
	assign \g63134/_0_  = _w5647_ ;
	assign \g63135/_0_  = _w5648_ ;
	assign \g63136/_0_  = _w5649_ ;
	assign \g63137/_0_  = _w5650_ ;
	assign \g63138/_0_  = _w5654_ ;
	assign \g63139/_0_  = _w5657_ ;
	assign \g63140/_0_  = _w5660_ ;
	assign \g63141/_0_  = _w5663_ ;
	assign \g63142/_0_  = _w5665_ ;
	assign \g63143/_0_  = _w5666_ ;
	assign \g63144/_0_  = _w5667_ ;
	assign \g63145/_0_  = _w5668_ ;
	assign \g63146/_0_  = _w5669_ ;
	assign \g63147/_0_  = _w5670_ ;
	assign \g63148/_0_  = _w5672_ ;
	assign \g63149/_0_  = _w5673_ ;
	assign \g63150/_0_  = _w5674_ ;
	assign \g63151/_0_  = _w5675_ ;
	assign \g63152/_0_  = _w5676_ ;
	assign \g63153/_0_  = _w5677_ ;
	assign \g63154/_0_  = _w5679_ ;
	assign \g63155/_0_  = _w5680_ ;
	assign \g63156/_0_  = _w5681_ ;
	assign \g63157/_0_  = _w5682_ ;
	assign \g63159/_0_  = _w5683_ ;
	assign \g63160/_0_  = _w5684_ ;
	assign \g63161/_0_  = _w5686_ ;
	assign \g63162/_0_  = _w5687_ ;
	assign \g63163/_0_  = _w5688_ ;
	assign \g63164/_0_  = _w5689_ ;
	assign \g63165/_0_  = _w5691_ ;
	assign \g63166/_0_  = _w5692_ ;
	assign \g63167/_0_  = _w5693_ ;
	assign \g63168/_0_  = _w5694_ ;
	assign \g63169/_0_  = _w5695_ ;
	assign \g63170/_0_  = _w5696_ ;
	assign \g63171/_0_  = _w5699_ ;
	assign \g63172/_0_  = _w5700_ ;
	assign \g63173/_0_  = _w5701_ ;
	assign \g63174/_0_  = _w5702_ ;
	assign \g63175/_0_  = _w5703_ ;
	assign \g63176/_0_  = _w5704_ ;
	assign \g63177/_0_  = _w5706_ ;
	assign \g63178/_0_  = _w5707_ ;
	assign \g63179/_0_  = _w5708_ ;
	assign \g63180/_0_  = _w5709_ ;
	assign \g63181/_0_  = _w5710_ ;
	assign \g63182/_0_  = _w5711_ ;
	assign \g63183/_0_  = _w5712_ ;
	assign \g63184/_0_  = _w5714_ ;
	assign \g63185/_0_  = _w5715_ ;
	assign \g63186/_0_  = _w5716_ ;
	assign \g63187/_0_  = _w5717_ ;
	assign \g63188/_0_  = _w5719_ ;
	assign \g63189/_0_  = _w5720_ ;
	assign \g63190/_0_  = _w5721_ ;
	assign \g63191/_0_  = _w5722_ ;
	assign \g63192/_0_  = _w5723_ ;
	assign \g63193/_0_  = _w5724_ ;
	assign \g63194/_0_  = _w5726_ ;
	assign \g63195/_0_  = _w5727_ ;
	assign \g63196/_0_  = _w5728_ ;
	assign \g63197/_0_  = _w5729_ ;
	assign \g63198/_0_  = _w5730_ ;
	assign \g63199/_0_  = _w5731_ ;
	assign \g63200/_0_  = _w5733_ ;
	assign \g63201/_0_  = _w5734_ ;
	assign \g63202/_0_  = _w5735_ ;
	assign \g63203/_0_  = _w5736_ ;
	assign \g63204/_0_  = _w5737_ ;
	assign \g63205/_0_  = _w5738_ ;
	assign \g63206/_0_  = _w5739_ ;
	assign \g63207/_0_  = _w5741_ ;
	assign \g63208/_0_  = _w5742_ ;
	assign \g63209/_0_  = _w5743_ ;
	assign \g63210/_0_  = _w5744_ ;
	assign \g63211/_0_  = _w5746_ ;
	assign \g63212/_0_  = _w5747_ ;
	assign \g63213/_0_  = _w5748_ ;
	assign \g63214/_0_  = _w5756_ ;
	assign \g63215/_0_  = _w5757_ ;
	assign \g63216/_0_  = _w5758_ ;
	assign \g63217/_0_  = _w5759_ ;
	assign \g63218/_0_  = _w5766_ ;
	assign \g63219/_0_  = _w5769_ ;
	assign \g63220/_0_  = _w5770_ ;
	assign \g63221/_0_  = _w5771_ ;
	assign \g63222/_0_  = _w5772_ ;
	assign \g63223/_0_  = _w5773_ ;
	assign \g63224/_0_  = _w5774_ ;
	assign \g63225/_0_  = _w5776_ ;
	assign \g63226/_0_  = _w5777_ ;
	assign \g63228/_0_  = _w5778_ ;
	assign \g63229/_0_  = _w5779_ ;
	assign \g63231/_0_  = _w5780_ ;
	assign \g63232/_0_  = _w5782_ ;
	assign \g63233/_0_  = _w5783_ ;
	assign \g63234/_0_  = _w5784_ ;
	assign \g63235/_0_  = _w5785_ ;
	assign \g63236/_0_  = _w5787_ ;
	assign \g63237/_0_  = _w5788_ ;
	assign \g63238/_0_  = _w5789_ ;
	assign \g63239/_0_  = _w5790_ ;
	assign \g63240/_0_  = _w5791_ ;
	assign \g63241/_0_  = _w5792_ ;
	assign \g63242/_0_  = _w5799_ ;
	assign \g63244/_0_  = _w5808_ ;
	assign \g63246/_0_  = _w5816_ ;
	assign \g63247/_0_  = _w5818_ ;
	assign \g63248/_0_  = _w5819_ ;
	assign \g63249/_0_  = _w5820_ ;
	assign \g63250/_0_  = _w5821_ ;
	assign \g63251/_0_  = _w5822_ ;
	assign \g63252/_0_  = _w5823_ ;
	assign \g63253/_0_  = _w5825_ ;
	assign \g63254/_0_  = _w5826_ ;
	assign \g63255/_0_  = _w5827_ ;
	assign \g63256/_0_  = _w5828_ ;
	assign \g63257/_0_  = _w5829_ ;
	assign \g63258/_0_  = _w5830_ ;
	assign \g63259/_0_  = _w5831_ ;
	assign \g63260/_0_  = _w5833_ ;
	assign \g63261/_0_  = _w5834_ ;
	assign \g63262/_0_  = _w5835_ ;
	assign \g63263/_0_  = _w5836_ ;
	assign \g63264/_0_  = _w5838_ ;
	assign \g63265/_0_  = _w5839_ ;
	assign \g63266/_0_  = _w5840_ ;
	assign \g63267/_0_  = _w5841_ ;
	assign \g63268/_0_  = _w5842_ ;
	assign \g63269/_0_  = _w5843_ ;
	assign \g63270/_0_  = _w5851_ ;
	assign \g63272/_0_  = _w5859_ ;
	assign \g63291/_0_  = _w5860_ ;
	assign \g63292/_0_  = _w5862_ ;
	assign \g63293/_0_  = _w5863_ ;
	assign \g63294/_0_  = _w5864_ ;
	assign \g63295/_0_  = _w5865_ ;
	assign \g63298/_0_  = _w5867_ ;
	assign \g63299/_0_  = _w5869_ ;
	assign \g63300/_0_  = _w5870_ ;
	assign \g63301/_0_  = _w5871_ ;
	assign \g63302/_0_  = _w5872_ ;
	assign \g63303/_0_  = _w5873_ ;
	assign \g63304/_0_  = _w5875_ ;
	assign \g63305/_0_  = _w5876_ ;
	assign \g63306/_0_  = _w5877_ ;
	assign \g63307/_0_  = _w5878_ ;
	assign \g63308/_0_  = _w5880_ ;
	assign \g63309/_0_  = _w5881_ ;
	assign \g63310/_0_  = _w5883_ ;
	assign \g63311/_0_  = _w5885_ ;
	assign \g63312/_0_  = _w5886_ ;
	assign \g63313/_0_  = _w5887_ ;
	assign \g63314/_0_  = _w5888_ ;
	assign \g63315/_0_  = _w5889_ ;
	assign \g63316/_0_  = _w5904_ ;
	assign \g63317/_0_  = _w5905_ ;
	assign \g63318/_0_  = _w5906_ ;
	assign \g63320/_0_  = _w5908_ ;
	assign \g63322/_0_  = _w5909_ ;
	assign \g63323/_0_  = _w5910_ ;
	assign \g63324/_0_  = _w5911_ ;
	assign \g63325/_0_  = _w5912_ ;
	assign \g63326/_0_  = _w5913_ ;
	assign \g63327/_0_  = _w5914_ ;
	assign \g63328/_0_  = _w5915_ ;
	assign \g63329/_0_  = _w5918_ ;
	assign \g63330/_0_  = _w5919_ ;
	assign \g63331/_0_  = _w5922_ ;
	assign \g63332/_0_  = _w5923_ ;
	assign \g63333/_0_  = _w5924_ ;
	assign \g63334/_0_  = _w5925_ ;
	assign \g63335/_0_  = _w5926_ ;
	assign \g63336/_0_  = _w5927_ ;
	assign \g63337/_0_  = _w5928_ ;
	assign \g63338/_0_  = _w5929_ ;
	assign \g63339/_0_  = _w5930_ ;
	assign \g63340/_0_  = _w5931_ ;
	assign \g63341/_0_  = _w5932_ ;
	assign \g63342/_0_  = _w5933_ ;
	assign \g63343/_0_  = _w5934_ ;
	assign \g63344/_0_  = _w5935_ ;
	assign \g63345/_0_  = _w5936_ ;
	assign \g63346/_0_  = _w5937_ ;
	assign \g63347/_0_  = _w5938_ ;
	assign \g63348/_0_  = _w5939_ ;
	assign \g63349/_0_  = _w5940_ ;
	assign \g63350/_0_  = _w5941_ ;
	assign \g63351/_0_  = _w5942_ ;
	assign \g63352/_0_  = _w5943_ ;
	assign \g63353/_0_  = _w5944_ ;
	assign \g63354/_0_  = _w5945_ ;
	assign \g63355/_0_  = _w5946_ ;
	assign \g63356/_0_  = _w5947_ ;
	assign \g63357/_0_  = _w5948_ ;
	assign \g63358/_0_  = _w5949_ ;
	assign \g63359/_0_  = _w5950_ ;
	assign \g63360/_0_  = _w5951_ ;
	assign \g63361/_0_  = _w5952_ ;
	assign \g63362/_0_  = _w5953_ ;
	assign \g63363/_0_  = _w5954_ ;
	assign \g63364/_0_  = _w5955_ ;
	assign \g63365/_0_  = _w5956_ ;
	assign \g63366/_0_  = _w5957_ ;
	assign \g63367/_0_  = _w5958_ ;
	assign \g63368/_0_  = _w5959_ ;
	assign \g63369/_0_  = _w5960_ ;
	assign \g63370/_0_  = _w5961_ ;
	assign \g63371/_0_  = _w5962_ ;
	assign \g63372/_0_  = _w5963_ ;
	assign \g63373/_0_  = _w5964_ ;
	assign \g63374/_0_  = _w5965_ ;
	assign \g63375/_0_  = _w5966_ ;
	assign \g63376/_0_  = _w5967_ ;
	assign \g63377/_0_  = _w5968_ ;
	assign \g63378/_0_  = _w5969_ ;
	assign \g63379/_0_  = _w5970_ ;
	assign \g63380/_0_  = _w5971_ ;
	assign \g63383/_3_  = _w5976_ ;
	assign \g63386/_0_  = _w5977_ ;
	assign \g63387/_0_  = _w5978_ ;
	assign \g63388/_0_  = _w5979_ ;
	assign \g63389/_0_  = _w5980_ ;
	assign \g63390/_0_  = _w5981_ ;
	assign \g63391/_0_  = _w5982_ ;
	assign \g63392/_0_  = _w5983_ ;
	assign \g63419/_0_  = _w5984_ ;
	assign \g63421/_0_  = _w5985_ ;
	assign \g63422/_0_  = _w5986_ ;
	assign \g63423/_0_  = _w5987_ ;
	assign \g63424/_0_  = _w5988_ ;
	assign \g63425/_0_  = _w5989_ ;
	assign \g63536/_3_  = _w5997_ ;
	assign \g63625/_0_  = _w5998_ ;
	assign \g63628/_0_  = _w5618_ ;
	assign \g63871/_0_  = _w6006_ ;
	assign \g63874/_0_  = _w2573_ ;
	assign \g63889/_0_  = _w6010_ ;
	assign \g63933/_0_  = _w6018_ ;
	assign \g63945/_0_  = _w6026_ ;
	assign \g63959/_0_  = _w6035_ ;
	assign \g63962/_0_  = _w6043_ ;
	assign \g63974/_0_  = _w6051_ ;
	assign \g63977/_0_  = _w6058_ ;
	assign \g64035/_0_  = _w6066_ ;
	assign \g64435/_3_  = _w6071_ ;
	assign \g64939/_0_  = _w6079_ ;
	assign \g65149/_0_  = _w6087_ ;
	assign \g65632/_3_  = _w6091_ ;
	assign \g65633/_0_  = _w6094_ ;
	assign \g65634/_0_  = _w6097_ ;
	assign \g65635/_0_  = _w6099_ ;
	assign \g65636/_0_  = _w6101_ ;
	assign \g65638/_3_  = _w6103_ ;
	assign \g65640/_3_  = _w6105_ ;
	assign \g65999/_0_  = _w6110_ ;
	assign \g66912/_0_  = _w6115_ ;
	assign \g66914/_0_  = _w6124_ ;
	assign \g67555/_3_  = _w6125_ ;
	assign \g67564/_3_  = _w6126_ ;
	assign \g67567/_3_  = _w6127_ ;
	assign \g67735/_0_  = _w6132_ ;
	assign \g67736/_0_  = _w6136_ ;
	assign \g67737/_0_  = _w6140_ ;
	assign \g67738/_0_  = _w6144_ ;
	assign \g67758/_0_  = _w6148_ ;
	assign \g67760/_0_  = _w6152_ ;
	assign \g67761/_0_  = _w6156_ ;
	assign \g67763/_0_  = _w6160_ ;
	assign \g67766/_0_  = _w6164_ ;
	assign \g67810/_0_  = _w6181_ ;
	assign \g67816/_0_  = _w6188_ ;
	assign \g67902/_0_  = _w6190_ ;
	assign \g67927/_0_  = _w6195_ ;
	assign \g67936/_0_  = _w6198_ ;
	assign \g68067/_0_  = _w6209_ ;
	assign \g68068/_0_  = _w6213_ ;
	assign \g68069/_0_  = _w6224_ ;
	assign \g68070/_0_  = _w6228_ ;
	assign \g68071/_0_  = _w6239_ ;
	assign \g68072/_0_  = _w6243_ ;
	assign \g68073/_0_  = _w6254_ ;
	assign \g68074/_0_  = _w6258_ ;
	assign \g68075/_0_  = _w6269_ ;
	assign \g68076/_0_  = _w6273_ ;
	assign \g68077/_0_  = _w6284_ ;
	assign \g68078/_0_  = _w6288_ ;
	assign \g68079/_0_  = _w6299_ ;
	assign \g68080/_0_  = _w6303_ ;
	assign \g68081/_0_  = _w6314_ ;
	assign \g68082/_0_  = _w6318_ ;
	assign \g68083/_0_  = _w6322_ ;
	assign \g68084/_0_  = _w6324_ ;
	assign \g68085/_0_  = _w6326_ ;
	assign \g68086/_0_  = _w6328_ ;
	assign \g68087/_0_  = _w6330_ ;
	assign \g68088/_0_  = _w6332_ ;
	assign \g68089/_0_  = _w6334_ ;
	assign \g68090/_0_  = _w6336_ ;
	assign \g68091/_0_  = _w6338_ ;
	assign \g68096/_0_  = _w6340_ ;
	assign \g68160/_0_  = _w6342_ ;
	assign \g68218/_0_  = _w6344_ ;
	assign \g68219/_0_  = _w6346_ ;
	assign \g68220/_0_  = _w6348_ ;
	assign \g68221/_0_  = _w6350_ ;
	assign \g68222/_0_  = _w6352_ ;
	assign \g68226/_0_  = _w6354_ ;
	assign \g68247/_0_  = _w6358_ ;
	assign \g68252/_0_  = _w6359_ ;
	assign \g68632/_0_  = _w6366_ ;
	assign \g68633/_0_  = _w6370_ ;
	assign \g68635/_0_  = _w6374_ ;
	assign \g68640/_0_  = _w6378_ ;
	assign \g68642/_0_  = _w6382_ ;
	assign \g68643/_0_  = _w6386_ ;
	assign \g68644/_0_  = _w6390_ ;
	assign \g68645/_0_  = _w6394_ ;
	assign \g68649/_0_  = _w6400_ ;
	assign \g68668/_2_  = _w6402_ ;
	assign \g68670/_0_  = _w6407_ ;
	assign \g68681/_3_  = _w6414_ ;
	assign \g68689/_0_  = _w6420_ ;
	assign \g68690/_0_  = _w6426_ ;
	assign \g68691/_0_  = _w6432_ ;
	assign \g68692/_0_  = _w6438_ ;
	assign \g68693/_0_  = _w6444_ ;
	assign \g68694/_0_  = _w6450_ ;
	assign \g68695/_0_  = _w6456_ ;
	assign \g68737/_0_  = _w6469_ ;
	assign \g68742/_0_  = _w6482_ ;
	assign \g68745/_0_  = _w6495_ ;
	assign \g68750/_0_  = _w6508_ ;
	assign \g68759/_0_  = _w6521_ ;
	assign \g68761/_0_  = _w6534_ ;
	assign \g68774/_0_  = _w3239_ ;
	assign \g68775/_0_  = _w3338_ ;
	assign \g68776/_0_  = _w3310_ ;
	assign \g68777/_0_  = _w3211_ ;
	assign \g68778/_0_  = _w3254_ ;
	assign \g68780/_0_  = _w3352_ ;
	assign \g68781/_0_  = _w3324_ ;
	assign \g68782/_0_  = _w3370_ ;
	assign \g68783/_0_  = _w3295_ ;
	assign \g68784/_0_  = _w3281_ ;
	assign \g68785/_0_  = _w3225_ ;
	assign \g68786/_0_  = _w3197_ ;
	assign \g68787/_0_  = _w6547_ ;
	assign \g68790/_0_  = _w6560_ ;
	assign \g68791/_0_  = _w6573_ ;
	assign \g68793/_0_  = _w6586_ ;
	assign \g68794/_0_  = _w6599_ ;
	assign \g68795/_0_  = _w6612_ ;
	assign \g68796/_0_  = _w6625_ ;
	assign \g68797/_0_  = _w6638_ ;
	assign \g68804/_0_  = _w6651_ ;
	assign \g68805/_0_  = _w6664_ ;
	assign \g68807/_0_  = _w6677_ ;
	assign \g68809/_0_  = _w6690_ ;
	assign \g68864/_3_  = _w6730_ ;
	assign \g68865/_3_  = _w6764_ ;
	assign \g68866/_3_  = _w6798_ ;
	assign \g68867/_3_  = _w6832_ ;
	assign \g68868/_3_  = _w6866_ ;
	assign \g68869/_3_  = _w6900_ ;
	assign \g68870/_3_  = _w6934_ ;
	assign \g68871/_3_  = _w6948_ ;
	assign \g68872/_3_  = _w6982_ ;
	assign \g68873/_3_  = _w6996_ ;
	assign \g68874/_3_  = _w7010_ ;
	assign \g68875/_3_  = _w7024_ ;
	assign \g68876/_3_  = _w7038_ ;
	assign \g68877/_3_  = _w7042_ ;
	assign \g68878/_3_  = _w7056_ ;
	assign \g68879/_3_  = _w7070_ ;
	assign \g68880/_3_  = _w7084_ ;
	assign \g68881/_3_  = _w7088_ ;
	assign \g68882/_3_  = _w7092_ ;
	assign \g68883/_3_  = _w7096_ ;
	assign \g68884/_3_  = _w7100_ ;
	assign \g68885/_3_  = _w7104_ ;
	assign \g68886/_3_  = _w7108_ ;
	assign \g68887/_3_  = _w7112_ ;
	assign \g68888/_3_  = _w7116_ ;
	assign \g68889/_3_  = _w7120_ ;
	assign \g68890/_3_  = _w7124_ ;
	assign \g68891/_3_  = _w7128_ ;
	assign \g68892/_3_  = _w7132_ ;
	assign \g68893/_3_  = _w7136_ ;
	assign \g68894/_3_  = _w7140_ ;
	assign \g68895/_3_  = _w7144_ ;
	assign \g69037/_1__syn_2  = _w6403_ ;
	assign \g69077/_0_  = _w7149_ ;
	assign \g69081/_0_  = _w7154_ ;
	assign \g69084/_0_  = _w7157_ ;
	assign \g69085/_0_  = _w7162_ ;
	assign \g69086/_0_  = _w7167_ ;
	assign \g69088/_0_  = _w7172_ ;
	assign \g69094/_0_  = _w7177_ ;
	assign \g69095/_0_  = _w7182_ ;
	assign \g69097/_0_  = _w7187_ ;
	assign \g69114/_3_  = _w7192_ ;
	assign \g69116/_3_  = _w7197_ ;
	assign \g69118/_3_  = _w7202_ ;
	assign \g69120/_3_  = _w7207_ ;
	assign \g69122/_3_  = _w7212_ ;
	assign \g69124/_3_  = _w7217_ ;
	assign \g69126/_3_  = _w7222_ ;
	assign \g69128/_3_  = _w7227_ ;
	assign \g69581/_3_  = _w5535_ ;
	assign \g70303/_1__syn_2  = _w7228_ ;
	assign \g70304/_1__syn_2  = _w7229_ ;
	assign \g70305/_1__syn_2  = _w7230_ ;
	assign \g70306/_1__syn_2  = _w7231_ ;
	assign \g70353/_1__syn_2  = _w7232_ ;
	assign \g70359/_2_  = _w7233_ ;
	assign \g70364/_1__syn_2  = _w7234_ ;
	assign \g70375/_1__syn_2  = _w7235_ ;
	assign \g70380/_2_  = _w7236_ ;
	assign \g70383/_1__syn_2  = _w7237_ ;
	assign \g70394/_2_  = _w7238_ ;
	assign \g70395/_2_  = _w3119_ ;
	assign \g70396/_1__syn_2  = _w7239_ ;
	assign \g70398/_1__syn_2  = _w7240_ ;
	assign \g70407/_1_  = _w7241_ ;
	assign \g70416/_1__syn_2  = _w7242_ ;
	assign \g70418/_1__syn_2  = _w7243_ ;
	assign \g70419/_2_  = _w3140_ ;
	assign \g70424/_1_  = _w7244_ ;
	assign \g70465/_2_  = _w7245_ ;
	assign \g70511/_1_  = _w7246_ ;
	assign \g70512/_1_  = _w7247_ ;
	assign \g70513/_2_  = _w7248_ ;
	assign \g70514/_2_  = _w3107_ ;
	assign \g70516/_2_  = _w7249_ ;
	assign \g70518/_2_  = _w7250_ ;
	assign \g70519/_2_  = _w3130_ ;
	assign \g70520/_2_  = _w7251_ ;
	assign \g70530/_2_  = _w7252_ ;
	assign \g70534/_3_  = _w5606_ ;
	assign \g70536/_3_  = _w5614_ ;
	assign \g70540/_3_  = _w5502_ ;
	assign \g70541/_2_  = _w7253_ ;
	assign \g70545/_3_  = _w5527_ ;
	assign \g70546/_2_  = _w7254_ ;
	assign \g70547/_2_  = _w3150_ ;
	assign \g70550/_3_  = _w5570_ ;
	assign \g70551/_2_  = _w7255_ ;
	assign \g70552/_2_  = _w3160_ ;
	assign \g70558/_3_  = _w5562_ ;
	assign \g70559/_2_  = _w3170_ ;
	assign \g70560/_2_  = _w7256_ ;
	assign \g70562/_3_  = _w5493_ ;
	assign \g70564/_3_  = _w5553_ ;
	assign \g70567/_3_  = _w5581_ ;
	assign \g70568/_2_  = _w7257_ ;
	assign \g70571/_3_  = _w5510_ ;
	assign \g70577/_0_  = _w7269_ ;
	assign \g70578/_2_  = _w7270_ ;
	assign \g70585/_3_  = _w5598_ ;
	assign \g70586/_2_  = _w7271_ ;
	assign \g70587/_2_  = _w3180_ ;
	assign \g70588/_3_  = _w7272_ ;
	assign \g70602/_3_  = _w7273_ ;
	assign \g70841/_0_  = _w7279_ ;
	assign \g70842/_0_  = _w7285_ ;
	assign \g70843/_0_  = _w7291_ ;
	assign \g70844/_0_  = _w7297_ ;
	assign \g70845/_0_  = _w7303_ ;
	assign \g70846/_0_  = _w7309_ ;
	assign \g70847/_0_  = _w7315_ ;
	assign \g70848/_0_  = _w7321_ ;
	assign \g70849/_0_  = _w7327_ ;
	assign \g70850/_0_  = _w7333_ ;
	assign \g70851/_0_  = _w7339_ ;
	assign \g70852/_0_  = _w7345_ ;
	assign \g70853/_0_  = _w7351_ ;
	assign \g70854/_0_  = _w7357_ ;
	assign \g70855/_0_  = _w7363_ ;
	assign \g70856/_0_  = _w7369_ ;
	assign \g70857/_0_  = _w7375_ ;
	assign \g70858/_0_  = _w7381_ ;
	assign \g70859/_0_  = _w7387_ ;
	assign \g70860/_0_  = _w7393_ ;
	assign \g70861/_0_  = _w7399_ ;
	assign \g70862/_0_  = _w7405_ ;
	assign \g70863/_0_  = _w7411_ ;
	assign \g70864/_0_  = _w7417_ ;
	assign \g70865/_0_  = _w7423_ ;
	assign \g70866/_0_  = _w7429_ ;
	assign \g70867/_0_  = _w7435_ ;
	assign \g70868/_0_  = _w7441_ ;
	assign \g70869/_0_  = _w7447_ ;
	assign \g70870/_0_  = _w7453_ ;
	assign \g70871/_0_  = _w7459_ ;
	assign \g70872/_0_  = _w7465_ ;
	assign \g70944/_1__syn_2  = _w7469_ ;
	assign \g71042/_1__syn_2  = _w7472_ ;
	assign \g71064/_1__syn_2  = _w7475_ ;
	assign \g71065/_1__syn_2  = _w7477_ ;
	assign \g71076/_1__syn_2  = _w7479_ ;
	assign \g71077/_1__syn_2  = _w7481_ ;
	assign \g71202/_1__syn_2  = _w7483_ ;
	assign \g71204/_1__syn_2  = _w7485_ ;
	assign \g71236/_0_  = _w7486_ ;
	assign \g71237/_0_  = _w7487_ ;
	assign \g71241/_0_  = _w7488_ ;
	assign \g71242/_0_  = _w7489_ ;
	assign \g71245/_0_  = _w7490_ ;
	assign \g71246/_0_  = _w7491_ ;
	assign \g71306/_0_  = _w7492_ ;
	assign \g71308/_0_  = _w7493_ ;
	assign \g71309/_0_  = _w7494_ ;
	assign \g71310/_0_  = _w7495_ ;
	assign \g71355/_0_  = _w7496_ ;
	assign \g71416/_0_  = _w7497_ ;
	assign \g71417/_0_  = _w7498_ ;
	assign \g71420/_0_  = _w7499_ ;
	assign \g71432/_0_  = _w7500_ ;
	assign \g71434/_0_  = _w7501_ ;
	assign \g71435/_0_  = _w7502_ ;
	assign \g71436/_0_  = _w7503_ ;
	assign \g71446/_0_  = _w7504_ ;
	assign \g71449/_0_  = _w7505_ ;
	assign \g71451/_0_  = _w7506_ ;
	assign \g71452/_0_  = _w7507_ ;
	assign \g71485/_0_  = _w7508_ ;
	assign \g71494/_0_  = _w7509_ ;
	assign \g71499/_0_  = _w7510_ ;
	assign \g71500/_0_  = _w7511_ ;
	assign \g71501/_0_  = _w7512_ ;
	assign \g71502/_0_  = _w7513_ ;
	assign \g71503/_0_  = _w7514_ ;
	assign \g71504/_0_  = _w7515_ ;
	assign \g71505/_0_  = _w7516_ ;
	assign \g71506/_0_  = _w7517_ ;
	assign \g71815/_0_  = _w7518_ ;
	assign \g71823/_0_  = _w5868_ ;
	assign \g71832/_0_  = _w5407_ ;
	assign \g71833/_0__syn_2  = _w7519_ ;
	assign \g71837/_0_  = _w5271_ ;
	assign \g71838/_0_  = _w7520_ ;
	assign \g71846/_1__syn_2  = _w7521_ ;
	assign \g71847/_1__syn_2  = _w7522_ ;
	assign \g71849/_0_  = _w5418_ ;
	assign \g71854/_0_  = _w5288_ ;
	assign \g71858/_1__syn_2  = _w2240_ ;
	assign \g71859/_1__syn_2  = _w7523_ ;
	assign \g71863/_0_  = _w5308_ ;
	assign \g71867/_0_  = _w5424_ ;
	assign \g71869/_0_  = _w5428_ ;
	assign \g71872/_1_  = _w2271_ ;
	assign \g71873/_1__syn_2  = _w7524_ ;
	assign \g71874/_1__syn_2  = _w7526_ ;
	assign \g71875/_0_  = _w7527_ ;
	assign \g71877/_1__syn_2  = _w7529_ ;
	assign \g71881/_0_  = _w5884_ ;
	assign \g71906/_0_  = _w2273_ ;
	assign \g71907/_1__syn_2  = _w7530_ ;
	assign \g71910/_0_  = _w5280_ ;
	assign \g71911/_0_  = _w7531_ ;
	assign \g71912/_1__syn_2  = _w7533_ ;
	assign \g71913/_1__syn_2  = _w7535_ ;
	assign \g71914/_1__syn_2  = _w7536_ ;
	assign \g71918/_0_  = _w5445_ ;
	assign \g71921/_0_  = _w2245_ ;
	assign \g71922/_0_  = _w7537_ ;
	assign \g71929/_1__syn_2  = _w7538_ ;
	assign \g71931/_1__syn_2  = _w7539_ ;
	assign \g71938/_1__syn_2  = _w7540_ ;
	assign \g71942/_0_  = _w5328_ ;
	assign \g71946/_1__syn_2  = _w5265_ ;
	assign \g71947/_0_  = _w7541_ ;
	assign \g71951/_0_  = _w5745_ ;
	assign \g71958/_1__syn_2  = _w7542_ ;
	assign \g71965/_0_  = _w5330_ ;
	assign \g71970/_1__syn_2  = _w7543_ ;
	assign \g71972/_1__syn_2  = _w7544_ ;
	assign \g71973/_1__syn_2  = _w7545_ ;
	assign \g71986/_1__syn_2  = _w5259_ ;
	assign \g71987/_1__syn_2  = _w7546_ ;
	assign \g71990/_1__syn_2  = _w7548_ ;
	assign \g71991/_1__syn_2  = _w7549_ ;
	assign \g71992/_1__syn_2  = _w7550_ ;
	assign \g71994/_1__syn_2  = _w5459_ ;
	assign \g71997/_1__syn_2  = _w5348_ ;
	assign \g72001/_1__syn_2  = _w7551_ ;
	assign \g72013/_1__syn_2  = _w5352_ ;
	assign \g72021/_1__syn_2  = _w7552_ ;
	assign \g72030/_0_  = _w2252_ ;
	assign \g72031/_0__syn_2  = _w7553_ ;
	assign \g72036/_1__syn_2  = _w7554_ ;
	assign \g72038/_0_  = _w2269_ ;
	assign \g72042/_1__syn_2  = _w7555_ ;
	assign \g72047/_1__syn_2  = _w2277_ ;
	assign \g72048/_1__syn_2  = _w7556_ ;
	assign \g72049/_1__syn_2  = _w7557_ ;
	assign \g72056/_0_  = _w2275_ ;
	assign \g72064/_1__syn_2  = _w5837_ ;
	assign \g72073/_1__syn_2  = _w7558_ ;
	assign \g72075/_0_  = _w5401_ ;
	assign \g72078/_0_  = _w5404_ ;
	assign \g72081/_0_  = _w2279_ ;
	assign \g72091/_0_  = _w7559_ ;
	assign \g72096/_0_  = _w7560_ ;
	assign \g72100/_1__syn_2  = _w5664_ ;
	assign \g72113/_0_  = _w5299_ ;
	assign \g72118/_0_  = _w2259_ ;
	assign \g72121/_1__syn_2  = _w5232_ ;
	assign \g72122/_1__syn_2  = _w7561_ ;
	assign \g72125/_1__syn_2  = _w5338_ ;
	assign \g72128/_0_  = _w7562_ ;
	assign \g72140/_0_  = _w7563_ ;
	assign \g72144/_1__syn_2  = _w5690_ ;
	assign \g72154/_1__syn_2  = _w5379_ ;
	assign \g72159/_0_  = _w2263_ ;
	assign \g72164/_1__syn_2  = _w5242_ ;
	assign \g72165/_1__syn_2  = _w7564_ ;
	assign \g72167/_1__syn_2  = _w5318_ ;
	assign \g72170/_1__syn_2  = _w2250_ ;
	assign \g72172/_1__syn_2  = _w7565_ ;
	assign \g72173/_0_  = _w7566_ ;
	assign \g72177/_1__syn_2  = _w5718_ ;
	assign \g72189/_0_  = _w5320_ ;
	assign \g72194/_0_  = _w2265_ ;
	assign \g72196/_0_  = _w5316_ ;
	assign \g72198/_0_  = _w7567_ ;
	assign \g72206/_1__syn_2  = _w5390_ ;
	assign \g72209/_1__syn_2  = _w2255_ ;
	assign \g72210/_1__syn_2  = _w7568_ ;
	assign \g72211/_0_  = _w7569_ ;
	assign \g72215/_0_  = _w5786_ ;
	assign \g72227/_1__syn_2  = _w5341_ ;
	assign \g72229/_1__syn_2  = _w2267_ ;
	assign \g72230/_0_  = _w7570_ ;
	assign \g72239/_0_  = _w7573_ ;
	assign \g72250/_3_  = _w7574_ ;
	assign \g72251/_3_  = _w7575_ ;
	assign \g72252/_3_  = _w7576_ ;
	assign \g72253/_3_  = _w7577_ ;
	assign \g72254/_3_  = _w7578_ ;
	assign \g72255/_3_  = _w7579_ ;
	assign \g72256/_3_  = _w7580_ ;
	assign \g72257/_3_  = _w7581_ ;
	assign \g72259/_3_  = _w7582_ ;
	assign \g72260/_3_  = _w7583_ ;
	assign \g72261/_3_  = _w7584_ ;
	assign \g72262/_3_  = _w7585_ ;
	assign \g72263/_3_  = _w7586_ ;
	assign \g72264/_3_  = _w7587_ ;
	assign \g72265/_3_  = _w7588_ ;
	assign \g72266/_3_  = _w7589_ ;
	assign \g72267/_3_  = _w7590_ ;
	assign \g72273/_3_  = _w7591_ ;
	assign \g72275/_3_  = _w7592_ ;
	assign \g72282/_3_  = _w7593_ ;
	assign \g72285/_3_  = _w7594_ ;
	assign \g72293/_3_  = _w7595_ ;
	assign \g72304/_3_  = _w7596_ ;
	assign \g72305/_3_  = _w7597_ ;
	assign \g72306/_3_  = _w7598_ ;
	assign \g72307/_3_  = _w7599_ ;
	assign \g72309/_3_  = _w6128_ ;
	assign \g72310/_3_  = _w7600_ ;
	assign \g72324/_3_  = _w2998_ ;
	assign \g72325/_3_  = _w7601_ ;
	assign \g72326/_3_  = _w7602_ ;
	assign \g72327/_3_  = _w7603_ ;
	assign \g72711/_0_  = _w7616_ ;
	assign \g72763/_0_  = _w7619_ ;
	assign \g72966/_0_  = _w7623_ ;
	assign \g72967/_0_  = _w7625_ ;
	assign \g73018/_0_  = _w2510_ ;
	assign \g73058/_0_  = _w2519_ ;
	assign \g73062/_0_  = _w2515_ ;
	assign \g73067/_0_  = _w7628_ ;
	assign \g73068/_0_  = _w7629_ ;
	assign \g73207/_0_  = _w7263_ ;
	assign \g75007/_1__syn_2  = _w7630_ ;
	assign \g75568/_1_  = _w7606_ ;
	assign \g75792/_0_  = _w7631_ ;
	assign \g75836/_0_  = _w7632_ ;
	assign \g76027/_0_  = _w7633_ ;
	assign \g76034/_0_  = _w7634_ ;
	assign \g76108/_0_  = _w7635_ ;
	assign \g76130/_0_  = _w7636_ ;
	assign \g76266/_0_  = _w7637_ ;
	assign \g76315/_0_  = _w7638_ ;
	assign \g76569/_0_  = _w7639_ ;
	assign \g76714/_0_  = _w7640_ ;
	assign \g77122/_1__syn_2  = _w3386_ ;
	assign \g77709/_1_  = _w5972_ ;
	assign \g81909/_0_  = _w7641_ ;
	assign \g81922/_0_  = _w7642_ ;
	assign \g81926/_1__syn_2  = _w2257_ ;
	assign \g82197/_1_  = _w2435_ ;
	assign \g82272/_0_  = _w7643_ ;
	assign \g82291/_0_  = _w7644_ ;
	assign \g82716/_0_  = _w7645_ ;
	assign \g82718/_0_  = _w5449_ ;
	assign \g82738/_0_  = _w7646_ ;
	assign \g82769/_0_  = _w7647_ ;
	assign \g82775/_0_  = _w7648_ ;
	assign \g82779/_1__syn_2  = _w5254_ ;
	assign \g82804/_0_  = _w7649_ ;
	assign \g82810/_0_  = _w7650_ ;
	assign \g82817/_0_  = _w7651_ ;
	assign \g82823/_0_  = _w7652_ ;
	assign \g82835/_0_  = _w7653_ ;
	assign \g82841/_0_  = _w7654_ ;
	assign \g82847/_0_  = _w7655_ ;
	assign \g82853/_0_  = _w7656_ ;
	assign \g82859/_0_  = _w7657_ ;
	assign \g82862/_1__syn_2  = _w5249_ ;
	assign \g82956/_0_  = _w7658_ ;
	assign \g82959/_1_  = _w5430_ ;
	assign \g83020/_0_  = _w7659_ ;
	assign \g83025/_0_  = _w7660_ ;
	assign \g83078/_0_  = _w7661_ ;
	assign \g83083/_0_  = _w7662_ ;
	assign \g83121/_0_  = _w7663_ ;
	assign \g83135/_0_  = _w7664_ ;
	assign \g83205/_0_  = _w7665_ ;
	assign \g83240/_0_  = _w7666_ ;
	assign \g83509/_1__syn_2  = _w5573_ ;
	assign \g83769/_0_  = _w7667_ ;
	assign \h0lock_pad  = 1'b0;
	assign \h1sel_br[7]_pad  = _w5589_ ;
	assign \h1sel_dma[0]_pad  = _w5545_ ;
	assign \h1sel_dma[4]_pad  = _w5485_ ;
	assign \h1sel_dma[7]_pad  = _w5518_ ;
endmodule;