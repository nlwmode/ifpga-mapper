module top( \S1_reg[0]/NET0131  , \S1_reg[1]/NET0131  , \S1_reg[2]/NET0131  , \S2_reg[0]/NET0131  , \S2_reg[1]/NET0131  , \add_mpx2_pad  , \canale[0]_pad  , \canale[1]_pad  , \canale[2]_pad  , \confirm_reg/NET0131  , dsr_pad , eoc_pad , error_pad , \itfc_state_reg[0]/NET0131  , \itfc_state_reg[1]/NET0131  , load_dato_pad , \load_reg/NET0131  , \mpx_reg/NET0131  , \mux_en_reg/NET0131  , \next_bit_reg[0]/NET0131  , \next_bit_reg[1]/NET0131  , \next_bit_reg[2]/NET0131  , \next_bit_reg[3]/NET0131  , \out_reg_reg[0]/NET0131  , \out_reg_reg[1]/NET0131  , \out_reg_reg[2]/NET0131  , \out_reg_reg[3]/NET0131  , \out_reg_reg[4]/NET0131  , \out_reg_reg[5]/NET0131  , \out_reg_reg[6]/NET0131  , \out_reg_reg[7]/NET0131  , \rdy_reg/NET0131  , \send_data_reg/NET0131  , \send_en_reg/NET0131  , \send_reg/NET0131  , \shot_reg/NET0131  , \soc_reg/NET0131  , \tre_reg/NET0131  , \tx_conta_reg[0]/NET0131  , \tx_conta_reg[1]/NET0131  , \tx_conta_reg[2]/NET0131  , \tx_conta_reg[3]/NET0131  , \tx_conta_reg[4]/NET0131  , \tx_conta_reg[5]/NET0131  , \tx_conta_reg[6]/NET0131  , \tx_end_reg/NET0131  , \_al_n0  , \_al_n1  , \g1515/_0_  , \g1518/_0_  , \g1524/_0_  , \g1525/_0_  , \g1534/_0_  , \g1535/_0_  , \g1557/_0_  , \g1558/_0_  , \g1559/_0_  , \g1560/_0_  , \g1561/_0_  , \g1562/_0_  , \g1563/_0_  , \g1575/_0_  , \g1577/_0_  , \g1579/_0_  , \g1581/_0_  , \g1583/_3_  , \g1588/_1_  , \g1589/_0_  , \g1601/_0_  , \g1604/_0_  , \g1608/_0_  , \g1626/_0_  , \g1668/_0_  , \g1669/_0_  , \g1672/_0_  , \g1673/_0_  , \g1675/_3_  , \g1690/_0_  , \g1693/_0_  , \g1701/_0_  , \g1703/_0_  , \g1706/_3_  , \g1707/u3_syn_4  , \g1733/_0_  , \g1743/_0_  , \g1760/_0_  , \g2093/_0_  );
  input \S1_reg[0]/NET0131  ;
  input \S1_reg[1]/NET0131  ;
  input \S1_reg[2]/NET0131  ;
  input \S2_reg[0]/NET0131  ;
  input \S2_reg[1]/NET0131  ;
  input \add_mpx2_pad  ;
  input \canale[0]_pad  ;
  input \canale[1]_pad  ;
  input \canale[2]_pad  ;
  input \confirm_reg/NET0131  ;
  input dsr_pad ;
  input eoc_pad ;
  input error_pad ;
  input \itfc_state_reg[0]/NET0131  ;
  input \itfc_state_reg[1]/NET0131  ;
  input load_dato_pad ;
  input \load_reg/NET0131  ;
  input \mpx_reg/NET0131  ;
  input \mux_en_reg/NET0131  ;
  input \next_bit_reg[0]/NET0131  ;
  input \next_bit_reg[1]/NET0131  ;
  input \next_bit_reg[2]/NET0131  ;
  input \next_bit_reg[3]/NET0131  ;
  input \out_reg_reg[0]/NET0131  ;
  input \out_reg_reg[1]/NET0131  ;
  input \out_reg_reg[2]/NET0131  ;
  input \out_reg_reg[3]/NET0131  ;
  input \out_reg_reg[4]/NET0131  ;
  input \out_reg_reg[5]/NET0131  ;
  input \out_reg_reg[6]/NET0131  ;
  input \out_reg_reg[7]/NET0131  ;
  input \rdy_reg/NET0131  ;
  input \send_data_reg/NET0131  ;
  input \send_en_reg/NET0131  ;
  input \send_reg/NET0131  ;
  input \shot_reg/NET0131  ;
  input \soc_reg/NET0131  ;
  input \tre_reg/NET0131  ;
  input \tx_conta_reg[0]/NET0131  ;
  input \tx_conta_reg[1]/NET0131  ;
  input \tx_conta_reg[2]/NET0131  ;
  input \tx_conta_reg[3]/NET0131  ;
  input \tx_conta_reg[4]/NET0131  ;
  input \tx_conta_reg[5]/NET0131  ;
  input \tx_conta_reg[6]/NET0131  ;
  input \tx_end_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1515/_0_  ;
  output \g1518/_0_  ;
  output \g1524/_0_  ;
  output \g1525/_0_  ;
  output \g1534/_0_  ;
  output \g1535/_0_  ;
  output \g1557/_0_  ;
  output \g1558/_0_  ;
  output \g1559/_0_  ;
  output \g1560/_0_  ;
  output \g1561/_0_  ;
  output \g1562/_0_  ;
  output \g1563/_0_  ;
  output \g1575/_0_  ;
  output \g1577/_0_  ;
  output \g1579/_0_  ;
  output \g1581/_0_  ;
  output \g1583/_3_  ;
  output \g1588/_1_  ;
  output \g1589/_0_  ;
  output \g1601/_0_  ;
  output \g1604/_0_  ;
  output \g1608/_0_  ;
  output \g1626/_0_  ;
  output \g1668/_0_  ;
  output \g1669/_0_  ;
  output \g1672/_0_  ;
  output \g1673/_0_  ;
  output \g1675/_3_  ;
  output \g1690/_0_  ;
  output \g1693/_0_  ;
  output \g1701/_0_  ;
  output \g1703/_0_  ;
  output \g1706/_3_  ;
  output \g1707/u3_syn_4  ;
  output \g1733/_0_  ;
  output \g1743/_0_  ;
  output \g1760/_0_  ;
  output \g2093/_0_  ;
  wire n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
  assign n47 = ~\send_en_reg/NET0131  & \tx_conta_reg[4]/NET0131  ;
  assign n56 = \tx_conta_reg[0]/NET0131  & \tx_conta_reg[1]/NET0131  ;
  assign n57 = \tx_conta_reg[2]/NET0131  & n56 ;
  assign n58 = \tx_conta_reg[3]/NET0131  & n57 ;
  assign n59 = ~\tx_conta_reg[4]/NET0131  & ~n58 ;
  assign n48 = ~\tx_conta_reg[3]/NET0131  & ~\tx_conta_reg[4]/NET0131  ;
  assign n49 = \tx_conta_reg[5]/NET0131  & \tx_conta_reg[6]/NET0131  ;
  assign n50 = ~n48 & n49 ;
  assign n51 = ~\tx_conta_reg[0]/NET0131  & ~\tx_conta_reg[1]/NET0131  ;
  assign n52 = ~\tx_conta_reg[2]/NET0131  & ~\tx_conta_reg[4]/NET0131  ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & ~n53 ;
  assign n55 = \send_en_reg/NET0131  & ~n54 ;
  assign n60 = \tx_conta_reg[3]/NET0131  & \tx_conta_reg[4]/NET0131  ;
  assign n61 = n57 & n60 ;
  assign n62 = n55 & ~n61 ;
  assign n63 = ~n59 & n62 ;
  assign n64 = ~n47 & ~n63 ;
  assign n65 = ~\S1_reg[0]/NET0131  & \S1_reg[1]/NET0131  ;
  assign n66 = \S1_reg[2]/NET0131  & n65 ;
  assign n67 = ~\canale[0]_pad  & ~n66 ;
  assign n68 = \canale[0]_pad  & n66 ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = ~\canale[1]_pad  & ~n68 ;
  assign n71 = \canale[1]_pad  & n68 ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = \canale[2]_pad  & ~n71 ;
  assign n74 = ~\canale[2]_pad  & n71 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = \send_en_reg/NET0131  & n54 ;
  assign n77 = \next_bit_reg[0]/NET0131  & n76 ;
  assign n78 = \next_bit_reg[3]/NET0131  & ~n77 ;
  assign n79 = \next_bit_reg[0]/NET0131  & \next_bit_reg[1]/NET0131  ;
  assign n80 = \next_bit_reg[2]/NET0131  & n79 ;
  assign n81 = n76 & n80 ;
  assign n82 = ~n78 & ~n81 ;
  assign n83 = ~\send_en_reg/NET0131  & \tx_conta_reg[3]/NET0131  ;
  assign n84 = ~\tx_conta_reg[3]/NET0131  & ~n57 ;
  assign n85 = ~n58 & ~n84 ;
  assign n86 = n55 & n85 ;
  assign n87 = ~n83 & ~n86 ;
  assign n88 = ~\next_bit_reg[1]/NET0131  & ~\next_bit_reg[2]/NET0131  ;
  assign n89 = n76 & ~n88 ;
  assign n90 = ~\next_bit_reg[0]/NET0131  & ~n89 ;
  assign n91 = ~n77 & ~n90 ;
  assign n92 = \next_bit_reg[3]/NET0131  & n76 ;
  assign n93 = ~n91 & ~n92 ;
  assign n106 = \next_bit_reg[0]/NET0131  & ~\out_reg_reg[2]/NET0131  ;
  assign n105 = ~\next_bit_reg[0]/NET0131  & ~\out_reg_reg[3]/NET0131  ;
  assign n107 = \next_bit_reg[1]/NET0131  & ~n105 ;
  assign n108 = ~n106 & n107 ;
  assign n110 = \next_bit_reg[0]/NET0131  & ~\out_reg_reg[4]/NET0131  ;
  assign n109 = ~\next_bit_reg[0]/NET0131  & ~\out_reg_reg[5]/NET0131  ;
  assign n111 = ~\next_bit_reg[1]/NET0131  & ~n109 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ~n108 & ~n112 ;
  assign n114 = \next_bit_reg[2]/NET0131  & ~\next_bit_reg[3]/NET0131  ;
  assign n115 = ~n113 & n114 ;
  assign n101 = ~\out_reg_reg[6]/NET0131  & n79 ;
  assign n99 = \next_bit_reg[1]/NET0131  & \out_reg_reg[7]/NET0131  ;
  assign n100 = ~\next_bit_reg[0]/NET0131  & ~n99 ;
  assign n102 = ~\next_bit_reg[2]/NET0131  & ~\next_bit_reg[3]/NET0131  ;
  assign n103 = ~n100 & n102 ;
  assign n104 = ~n101 & n103 ;
  assign n94 = ~\next_bit_reg[0]/NET0131  & \out_reg_reg[1]/NET0131  ;
  assign n95 = \next_bit_reg[0]/NET0131  & \out_reg_reg[0]/NET0131  ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = \next_bit_reg[3]/NET0131  & n88 ;
  assign n98 = ~n96 & n97 ;
  assign n116 = n76 & ~n98 ;
  assign n117 = ~n104 & n116 ;
  assign n118 = ~n115 & n117 ;
  assign n119 = \next_bit_reg[1]/NET0131  & ~n77 ;
  assign n120 = \next_bit_reg[0]/NET0131  & ~\next_bit_reg[1]/NET0131  ;
  assign n121 = ~n102 & ~n120 ;
  assign n122 = \next_bit_reg[0]/NET0131  & ~\next_bit_reg[2]/NET0131  ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = n76 & n123 ;
  assign n125 = ~n119 & ~n124 ;
  assign n128 = \send_en_reg/NET0131  & n50 ;
  assign n126 = \send_en_reg/NET0131  & \tx_conta_reg[0]/NET0131  ;
  assign n127 = ~\tx_conta_reg[1]/NET0131  & ~n126 ;
  assign n129 = \tx_conta_reg[1]/NET0131  & n126 ;
  assign n130 = ~n127 & ~n129 ;
  assign n131 = ~n128 & n130 ;
  assign n132 = ~n50 & ~n57 ;
  assign n133 = \send_en_reg/NET0131  & ~n132 ;
  assign n134 = ~\tx_conta_reg[2]/NET0131  & ~n129 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = ~\send_en_reg/NET0131  & \tx_conta_reg[5]/NET0131  ;
  assign n138 = ~\tx_conta_reg[5]/NET0131  & ~n61 ;
  assign n137 = \tx_conta_reg[5]/NET0131  & n61 ;
  assign n139 = n55 & ~n137 ;
  assign n140 = ~n138 & n139 ;
  assign n141 = ~n136 & ~n140 ;
  assign n142 = \send_en_reg/NET0131  & n137 ;
  assign n144 = ~\tx_conta_reg[6]/NET0131  & ~n142 ;
  assign n143 = \tx_conta_reg[6]/NET0131  & n142 ;
  assign n145 = ~n76 & ~n143 ;
  assign n146 = ~n144 & n145 ;
  assign n147 = \S1_reg[0]/NET0131  & ~\S1_reg[1]/NET0131  ;
  assign n148 = \S1_reg[2]/NET0131  & n147 ;
  assign n149 = ~eoc_pad & n148 ;
  assign n150 = \S1_reg[0]/NET0131  & \S1_reg[1]/NET0131  ;
  assign n151 = \rdy_reg/NET0131  & n150 ;
  assign n152 = ~\S1_reg[0]/NET0131  & \S1_reg[2]/NET0131  ;
  assign n153 = \S1_reg[0]/NET0131  & ~\S1_reg[2]/NET0131  ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = ~n151 & ~n154 ;
  assign n156 = ~n149 & ~n155 ;
  assign n157 = ~\S2_reg[0]/NET0131  & ~\S2_reg[1]/NET0131  ;
  assign n158 = \send_data_reg/NET0131  & n157 ;
  assign n159 = ~\S2_reg[0]/NET0131  & \S2_reg[1]/NET0131  ;
  assign n160 = \confirm_reg/NET0131  & n159 ;
  assign n161 = \mpx_reg/NET0131  & n160 ;
  assign n162 = \rdy_reg/NET0131  & ~n161 ;
  assign n163 = ~n158 & ~n162 ;
  assign n164 = ~\S1_reg[0]/NET0131  & ~\S1_reg[1]/NET0131  ;
  assign n165 = ~\S1_reg[2]/NET0131  & n164 ;
  assign n166 = ~\mux_en_reg/NET0131  & ~n165 ;
  assign n167 = ~n149 & ~n166 ;
  assign n168 = ~\tx_conta_reg[0]/NET0131  & ~n55 ;
  assign n169 = ~n126 & ~n168 ;
  assign n170 = n102 & n120 ;
  assign n171 = n76 & n170 ;
  assign n172 = ~\soc_reg/NET0131  & ~n65 ;
  assign n173 = ~n66 & ~n172 ;
  assign n174 = load_dato_pad & ~n66 ;
  assign n175 = ~n149 & ~n174 ;
  assign n176 = ~n153 & ~n164 ;
  assign n177 = \S1_reg[2]/NET0131  & n150 ;
  assign n178 = \send_data_reg/NET0131  & ~n151 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = \confirm_reg/NET0131  & ~\mpx_reg/NET0131  ;
  assign n181 = n159 & n180 ;
  assign n182 = ~\add_mpx2_pad  & ~n181 ;
  assign n183 = ~\confirm_reg/NET0131  & n159 ;
  assign n184 = \S2_reg[0]/NET0131  & ~\S2_reg[1]/NET0131  ;
  assign n185 = ~\shot_reg/NET0131  & ~n184 ;
  assign n186 = ~n183 & ~n185 ;
  assign n187 = \itfc_state_reg[0]/NET0131  & ~\itfc_state_reg[1]/NET0131  ;
  assign n188 = \load_reg/NET0131  & ~n187 ;
  assign n189 = ~\itfc_state_reg[0]/NET0131  & ~\itfc_state_reg[1]/NET0131  ;
  assign n190 = \shot_reg/NET0131  & n189 ;
  assign n191 = ~n188 & ~n190 ;
  assign n192 = ~\mpx_reg/NET0131  & ~n160 ;
  assign n193 = ~n161 & ~n192 ;
  assign n194 = n159 & ~n180 ;
  assign n195 = ~n184 & ~n194 ;
  assign n196 = \itfc_state_reg[0]/NET0131  & \itfc_state_reg[1]/NET0131  ;
  assign n197 = \tx_end_reg/NET0131  & n196 ;
  assign n198 = \confirm_reg/NET0131  & ~n189 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = ~\next_bit_reg[2]/NET0131  & ~n79 ;
  assign n201 = ~n80 & ~n200 ;
  assign n202 = n189 & ~n196 ;
  assign n203 = ~n197 & ~n202 ;
  assign n204 = ~\itfc_state_reg[0]/NET0131  & \itfc_state_reg[1]/NET0131  ;
  assign n205 = \send_reg/NET0131  & ~n204 ;
  assign n206 = ~n187 & ~n205 ;
  assign n207 = ~\tx_end_reg/NET0131  & n196 ;
  assign n208 = ~n190 & ~n204 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = dsr_pad & \send_reg/NET0131  ;
  assign n211 = \tre_reg/NET0131  & n210 ;
  assign n212 = \load_reg/NET0131  & ~\tre_reg/NET0131  ;
  assign n213 = ~error_pad & ~\load_reg/NET0131  ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = ~\send_reg/NET0131  & ~n214 ;
  assign n216 = ~n211 & ~n215 ;
  assign n217 = ~n158 & ~n160 ;
  assign n218 = \send_en_reg/NET0131  & ~\tx_end_reg/NET0131  ;
  assign n219 = ~n211 & ~n218 ;
  assign n220 = ~\load_reg/NET0131  & ~\tre_reg/NET0131  ;
  assign n221 = ~\tx_end_reg/NET0131  & n220 ;
  assign n224 = eoc_pad & n148 ;
  assign n222 = \S1_reg[1]/NET0131  & ~\S1_reg[2]/NET0131  ;
  assign n223 = ~\rdy_reg/NET0131  & n222 ;
  assign n225 = \S1_reg[0]/NET0131  & ~n223 ;
  assign n226 = ~n224 & n225 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1515/_0_  = ~n64 ;
  assign \g1518/_0_  = n69 ;
  assign \g1524/_0_  = n72 ;
  assign \g1525/_0_  = ~n75 ;
  assign \g1534/_0_  = ~n82 ;
  assign \g1535/_0_  = ~n87 ;
  assign \g1557/_0_  = ~n93 ;
  assign \g1558/_0_  = ~n118 ;
  assign \g1559/_0_  = ~n125 ;
  assign \g1560/_0_  = n131 ;
  assign \g1561/_0_  = n135 ;
  assign \g1562/_0_  = ~n141 ;
  assign \g1563/_0_  = n146 ;
  assign \g1575/_0_  = ~n156 ;
  assign \g1577/_0_  = ~n163 ;
  assign \g1579/_0_  = n167 ;
  assign \g1581/_0_  = n169 ;
  assign \g1583/_3_  = n171 ;
  assign \g1588/_1_  = n76 ;
  assign \g1589/_0_  = n173 ;
  assign \g1601/_0_  = ~n175 ;
  assign \g1604/_0_  = n176 ;
  assign \g1608/_0_  = ~n179 ;
  assign \g1626/_0_  = ~n182 ;
  assign \g1668/_0_  = n186 ;
  assign \g1669/_0_  = ~n191 ;
  assign \g1672/_0_  = n193 ;
  assign \g1673/_0_  = ~n195 ;
  assign \g1675/_3_  = ~n199 ;
  assign \g1690/_0_  = n201 ;
  assign \g1693/_0_  = n203 ;
  assign \g1701/_0_  = ~n206 ;
  assign \g1703/_0_  = ~n209 ;
  assign \g1706/_3_  = n216 ;
  assign \g1707/u3_syn_4  = n212 ;
  assign \g1733/_0_  = ~n217 ;
  assign \g1743/_0_  = ~n219 ;
  assign \g1760/_0_  = ~n221 ;
  assign \g2093/_0_  = ~n226 ;
endmodule
