module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , a_pad, \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , d_pad, \e0_pad , \e1_pad , \e2_pad , \e3_pad , \e4_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , \i3_pad , \i4_pad , i_pad, \j0_pad , \j1_pad , \j2_pad , \j3_pad , \j4_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , \l4_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , \m6_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , \n4_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , o_pad, \p0_pad , \p1_pad , \p2_pad , \p3_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , \q3_pad , q_pad, \r1_pad , \r2_pad , \r3_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , \t4_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u4_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , x_pad, \y0_pad , \y1_pad , \y2_pad , \y3_pad , y_pad, \z0_pad , \z1_pad , \z2_pad , \z3_pad , z_pad, \a5_pad , \a6_pad , \a7_pad , \a8_pad , \a9_pad , \b5_pad , \b6_pad , \b7_pad , \b8_pad , \b9_pad , \c5_pad , \c6_pad , \c7_pad , \c8_pad , \c9_pad , \d5_pad , \d6_pad , \d7_pad , \d8_pad , \d9_pad , \e5_pad , \e6_pad , \e7_pad , \e8_pad , \e9_pad , \f5_pad , \f6_pad , \f7_pad , \f8_pad , \f9_pad , \g5_pad , \g6_pad , \g7_pad , \g8_pad , \g9_pad , \h5_pad , \h6_pad , \h7_pad , \h8_pad , \h9_pad , \i5_pad , \i6_pad , \i7_pad , \i8_pad , \i9_pad , \j5_pad , \j6_pad , \j7_pad , \j8_pad , \j9_pad , \k5_pad , \k6_pad , \k7_pad , \k8_pad , \k9_pad , \l5_pad , \l6_pad , \l7_pad , \l8_pad , \l9_pad , \m7_pad , \m8_pad , \m9_pad , \n5_pad , \n6_pad , \n7_pad , \n8_pad , \n9_pad , \o4_pad , \o5_pad , \o6_pad , \o7_pad , \o8_pad , \o9_pad , \p4_pad , \p5_pad , \p6_pad , \p7_pad , \p8_pad , \p9_pad , \q4_pad , \q5_pad , \q6_pad , \q7_pad , \q8_pad , \q9_pad , \r4_pad , \r5_pad , \r6_pad , \r7_pad , \r8_pad , \r9_pad , \s4_pad , \s6_pad , \s7_pad , \s8_pad , \s9_pad , \t6_pad , \t7_pad , \t8_pad , \t9_pad , \u6_pad , \u7_pad , \u8_pad , \u9_pad , \v4_pad , \v6_pad , \v7_pad , \v8_pad , \v9_pad , \w4_pad , \w5_pad , \w6_pad , \w7_pad , \w8_pad , \w9_pad , \x4_pad , \x5_pad , \x6_pad , \x7_pad , \x8_pad , \y4_pad , \y5_pad , \y6_pad , \y7_pad , \y8_pad , \z4_pad , \z5_pad , \z6_pad , \z7_pad , \z8_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input \i4_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input \j4_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input \l4_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input \m6_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input \n4_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input q_pad ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input \t4_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u4_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input z_pad ;
	output \a5_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \a9_pad  ;
	output \b5_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \b9_pad  ;
	output \c5_pad  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \c9_pad  ;
	output \d5_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \d8_pad  ;
	output \d9_pad  ;
	output \e5_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \e8_pad  ;
	output \e9_pad  ;
	output \f5_pad  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \f8_pad  ;
	output \f9_pad  ;
	output \g5_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \g8_pad  ;
	output \g9_pad  ;
	output \h5_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \h8_pad  ;
	output \h9_pad  ;
	output \i5_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \i8_pad  ;
	output \i9_pad  ;
	output \j5_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \j8_pad  ;
	output \j9_pad  ;
	output \k5_pad  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \k8_pad  ;
	output \k9_pad  ;
	output \l5_pad  ;
	output \l6_pad  ;
	output \l7_pad  ;
	output \l8_pad  ;
	output \l9_pad  ;
	output \m7_pad  ;
	output \m8_pad  ;
	output \m9_pad  ;
	output \n5_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \n8_pad  ;
	output \n9_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \o8_pad  ;
	output \o9_pad  ;
	output \p4_pad  ;
	output \p5_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \p8_pad  ;
	output \p9_pad  ;
	output \q4_pad  ;
	output \q5_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \q8_pad  ;
	output \q9_pad  ;
	output \r4_pad  ;
	output \r5_pad  ;
	output \r6_pad  ;
	output \r7_pad  ;
	output \r8_pad  ;
	output \r9_pad  ;
	output \s4_pad  ;
	output \s6_pad  ;
	output \s7_pad  ;
	output \s8_pad  ;
	output \s9_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \t8_pad  ;
	output \t9_pad  ;
	output \u6_pad  ;
	output \u7_pad  ;
	output \u8_pad  ;
	output \u9_pad  ;
	output \v4_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \v8_pad  ;
	output \v9_pad  ;
	output \w4_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \w8_pad  ;
	output \w9_pad  ;
	output \x4_pad  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \x8_pad  ;
	output \y4_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \y8_pad  ;
	output \z4_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	output \z8_pad  ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\k0_pad ,
		\l0_pad ,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\k0_pad ,
		\l0_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\r3_pad ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\j3_pad ,
		_w145_,
		_w147_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\m0_pad ,
		_w146_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\m1_pad ,
		\m6_pad ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\k1_pad ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\o0_pad ,
		\q0_pad ,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\k1_pad ,
		\l1_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\j1_pad ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\h1_pad ,
		\i1_pad ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\n0_pad ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\f0_pad ,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\y3_pad ,
		\z3_pad ,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\a4_pad ,
		\b4_pad ,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\c4_pad ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w159_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\x3_pad ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\l4_pad ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\r1_pad ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\s1_pad ,
		_w164_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w157_,
		_w165_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w158_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w152_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\m0_pad ,
		_w157_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		h_pad,
		_w143_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		p_pad,
		_w143_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w171_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\r2_pad ,
		_w164_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\s2_pad ,
		_w164_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w171_,
		_w176_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w175_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		_w152_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\k1_pad ,
		\l1_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\j1_pad ,
		_w153_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w155_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w154_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\e4_pad ,
		\f4_pad ,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\g4_pad ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		\h4_pad ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\h1_pad ,
		\x0_pad ,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\j1_pad ,
		\z0_pad ,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		\b1_pad ,
		\l1_pad ,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\i1_pad ,
		\y0_pad ,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\a1_pad ,
		\k1_pad ,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w190_,
		_w191_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w192_,
		_w193_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w194_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w195_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w189_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\m6_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\h1_pad ,
		\i1_pad ,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w156_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w186_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w200_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\r3_pad ,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\s3_pad ,
		_w204_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w152_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\s3_pad ,
		_w145_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\k3_pad ,
		_w145_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\m0_pad ,
		_w209_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\l1_pad ,
		_w150_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\e0_pad ,
		_w157_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\s1_pad ,
		_w164_,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\t1_pad ,
		_w164_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w157_,
		_w215_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w214_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w152_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w145_,
		_w171_,
		_w221_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		i_pad,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\s2_pad ,
		_w164_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		\t2_pad ,
		_w164_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w221_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		_w152_,
		_w222_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\s3_pad ,
		_w204_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		\t3_pad ,
		_w204_,
		_w230_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w152_,
		_w229_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\t3_pad ,
		_w145_,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		\l3_pad ,
		_w145_,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\m0_pad ,
		_w233_,
		_w235_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\h1_pad ,
		\l4_pad ,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\d0_pad ,
		_w157_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\t1_pad ,
		_w164_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\u1_pad ,
		_w164_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w157_,
		_w239_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w238_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		_w152_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		j_pad,
		_w221_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\t2_pad ,
		_w164_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\u2_pad ,
		_w164_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w246_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w221_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		_w152_,
		_w245_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\t3_pad ,
		_w204_,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\t4_pad ,
		_w204_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		_w152_,
		_w252_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\m0_pad ,
		\m3_pad ,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\i1_pad ,
		\l4_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w152_,
		_w171_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\u1_pad ,
		_w164_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\v1_pad ,
		_w164_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w157_,
		_w259_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w258_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		k_pad,
		_w221_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\u2_pad ,
		_w164_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\v2_pad ,
		_w164_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w265_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w221_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		_w152_,
		_w264_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		\t4_pad ,
		_w204_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		\u4_pad ,
		_w204_,
		_w272_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		_w152_,
		_w271_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\m0_pad ,
		\n3_pad ,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\j1_pad ,
		\l4_pad ,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\k0_pad ,
		_w157_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		\v1_pad ,
		_w164_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		\w1_pad ,
		_w164_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w157_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		_w152_,
		_w277_,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		l_pad,
		_w221_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\v2_pad ,
		_w164_,
		_w285_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\w2_pad ,
		_w164_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w221_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		_w152_,
		_w284_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\u4_pad ,
		_w204_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		\w3_pad ,
		_w204_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w152_,
		_w291_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w292_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\m0_pad ,
		\o3_pad ,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\k1_pad ,
		\l4_pad ,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		\l0_pad ,
		_w157_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\w1_pad ,
		_w164_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\x1_pad ,
		_w164_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w157_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		_w152_,
		_w297_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		m_pad,
		_w221_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\w2_pad ,
		_w164_,
		_w305_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\x2_pad ,
		_w164_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w221_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		_w152_,
		_w304_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\w3_pad ,
		_w204_,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		\h1_pad ,
		\i1_pad ,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\s0_pad ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w154_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\j1_pad ,
		\l1_pad ,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\k1_pad ,
		\v0_pad ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\l1_pad ,
		\u0_pad ,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		\j1_pad ,
		\w0_pad ,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\k1_pad ,
		_w315_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\i1_pad ,
		_w317_,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\t0_pad ,
		_w154_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		\i1_pad ,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\h1_pad ,
		_w324_,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w314_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		_w200_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w311_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		_w152_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\m0_pad ,
		\p3_pad ,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\l1_pad ,
		\l4_pad ,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		q_pad,
		_w157_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		\x1_pad ,
		_w164_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		\y1_pad ,
		_w164_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w157_,
		_w336_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w335_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		_w152_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		n_pad,
		_w221_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		\x2_pad ,
		_w164_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\y2_pad ,
		_w164_,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w221_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		_w152_,
		_w342_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		_w152_,
		_w157_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		\l4_pad ,
		\x3_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\l4_pad ,
		\x3_pad ,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w162_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w350_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w349_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\m0_pad ,
		\q3_pad ,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		r_pad,
		_w157_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\y1_pad ,
		_w164_,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\z1_pad ,
		_w164_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w157_,
		_w357_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w356_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w152_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		o_pad,
		_w221_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		\y2_pad ,
		_w164_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		\z2_pad ,
		_w164_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w221_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w152_,
		_w363_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\y3_pad ,
		_w352_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\y3_pad ,
		_w351_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w370_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		_w349_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\m0_pad ,
		\r3_pad ,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		s_pad,
		_w157_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\z1_pad ,
		_w164_,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\a2_pad ,
		_w164_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w157_,
		_w376_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w375_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		_w152_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		p_pad,
		_w221_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\z2_pad ,
		_w164_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w221_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w382_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		_w152_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\z3_pad ,
		_w370_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w159_,
		_w351_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w161_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w387_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		_w349_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\m0_pad ,
		\s3_pad ,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		t_pad,
		_w157_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\a2_pad ,
		_w164_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\b2_pad ,
		_w164_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w157_,
		_w394_,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w393_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w152_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\a3_pad ,
		_w204_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		\b3_pad ,
		_w204_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		_w152_,
		_w400_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		\a4_pad ,
		_w389_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		\a4_pad ,
		_w388_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w157_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w404_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w145_,
		_w171_,
		_w408_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		_w152_,
		_w407_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w408_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\m0_pad ,
		\t3_pad ,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		u_pad,
		_w157_,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		\b2_pad ,
		_w164_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name271 (
		\c2_pad ,
		_w164_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w157_,
		_w413_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w414_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w412_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w152_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		\b3_pad ,
		_w204_,
		_w419_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		\c3_pad ,
		_w204_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		_w152_,
		_w419_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w420_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\b4_pad ,
		_w404_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w160_,
		_w389_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w157_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w423_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w258_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\g1_pad ,
		\j4_pad ,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		v_pad,
		_w157_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		\c2_pad ,
		_w164_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		\d2_pad ,
		_w164_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w157_,
		_w430_,
		_w432_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w431_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w429_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w152_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\c3_pad ,
		_w204_,
		_w436_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\d3_pad ,
		_w204_,
		_w437_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w152_,
		_w436_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\c4_pad ,
		_w425_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w171_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w152_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		w_pad,
		_w157_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		\d2_pad ,
		_w164_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\e2_pad ,
		_w164_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w157_,
		_w444_,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w443_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w152_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\d3_pad ,
		_w204_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		\e3_pad ,
		_w204_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w152_,
		_w450_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\q0_pad ,
		_w157_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\g1_pad ,
		\q0_pad ,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		\d4_pad ,
		_w200_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		\d4_pad ,
		_w200_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w455_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w454_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		\o0_pad ,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\h1_pad ,
		\m6_pad ,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		\n0_pad ,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\f1_pad ,
		\i4_pad ,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\f1_pad ,
		\i4_pad ,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w464_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		x_pad,
		_w157_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		\e2_pad ,
		_w164_,
		_w468_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		\f2_pad ,
		_w164_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w157_,
		_w468_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w469_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w467_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		_w152_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		\e3_pad ,
		_w204_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		\f3_pad ,
		_w204_,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		_w152_,
		_w474_,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\e4_pad ,
		_w457_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\d4_pad ,
		_w157_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w200_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		\e4_pad ,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w478_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\o0_pad ,
		_w455_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w157_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w482_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\i1_pad ,
		\m6_pad ,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		\n0_pad ,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\x3_pad ,
		_w162_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		y_pad,
		_w157_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\f2_pad ,
		_w164_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		\g2_pad ,
		_w164_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w157_,
		_w490_,
		_w492_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w489_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w152_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\f3_pad ,
		_w204_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\g3_pad ,
		_w204_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		_w152_,
		_w496_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		\e4_pad ,
		\f4_pad ,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w480_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\f4_pad ,
		_w478_,
		_w502_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		_w484_,
		_w501_,
		_w503_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		\l3_pad ,
		_w145_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\d3_pad ,
		_w145_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w505_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		\m0_pad ,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		\m0_pad ,
		\t3_pad ,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w508_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		\j1_pad ,
		\m6_pad ,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		\n0_pad ,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\n4_pad ,
		_w189_,
		_w513_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w198_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\d4_pad ,
		\g1_pad ,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w189_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w514_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w152_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		z_pad,
		_w157_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\g2_pad ,
		_w164_,
		_w520_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		\h2_pad ,
		_w164_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w157_,
		_w520_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w521_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w519_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		_w152_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\g3_pad ,
		_w204_,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		\h3_pad ,
		_w204_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		_w152_,
		_w526_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w527_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\m0_pad ,
		_w145_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		_w152_,
		_w157_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		\g1_pad ,
		\m6_pad ,
		_w533_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\d4_pad ,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		_w188_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w199_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		_w349_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w187_,
		_w480_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\g4_pad ,
		_w484_,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w532_,
		_w537_,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		\k3_pad ,
		_w145_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		\c3_pad ,
		_w145_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\m0_pad ,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		\m0_pad ,
		\s3_pad ,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\k1_pad ,
		\m6_pad ,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		\n0_pad ,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		\h1_pad ,
		_w483_,
		_w551_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		\e1_pad ,
		_w157_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\c1_pad ,
		\d1_pad ,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w152_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w552_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w551_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\a0_pad ,
		_w157_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		\h2_pad ,
		_w164_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		\i2_pad ,
		_w164_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w157_,
		_w558_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w557_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h2)
	) name420 (
		_w152_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		\h3_pad ,
		_w204_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		\i3_pad ,
		_w204_,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		_w152_,
		_w564_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		\m0_pad ,
		_w531_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		\g4_pad ,
		_w538_,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\h4_pad ,
		_w484_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w568_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		\j3_pad ,
		_w145_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		\b3_pad ,
		_w145_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w573_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\m0_pad ,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\m0_pad ,
		\r3_pad ,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w576_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\l1_pad ,
		\m6_pad ,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		\n0_pad ,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		\e1_pad ,
		_w553_,
		_w581_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		_w157_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		\g1_pad ,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		\i1_pad ,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		\c1_pad ,
		\d1_pad ,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w552_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w584_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		_w152_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		\b0_pad ,
		_w157_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\i2_pad ,
		_w164_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		\j2_pad ,
		_w164_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w157_,
		_w590_,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name450 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w589_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h2)
	) name452 (
		_w152_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		\i3_pad ,
		_w204_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\j3_pad ,
		_w204_,
		_w597_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		_w152_,
		_w596_,
		_w598_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w597_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		\i4_pad ,
		\n1_pad ,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		\i4_pad ,
		\n1_pad ,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w600_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		_w152_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w164_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		\i3_pad ,
		_w145_,
		_w605_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		\a3_pad ,
		_w145_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		\m0_pad ,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		\m0_pad ,
		\q3_pad ,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w608_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		\j1_pad ,
		_w583_,
		_w611_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		\c1_pad ,
		\d1_pad ,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w552_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		_w611_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h2)
	) name472 (
		_w152_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		\c0_pad ,
		_w157_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		\j2_pad ,
		_w164_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name475 (
		\k2_pad ,
		_w164_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w157_,
		_w617_,
		_w619_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w616_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		_w152_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\j3_pad ,
		_w204_,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		\k3_pad ,
		_w204_,
		_w624_
	);
	LUT2 #(
		.INIT('h2)
	) name482 (
		_w152_,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		\k1_pad ,
		\w0_pad ,
		_w627_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		\l1_pad ,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		\i1_pad ,
		\j1_pad ,
		_w629_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		_w316_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w628_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\h1_pad ,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w314_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		\u0_pad ,
		_w153_,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		_w155_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		\m6_pad ,
		\n4_pad ,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w184_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w635_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		_w326_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		_w199_,
		_w633_,
		_w640_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		\j4_pad ,
		_w483_,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		\j4_pad ,
		\n4_pad ,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name502 (
		_w152_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		_w533_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w199_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w329_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w643_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		\k1_pad ,
		_w552_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name508 (
		_w583_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		\c1_pad ,
		\d1_pad ,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w552_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w651_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		_w152_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		a_pad,
		_w143_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		i_pad,
		_w143_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w656_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		_w171_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		\k2_pad ,
		_w164_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		\l2_pad ,
		_w164_,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w171_,
		_w660_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w661_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w659_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		_w152_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		\k3_pad ,
		_w204_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		\l3_pad ,
		_w204_,
		_w667_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w152_,
		_w666_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		\m1_pad ,
		_w152_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w162_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		_w157_,
		_w553_,
		_w672_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		\g1_pad ,
		\l1_pad ,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w672_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		_w152_,
		_w552_,
		_w675_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		b_pad,
		_w143_,
		_w677_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		j_pad,
		_w143_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w677_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w171_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		\l2_pad ,
		_w164_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		\m2_pad ,
		_w164_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w171_,
		_w681_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w680_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w152_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		\l3_pad ,
		_w204_,
		_w687_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\m3_pad ,
		_w204_,
		_w688_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		_w152_,
		_w687_,
		_w689_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w688_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w163_,
		_w670_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\m3_pad ,
		_w145_,
		_w692_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\e3_pad ,
		_w145_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		\m0_pad ,
		_w692_,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		\n0_pad ,
		\p0_pad ,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		\m1_pad ,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		\m1_pad ,
		_w517_,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		_w152_,
		_w697_,
		_w699_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		c_pad,
		_w143_,
		_w701_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		k_pad,
		_w143_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w701_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		_w171_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		\m2_pad ,
		_w164_,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		\n2_pad ,
		_w164_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w171_,
		_w705_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w704_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		_w152_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\m3_pad ,
		_w204_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		\n3_pad ,
		_w204_,
		_w712_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		_w152_,
		_w711_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w198_,
		_w513_,
		_w715_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		_w518_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\n3_pad ,
		_w145_,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		\f3_pad ,
		_w145_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		\m0_pad ,
		_w717_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		_w162_,
		_w466_,
		_w721_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		\n1_pad ,
		_w162_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w721_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		\j0_pad ,
		_w157_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		\n1_pad ,
		_w164_,
		_w725_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		\o1_pad ,
		_w164_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w157_,
		_w725_,
		_w727_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w726_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w724_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w152_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		d_pad,
		_w143_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		l_pad,
		_w143_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w171_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		\n2_pad ,
		_w164_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		\o2_pad ,
		_w164_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w171_,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w734_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h2)
	) name597 (
		_w152_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		\n3_pad ,
		_w204_,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name599 (
		\o3_pad ,
		_w204_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		_w152_,
		_w741_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\m6_pad ,
		_w152_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w198_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		\o3_pad ,
		_w145_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		\g3_pad ,
		_w145_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\m0_pad ,
		_w747_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\h1_pad ,
		_w150_,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\i0_pad ,
		_w157_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		\o1_pad ,
		_w164_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		\p1_pad ,
		_w164_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		_w157_,
		_w753_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		_w754_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w752_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name615 (
		_w152_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		e_pad,
		_w143_,
		_w759_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		m_pad,
		_w143_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w759_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		_w171_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\o2_pad ,
		_w164_,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		\p2_pad ,
		_w164_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		_w171_,
		_w763_,
		_w765_
	);
	LUT2 #(
		.INIT('h4)
	) name623 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w762_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		_w152_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		\o3_pad ,
		_w204_,
		_w769_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		\p3_pad ,
		_w204_,
		_w770_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		_w152_,
		_w769_,
		_w771_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w770_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		\p3_pad ,
		_w145_,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		\h3_pad ,
		_w145_,
		_w774_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\m0_pad ,
		_w773_,
		_w775_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w774_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\i1_pad ,
		_w150_,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\h0_pad ,
		_w157_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\p1_pad ,
		_w164_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		\q1_pad ,
		_w164_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w157_,
		_w779_,
		_w781_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w780_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w778_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w152_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		f_pad,
		_w143_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		n_pad,
		_w143_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w171_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		\p2_pad ,
		_w164_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		\q2_pad ,
		_w164_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w171_,
		_w789_,
		_w791_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w790_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w788_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		_w152_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		\p3_pad ,
		_w204_,
		_w795_
	);
	LUT2 #(
		.INIT('h4)
	) name653 (
		\q3_pad ,
		_w204_,
		_w796_
	);
	LUT2 #(
		.INIT('h2)
	) name654 (
		_w152_,
		_w795_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		_w796_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		\q3_pad ,
		_w145_,
		_w799_
	);
	LUT2 #(
		.INIT('h4)
	) name657 (
		\i3_pad ,
		_w145_,
		_w800_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		\m0_pad ,
		_w799_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		_w800_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		\j1_pad ,
		_w150_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		\g0_pad ,
		_w157_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		\q1_pad ,
		_w164_,
		_w805_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		\r1_pad ,
		_w164_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w157_,
		_w805_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		_w806_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w804_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		_w152_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		g_pad,
		_w143_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		o_pad,
		_w143_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w171_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		\q2_pad ,
		_w164_,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		\r2_pad ,
		_w164_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w171_,
		_w815_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w816_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w814_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		_w152_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		\q3_pad ,
		_w204_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		\r3_pad ,
		_w204_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		_w152_,
		_w821_,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w822_,
		_w823_,
		_w824_
	);
	assign \a5_pad  = _w149_ ;
	assign \a6_pad  = _w151_ ;
	assign \a7_pad  = _w170_ ;
	assign \a8_pad  = _w181_ ;
	assign \a9_pad  = _w208_ ;
	assign \b5_pad  = _w212_ ;
	assign \b6_pad  = _w213_ ;
	assign \b7_pad  = _w220_ ;
	assign \b8_pad  = _w228_ ;
	assign \b9_pad  = _w232_ ;
	assign \c5_pad  = _w236_ ;
	assign \c6_pad  = _w237_ ;
	assign \c7_pad  = _w244_ ;
	assign \c8_pad  = _w251_ ;
	assign \c9_pad  = _w255_ ;
	assign \d5_pad  = _w256_ ;
	assign \d6_pad  = _w257_ ;
	assign \d7_pad  = _w263_ ;
	assign \d8_pad  = _w270_ ;
	assign \d9_pad  = _w274_ ;
	assign \e5_pad  = _w275_ ;
	assign \e6_pad  = _w276_ ;
	assign \e7_pad  = _w283_ ;
	assign \e8_pad  = _w290_ ;
	assign \e9_pad  = _w294_ ;
	assign \f5_pad  = _w295_ ;
	assign \f6_pad  = _w296_ ;
	assign \f7_pad  = _w303_ ;
	assign \f8_pad  = _w310_ ;
	assign \f9_pad  = _w332_ ;
	assign \g5_pad  = _w333_ ;
	assign \g6_pad  = _w334_ ;
	assign \g7_pad  = _w341_ ;
	assign \g8_pad  = _w348_ ;
	assign \g9_pad  = _w354_ ;
	assign \h5_pad  = _w355_ ;
	assign \h6_pad  = \h1_pad ;
	assign \h7_pad  = _w362_ ;
	assign \h8_pad  = _w369_ ;
	assign \h9_pad  = _w373_ ;
	assign \i5_pad  = _w374_ ;
	assign \i6_pad  = \i1_pad ;
	assign \i7_pad  = _w381_ ;
	assign \i8_pad  = _w386_ ;
	assign \i9_pad  = _w391_ ;
	assign \j5_pad  = _w392_ ;
	assign \j6_pad  = \j1_pad ;
	assign \j7_pad  = _w399_ ;
	assign \j8_pad  = _w403_ ;
	assign \j9_pad  = _w410_ ;
	assign \k5_pad  = _w411_ ;
	assign \k6_pad  = \k1_pad ;
	assign \k7_pad  = _w418_ ;
	assign \k8_pad  = _w422_ ;
	assign \k9_pad  = _w427_ ;
	assign \l5_pad  = _w428_ ;
	assign \l6_pad  = \l1_pad ;
	assign \l7_pad  = _w435_ ;
	assign \l8_pad  = _w439_ ;
	assign \l9_pad  = _w442_ ;
	assign \m7_pad  = _w449_ ;
	assign \m8_pad  = _w453_ ;
	assign \m9_pad  = _w461_ ;
	assign \n5_pad  = _w463_ ;
	assign \n6_pad  = _w466_ ;
	assign \n7_pad  = _w473_ ;
	assign \n8_pad  = _w477_ ;
	assign \n9_pad  = _w485_ ;
	assign \o4_pad  = \g1_pad ;
	assign \o5_pad  = _w487_ ;
	assign \o6_pad  = _w488_ ;
	assign \o7_pad  = _w495_ ;
	assign \o8_pad  = _w499_ ;
	assign \o9_pad  = _w504_ ;
	assign \p4_pad  = _w510_ ;
	assign \p5_pad  = _w512_ ;
	assign \p6_pad  = _w518_ ;
	assign \p7_pad  = _w525_ ;
	assign \p8_pad  = _w529_ ;
	assign \p9_pad  = _w542_ ;
	assign \q4_pad  = _w548_ ;
	assign \q5_pad  = _w550_ ;
	assign \q6_pad  = _w556_ ;
	assign \q7_pad  = _w563_ ;
	assign \q8_pad  = _w567_ ;
	assign \q9_pad  = _w572_ ;
	assign \r4_pad  = _w578_ ;
	assign \r5_pad  = _w580_ ;
	assign \r6_pad  = _w588_ ;
	assign \r7_pad  = _w595_ ;
	assign \r8_pad  = _w599_ ;
	assign \r9_pad  = _w604_ ;
	assign \s4_pad  = _w610_ ;
	assign \s6_pad  = _w615_ ;
	assign \s7_pad  = _w622_ ;
	assign \s8_pad  = _w626_ ;
	assign \s9_pad  = _w649_ ;
	assign \t6_pad  = _w655_ ;
	assign \t7_pad  = _w665_ ;
	assign \t8_pad  = _w669_ ;
	assign \t9_pad  = _w671_ ;
	assign \u6_pad  = _w676_ ;
	assign \u7_pad  = _w686_ ;
	assign \u8_pad  = _w690_ ;
	assign \u9_pad  = _w691_ ;
	assign \v4_pad  = _w695_ ;
	assign \v6_pad  = _w700_ ;
	assign \v7_pad  = _w710_ ;
	assign \v8_pad  = _w714_ ;
	assign \v9_pad  = _w716_ ;
	assign \w4_pad  = _w720_ ;
	assign \w5_pad  = _w723_ ;
	assign \w6_pad  = _w730_ ;
	assign \w7_pad  = _w740_ ;
	assign \w8_pad  = _w744_ ;
	assign \w9_pad  = _w746_ ;
	assign \x4_pad  = _w750_ ;
	assign \x5_pad  = _w751_ ;
	assign \x6_pad  = _w758_ ;
	assign \x7_pad  = _w768_ ;
	assign \x8_pad  = _w772_ ;
	assign \y4_pad  = _w776_ ;
	assign \y5_pad  = _w777_ ;
	assign \y6_pad  = _w784_ ;
	assign \y7_pad  = _w794_ ;
	assign \y8_pad  = _w798_ ;
	assign \z4_pad  = _w802_ ;
	assign \z5_pad  = _w803_ ;
	assign \z6_pad  = _w810_ ;
	assign \z7_pad  = _w820_ ;
	assign \z8_pad  = _w824_ ;
endmodule;