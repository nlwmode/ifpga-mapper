module top( \g100_reg/NET0131  , \g1037_reg/NET0131  , \g103_reg/NET0131  , \g1041_reg/NET0131  , \g1045_reg/NET0131  , \g1049_reg/NET0131  , \g104_reg/NET0131  , \g1053_reg/NET0131  , \g1057_reg/NET0131  , \g1061_reg/NET0131  , \g1065_reg/NET0131  , \g1069_reg/NET0131  , \g1073_reg/NET0131  , \g1077_reg/NET0131  , \g1080_pad  , \g1087_reg/NET0131  , \g1092_reg/NET0131  , \g1097_reg/NET0131  , \g1098_reg/NET0131  , \g1102_reg/NET0131  , \g1106_reg/NET0131  , \g1110_reg/NET0131  , \g1114_reg/NET0131  , \g1118_reg/NET0131  , \g1122_reg/NET0131  , \g1126_reg/NET0131  , \g1130_reg/NET0131  , \g1134_reg/NET0131  , \g1138_reg/NET0131  , \g1142_reg/NET0131  , \g1148_reg/NET0131  , \g1149_reg/NET0131  , \g1158_reg/NET0131  , \g1166_reg/NET0131  , \g1176_reg/NET0131  , \g1179_reg/NET0131  , \g1189_reg/NET0131  , \g1207_reg/NET0131  , \g1211_reg/NET0131  , \g1214_reg/NET0131  , \g1217_reg/NET0131  , \g1220_reg/NET0131  , \g1223_reg/NET0131  , \g1224_reg/NET0131  , \g1225_reg/NET0131  , \g1226_reg/NET0131  , \g1227_reg/NET0131  , \g1228_reg/NET0131  , \g1229_reg/NET0131  , \g1230_reg/NET0131  , \g1231_reg/NET0131  , \g1247_reg/NET0131  , \g1251_reg/NET0131  , \g1252_reg/NET0131  , \g1253_reg/NET0131  , \g1257_reg/NET0131  , \g1260_reg/NET0131  , \g1263_reg/NET0131  , \g1266_reg/NET0131  , \g1268_reg/NET0131  , \g1269_reg/NET0131  , \g1272_reg/NET0131  , \g1276_reg/NET0131  , \g1280_reg/NET0131  , \g1284_reg/NET0131  , \g1288_reg/NET0131  , \g1292_reg/NET0131  , \g1296_reg/NET0131  , \g1300_reg/NET0131  , \g1304_reg/NET0131  , \g1307_reg/NET0131  , \g1313_reg/NET0131  , \g1317_reg/NET0131  , \g1318_reg/NET0131  , \g1319_reg/NET0131  , \g1320_reg/NET0131  , \g1321_reg/NET0131  , \g1322_reg/NET0131  , \g1323_reg/NET0131  , \g1324_reg/NET0131  , \g1325_reg/NET0131  , \g1326_reg/NET0131  , \g1327_reg/NET0131  , \g1328_reg/NET0131  , \g1329_reg/NET0131  , \g1330_reg/NET0131  , \g1333_reg/NET0131  , \g1336_reg/NET0131  , \g1339_reg/NET0131  , \g1342_reg/NET0131  , \g1345_reg/NET0131  , \g1348_reg/NET0131  , \g1351_reg/NET0131  , \g1354_reg/NET0131  , \g1357_reg/NET0131  , \g1360_reg/NET0131  , \g1363_reg/NET0131  , \g1364_reg/NET0131  , \g1365_reg/NET0131  , \g1366_reg/NET0131  , \g1367_reg/NET0131  , \g1368_reg/NET0131  , \g1369_reg/NET0131  , \g1370_reg/NET0131  , \g1371_reg/NET0131  , \g1372_reg/NET0131  , \g1373_reg/NET0131  , \g1374_reg/NET0131  , \g1375_reg/NET0131  , \g1405_reg/NET0131  , \g1408_reg/NET0131  , \g1412_reg/NET0131  , \g1415_reg/NET0131  , \g1416_reg/NET0131  , \g1421_reg/NET0131  , \g1428_reg/NET0131  , \g1430_reg/NET0131  , \g1432_reg/NET0131  , \g1435_reg/NET0131  , \g1439_reg/NET0131  , \g1444_reg/NET0131  , \g1450_reg/NET0131  , \g1454_reg/NET0131  , \g1462_reg/NET0131  , \g1467_reg/NET0131  , \g1472_reg/NET0131  , \g1481_reg/NET0131  , \g1486_reg/NET0131  , \g1489_reg/NET0131  , \g1494_reg/NET0131  , \g1499_reg/NET0131  , \g1504_reg/NET0131  , \g1509_reg/NET0131  , \g1514_reg/NET0131  , \g1519_reg/NET0131  , \g1944_pad  , \g2662_pad  , \g2888_pad  , \g2_reg/NET0131  , \g4370_pad  , \g4371_pad  , \g4372_pad  , \g4373_pad  , \g43_pad  , \g652_reg/NET0131  , \g7423_pad  , \g7424_pad  , \g7425_pad  , \g7504_pad  , \g7505_pad  , \g7507_pad  , \g7508_pad  , \g785_pad  , \g866_reg/NET0131  , \g871_reg/NET0131  , \g889_reg/NET0131  , \g929_reg/NET0131  , \g933_reg/NET0131  , \g936_reg/NET0131  , \g940_reg/NET0131  , \g942_reg/NET0131  , \g943_reg/NET0131  , \g944_reg/NET0131  , \g950_reg/NET0131  , \g951_reg/NET0131  , \g952_reg/NET0131  , \g953_reg/NET0131  , \g954_reg/NET0131  , \g962_pad  , \g1006_pad  , \g1158_reg/P0001  , \g1252_reg/P0001  , \g1260_reg/P0001  , \g1416_reg/NET0131_syn_2  , \g17/_0_  , \g19189/_0_  , \g19252/_0_  , \g19253/_0_  , \g19273/_3_  , \g19284/_0_  , \g19285/_0_  , \g19295/_3_  , \g19302/_0_  , \g19303/_0_  , \g19304/_0_  , \g19308/_0_  , \g19309/_0_  , \g19310/_0_  , \g19321/_0_  , \g19326/_3_  , \g19331/_0_  , \g19341/_0_  , \g19366/_0_  , \g19372/_3_  , \g19385/_0_  , \g19386/_0_  , \g19387/_0_  , \g19388/_0_  , \g19389/_0_  , \g19390/_0_  , \g19392/_0_  , \g19393/_0_  , \g19394/_0_  , \g19398/_0_  , \g19399/_0_  , \g19400/_0_  , \g19401/_0_  , \g19403/_0_  , \g19405/_0_  , \g19406/_0_  , \g19437/_0_  , \g19438/_0_  , \g19445/_0_  , \g19446/_0_  , \g19450/_3_  , \g19472/_0_  , \g19473/_0_  , \g19474/_0_  , \g19476/_0_  , \g19484/_0_  , \g19485/_0_  , \g19492/_0_  , \g19493/_0_  , \g19499/_0_  , \g19500/_0_  , \g19501/_0_  , \g19502/_0_  , \g19503/_0_  , \g19504/_0_  , \g19507/_3_  , \g19508/_3_  , \g19512/_3_  , \g19513/_3_  , \g19514/_3_  , \g19528/_0_  , \g19529/_0_  , \g19534/_0_  , \g19535/_0_  , \g19536/_0_  , \g19538/_0_  , \g19542/_0_  , \g19560/_0_  , \g19563/_0_  , \g19565/_0_  , \g19567/_0_  , \g19569/_1_  , \g19572/_0_  , \g19574/_3_  , \g19614/_0_  , \g19615/_0_  , \g19620/_0_  , \g19626/_0_  , \g19629/_0_  , \g19631/_0_  , \g19666/_0_  , \g19667/_0_  , \g19669/_0_  , \g19677/_0_  , \g19690/_3_  , \g19721/_0_  , \g19723/_0_  , \g19723/_1_  , \g19725/_2_  , \g19751/_0_  , \g19752/_0_  , \g19753/_0_  , \g19755/_0_  , \g19815/_0_  , \g19821/_0_  , \g19822/_0_  , \g19833/_0_  , \g19877/_0_  , \g19898/_0_  , \g19899/_0_  , \g19900/_0_  , \g19901/_0_  , \g19908/_0_  , \g19927/_0_  , \g19928/_0_  , \g19930/_0_  , \g19931/_0_  , \g19932/_0_  , \g19934/_0_  , \g19992/_0_  , \g19993/_0_  , \g20002/_0_  , \g20008/_0_  , \g20010/_0_  , \g20016/_0_  , \g20110/_0_  , \g20117/_0_  , \g20118/_0_  , \g20131/_0_  , \g20246/_0_  , \g20704/_0_  , \g20722/_0_  , \g20731/_0_  , \g20732/_2_  , \g20870/_0_  , \g20883/_0_  , \g20931/_0_  , \g20951/_0_  , \g20969/_0_  , \g20989/_0_  , \g21/_2_  , \g21070/_0_  , \g21108/_0_  , \g21122/_0_  , \g21152/_0_  , \g21191/_0_  , \g21279/_0_  , \g21316/_0_  , \g21323/_0_  , \g21349/_3_  , \g21352/_3_  , \g21464/_0_  , \g21472/_0_  , \g21484/_0_  , \g21510/_0_  , \g21517/_0_  , \g21608/_0_  , \g21625/_0_  , \g21644/_1_  , \g4655_pad  , \g6850_pad  , \g6895_pad  , \g7048_pad  , \g7103_pad  , \g7731_pad  , \g7732_pad  , \g8219_pad  , \g8663_pad  );
  input \g100_reg/NET0131  ;
  input \g1037_reg/NET0131  ;
  input \g103_reg/NET0131  ;
  input \g1041_reg/NET0131  ;
  input \g1045_reg/NET0131  ;
  input \g1049_reg/NET0131  ;
  input \g104_reg/NET0131  ;
  input \g1053_reg/NET0131  ;
  input \g1057_reg/NET0131  ;
  input \g1061_reg/NET0131  ;
  input \g1065_reg/NET0131  ;
  input \g1069_reg/NET0131  ;
  input \g1073_reg/NET0131  ;
  input \g1077_reg/NET0131  ;
  input \g1080_pad  ;
  input \g1087_reg/NET0131  ;
  input \g1092_reg/NET0131  ;
  input \g1097_reg/NET0131  ;
  input \g1098_reg/NET0131  ;
  input \g1102_reg/NET0131  ;
  input \g1106_reg/NET0131  ;
  input \g1110_reg/NET0131  ;
  input \g1114_reg/NET0131  ;
  input \g1118_reg/NET0131  ;
  input \g1122_reg/NET0131  ;
  input \g1126_reg/NET0131  ;
  input \g1130_reg/NET0131  ;
  input \g1134_reg/NET0131  ;
  input \g1138_reg/NET0131  ;
  input \g1142_reg/NET0131  ;
  input \g1148_reg/NET0131  ;
  input \g1149_reg/NET0131  ;
  input \g1158_reg/NET0131  ;
  input \g1166_reg/NET0131  ;
  input \g1176_reg/NET0131  ;
  input \g1179_reg/NET0131  ;
  input \g1189_reg/NET0131  ;
  input \g1207_reg/NET0131  ;
  input \g1211_reg/NET0131  ;
  input \g1214_reg/NET0131  ;
  input \g1217_reg/NET0131  ;
  input \g1220_reg/NET0131  ;
  input \g1223_reg/NET0131  ;
  input \g1224_reg/NET0131  ;
  input \g1225_reg/NET0131  ;
  input \g1226_reg/NET0131  ;
  input \g1227_reg/NET0131  ;
  input \g1228_reg/NET0131  ;
  input \g1229_reg/NET0131  ;
  input \g1230_reg/NET0131  ;
  input \g1231_reg/NET0131  ;
  input \g1247_reg/NET0131  ;
  input \g1251_reg/NET0131  ;
  input \g1252_reg/NET0131  ;
  input \g1253_reg/NET0131  ;
  input \g1257_reg/NET0131  ;
  input \g1260_reg/NET0131  ;
  input \g1263_reg/NET0131  ;
  input \g1266_reg/NET0131  ;
  input \g1268_reg/NET0131  ;
  input \g1269_reg/NET0131  ;
  input \g1272_reg/NET0131  ;
  input \g1276_reg/NET0131  ;
  input \g1280_reg/NET0131  ;
  input \g1284_reg/NET0131  ;
  input \g1288_reg/NET0131  ;
  input \g1292_reg/NET0131  ;
  input \g1296_reg/NET0131  ;
  input \g1300_reg/NET0131  ;
  input \g1304_reg/NET0131  ;
  input \g1307_reg/NET0131  ;
  input \g1313_reg/NET0131  ;
  input \g1317_reg/NET0131  ;
  input \g1318_reg/NET0131  ;
  input \g1319_reg/NET0131  ;
  input \g1320_reg/NET0131  ;
  input \g1321_reg/NET0131  ;
  input \g1322_reg/NET0131  ;
  input \g1323_reg/NET0131  ;
  input \g1324_reg/NET0131  ;
  input \g1325_reg/NET0131  ;
  input \g1326_reg/NET0131  ;
  input \g1327_reg/NET0131  ;
  input \g1328_reg/NET0131  ;
  input \g1329_reg/NET0131  ;
  input \g1330_reg/NET0131  ;
  input \g1333_reg/NET0131  ;
  input \g1336_reg/NET0131  ;
  input \g1339_reg/NET0131  ;
  input \g1342_reg/NET0131  ;
  input \g1345_reg/NET0131  ;
  input \g1348_reg/NET0131  ;
  input \g1351_reg/NET0131  ;
  input \g1354_reg/NET0131  ;
  input \g1357_reg/NET0131  ;
  input \g1360_reg/NET0131  ;
  input \g1363_reg/NET0131  ;
  input \g1364_reg/NET0131  ;
  input \g1365_reg/NET0131  ;
  input \g1366_reg/NET0131  ;
  input \g1367_reg/NET0131  ;
  input \g1368_reg/NET0131  ;
  input \g1369_reg/NET0131  ;
  input \g1370_reg/NET0131  ;
  input \g1371_reg/NET0131  ;
  input \g1372_reg/NET0131  ;
  input \g1373_reg/NET0131  ;
  input \g1374_reg/NET0131  ;
  input \g1375_reg/NET0131  ;
  input \g1405_reg/NET0131  ;
  input \g1408_reg/NET0131  ;
  input \g1412_reg/NET0131  ;
  input \g1415_reg/NET0131  ;
  input \g1416_reg/NET0131  ;
  input \g1421_reg/NET0131  ;
  input \g1428_reg/NET0131  ;
  input \g1430_reg/NET0131  ;
  input \g1432_reg/NET0131  ;
  input \g1435_reg/NET0131  ;
  input \g1439_reg/NET0131  ;
  input \g1444_reg/NET0131  ;
  input \g1450_reg/NET0131  ;
  input \g1454_reg/NET0131  ;
  input \g1462_reg/NET0131  ;
  input \g1467_reg/NET0131  ;
  input \g1472_reg/NET0131  ;
  input \g1481_reg/NET0131  ;
  input \g1486_reg/NET0131  ;
  input \g1489_reg/NET0131  ;
  input \g1494_reg/NET0131  ;
  input \g1499_reg/NET0131  ;
  input \g1504_reg/NET0131  ;
  input \g1509_reg/NET0131  ;
  input \g1514_reg/NET0131  ;
  input \g1519_reg/NET0131  ;
  input \g1944_pad  ;
  input \g2662_pad  ;
  input \g2888_pad  ;
  input \g2_reg/NET0131  ;
  input \g4370_pad  ;
  input \g4371_pad  ;
  input \g4372_pad  ;
  input \g4373_pad  ;
  input \g43_pad  ;
  input \g652_reg/NET0131  ;
  input \g7423_pad  ;
  input \g7424_pad  ;
  input \g7425_pad  ;
  input \g7504_pad  ;
  input \g7505_pad  ;
  input \g7507_pad  ;
  input \g7508_pad  ;
  input \g785_pad  ;
  input \g866_reg/NET0131  ;
  input \g871_reg/NET0131  ;
  input \g889_reg/NET0131  ;
  input \g929_reg/NET0131  ;
  input \g933_reg/NET0131  ;
  input \g936_reg/NET0131  ;
  input \g940_reg/NET0131  ;
  input \g942_reg/NET0131  ;
  input \g943_reg/NET0131  ;
  input \g944_reg/NET0131  ;
  input \g950_reg/NET0131  ;
  input \g951_reg/NET0131  ;
  input \g952_reg/NET0131  ;
  input \g953_reg/NET0131  ;
  input \g954_reg/NET0131  ;
  input \g962_pad  ;
  output \g1006_pad  ;
  output \g1158_reg/P0001  ;
  output \g1252_reg/P0001  ;
  output \g1260_reg/P0001  ;
  output \g1416_reg/NET0131_syn_2  ;
  output \g17/_0_  ;
  output \g19189/_0_  ;
  output \g19252/_0_  ;
  output \g19253/_0_  ;
  output \g19273/_3_  ;
  output \g19284/_0_  ;
  output \g19285/_0_  ;
  output \g19295/_3_  ;
  output \g19302/_0_  ;
  output \g19303/_0_  ;
  output \g19304/_0_  ;
  output \g19308/_0_  ;
  output \g19309/_0_  ;
  output \g19310/_0_  ;
  output \g19321/_0_  ;
  output \g19326/_3_  ;
  output \g19331/_0_  ;
  output \g19341/_0_  ;
  output \g19366/_0_  ;
  output \g19372/_3_  ;
  output \g19385/_0_  ;
  output \g19386/_0_  ;
  output \g19387/_0_  ;
  output \g19388/_0_  ;
  output \g19389/_0_  ;
  output \g19390/_0_  ;
  output \g19392/_0_  ;
  output \g19393/_0_  ;
  output \g19394/_0_  ;
  output \g19398/_0_  ;
  output \g19399/_0_  ;
  output \g19400/_0_  ;
  output \g19401/_0_  ;
  output \g19403/_0_  ;
  output \g19405/_0_  ;
  output \g19406/_0_  ;
  output \g19437/_0_  ;
  output \g19438/_0_  ;
  output \g19445/_0_  ;
  output \g19446/_0_  ;
  output \g19450/_3_  ;
  output \g19472/_0_  ;
  output \g19473/_0_  ;
  output \g19474/_0_  ;
  output \g19476/_0_  ;
  output \g19484/_0_  ;
  output \g19485/_0_  ;
  output \g19492/_0_  ;
  output \g19493/_0_  ;
  output \g19499/_0_  ;
  output \g19500/_0_  ;
  output \g19501/_0_  ;
  output \g19502/_0_  ;
  output \g19503/_0_  ;
  output \g19504/_0_  ;
  output \g19507/_3_  ;
  output \g19508/_3_  ;
  output \g19512/_3_  ;
  output \g19513/_3_  ;
  output \g19514/_3_  ;
  output \g19528/_0_  ;
  output \g19529/_0_  ;
  output \g19534/_0_  ;
  output \g19535/_0_  ;
  output \g19536/_0_  ;
  output \g19538/_0_  ;
  output \g19542/_0_  ;
  output \g19560/_0_  ;
  output \g19563/_0_  ;
  output \g19565/_0_  ;
  output \g19567/_0_  ;
  output \g19569/_1_  ;
  output \g19572/_0_  ;
  output \g19574/_3_  ;
  output \g19614/_0_  ;
  output \g19615/_0_  ;
  output \g19620/_0_  ;
  output \g19626/_0_  ;
  output \g19629/_0_  ;
  output \g19631/_0_  ;
  output \g19666/_0_  ;
  output \g19667/_0_  ;
  output \g19669/_0_  ;
  output \g19677/_0_  ;
  output \g19690/_3_  ;
  output \g19721/_0_  ;
  output \g19723/_0_  ;
  output \g19723/_1_  ;
  output \g19725/_2_  ;
  output \g19751/_0_  ;
  output \g19752/_0_  ;
  output \g19753/_0_  ;
  output \g19755/_0_  ;
  output \g19815/_0_  ;
  output \g19821/_0_  ;
  output \g19822/_0_  ;
  output \g19833/_0_  ;
  output \g19877/_0_  ;
  output \g19898/_0_  ;
  output \g19899/_0_  ;
  output \g19900/_0_  ;
  output \g19901/_0_  ;
  output \g19908/_0_  ;
  output \g19927/_0_  ;
  output \g19928/_0_  ;
  output \g19930/_0_  ;
  output \g19931/_0_  ;
  output \g19932/_0_  ;
  output \g19934/_0_  ;
  output \g19992/_0_  ;
  output \g19993/_0_  ;
  output \g20002/_0_  ;
  output \g20008/_0_  ;
  output \g20010/_0_  ;
  output \g20016/_0_  ;
  output \g20110/_0_  ;
  output \g20117/_0_  ;
  output \g20118/_0_  ;
  output \g20131/_0_  ;
  output \g20246/_0_  ;
  output \g20704/_0_  ;
  output \g20722/_0_  ;
  output \g20731/_0_  ;
  output \g20732/_2_  ;
  output \g20870/_0_  ;
  output \g20883/_0_  ;
  output \g20931/_0_  ;
  output \g20951/_0_  ;
  output \g20969/_0_  ;
  output \g20989/_0_  ;
  output \g21/_2_  ;
  output \g21070/_0_  ;
  output \g21108/_0_  ;
  output \g21122/_0_  ;
  output \g21152/_0_  ;
  output \g21191/_0_  ;
  output \g21279/_0_  ;
  output \g21316/_0_  ;
  output \g21323/_0_  ;
  output \g21349/_3_  ;
  output \g21352/_3_  ;
  output \g21464/_0_  ;
  output \g21472/_0_  ;
  output \g21484/_0_  ;
  output \g21510/_0_  ;
  output \g21517/_0_  ;
  output \g21608/_0_  ;
  output \g21625/_0_  ;
  output \g21644/_1_  ;
  output \g4655_pad  ;
  output \g6850_pad  ;
  output \g6895_pad  ;
  output \g7048_pad  ;
  output \g7103_pad  ;
  output \g7731_pad  ;
  output \g7732_pad  ;
  output \g8219_pad  ;
  output \g8663_pad  ;
  wire n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 ;
  assign n170 = \g1330_reg/NET0131  & \g1333_reg/NET0131  ;
  assign n171 = \g1336_reg/NET0131  & \g1339_reg/NET0131  ;
  assign n172 = n170 & n171 ;
  assign n173 = \g1342_reg/NET0131  & \g1345_reg/NET0131  ;
  assign n174 = n172 & n173 ;
  assign n175 = ~\g1348_reg/NET0131  & ~n174 ;
  assign n176 = \g1348_reg/NET0131  & n173 ;
  assign n177 = n172 & n176 ;
  assign n178 = \g1247_reg/NET0131  & ~n177 ;
  assign n179 = ~n175 & n178 ;
  assign n180 = \g1073_reg/NET0131  & ~\g1158_reg/NET0131  ;
  assign n181 = \g1092_reg/NET0131  & \g1130_reg/NET0131  ;
  assign n182 = \g1134_reg/NET0131  & \g1138_reg/NET0131  ;
  assign n183 = n181 & n182 ;
  assign n184 = \g1045_reg/NET0131  & \g1149_reg/NET0131  ;
  assign n185 = \g1037_reg/NET0131  & \g1041_reg/NET0131  ;
  assign n186 = n184 & n185 ;
  assign n187 = n183 & n186 ;
  assign n188 = \g1049_reg/NET0131  & \g1053_reg/NET0131  ;
  assign n189 = \g1057_reg/NET0131  & \g1061_reg/NET0131  ;
  assign n190 = n188 & n189 ;
  assign n191 = \g1065_reg/NET0131  & n190 ;
  assign n192 = n187 & n191 ;
  assign n193 = ~\g1073_reg/NET0131  & \g1158_reg/NET0131  ;
  assign n194 = \g1069_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n195 = n193 & n194 ;
  assign n196 = n192 & n195 ;
  assign n197 = ~n180 & ~n196 ;
  assign n198 = \g936_reg/NET0131  & ~\g940_reg/NET0131  ;
  assign n199 = ~\g936_reg/NET0131  & \g940_reg/NET0131  ;
  assign n200 = ~\g943_reg/NET0131  & n199 ;
  assign n201 = ~n198 & ~n200 ;
  assign n202 = \g1158_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n203 = \g1073_reg/NET0131  & \g1158_reg/NET0131  ;
  assign n204 = ~n202 & ~n203 ;
  assign n205 = \g1049_reg/NET0131  & n204 ;
  assign n206 = \g1049_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n207 = n193 & n206 ;
  assign n208 = ~n187 & n207 ;
  assign n209 = ~\g1049_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n210 = n193 & n209 ;
  assign n211 = n187 & n210 ;
  assign n212 = ~n208 & ~n211 ;
  assign n213 = ~n205 & n212 ;
  assign n214 = \g954_reg/NET0131  & ~n198 ;
  assign n215 = \g2_reg/NET0131  & n198 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = ~\g1251_reg/NET0131  & \g1481_reg/NET0131  ;
  assign n218 = \g1489_reg/NET0131  & \g1494_reg/NET0131  ;
  assign n219 = n217 & n218 ;
  assign n220 = \g1499_reg/NET0131  & \g1504_reg/NET0131  ;
  assign n221 = \g1509_reg/NET0131  & n220 ;
  assign n222 = n219 & n221 ;
  assign n223 = ~\g1514_reg/NET0131  & ~n222 ;
  assign n224 = \g1462_reg/NET0131  & \g1467_reg/NET0131  ;
  assign n225 = \g1514_reg/NET0131  & \g1519_reg/NET0131  ;
  assign n226 = \g1472_reg/NET0131  & \g1499_reg/NET0131  ;
  assign n227 = n225 & n226 ;
  assign n228 = n224 & n227 ;
  assign n229 = n219 & n228 ;
  assign n230 = \g1509_reg/NET0131  & \g1514_reg/NET0131  ;
  assign n231 = n220 & n230 ;
  assign n232 = n219 & n231 ;
  assign n233 = ~n229 & ~n232 ;
  assign n234 = ~n223 & n233 ;
  assign n235 = \g1087_reg/NET0131  & \g1098_reg/NET0131  ;
  assign n236 = \g1102_reg/NET0131  & \g1106_reg/NET0131  ;
  assign n237 = n235 & n236 ;
  assign n238 = \g1110_reg/NET0131  & \g1148_reg/NET0131  ;
  assign n239 = \g1114_reg/NET0131  & n238 ;
  assign n240 = n237 & n239 ;
  assign n241 = ~\g1097_reg/NET0131  & ~\g1118_reg/NET0131  ;
  assign n242 = ~n240 & n241 ;
  assign n243 = ~\g1097_reg/NET0131  & \g1114_reg/NET0131  ;
  assign n244 = n238 & n243 ;
  assign n245 = n237 & n244 ;
  assign n246 = \g1118_reg/NET0131  & n245 ;
  assign n247 = ~n242 & ~n246 ;
  assign n248 = \g953_reg/NET0131  & ~n198 ;
  assign n249 = ~n215 & ~n248 ;
  assign n250 = \g1148_reg/NET0131  & n237 ;
  assign n251 = \g1102_reg/NET0131  & \g1148_reg/NET0131  ;
  assign n252 = n235 & n251 ;
  assign n253 = ~\g1106_reg/NET0131  & ~n252 ;
  assign n254 = ~n250 & ~n253 ;
  assign n255 = ~\g1097_reg/NET0131  & ~n254 ;
  assign n256 = ~\g1097_reg/NET0131  & ~\g1110_reg/NET0131  ;
  assign n257 = ~n250 & n256 ;
  assign n258 = ~\g1097_reg/NET0131  & \g1110_reg/NET0131  ;
  assign n259 = \g1148_reg/NET0131  & n258 ;
  assign n260 = n237 & n259 ;
  assign n261 = ~n257 & ~n260 ;
  assign n262 = n237 & n238 ;
  assign n263 = ~\g1097_reg/NET0131  & ~\g1114_reg/NET0131  ;
  assign n264 = ~n262 & n263 ;
  assign n265 = ~n245 & ~n264 ;
  assign n266 = n219 & n220 ;
  assign n267 = ~\g1509_reg/NET0131  & ~n266 ;
  assign n268 = ~n222 & ~n267 ;
  assign n269 = ~n229 & n268 ;
  assign n270 = ~\g1097_reg/NET0131  & ~\g1148_reg/NET0131  ;
  assign n271 = \g1098_reg/NET0131  & n270 ;
  assign n272 = ~\g1097_reg/NET0131  & \g1148_reg/NET0131  ;
  assign n273 = ~\g1087_reg/NET0131  & ~\g1098_reg/NET0131  ;
  assign n274 = ~n235 & ~n273 ;
  assign n275 = n272 & n274 ;
  assign n276 = ~n271 & ~n275 ;
  assign n277 = ~\g1102_reg/NET0131  & ~n235 ;
  assign n278 = ~\g1102_reg/NET0131  & ~\g1148_reg/NET0131  ;
  assign n279 = ~\g1097_reg/NET0131  & ~n278 ;
  assign n280 = ~n252 & n279 ;
  assign n281 = ~n277 & n280 ;
  assign n282 = \g1037_reg/NET0131  & n204 ;
  assign n283 = \g1149_reg/NET0131  & n183 ;
  assign n284 = ~\g1037_reg/NET0131  & ~n283 ;
  assign n285 = ~\g1251_reg/NET0131  & n193 ;
  assign n286 = \g1037_reg/NET0131  & \g1149_reg/NET0131  ;
  assign n287 = n183 & n286 ;
  assign n288 = n285 & ~n287 ;
  assign n289 = ~n284 & n288 ;
  assign n290 = ~n282 & ~n289 ;
  assign n291 = \g952_reg/NET0131  & ~n198 ;
  assign n292 = ~n215 & ~n291 ;
  assign n293 = \g1087_reg/NET0131  & ~\g1148_reg/NET0131  ;
  assign n294 = ~\g1087_reg/NET0131  & \g1148_reg/NET0131  ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = ~\g1097_reg/NET0131  & ~n295 ;
  assign n297 = \g1499_reg/NET0131  & n219 ;
  assign n298 = ~\g1504_reg/NET0131  & ~n297 ;
  assign n299 = ~n229 & ~n298 ;
  assign n300 = ~n266 & n299 ;
  assign n301 = ~\g1149_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n302 = n193 & n301 ;
  assign n303 = n183 & n302 ;
  assign n304 = \g1149_reg/NET0131  & n204 ;
  assign n305 = ~\g1073_reg/NET0131  & \g1149_reg/NET0131  ;
  assign n306 = n202 & n305 ;
  assign n307 = ~n183 & n306 ;
  assign n308 = ~n304 & ~n307 ;
  assign n309 = ~n303 & n308 ;
  assign n310 = \g951_reg/NET0131  & ~n198 ;
  assign n311 = ~n215 & ~n310 ;
  assign n312 = ~\g1092_reg/NET0131  & n202 ;
  assign n313 = \g1092_reg/NET0131  & ~n202 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n203 & ~n314 ;
  assign n316 = \g1313_reg/NET0131  & \g1317_reg/NET0131  ;
  assign n317 = ~\g1318_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n318 = n316 & n317 ;
  assign n319 = \g100_reg/NET0131  & \g1329_reg/NET0131  ;
  assign n320 = \g1318_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n321 = ~n316 & n320 ;
  assign n322 = ~n319 & ~n321 ;
  assign n323 = ~n318 & n322 ;
  assign n324 = \g1251_reg/NET0131  & ~\g1481_reg/NET0131  ;
  assign n325 = ~n217 & ~n324 ;
  assign n326 = \g1489_reg/NET0131  & n217 ;
  assign n327 = ~\g1489_reg/NET0131  & ~n217 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = \g1318_reg/NET0131  & \g1319_reg/NET0131  ;
  assign n330 = n316 & n329 ;
  assign n331 = \g1320_reg/NET0131  & \g1321_reg/NET0131  ;
  assign n332 = \g1322_reg/NET0131  & \g1323_reg/NET0131  ;
  assign n333 = n331 & n332 ;
  assign n334 = n330 & n333 ;
  assign n335 = ~\g1324_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n336 = n334 & n335 ;
  assign n337 = \g103_reg/NET0131  & \g1329_reg/NET0131  ;
  assign n338 = \g1324_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n339 = ~n334 & n338 ;
  assign n340 = ~n337 & ~n339 ;
  assign n341 = ~n336 & n340 ;
  assign n342 = \g1348_reg/NET0131  & \g1351_reg/NET0131  ;
  assign n343 = n173 & n342 ;
  assign n344 = n172 & n343 ;
  assign n345 = \g1247_reg/NET0131  & \g1354_reg/NET0131  ;
  assign n346 = ~n344 & n345 ;
  assign n347 = \g1247_reg/NET0131  & ~\g1354_reg/NET0131  ;
  assign n348 = n344 & n347 ;
  assign n349 = ~n346 & ~n348 ;
  assign n350 = ~\g1371_reg/NET0131  & ~\g1372_reg/NET0131  ;
  assign n351 = ~\g1369_reg/NET0131  & n350 ;
  assign n352 = ~\g1373_reg/NET0131  & ~\g1374_reg/NET0131  ;
  assign n353 = ~\g1370_reg/NET0131  & ~\g1375_reg/NET0131  ;
  assign n354 = n352 & n353 ;
  assign n355 = n351 & n354 ;
  assign n356 = ~\g1363_reg/NET0131  & ~\g1364_reg/NET0131  ;
  assign n357 = ~\g1367_reg/NET0131  & ~\g1368_reg/NET0131  ;
  assign n358 = ~\g1365_reg/NET0131  & ~\g1366_reg/NET0131  ;
  assign n359 = n357 & n358 ;
  assign n360 = n356 & n359 ;
  assign n361 = n355 & n360 ;
  assign n362 = \g1324_reg/NET0131  & \g1328_reg/NET0131  ;
  assign n363 = \g1325_reg/NET0131  & \g1326_reg/NET0131  ;
  assign n364 = \g1327_reg/NET0131  & n363 ;
  assign n365 = n362 & n364 ;
  assign n366 = n334 & n365 ;
  assign n367 = ~\g7504_pad  & ~n366 ;
  assign n368 = ~\g1329_reg/NET0131  & ~n367 ;
  assign n369 = \g929_reg/NET0131  & \g933_reg/NET0131  ;
  assign n370 = \g871_reg/NET0131  & ~\g889_reg/NET0131  ;
  assign n371 = n369 & n370 ;
  assign n372 = ~\g785_pad  & ~n371 ;
  assign n373 = \g1324_reg/NET0131  & \g1325_reg/NET0131  ;
  assign n374 = n334 & n373 ;
  assign n375 = \g1326_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n376 = ~n374 & n375 ;
  assign n377 = \g1325_reg/NET0131  & ~\g1326_reg/NET0131  ;
  assign n378 = n338 & n377 ;
  assign n379 = n334 & n378 ;
  assign n380 = ~n337 & ~n379 ;
  assign n381 = ~n376 & n380 ;
  assign n382 = \g1134_reg/NET0131  & n204 ;
  assign n383 = ~\g1134_reg/NET0131  & ~n181 ;
  assign n384 = \g1134_reg/NET0131  & n181 ;
  assign n385 = ~n383 & ~n384 ;
  assign n386 = n285 & n385 ;
  assign n387 = ~n382 & ~n386 ;
  assign n388 = n330 & n331 ;
  assign n389 = ~n319 & n388 ;
  assign n390 = \g1320_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n391 = n330 & n390 ;
  assign n392 = \g1321_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n393 = ~n319 & ~n392 ;
  assign n394 = ~n391 & n393 ;
  assign n395 = ~n389 & ~n394 ;
  assign n396 = \g1138_reg/NET0131  & n204 ;
  assign n397 = ~\g1138_reg/NET0131  & ~n384 ;
  assign n398 = ~n183 & n285 ;
  assign n399 = ~n397 & n398 ;
  assign n400 = ~n396 & ~n399 ;
  assign n401 = \g1130_reg/NET0131  & n204 ;
  assign n402 = ~\g1092_reg/NET0131  & ~\g1130_reg/NET0131  ;
  assign n403 = ~n181 & ~n402 ;
  assign n404 = n285 & n403 ;
  assign n405 = ~n401 & ~n404 ;
  assign n406 = \g1405_reg/NET0131  & \g1408_reg/NET0131  ;
  assign n407 = ~\g1231_reg/NET0131  & ~\g1428_reg/NET0131  ;
  assign n408 = ~n406 & n407 ;
  assign n409 = \g1412_reg/NET0131  & \g1415_reg/NET0131  ;
  assign n410 = ~\g1231_reg/NET0131  & ~\g1430_reg/NET0131  ;
  assign n411 = ~n409 & n410 ;
  assign n412 = \g1272_reg/NET0131  & \g1307_reg/NET0131  ;
  assign n413 = \g1276_reg/NET0131  & n412 ;
  assign n414 = ~\g1280_reg/NET0131  & ~n413 ;
  assign n415 = \g1276_reg/NET0131  & \g1280_reg/NET0131  ;
  assign n416 = n412 & n415 ;
  assign n417 = ~\g1304_reg/NET0131  & ~n416 ;
  assign n418 = ~n414 & n417 ;
  assign n419 = \g1280_reg/NET0131  & \g1284_reg/NET0131  ;
  assign n420 = \g1272_reg/NET0131  & \g1276_reg/NET0131  ;
  assign n421 = n419 & n420 ;
  assign n422 = \g1288_reg/NET0131  & \g1307_reg/NET0131  ;
  assign n423 = n421 & n422 ;
  assign n424 = ~\g1292_reg/NET0131  & ~n423 ;
  assign n425 = \g1292_reg/NET0131  & n422 ;
  assign n426 = n421 & n425 ;
  assign n427 = ~\g1304_reg/NET0131  & ~n426 ;
  assign n428 = ~n424 & n427 ;
  assign n429 = \g1296_reg/NET0131  & \g1300_reg/NET0131  ;
  assign n430 = n426 & n429 ;
  assign n431 = \g1296_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n432 = \g1300_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n433 = n426 & n432 ;
  assign n434 = ~n431 & ~n433 ;
  assign n435 = ~n430 & ~n434 ;
  assign n436 = ~n426 & n432 ;
  assign n437 = \g1292_reg/NET0131  & ~\g1300_reg/NET0131  ;
  assign n438 = n422 & n437 ;
  assign n439 = n421 & n438 ;
  assign n440 = ~\g1304_reg/NET0131  & n439 ;
  assign n441 = ~n436 & ~n440 ;
  assign n442 = \g1276_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n443 = ~n412 & n442 ;
  assign n444 = ~\g1276_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n445 = n412 & n444 ;
  assign n446 = ~n443 & ~n445 ;
  assign n447 = \g1432_reg/NET0131  & \g1439_reg/NET0131  ;
  assign n448 = ~\g1430_reg/NET0131  & \g1435_reg/NET0131  ;
  assign n449 = ~n447 & n448 ;
  assign n450 = ~\g1430_reg/NET0131  & ~n447 ;
  assign n451 = \g1435_reg/NET0131  & \g1439_reg/NET0131  ;
  assign n452 = ~\g1435_reg/NET0131  & ~\g1439_reg/NET0131  ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = n450 & n453 ;
  assign n455 = ~\g1430_reg/NET0131  & ~\g7507_pad  ;
  assign n456 = ~n447 & n455 ;
  assign n457 = ~\g1430_reg/NET0131  & \g7507_pad  ;
  assign n458 = n447 & n457 ;
  assign n459 = ~n456 & ~n458 ;
  assign n460 = ~\g1432_reg/NET0131  & ~n451 ;
  assign n461 = n450 & ~n460 ;
  assign n462 = ~\g1284_reg/NET0131  & ~n416 ;
  assign n463 = \g1307_reg/NET0131  & n421 ;
  assign n464 = ~\g1304_reg/NET0131  & ~n463 ;
  assign n465 = ~n462 & n464 ;
  assign n466 = ~\g1288_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n467 = ~n463 & n466 ;
  assign n468 = \g1288_reg/NET0131  & \g1292_reg/NET0131  ;
  assign n469 = n429 & n468 ;
  assign n470 = \g1288_reg/NET0131  & ~\g1304_reg/NET0131  ;
  assign n471 = ~n469 & n470 ;
  assign n472 = n463 & n471 ;
  assign n473 = ~n467 & ~n472 ;
  assign n474 = \g1211_reg/NET0131  & \g1214_reg/NET0131  ;
  assign n475 = \g1207_reg/NET0131  & \g1217_reg/NET0131  ;
  assign n476 = n474 & n475 ;
  assign n477 = \g1220_reg/NET0131  & n476 ;
  assign n478 = ~\g1223_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n479 = ~n477 & n478 ;
  assign n480 = \g1223_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n481 = \g1220_reg/NET0131  & n480 ;
  assign n482 = n476 & n481 ;
  assign n483 = ~n479 & ~n482 ;
  assign n484 = ~\g1304_reg/NET0131  & ~n412 ;
  assign n485 = ~\g1272_reg/NET0131  & ~\g1307_reg/NET0131  ;
  assign n486 = n484 & ~n485 ;
  assign n487 = ~\g1313_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n488 = ~n319 & ~n487 ;
  assign n489 = ~\g1322_reg/NET0131  & ~n388 ;
  assign n490 = \g1322_reg/NET0131  & n331 ;
  assign n491 = n330 & n490 ;
  assign n492 = ~\g1329_reg/NET0131  & ~n491 ;
  assign n493 = ~n489 & n492 ;
  assign n494 = ~n319 & ~n493 ;
  assign n495 = ~\g1323_reg/NET0131  & ~n491 ;
  assign n496 = ~\g1329_reg/NET0131  & ~n334 ;
  assign n497 = ~n495 & n496 ;
  assign n498 = ~n319 & ~n497 ;
  assign n499 = ~\g1329_reg/NET0131  & ~n374 ;
  assign n500 = \g1324_reg/NET0131  & n334 ;
  assign n501 = ~\g1325_reg/NET0131  & ~n500 ;
  assign n502 = n499 & ~n501 ;
  assign n503 = ~n337 & ~n502 ;
  assign n504 = \g1318_reg/NET0131  & n316 ;
  assign n505 = ~\g1319_reg/NET0131  & ~n504 ;
  assign n506 = ~\g1329_reg/NET0131  & ~n330 ;
  assign n507 = ~n505 & n506 ;
  assign n508 = ~n319 & ~n507 ;
  assign n509 = \g1324_reg/NET0131  & n363 ;
  assign n510 = n334 & n509 ;
  assign n511 = ~\g1327_reg/NET0131  & ~n510 ;
  assign n512 = \g1324_reg/NET0131  & \g1327_reg/NET0131  ;
  assign n513 = n363 & n512 ;
  assign n514 = n334 & n513 ;
  assign n515 = ~\g1329_reg/NET0131  & ~n514 ;
  assign n516 = ~n511 & n515 ;
  assign n517 = ~n337 & ~n516 ;
  assign n518 = ~\g1494_reg/NET0131  & ~n326 ;
  assign n519 = ~n219 & ~n518 ;
  assign n520 = ~\g1499_reg/NET0131  & ~n219 ;
  assign n521 = ~n297 & ~n520 ;
  assign n522 = ~\g1313_reg/NET0131  & ~\g1317_reg/NET0131  ;
  assign n523 = ~\g1329_reg/NET0131  & ~n316 ;
  assign n524 = ~n522 & n523 ;
  assign n525 = ~n319 & ~n524 ;
  assign n526 = \g950_reg/NET0131  & ~n198 ;
  assign n527 = ~n215 & ~n526 ;
  assign n528 = ~\g1320_reg/NET0131  & ~\g1329_reg/NET0131  ;
  assign n529 = n330 & n528 ;
  assign n530 = ~n330 & n390 ;
  assign n531 = ~n319 & ~n530 ;
  assign n532 = ~n529 & n531 ;
  assign n533 = \g1450_reg/NET0131  & \g1454_reg/NET0131  ;
  assign n534 = ~\g1307_reg/NET0131  & \g1444_reg/NET0131  ;
  assign n535 = ~n533 & n534 ;
  assign n536 = \g1444_reg/NET0131  & ~\g1450_reg/NET0131  ;
  assign n537 = ~\g1307_reg/NET0131  & n536 ;
  assign n538 = ~\g1444_reg/NET0131  & \g1450_reg/NET0131  ;
  assign n539 = ~\g1307_reg/NET0131  & ~\g1454_reg/NET0131  ;
  assign n540 = n538 & n539 ;
  assign n541 = ~n537 & ~n540 ;
  assign n542 = ~\g1405_reg/NET0131  & n407 ;
  assign n543 = ~\g1412_reg/NET0131  & n410 ;
  assign n544 = ~\g1307_reg/NET0131  & \g1416_reg/NET0131  ;
  assign n545 = ~\g1421_reg/NET0131  & n544 ;
  assign n546 = ~\g1307_reg/NET0131  & ~n533 ;
  assign n547 = \g1444_reg/NET0131  & \g1450_reg/NET0131  ;
  assign n548 = ~\g1454_reg/NET0131  & ~n547 ;
  assign n549 = n546 & ~n548 ;
  assign n550 = ~\g7507_pad  & ~\g7508_pad  ;
  assign n551 = n447 & n550 ;
  assign n552 = ~\g1430_reg/NET0131  & ~\g7508_pad  ;
  assign n553 = n447 & n455 ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~n551 & ~n554 ;
  assign n556 = ~\g1354_reg/NET0131  & ~\g1357_reg/NET0131  ;
  assign n557 = ~\g1348_reg/NET0131  & ~\g1351_reg/NET0131  ;
  assign n558 = ~\g1342_reg/NET0131  & n557 ;
  assign n559 = ~\g104_reg/NET0131  & ~\g1336_reg/NET0131  ;
  assign n560 = ~\g1345_reg/NET0131  & ~\g1360_reg/NET0131  ;
  assign n561 = n559 & n560 ;
  assign n562 = n558 & n561 ;
  assign n563 = n556 & n562 ;
  assign n564 = \g104_reg/NET0131  & \g1336_reg/NET0131  ;
  assign n565 = \g1354_reg/NET0131  & \g1357_reg/NET0131  ;
  assign n566 = \g1360_reg/NET0131  & n565 ;
  assign n567 = n564 & n566 ;
  assign n568 = n343 & n567 ;
  assign n569 = ~n563 & ~n568 ;
  assign n570 = ~\g1330_reg/NET0131  & ~\g1333_reg/NET0131  ;
  assign n571 = \g104_reg/NET0131  & \g1339_reg/NET0131  ;
  assign n572 = ~n570 & ~n571 ;
  assign n573 = ~\g104_reg/NET0131  & ~\g1339_reg/NET0131  ;
  assign n574 = ~n170 & ~n573 ;
  assign n575 = ~n572 & ~n574 ;
  assign n576 = ~n569 & n575 ;
  assign n577 = \g1077_reg/NET0131  & \g2888_pad  ;
  assign n578 = \g1158_reg/NET0131  & \g652_reg/NET0131  ;
  assign n579 = \g1176_reg/NET0131  & n578 ;
  assign n580 = ~n577 & ~n579 ;
  assign n581 = \g1247_reg/NET0131  & ~n170 ;
  assign n582 = ~n570 & n581 ;
  assign n583 = ~\g1351_reg/NET0131  & ~n177 ;
  assign n584 = \g1247_reg/NET0131  & ~n344 ;
  assign n585 = ~n583 & n584 ;
  assign n586 = ~\g785_pad  & \g866_reg/NET0131  ;
  assign n587 = \g889_reg/NET0131  & n586 ;
  assign n588 = \g1179_reg/NET0131  & n578 ;
  assign n589 = ~\g2888_pad  & ~n588 ;
  assign n590 = \g1179_reg/NET0131  & \g2888_pad  ;
  assign n591 = n578 & n590 ;
  assign n592 = ~n577 & ~n591 ;
  assign n593 = ~n589 & n592 ;
  assign n594 = ~\g1176_reg/NET0131  & \g1944_pad  ;
  assign n595 = \g1080_pad  & ~\g1944_pad  ;
  assign n596 = ~n594 & ~n595 ;
  assign n597 = \g1223_reg/NET0131  & \g1224_reg/NET0131  ;
  assign n598 = \g1220_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n599 = n597 & n598 ;
  assign n600 = n476 & n599 ;
  assign n601 = ~\g1224_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n602 = \g1220_reg/NET0131  & \g1223_reg/NET0131  ;
  assign n603 = n476 & n602 ;
  assign n604 = n601 & ~n603 ;
  assign n605 = ~n600 & ~n604 ;
  assign n606 = ~n571 & ~n573 ;
  assign n607 = n570 & ~n606 ;
  assign n608 = ~n569 & n607 ;
  assign n609 = \g1226_reg/NET0131  & ~\g1229_reg/NET0131  ;
  assign n610 = \g1227_reg/NET0131  & \g1228_reg/NET0131  ;
  assign n611 = \g1230_reg/NET0131  & n610 ;
  assign n612 = n609 & n611 ;
  assign n613 = ~\g1257_reg/NET0131  & ~\g1263_reg/NET0131  ;
  assign n614 = \g1225_reg/NET0131  & n597 ;
  assign n615 = ~n613 & n614 ;
  assign n616 = n612 & n615 ;
  assign n617 = \g1247_reg/NET0131  & ~n616 ;
  assign n618 = \g1253_reg/NET0131  & ~n617 ;
  assign n619 = \g1336_reg/NET0131  & n170 ;
  assign n620 = ~\g1339_reg/NET0131  & ~n619 ;
  assign n621 = \g1247_reg/NET0131  & ~n172 ;
  assign n622 = ~n620 & n621 ;
  assign n623 = ~\g1220_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n624 = ~n476 & n623 ;
  assign n625 = n476 & n598 ;
  assign n626 = ~n624 & ~n625 ;
  assign n627 = ~\g1416_reg/NET0131  & ~\g1421_reg/NET0131  ;
  assign n628 = ~\g1307_reg/NET0131  & ~n627 ;
  assign n629 = \g1247_reg/NET0131  & ~\g1330_reg/NET0131  ;
  assign n630 = \g1247_reg/NET0131  & \g1336_reg/NET0131  ;
  assign n631 = ~n170 & n630 ;
  assign n632 = \g1247_reg/NET0131  & ~\g1336_reg/NET0131  ;
  assign n633 = n170 & n632 ;
  assign n634 = ~n631 & ~n633 ;
  assign n635 = \g1247_reg/NET0131  & \g1342_reg/NET0131  ;
  assign n636 = ~n172 & n635 ;
  assign n637 = \g1247_reg/NET0131  & ~\g1342_reg/NET0131  ;
  assign n638 = n172 & n637 ;
  assign n639 = ~n636 & ~n638 ;
  assign n640 = n421 & n469 ;
  assign n641 = \g104_reg/NET0131  & n640 ;
  assign n642 = ~\g1292_reg/NET0131  & ~\g1296_reg/NET0131  ;
  assign n643 = ~\g1284_reg/NET0131  & ~\g1288_reg/NET0131  ;
  assign n644 = ~\g1276_reg/NET0131  & n643 ;
  assign n645 = ~\g104_reg/NET0131  & ~\g1272_reg/NET0131  ;
  assign n646 = ~\g1280_reg/NET0131  & ~\g1300_reg/NET0131  ;
  assign n647 = n645 & n646 ;
  assign n648 = n644 & n647 ;
  assign n649 = n642 & n648 ;
  assign n650 = ~n641 & ~n649 ;
  assign n651 = \g104_reg/NET0131  & ~n198 ;
  assign n652 = ~n215 & ~n651 ;
  assign n653 = ~\g1268_reg/NET0131  & ~\g1269_reg/NET0131  ;
  assign n654 = \g871_reg/NET0131  & n369 ;
  assign n655 = ~n198 & ~n199 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~\g4372_pad  & ~\g4373_pad  ;
  assign n658 = ~\g4370_pad  & n657 ;
  assign n659 = ~\g1073_reg/NET0131  & ~\g1179_reg/NET0131  ;
  assign n660 = ~\g4371_pad  & n659 ;
  assign n661 = n658 & n660 ;
  assign n662 = \g1225_reg/NET0131  & \g1263_reg/NET0131  ;
  assign n663 = n597 & n662 ;
  assign n664 = n612 & n663 ;
  assign n665 = \g1225_reg/NET0131  & \g1257_reg/NET0131  ;
  assign n666 = n597 & n665 ;
  assign n667 = n612 & n666 ;
  assign n668 = \g1225_reg/NET0131  & \g1266_reg/NET0131  ;
  assign n669 = n597 & n668 ;
  assign n670 = n612 & n669 ;
  assign n671 = \g1207_reg/NET0131  & n474 ;
  assign n672 = ~\g1217_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n673 = ~n671 & n672 ;
  assign n674 = \g1217_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n675 = n671 & n674 ;
  assign n676 = ~n673 & ~n675 ;
  assign n677 = ~\g1229_reg/NET0131  & ~\g1230_reg/NET0131  ;
  assign n678 = ~\g1227_reg/NET0131  & ~\g1228_reg/NET0131  ;
  assign n679 = n677 & n678 ;
  assign n680 = ~\g1225_reg/NET0131  & ~\g1226_reg/NET0131  ;
  assign n681 = ~\g1223_reg/NET0131  & ~\g1224_reg/NET0131  ;
  assign n682 = n680 & n681 ;
  assign n683 = n679 & n682 ;
  assign n684 = \g1207_reg/NET0131  & \g1211_reg/NET0131  ;
  assign n685 = ~\g1207_reg/NET0131  & ~\g1211_reg/NET0131  ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = ~\g1231_reg/NET0131  & ~n686 ;
  assign n688 = ~\g1214_reg/NET0131  & ~n684 ;
  assign n689 = ~\g1231_reg/NET0131  & \g2662_pad  ;
  assign n690 = ~n671 & n689 ;
  assign n691 = ~n688 & n690 ;
  assign n692 = ~\g871_reg/NET0131  & ~n369 ;
  assign n693 = ~n654 & ~n692 ;
  assign n694 = \g1207_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n695 = \g104_reg/NET0131  & ~\g1211_reg/NET0131  ;
  assign n696 = ~\g104_reg/NET0131  & \g1211_reg/NET0131  ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = \g104_reg/NET0131  & ~\g1214_reg/NET0131  ;
  assign n699 = ~\g104_reg/NET0131  & \g1214_reg/NET0131  ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = \g104_reg/NET0131  & ~\g1220_reg/NET0131  ;
  assign n702 = ~\g104_reg/NET0131  & \g1220_reg/NET0131  ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = \g104_reg/NET0131  & ~\g1207_reg/NET0131  ;
  assign n705 = ~\g104_reg/NET0131  & \g1207_reg/NET0131  ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = \g104_reg/NET0131  & ~\g1225_reg/NET0131  ;
  assign n708 = ~\g104_reg/NET0131  & \g1225_reg/NET0131  ;
  assign n709 = ~n707 & ~n708 ;
  assign n710 = \g104_reg/NET0131  & ~\g1227_reg/NET0131  ;
  assign n711 = ~\g104_reg/NET0131  & \g1227_reg/NET0131  ;
  assign n712 = ~n710 & ~n711 ;
  assign n713 = \g104_reg/NET0131  & ~\g1228_reg/NET0131  ;
  assign n714 = ~\g104_reg/NET0131  & \g1228_reg/NET0131  ;
  assign n715 = ~n713 & ~n714 ;
  assign n716 = \g104_reg/NET0131  & ~\g1230_reg/NET0131  ;
  assign n717 = ~\g104_reg/NET0131  & \g1230_reg/NET0131  ;
  assign n718 = ~n716 & ~n717 ;
  assign n719 = \g104_reg/NET0131  & ~\g1223_reg/NET0131  ;
  assign n720 = ~\g104_reg/NET0131  & \g1223_reg/NET0131  ;
  assign n721 = ~n719 & ~n720 ;
  assign n722 = \g104_reg/NET0131  & ~\g1224_reg/NET0131  ;
  assign n723 = ~\g104_reg/NET0131  & \g1224_reg/NET0131  ;
  assign n724 = ~n722 & ~n723 ;
  assign n725 = \g104_reg/NET0131  & ~\g1226_reg/NET0131  ;
  assign n726 = ~\g104_reg/NET0131  & \g1226_reg/NET0131  ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = \g1217_reg/NET0131  & \g1220_reg/NET0131  ;
  assign n729 = ~\g1211_reg/NET0131  & n728 ;
  assign n730 = \g1207_reg/NET0131  & \g1214_reg/NET0131  ;
  assign n731 = n729 & n730 ;
  assign n732 = ~\g1207_reg/NET0131  & \g1214_reg/NET0131  ;
  assign n733 = n729 & n732 ;
  assign n734 = \g1211_reg/NET0131  & n728 ;
  assign n735 = n732 & n734 ;
  assign n736 = \g104_reg/NET0131  & ~\g1217_reg/NET0131  ;
  assign n737 = ~\g104_reg/NET0131  & \g1217_reg/NET0131  ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = \g104_reg/NET0131  & ~\g1229_reg/NET0131  ;
  assign n740 = ~\g104_reg/NET0131  & \g1229_reg/NET0131  ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = ~\g929_reg/NET0131  & ~\g933_reg/NET0131  ;
  assign n743 = ~n369 & ~n742 ;
  assign n744 = ~\g1217_reg/NET0131  & ~\g1220_reg/NET0131  ;
  assign n745 = n474 & n744 ;
  assign n746 = ~\g1454_reg/NET0131  & n538 ;
  assign n747 = \g1454_reg/NET0131  & n536 ;
  assign n748 = \g942_reg/NET0131  & ~n199 ;
  assign n749 = \g1114_reg/NET0131  & \g1118_reg/NET0131  ;
  assign n750 = \g1122_reg/NET0131  & n749 ;
  assign n751 = ~\g1097_reg/NET0131  & n750 ;
  assign n752 = n262 & n751 ;
  assign n753 = n238 & n749 ;
  assign n754 = n237 & n753 ;
  assign n755 = ~\g1097_reg/NET0131  & ~\g1122_reg/NET0131  ;
  assign n756 = ~n754 & n755 ;
  assign n757 = ~n752 & ~n756 ;
  assign n758 = n262 & n750 ;
  assign n759 = ~\g1097_reg/NET0131  & ~\g1126_reg/NET0131  ;
  assign n760 = ~n758 & n759 ;
  assign n761 = ~\g1097_reg/NET0131  & \g1126_reg/NET0131  ;
  assign n762 = n750 & n761 ;
  assign n763 = n262 & n762 ;
  assign n764 = ~n760 & ~n763 ;
  assign n765 = \g1110_reg/NET0131  & \g1126_reg/NET0131  ;
  assign n766 = \g1142_reg/NET0131  & n765 ;
  assign n767 = n750 & n766 ;
  assign n768 = n237 & n767 ;
  assign n769 = ~\g7424_pad  & ~\g7425_pad  ;
  assign n770 = ~\g1166_reg/NET0131  & n769 ;
  assign n771 = ~\g7423_pad  & n770 ;
  assign n772 = ~n768 & n771 ;
  assign n773 = \g1211_reg/NET0131  & \g1226_reg/NET0131  ;
  assign n774 = n728 & n773 ;
  assign n775 = n610 & n730 ;
  assign n776 = n774 & n775 ;
  assign n777 = ~\g1231_reg/NET0131  & n614 ;
  assign n778 = n776 & n777 ;
  assign n779 = \g1226_reg/NET0131  & \g1227_reg/NET0131  ;
  assign n780 = n730 & n779 ;
  assign n781 = n614 & n780 ;
  assign n782 = n734 & n781 ;
  assign n783 = ~\g1228_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n784 = ~n782 & n783 ;
  assign n785 = ~n778 & ~n784 ;
  assign n786 = n614 & n776 ;
  assign n787 = ~\g1229_reg/NET0131  & ~n786 ;
  assign n788 = n614 & n730 ;
  assign n789 = \g1229_reg/NET0131  & n610 ;
  assign n790 = n774 & n789 ;
  assign n791 = n788 & n790 ;
  assign n792 = n689 & ~n791 ;
  assign n793 = ~n787 & n792 ;
  assign n794 = \g1462_reg/NET0131  & n225 ;
  assign n795 = n222 & n794 ;
  assign n796 = ~\g1467_reg/NET0131  & ~n795 ;
  assign n797 = \g1467_reg/NET0131  & n794 ;
  assign n798 = n222 & n797 ;
  assign n799 = ~n229 & ~n798 ;
  assign n800 = ~n796 & n799 ;
  assign n801 = \g1486_reg/NET0131  & ~n229 ;
  assign n802 = ~\g1486_reg/NET0131  & n219 ;
  assign n803 = n228 & n802 ;
  assign n804 = ~n801 & ~n803 ;
  assign n805 = n774 & n788 ;
  assign n806 = ~\g1227_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n807 = ~n805 & n806 ;
  assign n808 = \g1227_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n809 = n774 & n808 ;
  assign n810 = n788 & n809 ;
  assign n811 = ~n807 & ~n810 ;
  assign n812 = ~\g1519_reg/NET0131  & ~n232 ;
  assign n813 = n222 & n225 ;
  assign n814 = ~n229 & ~n813 ;
  assign n815 = ~n812 & n814 ;
  assign n816 = ~\g1462_reg/NET0131  & ~n813 ;
  assign n817 = ~n229 & ~n795 ;
  assign n818 = ~n816 & n817 ;
  assign n819 = n734 & n788 ;
  assign n820 = ~\g1226_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n821 = ~n819 & n820 ;
  assign n822 = \g1226_reg/NET0131  & ~\g1231_reg/NET0131  ;
  assign n823 = n734 & n822 ;
  assign n824 = n788 & n823 ;
  assign n825 = ~n821 & ~n824 ;
  assign n826 = \g1220_reg/NET0131  & n597 ;
  assign n827 = n476 & n826 ;
  assign n828 = \g1225_reg/NET0131  & ~n827 ;
  assign n829 = \g1220_reg/NET0131  & ~\g1225_reg/NET0131  ;
  assign n830 = n597 & n829 ;
  assign n831 = n476 & n830 ;
  assign n832 = ~\g1231_reg/NET0131  & ~n831 ;
  assign n833 = ~n828 & n832 ;
  assign n834 = \g1229_reg/NET0131  & \g1230_reg/NET0131  ;
  assign n835 = n610 & n834 ;
  assign n836 = n774 & n835 ;
  assign n837 = n788 & n836 ;
  assign n838 = ~\g1231_reg/NET0131  & n837 ;
  assign n839 = \g1229_reg/NET0131  & \g2662_pad  ;
  assign n840 = n610 & n839 ;
  assign n841 = n774 & n840 ;
  assign n842 = n788 & n841 ;
  assign n843 = \g1230_reg/NET0131  & \g2662_pad  ;
  assign n844 = ~\g1231_reg/NET0131  & ~n843 ;
  assign n845 = ~n842 & n844 ;
  assign n846 = ~n838 & ~n845 ;
  assign n847 = \g1354_reg/NET0131  & n344 ;
  assign n848 = ~\g1357_reg/NET0131  & ~n847 ;
  assign n849 = n344 & n565 ;
  assign n850 = \g1247_reg/NET0131  & ~n849 ;
  assign n851 = ~n848 & n850 ;
  assign n852 = \g1041_reg/NET0131  & n286 ;
  assign n853 = n183 & n852 ;
  assign n854 = \g1045_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n855 = n193 & n854 ;
  assign n856 = ~n853 & n855 ;
  assign n857 = \g1045_reg/NET0131  & n204 ;
  assign n858 = \g1041_reg/NET0131  & ~\g1045_reg/NET0131  ;
  assign n859 = n286 & n858 ;
  assign n860 = n183 & n859 ;
  assign n861 = n285 & n860 ;
  assign n862 = ~n857 & ~n861 ;
  assign n863 = ~n856 & n862 ;
  assign n864 = \g1065_reg/NET0131  & n204 ;
  assign n865 = n187 & n190 ;
  assign n866 = ~\g1065_reg/NET0131  & ~n865 ;
  assign n867 = ~n192 & n285 ;
  assign n868 = ~n866 & n867 ;
  assign n869 = ~n864 & ~n868 ;
  assign n870 = \g1053_reg/NET0131  & n204 ;
  assign n871 = \g1049_reg/NET0131  & n187 ;
  assign n872 = ~\g1053_reg/NET0131  & ~n871 ;
  assign n873 = n187 & n188 ;
  assign n874 = n285 & ~n873 ;
  assign n875 = ~n872 & n874 ;
  assign n876 = ~n870 & ~n875 ;
  assign n877 = \g1342_reg/NET0131  & n172 ;
  assign n878 = ~\g1345_reg/NET0131  & ~n877 ;
  assign n879 = \g1247_reg/NET0131  & ~n174 ;
  assign n880 = ~n878 & n879 ;
  assign n881 = \g1122_reg/NET0131  & \g1126_reg/NET0131  ;
  assign n882 = n749 & n881 ;
  assign n883 = n262 & n882 ;
  assign n884 = ~\g1142_reg/NET0131  & ~n883 ;
  assign n885 = \g1122_reg/NET0131  & \g1142_reg/NET0131  ;
  assign n886 = n749 & n885 ;
  assign n887 = \g1126_reg/NET0131  & n886 ;
  assign n888 = n262 & n887 ;
  assign n889 = ~\g1097_reg/NET0131  & ~n888 ;
  assign n890 = ~n884 & n889 ;
  assign n891 = n192 & n285 ;
  assign n892 = ~\g1069_reg/NET0131  & ~n891 ;
  assign n893 = \g1069_reg/NET0131  & ~n204 ;
  assign n894 = ~n867 & n893 ;
  assign n895 = ~n892 & ~n894 ;
  assign n896 = \g1049_reg/NET0131  & \g1057_reg/NET0131  ;
  assign n897 = \g1053_reg/NET0131  & n896 ;
  assign n898 = n187 & n897 ;
  assign n899 = \g1061_reg/NET0131  & n285 ;
  assign n900 = ~n898 & n899 ;
  assign n901 = \g1061_reg/NET0131  & n204 ;
  assign n902 = \g1057_reg/NET0131  & ~\g1061_reg/NET0131  ;
  assign n903 = n188 & n902 ;
  assign n904 = n285 & n903 ;
  assign n905 = n187 & n904 ;
  assign n906 = ~n901 & ~n905 ;
  assign n907 = ~n900 & n906 ;
  assign n908 = n344 & n566 ;
  assign n909 = \g1247_reg/NET0131  & \g1360_reg/NET0131  ;
  assign n910 = \g1247_reg/NET0131  & n565 ;
  assign n911 = n344 & n910 ;
  assign n912 = ~n909 & ~n911 ;
  assign n913 = ~n908 & ~n912 ;
  assign n914 = n188 & n285 ;
  assign n915 = n187 & n914 ;
  assign n916 = ~\g1057_reg/NET0131  & ~n915 ;
  assign n917 = \g1057_reg/NET0131  & ~n204 ;
  assign n918 = ~n874 & n917 ;
  assign n919 = ~n916 & ~n918 ;
  assign n920 = ~\g1328_reg/NET0131  & ~n514 ;
  assign n921 = ~\g1329_reg/NET0131  & ~n366 ;
  assign n922 = ~n920 & n921 ;
  assign n923 = ~n337 & ~n922 ;
  assign n924 = \g1041_reg/NET0131  & n204 ;
  assign n925 = \g1041_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n926 = n193 & n925 ;
  assign n927 = ~n287 & n926 ;
  assign n928 = ~n924 & ~n927 ;
  assign n929 = ~\g1041_reg/NET0131  & ~\g1251_reg/NET0131  ;
  assign n930 = n193 & n929 ;
  assign n931 = n287 & n930 ;
  assign n932 = n928 & ~n931 ;
  assign n933 = ~\g1472_reg/NET0131  & ~n798 ;
  assign n934 = \g1467_reg/NET0131  & \g1472_reg/NET0131  ;
  assign n935 = n794 & n934 ;
  assign n936 = n222 & n935 ;
  assign n937 = ~n229 & ~n936 ;
  assign n938 = ~n933 & n937 ;
  assign n939 = ~\g2_reg/NET0131  & ~\g962_pad  ;
  assign n940 = ~\g1189_reg/NET0131  & ~\g7505_pad  ;
  assign n941 = \g1405_reg/NET0131  & \g1412_reg/NET0131  ;
  assign \g1006_pad  = 1'b0 ;
  assign \g1158_reg/P0001  = ~\g1158_reg/NET0131  ;
  assign \g1252_reg/P0001  = ~\g1252_reg/NET0131  ;
  assign \g1260_reg/P0001  = ~\g1260_reg/NET0131  ;
  assign \g1416_reg/NET0131_syn_2  = ~\g1416_reg/NET0131  ;
  assign \g17/_0_  = n179 ;
  assign \g19189/_0_  = ~n197 ;
  assign \g19252/_0_  = ~n201 ;
  assign \g19253/_0_  = ~n213 ;
  assign \g19273/_3_  = ~n216 ;
  assign \g19284/_0_  = n234 ;
  assign \g19285/_0_  = n247 ;
  assign \g19295/_3_  = ~n249 ;
  assign \g19302/_0_  = ~n255 ;
  assign \g19303/_0_  = n261 ;
  assign \g19304/_0_  = n265 ;
  assign \g19308/_0_  = n269 ;
  assign \g19309/_0_  = ~n276 ;
  assign \g19310/_0_  = n281 ;
  assign \g19321/_0_  = ~n290 ;
  assign \g19326/_3_  = ~n292 ;
  assign \g19331/_0_  = n296 ;
  assign \g19341/_0_  = n300 ;
  assign \g19366/_0_  = ~n309 ;
  assign \g19372/_3_  = ~n311 ;
  assign \g19385/_0_  = n315 ;
  assign \g19386/_0_  = ~n323 ;
  assign \g19387/_0_  = n325 ;
  assign \g19388/_0_  = n328 ;
  assign \g19389/_0_  = ~n341 ;
  assign \g19390/_0_  = ~n349 ;
  assign \g19392/_0_  = n361 ;
  assign \g19393/_0_  = n368 ;
  assign \g19394/_0_  = n372 ;
  assign \g19398/_0_  = ~n381 ;
  assign \g19399/_0_  = ~n387 ;
  assign \g19400/_0_  = n395 ;
  assign \g19401/_0_  = ~n400 ;
  assign \g19403/_0_  = ~n405 ;
  assign \g19405/_0_  = n408 ;
  assign \g19406/_0_  = n411 ;
  assign \g19437/_0_  = n418 ;
  assign \g19438/_0_  = n428 ;
  assign \g19445/_0_  = n435 ;
  assign \g19446/_0_  = ~n441 ;
  assign \g19450/_3_  = ~n446 ;
  assign \g19472/_0_  = ~n449 ;
  assign \g19473/_0_  = n454 ;
  assign \g19474/_0_  = n459 ;
  assign \g19476/_0_  = n461 ;
  assign \g19484/_0_  = n465 ;
  assign \g19485/_0_  = n473 ;
  assign \g19492/_0_  = n483 ;
  assign \g19493/_0_  = n486 ;
  assign \g19499/_0_  = ~n488 ;
  assign \g19500/_0_  = ~n494 ;
  assign \g19501/_0_  = ~n498 ;
  assign \g19502/_0_  = ~n503 ;
  assign \g19503/_0_  = ~n508 ;
  assign \g19504/_0_  = ~n517 ;
  assign \g19507/_3_  = n519 ;
  assign \g19508/_3_  = n521 ;
  assign \g19512/_3_  = ~n525 ;
  assign \g19513/_3_  = ~n527 ;
  assign \g19514/_3_  = ~n532 ;
  assign \g19528/_0_  = ~n535 ;
  assign \g19529/_0_  = ~n541 ;
  assign \g19534/_0_  = ~n542 ;
  assign \g19535/_0_  = ~n543 ;
  assign \g19536/_0_  = n545 ;
  assign \g19538/_0_  = n549 ;
  assign \g19542/_0_  = ~n555 ;
  assign \g19560/_0_  = ~n576 ;
  assign \g19563/_0_  = ~n580 ;
  assign \g19565/_0_  = n582 ;
  assign \g19567/_0_  = n585 ;
  assign \g19569/_1_  = n587 ;
  assign \g19572/_0_  = n593 ;
  assign \g19574/_3_  = ~n596 ;
  assign \g19614/_0_  = n605 ;
  assign \g19615/_0_  = ~n608 ;
  assign \g19620/_0_  = ~n618 ;
  assign \g19626/_0_  = n622 ;
  assign \g19629/_0_  = n626 ;
  assign \g19631/_0_  = ~n628 ;
  assign \g19666/_0_  = n629 ;
  assign \g19667/_0_  = ~n634 ;
  assign \g19669/_0_  = ~n639 ;
  assign \g19677/_0_  = n650 ;
  assign \g19690/_3_  = ~n652 ;
  assign \g19721/_0_  = n653 ;
  assign \g19723/_0_  = n656 ;
  assign \g19723/_1_  = n654 ;
  assign \g19725/_2_  = ~n661 ;
  assign \g19751/_0_  = ~n664 ;
  assign \g19752/_0_  = ~n667 ;
  assign \g19753/_0_  = ~n670 ;
  assign \g19755/_0_  = n676 ;
  assign \g19815/_0_  = ~n683 ;
  assign \g19821/_0_  = ~n687 ;
  assign \g19822/_0_  = n691 ;
  assign \g19833/_0_  = n693 ;
  assign \g19877/_0_  = ~n694 ;
  assign \g19898/_0_  = ~n697 ;
  assign \g19899/_0_  = ~n700 ;
  assign \g19900/_0_  = ~n703 ;
  assign \g19901/_0_  = ~n706 ;
  assign \g19908/_0_  = ~n709 ;
  assign \g19927/_0_  = ~n712 ;
  assign \g19928/_0_  = ~n715 ;
  assign \g19930/_0_  = ~n718 ;
  assign \g19931/_0_  = ~n721 ;
  assign \g19932/_0_  = ~n724 ;
  assign \g19934/_0_  = ~n727 ;
  assign \g19992/_0_  = n731 ;
  assign \g19993/_0_  = n733 ;
  assign \g20002/_0_  = n735 ;
  assign \g20008/_0_  = ~n738 ;
  assign \g20010/_0_  = ~n741 ;
  assign \g20016/_0_  = n743 ;
  assign \g20110/_0_  = ~n745 ;
  assign \g20117/_0_  = n746 ;
  assign \g20118/_0_  = n747 ;
  assign \g20131/_0_  = n748 ;
  assign \g20246/_0_  = ~\g929_reg/NET0131  ;
  assign \g20704/_0_  = n757 ;
  assign \g20722/_0_  = n764 ;
  assign \g20731/_0_  = ~n772 ;
  assign \g20732/_2_  = n768 ;
  assign \g20870/_0_  = n785 ;
  assign \g20883/_0_  = n793 ;
  assign \g20931/_0_  = n800 ;
  assign \g20951/_0_  = ~n804 ;
  assign \g20969/_0_  = n811 ;
  assign \g20989/_0_  = n617 ;
  assign \g21/_2_  = n815 ;
  assign \g21070/_0_  = n818 ;
  assign \g21108/_0_  = n825 ;
  assign \g21122/_0_  = ~n833 ;
  assign \g21152/_0_  = n846 ;
  assign \g21191/_0_  = n851 ;
  assign \g21279/_0_  = ~n863 ;
  assign \g21316/_0_  = ~n869 ;
  assign \g21323/_0_  = ~n876 ;
  assign \g21349/_3_  = n640 ;
  assign \g21352/_3_  = n880 ;
  assign \g21464/_0_  = n890 ;
  assign \g21472/_0_  = n895 ;
  assign \g21484/_0_  = ~n907 ;
  assign \g21510/_0_  = n913 ;
  assign \g21517/_0_  = n919 ;
  assign \g21608/_0_  = ~n923 ;
  assign \g21625/_0_  = ~n932 ;
  assign \g21644/_1_  = n938 ;
  assign \g4655_pad  = ~n655 ;
  assign \g6850_pad  = ~\g43_pad  ;
  assign \g6895_pad  = ~1'b0 ;
  assign \g7048_pad  = ~\g944_reg/NET0131  ;
  assign \g7103_pad  = ~n939 ;
  assign \g7731_pad  = ~n940 ;
  assign \g7732_pad  = ~\g1486_reg/NET0131  ;
  assign \g8219_pad  = ~\g1432_reg/NET0131  ;
  assign \g8663_pad  = ~n941 ;
endmodule
