module top( \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G14_pad  , \G15_pad  , \G16_pad  , \G18_pad  , \G19_pad  , \G20_pad  , \G22_pad  , \G23_pad  , \G24_pad  , \G25_pad  , \G26_pad  , \G28_pad  , \G2_pad  , \G30_pad  , \G31_pad  , \G32_pad  , \G33_pad  , \G34_pad  , \G35_pad  , \G3_pad  , \G4_pad  , \G5_pad  , \G64_reg/NET0131  , \G65_reg/NET0131  , \G66_reg/NET0131  , \G69_reg/NET0131  , \G6_pad  , \G70_reg/NET0131  , \G71_reg/NET0131  , \G72_reg/NET0131  , \G73_reg/NET0131  , \G74_reg/NET0131  , \G75_reg/NET0131  , \G76_reg/NET0131  , \G77_reg/NET0131  , \G79_reg/NET0131  , \G81_reg/NET0131  , \G8_pad  , \G9_pad  , \G100BF_pad  , \G103BF_pad  , \G104BF_pad  , \G105BF_pad  , \G107_pad  , \G83_pad  , \G84_pad  , \G86BF_pad  , \G89BF_pad  , \G95BF_pad  , \G96BF_pad  , \G97BF_pad  , \G98BF_pad  , \G99BF_pad  , \_al_n0  , \_al_n1  , \g1017/_3_  , \g1150/_0_  , \g1168/_0_  , \g1308/_1_  , \g1318/_0_  , \g1337/_2_  , \g1339/_1_  , \g16/_0_  , \g26/_2_  , \g27/_0_  , \g29/_0_  , \g867/_3_  , \g875/_0_  , \g898/_0_  , \g931/_0_  , \g938/_0_  , \g967/_0_  , \g987/_0_  );
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G14_pad  ;
  input \G15_pad  ;
  input \G16_pad  ;
  input \G18_pad  ;
  input \G19_pad  ;
  input \G20_pad  ;
  input \G22_pad  ;
  input \G23_pad  ;
  input \G24_pad  ;
  input \G25_pad  ;
  input \G26_pad  ;
  input \G28_pad  ;
  input \G2_pad  ;
  input \G30_pad  ;
  input \G31_pad  ;
  input \G32_pad  ;
  input \G33_pad  ;
  input \G34_pad  ;
  input \G35_pad  ;
  input \G3_pad  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G64_reg/NET0131  ;
  input \G65_reg/NET0131  ;
  input \G66_reg/NET0131  ;
  input \G69_reg/NET0131  ;
  input \G6_pad  ;
  input \G70_reg/NET0131  ;
  input \G71_reg/NET0131  ;
  input \G72_reg/NET0131  ;
  input \G73_reg/NET0131  ;
  input \G74_reg/NET0131  ;
  input \G75_reg/NET0131  ;
  input \G76_reg/NET0131  ;
  input \G77_reg/NET0131  ;
  input \G79_reg/NET0131  ;
  input \G81_reg/NET0131  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G100BF_pad  ;
  output \G103BF_pad  ;
  output \G104BF_pad  ;
  output \G105BF_pad  ;
  output \G107_pad  ;
  output \G83_pad  ;
  output \G84_pad  ;
  output \G86BF_pad  ;
  output \G89BF_pad  ;
  output \G95BF_pad  ;
  output \G96BF_pad  ;
  output \G97BF_pad  ;
  output \G98BF_pad  ;
  output \G99BF_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1017/_3_  ;
  output \g1150/_0_  ;
  output \g1168/_0_  ;
  output \g1308/_1_  ;
  output \g1318/_0_  ;
  output \g1337/_2_  ;
  output \g1339/_1_  ;
  output \g16/_0_  ;
  output \g26/_2_  ;
  output \g27/_0_  ;
  output \g29/_0_  ;
  output \g867/_3_  ;
  output \g875/_0_  ;
  output \g898/_0_  ;
  output \g931/_0_  ;
  output \g938/_0_  ;
  output \g967/_0_  ;
  output \g987/_0_  ;
  wire n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 ;
  assign n44 = ~\G4_pad  & \G69_reg/NET0131  ;
  assign n45 = \G35_pad  & n44 ;
  assign n46 = \G3_pad  & \G75_reg/NET0131  ;
  assign n47 = \G14_pad  & n46 ;
  assign n48 = \G3_pad  & \G77_reg/NET0131  ;
  assign n49 = ~\G11_pad  & ~\G3_pad  ;
  assign n50 = ~\G2_pad  & \G66_reg/NET0131  ;
  assign n51 = \G24_pad  & ~n50 ;
  assign n52 = ~n49 & n51 ;
  assign n53 = ~\G10_pad  & ~\G13_pad  ;
  assign n54 = ~\G3_pad  & \G9_pad  ;
  assign n55 = n53 & n54 ;
  assign n56 = \G77_reg/NET0131  & ~n55 ;
  assign n57 = n52 & n56 ;
  assign n58 = ~n48 & ~n57 ;
  assign n59 = ~\G2_pad  & \G64_reg/NET0131  ;
  assign n60 = ~\G76_reg/NET0131  & n59 ;
  assign n61 = ~\G13_pad  & ~\G3_pad  ;
  assign n62 = \G10_pad  & ~\G9_pad  ;
  assign n63 = n61 & n62 ;
  assign n64 = \G23_pad  & ~\G65_reg/NET0131  ;
  assign n65 = ~n49 & n64 ;
  assign n66 = ~n63 & n65 ;
  assign n67 = ~\G3_pad  & n59 ;
  assign n68 = ~n66 & n67 ;
  assign n69 = ~n60 & ~n68 ;
  assign n70 = n58 & ~n69 ;
  assign n71 = ~\G10_pad  & ~\G9_pad  ;
  assign n72 = n61 & n71 ;
  assign n73 = \G22_pad  & \G75_reg/NET0131  ;
  assign n74 = ~n49 & n73 ;
  assign n75 = ~n72 & n74 ;
  assign n76 = \G14_pad  & n75 ;
  assign n77 = ~n70 & n76 ;
  assign n78 = ~n47 & ~n77 ;
  assign n79 = ~\G3_pad  & ~n66 ;
  assign n80 = \G15_pad  & \G76_reg/NET0131  ;
  assign n81 = ~n79 & n80 ;
  assign n82 = \G16_pad  & ~n58 ;
  assign n83 = \G18_pad  & ~\G4_pad  ;
  assign n84 = \G79_reg/NET0131  & n83 ;
  assign n85 = \G19_pad  & ~\G4_pad  ;
  assign n86 = \G65_reg/NET0131  & n85 ;
  assign n87 = \G20_pad  & ~\G4_pad  ;
  assign n88 = \G81_reg/NET0131  & n87 ;
  assign n89 = \G22_pad  & ~n49 ;
  assign n90 = ~n72 & n89 ;
  assign n91 = ~n70 & n90 ;
  assign n92 = \G10_pad  & \G9_pad  ;
  assign n93 = n61 & n92 ;
  assign n94 = \G25_pad  & ~n49 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = \G30_pad  & \G74_reg/NET0131  ;
  assign n97 = n90 & n96 ;
  assign n98 = ~n70 & n97 ;
  assign n99 = ~\G4_pad  & \G73_reg/NET0131  ;
  assign n100 = \G31_pad  & n99 ;
  assign n101 = \G32_pad  & \G72_reg/NET0131  ;
  assign n102 = n66 & n101 ;
  assign n103 = ~\G4_pad  & \G71_reg/NET0131  ;
  assign n104 = \G33_pad  & n103 ;
  assign n105 = \G34_pad  & \G70_reg/NET0131  ;
  assign n106 = ~n55 & n105 ;
  assign n107 = n52 & n106 ;
  assign n108 = \G13_pad  & \G28_pad  ;
  assign n109 = \G11_pad  & \G12_pad  ;
  assign n110 = n108 & n109 ;
  assign n111 = \G22_pad  & \G74_reg/NET0131  ;
  assign n112 = ~n49 & n111 ;
  assign n113 = ~n72 & n112 ;
  assign n114 = ~n70 & n113 ;
  assign n115 = n99 & ~n114 ;
  assign n116 = \G2_pad  & ~\G5_pad  ;
  assign n117 = \G76_reg/NET0131  & ~n116 ;
  assign n118 = ~n79 & n117 ;
  assign n119 = ~n70 & n75 ;
  assign n120 = \G5_pad  & \G72_reg/NET0131  ;
  assign n121 = n103 & n120 ;
  assign n122 = n66 & n121 ;
  assign n123 = n58 & n122 ;
  assign n124 = ~n46 & n123 ;
  assign n125 = ~n119 & n124 ;
  assign n126 = ~n118 & ~n125 ;
  assign n127 = ~n46 & ~n119 ;
  assign n128 = n52 & ~n55 ;
  assign n129 = ~\G2_pad  & ~n58 ;
  assign n130 = ~\G2_pad  & \G76_reg/NET0131  ;
  assign n131 = ~n79 & n130 ;
  assign n132 = n58 & n131 ;
  assign n133 = ~\G2_pad  & ~\G76_reg/NET0131  ;
  assign n134 = ~\G2_pad  & ~\G3_pad  ;
  assign n135 = ~n66 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = n46 & ~n136 ;
  assign n138 = n75 & ~n136 ;
  assign n139 = ~n70 & n138 ;
  assign n140 = ~n137 & ~n139 ;
  assign n141 = n58 & ~n140 ;
  assign n142 = \G2_pad  & ~\G8_pad  ;
  assign n143 = n46 & ~n142 ;
  assign n144 = n75 & ~n142 ;
  assign n145 = ~n70 & n144 ;
  assign n146 = ~n143 & ~n145 ;
  assign n147 = n58 & n113 ;
  assign n148 = ~\G76_reg/NET0131  & \G8_pad  ;
  assign n149 = n99 & n148 ;
  assign n150 = ~\G3_pad  & \G8_pad  ;
  assign n151 = n99 & n150 ;
  assign n152 = ~n66 & n151 ;
  assign n153 = ~n149 & ~n152 ;
  assign n154 = n69 & ~n153 ;
  assign n155 = n147 & n154 ;
  assign n156 = n146 & ~n155 ;
  assign n157 = ~\G13_pad  & \G72_reg/NET0131  ;
  assign n158 = n62 & n157 ;
  assign n159 = n103 & n158 ;
  assign n160 = n66 & n159 ;
  assign n161 = \G12_pad  & \G26_pad  ;
  assign n162 = ~n160 & n161 ;
  assign n163 = \G70_reg/NET0131  & ~n55 ;
  assign n164 = n44 & ~n49 ;
  assign n165 = n51 & n164 ;
  assign n166 = n163 & n165 ;
  assign n167 = \G9_pad  & n166 ;
  assign n168 = n53 & n167 ;
  assign n169 = \G74_reg/NET0131  & ~\G9_pad  ;
  assign n170 = n99 & n169 ;
  assign n171 = n90 & n170 ;
  assign n172 = n53 & n171 ;
  assign n173 = ~n70 & n172 ;
  assign n174 = ~n168 & ~n173 ;
  assign n175 = n162 & n174 ;
  assign n176 = \G2_pad  & ~\G6_pad  ;
  assign n177 = ~n58 & ~n176 ;
  assign n178 = \G6_pad  & ~\G76_reg/NET0131  ;
  assign n179 = ~\G3_pad  & \G6_pad  ;
  assign n180 = ~n66 & n179 ;
  assign n181 = ~n178 & ~n180 ;
  assign n182 = n166 & ~n181 ;
  assign n183 = ~n46 & n182 ;
  assign n184 = ~n119 & n183 ;
  assign n185 = ~n177 & ~n184 ;
  assign n186 = ~n91 & n99 ;
  assign n187 = ~n114 & ~n186 ;
  assign n188 = n52 & n163 ;
  assign n189 = n44 & ~n188 ;
  assign n190 = n44 & ~n128 ;
  assign n191 = ~n188 & ~n190 ;
  assign n192 = \G72_reg/NET0131  & n66 ;
  assign n193 = n103 & ~n192 ;
  assign n194 = ~n66 & n103 ;
  assign n195 = ~n192 & ~n194 ;
  assign \G100BF_pad  = ~n45 ;
  assign \G103BF_pad  = n78 ;
  assign \G104BF_pad  = ~n81 ;
  assign \G105BF_pad  = ~n82 ;
  assign \G107_pad  = n84 ;
  assign \G83_pad  = n86 ;
  assign \G84_pad  = n88 ;
  assign \G86BF_pad  = ~n91 ;
  assign \G89BF_pad  = ~n95 ;
  assign \G95BF_pad  = ~n98 ;
  assign \G96BF_pad  = ~n100 ;
  assign \G97BF_pad  = ~n102 ;
  assign \G98BF_pad  = ~n104 ;
  assign \G99BF_pad  = ~n107 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1017/_3_  = n110 ;
  assign \g1150/_0_  = ~n115 ;
  assign \g1168/_0_  = ~n126 ;
  assign \g1308/_1_  = ~n127 ;
  assign \g1318/_0_  = ~n128 ;
  assign \g1337/_2_  = n129 ;
  assign \g1339/_1_  = ~n58 ;
  assign \g16/_0_  = n132 ;
  assign \g26/_2_  = n141 ;
  assign \g27/_0_  = ~n156 ;
  assign \g29/_0_  = ~n66 ;
  assign \g867/_3_  = n175 ;
  assign \g875/_0_  = ~n185 ;
  assign \g898/_0_  = ~n187 ;
  assign \g931/_0_  = ~n189 ;
  assign \g938/_0_  = ~n191 ;
  assign \g967/_0_  = ~n193 ;
  assign \g987/_0_  = ~n195 ;
endmodule
