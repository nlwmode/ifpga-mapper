module top (\configuration_cache_line_size_reg_reg[0]/NET0131 , \configuration_cache_line_size_reg_reg[1]/NET0131 , \configuration_cache_line_size_reg_reg[2]/NET0131 , \configuration_cache_line_size_reg_reg[3]/NET0131 , \configuration_cache_line_size_reg_reg[4]/NET0131 , \configuration_cache_line_size_reg_reg[5]/NET0131 , \configuration_cache_line_size_reg_reg[6]/NET0131 , \configuration_cache_line_size_reg_reg[7]/NET0131 , \configuration_command_bit2_0_reg[0]/NET0131 , \configuration_command_bit2_0_reg[1]/NET0131 , \configuration_command_bit2_0_reg[2]/NET0131 , \configuration_command_bit6_reg/NET0131 , \configuration_command_bit8_reg/NET0131 , \configuration_icr_bit2_0_reg[0]/NET0131 , \configuration_icr_bit2_0_reg[1]/NET0131 , \configuration_icr_bit2_0_reg[2]/NET0131 , \configuration_icr_bit31_reg/NET0131 , \configuration_init_complete_reg/NET0131 , \configuration_interrupt_line_reg[0]/NET0131 , \configuration_interrupt_line_reg[1]/NET0131 , \configuration_interrupt_line_reg[2]/NET0131 , \configuration_interrupt_line_reg[3]/NET0131 , \configuration_interrupt_line_reg[4]/NET0131 , \configuration_interrupt_line_reg[5]/NET0131 , \configuration_interrupt_line_reg[6]/NET0131 , \configuration_interrupt_line_reg[7]/NET0131 , \configuration_interrupt_out_reg/NET0131 , \configuration_isr_bit2_0_reg[0]/NET0131 , \configuration_isr_bit2_0_reg[1]/NET0131 , \configuration_isr_bit2_0_reg[2]/NET0131 , \configuration_latency_timer_reg[0]/NET0131 , \configuration_latency_timer_reg[1]/NET0131 , \configuration_latency_timer_reg[2]/NET0131 , \configuration_latency_timer_reg[3]/NET0131 , \configuration_latency_timer_reg[4]/NET0131 , \configuration_latency_timer_reg[5]/NET0131 , \configuration_latency_timer_reg[6]/NET0131 , \configuration_latency_timer_reg[7]/NET0131 , \configuration_pci_am1_reg[10]/NET0131 , \configuration_pci_am1_reg[11]/NET0131 , \configuration_pci_am1_reg[12]/NET0131 , \configuration_pci_am1_reg[13]/NET0131 , \configuration_pci_am1_reg[14]/NET0131 , \configuration_pci_am1_reg[15]/NET0131 , \configuration_pci_am1_reg[16]/NET0131 , \configuration_pci_am1_reg[17]/NET0131 , \configuration_pci_am1_reg[18]/NET0131 , \configuration_pci_am1_reg[19]/NET0131 , \configuration_pci_am1_reg[20]/NET0131 , \configuration_pci_am1_reg[21]/NET0131 , \configuration_pci_am1_reg[22]/NET0131 , \configuration_pci_am1_reg[23]/NET0131 , \configuration_pci_am1_reg[24]/NET0131 , \configuration_pci_am1_reg[25]/NET0131 , \configuration_pci_am1_reg[26]/NET0131 , \configuration_pci_am1_reg[27]/NET0131 , \configuration_pci_am1_reg[28]/NET0131 , \configuration_pci_am1_reg[29]/NET0131 , \configuration_pci_am1_reg[30]/NET0131 , \configuration_pci_am1_reg[31]/NET0131 , \configuration_pci_am1_reg[8]/NET0131 , \configuration_pci_am1_reg[9]/NET0131 , \configuration_pci_ba0_bit31_8_reg[12]/NET0131 , \configuration_pci_ba0_bit31_8_reg[13]/NET0131 , \configuration_pci_ba0_bit31_8_reg[14]/NET0131 , \configuration_pci_ba0_bit31_8_reg[15]/NET0131 , \configuration_pci_ba0_bit31_8_reg[16]/NET0131 , \configuration_pci_ba0_bit31_8_reg[17]/NET0131 , \configuration_pci_ba0_bit31_8_reg[18]/NET0131 , \configuration_pci_ba0_bit31_8_reg[19]/NET0131 , \configuration_pci_ba0_bit31_8_reg[20]/NET0131 , \configuration_pci_ba0_bit31_8_reg[21]/NET0131 , \configuration_pci_ba0_bit31_8_reg[22]/NET0131 , \configuration_pci_ba0_bit31_8_reg[23]/NET0131 , \configuration_pci_ba0_bit31_8_reg[24]/NET0131 , \configuration_pci_ba0_bit31_8_reg[25]/NET0131 , \configuration_pci_ba0_bit31_8_reg[26]/NET0131 , \configuration_pci_ba0_bit31_8_reg[27]/NET0131 , \configuration_pci_ba0_bit31_8_reg[28]/NET0131 , \configuration_pci_ba0_bit31_8_reg[29]/NET0131 , \configuration_pci_ba0_bit31_8_reg[30]/NET0131 , \configuration_pci_ba0_bit31_8_reg[31]/NET0131 , \configuration_pci_ba1_bit31_8_reg[10]/NET0131 , \configuration_pci_ba1_bit31_8_reg[11]/NET0131 , \configuration_pci_ba1_bit31_8_reg[12]/NET0131 , \configuration_pci_ba1_bit31_8_reg[13]/NET0131 , \configuration_pci_ba1_bit31_8_reg[14]/NET0131 , \configuration_pci_ba1_bit31_8_reg[15]/NET0131 , \configuration_pci_ba1_bit31_8_reg[16]/NET0131 , \configuration_pci_ba1_bit31_8_reg[17]/NET0131 , \configuration_pci_ba1_bit31_8_reg[18]/NET0131 , \configuration_pci_ba1_bit31_8_reg[19]/NET0131 , \configuration_pci_ba1_bit31_8_reg[20]/NET0131 , \configuration_pci_ba1_bit31_8_reg[21]/NET0131 , \configuration_pci_ba1_bit31_8_reg[22]/NET0131 , \configuration_pci_ba1_bit31_8_reg[23]/NET0131 , \configuration_pci_ba1_bit31_8_reg[24]/NET0131 , \configuration_pci_ba1_bit31_8_reg[25]/NET0131 , \configuration_pci_ba1_bit31_8_reg[26]/NET0131 , \configuration_pci_ba1_bit31_8_reg[27]/NET0131 , \configuration_pci_ba1_bit31_8_reg[28]/NET0131 , \configuration_pci_ba1_bit31_8_reg[29]/NET0131 , \configuration_pci_ba1_bit31_8_reg[30]/NET0131 , \configuration_pci_ba1_bit31_8_reg[31]/NET0131 , \configuration_pci_ba1_bit31_8_reg[8]/NET0131 , \configuration_pci_ba1_bit31_8_reg[9]/NET0131 , \configuration_pci_err_addr_reg[0]/NET0131 , \configuration_pci_err_addr_reg[10]/NET0131 , \configuration_pci_err_addr_reg[11]/NET0131 , \configuration_pci_err_addr_reg[12]/NET0131 , \configuration_pci_err_addr_reg[13]/NET0131 , \configuration_pci_err_addr_reg[14]/NET0131 , \configuration_pci_err_addr_reg[15]/NET0131 , \configuration_pci_err_addr_reg[16]/NET0131 , \configuration_pci_err_addr_reg[17]/NET0131 , \configuration_pci_err_addr_reg[18]/NET0131 , \configuration_pci_err_addr_reg[19]/NET0131 , \configuration_pci_err_addr_reg[1]/NET0131 , \configuration_pci_err_addr_reg[20]/NET0131 , \configuration_pci_err_addr_reg[21]/NET0131 , \configuration_pci_err_addr_reg[22]/NET0131 , \configuration_pci_err_addr_reg[23]/NET0131 , \configuration_pci_err_addr_reg[24]/NET0131 , \configuration_pci_err_addr_reg[25]/NET0131 , \configuration_pci_err_addr_reg[26]/NET0131 , \configuration_pci_err_addr_reg[27]/NET0131 , \configuration_pci_err_addr_reg[28]/NET0131 , \configuration_pci_err_addr_reg[29]/NET0131 , \configuration_pci_err_addr_reg[2]/NET0131 , \configuration_pci_err_addr_reg[30]/NET0131 , \configuration_pci_err_addr_reg[31]/NET0131 , \configuration_pci_err_addr_reg[3]/NET0131 , \configuration_pci_err_addr_reg[4]/NET0131 , \configuration_pci_err_addr_reg[5]/NET0131 , \configuration_pci_err_addr_reg[6]/NET0131 , \configuration_pci_err_addr_reg[7]/NET0131 , \configuration_pci_err_addr_reg[8]/NET0131 , \configuration_pci_err_addr_reg[9]/NET0131 , \configuration_pci_err_cs_bit0_reg/NET0131 , \configuration_pci_err_cs_bit10_reg/NET0131 , \configuration_pci_err_cs_bit31_24_reg[24]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[25]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[26]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[27]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[28]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[29]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[30]/NET0131 , \configuration_pci_err_cs_bit31_24_reg[31]/NET0131 , \configuration_pci_err_cs_bit8_reg/NET0131 , \configuration_pci_err_data_reg[0]/NET0131 , \configuration_pci_err_data_reg[10]/NET0131 , \configuration_pci_err_data_reg[11]/NET0131 , \configuration_pci_err_data_reg[12]/NET0131 , \configuration_pci_err_data_reg[13]/NET0131 , \configuration_pci_err_data_reg[14]/NET0131 , \configuration_pci_err_data_reg[15]/NET0131 , \configuration_pci_err_data_reg[16]/NET0131 , \configuration_pci_err_data_reg[17]/NET0131 , \configuration_pci_err_data_reg[18]/NET0131 , \configuration_pci_err_data_reg[19]/NET0131 , \configuration_pci_err_data_reg[1]/NET0131 , \configuration_pci_err_data_reg[20]/NET0131 , \configuration_pci_err_data_reg[21]/NET0131 , \configuration_pci_err_data_reg[22]/NET0131 , \configuration_pci_err_data_reg[23]/NET0131 , \configuration_pci_err_data_reg[24]/NET0131 , \configuration_pci_err_data_reg[25]/NET0131 , \configuration_pci_err_data_reg[26]/NET0131 , \configuration_pci_err_data_reg[27]/NET0131 , \configuration_pci_err_data_reg[28]/NET0131 , \configuration_pci_err_data_reg[29]/NET0131 , \configuration_pci_err_data_reg[2]/NET0131 , \configuration_pci_err_data_reg[30]/NET0131 , \configuration_pci_err_data_reg[31]/NET0131 , \configuration_pci_err_data_reg[3]/NET0131 , \configuration_pci_err_data_reg[4]/NET0131 , \configuration_pci_err_data_reg[5]/NET0131 , \configuration_pci_err_data_reg[6]/NET0131 , \configuration_pci_err_data_reg[7]/NET0131 , \configuration_pci_err_data_reg[8]/NET0131 , \configuration_pci_err_data_reg[9]/NET0131 , \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131 , \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131 , \configuration_pci_ta1_reg[10]/NET0131 , \configuration_pci_ta1_reg[11]/NET0131 , \configuration_pci_ta1_reg[12]/NET0131 , \configuration_pci_ta1_reg[13]/NET0131 , \configuration_pci_ta1_reg[14]/NET0131 , \configuration_pci_ta1_reg[15]/NET0131 , \configuration_pci_ta1_reg[16]/NET0131 , \configuration_pci_ta1_reg[17]/NET0131 , \configuration_pci_ta1_reg[18]/NET0131 , \configuration_pci_ta1_reg[19]/NET0131 , \configuration_pci_ta1_reg[20]/NET0131 , \configuration_pci_ta1_reg[21]/NET0131 , \configuration_pci_ta1_reg[22]/NET0131 , \configuration_pci_ta1_reg[23]/NET0131 , \configuration_pci_ta1_reg[24]/NET0131 , \configuration_pci_ta1_reg[25]/NET0131 , \configuration_pci_ta1_reg[26]/NET0131 , \configuration_pci_ta1_reg[27]/NET0131 , \configuration_pci_ta1_reg[28]/NET0131 , \configuration_pci_ta1_reg[29]/NET0131 , \configuration_pci_ta1_reg[30]/NET0131 , \configuration_pci_ta1_reg[31]/NET0131 , \configuration_pci_ta1_reg[8]/NET0131 , \configuration_pci_ta1_reg[9]/NET0131 , \configuration_rst_inactive_reg/NET0131 , \configuration_set_isr_bit2_reg/NET0131 , \configuration_set_pci_err_cs_bit8_reg/NET0131 , \configuration_status_bit15_11_reg[11]/NET0131 , \configuration_status_bit15_11_reg[12]/NET0131 , \configuration_status_bit15_11_reg[13]/NET0131 , \configuration_status_bit15_11_reg[14]/NET0131 , \configuration_status_bit15_11_reg[15]/NET0131 , \configuration_status_bit8_reg/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131 , \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 , \configuration_sync_command_bit_reg/NET0131 , \configuration_sync_isr_2_del_bit_reg/NET0131 , \configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131 , \configuration_sync_isr_2_delayed_del_bit_reg/NET0131 , \configuration_sync_isr_2_sync_bckp_bit_reg/NET0131 , \configuration_sync_isr_2_sync_del_bit_reg/NET0131 , \configuration_sync_pci_err_cs_8_del_bit_reg/NET0131 , \configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131 , \configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131 , \configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131 , \configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131 , \configuration_wb_am1_reg[31]/NET0131 , \configuration_wb_am2_reg[31]/NET0131 , \configuration_wb_ba1_bit0_reg/NET0131 , \configuration_wb_ba1_bit31_12_reg[31]/NET0131 , \configuration_wb_ba2_bit0_reg/NET0131 , \configuration_wb_ba2_bit31_12_reg[31]/NET0131 , \configuration_wb_err_addr_reg[0]/NET0131 , \configuration_wb_err_addr_reg[10]/NET0131 , \configuration_wb_err_addr_reg[11]/NET0131 , \configuration_wb_err_addr_reg[12]/NET0131 , \configuration_wb_err_addr_reg[13]/NET0131 , \configuration_wb_err_addr_reg[14]/NET0131 , \configuration_wb_err_addr_reg[15]/NET0131 , \configuration_wb_err_addr_reg[16]/NET0131 , \configuration_wb_err_addr_reg[17]/NET0131 , \configuration_wb_err_addr_reg[18]/NET0131 , \configuration_wb_err_addr_reg[19]/NET0131 , \configuration_wb_err_addr_reg[1]/NET0131 , \configuration_wb_err_addr_reg[20]/NET0131 , \configuration_wb_err_addr_reg[21]/NET0131 , \configuration_wb_err_addr_reg[22]/NET0131 , \configuration_wb_err_addr_reg[23]/NET0131 , \configuration_wb_err_addr_reg[24]/NET0131 , \configuration_wb_err_addr_reg[25]/NET0131 , \configuration_wb_err_addr_reg[26]/NET0131 , \configuration_wb_err_addr_reg[27]/NET0131 , \configuration_wb_err_addr_reg[28]/NET0131 , \configuration_wb_err_addr_reg[29]/NET0131 , \configuration_wb_err_addr_reg[2]/NET0131 , \configuration_wb_err_addr_reg[30]/NET0131 , \configuration_wb_err_addr_reg[31]/NET0131 , \configuration_wb_err_addr_reg[3]/NET0131 , \configuration_wb_err_addr_reg[4]/NET0131 , \configuration_wb_err_addr_reg[5]/NET0131 , \configuration_wb_err_addr_reg[6]/NET0131 , \configuration_wb_err_addr_reg[7]/NET0131 , \configuration_wb_err_addr_reg[8]/NET0131 , \configuration_wb_err_addr_reg[9]/NET0131 , \configuration_wb_err_cs_bit0_reg/NET0131 , \configuration_wb_err_cs_bit31_24_reg[24]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[25]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[26]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[27]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[28]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[29]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[30]/NET0131 , \configuration_wb_err_cs_bit31_24_reg[31]/NET0131 , \configuration_wb_err_cs_bit8_reg/NET0131 , \configuration_wb_err_cs_bit9_reg/NET0131 , \configuration_wb_err_data_reg[0]/NET0131 , \configuration_wb_err_data_reg[10]/NET0131 , \configuration_wb_err_data_reg[11]/NET0131 , \configuration_wb_err_data_reg[12]/NET0131 , \configuration_wb_err_data_reg[13]/NET0131 , \configuration_wb_err_data_reg[14]/NET0131 , \configuration_wb_err_data_reg[15]/NET0131 , \configuration_wb_err_data_reg[16]/NET0131 , \configuration_wb_err_data_reg[17]/NET0131 , \configuration_wb_err_data_reg[18]/NET0131 , \configuration_wb_err_data_reg[19]/NET0131 , \configuration_wb_err_data_reg[1]/NET0131 , \configuration_wb_err_data_reg[20]/NET0131 , \configuration_wb_err_data_reg[21]/NET0131 , \configuration_wb_err_data_reg[22]/NET0131 , \configuration_wb_err_data_reg[23]/NET0131 , \configuration_wb_err_data_reg[24]/NET0131 , \configuration_wb_err_data_reg[25]/NET0131 , \configuration_wb_err_data_reg[26]/NET0131 , \configuration_wb_err_data_reg[27]/NET0131 , \configuration_wb_err_data_reg[28]/NET0131 , \configuration_wb_err_data_reg[29]/NET0131 , \configuration_wb_err_data_reg[2]/NET0131 , \configuration_wb_err_data_reg[30]/NET0131 , \configuration_wb_err_data_reg[31]/NET0131 , \configuration_wb_err_data_reg[3]/NET0131 , \configuration_wb_err_data_reg[4]/NET0131 , \configuration_wb_err_data_reg[5]/NET0131 , \configuration_wb_err_data_reg[6]/NET0131 , \configuration_wb_err_data_reg[7]/NET0131 , \configuration_wb_err_data_reg[8]/NET0131 , \configuration_wb_err_data_reg[9]/NET0131 , \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131 , \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131 , \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131 , \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131 , \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131 , \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131 , \configuration_wb_init_complete_out_reg/NET0131 , \configuration_wb_ta1_reg[31]/NET0131 , \configuration_wb_ta2_reg[31]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131 , \i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 , \input_register_pci_ad_reg_out_reg[0]/NET0131 , \input_register_pci_ad_reg_out_reg[10]/NET0131 , \input_register_pci_ad_reg_out_reg[11]/NET0131 , \input_register_pci_ad_reg_out_reg[12]/NET0131 , \input_register_pci_ad_reg_out_reg[13]/NET0131 , \input_register_pci_ad_reg_out_reg[14]/NET0131 , \input_register_pci_ad_reg_out_reg[15]/NET0131 , \input_register_pci_ad_reg_out_reg[16]/NET0131 , \input_register_pci_ad_reg_out_reg[17]/NET0131 , \input_register_pci_ad_reg_out_reg[18]/NET0131 , \input_register_pci_ad_reg_out_reg[19]/NET0131 , \input_register_pci_ad_reg_out_reg[1]/NET0131 , \input_register_pci_ad_reg_out_reg[20]/NET0131 , \input_register_pci_ad_reg_out_reg[21]/NET0131 , \input_register_pci_ad_reg_out_reg[22]/NET0131 , \input_register_pci_ad_reg_out_reg[23]/NET0131 , \input_register_pci_ad_reg_out_reg[24]/NET0131 , \input_register_pci_ad_reg_out_reg[25]/NET0131 , \input_register_pci_ad_reg_out_reg[26]/NET0131 , \input_register_pci_ad_reg_out_reg[27]/NET0131 , \input_register_pci_ad_reg_out_reg[28]/NET0131 , \input_register_pci_ad_reg_out_reg[29]/NET0131 , \input_register_pci_ad_reg_out_reg[2]/NET0131 , \input_register_pci_ad_reg_out_reg[30]/NET0131 , \input_register_pci_ad_reg_out_reg[31]/NET0131 , \input_register_pci_ad_reg_out_reg[3]/NET0131 , \input_register_pci_ad_reg_out_reg[4]/NET0131 , \input_register_pci_ad_reg_out_reg[5]/NET0131 , \input_register_pci_ad_reg_out_reg[6]/NET0131 , \input_register_pci_ad_reg_out_reg[7]/NET0131 , \input_register_pci_ad_reg_out_reg[8]/NET0131 , \input_register_pci_ad_reg_out_reg[9]/NET0131 , \input_register_pci_cbe_reg_out_reg[0]/NET0131 , \input_register_pci_cbe_reg_out_reg[1]/NET0131 , \input_register_pci_cbe_reg_out_reg[2]/NET0131 , \input_register_pci_cbe_reg_out_reg[3]/NET0131 , \input_register_pci_devsel_reg_out_reg/NET0131 , \input_register_pci_frame_reg_out_reg/NET0131 , \input_register_pci_idsel_reg_out_reg/NET0131 , \input_register_pci_irdy_reg_out_reg/NET0131 , \input_register_pci_stop_reg_out_reg/NET0131 , \input_register_pci_trdy_reg_out_reg/NET0131 , \output_backup_ad_out_reg[0]/NET0131 , \output_backup_ad_out_reg[10]/NET0131 , \output_backup_ad_out_reg[11]/NET0131 , \output_backup_ad_out_reg[12]/NET0131 , \output_backup_ad_out_reg[13]/NET0131 , \output_backup_ad_out_reg[14]/NET0131 , \output_backup_ad_out_reg[15]/NET0131 , \output_backup_ad_out_reg[16]/NET0131 , \output_backup_ad_out_reg[17]/NET0131 , \output_backup_ad_out_reg[18]/NET0131 , \output_backup_ad_out_reg[19]/NET0131 , \output_backup_ad_out_reg[1]/NET0131 , \output_backup_ad_out_reg[20]/NET0131 , \output_backup_ad_out_reg[21]/NET0131 , \output_backup_ad_out_reg[22]/NET0131 , \output_backup_ad_out_reg[23]/NET0131 , \output_backup_ad_out_reg[24]/NET0131 , \output_backup_ad_out_reg[25]/NET0131 , \output_backup_ad_out_reg[26]/NET0131 , \output_backup_ad_out_reg[27]/NET0131 , \output_backup_ad_out_reg[28]/NET0131 , \output_backup_ad_out_reg[29]/NET0131 , \output_backup_ad_out_reg[2]/NET0131 , \output_backup_ad_out_reg[30]/NET0131 , \output_backup_ad_out_reg[31]/NET0131 , \output_backup_ad_out_reg[3]/NET0131 , \output_backup_ad_out_reg[4]/NET0131 , \output_backup_ad_out_reg[5]/NET0131 , \output_backup_ad_out_reg[6]/NET0131 , \output_backup_ad_out_reg[7]/NET0131 , \output_backup_ad_out_reg[8]/NET0131 , \output_backup_ad_out_reg[9]/NET0131 , \output_backup_cbe_en_out_reg/NET0131 , \output_backup_cbe_out_reg[0]/NET0131 , \output_backup_cbe_out_reg[1]/NET0131 , \output_backup_cbe_out_reg[2]/NET0131 , \output_backup_cbe_out_reg[3]/NET0131 , \output_backup_devsel_out_reg/NET0131 , \output_backup_frame_en_out_reg/NET0131 , \output_backup_frame_out_reg/NET0131 , \output_backup_irdy_en_out_reg/NET0131 , \output_backup_irdy_out_reg/NET0131 , \output_backup_mas_ad_en_out_reg/NET0131 , \output_backup_par_en_out_reg/NET0131 , \output_backup_par_out_reg/NET0131 , \output_backup_perr_en_out_reg/NET0131 , \output_backup_perr_out_reg/NET0131 , \output_backup_serr_en_out_reg/NET0131 , \output_backup_serr_out_reg/NET0131 , \output_backup_stop_out_reg/NET0131 , \output_backup_tar_ad_en_out_reg/NET0131 , \output_backup_trdy_en_out_reg/NET0131 , \output_backup_trdy_out_reg/NET0131 , \parity_checker_check_for_serr_on_second_reg/NET0131 , \parity_checker_check_perr_reg/NET0131 , \parity_checker_frame_dec2_reg/NET0131 , \parity_checker_master_perr_report_reg/NET0131 , \parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131 , \parity_checker_perr_sampled_reg/NET0131 , \pci_cbe_i[0]_pad , \pci_cbe_i[1]_pad , \pci_cbe_i[2]_pad , \pci_cbe_i[3]_pad , pci_devsel_i_pad, pci_frame_i_pad, pci_frame_o_pad, pci_gnt_i_pad, pci_irdy_i_pad, pci_par_i_pad, pci_perr_i_pad, pci_rst_i_pad, pci_stop_i_pad, \pci_target_unit_del_sync_addr_out_reg[0]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[10]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[11]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[12]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[13]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[14]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[15]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[16]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[17]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[18]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[19]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[1]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[20]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[21]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[22]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[23]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[24]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[25]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[26]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[27]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[28]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[29]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[2]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[30]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[31]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[3]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[4]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[5]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[6]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[7]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[8]/NET0131 , \pci_target_unit_del_sync_addr_out_reg[9]/NET0131 , \pci_target_unit_del_sync_bc_out_reg[0]/NET0131 , \pci_target_unit_del_sync_bc_out_reg[1]/NET0131 , \pci_target_unit_del_sync_bc_out_reg[2]/NET0131 , \pci_target_unit_del_sync_bc_out_reg[3]/NET0131 , \pci_target_unit_del_sync_be_out_reg[0]/NET0131 , \pci_target_unit_del_sync_be_out_reg[1]/NET0131 , \pci_target_unit_del_sync_be_out_reg[2]/NET0131 , \pci_target_unit_del_sync_be_out_reg[3]/NET0131 , \pci_target_unit_del_sync_burst_out_reg/NET0131 , \pci_target_unit_del_sync_comp_comp_pending_reg/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131 , \pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131 , \pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131 , \pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131 , \pci_target_unit_del_sync_comp_flush_out_reg/NET0131 , \pci_target_unit_del_sync_comp_req_pending_reg/NET0131 , \pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131 , \pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131 , \pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131 , \pci_target_unit_del_sync_req_comp_pending_reg/NET0131 , \pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131 , \pci_target_unit_del_sync_req_done_reg_reg/NET0131 , \pci_target_unit_del_sync_req_req_pending_reg/NET0131 , \pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131 , \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131 , \pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131 , \pci_target_unit_fifos_inGreyCount_reg[0]/NET0131 , \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131 , \pci_target_unit_fifos_outGreyCount_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131 , \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001 , \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131 , \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001 , \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001 , \pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131 , \pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131 , \pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131 , \pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131 , \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 , \pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 , \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 , \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 , \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131 , \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 , \pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 , \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131 , \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131 , \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 , \pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131 , \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 , \pci_target_unit_pci_target_if_target_rd_reg/NET0131 , \pci_target_unit_pci_target_sm_backoff_reg/NET0131 , \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 , \pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 , \pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 , \pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 , \pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 , \pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131 , \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 , \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131 , \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131 , \pci_target_unit_pci_target_sm_rd_request_reg/NET0131 , \pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131 , \pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131 , \pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131 , \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131 , \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131 , \pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 , \pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131 , \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131 , \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 , \pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 , \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 , \pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131 , \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131 , \pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131 , \pci_target_unit_wishbone_master_read_bound_reg/NET0131 , \pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 , \pci_target_unit_wishbone_master_read_count_reg[1]/NET0131 , \pci_target_unit_wishbone_master_read_count_reg[2]/NET0131 , \pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 , \pci_target_unit_wishbone_master_retried_reg/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131 , \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131 , \pci_target_unit_wishbone_master_w_attempt_reg/NET0131 , \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131 , \pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131 , pci_trdy_i_pad, wb_int_i_pad, wbm_ack_i_pad, \wbm_adr_o[0]_pad , \wbm_adr_o[10]_pad , \wbm_adr_o[11]_pad , \wbm_adr_o[12]_pad , \wbm_adr_o[13]_pad , \wbm_adr_o[14]_pad , \wbm_adr_o[15]_pad , \wbm_adr_o[16]_pad , \wbm_adr_o[17]_pad , \wbm_adr_o[18]_pad , \wbm_adr_o[19]_pad , \wbm_adr_o[1]_pad , \wbm_adr_o[20]_pad , \wbm_adr_o[21]_pad , \wbm_adr_o[22]_pad , \wbm_adr_o[23]_pad , \wbm_adr_o[24]_pad , \wbm_adr_o[25]_pad , \wbm_adr_o[26]_pad , \wbm_adr_o[27]_pad , \wbm_adr_o[28]_pad , \wbm_adr_o[29]_pad , \wbm_adr_o[2]_pad , \wbm_adr_o[30]_pad , \wbm_adr_o[31]_pad , \wbm_adr_o[3]_pad , \wbm_adr_o[4]_pad , \wbm_adr_o[5]_pad , \wbm_adr_o[6]_pad , \wbm_adr_o[7]_pad , \wbm_adr_o[8]_pad , \wbm_adr_o[9]_pad , \wbm_cti_o[0]_pad , \wbm_dat_o[0]_pad , \wbm_dat_o[10]_pad , \wbm_dat_o[11]_pad , \wbm_dat_o[12]_pad , \wbm_dat_o[13]_pad , \wbm_dat_o[14]_pad , \wbm_dat_o[15]_pad , \wbm_dat_o[16]_pad , \wbm_dat_o[17]_pad , \wbm_dat_o[18]_pad , \wbm_dat_o[19]_pad , \wbm_dat_o[1]_pad , \wbm_dat_o[20]_pad , \wbm_dat_o[21]_pad , \wbm_dat_o[22]_pad , \wbm_dat_o[23]_pad , \wbm_dat_o[24]_pad , \wbm_dat_o[25]_pad , \wbm_dat_o[26]_pad , \wbm_dat_o[27]_pad , \wbm_dat_o[28]_pad , \wbm_dat_o[29]_pad , \wbm_dat_o[2]_pad , \wbm_dat_o[30]_pad , \wbm_dat_o[31]_pad , \wbm_dat_o[3]_pad , \wbm_dat_o[4]_pad , \wbm_dat_o[5]_pad , \wbm_dat_o[6]_pad , \wbm_dat_o[7]_pad , \wbm_dat_o[8]_pad , \wbm_dat_o[9]_pad , wbm_err_i_pad, wbm_rty_i_pad, \wbm_sel_o[0]_pad , \wbm_sel_o[1]_pad , \wbm_sel_o[2]_pad , \wbm_sel_o[3]_pad , \wbs_adr_i[10]_pad , \wbs_adr_i[11]_pad , \wbs_adr_i[12]_pad , \wbs_adr_i[13]_pad , \wbs_adr_i[14]_pad , \wbs_adr_i[15]_pad , \wbs_adr_i[16]_pad , \wbs_adr_i[17]_pad , \wbs_adr_i[18]_pad , \wbs_adr_i[19]_pad , \wbs_adr_i[20]_pad , \wbs_adr_i[21]_pad , \wbs_adr_i[22]_pad , \wbs_adr_i[23]_pad , \wbs_adr_i[24]_pad , \wbs_adr_i[25]_pad , \wbs_adr_i[26]_pad , \wbs_adr_i[27]_pad , \wbs_adr_i[28]_pad , \wbs_adr_i[29]_pad , \wbs_adr_i[2]_pad , \wbs_adr_i[30]_pad , \wbs_adr_i[31]_pad , \wbs_adr_i[3]_pad , \wbs_adr_i[4]_pad , \wbs_adr_i[5]_pad , \wbs_adr_i[6]_pad , \wbs_adr_i[7]_pad , \wbs_adr_i[8]_pad , \wbs_adr_i[9]_pad , \wbs_bte_i[0]_pad , \wbs_bte_i[1]_pad , \wbs_cti_i[0]_pad , \wbs_cti_i[1]_pad , \wbs_cti_i[2]_pad , wbs_cyc_i_pad, wbs_stb_i_pad, wbs_we_i_pad, \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131 , \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131 , \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 , \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131 , \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131 , \wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131 , \wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131 , \wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131 , \wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131 , \wishbone_slave_unit_del_sync_burst_out_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131 , \wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131 , \wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131 , \wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131 , \wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 , \wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131 , \wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131 , \wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 , \wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131 , \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131 , \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131 , \wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131 , \wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131 , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131 , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131 , \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001 , \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001 , \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001 , \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131 , \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131 , \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131 , \wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131 , \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131 , \wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131 , \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131 , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 , \wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 , \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 , \wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131 , \wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131 , \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 , \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131 , \wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131 , \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131 , \wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131 , \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_map_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131 , \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 , \configuration_init_complete_reg/P0001 , \configuration_interrupt_out_reg/P0001 , \g21/_0_ , \g52241/_0_ , \g52244/_0_ , \g52348/_0_ , \g52349/_0_ , \g52350/_0_ , \g52351/_0_ , \g52352/_0_ , \g52390/_0_ , \g52391/_0_ , \g52393/_3_ , \g52394/_3_ , \g52395/_3_ , \g52396/_3_ , \g52397/_3_ , \g52398/_3_ , \g52399/_3_ , \g52400/_3_ , \g52401/_3_ , \g52402/_3_ , \g52403/_3_ , \g52404/_3_ , \g52405/_3_ , \g52406/_0_ , \g52408/_0_ , \g52409/_0_ , \g52410/_0_ , \g52411/_0_ , \g52412/_0_ , \g52413/_0_ , \g52414/_0_ , \g52415/_0_ , \g52416/_0_ , \g52417/_0_ , \g52418/_0_ , \g52419/_0_ , \g52421/_0_ , \g52422/_0_ , \g52423/_0_ , \g52424/_0_ , \g52425/_0_ , \g52426/_0_ , \g52427/_0_ , \g52428/_0_ , \g52429/_0_ , \g52430/_0_ , \g52431/_0_ , \g52432/_0_ , \g52433/_0_ , \g52434/_0_ , \g52435/_0_ , \g52436/_0_ , \g52437/_0_ , \g52439/_3_ , \g52440/_3_ , \g52441/_3_ , \g52442/_3_ , \g52443/_3_ , \g52444/_3_ , \g52445/_3_ , \g52446/_3_ , \g52447/_3_ , \g52448/_3_ , \g52449/_3_ , \g52450/_3_ , \g52451/_3_ , \g52452/_3_ , \g52453/_3_ , \g52454/_3_ , \g52455/_3_ , \g52456/_3_ , \g52457/_3_ , \g52458/_3_ , \g52459/_3_ , \g52460/_3_ , \g52461/_3_ , \g52462/_3_ , \g52463/_3_ , \g52464/_3_ , \g52465/_3_ , \g52466/_3_ , \g52467/_3_ , \g52468/_3_ , \g52469/_3_ , \g52470/_3_ , \g52471/_3_ , \g52472/_3_ , \g52473/_3_ , \g52474/_3_ , \g52475/_3_ , \g52476/_3_ , \g52477/_3_ , \g52478/_3_ , \g52479/_3_ , \g52480/_3_ , \g52481/_3_ , \g52482/_3_ , \g52483/_3_ , \g52484/_3_ , \g52485/_3_ , \g52499/_0_ , \g52500/_0_ , \g52501/_0_ , \g52547/_0_ , \g52550/_0_ , \g52553/_0_ , \g52675/_0__syn_2 , \g52714/_0_ , \g52715/_0_ , \g52716/_0_ , \g52717/_0_ , \g52718/_0_ , \g52720/_0_ , \g52865/_0_ , \g52867/_0_ , \g52867/_1_ , \g52868/_0_ , \g52871/_2_ , \g52897/_0_ , \g52898/_0_ , \g52899/_0_ , \g52900/_0_ , \g52901/_0_ , \g52902/_0_ , \g52903/_0_ , \g52904/_0_ , \g52905/_0_ , \g52906/_0_ , \g52907/_0_ , \g52908/_0_ , \g52909/_0_ , \g52910/_0_ , \g52911/_0_ , \g52912/_0_ , \g52913/_0_ , \g52914/_0_ , \g52915/_0_ , \g52916/_0_ , \g52917/_0_ , \g52918/_0_ , \g52920/_0_ , \g52921/_0_ , \g52922/_0_ , \g52923/_0_ , \g52924/_0_ , \g52925/_0_ , \g52948/_0_ , \g52958/_0_ , \g52959/_0_ , \g52960/_0_ , \g52961/_0_ , \g52962/_0_ , \g52963/_0_ , \g52965/_0_ , \g52966/_0_ , \g52969/_0_ , \g52970/_0_ , \g52971/_0_ , \g52972/_0_ , \g52973/_0_ , \g52975/_0_ , \g52976/_0_ , \g52977/_0_ , \g52978/_0_ , \g52979/_0_ , \g52980/_0_ , \g52981/_0_ , \g52982/_0_ , \g52983/_0_ , \g52984/_0_ , \g52985/_0_ , \g52986/_0_ , \g52988/_0_ , \g52990/_0_ , \g52991/_0_ , \g52993/_0_ , \g52994/_0_ , \g52996/_0_ , \g52997/_0_ , \g53068/_0_ , \g53085/_0_ , \g53086/_0_ , \g53088/_0_ , \g53089/_0_ , \g53090/_0_ , \g53091/_0_ , \g53096/_0_ , \g53123/_0_ , \g53124/_0_ , \g53137/_0_ , \g53137/_1_ , \g53145/_0_ , \g53146/_0_ , \g53147/_0_ , \g53870/_0_ , \g53871/_0_ , \g53872/_0_ , \g53873/_0_ , \g53874/_0_ , \g53875/_0_ , \g53876/_0_ , \g53877/_0_ , \g53878/_0_ , \g53879/_0_ , \g53880/_0_ , \g53881/_0_ , \g53882/_0_ , \g53883/_0_ , \g53884/_0_ , \g53885/_0_ , \g53886/_0_ , \g53887/_0_ , \g53888/_0_ , \g53889/_0_ , \g53890/_3_ , \g53897/_3_ , \g53935/_3_ , \g53936/_3_ , \g53937/_3_ , \g53938/_3_ , \g53939/_3_ , \g53940/_3_ , \g53941/_3_ , \g53942/_3_ , \g54022/_0_ , \g54160/_3_ , \g54163/_3_ , \g54166/_3_ , \g54167/_2_ , \g54168/_3_ , \g54169/_3_ , \g54170/_3_ , \g54171/_2_ , \g54172/_3_ , \g54173/_3_ , \g54204/_2_ , \g54205/_2_ , \g54206/_2_ , \g54207/_2_ , \g54208/_2_ , \g54209/_2_ , \g54210/_2_ , \g54211/_2_ , \g54212/_2_ , \g54213/_2_ , \g54214/_2_ , \g54215/_2_ , \g54216/_2_ , \g54217/_2_ , \g54218/_2_ , \g54219/_2_ , \g54220/_2_ , \g54221/_2_ , \g54222/_2_ , \g54223/_2_ , \g54224/_2_ , \g54225/_2_ , \g54226/_2_ , \g54227/_2_ , \g54228/_2_ , \g54229/_2_ , \g54230/_2_ , \g54231/_2_ , \g54232/_2_ , \g54233/_2_ , \g54267/_0_ , \g54268/_0_ , \g54269/_0_ , \g54270/_0_ , \g54271/_0_ , \g54272/_0_ , \g54273/_0_ , \g54274/_0_ , \g54275/_0_ , \g54276/_0_ , \g54278/_0_ , \g54279/_0_ , \g54280/_0_ , \g54281/_0_ , \g54282/_0_ , \g54283/_0_ , \g54284/_0_ , \g54285/_0_ , \g54286/_0_ , \g54287/_0_ , \g54288/_0_ , \g54289/_0_ , \g54290/_0_ , \g54291/_0_ , \g54292/_0_ , \g54293/_0_ , \g54294/_0_ , \g54296/_0_ , \g54297/_0_ , \g54298/_0_ , \g54299/_0_ , \g54300/_0_ , \g54301/_0_ , \g54302/_0_ , \g54303/_0_ , \g54329/_0_ , \g54453/_0_ , \g54466/_0_ , \g54470/_0_ , \g54470/_1_ , \g54496/_0_ , \g54597/_0_ , \g54628/_0_ , \g54629/_0_ , \g54630/_0_ , \g54631/_0_ , \g54632/_0_ , \g54633/_0_ , \g54634/_0_ , \g54635/_0_ , \g54636/_0_ , \g54638/_0_ , \g54639/_0_ , \g54640/_0_ , \g54641/_0_ , \g54642/_0_ , \g54643/_0_ , \g54645/_0_ , \g54646/_0_ , \g54647/_0_ , \g54648/_0_ , \g54649/_0_ , \g54650/_0_ , \g54651/_0_ , \g54652/_0_ , \g54653/_0_ , \g54654/_0_ , \g54655/_0_ , \g54656/_0_ , \g54657/_0_ , \g54658/_0_ , \g54659/_0_ , \g54660/_0_ , \g54661/_0_ , \g54662/_0_ , \g54663/_0_ , \g54664/_0_ , \g54669/_0_ , \g54832/_0_ , \g54833/_0_ , \g54867/_0_ , \g54868/_0_ , \g54869/_0_ , \g54870/_0_ , \g54871/_0_ , \g54872/_0_ , \g54873/_0_ , \g54874/_0_ , \g54875/_0_ , \g54876/_0_ , \g54877/_0_ , \g54878/_0_ , \g54879/_0_ , \g54880/_0_ , \g54881/_0_ , \g54882/_0_ , \g54883/_0_ , \g54884/_0_ , \g54885/_0_ , \g54886/_0_ , \g54887/_0_ , \g54888/_0_ , \g54889/_0_ , \g54890/_0_ , \g54891/_0_ , \g54892/_0_ , \g54893/_0_ , \g54894/_0_ , \g54895/_0_ , \g54896/_0_ , \g54897/_0_ , \g54898/_0_ , \g54899/_0_ , \g56438/_0_ , \g56439/_0_ , \g56933/_3_ , \g56934/_3_ , \g56960/_0_ , \g56960/_1_ , \g56961/_3__syn_2 , \g57019/_0_ , \g57020/_0_ , \g57021/_0_ , \g57022/_0_ , \g57023/_0_ , \g57024/_0_ , \g57025/_0_ , \g57026/_0_ , \g57027/_0_ , \g57028/_0_ , \g57029/_0_ , \g57031/_0_ , \g57032/_0_ , \g57034/u3_syn_4 , \g57069/u3_syn_4 , \g57104/u3_syn_4 , \g57139/u3_syn_4 , \g57174/u3_syn_4 , \g57209/u3_syn_4 , \g57244/u3_syn_4 , \g57276/u3_syn_4 , \g57308/u3_syn_4 , \g57340/u3_syn_4 , \g57372/u3_syn_4 , \g57404/u3_syn_4 , \g57408/u3_syn_4 , \g57444/u3_syn_4 , \g57480/u3_syn_4 , \g57516/u3_syn_4 , \g57646/_0_ , \g57649/_0_ , \g57779/_3_ , \g57780/_3_ , \g57781/_3_ , \g57782/_3_ , \g57783/_3_ , \g57784/_3_ , \g57785/_3_ , \g57786/_3_ , \g57787/_3_ , \g57788/_3_ , \g57789/_3_ , \g57791/_3_ , \g57795/_3_ , \g57796/_3_ , \g57797/_3_ , \g57798/_3_ , \g57799/_3_ , \g57800/_3_ , \g57801/_3_ , \g57802/_3_ , \g57850/_0_ , \g57852/_0_ , \g57871/_0_ , \g57872/_0_ , \g57873/_0_ , \g58/_0_ , \g58490/_0_ , \g58564/_0_ , \g58569/_0_ , \g58571/_0_ , \g58573/_0_ , \g58577/_0_ , \g58578/_0_ , \g58579/_0_ , \g58580/_0_ , \g58583/_0_ , \g58584/_0_ , \g58603/_0_ , \g58611/_3_ , \g58637/_0_ , \g58638/_0_ , \g58639/_0_ , \g58691/_0_ , \g58693/_0_ , \g58696/_0_ , \g58700/_0_ , \g58701/_0_ , \g58708/_1_ , \g58730/_0_ , \g58731/_0_ , \g58732/_0_ , \g58733/_0_ , \g58734/_0_ , \g58735/_0_ , \g58736/_0_ , \g58737/_0_ , \g58738/_0_ , \g58739/_0_ , \g58740/_0_ , \g58741/_1__syn_2 , \g58748/_0_ , \g58751/_0_ , \g58752/_0_ , \g58753/_0_ , \g58754/_0_ , \g58756/_0_ , \g58767/_3_ , \g58768/_3_ , \g58769/_3_ , \g58770/_3_ , \g58771/_3_ , \g58772/_3_ , \g58773/_3_ , \g58774/_3_ , \g58775/_3_ , \g58776/_3_ , \g58777/_3_ , \g58778/_3_ , \g58779/_3_ , \g58780/_3_ , \g58781/_3_ , \g58782/_3_ , \g58783/_3_ , \g58784/_3_ , \g58785/_3_ , \g58786/_3_ , \g58787/_3_ , \g58788/_3_ , \g58789/_3_ , \g58790/_3_ , \g58791/_3_ , \g58792/_3_ , \g58793/_3_ , \g58794/_3_ , \g58795/_3_ , \g58796/_3_ , \g58797/_3_ , \g58798/_3_ , \g58874/_0_ , \g59064/_1_ , \g59072/_0_ , \g59080/_0_ , \g59083/_0_ , \g59084/_0_ , \g59085/_0_ , \g59088/_0_ , \g59094/_0_ , \g59095/_0_ , \g59126/_3_ , \g59128/_0_ , \g59174/_2_ , \g59180/_0_ , \g59181/_0_ , \g59182/_0_ , \g59190/_0_ , \g59191/_0_ , \g59192/_0_ , \g59204/_0_ , \g59205/_0_ , \g59210/_3_ , \g59213/_0_ , \g59214/_0_ , \g59215/_0_ , \g59216/_0_ , \g59217/_0_ , \g59218/_0_ , \g59219/_0_ , \g59220/_0_ , \g59221/_0_ , \g59222/_0_ , \g59223/_0_ , \g59226/_3_ , \g59232/_00_ , \g59233/_0_ , \g59235/_0_ , \g59236/_0_ , \g59237/_0_ , \g59238/_0_ , \g59318/_0_ , \g59331/_0_ , \g59336/_0_ , \g59351/_0_ , \g59354/_0_ , \g59358/_0_ , \g59363/_0_ , \g59366/_0_ , \g59370/u3_syn_4 , \g59371/u3_syn_4 , \g59372/u3_syn_4 , \g59373/u3_syn_4 , \g59378/u3_syn_4 , \g59379/u3_syn_4 , \g59380/u3_syn_4 , \g59381/u3_syn_4 , \g59589/_0_ , \g59655/_0_ , \g59662/_0_ , \g59735/_0_ , \g59739/_0_ , \g59740/_0_ , \g59741/_0_ , \g59742/_0_ , \g59743/_0_ , \g59744/_0_ , \g59745/_0_ , \g59746/_0_ , \g59747/_0_ , \g59748/_0_ , \g59749/_0_ , \g59750/_0_ , \g59751/_0_ , \g59752/_0_ , \g59753/_0_ , \g59754/_0_ , \g59755/_0_ , \g59756/_0_ , \g59757/_0_ , \g59758/_0_ , \g59759/_0_ , \g59760/_0_ , \g59764/_0_ , \g59766/_0_ , \g59774/_0_ , \g59775/_0_ , \g59776/_0_ , \g59777/_0_ , \g59778/_0_ , \g59779/_0_ , \g59780/_0_ , \g59781/_0_ , \g59789/_3_ , \g59799/_3_ , \g60311/_0_ , \g60326/_0_ , \g60333/_0_ , \g60336/_3_ , \g60341/_0_ , \g60343/_0_ , \g60344/_0_ , \g60345/_0_ , \g60354/_0_ , \g60355/_0_ , \g60356/_0_ , \g60357/_0_ , \g60358/_0_ , \g60359/_0_ , \g60360/_0_ , \g60361/_0_ , \g60362/_0_ , \g60363/_0_ , \g60364/_0_ , \g60398/_2_ , \g60399/_0_ , \g60400/_0_ , \g60401/_0_ , \g60402/_0_ , \g60403/_0_ , \g60406/_0_ , \g60410/_0_ , \g60411/_0_ , \g60417/_3_ , \g60419/_3_ , \g60421/_3_ , \g60423/_3_ , \g60425/_3_ , \g60427/_3_ , \g60429/_3_ , \g60431/_3_ , \g60433/_3_ , \g60435/_3_ , \g60437/_3_ , \g60439/_3_ , \g60441/_3_ , \g60443/_3_ , \g60445/_3_ , \g60447/_3_ , \g60449/_3_ , \g60451/_3_ , \g60453/_3_ , \g60455/_3_ , \g60457/_3_ , \g60459/_3_ , \g60461/_3_ , \g60463/_3_ , \g60465/_3_ , \g60467/_3_ , \g60469/_3_ , \g60471/_3_ , \g60473/_3_ , \g60475/_3_ , \g60477/_3_ , \g60479/_3_ , \g60481/_3_ , \g60483/_3_ , \g60485/_3_ , \g60487/_3_ , \g60489/_3_ , \g60491/_3_ , \g60493/_3_ , \g60495/_3_ , \g60497/_3_ , \g60499/_3_ , \g60501/_3_ , \g60503/_3_ , \g60505/_3_ , \g60507/_3_ , \g60509/_3_ , \g60511/_3_ , \g60513/_3_ , \g60515/_3_ , \g60517/_3_ , \g60519/_3_ , \g60521/_3_ , \g60523/_3_ , \g60525/_3_ , \g60527/_3_ , \g60529/_3_ , \g60531/_3_ , \g60533/_3_ , \g60535/_3_ , \g60537/_3_ , \g60539/_3_ , \g60541/_3_ , \g60544/_3_ , \g60546/_3_ , \g60548/_3_ , \g60550/_3_ , \g60552/_3_ , \g60554/_3_ , \g60556/_3_ , \g60559/_3_ , \g60561/_3_ , \g60563/_3_ , \g60565/_3_ , \g60567/_3_ , \g60569/_3_ , \g60571/_3_ , \g60573/_3_ , \g60575/_3_ , \g60577/_3_ , \g60579/_3_ , \g60581/_3_ , \g60583/_3_ , \g60585/_3_ , \g60588/_3_ , \g60590/_3_ , \g60593/_3_ , \g60596/_3_ , \g60598/_3_ , \g60600/_3_ , \g60602/_3_ , \g60603/_3_ , \g60671/_3_ , \g60672/_3_ , \g60674/_3_ , \g60680/_0_ , \g60682/_3_ , \g60690/_3_ , \g60692/_3_ , \g61594/_0_ , \g61614/_0_ , \g61618/_00_ , \g61649/_0_ , \g61651/_0_ , \g61656/_0_ , \g61657/_0_ , \g61659/_0_ , \g61662/_0_ , \g61663/_0_ , \g61664/_0_ , \g61665/_0_ , \g61667/_2_ , \g61669/_3__syn_2 , \g61678/_0_ , \g61679/_0_ , \g61680/_0_ , \g61681/_0_ , \g61684/_0_ , \g61685/_0_ , \g61686/_0_ , \g61690/_0_ , \g61692/_0_ , \g61694/_0_ , \g61695/_0_ , \g61696/_0_ , \g61699/u3_syn_4 , \g61732/u3_syn_4 , \g61765/u3_syn_4 , \g61798/u3_syn_4 , \g61848/_0_ , \g61848/_3_ , \g61853/_0_ , \g61854/_1__syn_2 , \g61858/u3_syn_4 , \g61880/u3_syn_4 , \g61887/u3_syn_4 , \g61920/u3_syn_4 , \g61990/u3_syn_4 , \g62254/_0__syn_2 , \g62260/_0_ , \g62262/_1__syn_2 , \g62290/_0_ , \g62317/_0_ , \g62319/_0_ , \g62324/_0_ , \g62329/_0_ , \g62331/_0_ , \g62331/_1_ , \g62333/u3_syn_4 , \g62335/u3_syn_4 , \g62336/u3_syn_4 , \g62428/u3_syn_4 , \g62454/u3_syn_4 , \g62487/u3_syn_4 , \g62520/u3_syn_4 , \g62552/u3_syn_4 , \g62584/u3_syn_4 , \g62619/u3_syn_4 , \g62651/u3_syn_4 , \g62692/_0_ , \g62873/_0_ , \g62882/_0_ , \g62883/u3_syn_4 , \g62886/u3_syn_4 , \g62908/u3_syn_4 , \g62952/u3_syn_4 , \g62974/u3_syn_4 , \g63207/_0_ , \g63214/_3_ , \g63227/_0_ , \g63250/_1__syn_2 , \g63315/_0__syn_2 , \g63320/_0_ , \g63322/_0_ , \g63324/_2_ , \g63338/_0__syn_2 , \g63340/_0_ , \g63376/_0_ , \g63395/_2_ , \g63398/_0_ , \g63419/_0_ , \g63524/_3_ , \g63540/_0_ , \g63541/_0_ , \g63682/_0_ , \g63890/_1_ , \g63892/_0_ , \g63894/_0_ , \g63897/_1_ , \g63908/_0_ , \g63913/_0_ , \g63914/_0_ , \g63927/_1__syn_2 , \g63934/_0_ , \g63942/_0_ , \g63952/_0_ , \g63965/_0_ , \g63969/_0_ , \g63985/_0_ , \g63986/_0_ , \g63987/_0_ , \g63988/_0_ , \g63990/_0_ , \g63991/_0_ , \g63992/_0_ , \g63993/_0_ , \g64016/_0_ , \g64017/_0_ , \g64018/_0_ , \g64019/_0_ , \g64020/_0_ , \g64021/_0_ , \g64023/_0_ , \g64024/_0_ , \g64101/_0_ , \g64104/_0_ , \g64121/_0_ , \g64174/_0_ , \g64249/_0_ , \g64299/_0_ , \g64338/_0_ , \g64364/_0_ , \g64459/_0_ , \g64461/_0_ , \g64466/_0_ , \g64577/_0_ , \g64583/_0_ , \g64589/_1_ , \g64595/_0_ , \g64598/_0_ , \g64649/_0_ , \g64678/_0_ , \g64688/_3_ , \g64689/_0_ , \g64694/_0_ , \g64695/_0_ , \g64700/_0_ , \g64714/_0_ , \g64744/_2_ , \g65255/_0_ , \g65258/_0_ , \g65269/_3_ , \g65489/_0_ , \g65513/_0_ , \g65530/_0_ , \g65561/_0_ , \g65563/_0_ , \g65564/_0_ , \g65573/_0_ , \g65578/_2_ , \g65597/_0_ , \g65605/_0_ , \g65606/_0_ , \g65609/_0_ , \g65611/_0_ , \g65612/_0_ , \g65613/_0_ , \g65615/_0_ , \g65618/_0_ , \g65631/_0_ , \g65634/_0_ , \g65635/_0_ , \g65639/_0_ , \g65644/_0_ , \g65648/_0_ , \g65650/_0_ , \g65662/_3_ , \g65665/_3_ , \g65729/_0_ , \g65801/_0_ , \g66072/_0_ , \g66074/_0_ , \g66075/_0_ , \g66076/_0_ , \g66077/_0_ , \g66078/_0_ , \g66079/_0_ , \g66080/_0_ , \g66081/_0_ , \g66082/_0_ , \g66085/_0_ , \g66086/_0_ , \g66087/_0_ , \g66089/_0_ , \g66090/_0_ , \g66093/_0_ , \g66094/_0_ , \g66095/_0_ , \g66098/_0_ , \g66100/_0_ , \g66106/_1_ , \g66107/_0_ , \g66108/_0_ , \g66110/_0_ , \g66114/_0_ , \g66124/_0_ , \g66125/_0_ , \g66127/_0_ , \g66128/_0_ , \g66129/_0_ , \g66130/_0_ , \g66133/_0_ , \g66134/_0_ , \g66136/_0_ , \g66141/_1_ , \g66153/_0_ , \g66182/_0_ , \g66187/_0_ , \g66240/_0_ , \g66268/_0_ , \g66354/_0_ , \g66397/_3_ , \g66398/_3_ , \g66399/_3_ , \g66400/_3_ , \g66401/_3_ , \g66402/_3_ , \g66403/_3_ , \g66404/_3_ , \g66405/_3_ , \g66406/_3_ , \g66407/_3_ , \g66408/_3_ , \g66409/_3_ , \g66410/_3_ , \g66411/_3_ , \g66412/_3_ , \g66413/_3_ , \g66414/_3_ , \g66415/_3_ , \g66416/_3_ , \g66417/_3_ , \g66418/_3_ , \g66419/_3_ , \g66420/_3_ , \g66421/_3_ , \g66422/_3_ , \g66423/_3_ , \g66424/_3_ , \g66425/_3_ , \g66426/_3_ , \g66427/_3_ , \g66428/_3_ , \g66429/_3_ , \g66430/_3_ , \g66464/_0_ , \g66465/_0_ , \g66477/_3_ , \g66643/_0_ , \g66733/_2_ , \g66735/_1_ , \g66801/_0_ , \g66866/_0_ , \g66875/_0_ , \g66885/_1_ , \g66890/_0_ , \g66939/_0_ , \g66950/_0_ , \g67035/_0_ , \g67038/_0_ , \g67044/_3_ , \g67045/_3_ , \g67046/_3_ , \g67070/_3_ , \g67082/_3_ , \g67090/_3_ , \g67106/_0_ , \g67107/_0_ , \g67108/_0_ , \g67109/_0_ , \g67117/_0_ , \g67131/_0_ , \g67142/_0_ , \g67421/_0_ , \g67456/_0_ , \g67464/_0_ , \g67617/_1_ , \g67772/_0_ , \g68523/_0_ , \g73970/_0_ , \g73976/_0_ , \g74120/_1_ , \g74148/_2_ , \g74245/_0_ , \g74426/_0_ , \g74434/_3_ , \g74589/_0_ , \g74626/_1__syn_2 , \g74790/_0_ , \g74801/_0_ , \g74838/_0_ , \g74850/_0_ , \g74855/_0_ , \g74862/_0_ , \g74871/_0_ , \g74878/_0_ , \g74885/_0_ , \g74922/_0_ , \g75066/_1__syn_2 , \g75100/_1_ , \g75201/_1_ , \g75205/_1_ , \g75420/_1_ , pci_rst_oe_o_pad, wb_int_o_pad, wb_rst_o_pad);
	input \configuration_cache_line_size_reg_reg[0]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[1]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[2]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[3]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[4]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[5]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[6]/NET0131  ;
	input \configuration_cache_line_size_reg_reg[7]/NET0131  ;
	input \configuration_command_bit2_0_reg[0]/NET0131  ;
	input \configuration_command_bit2_0_reg[1]/NET0131  ;
	input \configuration_command_bit2_0_reg[2]/NET0131  ;
	input \configuration_command_bit6_reg/NET0131  ;
	input \configuration_command_bit8_reg/NET0131  ;
	input \configuration_icr_bit2_0_reg[0]/NET0131  ;
	input \configuration_icr_bit2_0_reg[1]/NET0131  ;
	input \configuration_icr_bit2_0_reg[2]/NET0131  ;
	input \configuration_icr_bit31_reg/NET0131  ;
	input \configuration_init_complete_reg/NET0131  ;
	input \configuration_interrupt_line_reg[0]/NET0131  ;
	input \configuration_interrupt_line_reg[1]/NET0131  ;
	input \configuration_interrupt_line_reg[2]/NET0131  ;
	input \configuration_interrupt_line_reg[3]/NET0131  ;
	input \configuration_interrupt_line_reg[4]/NET0131  ;
	input \configuration_interrupt_line_reg[5]/NET0131  ;
	input \configuration_interrupt_line_reg[6]/NET0131  ;
	input \configuration_interrupt_line_reg[7]/NET0131  ;
	input \configuration_interrupt_out_reg/NET0131  ;
	input \configuration_isr_bit2_0_reg[0]/NET0131  ;
	input \configuration_isr_bit2_0_reg[1]/NET0131  ;
	input \configuration_isr_bit2_0_reg[2]/NET0131  ;
	input \configuration_latency_timer_reg[0]/NET0131  ;
	input \configuration_latency_timer_reg[1]/NET0131  ;
	input \configuration_latency_timer_reg[2]/NET0131  ;
	input \configuration_latency_timer_reg[3]/NET0131  ;
	input \configuration_latency_timer_reg[4]/NET0131  ;
	input \configuration_latency_timer_reg[5]/NET0131  ;
	input \configuration_latency_timer_reg[6]/NET0131  ;
	input \configuration_latency_timer_reg[7]/NET0131  ;
	input \configuration_pci_am1_reg[10]/NET0131  ;
	input \configuration_pci_am1_reg[11]/NET0131  ;
	input \configuration_pci_am1_reg[12]/NET0131  ;
	input \configuration_pci_am1_reg[13]/NET0131  ;
	input \configuration_pci_am1_reg[14]/NET0131  ;
	input \configuration_pci_am1_reg[15]/NET0131  ;
	input \configuration_pci_am1_reg[16]/NET0131  ;
	input \configuration_pci_am1_reg[17]/NET0131  ;
	input \configuration_pci_am1_reg[18]/NET0131  ;
	input \configuration_pci_am1_reg[19]/NET0131  ;
	input \configuration_pci_am1_reg[20]/NET0131  ;
	input \configuration_pci_am1_reg[21]/NET0131  ;
	input \configuration_pci_am1_reg[22]/NET0131  ;
	input \configuration_pci_am1_reg[23]/NET0131  ;
	input \configuration_pci_am1_reg[24]/NET0131  ;
	input \configuration_pci_am1_reg[25]/NET0131  ;
	input \configuration_pci_am1_reg[26]/NET0131  ;
	input \configuration_pci_am1_reg[27]/NET0131  ;
	input \configuration_pci_am1_reg[28]/NET0131  ;
	input \configuration_pci_am1_reg[29]/NET0131  ;
	input \configuration_pci_am1_reg[30]/NET0131  ;
	input \configuration_pci_am1_reg[31]/NET0131  ;
	input \configuration_pci_am1_reg[8]/NET0131  ;
	input \configuration_pci_am1_reg[9]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[12]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[13]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[14]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[15]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[16]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[17]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[18]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[19]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[20]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[21]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[22]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[23]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[24]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[25]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[26]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[27]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[28]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[29]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[30]/NET0131  ;
	input \configuration_pci_ba0_bit31_8_reg[31]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[10]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[11]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[12]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[13]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[14]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[15]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[16]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[17]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[18]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[19]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[20]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[21]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[22]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[23]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[24]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[25]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[26]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[27]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[28]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[29]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[30]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[31]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[8]/NET0131  ;
	input \configuration_pci_ba1_bit31_8_reg[9]/NET0131  ;
	input \configuration_pci_err_addr_reg[0]/NET0131  ;
	input \configuration_pci_err_addr_reg[10]/NET0131  ;
	input \configuration_pci_err_addr_reg[11]/NET0131  ;
	input \configuration_pci_err_addr_reg[12]/NET0131  ;
	input \configuration_pci_err_addr_reg[13]/NET0131  ;
	input \configuration_pci_err_addr_reg[14]/NET0131  ;
	input \configuration_pci_err_addr_reg[15]/NET0131  ;
	input \configuration_pci_err_addr_reg[16]/NET0131  ;
	input \configuration_pci_err_addr_reg[17]/NET0131  ;
	input \configuration_pci_err_addr_reg[18]/NET0131  ;
	input \configuration_pci_err_addr_reg[19]/NET0131  ;
	input \configuration_pci_err_addr_reg[1]/NET0131  ;
	input \configuration_pci_err_addr_reg[20]/NET0131  ;
	input \configuration_pci_err_addr_reg[21]/NET0131  ;
	input \configuration_pci_err_addr_reg[22]/NET0131  ;
	input \configuration_pci_err_addr_reg[23]/NET0131  ;
	input \configuration_pci_err_addr_reg[24]/NET0131  ;
	input \configuration_pci_err_addr_reg[25]/NET0131  ;
	input \configuration_pci_err_addr_reg[26]/NET0131  ;
	input \configuration_pci_err_addr_reg[27]/NET0131  ;
	input \configuration_pci_err_addr_reg[28]/NET0131  ;
	input \configuration_pci_err_addr_reg[29]/NET0131  ;
	input \configuration_pci_err_addr_reg[2]/NET0131  ;
	input \configuration_pci_err_addr_reg[30]/NET0131  ;
	input \configuration_pci_err_addr_reg[31]/NET0131  ;
	input \configuration_pci_err_addr_reg[3]/NET0131  ;
	input \configuration_pci_err_addr_reg[4]/NET0131  ;
	input \configuration_pci_err_addr_reg[5]/NET0131  ;
	input \configuration_pci_err_addr_reg[6]/NET0131  ;
	input \configuration_pci_err_addr_reg[7]/NET0131  ;
	input \configuration_pci_err_addr_reg[8]/NET0131  ;
	input \configuration_pci_err_addr_reg[9]/NET0131  ;
	input \configuration_pci_err_cs_bit0_reg/NET0131  ;
	input \configuration_pci_err_cs_bit10_reg/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[24]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[25]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[26]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[27]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[28]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[29]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[30]/NET0131  ;
	input \configuration_pci_err_cs_bit31_24_reg[31]/NET0131  ;
	input \configuration_pci_err_cs_bit8_reg/NET0131  ;
	input \configuration_pci_err_data_reg[0]/NET0131  ;
	input \configuration_pci_err_data_reg[10]/NET0131  ;
	input \configuration_pci_err_data_reg[11]/NET0131  ;
	input \configuration_pci_err_data_reg[12]/NET0131  ;
	input \configuration_pci_err_data_reg[13]/NET0131  ;
	input \configuration_pci_err_data_reg[14]/NET0131  ;
	input \configuration_pci_err_data_reg[15]/NET0131  ;
	input \configuration_pci_err_data_reg[16]/NET0131  ;
	input \configuration_pci_err_data_reg[17]/NET0131  ;
	input \configuration_pci_err_data_reg[18]/NET0131  ;
	input \configuration_pci_err_data_reg[19]/NET0131  ;
	input \configuration_pci_err_data_reg[1]/NET0131  ;
	input \configuration_pci_err_data_reg[20]/NET0131  ;
	input \configuration_pci_err_data_reg[21]/NET0131  ;
	input \configuration_pci_err_data_reg[22]/NET0131  ;
	input \configuration_pci_err_data_reg[23]/NET0131  ;
	input \configuration_pci_err_data_reg[24]/NET0131  ;
	input \configuration_pci_err_data_reg[25]/NET0131  ;
	input \configuration_pci_err_data_reg[26]/NET0131  ;
	input \configuration_pci_err_data_reg[27]/NET0131  ;
	input \configuration_pci_err_data_reg[28]/NET0131  ;
	input \configuration_pci_err_data_reg[29]/NET0131  ;
	input \configuration_pci_err_data_reg[2]/NET0131  ;
	input \configuration_pci_err_data_reg[30]/NET0131  ;
	input \configuration_pci_err_data_reg[31]/NET0131  ;
	input \configuration_pci_err_data_reg[3]/NET0131  ;
	input \configuration_pci_err_data_reg[4]/NET0131  ;
	input \configuration_pci_err_data_reg[5]/NET0131  ;
	input \configuration_pci_err_data_reg[6]/NET0131  ;
	input \configuration_pci_err_data_reg[7]/NET0131  ;
	input \configuration_pci_err_data_reg[8]/NET0131  ;
	input \configuration_pci_err_data_reg[9]/NET0131  ;
	input \configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131  ;
	input \configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131  ;
	input \configuration_pci_ta1_reg[10]/NET0131  ;
	input \configuration_pci_ta1_reg[11]/NET0131  ;
	input \configuration_pci_ta1_reg[12]/NET0131  ;
	input \configuration_pci_ta1_reg[13]/NET0131  ;
	input \configuration_pci_ta1_reg[14]/NET0131  ;
	input \configuration_pci_ta1_reg[15]/NET0131  ;
	input \configuration_pci_ta1_reg[16]/NET0131  ;
	input \configuration_pci_ta1_reg[17]/NET0131  ;
	input \configuration_pci_ta1_reg[18]/NET0131  ;
	input \configuration_pci_ta1_reg[19]/NET0131  ;
	input \configuration_pci_ta1_reg[20]/NET0131  ;
	input \configuration_pci_ta1_reg[21]/NET0131  ;
	input \configuration_pci_ta1_reg[22]/NET0131  ;
	input \configuration_pci_ta1_reg[23]/NET0131  ;
	input \configuration_pci_ta1_reg[24]/NET0131  ;
	input \configuration_pci_ta1_reg[25]/NET0131  ;
	input \configuration_pci_ta1_reg[26]/NET0131  ;
	input \configuration_pci_ta1_reg[27]/NET0131  ;
	input \configuration_pci_ta1_reg[28]/NET0131  ;
	input \configuration_pci_ta1_reg[29]/NET0131  ;
	input \configuration_pci_ta1_reg[30]/NET0131  ;
	input \configuration_pci_ta1_reg[31]/NET0131  ;
	input \configuration_pci_ta1_reg[8]/NET0131  ;
	input \configuration_pci_ta1_reg[9]/NET0131  ;
	input \configuration_rst_inactive_reg/NET0131  ;
	input \configuration_set_isr_bit2_reg/NET0131  ;
	input \configuration_set_pci_err_cs_bit8_reg/NET0131  ;
	input \configuration_status_bit15_11_reg[11]/NET0131  ;
	input \configuration_status_bit15_11_reg[12]/NET0131  ;
	input \configuration_status_bit15_11_reg[13]/NET0131  ;
	input \configuration_status_bit15_11_reg[14]/NET0131  ;
	input \configuration_status_bit15_11_reg[15]/NET0131  ;
	input \configuration_status_bit8_reg/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131  ;
	input \configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131  ;
	input \configuration_sync_command_bit_reg/NET0131  ;
	input \configuration_sync_isr_2_del_bit_reg/NET0131  ;
	input \configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131  ;
	input \configuration_sync_isr_2_delayed_del_bit_reg/NET0131  ;
	input \configuration_sync_isr_2_sync_bckp_bit_reg/NET0131  ;
	input \configuration_sync_isr_2_sync_del_bit_reg/NET0131  ;
	input \configuration_sync_pci_err_cs_8_del_bit_reg/NET0131  ;
	input \configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131  ;
	input \configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131  ;
	input \configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131  ;
	input \configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131  ;
	input \configuration_wb_am1_reg[31]/NET0131  ;
	input \configuration_wb_am2_reg[31]/NET0131  ;
	input \configuration_wb_ba1_bit0_reg/NET0131  ;
	input \configuration_wb_ba1_bit31_12_reg[31]/NET0131  ;
	input \configuration_wb_ba2_bit0_reg/NET0131  ;
	input \configuration_wb_ba2_bit31_12_reg[31]/NET0131  ;
	input \configuration_wb_err_addr_reg[0]/NET0131  ;
	input \configuration_wb_err_addr_reg[10]/NET0131  ;
	input \configuration_wb_err_addr_reg[11]/NET0131  ;
	input \configuration_wb_err_addr_reg[12]/NET0131  ;
	input \configuration_wb_err_addr_reg[13]/NET0131  ;
	input \configuration_wb_err_addr_reg[14]/NET0131  ;
	input \configuration_wb_err_addr_reg[15]/NET0131  ;
	input \configuration_wb_err_addr_reg[16]/NET0131  ;
	input \configuration_wb_err_addr_reg[17]/NET0131  ;
	input \configuration_wb_err_addr_reg[18]/NET0131  ;
	input \configuration_wb_err_addr_reg[19]/NET0131  ;
	input \configuration_wb_err_addr_reg[1]/NET0131  ;
	input \configuration_wb_err_addr_reg[20]/NET0131  ;
	input \configuration_wb_err_addr_reg[21]/NET0131  ;
	input \configuration_wb_err_addr_reg[22]/NET0131  ;
	input \configuration_wb_err_addr_reg[23]/NET0131  ;
	input \configuration_wb_err_addr_reg[24]/NET0131  ;
	input \configuration_wb_err_addr_reg[25]/NET0131  ;
	input \configuration_wb_err_addr_reg[26]/NET0131  ;
	input \configuration_wb_err_addr_reg[27]/NET0131  ;
	input \configuration_wb_err_addr_reg[28]/NET0131  ;
	input \configuration_wb_err_addr_reg[29]/NET0131  ;
	input \configuration_wb_err_addr_reg[2]/NET0131  ;
	input \configuration_wb_err_addr_reg[30]/NET0131  ;
	input \configuration_wb_err_addr_reg[31]/NET0131  ;
	input \configuration_wb_err_addr_reg[3]/NET0131  ;
	input \configuration_wb_err_addr_reg[4]/NET0131  ;
	input \configuration_wb_err_addr_reg[5]/NET0131  ;
	input \configuration_wb_err_addr_reg[6]/NET0131  ;
	input \configuration_wb_err_addr_reg[7]/NET0131  ;
	input \configuration_wb_err_addr_reg[8]/NET0131  ;
	input \configuration_wb_err_addr_reg[9]/NET0131  ;
	input \configuration_wb_err_cs_bit0_reg/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[24]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[25]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[26]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[27]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[28]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[29]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[30]/NET0131  ;
	input \configuration_wb_err_cs_bit31_24_reg[31]/NET0131  ;
	input \configuration_wb_err_cs_bit8_reg/NET0131  ;
	input \configuration_wb_err_cs_bit9_reg/NET0131  ;
	input \configuration_wb_err_data_reg[0]/NET0131  ;
	input \configuration_wb_err_data_reg[10]/NET0131  ;
	input \configuration_wb_err_data_reg[11]/NET0131  ;
	input \configuration_wb_err_data_reg[12]/NET0131  ;
	input \configuration_wb_err_data_reg[13]/NET0131  ;
	input \configuration_wb_err_data_reg[14]/NET0131  ;
	input \configuration_wb_err_data_reg[15]/NET0131  ;
	input \configuration_wb_err_data_reg[16]/NET0131  ;
	input \configuration_wb_err_data_reg[17]/NET0131  ;
	input \configuration_wb_err_data_reg[18]/NET0131  ;
	input \configuration_wb_err_data_reg[19]/NET0131  ;
	input \configuration_wb_err_data_reg[1]/NET0131  ;
	input \configuration_wb_err_data_reg[20]/NET0131  ;
	input \configuration_wb_err_data_reg[21]/NET0131  ;
	input \configuration_wb_err_data_reg[22]/NET0131  ;
	input \configuration_wb_err_data_reg[23]/NET0131  ;
	input \configuration_wb_err_data_reg[24]/NET0131  ;
	input \configuration_wb_err_data_reg[25]/NET0131  ;
	input \configuration_wb_err_data_reg[26]/NET0131  ;
	input \configuration_wb_err_data_reg[27]/NET0131  ;
	input \configuration_wb_err_data_reg[28]/NET0131  ;
	input \configuration_wb_err_data_reg[29]/NET0131  ;
	input \configuration_wb_err_data_reg[2]/NET0131  ;
	input \configuration_wb_err_data_reg[30]/NET0131  ;
	input \configuration_wb_err_data_reg[31]/NET0131  ;
	input \configuration_wb_err_data_reg[3]/NET0131  ;
	input \configuration_wb_err_data_reg[4]/NET0131  ;
	input \configuration_wb_err_data_reg[5]/NET0131  ;
	input \configuration_wb_err_data_reg[6]/NET0131  ;
	input \configuration_wb_err_data_reg[7]/NET0131  ;
	input \configuration_wb_err_data_reg[8]/NET0131  ;
	input \configuration_wb_err_data_reg[9]/NET0131  ;
	input \configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131  ;
	input \configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131  ;
	input \configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131  ;
	input \configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131  ;
	input \configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131  ;
	input \configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131  ;
	input \configuration_wb_init_complete_out_reg/NET0131  ;
	input \configuration_wb_ta1_reg[31]/NET0131  ;
	input \configuration_wb_ta2_reg[31]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131  ;
	input \i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[0]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[10]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[11]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[12]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[13]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[14]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[15]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[16]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[17]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[18]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[19]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[1]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[20]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[21]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[22]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[23]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[24]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[25]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[26]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[27]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[28]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[29]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[2]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[30]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[31]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[3]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[4]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[5]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[6]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[7]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[8]/NET0131  ;
	input \input_register_pci_ad_reg_out_reg[9]/NET0131  ;
	input \input_register_pci_cbe_reg_out_reg[0]/NET0131  ;
	input \input_register_pci_cbe_reg_out_reg[1]/NET0131  ;
	input \input_register_pci_cbe_reg_out_reg[2]/NET0131  ;
	input \input_register_pci_cbe_reg_out_reg[3]/NET0131  ;
	input \input_register_pci_devsel_reg_out_reg/NET0131  ;
	input \input_register_pci_frame_reg_out_reg/NET0131  ;
	input \input_register_pci_idsel_reg_out_reg/NET0131  ;
	input \input_register_pci_irdy_reg_out_reg/NET0131  ;
	input \input_register_pci_stop_reg_out_reg/NET0131  ;
	input \input_register_pci_trdy_reg_out_reg/NET0131  ;
	input \output_backup_ad_out_reg[0]/NET0131  ;
	input \output_backup_ad_out_reg[10]/NET0131  ;
	input \output_backup_ad_out_reg[11]/NET0131  ;
	input \output_backup_ad_out_reg[12]/NET0131  ;
	input \output_backup_ad_out_reg[13]/NET0131  ;
	input \output_backup_ad_out_reg[14]/NET0131  ;
	input \output_backup_ad_out_reg[15]/NET0131  ;
	input \output_backup_ad_out_reg[16]/NET0131  ;
	input \output_backup_ad_out_reg[17]/NET0131  ;
	input \output_backup_ad_out_reg[18]/NET0131  ;
	input \output_backup_ad_out_reg[19]/NET0131  ;
	input \output_backup_ad_out_reg[1]/NET0131  ;
	input \output_backup_ad_out_reg[20]/NET0131  ;
	input \output_backup_ad_out_reg[21]/NET0131  ;
	input \output_backup_ad_out_reg[22]/NET0131  ;
	input \output_backup_ad_out_reg[23]/NET0131  ;
	input \output_backup_ad_out_reg[24]/NET0131  ;
	input \output_backup_ad_out_reg[25]/NET0131  ;
	input \output_backup_ad_out_reg[26]/NET0131  ;
	input \output_backup_ad_out_reg[27]/NET0131  ;
	input \output_backup_ad_out_reg[28]/NET0131  ;
	input \output_backup_ad_out_reg[29]/NET0131  ;
	input \output_backup_ad_out_reg[2]/NET0131  ;
	input \output_backup_ad_out_reg[30]/NET0131  ;
	input \output_backup_ad_out_reg[31]/NET0131  ;
	input \output_backup_ad_out_reg[3]/NET0131  ;
	input \output_backup_ad_out_reg[4]/NET0131  ;
	input \output_backup_ad_out_reg[5]/NET0131  ;
	input \output_backup_ad_out_reg[6]/NET0131  ;
	input \output_backup_ad_out_reg[7]/NET0131  ;
	input \output_backup_ad_out_reg[8]/NET0131  ;
	input \output_backup_ad_out_reg[9]/NET0131  ;
	input \output_backup_cbe_en_out_reg/NET0131  ;
	input \output_backup_cbe_out_reg[0]/NET0131  ;
	input \output_backup_cbe_out_reg[1]/NET0131  ;
	input \output_backup_cbe_out_reg[2]/NET0131  ;
	input \output_backup_cbe_out_reg[3]/NET0131  ;
	input \output_backup_devsel_out_reg/NET0131  ;
	input \output_backup_frame_en_out_reg/NET0131  ;
	input \output_backup_frame_out_reg/NET0131  ;
	input \output_backup_irdy_en_out_reg/NET0131  ;
	input \output_backup_irdy_out_reg/NET0131  ;
	input \output_backup_mas_ad_en_out_reg/NET0131  ;
	input \output_backup_par_en_out_reg/NET0131  ;
	input \output_backup_par_out_reg/NET0131  ;
	input \output_backup_perr_en_out_reg/NET0131  ;
	input \output_backup_perr_out_reg/NET0131  ;
	input \output_backup_serr_en_out_reg/NET0131  ;
	input \output_backup_serr_out_reg/NET0131  ;
	input \output_backup_stop_out_reg/NET0131  ;
	input \output_backup_tar_ad_en_out_reg/NET0131  ;
	input \output_backup_trdy_en_out_reg/NET0131  ;
	input \output_backup_trdy_out_reg/NET0131  ;
	input \parity_checker_check_for_serr_on_second_reg/NET0131  ;
	input \parity_checker_check_perr_reg/NET0131  ;
	input \parity_checker_frame_dec2_reg/NET0131  ;
	input \parity_checker_master_perr_report_reg/NET0131  ;
	input \parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131  ;
	input \parity_checker_perr_sampled_reg/NET0131  ;
	input \pci_cbe_i[0]_pad  ;
	input \pci_cbe_i[1]_pad  ;
	input \pci_cbe_i[2]_pad  ;
	input \pci_cbe_i[3]_pad  ;
	input pci_devsel_i_pad ;
	input pci_frame_i_pad ;
	input pci_frame_o_pad ;
	input pci_gnt_i_pad ;
	input pci_irdy_i_pad ;
	input pci_par_i_pad ;
	input pci_perr_i_pad ;
	input pci_rst_i_pad ;
	input pci_stop_i_pad ;
	input \pci_target_unit_del_sync_addr_out_reg[0]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[10]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[11]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[12]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[13]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[14]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[15]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[16]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[17]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[18]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[19]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[1]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[20]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[21]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[22]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[23]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[24]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[25]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[26]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[27]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[28]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[29]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[2]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[30]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[31]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[3]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[4]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[5]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[6]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[7]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[8]/NET0131  ;
	input \pci_target_unit_del_sync_addr_out_reg[9]/NET0131  ;
	input \pci_target_unit_del_sync_bc_out_reg[0]/NET0131  ;
	input \pci_target_unit_del_sync_bc_out_reg[1]/NET0131  ;
	input \pci_target_unit_del_sync_bc_out_reg[2]/NET0131  ;
	input \pci_target_unit_del_sync_bc_out_reg[3]/NET0131  ;
	input \pci_target_unit_del_sync_be_out_reg[0]/NET0131  ;
	input \pci_target_unit_del_sync_be_out_reg[1]/NET0131  ;
	input \pci_target_unit_del_sync_be_out_reg[2]/NET0131  ;
	input \pci_target_unit_del_sync_be_out_reg[3]/NET0131  ;
	input \pci_target_unit_del_sync_burst_out_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_comp_pending_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131  ;
	input \pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131  ;
	input \pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_flush_out_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_req_pending_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131  ;
	input \pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  ;
	input \pci_target_unit_del_sync_req_comp_pending_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_done_reg_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_req_pending_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131  ;
	input \pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_inGreyCount_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_outGreyCount_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_outGreyCount_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001  ;
	input \pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001  ;
	input \pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001  ;
	input \pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131  ;
	input \pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131  ;
	input \pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131  ;
	input \pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131  ;
	input \pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131  ;
	input \pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131  ;
	input \pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131  ;
	input \pci_target_unit_pci_target_if_same_read_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_if_target_rd_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_backoff_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131  ;
	input \pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131  ;
	input \pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131  ;
	input \pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_rd_progress_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_rd_request_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_wr_progress_reg/NET0131  ;
	input \pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_burst_chopped_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_c_state_reg[0]/NET0131  ;
	input \pci_target_unit_wishbone_master_c_state_reg[1]/NET0131  ;
	input \pci_target_unit_wishbone_master_c_state_reg[2]/NET0131  ;
	input \pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_read_bound_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_read_count_reg[0]/NET0131  ;
	input \pci_target_unit_wishbone_master_read_count_reg[1]/NET0131  ;
	input \pci_target_unit_wishbone_master_read_count_reg[2]/NET0131  ;
	input \pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_retried_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131  ;
	input \pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131  ;
	input \pci_target_unit_wishbone_master_w_attempt_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131  ;
	input \pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131  ;
	input pci_trdy_i_pad ;
	input wb_int_i_pad ;
	input wbm_ack_i_pad ;
	input \wbm_adr_o[0]_pad  ;
	input \wbm_adr_o[10]_pad  ;
	input \wbm_adr_o[11]_pad  ;
	input \wbm_adr_o[12]_pad  ;
	input \wbm_adr_o[13]_pad  ;
	input \wbm_adr_o[14]_pad  ;
	input \wbm_adr_o[15]_pad  ;
	input \wbm_adr_o[16]_pad  ;
	input \wbm_adr_o[17]_pad  ;
	input \wbm_adr_o[18]_pad  ;
	input \wbm_adr_o[19]_pad  ;
	input \wbm_adr_o[1]_pad  ;
	input \wbm_adr_o[20]_pad  ;
	input \wbm_adr_o[21]_pad  ;
	input \wbm_adr_o[22]_pad  ;
	input \wbm_adr_o[23]_pad  ;
	input \wbm_adr_o[24]_pad  ;
	input \wbm_adr_o[25]_pad  ;
	input \wbm_adr_o[26]_pad  ;
	input \wbm_adr_o[27]_pad  ;
	input \wbm_adr_o[28]_pad  ;
	input \wbm_adr_o[29]_pad  ;
	input \wbm_adr_o[2]_pad  ;
	input \wbm_adr_o[30]_pad  ;
	input \wbm_adr_o[31]_pad  ;
	input \wbm_adr_o[3]_pad  ;
	input \wbm_adr_o[4]_pad  ;
	input \wbm_adr_o[5]_pad  ;
	input \wbm_adr_o[6]_pad  ;
	input \wbm_adr_o[7]_pad  ;
	input \wbm_adr_o[8]_pad  ;
	input \wbm_adr_o[9]_pad  ;
	input \wbm_cti_o[0]_pad  ;
	input \wbm_dat_o[0]_pad  ;
	input \wbm_dat_o[10]_pad  ;
	input \wbm_dat_o[11]_pad  ;
	input \wbm_dat_o[12]_pad  ;
	input \wbm_dat_o[13]_pad  ;
	input \wbm_dat_o[14]_pad  ;
	input \wbm_dat_o[15]_pad  ;
	input \wbm_dat_o[16]_pad  ;
	input \wbm_dat_o[17]_pad  ;
	input \wbm_dat_o[18]_pad  ;
	input \wbm_dat_o[19]_pad  ;
	input \wbm_dat_o[1]_pad  ;
	input \wbm_dat_o[20]_pad  ;
	input \wbm_dat_o[21]_pad  ;
	input \wbm_dat_o[22]_pad  ;
	input \wbm_dat_o[23]_pad  ;
	input \wbm_dat_o[24]_pad  ;
	input \wbm_dat_o[25]_pad  ;
	input \wbm_dat_o[26]_pad  ;
	input \wbm_dat_o[27]_pad  ;
	input \wbm_dat_o[28]_pad  ;
	input \wbm_dat_o[29]_pad  ;
	input \wbm_dat_o[2]_pad  ;
	input \wbm_dat_o[30]_pad  ;
	input \wbm_dat_o[31]_pad  ;
	input \wbm_dat_o[3]_pad  ;
	input \wbm_dat_o[4]_pad  ;
	input \wbm_dat_o[5]_pad  ;
	input \wbm_dat_o[6]_pad  ;
	input \wbm_dat_o[7]_pad  ;
	input \wbm_dat_o[8]_pad  ;
	input \wbm_dat_o[9]_pad  ;
	input wbm_err_i_pad ;
	input wbm_rty_i_pad ;
	input \wbm_sel_o[0]_pad  ;
	input \wbm_sel_o[1]_pad  ;
	input \wbm_sel_o[2]_pad  ;
	input \wbm_sel_o[3]_pad  ;
	input \wbs_adr_i[10]_pad  ;
	input \wbs_adr_i[11]_pad  ;
	input \wbs_adr_i[12]_pad  ;
	input \wbs_adr_i[13]_pad  ;
	input \wbs_adr_i[14]_pad  ;
	input \wbs_adr_i[15]_pad  ;
	input \wbs_adr_i[16]_pad  ;
	input \wbs_adr_i[17]_pad  ;
	input \wbs_adr_i[18]_pad  ;
	input \wbs_adr_i[19]_pad  ;
	input \wbs_adr_i[20]_pad  ;
	input \wbs_adr_i[21]_pad  ;
	input \wbs_adr_i[22]_pad  ;
	input \wbs_adr_i[23]_pad  ;
	input \wbs_adr_i[24]_pad  ;
	input \wbs_adr_i[25]_pad  ;
	input \wbs_adr_i[26]_pad  ;
	input \wbs_adr_i[27]_pad  ;
	input \wbs_adr_i[28]_pad  ;
	input \wbs_adr_i[29]_pad  ;
	input \wbs_adr_i[2]_pad  ;
	input \wbs_adr_i[30]_pad  ;
	input \wbs_adr_i[31]_pad  ;
	input \wbs_adr_i[3]_pad  ;
	input \wbs_adr_i[4]_pad  ;
	input \wbs_adr_i[5]_pad  ;
	input \wbs_adr_i[6]_pad  ;
	input \wbs_adr_i[7]_pad  ;
	input \wbs_adr_i[8]_pad  ;
	input \wbs_adr_i[9]_pad  ;
	input \wbs_bte_i[0]_pad  ;
	input \wbs_bte_i[1]_pad  ;
	input \wbs_cti_i[0]_pad  ;
	input \wbs_cti_i[1]_pad  ;
	input \wbs_cti_i[2]_pad  ;
	input wbs_cyc_i_pad ;
	input wbs_stb_i_pad ;
	input wbs_we_i_pad ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131  ;
	input \wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131  ;
	input \wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_del_sync_burst_out_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131  ;
	input \wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001  ;
	input \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131  ;
	input \wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131  ;
	input \wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_map_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131  ;
	input \wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131  ;
	output \configuration_init_complete_reg/P0001  ;
	output \configuration_interrupt_out_reg/P0001  ;
	output \g21/_0_  ;
	output \g52241/_0_  ;
	output \g52244/_0_  ;
	output \g52348/_0_  ;
	output \g52349/_0_  ;
	output \g52350/_0_  ;
	output \g52351/_0_  ;
	output \g52352/_0_  ;
	output \g52390/_0_  ;
	output \g52391/_0_  ;
	output \g52393/_3_  ;
	output \g52394/_3_  ;
	output \g52395/_3_  ;
	output \g52396/_3_  ;
	output \g52397/_3_  ;
	output \g52398/_3_  ;
	output \g52399/_3_  ;
	output \g52400/_3_  ;
	output \g52401/_3_  ;
	output \g52402/_3_  ;
	output \g52403/_3_  ;
	output \g52404/_3_  ;
	output \g52405/_3_  ;
	output \g52406/_0_  ;
	output \g52408/_0_  ;
	output \g52409/_0_  ;
	output \g52410/_0_  ;
	output \g52411/_0_  ;
	output \g52412/_0_  ;
	output \g52413/_0_  ;
	output \g52414/_0_  ;
	output \g52415/_0_  ;
	output \g52416/_0_  ;
	output \g52417/_0_  ;
	output \g52418/_0_  ;
	output \g52419/_0_  ;
	output \g52421/_0_  ;
	output \g52422/_0_  ;
	output \g52423/_0_  ;
	output \g52424/_0_  ;
	output \g52425/_0_  ;
	output \g52426/_0_  ;
	output \g52427/_0_  ;
	output \g52428/_0_  ;
	output \g52429/_0_  ;
	output \g52430/_0_  ;
	output \g52431/_0_  ;
	output \g52432/_0_  ;
	output \g52433/_0_  ;
	output \g52434/_0_  ;
	output \g52435/_0_  ;
	output \g52436/_0_  ;
	output \g52437/_0_  ;
	output \g52439/_3_  ;
	output \g52440/_3_  ;
	output \g52441/_3_  ;
	output \g52442/_3_  ;
	output \g52443/_3_  ;
	output \g52444/_3_  ;
	output \g52445/_3_  ;
	output \g52446/_3_  ;
	output \g52447/_3_  ;
	output \g52448/_3_  ;
	output \g52449/_3_  ;
	output \g52450/_3_  ;
	output \g52451/_3_  ;
	output \g52452/_3_  ;
	output \g52453/_3_  ;
	output \g52454/_3_  ;
	output \g52455/_3_  ;
	output \g52456/_3_  ;
	output \g52457/_3_  ;
	output \g52458/_3_  ;
	output \g52459/_3_  ;
	output \g52460/_3_  ;
	output \g52461/_3_  ;
	output \g52462/_3_  ;
	output \g52463/_3_  ;
	output \g52464/_3_  ;
	output \g52465/_3_  ;
	output \g52466/_3_  ;
	output \g52467/_3_  ;
	output \g52468/_3_  ;
	output \g52469/_3_  ;
	output \g52470/_3_  ;
	output \g52471/_3_  ;
	output \g52472/_3_  ;
	output \g52473/_3_  ;
	output \g52474/_3_  ;
	output \g52475/_3_  ;
	output \g52476/_3_  ;
	output \g52477/_3_  ;
	output \g52478/_3_  ;
	output \g52479/_3_  ;
	output \g52480/_3_  ;
	output \g52481/_3_  ;
	output \g52482/_3_  ;
	output \g52483/_3_  ;
	output \g52484/_3_  ;
	output \g52485/_3_  ;
	output \g52499/_0_  ;
	output \g52500/_0_  ;
	output \g52501/_0_  ;
	output \g52547/_0_  ;
	output \g52550/_0_  ;
	output \g52553/_0_  ;
	output \g52675/_0__syn_2  ;
	output \g52714/_0_  ;
	output \g52715/_0_  ;
	output \g52716/_0_  ;
	output \g52717/_0_  ;
	output \g52718/_0_  ;
	output \g52720/_0_  ;
	output \g52865/_0_  ;
	output \g52867/_0_  ;
	output \g52867/_1_  ;
	output \g52868/_0_  ;
	output \g52871/_2_  ;
	output \g52897/_0_  ;
	output \g52898/_0_  ;
	output \g52899/_0_  ;
	output \g52900/_0_  ;
	output \g52901/_0_  ;
	output \g52902/_0_  ;
	output \g52903/_0_  ;
	output \g52904/_0_  ;
	output \g52905/_0_  ;
	output \g52906/_0_  ;
	output \g52907/_0_  ;
	output \g52908/_0_  ;
	output \g52909/_0_  ;
	output \g52910/_0_  ;
	output \g52911/_0_  ;
	output \g52912/_0_  ;
	output \g52913/_0_  ;
	output \g52914/_0_  ;
	output \g52915/_0_  ;
	output \g52916/_0_  ;
	output \g52917/_0_  ;
	output \g52918/_0_  ;
	output \g52920/_0_  ;
	output \g52921/_0_  ;
	output \g52922/_0_  ;
	output \g52923/_0_  ;
	output \g52924/_0_  ;
	output \g52925/_0_  ;
	output \g52948/_0_  ;
	output \g52958/_0_  ;
	output \g52959/_0_  ;
	output \g52960/_0_  ;
	output \g52961/_0_  ;
	output \g52962/_0_  ;
	output \g52963/_0_  ;
	output \g52965/_0_  ;
	output \g52966/_0_  ;
	output \g52969/_0_  ;
	output \g52970/_0_  ;
	output \g52971/_0_  ;
	output \g52972/_0_  ;
	output \g52973/_0_  ;
	output \g52975/_0_  ;
	output \g52976/_0_  ;
	output \g52977/_0_  ;
	output \g52978/_0_  ;
	output \g52979/_0_  ;
	output \g52980/_0_  ;
	output \g52981/_0_  ;
	output \g52982/_0_  ;
	output \g52983/_0_  ;
	output \g52984/_0_  ;
	output \g52985/_0_  ;
	output \g52986/_0_  ;
	output \g52988/_0_  ;
	output \g52990/_0_  ;
	output \g52991/_0_  ;
	output \g52993/_0_  ;
	output \g52994/_0_  ;
	output \g52996/_0_  ;
	output \g52997/_0_  ;
	output \g53068/_0_  ;
	output \g53085/_0_  ;
	output \g53086/_0_  ;
	output \g53088/_0_  ;
	output \g53089/_0_  ;
	output \g53090/_0_  ;
	output \g53091/_0_  ;
	output \g53096/_0_  ;
	output \g53123/_0_  ;
	output \g53124/_0_  ;
	output \g53137/_0_  ;
	output \g53137/_1_  ;
	output \g53145/_0_  ;
	output \g53146/_0_  ;
	output \g53147/_0_  ;
	output \g53870/_0_  ;
	output \g53871/_0_  ;
	output \g53872/_0_  ;
	output \g53873/_0_  ;
	output \g53874/_0_  ;
	output \g53875/_0_  ;
	output \g53876/_0_  ;
	output \g53877/_0_  ;
	output \g53878/_0_  ;
	output \g53879/_0_  ;
	output \g53880/_0_  ;
	output \g53881/_0_  ;
	output \g53882/_0_  ;
	output \g53883/_0_  ;
	output \g53884/_0_  ;
	output \g53885/_0_  ;
	output \g53886/_0_  ;
	output \g53887/_0_  ;
	output \g53888/_0_  ;
	output \g53889/_0_  ;
	output \g53890/_3_  ;
	output \g53897/_3_  ;
	output \g53935/_3_  ;
	output \g53936/_3_  ;
	output \g53937/_3_  ;
	output \g53938/_3_  ;
	output \g53939/_3_  ;
	output \g53940/_3_  ;
	output \g53941/_3_  ;
	output \g53942/_3_  ;
	output \g54022/_0_  ;
	output \g54160/_3_  ;
	output \g54163/_3_  ;
	output \g54166/_3_  ;
	output \g54167/_2_  ;
	output \g54168/_3_  ;
	output \g54169/_3_  ;
	output \g54170/_3_  ;
	output \g54171/_2_  ;
	output \g54172/_3_  ;
	output \g54173/_3_  ;
	output \g54204/_2_  ;
	output \g54205/_2_  ;
	output \g54206/_2_  ;
	output \g54207/_2_  ;
	output \g54208/_2_  ;
	output \g54209/_2_  ;
	output \g54210/_2_  ;
	output \g54211/_2_  ;
	output \g54212/_2_  ;
	output \g54213/_2_  ;
	output \g54214/_2_  ;
	output \g54215/_2_  ;
	output \g54216/_2_  ;
	output \g54217/_2_  ;
	output \g54218/_2_  ;
	output \g54219/_2_  ;
	output \g54220/_2_  ;
	output \g54221/_2_  ;
	output \g54222/_2_  ;
	output \g54223/_2_  ;
	output \g54224/_2_  ;
	output \g54225/_2_  ;
	output \g54226/_2_  ;
	output \g54227/_2_  ;
	output \g54228/_2_  ;
	output \g54229/_2_  ;
	output \g54230/_2_  ;
	output \g54231/_2_  ;
	output \g54232/_2_  ;
	output \g54233/_2_  ;
	output \g54267/_0_  ;
	output \g54268/_0_  ;
	output \g54269/_0_  ;
	output \g54270/_0_  ;
	output \g54271/_0_  ;
	output \g54272/_0_  ;
	output \g54273/_0_  ;
	output \g54274/_0_  ;
	output \g54275/_0_  ;
	output \g54276/_0_  ;
	output \g54278/_0_  ;
	output \g54279/_0_  ;
	output \g54280/_0_  ;
	output \g54281/_0_  ;
	output \g54282/_0_  ;
	output \g54283/_0_  ;
	output \g54284/_0_  ;
	output \g54285/_0_  ;
	output \g54286/_0_  ;
	output \g54287/_0_  ;
	output \g54288/_0_  ;
	output \g54289/_0_  ;
	output \g54290/_0_  ;
	output \g54291/_0_  ;
	output \g54292/_0_  ;
	output \g54293/_0_  ;
	output \g54294/_0_  ;
	output \g54296/_0_  ;
	output \g54297/_0_  ;
	output \g54298/_0_  ;
	output \g54299/_0_  ;
	output \g54300/_0_  ;
	output \g54301/_0_  ;
	output \g54302/_0_  ;
	output \g54303/_0_  ;
	output \g54329/_0_  ;
	output \g54453/_0_  ;
	output \g54466/_0_  ;
	output \g54470/_0_  ;
	output \g54470/_1_  ;
	output \g54496/_0_  ;
	output \g54597/_0_  ;
	output \g54628/_0_  ;
	output \g54629/_0_  ;
	output \g54630/_0_  ;
	output \g54631/_0_  ;
	output \g54632/_0_  ;
	output \g54633/_0_  ;
	output \g54634/_0_  ;
	output \g54635/_0_  ;
	output \g54636/_0_  ;
	output \g54638/_0_  ;
	output \g54639/_0_  ;
	output \g54640/_0_  ;
	output \g54641/_0_  ;
	output \g54642/_0_  ;
	output \g54643/_0_  ;
	output \g54645/_0_  ;
	output \g54646/_0_  ;
	output \g54647/_0_  ;
	output \g54648/_0_  ;
	output \g54649/_0_  ;
	output \g54650/_0_  ;
	output \g54651/_0_  ;
	output \g54652/_0_  ;
	output \g54653/_0_  ;
	output \g54654/_0_  ;
	output \g54655/_0_  ;
	output \g54656/_0_  ;
	output \g54657/_0_  ;
	output \g54658/_0_  ;
	output \g54659/_0_  ;
	output \g54660/_0_  ;
	output \g54661/_0_  ;
	output \g54662/_0_  ;
	output \g54663/_0_  ;
	output \g54664/_0_  ;
	output \g54669/_0_  ;
	output \g54832/_0_  ;
	output \g54833/_0_  ;
	output \g54867/_0_  ;
	output \g54868/_0_  ;
	output \g54869/_0_  ;
	output \g54870/_0_  ;
	output \g54871/_0_  ;
	output \g54872/_0_  ;
	output \g54873/_0_  ;
	output \g54874/_0_  ;
	output \g54875/_0_  ;
	output \g54876/_0_  ;
	output \g54877/_0_  ;
	output \g54878/_0_  ;
	output \g54879/_0_  ;
	output \g54880/_0_  ;
	output \g54881/_0_  ;
	output \g54882/_0_  ;
	output \g54883/_0_  ;
	output \g54884/_0_  ;
	output \g54885/_0_  ;
	output \g54886/_0_  ;
	output \g54887/_0_  ;
	output \g54888/_0_  ;
	output \g54889/_0_  ;
	output \g54890/_0_  ;
	output \g54891/_0_  ;
	output \g54892/_0_  ;
	output \g54893/_0_  ;
	output \g54894/_0_  ;
	output \g54895/_0_  ;
	output \g54896/_0_  ;
	output \g54897/_0_  ;
	output \g54898/_0_  ;
	output \g54899/_0_  ;
	output \g56438/_0_  ;
	output \g56439/_0_  ;
	output \g56933/_3_  ;
	output \g56934/_3_  ;
	output \g56960/_0_  ;
	output \g56960/_1_  ;
	output \g56961/_3__syn_2  ;
	output \g57019/_0_  ;
	output \g57020/_0_  ;
	output \g57021/_0_  ;
	output \g57022/_0_  ;
	output \g57023/_0_  ;
	output \g57024/_0_  ;
	output \g57025/_0_  ;
	output \g57026/_0_  ;
	output \g57027/_0_  ;
	output \g57028/_0_  ;
	output \g57029/_0_  ;
	output \g57031/_0_  ;
	output \g57032/_0_  ;
	output \g57034/u3_syn_4  ;
	output \g57069/u3_syn_4  ;
	output \g57104/u3_syn_4  ;
	output \g57139/u3_syn_4  ;
	output \g57174/u3_syn_4  ;
	output \g57209/u3_syn_4  ;
	output \g57244/u3_syn_4  ;
	output \g57276/u3_syn_4  ;
	output \g57308/u3_syn_4  ;
	output \g57340/u3_syn_4  ;
	output \g57372/u3_syn_4  ;
	output \g57404/u3_syn_4  ;
	output \g57408/u3_syn_4  ;
	output \g57444/u3_syn_4  ;
	output \g57480/u3_syn_4  ;
	output \g57516/u3_syn_4  ;
	output \g57646/_0_  ;
	output \g57649/_0_  ;
	output \g57779/_3_  ;
	output \g57780/_3_  ;
	output \g57781/_3_  ;
	output \g57782/_3_  ;
	output \g57783/_3_  ;
	output \g57784/_3_  ;
	output \g57785/_3_  ;
	output \g57786/_3_  ;
	output \g57787/_3_  ;
	output \g57788/_3_  ;
	output \g57789/_3_  ;
	output \g57791/_3_  ;
	output \g57795/_3_  ;
	output \g57796/_3_  ;
	output \g57797/_3_  ;
	output \g57798/_3_  ;
	output \g57799/_3_  ;
	output \g57800/_3_  ;
	output \g57801/_3_  ;
	output \g57802/_3_  ;
	output \g57850/_0_  ;
	output \g57852/_0_  ;
	output \g57871/_0_  ;
	output \g57872/_0_  ;
	output \g57873/_0_  ;
	output \g58/_0_  ;
	output \g58490/_0_  ;
	output \g58564/_0_  ;
	output \g58569/_0_  ;
	output \g58571/_0_  ;
	output \g58573/_0_  ;
	output \g58577/_0_  ;
	output \g58578/_0_  ;
	output \g58579/_0_  ;
	output \g58580/_0_  ;
	output \g58583/_0_  ;
	output \g58584/_0_  ;
	output \g58603/_0_  ;
	output \g58611/_3_  ;
	output \g58637/_0_  ;
	output \g58638/_0_  ;
	output \g58639/_0_  ;
	output \g58691/_0_  ;
	output \g58693/_0_  ;
	output \g58696/_0_  ;
	output \g58700/_0_  ;
	output \g58701/_0_  ;
	output \g58708/_1_  ;
	output \g58730/_0_  ;
	output \g58731/_0_  ;
	output \g58732/_0_  ;
	output \g58733/_0_  ;
	output \g58734/_0_  ;
	output \g58735/_0_  ;
	output \g58736/_0_  ;
	output \g58737/_0_  ;
	output \g58738/_0_  ;
	output \g58739/_0_  ;
	output \g58740/_0_  ;
	output \g58741/_1__syn_2  ;
	output \g58748/_0_  ;
	output \g58751/_0_  ;
	output \g58752/_0_  ;
	output \g58753/_0_  ;
	output \g58754/_0_  ;
	output \g58756/_0_  ;
	output \g58767/_3_  ;
	output \g58768/_3_  ;
	output \g58769/_3_  ;
	output \g58770/_3_  ;
	output \g58771/_3_  ;
	output \g58772/_3_  ;
	output \g58773/_3_  ;
	output \g58774/_3_  ;
	output \g58775/_3_  ;
	output \g58776/_3_  ;
	output \g58777/_3_  ;
	output \g58778/_3_  ;
	output \g58779/_3_  ;
	output \g58780/_3_  ;
	output \g58781/_3_  ;
	output \g58782/_3_  ;
	output \g58783/_3_  ;
	output \g58784/_3_  ;
	output \g58785/_3_  ;
	output \g58786/_3_  ;
	output \g58787/_3_  ;
	output \g58788/_3_  ;
	output \g58789/_3_  ;
	output \g58790/_3_  ;
	output \g58791/_3_  ;
	output \g58792/_3_  ;
	output \g58793/_3_  ;
	output \g58794/_3_  ;
	output \g58795/_3_  ;
	output \g58796/_3_  ;
	output \g58797/_3_  ;
	output \g58798/_3_  ;
	output \g58874/_0_  ;
	output \g59064/_1_  ;
	output \g59072/_0_  ;
	output \g59080/_0_  ;
	output \g59083/_0_  ;
	output \g59084/_0_  ;
	output \g59085/_0_  ;
	output \g59088/_0_  ;
	output \g59094/_0_  ;
	output \g59095/_0_  ;
	output \g59126/_3_  ;
	output \g59128/_0_  ;
	output \g59174/_2_  ;
	output \g59180/_0_  ;
	output \g59181/_0_  ;
	output \g59182/_0_  ;
	output \g59190/_0_  ;
	output \g59191/_0_  ;
	output \g59192/_0_  ;
	output \g59204/_0_  ;
	output \g59205/_0_  ;
	output \g59210/_3_  ;
	output \g59213/_0_  ;
	output \g59214/_0_  ;
	output \g59215/_0_  ;
	output \g59216/_0_  ;
	output \g59217/_0_  ;
	output \g59218/_0_  ;
	output \g59219/_0_  ;
	output \g59220/_0_  ;
	output \g59221/_0_  ;
	output \g59222/_0_  ;
	output \g59223/_0_  ;
	output \g59226/_3_  ;
	output \g59232/_00_  ;
	output \g59233/_0_  ;
	output \g59235/_0_  ;
	output \g59236/_0_  ;
	output \g59237/_0_  ;
	output \g59238/_0_  ;
	output \g59318/_0_  ;
	output \g59331/_0_  ;
	output \g59336/_0_  ;
	output \g59351/_0_  ;
	output \g59354/_0_  ;
	output \g59358/_0_  ;
	output \g59363/_0_  ;
	output \g59366/_0_  ;
	output \g59370/u3_syn_4  ;
	output \g59371/u3_syn_4  ;
	output \g59372/u3_syn_4  ;
	output \g59373/u3_syn_4  ;
	output \g59378/u3_syn_4  ;
	output \g59379/u3_syn_4  ;
	output \g59380/u3_syn_4  ;
	output \g59381/u3_syn_4  ;
	output \g59589/_0_  ;
	output \g59655/_0_  ;
	output \g59662/_0_  ;
	output \g59735/_0_  ;
	output \g59739/_0_  ;
	output \g59740/_0_  ;
	output \g59741/_0_  ;
	output \g59742/_0_  ;
	output \g59743/_0_  ;
	output \g59744/_0_  ;
	output \g59745/_0_  ;
	output \g59746/_0_  ;
	output \g59747/_0_  ;
	output \g59748/_0_  ;
	output \g59749/_0_  ;
	output \g59750/_0_  ;
	output \g59751/_0_  ;
	output \g59752/_0_  ;
	output \g59753/_0_  ;
	output \g59754/_0_  ;
	output \g59755/_0_  ;
	output \g59756/_0_  ;
	output \g59757/_0_  ;
	output \g59758/_0_  ;
	output \g59759/_0_  ;
	output \g59760/_0_  ;
	output \g59764/_0_  ;
	output \g59766/_0_  ;
	output \g59774/_0_  ;
	output \g59775/_0_  ;
	output \g59776/_0_  ;
	output \g59777/_0_  ;
	output \g59778/_0_  ;
	output \g59779/_0_  ;
	output \g59780/_0_  ;
	output \g59781/_0_  ;
	output \g59789/_3_  ;
	output \g59799/_3_  ;
	output \g60311/_0_  ;
	output \g60326/_0_  ;
	output \g60333/_0_  ;
	output \g60336/_3_  ;
	output \g60341/_0_  ;
	output \g60343/_0_  ;
	output \g60344/_0_  ;
	output \g60345/_0_  ;
	output \g60354/_0_  ;
	output \g60355/_0_  ;
	output \g60356/_0_  ;
	output \g60357/_0_  ;
	output \g60358/_0_  ;
	output \g60359/_0_  ;
	output \g60360/_0_  ;
	output \g60361/_0_  ;
	output \g60362/_0_  ;
	output \g60363/_0_  ;
	output \g60364/_0_  ;
	output \g60398/_2_  ;
	output \g60399/_0_  ;
	output \g60400/_0_  ;
	output \g60401/_0_  ;
	output \g60402/_0_  ;
	output \g60403/_0_  ;
	output \g60406/_0_  ;
	output \g60410/_0_  ;
	output \g60411/_0_  ;
	output \g60417/_3_  ;
	output \g60419/_3_  ;
	output \g60421/_3_  ;
	output \g60423/_3_  ;
	output \g60425/_3_  ;
	output \g60427/_3_  ;
	output \g60429/_3_  ;
	output \g60431/_3_  ;
	output \g60433/_3_  ;
	output \g60435/_3_  ;
	output \g60437/_3_  ;
	output \g60439/_3_  ;
	output \g60441/_3_  ;
	output \g60443/_3_  ;
	output \g60445/_3_  ;
	output \g60447/_3_  ;
	output \g60449/_3_  ;
	output \g60451/_3_  ;
	output \g60453/_3_  ;
	output \g60455/_3_  ;
	output \g60457/_3_  ;
	output \g60459/_3_  ;
	output \g60461/_3_  ;
	output \g60463/_3_  ;
	output \g60465/_3_  ;
	output \g60467/_3_  ;
	output \g60469/_3_  ;
	output \g60471/_3_  ;
	output \g60473/_3_  ;
	output \g60475/_3_  ;
	output \g60477/_3_  ;
	output \g60479/_3_  ;
	output \g60481/_3_  ;
	output \g60483/_3_  ;
	output \g60485/_3_  ;
	output \g60487/_3_  ;
	output \g60489/_3_  ;
	output \g60491/_3_  ;
	output \g60493/_3_  ;
	output \g60495/_3_  ;
	output \g60497/_3_  ;
	output \g60499/_3_  ;
	output \g60501/_3_  ;
	output \g60503/_3_  ;
	output \g60505/_3_  ;
	output \g60507/_3_  ;
	output \g60509/_3_  ;
	output \g60511/_3_  ;
	output \g60513/_3_  ;
	output \g60515/_3_  ;
	output \g60517/_3_  ;
	output \g60519/_3_  ;
	output \g60521/_3_  ;
	output \g60523/_3_  ;
	output \g60525/_3_  ;
	output \g60527/_3_  ;
	output \g60529/_3_  ;
	output \g60531/_3_  ;
	output \g60533/_3_  ;
	output \g60535/_3_  ;
	output \g60537/_3_  ;
	output \g60539/_3_  ;
	output \g60541/_3_  ;
	output \g60544/_3_  ;
	output \g60546/_3_  ;
	output \g60548/_3_  ;
	output \g60550/_3_  ;
	output \g60552/_3_  ;
	output \g60554/_3_  ;
	output \g60556/_3_  ;
	output \g60559/_3_  ;
	output \g60561/_3_  ;
	output \g60563/_3_  ;
	output \g60565/_3_  ;
	output \g60567/_3_  ;
	output \g60569/_3_  ;
	output \g60571/_3_  ;
	output \g60573/_3_  ;
	output \g60575/_3_  ;
	output \g60577/_3_  ;
	output \g60579/_3_  ;
	output \g60581/_3_  ;
	output \g60583/_3_  ;
	output \g60585/_3_  ;
	output \g60588/_3_  ;
	output \g60590/_3_  ;
	output \g60593/_3_  ;
	output \g60596/_3_  ;
	output \g60598/_3_  ;
	output \g60600/_3_  ;
	output \g60602/_3_  ;
	output \g60603/_3_  ;
	output \g60671/_3_  ;
	output \g60672/_3_  ;
	output \g60674/_3_  ;
	output \g60680/_0_  ;
	output \g60682/_3_  ;
	output \g60690/_3_  ;
	output \g60692/_3_  ;
	output \g61594/_0_  ;
	output \g61614/_0_  ;
	output \g61618/_00_  ;
	output \g61649/_0_  ;
	output \g61651/_0_  ;
	output \g61656/_0_  ;
	output \g61657/_0_  ;
	output \g61659/_0_  ;
	output \g61662/_0_  ;
	output \g61663/_0_  ;
	output \g61664/_0_  ;
	output \g61665/_0_  ;
	output \g61667/_2_  ;
	output \g61669/_3__syn_2  ;
	output \g61678/_0_  ;
	output \g61679/_0_  ;
	output \g61680/_0_  ;
	output \g61681/_0_  ;
	output \g61684/_0_  ;
	output \g61685/_0_  ;
	output \g61686/_0_  ;
	output \g61690/_0_  ;
	output \g61692/_0_  ;
	output \g61694/_0_  ;
	output \g61695/_0_  ;
	output \g61696/_0_  ;
	output \g61699/u3_syn_4  ;
	output \g61732/u3_syn_4  ;
	output \g61765/u3_syn_4  ;
	output \g61798/u3_syn_4  ;
	output \g61848/_0_  ;
	output \g61848/_3_  ;
	output \g61853/_0_  ;
	output \g61854/_1__syn_2  ;
	output \g61858/u3_syn_4  ;
	output \g61880/u3_syn_4  ;
	output \g61887/u3_syn_4  ;
	output \g61920/u3_syn_4  ;
	output \g61990/u3_syn_4  ;
	output \g62254/_0__syn_2  ;
	output \g62260/_0_  ;
	output \g62262/_1__syn_2  ;
	output \g62290/_0_  ;
	output \g62317/_0_  ;
	output \g62319/_0_  ;
	output \g62324/_0_  ;
	output \g62329/_0_  ;
	output \g62331/_0_  ;
	output \g62331/_1_  ;
	output \g62333/u3_syn_4  ;
	output \g62335/u3_syn_4  ;
	output \g62336/u3_syn_4  ;
	output \g62428/u3_syn_4  ;
	output \g62454/u3_syn_4  ;
	output \g62487/u3_syn_4  ;
	output \g62520/u3_syn_4  ;
	output \g62552/u3_syn_4  ;
	output \g62584/u3_syn_4  ;
	output \g62619/u3_syn_4  ;
	output \g62651/u3_syn_4  ;
	output \g62692/_0_  ;
	output \g62873/_0_  ;
	output \g62882/_0_  ;
	output \g62883/u3_syn_4  ;
	output \g62886/u3_syn_4  ;
	output \g62908/u3_syn_4  ;
	output \g62952/u3_syn_4  ;
	output \g62974/u3_syn_4  ;
	output \g63207/_0_  ;
	output \g63214/_3_  ;
	output \g63227/_0_  ;
	output \g63250/_1__syn_2  ;
	output \g63315/_0__syn_2  ;
	output \g63320/_0_  ;
	output \g63322/_0_  ;
	output \g63324/_2_  ;
	output \g63338/_0__syn_2  ;
	output \g63340/_0_  ;
	output \g63376/_0_  ;
	output \g63395/_2_  ;
	output \g63398/_0_  ;
	output \g63419/_0_  ;
	output \g63524/_3_  ;
	output \g63540/_0_  ;
	output \g63541/_0_  ;
	output \g63682/_0_  ;
	output \g63890/_1_  ;
	output \g63892/_0_  ;
	output \g63894/_0_  ;
	output \g63897/_1_  ;
	output \g63908/_0_  ;
	output \g63913/_0_  ;
	output \g63914/_0_  ;
	output \g63927/_1__syn_2  ;
	output \g63934/_0_  ;
	output \g63942/_0_  ;
	output \g63952/_0_  ;
	output \g63965/_0_  ;
	output \g63969/_0_  ;
	output \g63985/_0_  ;
	output \g63986/_0_  ;
	output \g63987/_0_  ;
	output \g63988/_0_  ;
	output \g63990/_0_  ;
	output \g63991/_0_  ;
	output \g63992/_0_  ;
	output \g63993/_0_  ;
	output \g64016/_0_  ;
	output \g64017/_0_  ;
	output \g64018/_0_  ;
	output \g64019/_0_  ;
	output \g64020/_0_  ;
	output \g64021/_0_  ;
	output \g64023/_0_  ;
	output \g64024/_0_  ;
	output \g64101/_0_  ;
	output \g64104/_0_  ;
	output \g64121/_0_  ;
	output \g64174/_0_  ;
	output \g64249/_0_  ;
	output \g64299/_0_  ;
	output \g64338/_0_  ;
	output \g64364/_0_  ;
	output \g64459/_0_  ;
	output \g64461/_0_  ;
	output \g64466/_0_  ;
	output \g64577/_0_  ;
	output \g64583/_0_  ;
	output \g64589/_1_  ;
	output \g64595/_0_  ;
	output \g64598/_0_  ;
	output \g64649/_0_  ;
	output \g64678/_0_  ;
	output \g64688/_3_  ;
	output \g64689/_0_  ;
	output \g64694/_0_  ;
	output \g64695/_0_  ;
	output \g64700/_0_  ;
	output \g64714/_0_  ;
	output \g64744/_2_  ;
	output \g65255/_0_  ;
	output \g65258/_0_  ;
	output \g65269/_3_  ;
	output \g65489/_0_  ;
	output \g65513/_0_  ;
	output \g65530/_0_  ;
	output \g65561/_0_  ;
	output \g65563/_0_  ;
	output \g65564/_0_  ;
	output \g65573/_0_  ;
	output \g65578/_2_  ;
	output \g65597/_0_  ;
	output \g65605/_0_  ;
	output \g65606/_0_  ;
	output \g65609/_0_  ;
	output \g65611/_0_  ;
	output \g65612/_0_  ;
	output \g65613/_0_  ;
	output \g65615/_0_  ;
	output \g65618/_0_  ;
	output \g65631/_0_  ;
	output \g65634/_0_  ;
	output \g65635/_0_  ;
	output \g65639/_0_  ;
	output \g65644/_0_  ;
	output \g65648/_0_  ;
	output \g65650/_0_  ;
	output \g65662/_3_  ;
	output \g65665/_3_  ;
	output \g65729/_0_  ;
	output \g65801/_0_  ;
	output \g66072/_0_  ;
	output \g66074/_0_  ;
	output \g66075/_0_  ;
	output \g66076/_0_  ;
	output \g66077/_0_  ;
	output \g66078/_0_  ;
	output \g66079/_0_  ;
	output \g66080/_0_  ;
	output \g66081/_0_  ;
	output \g66082/_0_  ;
	output \g66085/_0_  ;
	output \g66086/_0_  ;
	output \g66087/_0_  ;
	output \g66089/_0_  ;
	output \g66090/_0_  ;
	output \g66093/_0_  ;
	output \g66094/_0_  ;
	output \g66095/_0_  ;
	output \g66098/_0_  ;
	output \g66100/_0_  ;
	output \g66106/_1_  ;
	output \g66107/_0_  ;
	output \g66108/_0_  ;
	output \g66110/_0_  ;
	output \g66114/_0_  ;
	output \g66124/_0_  ;
	output \g66125/_0_  ;
	output \g66127/_0_  ;
	output \g66128/_0_  ;
	output \g66129/_0_  ;
	output \g66130/_0_  ;
	output \g66133/_0_  ;
	output \g66134/_0_  ;
	output \g66136/_0_  ;
	output \g66141/_1_  ;
	output \g66153/_0_  ;
	output \g66182/_0_  ;
	output \g66187/_0_  ;
	output \g66240/_0_  ;
	output \g66268/_0_  ;
	output \g66354/_0_  ;
	output \g66397/_3_  ;
	output \g66398/_3_  ;
	output \g66399/_3_  ;
	output \g66400/_3_  ;
	output \g66401/_3_  ;
	output \g66402/_3_  ;
	output \g66403/_3_  ;
	output \g66404/_3_  ;
	output \g66405/_3_  ;
	output \g66406/_3_  ;
	output \g66407/_3_  ;
	output \g66408/_3_  ;
	output \g66409/_3_  ;
	output \g66410/_3_  ;
	output \g66411/_3_  ;
	output \g66412/_3_  ;
	output \g66413/_3_  ;
	output \g66414/_3_  ;
	output \g66415/_3_  ;
	output \g66416/_3_  ;
	output \g66417/_3_  ;
	output \g66418/_3_  ;
	output \g66419/_3_  ;
	output \g66420/_3_  ;
	output \g66421/_3_  ;
	output \g66422/_3_  ;
	output \g66423/_3_  ;
	output \g66424/_3_  ;
	output \g66425/_3_  ;
	output \g66426/_3_  ;
	output \g66427/_3_  ;
	output \g66428/_3_  ;
	output \g66429/_3_  ;
	output \g66430/_3_  ;
	output \g66464/_0_  ;
	output \g66465/_0_  ;
	output \g66477/_3_  ;
	output \g66643/_0_  ;
	output \g66733/_2_  ;
	output \g66735/_1_  ;
	output \g66801/_0_  ;
	output \g66866/_0_  ;
	output \g66875/_0_  ;
	output \g66885/_1_  ;
	output \g66890/_0_  ;
	output \g66939/_0_  ;
	output \g66950/_0_  ;
	output \g67035/_0_  ;
	output \g67038/_0_  ;
	output \g67044/_3_  ;
	output \g67045/_3_  ;
	output \g67046/_3_  ;
	output \g67070/_3_  ;
	output \g67082/_3_  ;
	output \g67090/_3_  ;
	output \g67106/_0_  ;
	output \g67107/_0_  ;
	output \g67108/_0_  ;
	output \g67109/_0_  ;
	output \g67117/_0_  ;
	output \g67131/_0_  ;
	output \g67142/_0_  ;
	output \g67421/_0_  ;
	output \g67456/_0_  ;
	output \g67464/_0_  ;
	output \g67617/_1_  ;
	output \g67772/_0_  ;
	output \g68523/_0_  ;
	output \g73970/_0_  ;
	output \g73976/_0_  ;
	output \g74120/_1_  ;
	output \g74148/_2_  ;
	output \g74245/_0_  ;
	output \g74426/_0_  ;
	output \g74434/_3_  ;
	output \g74589/_0_  ;
	output \g74626/_1__syn_2  ;
	output \g74790/_0_  ;
	output \g74801/_0_  ;
	output \g74838/_0_  ;
	output \g74850/_0_  ;
	output \g74855/_0_  ;
	output \g74862/_0_  ;
	output \g74871/_0_  ;
	output \g74878/_0_  ;
	output \g74885/_0_  ;
	output \g74922/_0_  ;
	output \g75066/_1__syn_2  ;
	output \g75100/_1_  ;
	output \g75201/_1_  ;
	output \g75205/_1_  ;
	output \g75420/_1_  ;
	output pci_rst_oe_o_pad ;
	output wb_int_o_pad ;
	output wb_rst_o_pad ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3779_ ;
	wire _w5539_ ;
	wire _w452_ ;
	wire _w5166_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3024_ ;
	wire _w3021_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3048_ ;
	wire _w3022_ ;
	wire _w3119_ ;
	wire _w3033_ ;
	wire _w3020_ ;
	wire _w3023_ ;
	wire _w3036_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3078_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3276_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w4734_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w4744_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w20_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w30_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\configuration_init_complete_reg/NET0131 ,
		_w20_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\configuration_interrupt_out_reg/NET0131 ,
		_w30_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\output_backup_frame_en_out_reg/NET0131 ,
		_w452_
	);
	LUT4 #(
		.INIT('h8421)
	) name3 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]/NET0131 ,
		_w3015_
	);
	LUT4 #(
		.INIT('h8421)
	) name4 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]/NET0131 ,
		_w3016_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\input_register_pci_devsel_reg_out_reg/NET0131 ,
		\input_register_pci_trdy_reg_out_reg/NET0131 ,
		_w3018_
	);
	LUT4 #(
		.INIT('h0110)
	) name7 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w3019_
	);
	LUT4 #(
		.INIT('h5111)
	) name8 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('ha2)
	) name9 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131 ,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3022_
	);
	LUT3 #(
		.INIT('h04)
	) name11 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3023_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name12 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131 ,
		_w3024_
	);
	LUT2 #(
		.INIT('h9)
	) name13 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]/NET0131 ,
		_w3025_
	);
	LUT4 #(
		.INIT('haf23)
	) name14 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_outGreyCount_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]/NET0131 ,
		_w3026_
	);
	LUT3 #(
		.INIT('h80)
	) name15 (
		_w3024_,
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT3 #(
		.INIT('h01)
	) name16 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3028_
	);
	LUT3 #(
		.INIT('h70)
	) name17 (
		_w3015_,
		_w3016_,
		_w3028_,
		_w3029_
	);
	LUT3 #(
		.INIT('h45)
	) name18 (
		_w3023_,
		_w3027_,
		_w3029_,
		_w3030_
	);
	LUT3 #(
		.INIT('h45)
	) name19 (
		_w3017_,
		_w3021_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h8a88)
	) name20 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w3032_
	);
	LUT4 #(
		.INIT('h2022)
	) name21 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w3033_
	);
	LUT2 #(
		.INIT('he)
	) name22 (
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\configuration_command_bit6_reg/NET0131 ,
		\configuration_init_complete_reg/NET0131 ,
		_w3035_
	);
	LUT4 #(
		.INIT('h070f)
	) name24 (
		\configuration_command_bit6_reg/NET0131 ,
		\configuration_init_complete_reg/NET0131 ,
		\parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131 ,
		\parity_checker_perr_sampled_reg/NET0131 ,
		_w3036_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\parity_checker_master_perr_report_reg/NET0131 ,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3039_
	);
	LUT3 #(
		.INIT('h01)
	) name28 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3040_
	);
	LUT3 #(
		.INIT('h02)
	) name29 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3041_
	);
	LUT4 #(
		.INIT('h0002)
	) name30 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3042_
	);
	LUT3 #(
		.INIT('h40)
	) name31 (
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w3045_
	);
	LUT4 #(
		.INIT('h0400)
	) name34 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131 ,
		_w3046_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w3044_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name36 (
		\configuration_status_bit8_reg/NET0131 ,
		_w3038_,
		_w3043_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('he)
	) name37 (
		_w3037_,
		_w3048_,
		_w3049_
	);
	LUT3 #(
		.INIT('h08)
	) name38 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		_w3051_
	);
	LUT3 #(
		.INIT('h10)
	) name40 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3052_
	);
	LUT4 #(
		.INIT('h8000)
	) name41 (
		\pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131 ,
		_w3053_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131 ,
		_w3054_
	);
	LUT4 #(
		.INIT('h4000)
	) name43 (
		\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131 ,
		_w3055_
	);
	LUT3 #(
		.INIT('h80)
	) name44 (
		_w3052_,
		_w3053_,
		_w3055_,
		_w3056_
	);
	LUT3 #(
		.INIT('h02)
	) name45 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\pci_target_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[3]/NET0131 ,
		_w3058_
	);
	LUT4 #(
		.INIT('h0040)
	) name47 (
		\pci_target_unit_del_sync_bc_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_burst_out_reg/NET0131 ,
		\pci_target_unit_wishbone_master_read_bound_reg/NET0131 ,
		_w3059_
	);
	LUT3 #(
		.INIT('h04)
	) name48 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3060_
	);
	LUT4 #(
		.INIT('hfecf)
	) name49 (
		\pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131 ,
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3061_
	);
	LUT4 #(
		.INIT('h7500)
	) name50 (
		_w3057_,
		_w3058_,
		_w3059_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h8c)
	) name51 (
		_w3056_,
		_w3050_,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h6)
	) name52 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		_w3064_
	);
	LUT4 #(
		.INIT('h8421)
	) name53 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		_w3065_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w3064_,
		_w3065_,
		_w3066_
	);
	LUT3 #(
		.INIT('h45)
	) name55 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		_w3064_,
		_w3065_,
		_w3067_
	);
	LUT3 #(
		.INIT('h02)
	) name56 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w3068_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w3060_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w3068_,
		_w3057_,
		_w3070_
	);
	LUT4 #(
		.INIT('h0200)
	) name59 (
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w3071_
	);
	LUT4 #(
		.INIT('h00ab)
	) name60 (
		_w3067_,
		_w3070_,
		_w3069_,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w3063_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('hb)
	) name62 (
		_w3063_,
		_w3072_,
		_w3074_
	);
	LUT3 #(
		.INIT('hf9)
	) name63 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3075_
	);
	LUT3 #(
		.INIT('he9)
	) name64 (
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3076_
	);
	LUT3 #(
		.INIT('h01)
	) name65 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w3077_
	);
	LUT4 #(
		.INIT('h0001)
	) name66 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		\pci_target_unit_wishbone_master_retried_reg/NET0131 ,
		_w3078_
	);
	LUT4 #(
		.INIT('h0082)
	) name67 (
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_wishbone_master_w_attempt_reg/NET0131 ,
		_w3079_
	);
	LUT3 #(
		.INIT('h20)
	) name68 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		\pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131 ,
		\pci_target_unit_wishbone_master_w_attempt_reg/NET0131 ,
		_w3080_
	);
	LUT4 #(
		.INIT('haa80)
	) name69 (
		_w3078_,
		_w3065_,
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]/NET0131 ,
		_w3082_
	);
	LUT3 #(
		.INIT('hb0)
	) name71 (
		_w3064_,
		_w3065_,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w3081_,
		_w3083_,
		_w3084_
	);
	LUT3 #(
		.INIT('h80)
	) name73 (
		_w3078_,
		_w3065_,
		_w3079_,
		_w3085_
	);
	LUT4 #(
		.INIT('h8000)
	) name74 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 ,
		_w3078_,
		_w3065_,
		_w3079_,
		_w3086_
	);
	LUT3 #(
		.INIT('h13)
	) name75 (
		\pci_target_unit_del_sync_burst_out_reg/NET0131 ,
		\pci_target_unit_wishbone_master_first_data_is_burst_reg_reg/NET0131 ,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h7500)
	) name76 (
		\pci_target_unit_wishbone_master_burst_chopped_reg/NET0131 ,
		_w3084_,
		_w3087_,
		_w3057_,
		_w3088_
	);
	LUT4 #(
		.INIT('h0c0e)
	) name77 (
		_w3067_,
		_w3075_,
		_w3076_,
		_w3088_,
		_w3089_
	);
	LUT3 #(
		.INIT('h80)
	) name78 (
		_w3077_,
		_w3065_,
		_w3079_,
		_w3090_
	);
	LUT4 #(
		.INIT('h0100)
	) name79 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		\pci_target_unit_wishbone_master_w_attempt_reg/NET0131 ,
		_w3091_
	);
	LUT3 #(
		.INIT('h70)
	) name80 (
		_w3065_,
		_w3079_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('h0200)
	) name81 (
		\pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131 ,
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3093_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w3050_,
		_w3093_,
		_w3094_
	);
	LUT3 #(
		.INIT('h01)
	) name83 (
		_w3092_,
		_w3094_,
		_w3090_,
		_w3095_
	);
	LUT3 #(
		.INIT('h2f)
	) name84 (
		_w3068_,
		_w3089_,
		_w3095_,
		_w3096_
	);
	LUT4 #(
		.INIT('h08cc)
	) name85 (
		_w3068_,
		_w3073_,
		_w3089_,
		_w3095_,
		_w3097_
	);
	LUT4 #(
		.INIT('h4500)
	) name86 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		_w3064_,
		_w3065_,
		_w3060_,
		_w3098_
	);
	LUT3 #(
		.INIT('hc8)
	) name87 (
		_w3056_,
		_w3068_,
		_w3098_,
		_w3099_
	);
	LUT4 #(
		.INIT('h00df)
	) name88 (
		_w3057_,
		_w3058_,
		_w3059_,
		_w3076_,
		_w3100_
	);
	LUT3 #(
		.INIT('h04)
	) name89 (
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w3101_
	);
	LUT4 #(
		.INIT('h4500)
	) name90 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		_w3064_,
		_w3065_,
		_w3101_,
		_w3102_
	);
	LUT4 #(
		.INIT('h0501)
	) name91 (
		_w3102_,
		_w3050_,
		_w3090_,
		_w3100_,
		_w3103_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w3099_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('hb)
	) name93 (
		_w3099_,
		_w3103_,
		_w3105_
	);
	LUT4 #(
		.INIT('haf23)
	) name94 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131 ,
		_w3106_
	);
	LUT2 #(
		.INIT('h9)
	) name95 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]/NET0131 ,
		_w3107_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name96 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]/NET0131 ,
		_w3108_
	);
	LUT4 #(
		.INIT('h1555)
	) name97 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 ,
		_w3106_,
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('h4000)
	) name98 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		_w3052_,
		_w3053_,
		_w3055_,
		_w3110_
	);
	LUT4 #(
		.INIT('h888a)
	) name99 (
		\pci_target_unit_wishbone_master_burst_chopped_reg/NET0131 ,
		_w3066_,
		_w3060_,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('hb0)
	) name100 (
		_w3084_,
		_w3087_,
		_w3111_,
		_w3112_
	);
	LUT4 #(
		.INIT('h4500)
	) name101 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]/NET0131 ,
		_w3064_,
		_w3065_,
		_w3057_,
		_w3113_
	);
	LUT4 #(
		.INIT('h00ab)
	) name102 (
		_w3066_,
		_w3060_,
		_w3110_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		_w3068_,
		_w3114_,
		_w3115_
	);
	LUT4 #(
		.INIT('h1500)
	) name104 (
		\pci_target_unit_wishbone_master_retried_reg/NET0131 ,
		_w3065_,
		_w3079_,
		_w3091_,
		_w3116_
	);
	LUT3 #(
		.INIT('h01)
	) name105 (
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		_w3102_,
		_w3116_,
		_w3117_
	);
	LUT4 #(
		.INIT('h1055)
	) name106 (
		_w3109_,
		_w3112_,
		_w3115_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\pci_target_unit_wishbone_master_burst_chopped_delayed_reg/NET0131 ,
		\pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131 ,
		_w3119_
	);
	LUT4 #(
		.INIT('h0151)
	) name108 (
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		\pci_target_unit_wishbone_master_retried_reg/NET0131 ,
		\pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131 ,
		wbm_ack_i_pad,
		_w3120_
	);
	LUT3 #(
		.INIT('h45)
	) name109 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT3 #(
		.INIT('hb0)
	) name110 (
		_w3084_,
		_w3087_,
		_w3121_,
		_w3122_
	);
	LUT3 #(
		.INIT('h10)
	) name111 (
		\wbm_cti_o[0]_pad ,
		_w3119_,
		_w3120_,
		_w3123_
	);
	LUT3 #(
		.INIT('h0b)
	) name112 (
		_w3118_,
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\wbm_cti_o[0]_pad ,
		_w3120_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131 ,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w3120_,
		_w3126_,
		_w3127_
	);
	LUT4 #(
		.INIT('h040f)
	) name116 (
		_w3084_,
		_w3087_,
		_w3125_,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('ha280)
	) name117 (
		_w3097_,
		_w3104_,
		_w3124_,
		_w3128_,
		_w3129_
	);
	LUT3 #(
		.INIT('h01)
	) name118 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131 ,
		_w3130_
	);
	LUT4 #(
		.INIT('h0002)
	) name119 (
		\configuration_wb_init_complete_out_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131 ,
		_w3131_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		wbs_cyc_i_pad,
		wbs_stb_i_pad,
		_w3132_
	);
	LUT3 #(
		.INIT('h40)
	) name121 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		wbs_cyc_i_pad,
		wbs_stb_i_pad,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w3131_,
		_w3133_,
		_w3134_
	);
	LUT3 #(
		.INIT('h80)
	) name123 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		_w3135_
	);
	LUT4 #(
		.INIT('h7f00)
	) name124 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3136_
	);
	LUT3 #(
		.INIT('h80)
	) name125 (
		\wbs_cti_i[0]_pad ,
		\wbs_cti_i[1]_pad ,
		\wbs_cti_i[2]_pad ,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		wbs_stb_i_pad,
		_w3138_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		_w3139_
	);
	LUT4 #(
		.INIT('hba00)
	) name128 (
		_w3130_,
		_w3137_,
		_w3138_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\wishbone_slave_unit_wishbone_slave_img_hit_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_img_hit_reg[1]/NET0131 ,
		_w3141_
	);
	LUT3 #(
		.INIT('h08)
	) name130 (
		\wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3142_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w3141_,
		_w3142_,
		_w3143_
	);
	LUT3 #(
		.INIT('he0)
	) name132 (
		_w3140_,
		_w3135_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		_w3145_
	);
	LUT3 #(
		.INIT('h80)
	) name134 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		_w3146_
	);
	LUT4 #(
		.INIT('h00e0)
	) name135 (
		_w3140_,
		_w3135_,
		_w3143_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_del_completion_allow_reg/NET0131 ,
		_w3148_
	);
	LUT3 #(
		.INIT('h31)
	) name137 (
		_w3140_,
		_w3135_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h50dc)
	) name138 (
		\wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3148_,
		_w3150_
	);
	LUT3 #(
		.INIT('h02)
	) name139 (
		_w3147_,
		_w3150_,
		_w3136_,
		_w3151_
	);
	LUT4 #(
		.INIT('h8421)
	) name140 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]/NET0131 ,
		_w3152_
	);
	LUT4 #(
		.INIT('h8421)
	) name141 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]/NET0131 ,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w3152_,
		_w3153_,
		_w3154_
	);
	LUT4 #(
		.INIT('h9009)
	) name143 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]/NET0131 ,
		_w3155_
	);
	LUT4 #(
		.INIT('h8421)
	) name144 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]/NET0131 ,
		_w3156_
	);
	LUT4 #(
		.INIT('h0777)
	) name145 (
		_w3152_,
		_w3153_,
		_w3155_,
		_w3156_,
		_w3157_
	);
	LUT3 #(
		.INIT('h10)
	) name146 (
		\wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3158_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w3145_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('hd0)
	) name148 (
		_w3135_,
		_w3157_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h80)
	) name149 (
		_w3135_,
		_w3157_,
		_w3159_,
		_w3161_
	);
	LUT4 #(
		.INIT('h7000)
	) name150 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3162_
	);
	LUT4 #(
		.INIT('h8421)
	) name151 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131 ,
		_w3163_
	);
	LUT4 #(
		.INIT('h8421)
	) name152 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		_w3164_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w3163_,
		_w3164_,
		_w3165_
	);
	LUT3 #(
		.INIT('h20)
	) name154 (
		\wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3166_
	);
	LUT4 #(
		.INIT('h2a00)
	) name155 (
		_w3145_,
		_w3163_,
		_w3164_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w3140_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h00bf)
	) name157 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3140_,
		_w3167_,
		_w3162_,
		_w3169_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w3161_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w3137_,
		_w3171_,
		_w3172_
	);
	LUT4 #(
		.INIT('h00ba)
	) name161 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		_w3151_,
		_w3170_,
		_w3172_,
		_w3173_
	);
	LUT4 #(
		.INIT('h0a02)
	) name162 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3140_,
		_w3135_,
		_w3148_,
		_w3174_
	);
	LUT4 #(
		.INIT('h8000)
	) name163 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3175_
	);
	LUT4 #(
		.INIT('h007f)
	) name164 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3140_,
		_w3167_,
		_w3175_,
		_w3176_
	);
	LUT4 #(
		.INIT('h5700)
	) name165 (
		_w3144_,
		_w3146_,
		_w3174_,
		_w3176_,
		_w3177_
	);
	LUT3 #(
		.INIT('h20)
	) name166 (
		_w3135_,
		_w3157_,
		_w3159_,
		_w3178_
	);
	LUT4 #(
		.INIT('h002a)
	) name167 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg/NET0131 ,
		_w3147_,
		_w3150_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w3177_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('hfdcc)
	) name169 (
		_w3132_,
		_w3134_,
		_w3173_,
		_w3180_,
		_w3181_
	);
	LUT4 #(
		.INIT('h1055)
	) name170 (
		_w3081_,
		_w3112_,
		_w3115_,
		_w3117_,
		_w3182_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h5574)
	) name172 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]/P0001 ,
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		\wbm_sel_o[0]_pad ,
		_w3182_,
		_w3184_
	);
	LUT3 #(
		.INIT('h80)
	) name173 (
		_w3097_,
		_w3104_,
		_w3184_,
		_w3185_
	);
	LUT3 #(
		.INIT('h20)
	) name174 (
		\pci_target_unit_del_sync_be_out_reg[0]/NET0131 ,
		_w3084_,
		_w3087_,
		_w3186_
	);
	LUT4 #(
		.INIT('hddd1)
	) name175 (
		\wbm_sel_o[0]_pad ,
		_w3097_,
		_w3104_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('hb)
	) name176 (
		_w3185_,
		_w3187_,
		_w3188_
	);
	LUT4 #(
		.INIT('h5574)
	) name177 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]/P0001 ,
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		\wbm_sel_o[2]_pad ,
		_w3182_,
		_w3189_
	);
	LUT3 #(
		.INIT('h80)
	) name178 (
		_w3097_,
		_w3104_,
		_w3189_,
		_w3190_
	);
	LUT3 #(
		.INIT('h20)
	) name179 (
		\pci_target_unit_del_sync_be_out_reg[2]/NET0131 ,
		_w3084_,
		_w3087_,
		_w3191_
	);
	LUT4 #(
		.INIT('hddd1)
	) name180 (
		\wbm_sel_o[2]_pad ,
		_w3097_,
		_w3104_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('hb)
	) name181 (
		_w3190_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('h5574)
	) name182 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]/P0001 ,
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		\wbm_sel_o[1]_pad ,
		_w3182_,
		_w3194_
	);
	LUT3 #(
		.INIT('h80)
	) name183 (
		_w3097_,
		_w3104_,
		_w3194_,
		_w3195_
	);
	LUT3 #(
		.INIT('h20)
	) name184 (
		\pci_target_unit_del_sync_be_out_reg[1]/NET0131 ,
		_w3084_,
		_w3087_,
		_w3196_
	);
	LUT4 #(
		.INIT('hddd1)
	) name185 (
		\wbm_sel_o[1]_pad ,
		_w3097_,
		_w3104_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('hb)
	) name186 (
		_w3195_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('h5574)
	) name187 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]/P0001 ,
		\pci_target_unit_wishbone_master_addr_into_cnt_reg_reg/NET0131 ,
		\wbm_sel_o[3]_pad ,
		_w3182_,
		_w3199_
	);
	LUT3 #(
		.INIT('h80)
	) name188 (
		_w3097_,
		_w3104_,
		_w3199_,
		_w3200_
	);
	LUT3 #(
		.INIT('h20)
	) name189 (
		\pci_target_unit_del_sync_be_out_reg[3]/NET0131 ,
		_w3084_,
		_w3087_,
		_w3201_
	);
	LUT4 #(
		.INIT('hddd1)
	) name190 (
		\wbm_sel_o[3]_pad ,
		_w3097_,
		_w3104_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('hb)
	) name191 (
		_w3200_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h02)
	) name192 (
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3204_
	);
	LUT3 #(
		.INIT('h10)
	) name193 (
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3205_
	);
	LUT3 #(
		.INIT('h27)
	) name194 (
		\output_backup_frame_en_out_reg/NET0131 ,
		\output_backup_frame_out_reg/NET0131 ,
		pci_frame_i_pad,
		_w3206_
	);
	LUT3 #(
		.INIT('hd8)
	) name195 (
		\output_backup_frame_en_out_reg/NET0131 ,
		\output_backup_frame_out_reg/NET0131 ,
		pci_frame_i_pad,
		_w3207_
	);
	LUT3 #(
		.INIT('h27)
	) name196 (
		\output_backup_irdy_en_out_reg/NET0131 ,
		\output_backup_irdy_out_reg/NET0131 ,
		pci_irdy_i_pad,
		_w3208_
	);
	LUT3 #(
		.INIT('hd8)
	) name197 (
		\output_backup_irdy_en_out_reg/NET0131 ,
		\output_backup_irdy_out_reg/NET0131 ,
		pci_irdy_i_pad,
		_w3209_
	);
	LUT3 #(
		.INIT('h80)
	) name198 (
		_w3205_,
		_w3206_,
		_w3208_,
		_w3210_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w3044_,
		_w3205_,
		_w3211_
	);
	LUT3 #(
		.INIT('h04)
	) name200 (
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3212_
	);
	LUT4 #(
		.INIT('h5277)
	) name201 (
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		_w3213_
	);
	LUT3 #(
		.INIT('h04)
	) name202 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		_w3214_
	);
	LUT4 #(
		.INIT('haa08)
	) name203 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT3 #(
		.INIT('h10)
	) name204 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w3216_
	);
	LUT4 #(
		.INIT('hef00)
	) name205 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131 ,
		_w3217_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		_w3219_
	);
	LUT3 #(
		.INIT('h01)
	) name208 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		_w3220_
	);
	LUT3 #(
		.INIT('h20)
	) name209 (
		_w3218_,
		_w3220_,
		_w3217_,
		_w3221_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		_w3215_,
		_w3221_,
		_w3222_
	);
	LUT3 #(
		.INIT('h8a)
	) name211 (
		_w3212_,
		_w3215_,
		_w3221_,
		_w3223_
	);
	LUT4 #(
		.INIT('h0200)
	) name212 (
		\pci_target_unit_pci_target_sm_backoff_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\pci_target_unit_pci_target_sm_state_backoff_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_state_transfere_reg_reg/NET0131 ,
		_w3225_
	);
	LUT3 #(
		.INIT('h8a)
	) name214 (
		_w3045_,
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT4 #(
		.INIT('h0075)
	) name215 (
		_w3212_,
		_w3215_,
		_w3221_,
		_w3226_,
		_w3227_
	);
	LUT4 #(
		.INIT('h0200)
	) name216 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131 ,
		_w3228_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w3227_,
		_w3228_,
		_w3229_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name218 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131 ,
		_w3230_
	);
	LUT2 #(
		.INIT('h9)
	) name219 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]/NET0131 ,
		_w3231_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name220 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]/NET0131 ,
		_w3232_
	);
	LUT3 #(
		.INIT('h80)
	) name221 (
		_w3230_,
		_w3231_,
		_w3232_,
		_w3233_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name222 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131 ,
		_w3234_
	);
	LUT2 #(
		.INIT('h9)
	) name223 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]/NET0131 ,
		_w3235_
	);
	LUT4 #(
		.INIT('haf23)
	) name224 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]/NET0131 ,
		_w3236_
	);
	LUT3 #(
		.INIT('h80)
	) name225 (
		_w3234_,
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name226 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131 ,
		_w3238_
	);
	LUT2 #(
		.INIT('h9)
	) name227 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]/NET0131 ,
		_w3239_
	);
	LUT4 #(
		.INIT('haf23)
	) name228 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]/NET0131 ,
		_w3240_
	);
	LUT3 #(
		.INIT('h80)
	) name229 (
		_w3238_,
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w3237_,
		_w3241_,
		_w3242_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name231 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		_w3243_
	);
	LUT2 #(
		.INIT('h9)
	) name232 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]/NET0131 ,
		_w3244_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name233 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		_w3245_
	);
	LUT3 #(
		.INIT('h80)
	) name234 (
		_w3243_,
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT4 #(
		.INIT('h1110)
	) name235 (
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		_w3247_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		\pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w3247_,
		_w3248_,
		_w3249_
	);
	LUT4 #(
		.INIT('h0100)
	) name238 (
		_w3237_,
		_w3241_,
		_w3246_,
		_w3249_,
		_w3250_
	);
	LUT4 #(
		.INIT('hbf00)
	) name239 (
		_w3227_,
		_w3228_,
		_w3233_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name240 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		_w3252_
	);
	LUT2 #(
		.INIT('h9)
	) name241 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131 ,
		_w3253_
	);
	LUT4 #(
		.INIT('haf23)
	) name242 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		_w3254_
	);
	LUT3 #(
		.INIT('h80)
	) name243 (
		_w3252_,
		_w3253_,
		_w3254_,
		_w3255_
	);
	LUT3 #(
		.INIT('h13)
	) name244 (
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131 ,
		_w3256_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		_w3219_,
		_w3256_,
		_w3257_
	);
	LUT3 #(
		.INIT('h04)
	) name246 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3219_,
		_w3256_,
		_w3258_
	);
	LUT3 #(
		.INIT('h45)
	) name247 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		_w3255_,
		_w3258_,
		_w3259_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name248 (
		_w3045_,
		_w3252_,
		_w3253_,
		_w3254_,
		_w3260_
	);
	LUT4 #(
		.INIT('ha0c0)
	) name249 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3261_,
		_w3262_
	);
	LUT4 #(
		.INIT('h0045)
	) name251 (
		_w3211_,
		_w3251_,
		_w3259_,
		_w3262_,
		_w3263_
	);
	LUT4 #(
		.INIT('h2232)
	) name252 (
		\pci_target_unit_pci_target_sm_backoff_reg/NET0131 ,
		_w3204_,
		_w3210_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_progress_reg/NET0131 ,
		_w3266_
	);
	LUT4 #(
		.INIT('h5150)
	) name255 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3261_,
		_w3265_,
		_w3266_,
		_w3267_
	);
	LUT3 #(
		.INIT('h13)
	) name256 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_wr_progress_reg/NET0131 ,
		_w3268_
	);
	LUT4 #(
		.INIT('h8a88)
	) name257 (
		_w3212_,
		_w3222_,
		_w3267_,
		_w3268_,
		_w3269_
	);
	LUT4 #(
		.INIT('h5551)
	) name258 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3270_
	);
	LUT4 #(
		.INIT('h8000)
	) name259 (
		_w3205_,
		_w3206_,
		_w3208_,
		_w3270_,
		_w3271_
	);
	LUT3 #(
		.INIT('h40)
	) name260 (
		_w3215_,
		_w3221_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w3269_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('hb)
	) name262 (
		_w3264_,
		_w3273_,
		_w3274_
	);
	LUT4 #(
		.INIT('h2070)
	) name263 (
		\output_backup_perr_en_out_reg/NET0131 ,
		\output_backup_perr_out_reg/NET0131 ,
		\parity_checker_check_perr_reg/NET0131 ,
		pci_perr_i_pad,
		_w3275_
	);
	LUT3 #(
		.INIT('h37)
	) name264 (
		_w3068_,
		_w3057_,
		_w3050_,
		_w3276_
	);
	LUT4 #(
		.INIT('h8000)
	) name265 (
		\wbm_adr_o[4]_pad ,
		\wbm_adr_o[5]_pad ,
		\wbm_adr_o[6]_pad ,
		\wbm_adr_o[9]_pad ,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\wbm_adr_o[7]_pad ,
		\wbm_adr_o[8]_pad ,
		_w3278_
	);
	LUT4 #(
		.INIT('h8000)
	) name267 (
		\wbm_adr_o[2]_pad ,
		\wbm_adr_o[3]_pad ,
		\wbm_adr_o[7]_pad ,
		\wbm_adr_o[8]_pad ,
		_w3279_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w3277_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\wbm_adr_o[10]_pad ,
		\wbm_adr_o[11]_pad ,
		_w3281_
	);
	LUT4 #(
		.INIT('h2000)
	) name270 (
		\wbm_adr_o[12]_pad ,
		_w3276_,
		_w3280_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h8000)
	) name271 (
		\wbm_adr_o[13]_pad ,
		\wbm_adr_o[14]_pad ,
		\wbm_adr_o[15]_pad ,
		_w3282_,
		_w3283_
	);
	LUT4 #(
		.INIT('h0903)
	) name272 (
		\wbm_adr_o[16]_pad ,
		\wbm_adr_o[17]_pad ,
		_w3081_,
		_w3283_,
		_w3284_
	);
	LUT4 #(
		.INIT('h5333)
	) name273 (
		\pci_target_unit_del_sync_addr_out_reg[17]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001 ,
		_w3065_,
		_w3079_,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w3081_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w3284_,
		_w3286_,
		_w3287_
	);
	LUT4 #(
		.INIT('haccc)
	) name276 (
		\pci_target_unit_del_sync_addr_out_reg[18]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001 ,
		_w3065_,
		_w3079_,
		_w3288_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w3081_,
		_w3288_,
		_w3289_
	);
	LUT4 #(
		.INIT('h070f)
	) name278 (
		\wbm_adr_o[16]_pad ,
		\wbm_adr_o[17]_pad ,
		\wbm_adr_o[18]_pad ,
		_w3283_,
		_w3290_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\wbm_adr_o[17]_pad ,
		\wbm_adr_o[18]_pad ,
		_w3291_
	);
	LUT4 #(
		.INIT('h1333)
	) name280 (
		\wbm_adr_o[16]_pad ,
		_w3081_,
		_w3283_,
		_w3291_,
		_w3292_
	);
	LUT3 #(
		.INIT('hba)
	) name281 (
		_w3289_,
		_w3290_,
		_w3292_,
		_w3293_
	);
	LUT4 #(
		.INIT('h8000)
	) name282 (
		\wbm_adr_o[16]_pad ,
		\wbm_adr_o[19]_pad ,
		_w3283_,
		_w3291_,
		_w3294_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name283 (
		\wbm_adr_o[16]_pad ,
		\wbm_adr_o[19]_pad ,
		_w3283_,
		_w3291_,
		_w3295_
	);
	LUT4 #(
		.INIT('h5333)
	) name284 (
		\pci_target_unit_del_sync_addr_out_reg[19]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001 ,
		_w3065_,
		_w3079_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w3081_,
		_w3296_,
		_w3297_
	);
	LUT3 #(
		.INIT('h0e)
	) name286 (
		_w3081_,
		_w3295_,
		_w3297_,
		_w3298_
	);
	LUT4 #(
		.INIT('haccc)
	) name287 (
		\pci_target_unit_del_sync_addr_out_reg[20]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001 ,
		_w3065_,
		_w3079_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w3081_,
		_w3299_,
		_w3300_
	);
	LUT4 #(
		.INIT('hff12)
	) name289 (
		\wbm_adr_o[20]_pad ,
		_w3081_,
		_w3294_,
		_w3300_,
		_w3301_
	);
	LUT4 #(
		.INIT('haccc)
	) name290 (
		\pci_target_unit_del_sync_addr_out_reg[22]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001 ,
		_w3065_,
		_w3079_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w3081_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h070f)
	) name292 (
		\wbm_adr_o[20]_pad ,
		\wbm_adr_o[21]_pad ,
		\wbm_adr_o[22]_pad ,
		_w3294_,
		_w3304_
	);
	LUT4 #(
		.INIT('h8000)
	) name293 (
		\wbm_adr_o[19]_pad ,
		\wbm_adr_o[20]_pad ,
		\wbm_adr_o[21]_pad ,
		\wbm_adr_o[22]_pad ,
		_w3305_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		\wbm_adr_o[16]_pad ,
		_w3283_,
		_w3291_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w3081_,
		_w3306_,
		_w3307_
	);
	LUT3 #(
		.INIT('hba)
	) name296 (
		_w3303_,
		_w3304_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('haccc)
	) name297 (
		\pci_target_unit_del_sync_addr_out_reg[24]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001 ,
		_w3065_,
		_w3079_,
		_w3309_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w3081_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		\wbm_adr_o[23]_pad ,
		\wbm_adr_o[24]_pad ,
		_w3311_
	);
	LUT4 #(
		.INIT('h060c)
	) name300 (
		\wbm_adr_o[23]_pad ,
		\wbm_adr_o[24]_pad ,
		_w3081_,
		_w3306_,
		_w3312_
	);
	LUT2 #(
		.INIT('he)
	) name301 (
		_w3310_,
		_w3312_,
		_w3313_
	);
	LUT4 #(
		.INIT('h2111)
	) name302 (
		\wbm_adr_o[25]_pad ,
		_w3081_,
		_w3306_,
		_w3311_,
		_w3314_
	);
	LUT4 #(
		.INIT('h5333)
	) name303 (
		\pci_target_unit_del_sync_addr_out_reg[25]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001 ,
		_w3065_,
		_w3079_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w3081_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w3314_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\wbm_adr_o[25]_pad ,
		\wbm_adr_o[26]_pad ,
		_w3318_
	);
	LUT4 #(
		.INIT('h8000)
	) name307 (
		\wbm_adr_o[27]_pad ,
		_w3306_,
		_w3311_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name308 (
		\wbm_adr_o[27]_pad ,
		_w3306_,
		_w3311_,
		_w3318_,
		_w3320_
	);
	LUT4 #(
		.INIT('h5333)
	) name309 (
		\pci_target_unit_del_sync_addr_out_reg[27]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001 ,
		_w3065_,
		_w3079_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w3081_,
		_w3321_,
		_w3322_
	);
	LUT3 #(
		.INIT('h0e)
	) name311 (
		_w3081_,
		_w3320_,
		_w3322_,
		_w3323_
	);
	LUT4 #(
		.INIT('h0903)
	) name312 (
		\wbm_adr_o[20]_pad ,
		\wbm_adr_o[21]_pad ,
		_w3081_,
		_w3294_,
		_w3324_
	);
	LUT4 #(
		.INIT('h5333)
	) name313 (
		\pci_target_unit_del_sync_addr_out_reg[21]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001 ,
		_w3065_,
		_w3079_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w3081_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w3324_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('haccc)
	) name316 (
		\pci_target_unit_del_sync_addr_out_reg[29]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001 ,
		_w3065_,
		_w3079_,
		_w3328_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w3081_,
		_w3328_,
		_w3329_
	);
	LUT4 #(
		.INIT('h060c)
	) name318 (
		\wbm_adr_o[28]_pad ,
		\wbm_adr_o[29]_pad ,
		_w3081_,
		_w3319_,
		_w3330_
	);
	LUT2 #(
		.INIT('he)
	) name319 (
		_w3329_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h070f)
	) name320 (
		\wbm_adr_o[28]_pad ,
		\wbm_adr_o[29]_pad ,
		\wbm_adr_o[30]_pad ,
		_w3319_,
		_w3332_
	);
	LUT3 #(
		.INIT('h80)
	) name321 (
		\wbm_adr_o[28]_pad ,
		\wbm_adr_o[29]_pad ,
		\wbm_adr_o[30]_pad ,
		_w3333_
	);
	LUT3 #(
		.INIT('h15)
	) name322 (
		_w3081_,
		_w3319_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('haccc)
	) name323 (
		\pci_target_unit_del_sync_addr_out_reg[30]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001 ,
		_w3065_,
		_w3079_,
		_w3335_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w3081_,
		_w3335_,
		_w3336_
	);
	LUT3 #(
		.INIT('hf4)
	) name325 (
		_w3332_,
		_w3334_,
		_w3336_,
		_w3337_
	);
	LUT4 #(
		.INIT('h5333)
	) name326 (
		\pci_target_unit_del_sync_addr_out_reg[28]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001 ,
		_w3065_,
		_w3079_,
		_w3338_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		_w3081_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h00de)
	) name328 (
		\wbm_adr_o[28]_pad ,
		_w3081_,
		_w3319_,
		_w3339_,
		_w3340_
	);
	LUT4 #(
		.INIT('haccc)
	) name329 (
		\pci_target_unit_del_sync_addr_out_reg[31]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001 ,
		_w3065_,
		_w3079_,
		_w3341_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w3081_,
		_w3341_,
		_w3342_
	);
	LUT4 #(
		.INIT('h1222)
	) name331 (
		\wbm_adr_o[31]_pad ,
		_w3081_,
		_w3319_,
		_w3333_,
		_w3343_
	);
	LUT2 #(
		.INIT('he)
	) name332 (
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT4 #(
		.INIT('haa2a)
	) name333 (
		\wbm_dat_o[0]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3345_
	);
	LUT4 #(
		.INIT('h0080)
	) name334 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3346_
	);
	LUT2 #(
		.INIT('he)
	) name335 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('haa2a)
	) name336 (
		\wbm_dat_o[11]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3348_
	);
	LUT4 #(
		.INIT('h0080)
	) name337 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3349_
	);
	LUT2 #(
		.INIT('he)
	) name338 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('haa2a)
	) name339 (
		\wbm_dat_o[12]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3351_
	);
	LUT4 #(
		.INIT('h0080)
	) name340 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3352_
	);
	LUT2 #(
		.INIT('he)
	) name341 (
		_w3351_,
		_w3352_,
		_w3353_
	);
	LUT4 #(
		.INIT('haa2a)
	) name342 (
		\wbm_dat_o[13]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3354_
	);
	LUT4 #(
		.INIT('h0080)
	) name343 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3355_
	);
	LUT2 #(
		.INIT('he)
	) name344 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT4 #(
		.INIT('haa2a)
	) name345 (
		\wbm_dat_o[14]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3357_
	);
	LUT4 #(
		.INIT('h0080)
	) name346 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3358_
	);
	LUT2 #(
		.INIT('he)
	) name347 (
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT4 #(
		.INIT('haa2a)
	) name348 (
		\wbm_dat_o[15]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3360_
	);
	LUT4 #(
		.INIT('h0080)
	) name349 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3361_
	);
	LUT2 #(
		.INIT('he)
	) name350 (
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT4 #(
		.INIT('haa2a)
	) name351 (
		\wbm_dat_o[17]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3363_
	);
	LUT4 #(
		.INIT('h0080)
	) name352 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3364_
	);
	LUT2 #(
		.INIT('he)
	) name353 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT4 #(
		.INIT('haa2a)
	) name354 (
		\wbm_dat_o[16]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3366_
	);
	LUT4 #(
		.INIT('h0080)
	) name355 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3367_
	);
	LUT2 #(
		.INIT('he)
	) name356 (
		_w3366_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('haa2a)
	) name357 (
		\wbm_dat_o[18]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3369_
	);
	LUT4 #(
		.INIT('h0080)
	) name358 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3370_
	);
	LUT2 #(
		.INIT('he)
	) name359 (
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT4 #(
		.INIT('haa2a)
	) name360 (
		\wbm_dat_o[19]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3372_
	);
	LUT4 #(
		.INIT('h0080)
	) name361 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3373_
	);
	LUT2 #(
		.INIT('he)
	) name362 (
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('haa2a)
	) name363 (
		\wbm_dat_o[1]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3375_
	);
	LUT4 #(
		.INIT('h0080)
	) name364 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3376_
	);
	LUT2 #(
		.INIT('he)
	) name365 (
		_w3375_,
		_w3376_,
		_w3377_
	);
	LUT4 #(
		.INIT('haa2a)
	) name366 (
		\wbm_dat_o[20]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3378_
	);
	LUT4 #(
		.INIT('h0080)
	) name367 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3379_
	);
	LUT2 #(
		.INIT('he)
	) name368 (
		_w3378_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('haa2a)
	) name369 (
		\wbm_dat_o[21]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3381_
	);
	LUT4 #(
		.INIT('h0080)
	) name370 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3382_
	);
	LUT2 #(
		.INIT('he)
	) name371 (
		_w3381_,
		_w3382_,
		_w3383_
	);
	LUT4 #(
		.INIT('haa2a)
	) name372 (
		\wbm_dat_o[23]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3384_
	);
	LUT4 #(
		.INIT('h0080)
	) name373 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3385_
	);
	LUT2 #(
		.INIT('he)
	) name374 (
		_w3384_,
		_w3385_,
		_w3386_
	);
	LUT4 #(
		.INIT('haa2a)
	) name375 (
		\wbm_dat_o[24]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3387_
	);
	LUT4 #(
		.INIT('h0080)
	) name376 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3388_
	);
	LUT2 #(
		.INIT('he)
	) name377 (
		_w3387_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('haa2a)
	) name378 (
		\wbm_dat_o[25]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3390_
	);
	LUT4 #(
		.INIT('h0080)
	) name379 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3391_
	);
	LUT2 #(
		.INIT('he)
	) name380 (
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT4 #(
		.INIT('haa2a)
	) name381 (
		\wbm_dat_o[26]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3393_
	);
	LUT4 #(
		.INIT('h0080)
	) name382 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3394_
	);
	LUT2 #(
		.INIT('he)
	) name383 (
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT4 #(
		.INIT('haa2a)
	) name384 (
		\wbm_dat_o[28]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3396_
	);
	LUT4 #(
		.INIT('h0080)
	) name385 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3397_
	);
	LUT2 #(
		.INIT('he)
	) name386 (
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('haa2a)
	) name387 (
		\wbm_dat_o[27]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3399_
	);
	LUT4 #(
		.INIT('h0080)
	) name388 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3400_
	);
	LUT2 #(
		.INIT('he)
	) name389 (
		_w3399_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('haa2a)
	) name390 (
		\wbm_dat_o[29]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3402_
	);
	LUT4 #(
		.INIT('h0080)
	) name391 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3403_
	);
	LUT2 #(
		.INIT('he)
	) name392 (
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT4 #(
		.INIT('haa2a)
	) name393 (
		\wbm_dat_o[2]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3405_
	);
	LUT4 #(
		.INIT('h0080)
	) name394 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3406_
	);
	LUT2 #(
		.INIT('he)
	) name395 (
		_w3405_,
		_w3406_,
		_w3407_
	);
	LUT4 #(
		.INIT('haa2a)
	) name396 (
		\wbm_dat_o[30]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3408_
	);
	LUT4 #(
		.INIT('h0080)
	) name397 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3409_
	);
	LUT2 #(
		.INIT('he)
	) name398 (
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('haa2a)
	) name399 (
		\wbm_dat_o[3]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3411_
	);
	LUT4 #(
		.INIT('h0080)
	) name400 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3412_
	);
	LUT2 #(
		.INIT('he)
	) name401 (
		_w3411_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('haa2a)
	) name402 (
		\wbm_dat_o[4]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3414_
	);
	LUT4 #(
		.INIT('h0080)
	) name403 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3415_
	);
	LUT2 #(
		.INIT('he)
	) name404 (
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT4 #(
		.INIT('haa2a)
	) name405 (
		\wbm_dat_o[31]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3417_
	);
	LUT4 #(
		.INIT('h0080)
	) name406 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3418_
	);
	LUT2 #(
		.INIT('he)
	) name407 (
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('haa2a)
	) name408 (
		\wbm_dat_o[5]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3420_
	);
	LUT4 #(
		.INIT('h0080)
	) name409 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3421_
	);
	LUT2 #(
		.INIT('he)
	) name410 (
		_w3420_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('haa2a)
	) name411 (
		\wbm_dat_o[6]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3423_
	);
	LUT4 #(
		.INIT('h0080)
	) name412 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3424_
	);
	LUT2 #(
		.INIT('he)
	) name413 (
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT4 #(
		.INIT('haa2a)
	) name414 (
		\wbm_dat_o[7]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3426_
	);
	LUT4 #(
		.INIT('h0080)
	) name415 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3427_
	);
	LUT2 #(
		.INIT('he)
	) name416 (
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('haa2a)
	) name417 (
		\wbm_dat_o[8]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3429_
	);
	LUT4 #(
		.INIT('h0080)
	) name418 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3430_
	);
	LUT2 #(
		.INIT('he)
	) name419 (
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('haa2a)
	) name420 (
		\wbm_dat_o[9]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3432_
	);
	LUT4 #(
		.INIT('h0080)
	) name421 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w3433_
	);
	LUT2 #(
		.INIT('he)
	) name422 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT4 #(
		.INIT('h1211)
	) name423 (
		\wbm_adr_o[10]_pad ,
		_w3081_,
		_w3276_,
		_w3280_,
		_w3435_
	);
	LUT4 #(
		.INIT('h5333)
	) name424 (
		\pci_target_unit_del_sync_addr_out_reg[10]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001 ,
		_w3065_,
		_w3079_,
		_w3436_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w3081_,
		_w3436_,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w3435_,
		_w3437_,
		_w3438_
	);
	LUT4 #(
		.INIT('haccc)
	) name427 (
		\pci_target_unit_del_sync_addr_out_reg[11]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]/P0001 ,
		_w3065_,
		_w3079_,
		_w3439_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w3081_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h3133)
	) name429 (
		\wbm_adr_o[10]_pad ,
		\wbm_adr_o[11]_pad ,
		_w3276_,
		_w3280_,
		_w3441_
	);
	LUT4 #(
		.INIT('h4555)
	) name430 (
		_w3081_,
		_w3276_,
		_w3280_,
		_w3281_,
		_w3442_
	);
	LUT3 #(
		.INIT('hba)
	) name431 (
		_w3440_,
		_w3441_,
		_w3442_,
		_w3443_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name432 (
		\wbm_adr_o[12]_pad ,
		_w3276_,
		_w3280_,
		_w3281_,
		_w3444_
	);
	LUT4 #(
		.INIT('h5333)
	) name433 (
		\pci_target_unit_del_sync_addr_out_reg[12]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]/P0001 ,
		_w3065_,
		_w3079_,
		_w3445_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w3081_,
		_w3445_,
		_w3446_
	);
	LUT3 #(
		.INIT('h0e)
	) name435 (
		_w3081_,
		_w3444_,
		_w3446_,
		_w3447_
	);
	LUT4 #(
		.INIT('h5333)
	) name436 (
		\pci_target_unit_del_sync_addr_out_reg[13]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]/P0001 ,
		_w3065_,
		_w3079_,
		_w3448_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		_w3081_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h00de)
	) name438 (
		\wbm_adr_o[13]_pad ,
		_w3081_,
		_w3282_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h78f0)
	) name439 (
		\wbm_adr_o[13]_pad ,
		\wbm_adr_o[14]_pad ,
		\wbm_adr_o[15]_pad ,
		_w3282_,
		_w3451_
	);
	LUT4 #(
		.INIT('h5333)
	) name440 (
		\pci_target_unit_del_sync_addr_out_reg[15]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]/P0001 ,
		_w3065_,
		_w3079_,
		_w3452_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w3081_,
		_w3452_,
		_w3453_
	);
	LUT3 #(
		.INIT('h0e)
	) name442 (
		_w3081_,
		_w3451_,
		_w3453_,
		_w3454_
	);
	LUT4 #(
		.INIT('h5333)
	) name443 (
		\pci_target_unit_del_sync_addr_out_reg[16]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]/P0001 ,
		_w3065_,
		_w3079_,
		_w3455_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w3081_,
		_w3455_,
		_w3456_
	);
	LUT4 #(
		.INIT('h00de)
	) name445 (
		\wbm_adr_o[16]_pad ,
		_w3081_,
		_w3283_,
		_w3456_,
		_w3457_
	);
	LUT4 #(
		.INIT('h0903)
	) name446 (
		\wbm_adr_o[13]_pad ,
		\wbm_adr_o[14]_pad ,
		_w3081_,
		_w3282_,
		_w3458_
	);
	LUT4 #(
		.INIT('h5333)
	) name447 (
		\pci_target_unit_del_sync_addr_out_reg[14]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]/P0001 ,
		_w3065_,
		_w3079_,
		_w3459_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w3081_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w3458_,
		_w3460_,
		_w3461_
	);
	LUT4 #(
		.INIT('h5333)
	) name450 (
		\pci_target_unit_del_sync_addr_out_reg[23]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]/P0001 ,
		_w3065_,
		_w3079_,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w3081_,
		_w3462_,
		_w3463_
	);
	LUT4 #(
		.INIT('h00de)
	) name452 (
		\wbm_adr_o[23]_pad ,
		_w3081_,
		_w3306_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name453 (
		\wbm_adr_o[25]_pad ,
		\wbm_adr_o[26]_pad ,
		_w3306_,
		_w3311_,
		_w3465_
	);
	LUT4 #(
		.INIT('h5333)
	) name454 (
		\pci_target_unit_del_sync_addr_out_reg[26]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]/P0001 ,
		_w3065_,
		_w3079_,
		_w3466_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w3081_,
		_w3466_,
		_w3467_
	);
	LUT3 #(
		.INIT('h0e)
	) name456 (
		_w3081_,
		_w3465_,
		_w3467_,
		_w3468_
	);
	LUT4 #(
		.INIT('ha080)
	) name457 (
		\wbm_adr_o[2]_pad ,
		_w3068_,
		_w3057_,
		_w3050_,
		_w3469_
	);
	LUT4 #(
		.INIT('h5a6a)
	) name458 (
		\wbm_adr_o[2]_pad ,
		_w3068_,
		_w3057_,
		_w3050_,
		_w3470_
	);
	LUT4 #(
		.INIT('h5333)
	) name459 (
		\pci_target_unit_del_sync_addr_out_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]/P0001 ,
		_w3065_,
		_w3079_,
		_w3471_
	);
	LUT3 #(
		.INIT('h4e)
	) name460 (
		_w3081_,
		_w3470_,
		_w3471_,
		_w3472_
	);
	LUT4 #(
		.INIT('h5333)
	) name461 (
		\pci_target_unit_del_sync_addr_out_reg[3]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]/P0001 ,
		_w3065_,
		_w3079_,
		_w3473_
	);
	LUT4 #(
		.INIT('h12de)
	) name462 (
		\wbm_adr_o[3]_pad ,
		_w3081_,
		_w3469_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h0903)
	) name463 (
		\wbm_adr_o[3]_pad ,
		\wbm_adr_o[4]_pad ,
		_w3081_,
		_w3469_,
		_w3475_
	);
	LUT4 #(
		.INIT('h5333)
	) name464 (
		\pci_target_unit_del_sync_addr_out_reg[4]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]/P0001 ,
		_w3065_,
		_w3079_,
		_w3476_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w3081_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w3475_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('h8000)
	) name467 (
		\wbm_adr_o[3]_pad ,
		\wbm_adr_o[4]_pad ,
		\wbm_adr_o[5]_pad ,
		_w3469_,
		_w3479_
	);
	LUT4 #(
		.INIT('h78f0)
	) name468 (
		\wbm_adr_o[3]_pad ,
		\wbm_adr_o[4]_pad ,
		\wbm_adr_o[5]_pad ,
		_w3469_,
		_w3480_
	);
	LUT4 #(
		.INIT('h5333)
	) name469 (
		\pci_target_unit_del_sync_addr_out_reg[5]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]/P0001 ,
		_w3065_,
		_w3079_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w3081_,
		_w3481_,
		_w3482_
	);
	LUT3 #(
		.INIT('h0e)
	) name471 (
		_w3081_,
		_w3480_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('h0903)
	) name472 (
		\wbm_adr_o[6]_pad ,
		\wbm_adr_o[7]_pad ,
		_w3081_,
		_w3479_,
		_w3484_
	);
	LUT4 #(
		.INIT('h5333)
	) name473 (
		\pci_target_unit_del_sync_addr_out_reg[7]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]/P0001 ,
		_w3065_,
		_w3079_,
		_w3485_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w3081_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w3484_,
		_w3486_,
		_w3487_
	);
	LUT4 #(
		.INIT('h5333)
	) name476 (
		\pci_target_unit_del_sync_addr_out_reg[6]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]/P0001 ,
		_w3065_,
		_w3079_,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w3081_,
		_w3488_,
		_w3489_
	);
	LUT4 #(
		.INIT('h00de)
	) name478 (
		\wbm_adr_o[6]_pad ,
		_w3081_,
		_w3479_,
		_w3489_,
		_w3490_
	);
	LUT4 #(
		.INIT('h78f0)
	) name479 (
		\wbm_adr_o[6]_pad ,
		\wbm_adr_o[7]_pad ,
		\wbm_adr_o[8]_pad ,
		_w3479_,
		_w3491_
	);
	LUT4 #(
		.INIT('h5333)
	) name480 (
		\pci_target_unit_del_sync_addr_out_reg[8]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]/P0001 ,
		_w3065_,
		_w3079_,
		_w3492_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		_w3081_,
		_w3492_,
		_w3493_
	);
	LUT3 #(
		.INIT('h0e)
	) name482 (
		_w3081_,
		_w3491_,
		_w3493_,
		_w3494_
	);
	LUT4 #(
		.INIT('haccc)
	) name483 (
		\pci_target_unit_del_sync_addr_out_reg[9]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]/P0001 ,
		_w3065_,
		_w3079_,
		_w3495_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		_w3081_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('h1333)
	) name485 (
		\wbm_adr_o[6]_pad ,
		\wbm_adr_o[9]_pad ,
		_w3278_,
		_w3479_,
		_w3497_
	);
	LUT3 #(
		.INIT('h45)
	) name486 (
		_w3081_,
		_w3276_,
		_w3280_,
		_w3498_
	);
	LUT3 #(
		.INIT('hba)
	) name487 (
		_w3496_,
		_w3497_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 ,
		_w3500_
	);
	LUT4 #(
		.INIT('h8000)
	) name489 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 ,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		_w3500_,
		_w3501_,
		_w3502_
	);
	LUT3 #(
		.INIT('hb0)
	) name491 (
		_w3151_,
		_w3170_,
		_w3502_,
		_w3503_
	);
	LUT4 #(
		.INIT('h8a00)
	) name492 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 ,
		_w3151_,
		_w3170_,
		_w3502_,
		_w3504_
	);
	LUT4 #(
		.INIT('h060a)
	) name493 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3134_,
		_w3504_,
		_w3505_
	);
	LUT3 #(
		.INIT('h80)
	) name494 (
		\wbs_adr_i[10]_pad ,
		_w3131_,
		_w3133_,
		_w3506_
	);
	LUT2 #(
		.INIT('he)
	) name495 (
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT3 #(
		.INIT('h80)
	) name496 (
		\wbs_adr_i[11]_pad ,
		_w3131_,
		_w3133_,
		_w3508_
	);
	LUT4 #(
		.INIT('h1333)
	) name497 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3504_,
		_w3509_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 ,
		_w3510_
	);
	LUT3 #(
		.INIT('h80)
	) name499 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3504_,
		_w3510_,
		_w3511_
	);
	LUT4 #(
		.INIT('h1333)
	) name500 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3134_,
		_w3504_,
		_w3510_,
		_w3512_
	);
	LUT3 #(
		.INIT('hba)
	) name501 (
		_w3508_,
		_w3509_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('h8000)
	) name502 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3504_,
		_w3510_,
		_w3514_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name503 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\wbs_adr_i[12]_pad ,
		_w3134_,
		_w3511_,
		_w3515_
	);
	LUT3 #(
		.INIT('h80)
	) name504 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w3510_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w3504_,
		_w3517_,
		_w3518_
	);
	LUT4 #(
		.INIT('h3301)
	) name507 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		_w3134_,
		_w3514_,
		_w3518_,
		_w3519_
	);
	LUT3 #(
		.INIT('h40)
	) name508 (
		\wbs_adr_i[13]_pad ,
		_w3131_,
		_w3133_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		_w3522_
	);
	LUT3 #(
		.INIT('h80)
	) name511 (
		_w3504_,
		_w3517_,
		_w3522_,
		_w3523_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name512 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		_w3504_,
		_w3517_,
		_w3524_
	);
	LUT3 #(
		.INIT('hb8)
	) name513 (
		\wbs_adr_i[15]_pad ,
		_w3134_,
		_w3524_,
		_w3525_
	);
	LUT4 #(
		.INIT('h1222)
	) name514 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		_w3134_,
		_w3504_,
		_w3517_,
		_w3526_
	);
	LUT3 #(
		.INIT('h80)
	) name515 (
		\wbs_adr_i[14]_pad ,
		_w3131_,
		_w3133_,
		_w3527_
	);
	LUT2 #(
		.INIT('he)
	) name516 (
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT4 #(
		.INIT('h8000)
	) name517 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		_w3504_,
		_w3517_,
		_w3522_,
		_w3529_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name518 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\wbs_adr_i[16]_pad ,
		_w3134_,
		_w3523_,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		_w3531_
	);
	LUT4 #(
		.INIT('h8000)
	) name520 (
		_w3504_,
		_w3517_,
		_w3522_,
		_w3531_,
		_w3532_
	);
	LUT4 #(
		.INIT('h0903)
	) name521 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		_w3134_,
		_w3523_,
		_w3533_
	);
	LUT3 #(
		.INIT('h40)
	) name522 (
		\wbs_adr_i[17]_pad ,
		_w3131_,
		_w3133_,
		_w3534_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name524 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\wbs_adr_i[18]_pad ,
		_w3134_,
		_w3532_,
		_w3536_
	);
	LUT3 #(
		.INIT('h80)
	) name525 (
		\wbs_adr_i[19]_pad ,
		_w3131_,
		_w3133_,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		_w3538_
	);
	LUT4 #(
		.INIT('h060c)
	) name527 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		_w3134_,
		_w3532_,
		_w3539_
	);
	LUT2 #(
		.INIT('he)
	) name528 (
		_w3537_,
		_w3539_,
		_w3540_
	);
	LUT4 #(
		.INIT('h1222)
	) name529 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		_w3134_,
		_w3532_,
		_w3538_,
		_w3541_
	);
	LUT3 #(
		.INIT('h80)
	) name530 (
		\wbs_adr_i[20]_pad ,
		_w3131_,
		_w3133_,
		_w3542_
	);
	LUT2 #(
		.INIT('he)
	) name531 (
		_w3541_,
		_w3542_,
		_w3543_
	);
	LUT3 #(
		.INIT('h80)
	) name532 (
		\wbs_adr_i[21]_pad ,
		_w3131_,
		_w3133_,
		_w3544_
	);
	LUT4 #(
		.INIT('h8000)
	) name533 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		_w3545_
	);
	LUT4 #(
		.INIT('h1222)
	) name534 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		_w3134_,
		_w3529_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('he)
	) name535 (
		_w3544_,
		_w3546_,
		_w3547_
	);
	LUT4 #(
		.INIT('h8000)
	) name536 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		_w3548_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w3538_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('h8000)
	) name538 (
		_w3504_,
		_w3517_,
		_w3522_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name539 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\wbs_adr_i[22]_pad ,
		_w3134_,
		_w3550_,
		_w3551_
	);
	LUT3 #(
		.INIT('h80)
	) name540 (
		\wbs_adr_i[23]_pad ,
		_w3131_,
		_w3133_,
		_w3552_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name542 (
		_w3545_,
		_w3553_,
		_w3554_
	);
	LUT4 #(
		.INIT('h1222)
	) name543 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		_w3134_,
		_w3529_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('he)
	) name544 (
		_w3552_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		_w3557_
	);
	LUT3 #(
		.INIT('h80)
	) name546 (
		_w3538_,
		_w3548_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('h8000)
	) name547 (
		_w3504_,
		_w3517_,
		_w3522_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		_w3561_
	);
	LUT3 #(
		.INIT('h80)
	) name550 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		_w3550_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('h888b)
	) name551 (
		\wbs_adr_i[24]_pad ,
		_w3134_,
		_w3560_,
		_w3562_,
		_w3563_
	);
	LUT3 #(
		.INIT('h80)
	) name552 (
		\wbs_adr_i[25]_pad ,
		_w3131_,
		_w3133_,
		_w3564_
	);
	LUT3 #(
		.INIT('h80)
	) name553 (
		_w3545_,
		_w3553_,
		_w3561_,
		_w3565_
	);
	LUT4 #(
		.INIT('h1222)
	) name554 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		_w3134_,
		_w3529_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('he)
	) name555 (
		_w3564_,
		_w3566_,
		_w3567_
	);
	LUT3 #(
		.INIT('h80)
	) name556 (
		\wbs_adr_i[26]_pad ,
		_w3131_,
		_w3133_,
		_w3568_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		_w3569_
	);
	LUT4 #(
		.INIT('h1222)
	) name558 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		_w3134_,
		_w3559_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('he)
	) name559 (
		_w3568_,
		_w3570_,
		_w3571_
	);
	LUT3 #(
		.INIT('h80)
	) name560 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		_w3573_
	);
	LUT3 #(
		.INIT('h80)
	) name562 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		_w3574_
	);
	LUT4 #(
		.INIT('h8000)
	) name563 (
		_w3545_,
		_w3553_,
		_w3572_,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h8000)
	) name564 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		_w3504_,
		_w3517_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name565 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\wbs_adr_i[27]_pad ,
		_w3134_,
		_w3576_,
		_w3577_
	);
	LUT3 #(
		.INIT('h80)
	) name566 (
		\wbs_adr_i[28]_pad ,
		_w3131_,
		_w3133_,
		_w3578_
	);
	LUT4 #(
		.INIT('h8000)
	) name567 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		_w3579_
	);
	LUT4 #(
		.INIT('h1222)
	) name568 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		_w3134_,
		_w3559_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('he)
	) name569 (
		_w3578_,
		_w3580_,
		_w3581_
	);
	LUT3 #(
		.INIT('h8a)
	) name570 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		_w3151_,
		_w3170_,
		_w3582_
	);
	LUT4 #(
		.INIT('h1211)
	) name571 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		_w3134_,
		_w3151_,
		_w3170_,
		_w3583_
	);
	LUT3 #(
		.INIT('h80)
	) name572 (
		\wbs_adr_i[2]_pad ,
		_w3131_,
		_w3133_,
		_w3584_
	);
	LUT2 #(
		.INIT('he)
	) name573 (
		_w3583_,
		_w3584_,
		_w3585_
	);
	LUT3 #(
		.INIT('h80)
	) name574 (
		\wbs_adr_i[30]_pad ,
		_w3131_,
		_w3133_,
		_w3586_
	);
	LUT3 #(
		.INIT('h80)
	) name575 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		_w3587_
	);
	LUT3 #(
		.INIT('h80)
	) name576 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		_w3588_
	);
	LUT3 #(
		.INIT('h80)
	) name577 (
		_w3569_,
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT4 #(
		.INIT('h1222)
	) name578 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 ,
		_w3134_,
		_w3550_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('he)
	) name579 (
		_w3586_,
		_w3590_,
		_w3591_
	);
	LUT3 #(
		.INIT('h80)
	) name580 (
		\wbs_adr_i[29]_pad ,
		_w3131_,
		_w3133_,
		_w3592_
	);
	LUT3 #(
		.INIT('h80)
	) name581 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		_w3593_
	);
	LUT3 #(
		.INIT('h80)
	) name582 (
		_w3573_,
		_w3587_,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w3565_,
		_w3594_,
		_w3595_
	);
	LUT4 #(
		.INIT('h1222)
	) name584 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		_w3134_,
		_w3514_,
		_w3595_,
		_w3596_
	);
	LUT2 #(
		.INIT('he)
	) name585 (
		_w3592_,
		_w3596_,
		_w3597_
	);
	LUT3 #(
		.INIT('h80)
	) name586 (
		\wbs_adr_i[31]_pad ,
		_w3131_,
		_w3133_,
		_w3598_
	);
	LUT4 #(
		.INIT('h8000)
	) name587 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 ,
		_w3599_
	);
	LUT4 #(
		.INIT('h1222)
	) name588 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w3134_,
		_w3576_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('he)
	) name589 (
		_w3598_,
		_w3600_,
		_w3601_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name590 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\wbs_adr_i[3]_pad ,
		_w3134_,
		_w3582_,
		_w3602_
	);
	LUT4 #(
		.INIT('h8a00)
	) name591 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		_w3151_,
		_w3170_,
		_w3500_,
		_w3603_
	);
	LUT4 #(
		.INIT('h060c)
	) name592 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 ,
		_w3134_,
		_w3582_,
		_w3604_
	);
	LUT3 #(
		.INIT('h80)
	) name593 (
		\wbs_adr_i[4]_pad ,
		_w3131_,
		_w3133_,
		_w3605_
	);
	LUT2 #(
		.INIT('he)
	) name594 (
		_w3604_,
		_w3605_,
		_w3606_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name595 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\wbs_adr_i[5]_pad ,
		_w3134_,
		_w3603_,
		_w3607_
	);
	LUT4 #(
		.INIT('h060c)
	) name596 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		_w3134_,
		_w3603_,
		_w3608_
	);
	LUT3 #(
		.INIT('h80)
	) name597 (
		\wbs_adr_i[6]_pad ,
		_w3131_,
		_w3133_,
		_w3609_
	);
	LUT2 #(
		.INIT('he)
	) name598 (
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT3 #(
		.INIT('h80)
	) name599 (
		\wbs_adr_i[7]_pad ,
		_w3131_,
		_w3133_,
		_w3611_
	);
	LUT4 #(
		.INIT('h070f)
	) name600 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 ,
		_w3603_,
		_w3612_
	);
	LUT4 #(
		.INIT('h1055)
	) name601 (
		_w3134_,
		_w3151_,
		_w3170_,
		_w3502_,
		_w3613_
	);
	LUT3 #(
		.INIT('hba)
	) name602 (
		_w3611_,
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name603 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 ,
		\wbs_adr_i[8]_pad ,
		_w3134_,
		_w3503_,
		_w3615_
	);
	LUT4 #(
		.INIT('hc5ca)
	) name604 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		\wbs_adr_i[9]_pad ,
		_w3134_,
		_w3504_,
		_w3616_
	);
	LUT4 #(
		.INIT('h4000)
	) name605 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131 ,
		wbs_cyc_i_pad,
		wbs_stb_i_pad,
		wbs_we_i_pad,
		_w3617_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w3131_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h002a)
	) name607 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg/NET0131 ,
		_w3147_,
		_w3150_,
		_w3178_,
		_w3619_
	);
	LUT4 #(
		.INIT('h2000)
	) name608 (
		_w3177_,
		_w3151_,
		_w3170_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('he)
	) name609 (
		_w3618_,
		_w3620_,
		_w3621_
	);
	LUT4 #(
		.INIT('h2a00)
	) name610 (
		_w3078_,
		_w3065_,
		_w3079_,
		_w3080_,
		_w3622_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]/P0001 ,
		_w3622_,
		_w3623_
	);
	LUT4 #(
		.INIT('h4000)
	) name612 (
		\pci_target_unit_del_sync_bc_out_reg[3]/NET0131 ,
		_w3078_,
		_w3065_,
		_w3079_,
		_w3624_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\pci_target_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[2]/NET0131 ,
		_w3625_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name614 (
		\wbm_adr_o[0]_pad ,
		_w3081_,
		_w3624_,
		_w3625_,
		_w3626_
	);
	LUT2 #(
		.INIT('hb)
	) name615 (
		_w3623_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]/P0001 ,
		_w3622_,
		_w3628_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\pci_target_unit_del_sync_addr_out_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[2]/NET0131 ,
		_w3629_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name618 (
		\wbm_adr_o[1]_pad ,
		_w3081_,
		_w3624_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('hb)
	) name619 (
		_w3628_,
		_w3630_,
		_w3631_
	);
	LUT4 #(
		.INIT('h8421)
	) name620 (
		\pci_target_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		\pci_target_unit_fifos_outGreyCount_reg[1]/NET0131 ,
		\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]/NET0131 ,
		\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]/NET0131 ,
		_w3632_
	);
	LUT4 #(
		.INIT('h0002)
	) name621 (
		\pci_target_unit_wishbone_master_burst_chopped_reg/NET0131 ,
		wbm_ack_i_pad,
		wbm_err_i_pad,
		wbm_rty_i_pad,
		_w3633_
	);
	LUT3 #(
		.INIT('h32)
	) name622 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w3135_,
		_w3635_,
		_w3636_
	);
	LUT3 #(
		.INIT('h20)
	) name625 (
		_w3147_,
		_w3150_,
		_w3636_,
		_w3637_
	);
	LUT3 #(
		.INIT('h70)
	) name626 (
		_w3163_,
		_w3164_,
		_w3635_,
		_w3638_
	);
	LUT4 #(
		.INIT('h50d0)
	) name627 (
		_w3145_,
		_w3140_,
		_w3166_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131 ,
		_w3639_,
		_w3640_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name629 (
		\wishbone_slave_unit_del_sync_req_comp_pending_sample_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131 ,
		_w3637_,
		_w3640_,
		_w3641_
	);
	LUT4 #(
		.INIT('h0105)
	) name630 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131 ,
		_w3642_
	);
	LUT3 #(
		.INIT('h08)
	) name631 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		_w3247_,
		_w3642_,
		_w3643_
	);
	LUT4 #(
		.INIT('h00ba)
	) name632 (
		_w3211_,
		_w3251_,
		_w3259_,
		_w3643_,
		_w3644_
	);
	LUT4 #(
		.INIT('h0100)
	) name633 (
		\pci_target_unit_pci_target_sm_backoff_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w3645_
	);
	LUT3 #(
		.INIT('h80)
	) name634 (
		_w3044_,
		_w3206_,
		_w3645_,
		_w3646_
	);
	LUT3 #(
		.INIT('hb0)
	) name635 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3261_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		_w3648_
	);
	LUT3 #(
		.INIT('h10)
	) name637 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3649_
	);
	LUT2 #(
		.INIT('h2)
	) name638 (
		_w3268_,
		_w3649_,
		_w3650_
	);
	LUT4 #(
		.INIT('hbf00)
	) name639 (
		_w3261_,
		_w3266_,
		_w3648_,
		_w3650_,
		_w3651_
	);
	LUT4 #(
		.INIT('h0207)
	) name640 (
		\output_backup_frame_en_out_reg/NET0131 ,
		\output_backup_frame_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		pci_frame_i_pad,
		_w3652_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w3208_,
		_w3652_,
		_w3653_
	);
	LUT3 #(
		.INIT('h0d)
	) name642 (
		_w3223_,
		_w3651_,
		_w3653_,
		_w3654_
	);
	LUT3 #(
		.INIT('hb0)
	) name643 (
		_w3644_,
		_w3647_,
		_w3654_,
		_w3655_
	);
	LUT3 #(
		.INIT('h45)
	) name644 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		_w3151_,
		_w3170_,
		_w3656_
	);
	LUT3 #(
		.INIT('hca)
	) name645 (
		\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_done_reg_reg/NET0131 ,
		_w3657_
	);
	LUT3 #(
		.INIT('h40)
	) name646 (
		_w3637_,
		_w3640_,
		_w3657_,
		_w3658_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg/NET0131 ,
		wbs_stb_i_pad,
		_w3659_
	);
	LUT3 #(
		.INIT('hfb)
	) name648 (
		_w3151_,
		_w3170_,
		_w3659_,
		_w3660_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w3135_,
		_w3635_,
		_w3661_
	);
	LUT3 #(
		.INIT('h20)
	) name650 (
		_w3147_,
		_w3150_,
		_w3661_,
		_w3662_
	);
	LUT4 #(
		.INIT('ha020)
	) name651 (
		_w3145_,
		_w3140_,
		_w3166_,
		_w3638_,
		_w3663_
	);
	LUT4 #(
		.INIT('h0002)
	) name652 (
		\configuration_wb_init_complete_out_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_c_state_reg[2]/NET0131 ,
		_w3664_
	);
	LUT3 #(
		.INIT('he0)
	) name653 (
		_w3140_,
		_w3135_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w3663_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('hb)
	) name655 (
		_w3662_,
		_w3666_,
		_w3667_
	);
	LUT3 #(
		.INIT('h02)
	) name656 (
		_w3147_,
		_w3150_,
		_w3636_,
		_w3668_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w3160_,
		_w3663_,
		_w3669_
	);
	LUT2 #(
		.INIT('hb)
	) name658 (
		_w3668_,
		_w3669_,
		_w3670_
	);
	LUT3 #(
		.INIT('h04)
	) name659 (
		\pci_target_unit_pci_target_sm_backoff_reg/NET0131 ,
		_w3210_,
		_w3263_,
		_w3671_
	);
	LUT4 #(
		.INIT('h0207)
	) name660 (
		\output_backup_frame_en_out_reg/NET0131 ,
		\output_backup_frame_out_reg/NET0131 ,
		\output_backup_stop_out_reg/NET0131 ,
		pci_frame_i_pad,
		_w3672_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w3224_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w3269_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w3671_,
		_w3674_,
		_w3675_
	);
	LUT3 #(
		.INIT('h27)
	) name664 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg/NET0131 ,
		wbs_stb_i_pad,
		_w3177_,
		_w3676_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		\output_backup_devsel_out_reg/NET0131 ,
		_w3224_,
		_w3677_
	);
	LUT4 #(
		.INIT('hbf00)
	) name666 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3208_,
		_w3261_,
		_w3645_,
		_w3678_
	);
	LUT3 #(
		.INIT('ha8)
	) name667 (
		_w3206_,
		_w3677_,
		_w3678_,
		_w3679_
	);
	LUT3 #(
		.INIT('h20)
	) name668 (
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_progress_reg/NET0131 ,
		_w3680_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name669 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3223_,
		_w3261_,
		_w3680_,
		_w3681_
	);
	LUT3 #(
		.INIT('h28)
	) name670 (
		\configuration_pci_am1_reg[10]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		_w3682_
	);
	LUT3 #(
		.INIT('h28)
	) name671 (
		\configuration_pci_am1_reg[21]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		_w3683_
	);
	LUT3 #(
		.INIT('h28)
	) name672 (
		\configuration_pci_am1_reg[11]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		_w3684_
	);
	LUT3 #(
		.INIT('h01)
	) name673 (
		_w3683_,
		_w3684_,
		_w3682_,
		_w3685_
	);
	LUT3 #(
		.INIT('h28)
	) name674 (
		\configuration_pci_am1_reg[22]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[22]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		_w3686_
	);
	LUT3 #(
		.INIT('h28)
	) name675 (
		\configuration_pci_am1_reg[19]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		_w3687_
	);
	LUT3 #(
		.INIT('h28)
	) name676 (
		\configuration_pci_am1_reg[26]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		_w3688_
	);
	LUT3 #(
		.INIT('h28)
	) name677 (
		\configuration_pci_am1_reg[23]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		_w3689_
	);
	LUT4 #(
		.INIT('h0001)
	) name678 (
		_w3686_,
		_w3687_,
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT3 #(
		.INIT('h28)
	) name679 (
		\configuration_pci_am1_reg[17]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[17]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		_w3691_
	);
	LUT3 #(
		.INIT('h28)
	) name680 (
		\configuration_pci_am1_reg[24]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		_w3692_
	);
	LUT3 #(
		.INIT('h28)
	) name681 (
		\configuration_pci_am1_reg[20]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		_w3693_
	);
	LUT3 #(
		.INIT('h28)
	) name682 (
		\configuration_pci_am1_reg[15]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		_w3694_
	);
	LUT4 #(
		.INIT('h0001)
	) name683 (
		_w3691_,
		_w3692_,
		_w3693_,
		_w3694_,
		_w3695_
	);
	LUT3 #(
		.INIT('h80)
	) name684 (
		_w3685_,
		_w3690_,
		_w3695_,
		_w3696_
	);
	LUT4 #(
		.INIT('h0080)
	) name685 (
		\configuration_command_bit2_0_reg[0]/NET0131 ,
		\configuration_init_complete_reg/NET0131 ,
		\configuration_pci_am1_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3697_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3698_
	);
	LUT4 #(
		.INIT('h0090)
	) name687 (
		\configuration_pci_ba1_bit31_8_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		_w3697_,
		_w3699_,
		_w3700_
	);
	LUT3 #(
		.INIT('h28)
	) name689 (
		\configuration_pci_am1_reg[27]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		_w3701_
	);
	LUT3 #(
		.INIT('h28)
	) name690 (
		\configuration_pci_am1_reg[8]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[8]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		_w3702_
	);
	LUT3 #(
		.INIT('h28)
	) name691 (
		\configuration_pci_am1_reg[29]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[29]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		_w3703_
	);
	LUT3 #(
		.INIT('h28)
	) name692 (
		\configuration_pci_am1_reg[9]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[9]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		_w3704_
	);
	LUT4 #(
		.INIT('h0001)
	) name693 (
		_w3701_,
		_w3702_,
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT3 #(
		.INIT('h28)
	) name694 (
		\configuration_pci_am1_reg[18]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		_w3706_
	);
	LUT3 #(
		.INIT('h28)
	) name695 (
		\configuration_pci_am1_reg[28]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[28]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		_w3707_
	);
	LUT3 #(
		.INIT('h28)
	) name696 (
		\configuration_pci_am1_reg[12]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		_w3708_
	);
	LUT3 #(
		.INIT('h28)
	) name697 (
		\configuration_pci_am1_reg[14]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		_w3709_
	);
	LUT4 #(
		.INIT('h0001)
	) name698 (
		_w3706_,
		_w3707_,
		_w3708_,
		_w3709_,
		_w3710_
	);
	LUT3 #(
		.INIT('h28)
	) name699 (
		\configuration_pci_am1_reg[25]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		_w3711_
	);
	LUT3 #(
		.INIT('h28)
	) name700 (
		\configuration_pci_am1_reg[16]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		_w3712_
	);
	LUT3 #(
		.INIT('h28)
	) name701 (
		\configuration_pci_am1_reg[13]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		_w3713_
	);
	LUT3 #(
		.INIT('h28)
	) name702 (
		\configuration_pci_am1_reg[30]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		_w3714_
	);
	LUT4 #(
		.INIT('h0001)
	) name703 (
		_w3711_,
		_w3712_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT4 #(
		.INIT('h8000)
	) name704 (
		_w3700_,
		_w3710_,
		_w3715_,
		_w3705_,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		_w3696_,
		_w3716_,
		_w3717_
	);
	LUT4 #(
		.INIT('haf23)
	) name706 (
		\configuration_pci_ba0_bit31_8_reg[16]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		_w3718_
	);
	LUT4 #(
		.INIT('h8caf)
	) name707 (
		\configuration_pci_ba0_bit31_8_reg[20]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		_w3719_
	);
	LUT4 #(
		.INIT('hf531)
	) name708 (
		\configuration_pci_ba0_bit31_8_reg[14]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		_w3720_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name709 (
		\configuration_pci_ba0_bit31_8_reg[13]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		_w3721_
	);
	LUT4 #(
		.INIT('h8000)
	) name710 (
		_w3720_,
		_w3721_,
		_w3718_,
		_w3719_,
		_w3722_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		\configuration_pci_ba0_bit31_8_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		_w3723_
	);
	LUT4 #(
		.INIT('hf531)
	) name712 (
		\configuration_pci_ba0_bit31_8_reg[20]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[28]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		_w3724_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name713 (
		\configuration_pci_ba0_bit31_8_reg[21]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		_w3725_
	);
	LUT4 #(
		.INIT('h8caf)
	) name714 (
		\configuration_pci_ba0_bit31_8_reg[15]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[28]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		_w3726_
	);
	LUT4 #(
		.INIT('h4000)
	) name715 (
		_w3723_,
		_w3725_,
		_w3726_,
		_w3724_,
		_w3727_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		_w3722_,
		_w3727_,
		_w3728_
	);
	LUT4 #(
		.INIT('h8caf)
	) name717 (
		\configuration_pci_ba0_bit31_8_reg[22]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w3729_
	);
	LUT4 #(
		.INIT('haf23)
	) name718 (
		\configuration_pci_ba0_bit31_8_reg[26]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[29]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		_w3730_
	);
	LUT4 #(
		.INIT('hf531)
	) name719 (
		\configuration_pci_ba0_bit31_8_reg[22]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		_w3731_
	);
	LUT4 #(
		.INIT('haf23)
	) name720 (
		\configuration_pci_ba0_bit31_8_reg[12]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		_w3732_
	);
	LUT4 #(
		.INIT('h8000)
	) name721 (
		_w3731_,
		_w3732_,
		_w3729_,
		_w3730_,
		_w3733_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name722 (
		\configuration_pci_ba0_bit31_8_reg[23]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[29]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		_w3734_
	);
	LUT4 #(
		.INIT('haf23)
	) name723 (
		\configuration_pci_ba0_bit31_8_reg[13]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w3735_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name724 (
		\configuration_pci_ba0_bit31_8_reg[15]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		_w3736_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name725 (
		\configuration_pci_ba0_bit31_8_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3737_
	);
	LUT4 #(
		.INIT('h8000)
	) name726 (
		_w3736_,
		_w3737_,
		_w3734_,
		_w3735_,
		_w3738_
	);
	LUT4 #(
		.INIT('h2000)
	) name727 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3739_
	);
	LUT4 #(
		.INIT('h8421)
	) name728 (
		\configuration_pci_ba0_bit31_8_reg[18]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		_w3740_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		_w3739_,
		_w3740_,
		_w3741_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name730 (
		\configuration_pci_ba0_bit31_8_reg[16]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		_w3742_
	);
	LUT4 #(
		.INIT('hf531)
	) name731 (
		\configuration_pci_ba0_bit31_8_reg[12]/NET0131 ,
		\configuration_pci_ba0_bit31_8_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		_w3743_
	);
	LUT2 #(
		.INIT('h6)
	) name732 (
		\configuration_pci_ba0_bit31_8_reg[17]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		_w3744_
	);
	LUT3 #(
		.INIT('h80)
	) name733 (
		\configuration_command_bit2_0_reg[1]/NET0131 ,
		\configuration_init_complete_reg/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3745_
	);
	LUT4 #(
		.INIT('h4000)
	) name734 (
		_w3744_,
		_w3745_,
		_w3742_,
		_w3743_,
		_w3746_
	);
	LUT4 #(
		.INIT('h8000)
	) name735 (
		_w3741_,
		_w3746_,
		_w3733_,
		_w3738_,
		_w3747_
	);
	LUT4 #(
		.INIT('h1000)
	) name736 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\input_register_pci_idsel_reg_out_reg/NET0131 ,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w3698_,
		_w3748_,
		_w3749_
	);
	LUT3 #(
		.INIT('h07)
	) name738 (
		_w3728_,
		_w3747_,
		_w3749_,
		_w3750_
	);
	LUT4 #(
		.INIT('h1311)
	) name739 (
		_w3216_,
		_w3681_,
		_w3717_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h4)
	) name740 (
		_w3679_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h9)
	) name741 (
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		_w3753_
	);
	LUT2 #(
		.INIT('h6)
	) name742 (
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3754_
	);
	LUT4 #(
		.INIT('h9669)
	) name743 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		_w3755_
	);
	LUT2 #(
		.INIT('h9)
	) name744 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		_w3756_
	);
	LUT4 #(
		.INIT('h6996)
	) name745 (
		_w3753_,
		_w3754_,
		_w3755_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h9)
	) name746 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		_w3758_
	);
	LUT3 #(
		.INIT('h27)
	) name747 (
		\output_backup_par_en_out_reg/NET0131 ,
		\output_backup_par_out_reg/NET0131 ,
		pci_par_i_pad,
		_w3759_
	);
	LUT2 #(
		.INIT('h9)
	) name748 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		_w3760_
	);
	LUT4 #(
		.INIT('h9669)
	) name749 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3761_
	);
	LUT4 #(
		.INIT('h6996)
	) name750 (
		_w3758_,
		_w3759_,
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h6)
	) name751 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		_w3763_
	);
	LUT2 #(
		.INIT('h6)
	) name752 (
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		_w3764_
	);
	LUT4 #(
		.INIT('h9669)
	) name753 (
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		_w3765_
	);
	LUT3 #(
		.INIT('h96)
	) name754 (
		_w3763_,
		_w3764_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h69)
	) name755 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		_w3767_
	);
	LUT2 #(
		.INIT('h9)
	) name756 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		_w3768_
	);
	LUT3 #(
		.INIT('h96)
	) name757 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		_w3769_
	);
	LUT2 #(
		.INIT('h9)
	) name758 (
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		_w3770_
	);
	LUT4 #(
		.INIT('h6996)
	) name759 (
		_w3767_,
		_w3768_,
		_w3769_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('h9669)
	) name760 (
		_w3757_,
		_w3762_,
		_w3766_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('h8acf)
	) name761 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\input_register_pci_trdy_reg_out_reg/NET0131 ,
		\output_backup_irdy_en_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		\output_backup_mas_ad_en_out_reg/NET0131 ,
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3774_
	);
	LUT2 #(
		.INIT('he)
	) name763 (
		\output_backup_mas_ad_en_out_reg/NET0131 ,
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3775_
	);
	LUT3 #(
		.INIT('h01)
	) name764 (
		\output_backup_mas_ad_en_out_reg/NET0131 ,
		\output_backup_par_en_out_reg/NET0131 ,
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3776_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w3773_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h7)
	) name766 (
		_w3772_,
		_w3777_,
		_w3778_
	);
	LUT3 #(
		.INIT('h80)
	) name767 (
		_w3035_,
		_w3772_,
		_w3777_,
		_w3779_
	);
	LUT4 #(
		.INIT('h1555)
	) name768 (
		\parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131 ,
		_w3035_,
		_w3772_,
		_w3777_,
		_w3780_
	);
	LUT4 #(
		.INIT('heaaa)
	) name769 (
		\parity_checker_perr_en_crit_gen_perr_en_reg_out_reg/NET0131 ,
		_w3035_,
		_w3772_,
		_w3777_,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name770 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3782_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name771 (
		\configuration_status_bit15_11_reg[15]/NET0131 ,
		_w3043_,
		_w3047_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		\output_backup_perr_out_reg/NET0131 ,
		\output_backup_serr_out_reg/NET0131 ,
		_w3784_
	);
	LUT2 #(
		.INIT('hb)
	) name773 (
		_w3783_,
		_w3784_,
		_w3785_
	);
	LUT4 #(
		.INIT('h0010)
	) name774 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name775 (
		\output_backup_trdy_en_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3787_
	);
	LUT3 #(
		.INIT('h07)
	) name776 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131 ,
		_w3786_,
		_w3787_,
		_w3788_
	);
	LUT3 #(
		.INIT('h27)
	) name777 (
		\output_backup_trdy_en_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		pci_trdy_i_pad,
		_w3789_
	);
	LUT3 #(
		.INIT('hd8)
	) name778 (
		\output_backup_trdy_en_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		pci_trdy_i_pad,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		_w3208_,
		_w3789_,
		_w3791_
	);
	LUT4 #(
		.INIT('h0004)
	) name780 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w3792_
	);
	LUT4 #(
		.INIT('h0002)
	) name781 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w3793_
	);
	LUT4 #(
		.INIT('hfffd)
	) name782 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		_w3795_
	);
	LUT3 #(
		.INIT('h08)
	) name784 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		pci_gnt_i_pad,
		_w3796_
	);
	LUT3 #(
		.INIT('hea)
	) name785 (
		_w3792_,
		_w3793_,
		_w3796_,
		_w3797_
	);
	LUT4 #(
		.INIT('h0111)
	) name786 (
		_w3212_,
		_w3792_,
		_w3793_,
		_w3796_,
		_w3798_
	);
	LUT3 #(
		.INIT('hb0)
	) name787 (
		_w3788_,
		_w3791_,
		_w3798_,
		_w3799_
	);
	LUT3 #(
		.INIT('h4f)
	) name788 (
		_w3788_,
		_w3791_,
		_w3798_,
		_w3800_
	);
	LUT3 #(
		.INIT('ha8)
	) name789 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3801_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3802_
	);
	LUT4 #(
		.INIT('h2000)
	) name791 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3803_
	);
	LUT4 #(
		.INIT('h0001)
	) name792 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3804_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name793 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		_w3042_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('h0008)
	) name794 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3806_
	);
	LUT4 #(
		.INIT('h0004)
	) name795 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3807_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name796 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		_w3806_,
		_w3807_,
		_w3808_
	);
	LUT4 #(
		.INIT('h0080)
	) name797 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		\configuration_wb_err_data_reg[31]/NET0131 ,
		_w3809_,
		_w3810_
	);
	LUT4 #(
		.INIT('haaa8)
	) name799 (
		_w3803_,
		_w3808_,
		_w3805_,
		_w3810_,
		_w3811_
	);
	LUT3 #(
		.INIT('h80)
	) name800 (
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3812_
	);
	LUT4 #(
		.INIT('h8000)
	) name801 (
		\configuration_icr_bit31_reg/NET0131 ,
		_w3041_,
		_w3802_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w3814_
	);
	LUT4 #(
		.INIT('h0040)
	) name803 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3815_
	);
	LUT3 #(
		.INIT('h80)
	) name804 (
		\configuration_wb_err_addr_reg[31]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3817_
	);
	LUT4 #(
		.INIT('h1000)
	) name806 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3818_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		_w3818_,
		_w3807_,
		_w3819_
	);
	LUT3 #(
		.INIT('h80)
	) name808 (
		\configuration_wb_ta1_reg[31]/NET0131 ,
		_w3818_,
		_w3807_,
		_w3820_
	);
	LUT3 #(
		.INIT('h01)
	) name809 (
		_w3813_,
		_w3816_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3822_
	);
	LUT3 #(
		.INIT('h02)
	) name811 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w3823_
	);
	LUT4 #(
		.INIT('h0200)
	) name812 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3824_
	);
	LUT3 #(
		.INIT('h80)
	) name813 (
		\configuration_pci_ta1_reg[31]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('h80)
	) name814 (
		\configuration_wb_err_cs_bit31_24_reg[31]/NET0131 ,
		_w3809_,
		_w3818_,
		_w3826_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w3825_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('h2000)
	) name816 (
		\configuration_status_bit15_11_reg[15]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w3828_
	);
	LUT4 #(
		.INIT('h0100)
	) name817 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3829_
	);
	LUT4 #(
		.INIT('h0001)
	) name818 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3830_
	);
	LUT4 #(
		.INIT('h0777)
	) name819 (
		_w3042_,
		_w3829_,
		_w3830_,
		_w3807_,
		_w3831_
	);
	LUT3 #(
		.INIT('h31)
	) name820 (
		\configuration_pci_ba0_bit31_8_reg[31]/NET0131 ,
		_w3828_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('h80)
	) name821 (
		_w3821_,
		_w3827_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		_w3824_,
		_w3807_,
		_w3834_
	);
	LUT3 #(
		.INIT('h80)
	) name823 (
		\configuration_pci_ba1_bit31_8_reg[31]/NET0131 ,
		_w3040_,
		_w3806_,
		_w3835_
	);
	LUT3 #(
		.INIT('ha8)
	) name824 (
		\configuration_pci_am1_reg[31]/NET0131 ,
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('h0040)
	) name825 (
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3837_
	);
	LUT4 #(
		.INIT('h8000)
	) name826 (
		\configuration_pci_err_data_reg[31]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3838_
	);
	LUT3 #(
		.INIT('h80)
	) name827 (
		\configuration_wb_ta2_reg[31]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3839_
	);
	LUT4 #(
		.INIT('he0a0)
	) name828 (
		_w3824_,
		_w3817_,
		_w3804_,
		_w3839_,
		_w3840_
	);
	LUT3 #(
		.INIT('h80)
	) name829 (
		_w3039_,
		_w3814_,
		_w3837_,
		_w3841_
	);
	LUT4 #(
		.INIT('h8000)
	) name830 (
		\configuration_pci_err_cs_bit31_24_reg[31]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w3842_
	);
	LUT4 #(
		.INIT('h8000)
	) name831 (
		\configuration_pci_err_addr_reg[31]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3843_
	);
	LUT4 #(
		.INIT('h0001)
	) name832 (
		_w3838_,
		_w3840_,
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		_w3836_,
		_w3844_,
		_w3845_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name834 (
		_w3801_,
		_w3811_,
		_w3833_,
		_w3845_,
		_w3846_
	);
	LUT3 #(
		.INIT('h40)
	) name835 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001 ,
		_w3018_,
		_w3019_,
		_w3847_
	);
	LUT4 #(
		.INIT('hc888)
	) name836 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3848_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3849_
	);
	LUT4 #(
		.INIT('hff53)
	) name838 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[31]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3850_
	);
	LUT4 #(
		.INIT('h1055)
	) name839 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3847_,
		_w3848_,
		_w3850_,
		_w3851_
	);
	LUT3 #(
		.INIT('h02)
	) name840 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3852_
	);
	LUT4 #(
		.INIT('hac00)
	) name841 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]/NET0131 ,
		_w3260_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w3851_,
		_w3853_,
		_w3854_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name843 (
		\output_backup_ad_out_reg[31]/NET0131 ,
		_w3799_,
		_w3846_,
		_w3854_,
		_w3855_
	);
	LUT3 #(
		.INIT('h40)
	) name844 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001 ,
		_w3018_,
		_w3019_,
		_w3856_
	);
	LUT4 #(
		.INIT('hc888)
	) name845 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3857_
	);
	LUT3 #(
		.INIT('h08)
	) name846 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3858_
	);
	LUT4 #(
		.INIT('h5551)
	) name847 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[16]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3859_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w3858_,
		_w3859_,
		_w3860_
	);
	LUT3 #(
		.INIT('hb0)
	) name849 (
		_w3856_,
		_w3857_,
		_w3860_,
		_w3861_
	);
	LUT4 #(
		.INIT('h5030)
	) name850 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3862_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		\configuration_pci_ba0_bit31_8_reg[16]/NET0131 ,
		_w3831_,
		_w3863_
	);
	LUT3 #(
		.INIT('h80)
	) name852 (
		\configuration_wb_err_data_reg[16]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3864_
	);
	LUT3 #(
		.INIT('h80)
	) name853 (
		\configuration_wb_err_addr_reg[16]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3865_
	);
	LUT4 #(
		.INIT('h8000)
	) name854 (
		\configuration_pci_err_data_reg[16]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3866_
	);
	LUT4 #(
		.INIT('h0008)
	) name855 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3867_
	);
	LUT4 #(
		.INIT('h153f)
	) name856 (
		_w3042_,
		_w3830_,
		_w3804_,
		_w3867_,
		_w3868_
	);
	LUT4 #(
		.INIT('h0100)
	) name857 (
		_w3864_,
		_w3866_,
		_w3865_,
		_w3868_,
		_w3869_
	);
	LUT3 #(
		.INIT('h80)
	) name858 (
		\configuration_pci_ba1_bit31_8_reg[16]/NET0131 ,
		_w3040_,
		_w3806_,
		_w3870_
	);
	LUT3 #(
		.INIT('ha8)
	) name859 (
		\configuration_pci_am1_reg[16]/NET0131 ,
		_w3834_,
		_w3870_,
		_w3871_
	);
	LUT3 #(
		.INIT('h80)
	) name860 (
		\configuration_pci_ta1_reg[16]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3872_
	);
	LUT4 #(
		.INIT('h8000)
	) name861 (
		\configuration_pci_err_addr_reg[16]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3873_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		_w3823_,
		_w3804_,
		_w3874_
	);
	LUT3 #(
		.INIT('h80)
	) name863 (
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3823_,
		_w3804_,
		_w3875_
	);
	LUT4 #(
		.INIT('h1333)
	) name864 (
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3044_,
		_w3823_,
		_w3804_,
		_w3876_
	);
	LUT3 #(
		.INIT('h04)
	) name865 (
		_w3873_,
		_w3876_,
		_w3872_,
		_w3877_
	);
	LUT4 #(
		.INIT('h1000)
	) name866 (
		_w3863_,
		_w3871_,
		_w3877_,
		_w3869_,
		_w3878_
	);
	LUT4 #(
		.INIT('h1113)
	) name867 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3861_,
		_w3862_,
		_w3878_,
		_w3879_
	);
	LUT3 #(
		.INIT('hb8)
	) name868 (
		\output_backup_ad_out_reg[16]/NET0131 ,
		_w3799_,
		_w3879_,
		_w3880_
	);
	LUT4 #(
		.INIT('h4500)
	) name869 (
		\output_backup_ad_out_reg[17]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w3881_
	);
	LUT3 #(
		.INIT('h40)
	) name870 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001 ,
		_w3018_,
		_w3019_,
		_w3882_
	);
	LUT4 #(
		.INIT('hc888)
	) name871 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3883_
	);
	LUT3 #(
		.INIT('h08)
	) name872 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3884_
	);
	LUT4 #(
		.INIT('h5551)
	) name873 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[17]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3885_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w3884_,
		_w3885_,
		_w3886_
	);
	LUT3 #(
		.INIT('hb0)
	) name875 (
		_w3882_,
		_w3883_,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('h5030)
	) name876 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3888_
	);
	LUT3 #(
		.INIT('h80)
	) name877 (
		\configuration_wb_err_data_reg[17]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3889_
	);
	LUT4 #(
		.INIT('h8000)
	) name878 (
		\configuration_pci_err_addr_reg[17]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3890_
	);
	LUT4 #(
		.INIT('h8000)
	) name879 (
		\configuration_pci_err_data_reg[17]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\configuration_pci_am1_reg[17]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[17]/NET0131 ,
		_w3892_
	);
	LUT3 #(
		.INIT('h80)
	) name881 (
		_w3040_,
		_w3806_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h0001)
	) name882 (
		_w3889_,
		_w3890_,
		_w3891_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('h2)
	) name883 (
		\configuration_pci_ba0_bit31_8_reg[17]/NET0131 ,
		_w3831_,
		_w3895_
	);
	LUT3 #(
		.INIT('h80)
	) name884 (
		\configuration_wb_err_addr_reg[17]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3896_
	);
	LUT3 #(
		.INIT('h80)
	) name885 (
		\configuration_pci_am1_reg[17]/NET0131 ,
		_w3824_,
		_w3807_,
		_w3897_
	);
	LUT3 #(
		.INIT('h80)
	) name886 (
		\configuration_pci_ta1_reg[17]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3898_
	);
	LUT4 #(
		.INIT('h0002)
	) name887 (
		_w3876_,
		_w3897_,
		_w3898_,
		_w3896_,
		_w3899_
	);
	LUT4 #(
		.INIT('h4555)
	) name888 (
		_w3888_,
		_w3895_,
		_w3894_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('h3032)
	) name889 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w3887_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w3881_,
		_w3901_,
		_w3902_
	);
	LUT4 #(
		.INIT('h4500)
	) name891 (
		\output_backup_ad_out_reg[18]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w3903_
	);
	LUT3 #(
		.INIT('h40)
	) name892 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001 ,
		_w3018_,
		_w3019_,
		_w3904_
	);
	LUT4 #(
		.INIT('hc888)
	) name893 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3905_
	);
	LUT3 #(
		.INIT('h08)
	) name894 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3906_
	);
	LUT4 #(
		.INIT('h5551)
	) name895 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT3 #(
		.INIT('hb0)
	) name897 (
		_w3904_,
		_w3905_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('h5030)
	) name898 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3910_
	);
	LUT3 #(
		.INIT('h80)
	) name899 (
		\configuration_wb_err_data_reg[18]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3911_
	);
	LUT4 #(
		.INIT('h8000)
	) name900 (
		\configuration_pci_err_addr_reg[18]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3912_
	);
	LUT4 #(
		.INIT('h8000)
	) name901 (
		\configuration_pci_err_data_reg[18]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3913_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		\configuration_pci_am1_reg[18]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[18]/NET0131 ,
		_w3914_
	);
	LUT3 #(
		.INIT('h80)
	) name903 (
		_w3040_,
		_w3806_,
		_w3914_,
		_w3915_
	);
	LUT4 #(
		.INIT('h0001)
	) name904 (
		_w3911_,
		_w3912_,
		_w3913_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\configuration_pci_ba0_bit31_8_reg[18]/NET0131 ,
		_w3831_,
		_w3917_
	);
	LUT3 #(
		.INIT('h80)
	) name906 (
		\configuration_wb_err_addr_reg[18]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3918_
	);
	LUT3 #(
		.INIT('h80)
	) name907 (
		\configuration_pci_am1_reg[18]/NET0131 ,
		_w3824_,
		_w3807_,
		_w3919_
	);
	LUT3 #(
		.INIT('h80)
	) name908 (
		\configuration_pci_ta1_reg[18]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3920_
	);
	LUT4 #(
		.INIT('h0002)
	) name909 (
		_w3876_,
		_w3919_,
		_w3920_,
		_w3918_,
		_w3921_
	);
	LUT4 #(
		.INIT('h4555)
	) name910 (
		_w3910_,
		_w3917_,
		_w3916_,
		_w3921_,
		_w3922_
	);
	LUT4 #(
		.INIT('h3032)
	) name911 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w3909_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w3903_,
		_w3923_,
		_w3924_
	);
	LUT3 #(
		.INIT('h40)
	) name913 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001 ,
		_w3018_,
		_w3019_,
		_w3925_
	);
	LUT4 #(
		.INIT('hc888)
	) name914 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3926_
	);
	LUT3 #(
		.INIT('h08)
	) name915 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3927_
	);
	LUT4 #(
		.INIT('h5551)
	) name916 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[19]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3928_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w3927_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('hb0)
	) name918 (
		_w3925_,
		_w3926_,
		_w3929_,
		_w3930_
	);
	LUT4 #(
		.INIT('h5030)
	) name919 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3931_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		\configuration_pci_ba0_bit31_8_reg[19]/NET0131 ,
		_w3831_,
		_w3932_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		_w3806_,
		_w3867_,
		_w3933_
	);
	LUT4 #(
		.INIT('h8000)
	) name922 (
		\configuration_pci_err_data_reg[19]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3934_
	);
	LUT3 #(
		.INIT('h80)
	) name923 (
		\configuration_wb_err_addr_reg[19]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3935_
	);
	LUT4 #(
		.INIT('h0002)
	) name924 (
		_w3876_,
		_w3933_,
		_w3934_,
		_w3935_,
		_w3936_
	);
	LUT3 #(
		.INIT('h80)
	) name925 (
		\configuration_pci_ba1_bit31_8_reg[19]/NET0131 ,
		_w3040_,
		_w3806_,
		_w3937_
	);
	LUT3 #(
		.INIT('ha8)
	) name926 (
		\configuration_pci_am1_reg[19]/NET0131 ,
		_w3834_,
		_w3937_,
		_w3938_
	);
	LUT3 #(
		.INIT('h80)
	) name927 (
		\configuration_pci_ta1_reg[19]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3939_
	);
	LUT4 #(
		.INIT('h8000)
	) name928 (
		\configuration_pci_err_addr_reg[19]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3940_
	);
	LUT3 #(
		.INIT('h80)
	) name929 (
		\configuration_wb_err_data_reg[19]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3941_
	);
	LUT3 #(
		.INIT('h01)
	) name930 (
		_w3940_,
		_w3941_,
		_w3939_,
		_w3942_
	);
	LUT4 #(
		.INIT('h1000)
	) name931 (
		_w3938_,
		_w3932_,
		_w3942_,
		_w3936_,
		_w3943_
	);
	LUT4 #(
		.INIT('h1113)
	) name932 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3930_,
		_w3931_,
		_w3943_,
		_w3944_
	);
	LUT3 #(
		.INIT('hb8)
	) name933 (
		\output_backup_ad_out_reg[19]/NET0131 ,
		_w3799_,
		_w3944_,
		_w3945_
	);
	LUT4 #(
		.INIT('h4500)
	) name934 (
		\output_backup_ad_out_reg[1]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w3946_
	);
	LUT4 #(
		.INIT('h5030)
	) name935 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3947_
	);
	LUT3 #(
		.INIT('h40)
	) name936 (
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w3948_
	);
	LUT4 #(
		.INIT('h2000)
	) name937 (
		\configuration_cache_line_size_reg_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w3949_
	);
	LUT4 #(
		.INIT('h2000)
	) name938 (
		\configuration_command_bit2_0_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w3950_
	);
	LUT3 #(
		.INIT('h80)
	) name939 (
		\configuration_wb_err_addr_reg[1]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3951_
	);
	LUT4 #(
		.INIT('h1333)
	) name940 (
		\configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131 ,
		_w3044_,
		_w3829_,
		_w3807_,
		_w3952_
	);
	LUT4 #(
		.INIT('h0100)
	) name941 (
		_w3950_,
		_w3951_,
		_w3949_,
		_w3952_,
		_w3953_
	);
	LUT3 #(
		.INIT('h80)
	) name942 (
		\configuration_wb_err_data_reg[1]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3954_
	);
	LUT3 #(
		.INIT('h08)
	) name943 (
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3955_
	);
	LUT4 #(
		.INIT('h0080)
	) name944 (
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w3956_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		_w3957_
	);
	LUT4 #(
		.INIT('h1000)
	) name946 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w3958_
	);
	LUT3 #(
		.INIT('h80)
	) name947 (
		\configuration_isr_bit2_0_reg[1]/NET0131 ,
		_w3956_,
		_w3958_,
		_w3959_
	);
	LUT4 #(
		.INIT('h8000)
	) name948 (
		\configuration_pci_err_data_reg[1]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3960_
	);
	LUT4 #(
		.INIT('h8000)
	) name949 (
		\configuration_icr_bit2_0_reg[1]/NET0131 ,
		_w3041_,
		_w3802_,
		_w3812_,
		_w3961_
	);
	LUT4 #(
		.INIT('h0001)
	) name950 (
		_w3954_,
		_w3959_,
		_w3960_,
		_w3961_,
		_w3962_
	);
	LUT3 #(
		.INIT('h80)
	) name951 (
		\configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131 ,
		_w3042_,
		_w3818_,
		_w3963_
	);
	LUT3 #(
		.INIT('h80)
	) name952 (
		\configuration_interrupt_line_reg[1]/NET0131 ,
		_w3806_,
		_w3867_,
		_w3964_
	);
	LUT4 #(
		.INIT('h8000)
	) name953 (
		\configuration_pci_err_addr_reg[1]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3965_
	);
	LUT3 #(
		.INIT('h80)
	) name954 (
		\configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131 ,
		_w3806_,
		_w3818_,
		_w3966_
	);
	LUT4 #(
		.INIT('h0001)
	) name955 (
		_w3963_,
		_w3964_,
		_w3965_,
		_w3966_,
		_w3967_
	);
	LUT4 #(
		.INIT('h1555)
	) name956 (
		_w3947_,
		_w3962_,
		_w3967_,
		_w3953_,
		_w3968_
	);
	LUT3 #(
		.INIT('h40)
	) name957 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001 ,
		_w3018_,
		_w3019_,
		_w3969_
	);
	LUT4 #(
		.INIT('hc888)
	) name958 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3970_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w3969_,
		_w3970_,
		_w3971_
	);
	LUT3 #(
		.INIT('h02)
	) name960 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131 ,
		_w3972_
	);
	LUT4 #(
		.INIT('h0888)
	) name961 (
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131 ,
		_w3973_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name962 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131 ,
		_w3974_
	);
	LUT4 #(
		.INIT('h0e02)
	) name963 (
		\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]/NET0131 ,
		_w3972_,
		_w3974_,
		_w3973_,
		_w3975_
	);
	LUT4 #(
		.INIT('h5551)
	) name964 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3976_
	);
	LUT3 #(
		.INIT('h70)
	) name965 (
		_w3849_,
		_w3975_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		_w3971_,
		_w3977_,
		_w3978_
	);
	LUT4 #(
		.INIT('h3302)
	) name967 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w3968_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w3946_,
		_w3979_,
		_w3980_
	);
	LUT4 #(
		.INIT('h4500)
	) name969 (
		\output_backup_ad_out_reg[20]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w3981_
	);
	LUT3 #(
		.INIT('h40)
	) name970 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001 ,
		_w3018_,
		_w3019_,
		_w3982_
	);
	LUT4 #(
		.INIT('hc888)
	) name971 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w3983_
	);
	LUT3 #(
		.INIT('h08)
	) name972 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3984_
	);
	LUT4 #(
		.INIT('h5551)
	) name973 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3985_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT3 #(
		.INIT('hb0)
	) name975 (
		_w3982_,
		_w3983_,
		_w3986_,
		_w3987_
	);
	LUT4 #(
		.INIT('h5030)
	) name976 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]/NET0131 ,
		_w3044_,
		_w3260_,
		_w3988_
	);
	LUT3 #(
		.INIT('h80)
	) name977 (
		\configuration_wb_err_data_reg[20]/NET0131 ,
		_w3809_,
		_w3803_,
		_w3989_
	);
	LUT4 #(
		.INIT('h8000)
	) name978 (
		\configuration_pci_err_addr_reg[20]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w3990_
	);
	LUT4 #(
		.INIT('h8000)
	) name979 (
		\configuration_pci_err_data_reg[20]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w3991_
	);
	LUT2 #(
		.INIT('h8)
	) name980 (
		\configuration_pci_am1_reg[20]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[20]/NET0131 ,
		_w3992_
	);
	LUT3 #(
		.INIT('h80)
	) name981 (
		_w3040_,
		_w3806_,
		_w3992_,
		_w3993_
	);
	LUT4 #(
		.INIT('h0001)
	) name982 (
		_w3989_,
		_w3990_,
		_w3991_,
		_w3993_,
		_w3994_
	);
	LUT2 #(
		.INIT('h2)
	) name983 (
		\configuration_pci_ba0_bit31_8_reg[20]/NET0131 ,
		_w3831_,
		_w3995_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		\configuration_wb_err_addr_reg[20]/NET0131 ,
		_w3803_,
		_w3815_,
		_w3996_
	);
	LUT3 #(
		.INIT('h80)
	) name985 (
		\configuration_pci_am1_reg[20]/NET0131 ,
		_w3824_,
		_w3807_,
		_w3997_
	);
	LUT3 #(
		.INIT('h80)
	) name986 (
		\configuration_pci_ta1_reg[20]/NET0131 ,
		_w3806_,
		_w3824_,
		_w3998_
	);
	LUT4 #(
		.INIT('h0002)
	) name987 (
		_w3876_,
		_w3997_,
		_w3998_,
		_w3996_,
		_w3999_
	);
	LUT4 #(
		.INIT('h4555)
	) name988 (
		_w3988_,
		_w3995_,
		_w3994_,
		_w3999_,
		_w4000_
	);
	LUT4 #(
		.INIT('h3032)
	) name989 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w3987_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w3981_,
		_w4001_,
		_w4002_
	);
	LUT4 #(
		.INIT('h4500)
	) name991 (
		\output_backup_ad_out_reg[21]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4003_
	);
	LUT3 #(
		.INIT('h40)
	) name992 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001 ,
		_w3018_,
		_w3019_,
		_w4004_
	);
	LUT4 #(
		.INIT('hc888)
	) name993 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4005_
	);
	LUT3 #(
		.INIT('h08)
	) name994 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4006_
	);
	LUT4 #(
		.INIT('h5551)
	) name995 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4007_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w4006_,
		_w4007_,
		_w4008_
	);
	LUT3 #(
		.INIT('hb0)
	) name997 (
		_w4004_,
		_w4005_,
		_w4008_,
		_w4009_
	);
	LUT3 #(
		.INIT('h80)
	) name998 (
		\configuration_pci_ba1_bit31_8_reg[21]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4010_
	);
	LUT3 #(
		.INIT('ha8)
	) name999 (
		\configuration_pci_am1_reg[21]/NET0131 ,
		_w3834_,
		_w4010_,
		_w4011_
	);
	LUT3 #(
		.INIT('h80)
	) name1000 (
		\configuration_wb_err_data_reg[21]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4012_
	);
	LUT4 #(
		.INIT('h8000)
	) name1001 (
		\configuration_pci_err_data_reg[21]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4013_
	);
	LUT3 #(
		.INIT('h80)
	) name1002 (
		\configuration_pci_ta1_reg[21]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4014_
	);
	LUT4 #(
		.INIT('h8000)
	) name1003 (
		\configuration_pci_err_addr_reg[21]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4015_
	);
	LUT4 #(
		.INIT('h0001)
	) name1004 (
		_w4012_,
		_w4013_,
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h80)
	) name1005 (
		\configuration_wb_err_addr_reg[21]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4017_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1006 (
		\configuration_pci_ba0_bit31_8_reg[21]/NET0131 ,
		_w3831_,
		_w3876_,
		_w4017_,
		_w4018_
	);
	LUT4 #(
		.INIT('h5030)
	) name1007 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4019_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1008 (
		_w4011_,
		_w4016_,
		_w4018_,
		_w4019_,
		_w4020_
	);
	LUT4 #(
		.INIT('h3032)
	) name1009 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w4009_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h1)
	) name1010 (
		_w4003_,
		_w4021_,
		_w4022_
	);
	LUT4 #(
		.INIT('h4500)
	) name1011 (
		\output_backup_ad_out_reg[22]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4023_
	);
	LUT3 #(
		.INIT('h40)
	) name1012 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001 ,
		_w3018_,
		_w3019_,
		_w4024_
	);
	LUT4 #(
		.INIT('hc888)
	) name1013 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4025_
	);
	LUT3 #(
		.INIT('h08)
	) name1014 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4026_
	);
	LUT4 #(
		.INIT('h5551)
	) name1015 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4027_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w4026_,
		_w4027_,
		_w4028_
	);
	LUT3 #(
		.INIT('hb0)
	) name1017 (
		_w4024_,
		_w4025_,
		_w4028_,
		_w4029_
	);
	LUT3 #(
		.INIT('h80)
	) name1018 (
		\configuration_pci_ba1_bit31_8_reg[22]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4030_
	);
	LUT3 #(
		.INIT('ha8)
	) name1019 (
		\configuration_pci_am1_reg[22]/NET0131 ,
		_w3834_,
		_w4030_,
		_w4031_
	);
	LUT3 #(
		.INIT('h80)
	) name1020 (
		\configuration_wb_err_data_reg[22]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4032_
	);
	LUT4 #(
		.INIT('h8000)
	) name1021 (
		\configuration_pci_err_data_reg[22]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4033_
	);
	LUT3 #(
		.INIT('h80)
	) name1022 (
		\configuration_pci_ta1_reg[22]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4034_
	);
	LUT4 #(
		.INIT('h8000)
	) name1023 (
		\configuration_pci_err_addr_reg[22]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4035_
	);
	LUT4 #(
		.INIT('h0001)
	) name1024 (
		_w4032_,
		_w4033_,
		_w4034_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h80)
	) name1025 (
		\configuration_wb_err_addr_reg[22]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4037_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1026 (
		\configuration_pci_ba0_bit31_8_reg[22]/NET0131 ,
		_w3831_,
		_w3876_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('h5030)
	) name1027 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4039_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1028 (
		_w4031_,
		_w4036_,
		_w4038_,
		_w4039_,
		_w4040_
	);
	LUT4 #(
		.INIT('h3032)
	) name1029 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w4029_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w4023_,
		_w4041_,
		_w4042_
	);
	LUT3 #(
		.INIT('h40)
	) name1031 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001 ,
		_w3018_,
		_w3019_,
		_w4043_
	);
	LUT4 #(
		.INIT('hc888)
	) name1032 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4044_
	);
	LUT3 #(
		.INIT('h08)
	) name1033 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4045_
	);
	LUT4 #(
		.INIT('h5551)
	) name1034 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4046_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w4045_,
		_w4046_,
		_w4047_
	);
	LUT3 #(
		.INIT('hb0)
	) name1036 (
		_w4043_,
		_w4044_,
		_w4047_,
		_w4048_
	);
	LUT4 #(
		.INIT('h5030)
	) name1037 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w3043_,
		_w3874_,
		_w4050_
	);
	LUT3 #(
		.INIT('h80)
	) name1039 (
		\configuration_wb_err_data_reg[23]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4051_
	);
	LUT4 #(
		.INIT('h1333)
	) name1040 (
		\configuration_wb_err_addr_reg[23]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4052_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1041 (
		\configuration_pci_ba0_bit31_8_reg[23]/NET0131 ,
		_w3831_,
		_w4051_,
		_w4052_,
		_w4053_
	);
	LUT3 #(
		.INIT('h80)
	) name1042 (
		\configuration_pci_ba1_bit31_8_reg[23]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4054_
	);
	LUT3 #(
		.INIT('ha8)
	) name1043 (
		\configuration_pci_am1_reg[23]/NET0131 ,
		_w3834_,
		_w4054_,
		_w4055_
	);
	LUT4 #(
		.INIT('h8000)
	) name1044 (
		\configuration_pci_err_addr_reg[23]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4056_
	);
	LUT3 #(
		.INIT('h80)
	) name1045 (
		\configuration_pci_ta1_reg[23]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4057_
	);
	LUT4 #(
		.INIT('h8000)
	) name1046 (
		\configuration_pci_err_data_reg[23]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4058_
	);
	LUT3 #(
		.INIT('h01)
	) name1047 (
		_w4057_,
		_w4058_,
		_w4056_,
		_w4059_
	);
	LUT4 #(
		.INIT('h2000)
	) name1048 (
		_w4050_,
		_w4055_,
		_w4059_,
		_w4053_,
		_w4060_
	);
	LUT4 #(
		.INIT('h1113)
	) name1049 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4048_,
		_w4049_,
		_w4060_,
		_w4061_
	);
	LUT3 #(
		.INIT('hb8)
	) name1050 (
		\output_backup_ad_out_reg[23]/NET0131 ,
		_w3799_,
		_w4061_,
		_w4062_
	);
	LUT3 #(
		.INIT('h40)
	) name1051 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001 ,
		_w3018_,
		_w3019_,
		_w4063_
	);
	LUT4 #(
		.INIT('hc888)
	) name1052 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4064_
	);
	LUT3 #(
		.INIT('h08)
	) name1053 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4065_
	);
	LUT4 #(
		.INIT('h5551)
	) name1054 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[24]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4066_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('hb0)
	) name1056 (
		_w4063_,
		_w4064_,
		_w4067_,
		_w4068_
	);
	LUT4 #(
		.INIT('h5030)
	) name1057 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4069_
	);
	LUT3 #(
		.INIT('h80)
	) name1058 (
		\configuration_wb_err_addr_reg[24]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4070_
	);
	LUT4 #(
		.INIT('h8000)
	) name1059 (
		\configuration_pci_err_addr_reg[24]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4071_
	);
	LUT4 #(
		.INIT('h8000)
	) name1060 (
		\configuration_pci_err_cs_bit31_24_reg[24]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4072_
	);
	LUT4 #(
		.INIT('h0002)
	) name1061 (
		_w3876_,
		_w4071_,
		_w4070_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('h2000)
	) name1062 (
		\configuration_status_bit8_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4074_
	);
	LUT3 #(
		.INIT('h0d)
	) name1063 (
		\configuration_pci_ba0_bit31_8_reg[24]/NET0131 ,
		_w3831_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h80)
	) name1064 (
		\configuration_pci_ba1_bit31_8_reg[24]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4076_
	);
	LUT3 #(
		.INIT('ha8)
	) name1065 (
		\configuration_pci_am1_reg[24]/NET0131 ,
		_w3834_,
		_w4076_,
		_w4077_
	);
	LUT4 #(
		.INIT('h8000)
	) name1066 (
		\configuration_pci_err_data_reg[24]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4078_
	);
	LUT3 #(
		.INIT('h80)
	) name1067 (
		\configuration_wb_err_data_reg[24]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4079_
	);
	LUT3 #(
		.INIT('h80)
	) name1068 (
		\configuration_wb_err_cs_bit31_24_reg[24]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4080_
	);
	LUT3 #(
		.INIT('h80)
	) name1069 (
		\configuration_pci_ta1_reg[24]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4081_
	);
	LUT4 #(
		.INIT('h0001)
	) name1070 (
		_w4078_,
		_w4079_,
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT4 #(
		.INIT('h4000)
	) name1071 (
		_w4077_,
		_w4082_,
		_w4073_,
		_w4075_,
		_w4083_
	);
	LUT4 #(
		.INIT('h1113)
	) name1072 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4068_,
		_w4069_,
		_w4083_,
		_w4084_
	);
	LUT3 #(
		.INIT('hb8)
	) name1073 (
		\output_backup_ad_out_reg[24]/NET0131 ,
		_w3799_,
		_w4084_,
		_w4085_
	);
	LUT3 #(
		.INIT('h40)
	) name1074 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001 ,
		_w3018_,
		_w3019_,
		_w4086_
	);
	LUT4 #(
		.INIT('hc888)
	) name1075 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4087_
	);
	LUT3 #(
		.INIT('h08)
	) name1076 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4088_
	);
	LUT4 #(
		.INIT('h5551)
	) name1077 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[27]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4089_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT3 #(
		.INIT('hb0)
	) name1079 (
		_w4086_,
		_w4087_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('h5030)
	) name1080 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4092_
	);
	LUT2 #(
		.INIT('h2)
	) name1081 (
		\configuration_pci_ba0_bit31_8_reg[27]/NET0131 ,
		_w3831_,
		_w4093_
	);
	LUT4 #(
		.INIT('h2000)
	) name1082 (
		\configuration_status_bit15_11_reg[11]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4094_
	);
	LUT3 #(
		.INIT('h02)
	) name1083 (
		_w3876_,
		_w3933_,
		_w4094_,
		_w4095_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w4093_,
		_w4095_,
		_w4096_
	);
	LUT3 #(
		.INIT('h80)
	) name1085 (
		\configuration_pci_ba1_bit31_8_reg[27]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4097_
	);
	LUT3 #(
		.INIT('ha8)
	) name1086 (
		\configuration_pci_am1_reg[27]/NET0131 ,
		_w3834_,
		_w4097_,
		_w4098_
	);
	LUT4 #(
		.INIT('h8000)
	) name1087 (
		\configuration_pci_err_cs_bit31_24_reg[27]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4099_
	);
	LUT3 #(
		.INIT('h80)
	) name1088 (
		\configuration_wb_err_data_reg[27]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4100_
	);
	LUT4 #(
		.INIT('h8000)
	) name1089 (
		\configuration_pci_err_addr_reg[27]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4101_
	);
	LUT3 #(
		.INIT('h01)
	) name1090 (
		_w4100_,
		_w4101_,
		_w4099_,
		_w4102_
	);
	LUT3 #(
		.INIT('h80)
	) name1091 (
		\configuration_pci_ta1_reg[27]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4103_
	);
	LUT3 #(
		.INIT('h80)
	) name1092 (
		\configuration_wb_err_addr_reg[27]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4104_
	);
	LUT4 #(
		.INIT('h8000)
	) name1093 (
		\configuration_pci_err_data_reg[27]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4105_
	);
	LUT3 #(
		.INIT('h80)
	) name1094 (
		\configuration_wb_err_cs_bit31_24_reg[27]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4106_
	);
	LUT4 #(
		.INIT('h0001)
	) name1095 (
		_w4103_,
		_w4105_,
		_w4104_,
		_w4106_,
		_w4107_
	);
	LUT3 #(
		.INIT('h40)
	) name1096 (
		_w4098_,
		_w4102_,
		_w4107_,
		_w4108_
	);
	LUT4 #(
		.INIT('ha888)
	) name1097 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4092_,
		_w4096_,
		_w4108_,
		_w4109_
	);
	LUT4 #(
		.INIT('h888b)
	) name1098 (
		\output_backup_ad_out_reg[27]/NET0131 ,
		_w3799_,
		_w4091_,
		_w4109_,
		_w4110_
	);
	LUT3 #(
		.INIT('h40)
	) name1099 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001 ,
		_w3018_,
		_w3019_,
		_w4111_
	);
	LUT4 #(
		.INIT('hc888)
	) name1100 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4112_
	);
	LUT3 #(
		.INIT('h08)
	) name1101 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4113_
	);
	LUT4 #(
		.INIT('h5551)
	) name1102 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[28]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4114_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT3 #(
		.INIT('hb0)
	) name1104 (
		_w4111_,
		_w4112_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h5030)
	) name1105 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4117_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		\configuration_pci_ba0_bit31_8_reg[28]/NET0131 ,
		_w3831_,
		_w4118_
	);
	LUT4 #(
		.INIT('h2000)
	) name1107 (
		\configuration_status_bit15_11_reg[12]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4119_
	);
	LUT3 #(
		.INIT('h02)
	) name1108 (
		_w3876_,
		_w3933_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h4)
	) name1109 (
		_w4118_,
		_w4120_,
		_w4121_
	);
	LUT3 #(
		.INIT('h80)
	) name1110 (
		\configuration_pci_ba1_bit31_8_reg[28]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4122_
	);
	LUT3 #(
		.INIT('ha8)
	) name1111 (
		\configuration_pci_am1_reg[28]/NET0131 ,
		_w3834_,
		_w4122_,
		_w4123_
	);
	LUT4 #(
		.INIT('h8000)
	) name1112 (
		\configuration_pci_err_addr_reg[28]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4124_
	);
	LUT3 #(
		.INIT('h80)
	) name1113 (
		\configuration_wb_err_data_reg[28]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4125_
	);
	LUT4 #(
		.INIT('h8000)
	) name1114 (
		\configuration_pci_err_data_reg[28]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4126_
	);
	LUT3 #(
		.INIT('h01)
	) name1115 (
		_w4125_,
		_w4126_,
		_w4124_,
		_w4127_
	);
	LUT4 #(
		.INIT('h8000)
	) name1116 (
		\configuration_pci_err_cs_bit31_24_reg[28]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4128_
	);
	LUT3 #(
		.INIT('h80)
	) name1117 (
		\configuration_wb_err_addr_reg[28]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4129_
	);
	LUT3 #(
		.INIT('h80)
	) name1118 (
		\configuration_pci_ta1_reg[28]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4130_
	);
	LUT3 #(
		.INIT('h80)
	) name1119 (
		\configuration_wb_err_cs_bit31_24_reg[28]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4131_
	);
	LUT4 #(
		.INIT('h0001)
	) name1120 (
		_w4128_,
		_w4130_,
		_w4129_,
		_w4131_,
		_w4132_
	);
	LUT3 #(
		.INIT('h40)
	) name1121 (
		_w4123_,
		_w4127_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('ha888)
	) name1122 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4117_,
		_w4121_,
		_w4133_,
		_w4134_
	);
	LUT4 #(
		.INIT('h888b)
	) name1123 (
		\output_backup_ad_out_reg[28]/NET0131 ,
		_w3799_,
		_w4116_,
		_w4134_,
		_w4135_
	);
	LUT3 #(
		.INIT('h40)
	) name1124 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001 ,
		_w3018_,
		_w3019_,
		_w4136_
	);
	LUT4 #(
		.INIT('hc888)
	) name1125 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4137_
	);
	LUT3 #(
		.INIT('h08)
	) name1126 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4138_
	);
	LUT4 #(
		.INIT('h5551)
	) name1127 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[29]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4139_
	);
	LUT2 #(
		.INIT('h4)
	) name1128 (
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT3 #(
		.INIT('hb0)
	) name1129 (
		_w4136_,
		_w4137_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('h5030)
	) name1130 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name1131 (
		\configuration_pci_ba0_bit31_8_reg[29]/NET0131 ,
		_w3831_,
		_w4143_
	);
	LUT3 #(
		.INIT('h80)
	) name1132 (
		\configuration_wb_err_addr_reg[29]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4144_
	);
	LUT4 #(
		.INIT('h8000)
	) name1133 (
		\configuration_pci_err_cs_bit31_24_reg[29]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4145_
	);
	LUT3 #(
		.INIT('h80)
	) name1134 (
		\configuration_pci_ta1_reg[29]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4146_
	);
	LUT4 #(
		.INIT('h0002)
	) name1135 (
		_w3876_,
		_w4145_,
		_w4146_,
		_w4144_,
		_w4147_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w4143_,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		\configuration_status_bit15_11_reg[13]/NET0131 ,
		_w3042_,
		_w4149_
	);
	LUT3 #(
		.INIT('h80)
	) name1138 (
		\configuration_pci_am1_reg[29]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[29]/NET0131 ,
		_w3806_,
		_w4150_
	);
	LUT3 #(
		.INIT('ha8)
	) name1139 (
		_w3830_,
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT3 #(
		.INIT('h80)
	) name1140 (
		\configuration_pci_ba1_bit31_8_reg[29]/NET0131 ,
		_w3806_,
		_w3829_,
		_w4152_
	);
	LUT3 #(
		.INIT('ha8)
	) name1141 (
		\configuration_pci_am1_reg[29]/NET0131 ,
		_w3834_,
		_w4152_,
		_w4153_
	);
	LUT4 #(
		.INIT('h8000)
	) name1142 (
		\configuration_pci_err_addr_reg[29]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4154_
	);
	LUT4 #(
		.INIT('h8000)
	) name1143 (
		\configuration_pci_err_data_reg[29]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4155_
	);
	LUT3 #(
		.INIT('h80)
	) name1144 (
		\configuration_wb_err_data_reg[29]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4156_
	);
	LUT3 #(
		.INIT('h80)
	) name1145 (
		\configuration_wb_err_cs_bit31_24_reg[29]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4157_
	);
	LUT4 #(
		.INIT('h0001)
	) name1146 (
		_w4154_,
		_w4155_,
		_w4156_,
		_w4157_,
		_w4158_
	);
	LUT3 #(
		.INIT('h10)
	) name1147 (
		_w4153_,
		_w4151_,
		_w4158_,
		_w4159_
	);
	LUT4 #(
		.INIT('ha888)
	) name1148 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4142_,
		_w4148_,
		_w4159_,
		_w4160_
	);
	LUT4 #(
		.INIT('h888b)
	) name1149 (
		\output_backup_ad_out_reg[29]/NET0131 ,
		_w3799_,
		_w4141_,
		_w4160_,
		_w4161_
	);
	LUT3 #(
		.INIT('h40)
	) name1150 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001 ,
		_w3018_,
		_w3019_,
		_w4162_
	);
	LUT4 #(
		.INIT('hc888)
	) name1151 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4163_
	);
	LUT3 #(
		.INIT('h08)
	) name1152 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4164_
	);
	LUT4 #(
		.INIT('h5551)
	) name1153 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4165_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		_w4164_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('hb0)
	) name1155 (
		_w4162_,
		_w4163_,
		_w4166_,
		_w4167_
	);
	LUT4 #(
		.INIT('h5030)
	) name1156 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4168_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		_w3044_,
		_w3868_,
		_w4169_
	);
	LUT3 #(
		.INIT('h80)
	) name1158 (
		\configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131 ,
		_w3806_,
		_w3818_,
		_w4170_
	);
	LUT3 #(
		.INIT('h80)
	) name1159 (
		\configuration_wb_err_addr_reg[2]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4171_
	);
	LUT3 #(
		.INIT('h80)
	) name1160 (
		\configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131 ,
		_w3829_,
		_w3807_,
		_w4172_
	);
	LUT3 #(
		.INIT('h01)
	) name1161 (
		_w4170_,
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('h2000)
	) name1162 (
		\configuration_command_bit2_0_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4174_
	);
	LUT4 #(
		.INIT('h2000)
	) name1163 (
		\configuration_cache_line_size_reg_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		_w4174_,
		_w4175_,
		_w4176_
	);
	LUT3 #(
		.INIT('h80)
	) name1165 (
		_w4169_,
		_w4173_,
		_w4176_,
		_w4177_
	);
	LUT3 #(
		.INIT('h80)
	) name1166 (
		\configuration_isr_bit2_0_reg[2]/NET0131 ,
		_w3956_,
		_w3958_,
		_w4178_
	);
	LUT4 #(
		.INIT('h8000)
	) name1167 (
		\configuration_pci_err_addr_reg[2]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4179_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		\configuration_interrupt_line_reg[2]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4180_
	);
	LUT3 #(
		.INIT('h01)
	) name1169 (
		_w4179_,
		_w4180_,
		_w4178_,
		_w4181_
	);
	LUT4 #(
		.INIT('h8000)
	) name1170 (
		\configuration_icr_bit2_0_reg[2]/NET0131 ,
		_w3041_,
		_w3802_,
		_w3812_,
		_w4182_
	);
	LUT3 #(
		.INIT('h80)
	) name1171 (
		\configuration_wb_err_data_reg[2]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4183_
	);
	LUT4 #(
		.INIT('h8000)
	) name1172 (
		\configuration_pci_err_data_reg[2]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4184_
	);
	LUT3 #(
		.INIT('h80)
	) name1173 (
		\configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131 ,
		_w3042_,
		_w3818_,
		_w4185_
	);
	LUT4 #(
		.INIT('h0001)
	) name1174 (
		_w4182_,
		_w4183_,
		_w4184_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w4181_,
		_w4186_,
		_w4187_
	);
	LUT4 #(
		.INIT('ha888)
	) name1176 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4168_,
		_w4177_,
		_w4187_,
		_w4188_
	);
	LUT4 #(
		.INIT('h888b)
	) name1177 (
		\output_backup_ad_out_reg[2]/NET0131 ,
		_w3799_,
		_w4167_,
		_w4188_,
		_w4189_
	);
	LUT3 #(
		.INIT('h40)
	) name1178 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001 ,
		_w3018_,
		_w3019_,
		_w4190_
	);
	LUT4 #(
		.INIT('hc888)
	) name1179 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4191_
	);
	LUT3 #(
		.INIT('h08)
	) name1180 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4192_
	);
	LUT4 #(
		.INIT('h5551)
	) name1181 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[30]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4193_
	);
	LUT2 #(
		.INIT('h4)
	) name1182 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT3 #(
		.INIT('hb0)
	) name1183 (
		_w4190_,
		_w4191_,
		_w4194_,
		_w4195_
	);
	LUT4 #(
		.INIT('h5030)
	) name1184 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4196_
	);
	LUT3 #(
		.INIT('h80)
	) name1185 (
		\configuration_wb_err_addr_reg[30]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4197_
	);
	LUT4 #(
		.INIT('h8000)
	) name1186 (
		\configuration_pci_err_cs_bit31_24_reg[30]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4198_
	);
	LUT3 #(
		.INIT('h80)
	) name1187 (
		\configuration_wb_err_data_reg[30]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4199_
	);
	LUT4 #(
		.INIT('h0002)
	) name1188 (
		_w3876_,
		_w4198_,
		_w4199_,
		_w4197_,
		_w4200_
	);
	LUT4 #(
		.INIT('h2000)
	) name1189 (
		\configuration_status_bit15_11_reg[14]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4201_
	);
	LUT3 #(
		.INIT('h0d)
	) name1190 (
		\configuration_pci_ba0_bit31_8_reg[30]/NET0131 ,
		_w3831_,
		_w4201_,
		_w4202_
	);
	LUT3 #(
		.INIT('h80)
	) name1191 (
		\configuration_pci_ba1_bit31_8_reg[30]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4203_
	);
	LUT3 #(
		.INIT('ha8)
	) name1192 (
		\configuration_pci_am1_reg[30]/NET0131 ,
		_w3834_,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('h8000)
	) name1193 (
		\configuration_pci_err_data_reg[30]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4205_
	);
	LUT4 #(
		.INIT('h8000)
	) name1194 (
		\configuration_pci_err_addr_reg[30]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4206_
	);
	LUT3 #(
		.INIT('h80)
	) name1195 (
		\configuration_wb_err_cs_bit31_24_reg[30]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4207_
	);
	LUT3 #(
		.INIT('h80)
	) name1196 (
		\configuration_pci_ta1_reg[30]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4208_
	);
	LUT4 #(
		.INIT('h0001)
	) name1197 (
		_w4205_,
		_w4206_,
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT4 #(
		.INIT('h4000)
	) name1198 (
		_w4204_,
		_w4209_,
		_w4200_,
		_w4202_,
		_w4210_
	);
	LUT4 #(
		.INIT('h1113)
	) name1199 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4195_,
		_w4196_,
		_w4210_,
		_w4211_
	);
	LUT3 #(
		.INIT('hb8)
	) name1200 (
		\output_backup_ad_out_reg[30]/NET0131 ,
		_w3799_,
		_w4211_,
		_w4212_
	);
	LUT3 #(
		.INIT('h40)
	) name1201 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001 ,
		_w3018_,
		_w3019_,
		_w4213_
	);
	LUT4 #(
		.INIT('hc888)
	) name1202 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4214_
	);
	LUT3 #(
		.INIT('h08)
	) name1203 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4215_
	);
	LUT4 #(
		.INIT('h5551)
	) name1204 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4216_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT3 #(
		.INIT('hb0)
	) name1206 (
		_w4213_,
		_w4214_,
		_w4217_,
		_w4218_
	);
	LUT4 #(
		.INIT('h5030)
	) name1207 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4219_
	);
	LUT4 #(
		.INIT('h8000)
	) name1208 (
		\configuration_pci_err_addr_reg[3]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4220_
	);
	LUT3 #(
		.INIT('h80)
	) name1209 (
		\configuration_wb_err_data_reg[3]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4221_
	);
	LUT4 #(
		.INIT('h8000)
	) name1210 (
		\configuration_pci_err_data_reg[3]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4222_
	);
	LUT3 #(
		.INIT('h01)
	) name1211 (
		_w4221_,
		_w4222_,
		_w4220_,
		_w4223_
	);
	LUT4 #(
		.INIT('h2000)
	) name1212 (
		\configuration_cache_line_size_reg_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4224_
	);
	LUT3 #(
		.INIT('h80)
	) name1213 (
		\configuration_interrupt_line_reg[3]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4225_
	);
	LUT4 #(
		.INIT('h1333)
	) name1214 (
		\configuration_wb_err_addr_reg[3]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4226_
	);
	LUT3 #(
		.INIT('h10)
	) name1215 (
		_w4225_,
		_w4224_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('ha888)
	) name1216 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4219_,
		_w4223_,
		_w4227_,
		_w4228_
	);
	LUT4 #(
		.INIT('h888b)
	) name1217 (
		\output_backup_ad_out_reg[3]/NET0131 ,
		_w3799_,
		_w4218_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h4500)
	) name1218 (
		\output_backup_ad_out_reg[4]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4230_
	);
	LUT4 #(
		.INIT('h8000)
	) name1219 (
		\configuration_pci_err_data_reg[4]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4231_
	);
	LUT3 #(
		.INIT('h80)
	) name1220 (
		\configuration_wb_err_data_reg[4]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4232_
	);
	LUT3 #(
		.INIT('h80)
	) name1221 (
		\configuration_interrupt_line_reg[4]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4233_
	);
	LUT3 #(
		.INIT('h01)
	) name1222 (
		_w4232_,
		_w4233_,
		_w4231_,
		_w4234_
	);
	LUT4 #(
		.INIT('h2000)
	) name1223 (
		\configuration_cache_line_size_reg_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4235_
	);
	LUT4 #(
		.INIT('h8000)
	) name1224 (
		\configuration_pci_err_addr_reg[4]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4236_
	);
	LUT3 #(
		.INIT('h80)
	) name1225 (
		\configuration_wb_err_addr_reg[4]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4237_
	);
	LUT4 #(
		.INIT('h0004)
	) name1226 (
		_w3044_,
		_w3868_,
		_w4236_,
		_w4237_,
		_w4238_
	);
	LUT4 #(
		.INIT('h5030)
	) name1227 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4239_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1228 (
		_w4235_,
		_w4234_,
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT3 #(
		.INIT('h40)
	) name1229 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001 ,
		_w3018_,
		_w3019_,
		_w4241_
	);
	LUT4 #(
		.INIT('hc888)
	) name1230 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4242_
	);
	LUT3 #(
		.INIT('h08)
	) name1231 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4243_
	);
	LUT4 #(
		.INIT('h5551)
	) name1232 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4244_
	);
	LUT2 #(
		.INIT('h4)
	) name1233 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT3 #(
		.INIT('hb0)
	) name1234 (
		_w4241_,
		_w4242_,
		_w4245_,
		_w4246_
	);
	LUT4 #(
		.INIT('h3302)
	) name1235 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w4240_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w4230_,
		_w4247_,
		_w4248_
	);
	LUT3 #(
		.INIT('h40)
	) name1237 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001 ,
		_w3018_,
		_w3019_,
		_w4249_
	);
	LUT4 #(
		.INIT('hc888)
	) name1238 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4250_
	);
	LUT3 #(
		.INIT('h08)
	) name1239 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4251_
	);
	LUT4 #(
		.INIT('h5551)
	) name1240 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4252_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		_w4251_,
		_w4252_,
		_w4253_
	);
	LUT3 #(
		.INIT('hb0)
	) name1242 (
		_w4249_,
		_w4250_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h5030)
	) name1243 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4255_
	);
	LUT4 #(
		.INIT('h8000)
	) name1244 (
		\configuration_pci_err_addr_reg[5]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4256_
	);
	LUT3 #(
		.INIT('h80)
	) name1245 (
		\configuration_wb_err_data_reg[5]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4257_
	);
	LUT4 #(
		.INIT('h8000)
	) name1246 (
		\configuration_pci_err_data_reg[5]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4258_
	);
	LUT3 #(
		.INIT('h01)
	) name1247 (
		_w4257_,
		_w4258_,
		_w4256_,
		_w4259_
	);
	LUT4 #(
		.INIT('h2000)
	) name1248 (
		\configuration_cache_line_size_reg_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4260_
	);
	LUT3 #(
		.INIT('h80)
	) name1249 (
		\configuration_interrupt_line_reg[5]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4261_
	);
	LUT4 #(
		.INIT('h1333)
	) name1250 (
		\configuration_wb_err_addr_reg[5]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4262_
	);
	LUT3 #(
		.INIT('h10)
	) name1251 (
		_w4261_,
		_w4260_,
		_w4262_,
		_w4263_
	);
	LUT4 #(
		.INIT('ha888)
	) name1252 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4255_,
		_w4259_,
		_w4263_,
		_w4264_
	);
	LUT4 #(
		.INIT('h888b)
	) name1253 (
		\output_backup_ad_out_reg[5]/NET0131 ,
		_w3799_,
		_w4254_,
		_w4264_,
		_w4265_
	);
	LUT3 #(
		.INIT('h40)
	) name1254 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001 ,
		_w3018_,
		_w3019_,
		_w4266_
	);
	LUT4 #(
		.INIT('hc888)
	) name1255 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4267_
	);
	LUT3 #(
		.INIT('h08)
	) name1256 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4268_
	);
	LUT4 #(
		.INIT('h5551)
	) name1257 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT3 #(
		.INIT('hb0)
	) name1259 (
		_w4266_,
		_w4267_,
		_w4270_,
		_w4271_
	);
	LUT4 #(
		.INIT('h5030)
	) name1260 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4272_
	);
	LUT3 #(
		.INIT('h80)
	) name1261 (
		\configuration_wb_err_data_reg[6]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4273_
	);
	LUT4 #(
		.INIT('h8000)
	) name1262 (
		\configuration_pci_err_data_reg[6]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4274_
	);
	LUT4 #(
		.INIT('h8000)
	) name1263 (
		\configuration_pci_err_addr_reg[6]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4275_
	);
	LUT3 #(
		.INIT('h01)
	) name1264 (
		_w4274_,
		_w4275_,
		_w4273_,
		_w4276_
	);
	LUT4 #(
		.INIT('h2000)
	) name1265 (
		\configuration_cache_line_size_reg_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4277_
	);
	LUT4 #(
		.INIT('h2000)
	) name1266 (
		\configuration_command_bit6_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4278_
	);
	LUT3 #(
		.INIT('h80)
	) name1267 (
		\configuration_interrupt_line_reg[6]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4279_
	);
	LUT4 #(
		.INIT('h1333)
	) name1268 (
		\configuration_wb_err_addr_reg[6]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4280_
	);
	LUT4 #(
		.INIT('h0100)
	) name1269 (
		_w4278_,
		_w4279_,
		_w4277_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('ha888)
	) name1270 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4272_,
		_w4276_,
		_w4281_,
		_w4282_
	);
	LUT4 #(
		.INIT('h888b)
	) name1271 (
		\output_backup_ad_out_reg[6]/NET0131 ,
		_w3799_,
		_w4271_,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('h4500)
	) name1272 (
		\output_backup_ad_out_reg[7]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4284_
	);
	LUT4 #(
		.INIT('h8000)
	) name1273 (
		\configuration_pci_err_data_reg[7]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4285_
	);
	LUT3 #(
		.INIT('h80)
	) name1274 (
		\configuration_wb_err_data_reg[7]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4286_
	);
	LUT3 #(
		.INIT('h80)
	) name1275 (
		\configuration_interrupt_line_reg[7]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4287_
	);
	LUT3 #(
		.INIT('h01)
	) name1276 (
		_w4286_,
		_w4287_,
		_w4285_,
		_w4288_
	);
	LUT4 #(
		.INIT('h2000)
	) name1277 (
		\configuration_cache_line_size_reg_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4289_
	);
	LUT4 #(
		.INIT('h8000)
	) name1278 (
		\configuration_pci_err_addr_reg[7]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4290_
	);
	LUT3 #(
		.INIT('h80)
	) name1279 (
		\configuration_wb_err_addr_reg[7]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4291_
	);
	LUT4 #(
		.INIT('h0004)
	) name1280 (
		_w3044_,
		_w3868_,
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT4 #(
		.INIT('h5030)
	) name1281 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4293_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1282 (
		_w4289_,
		_w4288_,
		_w4292_,
		_w4293_,
		_w4294_
	);
	LUT3 #(
		.INIT('h40)
	) name1283 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001 ,
		_w3018_,
		_w3019_,
		_w4295_
	);
	LUT4 #(
		.INIT('hc888)
	) name1284 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4296_
	);
	LUT3 #(
		.INIT('h08)
	) name1285 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4297_
	);
	LUT4 #(
		.INIT('h5551)
	) name1286 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[7]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4298_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT3 #(
		.INIT('hb0)
	) name1288 (
		_w4295_,
		_w4296_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('h3302)
	) name1289 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w4294_,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w4284_,
		_w4301_,
		_w4302_
	);
	LUT3 #(
		.INIT('h40)
	) name1291 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001 ,
		_w3018_,
		_w3019_,
		_w4303_
	);
	LUT4 #(
		.INIT('hc888)
	) name1292 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4304_
	);
	LUT3 #(
		.INIT('h08)
	) name1293 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4305_
	);
	LUT4 #(
		.INIT('h5551)
	) name1294 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4306_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT3 #(
		.INIT('hb0)
	) name1296 (
		_w4303_,
		_w4304_,
		_w4307_,
		_w4308_
	);
	LUT4 #(
		.INIT('h5030)
	) name1297 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4309_
	);
	LUT3 #(
		.INIT('h80)
	) name1298 (
		\configuration_wb_err_addr_reg[8]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4310_
	);
	LUT3 #(
		.INIT('h15)
	) name1299 (
		_w3044_,
		_w3806_,
		_w3867_,
		_w4311_
	);
	LUT3 #(
		.INIT('h80)
	) name1300 (
		\configuration_wb_err_cs_bit8_reg/NET0131 ,
		_w3809_,
		_w3818_,
		_w4312_
	);
	LUT3 #(
		.INIT('h80)
	) name1301 (
		\configuration_wb_err_data_reg[8]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4313_
	);
	LUT4 #(
		.INIT('h0100)
	) name1302 (
		_w4312_,
		_w4313_,
		_w4310_,
		_w4311_,
		_w4314_
	);
	LUT4 #(
		.INIT('h2000)
	) name1303 (
		\configuration_latency_timer_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4315_
	);
	LUT4 #(
		.INIT('h2000)
	) name1304 (
		\configuration_command_bit8_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4316_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w4315_,
		_w4316_,
		_w4317_
	);
	LUT3 #(
		.INIT('h80)
	) name1306 (
		\configuration_pci_ba1_bit31_8_reg[8]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4318_
	);
	LUT3 #(
		.INIT('ha8)
	) name1307 (
		\configuration_pci_am1_reg[8]/NET0131 ,
		_w3834_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h8000)
	) name1308 (
		\configuration_pci_err_addr_reg[8]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4320_
	);
	LUT4 #(
		.INIT('h8000)
	) name1309 (
		\configuration_pci_err_cs_bit8_reg/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4321_
	);
	LUT3 #(
		.INIT('h80)
	) name1310 (
		\configuration_pci_ta1_reg[8]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4322_
	);
	LUT4 #(
		.INIT('h8000)
	) name1311 (
		\configuration_pci_err_data_reg[8]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4323_
	);
	LUT4 #(
		.INIT('h0001)
	) name1312 (
		_w4320_,
		_w4321_,
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT4 #(
		.INIT('h4000)
	) name1313 (
		_w4319_,
		_w4324_,
		_w4314_,
		_w4317_,
		_w4325_
	);
	LUT4 #(
		.INIT('h1113)
	) name1314 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4308_,
		_w4309_,
		_w4325_,
		_w4326_
	);
	LUT3 #(
		.INIT('hb8)
	) name1315 (
		\output_backup_ad_out_reg[8]/NET0131 ,
		_w3799_,
		_w4326_,
		_w4327_
	);
	LUT3 #(
		.INIT('h40)
	) name1316 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001 ,
		_w3018_,
		_w3019_,
		_w4328_
	);
	LUT4 #(
		.INIT('hc888)
	) name1317 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4329_
	);
	LUT3 #(
		.INIT('h08)
	) name1318 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4330_
	);
	LUT4 #(
		.INIT('h5551)
	) name1319 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[9]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4331_
	);
	LUT2 #(
		.INIT('h4)
	) name1320 (
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT3 #(
		.INIT('hb0)
	) name1321 (
		_w4328_,
		_w4329_,
		_w4332_,
		_w4333_
	);
	LUT4 #(
		.INIT('h5030)
	) name1322 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4334_
	);
	LUT4 #(
		.INIT('h2000)
	) name1323 (
		\configuration_latency_timer_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4335_
	);
	LUT3 #(
		.INIT('h80)
	) name1324 (
		\configuration_pci_ta1_reg[9]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4336_
	);
	LUT4 #(
		.INIT('h1333)
	) name1325 (
		\configuration_wb_err_addr_reg[9]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4337_
	);
	LUT3 #(
		.INIT('h80)
	) name1326 (
		\configuration_wb_err_cs_bit9_reg/NET0131 ,
		_w3809_,
		_w3818_,
		_w4338_
	);
	LUT4 #(
		.INIT('h8000)
	) name1327 (
		\configuration_pci_err_data_reg[9]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4339_
	);
	LUT4 #(
		.INIT('h0100)
	) name1328 (
		_w4336_,
		_w4338_,
		_w4339_,
		_w4337_,
		_w4340_
	);
	LUT3 #(
		.INIT('h80)
	) name1329 (
		\configuration_pci_ba1_bit31_8_reg[9]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4341_
	);
	LUT3 #(
		.INIT('ha8)
	) name1330 (
		\configuration_pci_am1_reg[9]/NET0131 ,
		_w3834_,
		_w4341_,
		_w4342_
	);
	LUT3 #(
		.INIT('h80)
	) name1331 (
		\configuration_wb_err_data_reg[9]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4343_
	);
	LUT4 #(
		.INIT('h8000)
	) name1332 (
		\configuration_pci_err_addr_reg[9]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4344_
	);
	LUT4 #(
		.INIT('h8000)
	) name1333 (
		\configuration_pci_err_cs_bit10_reg/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4345_
	);
	LUT3 #(
		.INIT('h01)
	) name1334 (
		_w4344_,
		_w4345_,
		_w4343_,
		_w4346_
	);
	LUT4 #(
		.INIT('h1000)
	) name1335 (
		_w4342_,
		_w4335_,
		_w4346_,
		_w4340_,
		_w4347_
	);
	LUT4 #(
		.INIT('h1113)
	) name1336 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4333_,
		_w4334_,
		_w4347_,
		_w4348_
	);
	LUT3 #(
		.INIT('hb8)
	) name1337 (
		\output_backup_ad_out_reg[9]/NET0131 ,
		_w3799_,
		_w4348_,
		_w4349_
	);
	LUT4 #(
		.INIT('h4500)
	) name1338 (
		\output_backup_ad_out_reg[10]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4350_
	);
	LUT3 #(
		.INIT('h40)
	) name1339 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001 ,
		_w3018_,
		_w3019_,
		_w4351_
	);
	LUT4 #(
		.INIT('hc888)
	) name1340 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4352_
	);
	LUT3 #(
		.INIT('h08)
	) name1341 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4353_
	);
	LUT4 #(
		.INIT('h5551)
	) name1342 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4354_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT3 #(
		.INIT('hb0)
	) name1344 (
		_w4351_,
		_w4352_,
		_w4355_,
		_w4356_
	);
	LUT4 #(
		.INIT('h5030)
	) name1345 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4357_
	);
	LUT3 #(
		.INIT('h80)
	) name1346 (
		\configuration_pci_ba1_bit31_8_reg[10]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4358_
	);
	LUT3 #(
		.INIT('ha8)
	) name1347 (
		\configuration_pci_am1_reg[10]/NET0131 ,
		_w3834_,
		_w4358_,
		_w4359_
	);
	LUT3 #(
		.INIT('h80)
	) name1348 (
		\configuration_pci_ta1_reg[10]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4360_
	);
	LUT4 #(
		.INIT('h8000)
	) name1349 (
		\configuration_pci_err_addr_reg[10]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4361_
	);
	LUT4 #(
		.INIT('h8000)
	) name1350 (
		\configuration_pci_err_data_reg[10]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4362_
	);
	LUT3 #(
		.INIT('h80)
	) name1351 (
		\configuration_wb_err_data_reg[10]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4363_
	);
	LUT4 #(
		.INIT('h0001)
	) name1352 (
		_w4360_,
		_w4361_,
		_w4362_,
		_w4363_,
		_w4364_
	);
	LUT4 #(
		.INIT('h2000)
	) name1353 (
		\configuration_latency_timer_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4365_
	);
	LUT4 #(
		.INIT('h1333)
	) name1354 (
		\configuration_wb_err_addr_reg[10]/NET0131 ,
		_w3044_,
		_w3803_,
		_w3815_,
		_w4366_
	);
	LUT3 #(
		.INIT('h10)
	) name1355 (
		_w4345_,
		_w4365_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('h4555)
	) name1356 (
		_w4357_,
		_w4359_,
		_w4364_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h3032)
	) name1357 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3799_,
		_w4356_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w4350_,
		_w4369_,
		_w4370_
	);
	LUT3 #(
		.INIT('h40)
	) name1359 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001 ,
		_w3018_,
		_w3019_,
		_w4371_
	);
	LUT4 #(
		.INIT('hc888)
	) name1360 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4372_
	);
	LUT3 #(
		.INIT('h08)
	) name1361 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4373_
	);
	LUT4 #(
		.INIT('h5551)
	) name1362 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4374_
	);
	LUT2 #(
		.INIT('h4)
	) name1363 (
		_w4373_,
		_w4374_,
		_w4375_
	);
	LUT3 #(
		.INIT('hb0)
	) name1364 (
		_w4371_,
		_w4372_,
		_w4375_,
		_w4376_
	);
	LUT4 #(
		.INIT('h5030)
	) name1365 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4377_
	);
	LUT4 #(
		.INIT('h2000)
	) name1366 (
		\configuration_latency_timer_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4378_
	);
	LUT3 #(
		.INIT('h80)
	) name1367 (
		\configuration_pci_ta1_reg[11]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4379_
	);
	LUT3 #(
		.INIT('h80)
	) name1368 (
		\configuration_wb_err_addr_reg[11]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4380_
	);
	LUT4 #(
		.INIT('h0004)
	) name1369 (
		_w3044_,
		_w3868_,
		_w4379_,
		_w4380_,
		_w4381_
	);
	LUT3 #(
		.INIT('h80)
	) name1370 (
		\configuration_pci_ba1_bit31_8_reg[11]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4382_
	);
	LUT3 #(
		.INIT('ha8)
	) name1371 (
		\configuration_pci_am1_reg[11]/NET0131 ,
		_w3834_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('h8000)
	) name1372 (
		\configuration_pci_err_addr_reg[11]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4384_
	);
	LUT3 #(
		.INIT('h80)
	) name1373 (
		\configuration_wb_err_data_reg[11]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4385_
	);
	LUT4 #(
		.INIT('h8000)
	) name1374 (
		\configuration_pci_err_data_reg[11]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4386_
	);
	LUT3 #(
		.INIT('h01)
	) name1375 (
		_w4385_,
		_w4386_,
		_w4384_,
		_w4387_
	);
	LUT4 #(
		.INIT('h1000)
	) name1376 (
		_w4378_,
		_w4383_,
		_w4387_,
		_w4381_,
		_w4388_
	);
	LUT4 #(
		.INIT('h1113)
	) name1377 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4376_,
		_w4377_,
		_w4388_,
		_w4389_
	);
	LUT3 #(
		.INIT('hb8)
	) name1378 (
		\output_backup_ad_out_reg[11]/NET0131 ,
		_w3799_,
		_w4389_,
		_w4390_
	);
	LUT3 #(
		.INIT('h40)
	) name1379 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001 ,
		_w3018_,
		_w3019_,
		_w4391_
	);
	LUT4 #(
		.INIT('hc888)
	) name1380 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4392_
	);
	LUT3 #(
		.INIT('h08)
	) name1381 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4393_
	);
	LUT4 #(
		.INIT('h5551)
	) name1382 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[12]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4394_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		_w4393_,
		_w4394_,
		_w4395_
	);
	LUT3 #(
		.INIT('hb0)
	) name1384 (
		_w4391_,
		_w4392_,
		_w4395_,
		_w4396_
	);
	LUT4 #(
		.INIT('h5030)
	) name1385 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4397_
	);
	LUT4 #(
		.INIT('h2000)
	) name1386 (
		\configuration_latency_timer_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4398_
	);
	LUT4 #(
		.INIT('h3100)
	) name1387 (
		\configuration_pci_ba0_bit31_8_reg[12]/NET0131 ,
		_w3044_,
		_w3831_,
		_w3868_,
		_w4399_
	);
	LUT2 #(
		.INIT('h4)
	) name1388 (
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT3 #(
		.INIT('h80)
	) name1389 (
		\configuration_wb_err_data_reg[12]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4401_
	);
	LUT4 #(
		.INIT('h8000)
	) name1390 (
		\configuration_pci_err_addr_reg[12]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4402_
	);
	LUT4 #(
		.INIT('h8000)
	) name1391 (
		\configuration_pci_err_data_reg[12]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4403_
	);
	LUT3 #(
		.INIT('h01)
	) name1392 (
		_w4402_,
		_w4403_,
		_w4401_,
		_w4404_
	);
	LUT3 #(
		.INIT('h80)
	) name1393 (
		\configuration_pci_ta1_reg[12]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4405_
	);
	LUT3 #(
		.INIT('h80)
	) name1394 (
		\configuration_wb_err_addr_reg[12]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4406_
	);
	LUT3 #(
		.INIT('h01)
	) name1395 (
		_w3875_,
		_w4405_,
		_w4406_,
		_w4407_
	);
	LUT3 #(
		.INIT('h80)
	) name1396 (
		\configuration_pci_am1_reg[12]/NET0131 ,
		_w3824_,
		_w3807_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		\configuration_pci_am1_reg[12]/NET0131 ,
		\configuration_pci_ba1_bit31_8_reg[12]/NET0131 ,
		_w4409_
	);
	LUT3 #(
		.INIT('h80)
	) name1398 (
		_w3040_,
		_w3806_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w4408_,
		_w4410_,
		_w4411_
	);
	LUT3 #(
		.INIT('h80)
	) name1400 (
		_w4407_,
		_w4411_,
		_w4404_,
		_w4412_
	);
	LUT4 #(
		.INIT('ha888)
	) name1401 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4397_,
		_w4400_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('h888b)
	) name1402 (
		\output_backup_ad_out_reg[12]/NET0131 ,
		_w3799_,
		_w4396_,
		_w4413_,
		_w4414_
	);
	LUT3 #(
		.INIT('h40)
	) name1403 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001 ,
		_w3018_,
		_w3019_,
		_w4415_
	);
	LUT4 #(
		.INIT('hc888)
	) name1404 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4416_
	);
	LUT3 #(
		.INIT('h08)
	) name1405 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4417_
	);
	LUT4 #(
		.INIT('h5551)
	) name1406 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name1407 (
		_w4417_,
		_w4418_,
		_w4419_
	);
	LUT3 #(
		.INIT('hb0)
	) name1408 (
		_w4415_,
		_w4416_,
		_w4419_,
		_w4420_
	);
	LUT4 #(
		.INIT('h5030)
	) name1409 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4421_
	);
	LUT4 #(
		.INIT('h2000)
	) name1410 (
		\configuration_latency_timer_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4422_
	);
	LUT3 #(
		.INIT('h80)
	) name1411 (
		\configuration_wb_err_addr_reg[13]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4423_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1412 (
		\configuration_pci_ba0_bit31_8_reg[13]/NET0131 ,
		_w3831_,
		_w3876_,
		_w4423_,
		_w4424_
	);
	LUT3 #(
		.INIT('h80)
	) name1413 (
		\configuration_pci_ba1_bit31_8_reg[13]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4425_
	);
	LUT3 #(
		.INIT('ha8)
	) name1414 (
		\configuration_pci_am1_reg[13]/NET0131 ,
		_w3834_,
		_w4425_,
		_w4426_
	);
	LUT3 #(
		.INIT('h80)
	) name1415 (
		\configuration_pci_ta1_reg[13]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4427_
	);
	LUT3 #(
		.INIT('h80)
	) name1416 (
		\configuration_wb_err_data_reg[13]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4428_
	);
	LUT4 #(
		.INIT('h8000)
	) name1417 (
		\configuration_pci_err_addr_reg[13]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4429_
	);
	LUT4 #(
		.INIT('h8000)
	) name1418 (
		\configuration_pci_err_data_reg[13]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4430_
	);
	LUT4 #(
		.INIT('h0001)
	) name1419 (
		_w4427_,
		_w4428_,
		_w4429_,
		_w4430_,
		_w4431_
	);
	LUT4 #(
		.INIT('h1000)
	) name1420 (
		_w4426_,
		_w4422_,
		_w4431_,
		_w4424_,
		_w4432_
	);
	LUT4 #(
		.INIT('h1113)
	) name1421 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4420_,
		_w4421_,
		_w4432_,
		_w4433_
	);
	LUT3 #(
		.INIT('hb8)
	) name1422 (
		\output_backup_ad_out_reg[13]/NET0131 ,
		_w3799_,
		_w4433_,
		_w4434_
	);
	LUT3 #(
		.INIT('h40)
	) name1423 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001 ,
		_w3018_,
		_w3019_,
		_w4435_
	);
	LUT4 #(
		.INIT('hc888)
	) name1424 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4436_
	);
	LUT3 #(
		.INIT('h08)
	) name1425 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4437_
	);
	LUT4 #(
		.INIT('h5551)
	) name1426 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4438_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		_w4437_,
		_w4438_,
		_w4439_
	);
	LUT3 #(
		.INIT('hb0)
	) name1428 (
		_w4435_,
		_w4436_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h5030)
	) name1429 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4441_
	);
	LUT4 #(
		.INIT('h2000)
	) name1430 (
		\configuration_latency_timer_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4442_
	);
	LUT3 #(
		.INIT('h80)
	) name1431 (
		\configuration_wb_err_addr_reg[14]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4443_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1432 (
		\configuration_pci_ba0_bit31_8_reg[14]/NET0131 ,
		_w3831_,
		_w3876_,
		_w4443_,
		_w4444_
	);
	LUT3 #(
		.INIT('h80)
	) name1433 (
		\configuration_pci_ba1_bit31_8_reg[14]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4445_
	);
	LUT3 #(
		.INIT('ha8)
	) name1434 (
		\configuration_pci_am1_reg[14]/NET0131 ,
		_w3834_,
		_w4445_,
		_w4446_
	);
	LUT3 #(
		.INIT('h80)
	) name1435 (
		\configuration_pci_ta1_reg[14]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4447_
	);
	LUT4 #(
		.INIT('h8000)
	) name1436 (
		\configuration_pci_err_data_reg[14]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4448_
	);
	LUT4 #(
		.INIT('h8000)
	) name1437 (
		\configuration_pci_err_addr_reg[14]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4449_
	);
	LUT3 #(
		.INIT('h80)
	) name1438 (
		\configuration_wb_err_data_reg[14]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4450_
	);
	LUT4 #(
		.INIT('h0001)
	) name1439 (
		_w4447_,
		_w4448_,
		_w4449_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h1000)
	) name1440 (
		_w4446_,
		_w4442_,
		_w4451_,
		_w4444_,
		_w4452_
	);
	LUT4 #(
		.INIT('h1113)
	) name1441 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4440_,
		_w4441_,
		_w4452_,
		_w4453_
	);
	LUT3 #(
		.INIT('hb8)
	) name1442 (
		\output_backup_ad_out_reg[14]/NET0131 ,
		_w3799_,
		_w4453_,
		_w4454_
	);
	LUT3 #(
		.INIT('h40)
	) name1443 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001 ,
		_w3018_,
		_w3019_,
		_w4455_
	);
	LUT4 #(
		.INIT('hc888)
	) name1444 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4456_
	);
	LUT3 #(
		.INIT('h08)
	) name1445 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4457_
	);
	LUT4 #(
		.INIT('h5551)
	) name1446 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4458_
	);
	LUT2 #(
		.INIT('h4)
	) name1447 (
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('hb0)
	) name1448 (
		_w4455_,
		_w4456_,
		_w4459_,
		_w4460_
	);
	LUT4 #(
		.INIT('h5030)
	) name1449 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]/NET0131 ,
		_w3044_,
		_w3260_,
		_w4461_
	);
	LUT4 #(
		.INIT('h2000)
	) name1450 (
		\configuration_latency_timer_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4462_
	);
	LUT3 #(
		.INIT('h80)
	) name1451 (
		\configuration_wb_err_addr_reg[15]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4463_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1452 (
		\configuration_pci_ba0_bit31_8_reg[15]/NET0131 ,
		_w3831_,
		_w3876_,
		_w4463_,
		_w4464_
	);
	LUT3 #(
		.INIT('h80)
	) name1453 (
		\configuration_pci_ba1_bit31_8_reg[15]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4465_
	);
	LUT3 #(
		.INIT('ha8)
	) name1454 (
		\configuration_pci_am1_reg[15]/NET0131 ,
		_w3834_,
		_w4465_,
		_w4466_
	);
	LUT3 #(
		.INIT('h80)
	) name1455 (
		\configuration_pci_ta1_reg[15]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4467_
	);
	LUT4 #(
		.INIT('h8000)
	) name1456 (
		\configuration_pci_err_data_reg[15]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4468_
	);
	LUT3 #(
		.INIT('h80)
	) name1457 (
		\configuration_wb_err_data_reg[15]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4469_
	);
	LUT4 #(
		.INIT('h8000)
	) name1458 (
		\configuration_pci_err_addr_reg[15]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4470_
	);
	LUT4 #(
		.INIT('h0001)
	) name1459 (
		_w4467_,
		_w4468_,
		_w4469_,
		_w4470_,
		_w4471_
	);
	LUT4 #(
		.INIT('h1000)
	) name1460 (
		_w4466_,
		_w4462_,
		_w4471_,
		_w4464_,
		_w4472_
	);
	LUT4 #(
		.INIT('h1113)
	) name1461 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w4460_,
		_w4461_,
		_w4472_,
		_w4473_
	);
	LUT3 #(
		.INIT('hb8)
	) name1462 (
		\output_backup_ad_out_reg[15]/NET0131 ,
		_w3799_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w4475_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1464 (
		\configuration_status_bit15_11_reg[14]/NET0131 ,
		_w3043_,
		_w3047_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('he)
	) name1465 (
		\output_backup_serr_en_out_reg/NET0131 ,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h1055)
	) name1466 (
		_w3066_,
		_w3112_,
		_w3115_,
		_w3117_,
		_w4478_
	);
	LUT3 #(
		.INIT('h53)
	) name1467 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w4478_,
		_w4479_
	);
	LUT3 #(
		.INIT('hac)
	) name1468 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131 ,
		_w4478_,
		_w4480_
	);
	LUT3 #(
		.INIT('h53)
	) name1469 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w4478_,
		_w4481_
	);
	LUT4 #(
		.INIT('h0002)
	) name1470 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('h0008)
	) name1471 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4483_
	);
	LUT4 #(
		.INIT('h2000)
	) name1472 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4484_
	);
	LUT4 #(
		.INIT('h8000)
	) name1473 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4485_
	);
	LUT4 #(
		.INIT('h0001)
	) name1474 (
		_w4482_,
		_w4483_,
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT4 #(
		.INIT('h0200)
	) name1475 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4487_
	);
	LUT4 #(
		.INIT('h0800)
	) name1476 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4488_
	);
	LUT4 #(
		.INIT('h0080)
	) name1477 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4489_
	);
	LUT4 #(
		.INIT('h0020)
	) name1478 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4490_
	);
	LUT4 #(
		.INIT('h0001)
	) name1479 (
		_w4487_,
		_w4488_,
		_w4489_,
		_w4490_,
		_w4491_
	);
	LUT2 #(
		.INIT('h7)
	) name1480 (
		_w4486_,
		_w4491_,
		_w4492_
	);
	LUT4 #(
		.INIT('h0200)
	) name1481 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4493_
	);
	LUT4 #(
		.INIT('h0800)
	) name1482 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4494_
	);
	LUT4 #(
		.INIT('h0080)
	) name1483 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4495_
	);
	LUT4 #(
		.INIT('h0020)
	) name1484 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4496_
	);
	LUT4 #(
		.INIT('h0001)
	) name1485 (
		_w4493_,
		_w4494_,
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT4 #(
		.INIT('h2000)
	) name1486 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4498_
	);
	LUT4 #(
		.INIT('h8000)
	) name1487 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4499_
	);
	LUT4 #(
		.INIT('h0002)
	) name1488 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4500_
	);
	LUT4 #(
		.INIT('h0008)
	) name1489 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4501_
	);
	LUT4 #(
		.INIT('h0001)
	) name1490 (
		_w4498_,
		_w4499_,
		_w4500_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h7)
	) name1491 (
		_w4497_,
		_w4502_,
		_w4503_
	);
	LUT4 #(
		.INIT('h0200)
	) name1492 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4504_
	);
	LUT4 #(
		.INIT('h0800)
	) name1493 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4505_
	);
	LUT4 #(
		.INIT('h0002)
	) name1494 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4506_
	);
	LUT4 #(
		.INIT('h0008)
	) name1495 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4507_
	);
	LUT4 #(
		.INIT('h0001)
	) name1496 (
		_w4504_,
		_w4505_,
		_w4506_,
		_w4507_,
		_w4508_
	);
	LUT4 #(
		.INIT('h2000)
	) name1497 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4509_
	);
	LUT4 #(
		.INIT('h8000)
	) name1498 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4510_
	);
	LUT4 #(
		.INIT('h0080)
	) name1499 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4511_
	);
	LUT4 #(
		.INIT('h0020)
	) name1500 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4512_
	);
	LUT4 #(
		.INIT('h0001)
	) name1501 (
		_w4509_,
		_w4510_,
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h7)
	) name1502 (
		_w4508_,
		_w4513_,
		_w4514_
	);
	LUT4 #(
		.INIT('h0080)
	) name1503 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4515_
	);
	LUT4 #(
		.INIT('h0020)
	) name1504 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4516_
	);
	LUT4 #(
		.INIT('h2000)
	) name1505 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4517_
	);
	LUT4 #(
		.INIT('h8000)
	) name1506 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4518_
	);
	LUT4 #(
		.INIT('h0001)
	) name1507 (
		_w4515_,
		_w4516_,
		_w4517_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('h0800)
	) name1508 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4520_
	);
	LUT4 #(
		.INIT('h0200)
	) name1509 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4521_
	);
	LUT4 #(
		.INIT('h0008)
	) name1510 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4522_
	);
	LUT4 #(
		.INIT('h0002)
	) name1511 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4523_
	);
	LUT4 #(
		.INIT('h0001)
	) name1512 (
		_w4520_,
		_w4521_,
		_w4522_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h7)
	) name1513 (
		_w4519_,
		_w4524_,
		_w4525_
	);
	LUT4 #(
		.INIT('h0080)
	) name1514 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4526_
	);
	LUT4 #(
		.INIT('h0020)
	) name1515 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4527_
	);
	LUT4 #(
		.INIT('h2000)
	) name1516 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4528_
	);
	LUT4 #(
		.INIT('h8000)
	) name1517 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4529_
	);
	LUT4 #(
		.INIT('h0001)
	) name1518 (
		_w4526_,
		_w4527_,
		_w4528_,
		_w4529_,
		_w4530_
	);
	LUT4 #(
		.INIT('h0800)
	) name1519 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4531_
	);
	LUT4 #(
		.INIT('h0200)
	) name1520 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4532_
	);
	LUT4 #(
		.INIT('h0002)
	) name1521 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4533_
	);
	LUT4 #(
		.INIT('h0008)
	) name1522 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4534_
	);
	LUT4 #(
		.INIT('h0001)
	) name1523 (
		_w4531_,
		_w4532_,
		_w4533_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h7)
	) name1524 (
		_w4530_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h0080)
	) name1525 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4537_
	);
	LUT4 #(
		.INIT('h0020)
	) name1526 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4538_
	);
	LUT4 #(
		.INIT('h0200)
	) name1527 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4539_
	);
	LUT4 #(
		.INIT('h0800)
	) name1528 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4540_
	);
	LUT4 #(
		.INIT('h0001)
	) name1529 (
		_w4537_,
		_w4538_,
		_w4539_,
		_w4540_,
		_w4541_
	);
	LUT4 #(
		.INIT('h2000)
	) name1530 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4542_
	);
	LUT4 #(
		.INIT('h8000)
	) name1531 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4543_
	);
	LUT4 #(
		.INIT('h0002)
	) name1532 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4544_
	);
	LUT4 #(
		.INIT('h0008)
	) name1533 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4545_
	);
	LUT4 #(
		.INIT('h0001)
	) name1534 (
		_w4542_,
		_w4543_,
		_w4544_,
		_w4545_,
		_w4546_
	);
	LUT2 #(
		.INIT('h7)
	) name1535 (
		_w4541_,
		_w4546_,
		_w4547_
	);
	LUT4 #(
		.INIT('h0080)
	) name1536 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4548_
	);
	LUT4 #(
		.INIT('h0020)
	) name1537 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4549_
	);
	LUT4 #(
		.INIT('h2000)
	) name1538 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4550_
	);
	LUT4 #(
		.INIT('h8000)
	) name1539 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4551_
	);
	LUT4 #(
		.INIT('h0001)
	) name1540 (
		_w4548_,
		_w4549_,
		_w4550_,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('h0800)
	) name1541 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4553_
	);
	LUT4 #(
		.INIT('h0200)
	) name1542 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4554_
	);
	LUT4 #(
		.INIT('h0008)
	) name1543 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4555_
	);
	LUT4 #(
		.INIT('h0002)
	) name1544 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4556_
	);
	LUT4 #(
		.INIT('h0001)
	) name1545 (
		_w4553_,
		_w4554_,
		_w4555_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h7)
	) name1546 (
		_w4552_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('h0002)
	) name1547 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4559_
	);
	LUT4 #(
		.INIT('h0008)
	) name1548 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4560_
	);
	LUT4 #(
		.INIT('h2000)
	) name1549 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4561_
	);
	LUT4 #(
		.INIT('h8000)
	) name1550 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4562_
	);
	LUT4 #(
		.INIT('h0001)
	) name1551 (
		_w4559_,
		_w4560_,
		_w4561_,
		_w4562_,
		_w4563_
	);
	LUT4 #(
		.INIT('h0200)
	) name1552 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4564_
	);
	LUT4 #(
		.INIT('h0800)
	) name1553 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4565_
	);
	LUT4 #(
		.INIT('h0020)
	) name1554 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4566_
	);
	LUT4 #(
		.INIT('h0080)
	) name1555 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4567_
	);
	LUT4 #(
		.INIT('h0001)
	) name1556 (
		_w4564_,
		_w4565_,
		_w4566_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h7)
	) name1557 (
		_w4563_,
		_w4568_,
		_w4569_
	);
	LUT4 #(
		.INIT('h0200)
	) name1558 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4570_
	);
	LUT4 #(
		.INIT('h0800)
	) name1559 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4571_
	);
	LUT4 #(
		.INIT('h0002)
	) name1560 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4572_
	);
	LUT4 #(
		.INIT('h0008)
	) name1561 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4573_
	);
	LUT4 #(
		.INIT('h0001)
	) name1562 (
		_w4570_,
		_w4571_,
		_w4572_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('h2000)
	) name1563 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4575_
	);
	LUT4 #(
		.INIT('h8000)
	) name1564 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4576_
	);
	LUT4 #(
		.INIT('h0080)
	) name1565 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4577_
	);
	LUT4 #(
		.INIT('h0020)
	) name1566 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4578_
	);
	LUT4 #(
		.INIT('h0001)
	) name1567 (
		_w4575_,
		_w4576_,
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h7)
	) name1568 (
		_w4574_,
		_w4579_,
		_w4580_
	);
	LUT4 #(
		.INIT('h0080)
	) name1569 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4581_
	);
	LUT4 #(
		.INIT('h0020)
	) name1570 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4582_
	);
	LUT4 #(
		.INIT('h2000)
	) name1571 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4583_
	);
	LUT4 #(
		.INIT('h8000)
	) name1572 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4584_
	);
	LUT4 #(
		.INIT('h0001)
	) name1573 (
		_w4581_,
		_w4582_,
		_w4583_,
		_w4584_,
		_w4585_
	);
	LUT4 #(
		.INIT('h0800)
	) name1574 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4586_
	);
	LUT4 #(
		.INIT('h0200)
	) name1575 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4587_
	);
	LUT4 #(
		.INIT('h0002)
	) name1576 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4588_
	);
	LUT4 #(
		.INIT('h0008)
	) name1577 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4589_
	);
	LUT4 #(
		.INIT('h0001)
	) name1578 (
		_w4586_,
		_w4587_,
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT2 #(
		.INIT('h7)
	) name1579 (
		_w4585_,
		_w4590_,
		_w4591_
	);
	LUT4 #(
		.INIT('h0080)
	) name1580 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4592_
	);
	LUT4 #(
		.INIT('h0020)
	) name1581 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4593_
	);
	LUT4 #(
		.INIT('h0002)
	) name1582 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4594_
	);
	LUT4 #(
		.INIT('h0008)
	) name1583 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4595_
	);
	LUT4 #(
		.INIT('h0001)
	) name1584 (
		_w4592_,
		_w4593_,
		_w4594_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h0800)
	) name1585 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4597_
	);
	LUT4 #(
		.INIT('h0200)
	) name1586 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4598_
	);
	LUT4 #(
		.INIT('h2000)
	) name1587 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4599_
	);
	LUT4 #(
		.INIT('h8000)
	) name1588 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4600_
	);
	LUT4 #(
		.INIT('h0001)
	) name1589 (
		_w4597_,
		_w4598_,
		_w4599_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h7)
	) name1590 (
		_w4596_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('h0080)
	) name1591 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4603_
	);
	LUT4 #(
		.INIT('h0020)
	) name1592 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4604_
	);
	LUT4 #(
		.INIT('h2000)
	) name1593 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4605_
	);
	LUT4 #(
		.INIT('h8000)
	) name1594 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4606_
	);
	LUT4 #(
		.INIT('h0001)
	) name1595 (
		_w4603_,
		_w4604_,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT4 #(
		.INIT('h0002)
	) name1596 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4608_
	);
	LUT4 #(
		.INIT('h0008)
	) name1597 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4609_
	);
	LUT4 #(
		.INIT('h0200)
	) name1598 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4610_
	);
	LUT4 #(
		.INIT('h0800)
	) name1599 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4611_
	);
	LUT4 #(
		.INIT('h0001)
	) name1600 (
		_w4608_,
		_w4609_,
		_w4610_,
		_w4611_,
		_w4612_
	);
	LUT2 #(
		.INIT('h7)
	) name1601 (
		_w4607_,
		_w4612_,
		_w4613_
	);
	LUT4 #(
		.INIT('h0080)
	) name1602 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4614_
	);
	LUT4 #(
		.INIT('h0020)
	) name1603 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4615_
	);
	LUT4 #(
		.INIT('h0200)
	) name1604 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4616_
	);
	LUT4 #(
		.INIT('h0800)
	) name1605 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4617_
	);
	LUT4 #(
		.INIT('h0001)
	) name1606 (
		_w4614_,
		_w4615_,
		_w4616_,
		_w4617_,
		_w4618_
	);
	LUT4 #(
		.INIT('h0002)
	) name1607 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4619_
	);
	LUT4 #(
		.INIT('h0008)
	) name1608 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4620_
	);
	LUT4 #(
		.INIT('h2000)
	) name1609 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4621_
	);
	LUT4 #(
		.INIT('h8000)
	) name1610 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4622_
	);
	LUT4 #(
		.INIT('h0001)
	) name1611 (
		_w4619_,
		_w4620_,
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h7)
	) name1612 (
		_w4618_,
		_w4623_,
		_w4624_
	);
	LUT4 #(
		.INIT('h0080)
	) name1613 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4625_
	);
	LUT4 #(
		.INIT('h0020)
	) name1614 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4626_
	);
	LUT4 #(
		.INIT('h0200)
	) name1615 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4627_
	);
	LUT4 #(
		.INIT('h0800)
	) name1616 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4628_
	);
	LUT4 #(
		.INIT('h0001)
	) name1617 (
		_w4625_,
		_w4626_,
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT4 #(
		.INIT('h2000)
	) name1618 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4630_
	);
	LUT4 #(
		.INIT('h8000)
	) name1619 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4631_
	);
	LUT4 #(
		.INIT('h0008)
	) name1620 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4632_
	);
	LUT4 #(
		.INIT('h0002)
	) name1621 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4633_
	);
	LUT4 #(
		.INIT('h0001)
	) name1622 (
		_w4630_,
		_w4631_,
		_w4632_,
		_w4633_,
		_w4634_
	);
	LUT2 #(
		.INIT('h7)
	) name1623 (
		_w4629_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('h0200)
	) name1624 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4636_
	);
	LUT4 #(
		.INIT('h0800)
	) name1625 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4637_
	);
	LUT4 #(
		.INIT('h0002)
	) name1626 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4638_
	);
	LUT4 #(
		.INIT('h0008)
	) name1627 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4639_
	);
	LUT4 #(
		.INIT('h0001)
	) name1628 (
		_w4636_,
		_w4637_,
		_w4638_,
		_w4639_,
		_w4640_
	);
	LUT4 #(
		.INIT('h0080)
	) name1629 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4641_
	);
	LUT4 #(
		.INIT('h0020)
	) name1630 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4642_
	);
	LUT4 #(
		.INIT('h2000)
	) name1631 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4643_
	);
	LUT4 #(
		.INIT('h8000)
	) name1632 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4644_
	);
	LUT4 #(
		.INIT('h0001)
	) name1633 (
		_w4641_,
		_w4642_,
		_w4643_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h7)
	) name1634 (
		_w4640_,
		_w4645_,
		_w4646_
	);
	LUT4 #(
		.INIT('h0200)
	) name1635 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4647_
	);
	LUT4 #(
		.INIT('h0800)
	) name1636 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4648_
	);
	LUT4 #(
		.INIT('h0002)
	) name1637 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4649_
	);
	LUT4 #(
		.INIT('h0008)
	) name1638 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4650_
	);
	LUT4 #(
		.INIT('h0001)
	) name1639 (
		_w4647_,
		_w4648_,
		_w4649_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('h2000)
	) name1640 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4652_
	);
	LUT4 #(
		.INIT('h8000)
	) name1641 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4653_
	);
	LUT4 #(
		.INIT('h0080)
	) name1642 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4654_
	);
	LUT4 #(
		.INIT('h0020)
	) name1643 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4655_
	);
	LUT4 #(
		.INIT('h0001)
	) name1644 (
		_w4652_,
		_w4653_,
		_w4654_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h7)
	) name1645 (
		_w4651_,
		_w4656_,
		_w4657_
	);
	LUT4 #(
		.INIT('h0002)
	) name1646 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4658_
	);
	LUT4 #(
		.INIT('h0008)
	) name1647 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4659_
	);
	LUT4 #(
		.INIT('h0080)
	) name1648 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4660_
	);
	LUT4 #(
		.INIT('h0020)
	) name1649 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4661_
	);
	LUT4 #(
		.INIT('h0001)
	) name1650 (
		_w4658_,
		_w4659_,
		_w4660_,
		_w4661_,
		_w4662_
	);
	LUT4 #(
		.INIT('h0200)
	) name1651 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4663_
	);
	LUT4 #(
		.INIT('h0800)
	) name1652 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4664_
	);
	LUT4 #(
		.INIT('h2000)
	) name1653 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4665_
	);
	LUT4 #(
		.INIT('h8000)
	) name1654 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4666_
	);
	LUT4 #(
		.INIT('h0001)
	) name1655 (
		_w4663_,
		_w4664_,
		_w4665_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h7)
	) name1656 (
		_w4662_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h0080)
	) name1657 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4669_
	);
	LUT4 #(
		.INIT('h0020)
	) name1658 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4670_
	);
	LUT4 #(
		.INIT('h2000)
	) name1659 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4671_
	);
	LUT4 #(
		.INIT('h8000)
	) name1660 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4672_
	);
	LUT4 #(
		.INIT('h0001)
	) name1661 (
		_w4669_,
		_w4670_,
		_w4671_,
		_w4672_,
		_w4673_
	);
	LUT4 #(
		.INIT('h0200)
	) name1662 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4674_
	);
	LUT4 #(
		.INIT('h0800)
	) name1663 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4675_
	);
	LUT4 #(
		.INIT('h0002)
	) name1664 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4676_
	);
	LUT4 #(
		.INIT('h0008)
	) name1665 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4677_
	);
	LUT4 #(
		.INIT('h0001)
	) name1666 (
		_w4674_,
		_w4675_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h7)
	) name1667 (
		_w4673_,
		_w4678_,
		_w4679_
	);
	LUT4 #(
		.INIT('h0080)
	) name1668 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4680_
	);
	LUT4 #(
		.INIT('h0020)
	) name1669 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4681_
	);
	LUT4 #(
		.INIT('h2000)
	) name1670 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4682_
	);
	LUT4 #(
		.INIT('h8000)
	) name1671 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4683_
	);
	LUT4 #(
		.INIT('h0001)
	) name1672 (
		_w4680_,
		_w4681_,
		_w4682_,
		_w4683_,
		_w4684_
	);
	LUT4 #(
		.INIT('h0002)
	) name1673 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4685_
	);
	LUT4 #(
		.INIT('h0008)
	) name1674 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4686_
	);
	LUT4 #(
		.INIT('h0200)
	) name1675 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4687_
	);
	LUT4 #(
		.INIT('h0800)
	) name1676 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4688_
	);
	LUT4 #(
		.INIT('h0001)
	) name1677 (
		_w4685_,
		_w4686_,
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h7)
	) name1678 (
		_w4684_,
		_w4689_,
		_w4690_
	);
	LUT4 #(
		.INIT('h0200)
	) name1679 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4691_
	);
	LUT4 #(
		.INIT('h0800)
	) name1680 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4692_
	);
	LUT4 #(
		.INIT('h0080)
	) name1681 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4693_
	);
	LUT4 #(
		.INIT('h0020)
	) name1682 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4694_
	);
	LUT4 #(
		.INIT('h0001)
	) name1683 (
		_w4691_,
		_w4692_,
		_w4693_,
		_w4694_,
		_w4695_
	);
	LUT4 #(
		.INIT('h0002)
	) name1684 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4696_
	);
	LUT4 #(
		.INIT('h0008)
	) name1685 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4697_
	);
	LUT4 #(
		.INIT('h2000)
	) name1686 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4698_
	);
	LUT4 #(
		.INIT('h8000)
	) name1687 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4699_
	);
	LUT4 #(
		.INIT('h0001)
	) name1688 (
		_w4696_,
		_w4697_,
		_w4698_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h7)
	) name1689 (
		_w4695_,
		_w4700_,
		_w4701_
	);
	LUT4 #(
		.INIT('h0080)
	) name1690 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4702_
	);
	LUT4 #(
		.INIT('h0020)
	) name1691 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4703_
	);
	LUT4 #(
		.INIT('h0002)
	) name1692 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4704_
	);
	LUT4 #(
		.INIT('h0008)
	) name1693 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4705_
	);
	LUT4 #(
		.INIT('h0001)
	) name1694 (
		_w4702_,
		_w4703_,
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT4 #(
		.INIT('h2000)
	) name1695 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4707_
	);
	LUT4 #(
		.INIT('h8000)
	) name1696 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4708_
	);
	LUT4 #(
		.INIT('h0200)
	) name1697 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4709_
	);
	LUT4 #(
		.INIT('h0800)
	) name1698 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4710_
	);
	LUT4 #(
		.INIT('h0001)
	) name1699 (
		_w4707_,
		_w4708_,
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h7)
	) name1700 (
		_w4706_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('h0080)
	) name1701 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4713_
	);
	LUT4 #(
		.INIT('h0020)
	) name1702 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4714_
	);
	LUT4 #(
		.INIT('h0200)
	) name1703 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4715_
	);
	LUT4 #(
		.INIT('h0800)
	) name1704 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4716_
	);
	LUT4 #(
		.INIT('h0001)
	) name1705 (
		_w4713_,
		_w4714_,
		_w4715_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('h0002)
	) name1706 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4718_
	);
	LUT4 #(
		.INIT('h0008)
	) name1707 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4719_
	);
	LUT4 #(
		.INIT('h2000)
	) name1708 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4720_
	);
	LUT4 #(
		.INIT('h8000)
	) name1709 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4721_
	);
	LUT4 #(
		.INIT('h0001)
	) name1710 (
		_w4718_,
		_w4719_,
		_w4720_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h7)
	) name1711 (
		_w4717_,
		_w4722_,
		_w4723_
	);
	LUT4 #(
		.INIT('h0080)
	) name1712 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4724_
	);
	LUT4 #(
		.INIT('h0020)
	) name1713 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4725_
	);
	LUT4 #(
		.INIT('h2000)
	) name1714 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4726_
	);
	LUT4 #(
		.INIT('h8000)
	) name1715 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4727_
	);
	LUT4 #(
		.INIT('h0001)
	) name1716 (
		_w4724_,
		_w4725_,
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('h0800)
	) name1717 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4729_
	);
	LUT4 #(
		.INIT('h0200)
	) name1718 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4730_
	);
	LUT4 #(
		.INIT('h0002)
	) name1719 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4731_
	);
	LUT4 #(
		.INIT('h0008)
	) name1720 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4732_
	);
	LUT4 #(
		.INIT('h0001)
	) name1721 (
		_w4729_,
		_w4730_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h7)
	) name1722 (
		_w4728_,
		_w4733_,
		_w4734_
	);
	LUT4 #(
		.INIT('h0080)
	) name1723 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4735_
	);
	LUT4 #(
		.INIT('h0020)
	) name1724 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4736_
	);
	LUT4 #(
		.INIT('h2000)
	) name1725 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4737_
	);
	LUT4 #(
		.INIT('h8000)
	) name1726 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4738_
	);
	LUT4 #(
		.INIT('h0001)
	) name1727 (
		_w4735_,
		_w4736_,
		_w4737_,
		_w4738_,
		_w4739_
	);
	LUT4 #(
		.INIT('h0002)
	) name1728 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4740_
	);
	LUT4 #(
		.INIT('h0008)
	) name1729 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4741_
	);
	LUT4 #(
		.INIT('h0200)
	) name1730 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4742_
	);
	LUT4 #(
		.INIT('h0800)
	) name1731 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4743_
	);
	LUT4 #(
		.INIT('h0001)
	) name1732 (
		_w4740_,
		_w4741_,
		_w4742_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h7)
	) name1733 (
		_w4739_,
		_w4744_,
		_w4745_
	);
	LUT4 #(
		.INIT('h0002)
	) name1734 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4746_
	);
	LUT4 #(
		.INIT('h0008)
	) name1735 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4747_
	);
	LUT4 #(
		.INIT('h0200)
	) name1736 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4748_
	);
	LUT4 #(
		.INIT('h0800)
	) name1737 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4749_
	);
	LUT4 #(
		.INIT('h0001)
	) name1738 (
		_w4746_,
		_w4747_,
		_w4748_,
		_w4749_,
		_w4750_
	);
	LUT4 #(
		.INIT('h2000)
	) name1739 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4751_
	);
	LUT4 #(
		.INIT('h8000)
	) name1740 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4752_
	);
	LUT4 #(
		.INIT('h0080)
	) name1741 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4753_
	);
	LUT4 #(
		.INIT('h0020)
	) name1742 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4754_
	);
	LUT4 #(
		.INIT('h0001)
	) name1743 (
		_w4751_,
		_w4752_,
		_w4753_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h7)
	) name1744 (
		_w4750_,
		_w4755_,
		_w4756_
	);
	LUT4 #(
		.INIT('h0002)
	) name1745 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4757_
	);
	LUT4 #(
		.INIT('h0008)
	) name1746 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4758_
	);
	LUT4 #(
		.INIT('h2000)
	) name1747 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4759_
	);
	LUT4 #(
		.INIT('h8000)
	) name1748 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4760_
	);
	LUT4 #(
		.INIT('h0001)
	) name1749 (
		_w4757_,
		_w4758_,
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('h0080)
	) name1750 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4762_
	);
	LUT4 #(
		.INIT('h0020)
	) name1751 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4763_
	);
	LUT4 #(
		.INIT('h0200)
	) name1752 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4764_
	);
	LUT4 #(
		.INIT('h0800)
	) name1753 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4765_
	);
	LUT4 #(
		.INIT('h0001)
	) name1754 (
		_w4762_,
		_w4763_,
		_w4764_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h7)
	) name1755 (
		_w4761_,
		_w4766_,
		_w4767_
	);
	LUT4 #(
		.INIT('h0080)
	) name1756 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4768_
	);
	LUT4 #(
		.INIT('h0020)
	) name1757 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4769_
	);
	LUT4 #(
		.INIT('h0002)
	) name1758 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4770_
	);
	LUT4 #(
		.INIT('h0008)
	) name1759 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4771_
	);
	LUT4 #(
		.INIT('h0001)
	) name1760 (
		_w4768_,
		_w4769_,
		_w4770_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('h0200)
	) name1761 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4773_
	);
	LUT4 #(
		.INIT('h0800)
	) name1762 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4774_
	);
	LUT4 #(
		.INIT('h2000)
	) name1763 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4775_
	);
	LUT4 #(
		.INIT('h8000)
	) name1764 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4776_
	);
	LUT4 #(
		.INIT('h0001)
	) name1765 (
		_w4773_,
		_w4774_,
		_w4775_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h7)
	) name1766 (
		_w4772_,
		_w4777_,
		_w4778_
	);
	LUT4 #(
		.INIT('h0002)
	) name1767 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4779_
	);
	LUT4 #(
		.INIT('h0008)
	) name1768 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4780_
	);
	LUT4 #(
		.INIT('h2000)
	) name1769 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4781_
	);
	LUT4 #(
		.INIT('h8000)
	) name1770 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4782_
	);
	LUT4 #(
		.INIT('h0001)
	) name1771 (
		_w4779_,
		_w4780_,
		_w4781_,
		_w4782_,
		_w4783_
	);
	LUT4 #(
		.INIT('h0200)
	) name1772 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4784_
	);
	LUT4 #(
		.INIT('h0800)
	) name1773 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4785_
	);
	LUT4 #(
		.INIT('h0020)
	) name1774 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4786_
	);
	LUT4 #(
		.INIT('h0080)
	) name1775 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4787_
	);
	LUT4 #(
		.INIT('h0001)
	) name1776 (
		_w4784_,
		_w4785_,
		_w4786_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h7)
	) name1777 (
		_w4783_,
		_w4788_,
		_w4789_
	);
	LUT4 #(
		.INIT('h0200)
	) name1778 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4790_
	);
	LUT4 #(
		.INIT('h0800)
	) name1779 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4791_
	);
	LUT4 #(
		.INIT('h0002)
	) name1780 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4792_
	);
	LUT4 #(
		.INIT('h0008)
	) name1781 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4793_
	);
	LUT4 #(
		.INIT('h0001)
	) name1782 (
		_w4790_,
		_w4791_,
		_w4792_,
		_w4793_,
		_w4794_
	);
	LUT4 #(
		.INIT('h2000)
	) name1783 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4795_
	);
	LUT4 #(
		.INIT('h8000)
	) name1784 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4796_
	);
	LUT4 #(
		.INIT('h0080)
	) name1785 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4797_
	);
	LUT4 #(
		.INIT('h0020)
	) name1786 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4798_
	);
	LUT4 #(
		.INIT('h0001)
	) name1787 (
		_w4795_,
		_w4796_,
		_w4797_,
		_w4798_,
		_w4799_
	);
	LUT2 #(
		.INIT('h7)
	) name1788 (
		_w4794_,
		_w4799_,
		_w4800_
	);
	LUT4 #(
		.INIT('h0002)
	) name1789 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4801_
	);
	LUT4 #(
		.INIT('h0008)
	) name1790 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4802_
	);
	LUT4 #(
		.INIT('h0200)
	) name1791 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4803_
	);
	LUT4 #(
		.INIT('h0800)
	) name1792 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4804_
	);
	LUT4 #(
		.INIT('h0001)
	) name1793 (
		_w4801_,
		_w4802_,
		_w4803_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('h2000)
	) name1794 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4806_
	);
	LUT4 #(
		.INIT('h8000)
	) name1795 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4807_
	);
	LUT4 #(
		.INIT('h0080)
	) name1796 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4808_
	);
	LUT4 #(
		.INIT('h0020)
	) name1797 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4809_
	);
	LUT4 #(
		.INIT('h0001)
	) name1798 (
		_w4806_,
		_w4807_,
		_w4808_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h7)
	) name1799 (
		_w4805_,
		_w4810_,
		_w4811_
	);
	LUT4 #(
		.INIT('h0200)
	) name1800 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4812_
	);
	LUT4 #(
		.INIT('h0800)
	) name1801 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4813_
	);
	LUT4 #(
		.INIT('h0002)
	) name1802 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4814_
	);
	LUT4 #(
		.INIT('h0008)
	) name1803 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4815_
	);
	LUT4 #(
		.INIT('h0001)
	) name1804 (
		_w4812_,
		_w4813_,
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT4 #(
		.INIT('h2000)
	) name1805 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4817_
	);
	LUT4 #(
		.INIT('h8000)
	) name1806 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4818_
	);
	LUT4 #(
		.INIT('h0080)
	) name1807 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4819_
	);
	LUT4 #(
		.INIT('h0020)
	) name1808 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4820_
	);
	LUT4 #(
		.INIT('h0001)
	) name1809 (
		_w4817_,
		_w4818_,
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h7)
	) name1810 (
		_w4816_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h0002)
	) name1811 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4823_
	);
	LUT4 #(
		.INIT('h0008)
	) name1812 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4824_
	);
	LUT4 #(
		.INIT('h2000)
	) name1813 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4825_
	);
	LUT4 #(
		.INIT('h8000)
	) name1814 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4826_
	);
	LUT4 #(
		.INIT('h0001)
	) name1815 (
		_w4823_,
		_w4824_,
		_w4825_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('h0200)
	) name1816 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4828_
	);
	LUT4 #(
		.INIT('h0800)
	) name1817 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4829_
	);
	LUT4 #(
		.INIT('h0020)
	) name1818 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4830_
	);
	LUT4 #(
		.INIT('h0080)
	) name1819 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w4831_
	);
	LUT4 #(
		.INIT('h0001)
	) name1820 (
		_w4828_,
		_w4829_,
		_w4830_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h7)
	) name1821 (
		_w4827_,
		_w4832_,
		_w4833_
	);
	LUT3 #(
		.INIT('h80)
	) name1822 (
		\configuration_pci_ta1_reg[25]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4834_
	);
	LUT3 #(
		.INIT('h80)
	) name1823 (
		\configuration_wb_err_addr_reg[25]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4835_
	);
	LUT3 #(
		.INIT('h01)
	) name1824 (
		_w3933_,
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT3 #(
		.INIT('h80)
	) name1825 (
		\configuration_wb_err_cs_bit31_24_reg[25]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4837_
	);
	LUT4 #(
		.INIT('h8000)
	) name1826 (
		\configuration_pci_err_addr_reg[25]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h0031)
	) name1828 (
		\configuration_pci_ba0_bit31_8_reg[25]/NET0131 ,
		_w3043_,
		_w3831_,
		_w3874_,
		_w4840_
	);
	LUT3 #(
		.INIT('h80)
	) name1829 (
		_w4836_,
		_w4839_,
		_w4840_,
		_w4841_
	);
	LUT3 #(
		.INIT('h80)
	) name1830 (
		\configuration_pci_ba1_bit31_8_reg[25]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4842_
	);
	LUT3 #(
		.INIT('ha8)
	) name1831 (
		\configuration_pci_am1_reg[25]/NET0131 ,
		_w3834_,
		_w4842_,
		_w4843_
	);
	LUT4 #(
		.INIT('h8000)
	) name1832 (
		\configuration_pci_err_cs_bit31_24_reg[25]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4844_
	);
	LUT4 #(
		.INIT('h8000)
	) name1833 (
		\configuration_pci_err_data_reg[25]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4845_
	);
	LUT3 #(
		.INIT('h80)
	) name1834 (
		\configuration_wb_err_data_reg[25]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4846_
	);
	LUT3 #(
		.INIT('h01)
	) name1835 (
		_w4845_,
		_w4846_,
		_w4844_,
		_w4847_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w4843_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('hac00)
	) name1837 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]/NET0131 ,
		_w3260_,
		_w3852_,
		_w4849_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1838 (
		_w3801_,
		_w4841_,
		_w4848_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1839 (
		\output_backup_ad_out_reg[25]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4851_
	);
	LUT4 #(
		.INIT('h1055)
	) name1840 (
		\output_backup_tar_ad_en_out_reg/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4852_
	);
	LUT3 #(
		.INIT('h40)
	) name1841 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001 ,
		_w3018_,
		_w3019_,
		_w4853_
	);
	LUT4 #(
		.INIT('hc888)
	) name1842 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4854_
	);
	LUT4 #(
		.INIT('hff53)
	) name1843 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4855_
	);
	LUT3 #(
		.INIT('hb0)
	) name1844 (
		_w4853_,
		_w4854_,
		_w4855_,
		_w4856_
	);
	LUT3 #(
		.INIT('h51)
	) name1845 (
		_w4851_,
		_w4852_,
		_w4856_,
		_w4857_
	);
	LUT3 #(
		.INIT('h1f)
	) name1846 (
		_w3799_,
		_w4850_,
		_w4857_,
		_w4858_
	);
	LUT2 #(
		.INIT('h2)
	) name1847 (
		\configuration_pci_ba0_bit31_8_reg[26]/NET0131 ,
		_w3831_,
		_w4859_
	);
	LUT4 #(
		.INIT('h8000)
	) name1848 (
		\configuration_pci_err_addr_reg[26]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4860_
	);
	LUT3 #(
		.INIT('h80)
	) name1849 (
		\configuration_wb_err_addr_reg[26]/NET0131 ,
		_w3803_,
		_w3815_,
		_w4861_
	);
	LUT3 #(
		.INIT('h01)
	) name1850 (
		_w3874_,
		_w4860_,
		_w4861_,
		_w4862_
	);
	LUT4 #(
		.INIT('h8000)
	) name1851 (
		\configuration_pci_err_cs_bit31_24_reg[26]/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4863_
	);
	LUT3 #(
		.INIT('h80)
	) name1852 (
		\configuration_wb_err_data_reg[26]/NET0131 ,
		_w3809_,
		_w3803_,
		_w4864_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w4863_,
		_w4864_,
		_w4865_
	);
	LUT3 #(
		.INIT('h40)
	) name1854 (
		_w4859_,
		_w4862_,
		_w4865_,
		_w4866_
	);
	LUT3 #(
		.INIT('h80)
	) name1855 (
		\configuration_pci_ba1_bit31_8_reg[26]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4867_
	);
	LUT3 #(
		.INIT('ha8)
	) name1856 (
		\configuration_pci_am1_reg[26]/NET0131 ,
		_w3834_,
		_w4867_,
		_w4868_
	);
	LUT3 #(
		.INIT('h80)
	) name1857 (
		\configuration_pci_ta1_reg[26]/NET0131 ,
		_w3806_,
		_w3824_,
		_w4869_
	);
	LUT4 #(
		.INIT('h8000)
	) name1858 (
		\configuration_pci_err_data_reg[26]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4870_
	);
	LUT3 #(
		.INIT('h80)
	) name1859 (
		\configuration_wb_err_cs_bit31_24_reg[26]/NET0131 ,
		_w3809_,
		_w3818_,
		_w4871_
	);
	LUT3 #(
		.INIT('h01)
	) name1860 (
		_w4870_,
		_w4871_,
		_w4869_,
		_w4872_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w4868_,
		_w4872_,
		_w4873_
	);
	LUT4 #(
		.INIT('hac00)
	) name1862 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]/NET0131 ,
		_w3260_,
		_w3852_,
		_w4874_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1863 (
		_w3801_,
		_w4866_,
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1864 (
		\output_backup_ad_out_reg[26]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4876_
	);
	LUT3 #(
		.INIT('h40)
	) name1865 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001 ,
		_w3018_,
		_w3019_,
		_w4877_
	);
	LUT4 #(
		.INIT('hc888)
	) name1866 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4878_
	);
	LUT4 #(
		.INIT('hff53)
	) name1867 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4879_
	);
	LUT3 #(
		.INIT('hb0)
	) name1868 (
		_w4877_,
		_w4878_,
		_w4879_,
		_w4880_
	);
	LUT3 #(
		.INIT('h31)
	) name1869 (
		_w4852_,
		_w4876_,
		_w4880_,
		_w4881_
	);
	LUT3 #(
		.INIT('h1f)
	) name1870 (
		_w3799_,
		_w4875_,
		_w4881_,
		_w4882_
	);
	LUT4 #(
		.INIT('hee0f)
	) name1871 (
		\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4883_
	);
	LUT4 #(
		.INIT('h11f0)
	) name1872 (
		\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4884_
	);
	LUT2 #(
		.INIT('h2)
	) name1873 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w4883_,
		_w4885_
	);
	LUT3 #(
		.INIT('h40)
	) name1874 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001 ,
		_w3018_,
		_w3019_,
		_w4886_
	);
	LUT4 #(
		.INIT('h5444)
	) name1875 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4887_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1876 (
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4885_,
		_w4886_,
		_w4887_,
		_w4888_
	);
	LUT4 #(
		.INIT('hff53)
	) name1877 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4889_
	);
	LUT2 #(
		.INIT('hb)
	) name1878 (
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT4 #(
		.INIT('hee0f)
	) name1879 (
		\wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4891_
	);
	LUT4 #(
		.INIT('h11f0)
	) name1880 (
		\wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4892_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w4891_,
		_w4893_
	);
	LUT3 #(
		.INIT('h40)
	) name1882 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001 ,
		_w3018_,
		_w3019_,
		_w4894_
	);
	LUT4 #(
		.INIT('h5444)
	) name1883 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4895_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1884 (
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4893_,
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT4 #(
		.INIT('hff53)
	) name1885 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4897_
	);
	LUT2 #(
		.INIT('hb)
	) name1886 (
		_w4896_,
		_w4897_,
		_w4898_
	);
	LUT4 #(
		.INIT('hee0f)
	) name1887 (
		\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4899_
	);
	LUT4 #(
		.INIT('h11f0)
	) name1888 (
		\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w4900_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w4899_,
		_w4901_
	);
	LUT3 #(
		.INIT('h40)
	) name1890 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001 ,
		_w3018_,
		_w3019_,
		_w4902_
	);
	LUT4 #(
		.INIT('h5444)
	) name1891 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4903_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1892 (
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4901_,
		_w4902_,
		_w4903_,
		_w4904_
	);
	LUT4 #(
		.INIT('hff53)
	) name1893 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4905_
	);
	LUT2 #(
		.INIT('hb)
	) name1894 (
		_w4904_,
		_w4905_,
		_w4906_
	);
	LUT3 #(
		.INIT('h40)
	) name1895 (
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3823_,
		_w3804_,
		_w4907_
	);
	LUT4 #(
		.INIT('h8000)
	) name1896 (
		\configuration_pci_err_cs_bit0_reg/NET0131 ,
		_w3039_,
		_w3814_,
		_w3837_,
		_w4908_
	);
	LUT3 #(
		.INIT('h80)
	) name1897 (
		\configuration_interrupt_line_reg[0]/NET0131 ,
		_w3806_,
		_w3867_,
		_w4909_
	);
	LUT4 #(
		.INIT('h0002)
	) name1898 (
		_w3868_,
		_w4908_,
		_w4909_,
		_w4907_,
		_w4910_
	);
	LUT4 #(
		.INIT('h2000)
	) name1899 (
		\configuration_cache_line_size_reg_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3042_,
		_w3823_,
		_w4911_
	);
	LUT4 #(
		.INIT('h2000)
	) name1900 (
		\configuration_command_bit2_0_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w3040_,
		_w3042_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w4911_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		_w4910_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		\configuration_wb_err_data_reg[0]/NET0131 ,
		_w3809_,
		_w4915_
	);
	LUT2 #(
		.INIT('h8)
	) name1904 (
		\configuration_wb_ba2_bit0_reg/NET0131 ,
		_w3807_,
		_w4916_
	);
	LUT4 #(
		.INIT('h153f)
	) name1905 (
		\configuration_wb_ba1_bit0_reg/NET0131 ,
		\configuration_wb_err_addr_reg[0]/NET0131 ,
		_w3815_,
		_w3804_,
		_w4917_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1906 (
		_w3803_,
		_w4915_,
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT4 #(
		.INIT('h8000)
	) name1907 (
		\configuration_pci_err_data_reg[0]/NET0131 ,
		_w3822_,
		_w3814_,
		_w3837_,
		_w4919_
	);
	LUT3 #(
		.INIT('h80)
	) name1908 (
		\configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131 ,
		_w3806_,
		_w3818_,
		_w4920_
	);
	LUT3 #(
		.INIT('h80)
	) name1909 (
		\configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131 ,
		_w3042_,
		_w3818_,
		_w4921_
	);
	LUT3 #(
		.INIT('h80)
	) name1910 (
		\configuration_isr_bit2_0_reg[0]/NET0131 ,
		_w3956_,
		_w3958_,
		_w4922_
	);
	LUT4 #(
		.INIT('h0001)
	) name1911 (
		_w4919_,
		_w4920_,
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT3 #(
		.INIT('h80)
	) name1912 (
		\configuration_pci_am1_reg[31]/NET0131 ,
		_w3040_,
		_w3806_,
		_w4924_
	);
	LUT3 #(
		.INIT('h80)
	) name1913 (
		\configuration_wb_err_cs_bit0_reg/NET0131 ,
		_w3809_,
		_w3818_,
		_w4925_
	);
	LUT4 #(
		.INIT('h8000)
	) name1914 (
		\configuration_pci_err_addr_reg[0]/NET0131 ,
		_w3039_,
		_w3041_,
		_w3812_,
		_w4926_
	);
	LUT4 #(
		.INIT('h8000)
	) name1915 (
		\configuration_icr_bit2_0_reg[0]/NET0131 ,
		_w3041_,
		_w3802_,
		_w3812_,
		_w4927_
	);
	LUT4 #(
		.INIT('h0001)
	) name1916 (
		_w4924_,
		_w4925_,
		_w4926_,
		_w4927_,
		_w4928_
	);
	LUT3 #(
		.INIT('h40)
	) name1917 (
		_w4918_,
		_w4923_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('hac00)
	) name1918 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]/P0001 ,
		\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]/NET0131 ,
		_w3260_,
		_w3852_,
		_w4930_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1919 (
		_w3801_,
		_w4914_,
		_w4929_,
		_w4930_,
		_w4931_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1920 (
		\output_backup_ad_out_reg[0]/NET0131 ,
		_w3788_,
		_w3791_,
		_w3798_,
		_w4932_
	);
	LUT3 #(
		.INIT('h40)
	) name1921 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001 ,
		_w3018_,
		_w3019_,
		_w4933_
	);
	LUT4 #(
		.INIT('hc888)
	) name1922 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w4934_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT4 #(
		.INIT('h22a2)
	) name1924 (
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131 ,
		_w4936_
	);
	LUT4 #(
		.INIT('h0e02)
	) name1925 (
		\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]/NET0131 ,
		_w3972_,
		_w3974_,
		_w4936_,
		_w4937_
	);
	LUT3 #(
		.INIT('h02)
	) name1926 (
		\wishbone_slave_unit_pci_initiator_if_data_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w4938_
	);
	LUT3 #(
		.INIT('h07)
	) name1927 (
		_w3849_,
		_w4937_,
		_w4938_,
		_w4939_
	);
	LUT4 #(
		.INIT('h1311)
	) name1928 (
		_w4852_,
		_w4932_,
		_w4935_,
		_w4939_,
		_w4940_
	);
	LUT3 #(
		.INIT('h1f)
	) name1929 (
		_w3799_,
		_w4931_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w3165_,
		_w3639_,
		_w4942_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1931 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_check_for_serr_on_second_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w4943_
	);
	LUT2 #(
		.INIT('hd)
	) name1932 (
		_w3772_,
		_w4943_,
		_w4944_
	);
	LUT3 #(
		.INIT('h80)
	) name1933 (
		\configuration_command_bit6_reg/NET0131 ,
		\configuration_command_bit8_reg/NET0131 ,
		\configuration_init_complete_reg/NET0131 ,
		_w4945_
	);
	LUT3 #(
		.INIT('h20)
	) name1934 (
		_w3772_,
		_w4943_,
		_w4945_,
		_w4946_
	);
	LUT3 #(
		.INIT('hdf)
	) name1935 (
		_w3772_,
		_w4943_,
		_w4945_,
		_w4947_
	);
	LUT3 #(
		.INIT('h0e)
	) name1936 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 ,
		_w4948_
	);
	LUT4 #(
		.INIT('h007f)
	) name1937 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w4948_,
		_w4949_
	);
	LUT4 #(
		.INIT('hff80)
	) name1938 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w4948_,
		_w4950_
	);
	LUT3 #(
		.INIT('h74)
	) name1939 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w4891_,
		_w4951_
	);
	LUT3 #(
		.INIT('h8b)
	) name1940 (
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]/NET0131 ,
		_w4949_,
		_w4951_,
		_w4952_
	);
	LUT3 #(
		.INIT('h74)
	) name1941 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w4899_,
		_w4953_
	);
	LUT3 #(
		.INIT('h8b)
	) name1942 (
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]/NET0131 ,
		_w4949_,
		_w4953_,
		_w4954_
	);
	LUT3 #(
		.INIT('h74)
	) name1943 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w4883_,
		_w4955_
	);
	LUT3 #(
		.INIT('h8b)
	) name1944 (
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]/NET0131 ,
		_w4949_,
		_w4955_,
		_w4956_
	);
	LUT4 #(
		.INIT('h8000)
	) name1945 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w4957_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131 ,
		_w4958_
	);
	LUT4 #(
		.INIT('h8000)
	) name1947 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131 ,
		_w4957_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131 ,
		_w4960_
	);
	LUT4 #(
		.INIT('h8000)
	) name1949 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131 ,
		_w4961_
	);
	LUT2 #(
		.INIT('h8)
	) name1950 (
		_w4960_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		_w4959_,
		_w4962_,
		_w4963_
	);
	LUT4 #(
		.INIT('h8000)
	) name1952 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131 ,
		_w4959_,
		_w4962_,
		_w4964_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1953 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131 ,
		_w4959_,
		_w4962_,
		_w4965_
	);
	LUT3 #(
		.INIT('h8a)
	) name1954 (
		\wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131 ,
		_w3027_,
		_w3029_,
		_w4966_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1955 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4967_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT3 #(
		.INIT('h0e)
	) name1957 (
		_w3022_,
		_w4965_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('h10)
	) name1958 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001 ,
		_w3027_,
		_w3029_,
		_w4970_
	);
	LUT4 #(
		.INIT('h8c88)
	) name1959 (
		\wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4971_
	);
	LUT2 #(
		.INIT('h4)
	) name1960 (
		_w4970_,
		_w4971_,
		_w4972_
	);
	LUT4 #(
		.INIT('h8000)
	) name1961 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131 ,
		_w4959_,
		_w4973_
	);
	LUT4 #(
		.INIT('h8000)
	) name1962 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w4974_
	);
	LUT3 #(
		.INIT('h80)
	) name1963 (
		_w4960_,
		_w4973_,
		_w4974_,
		_w4975_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name1964 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		_w3022_,
		_w4972_,
		_w4975_,
		_w4976_
	);
	LUT3 #(
		.INIT('h80)
	) name1965 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131 ,
		_w4977_
	);
	LUT4 #(
		.INIT('h8000)
	) name1966 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 ,
		_w4964_,
		_w4977_,
		_w4978_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1967 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 ,
		_w4964_,
		_w4977_,
		_w4979_
	);
	LUT3 #(
		.INIT('h8a)
	) name1968 (
		\wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131 ,
		_w3027_,
		_w3029_,
		_w4980_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1969 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4981_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w4980_,
		_w4981_,
		_w4982_
	);
	LUT3 #(
		.INIT('h0e)
	) name1971 (
		_w3022_,
		_w4979_,
		_w4982_,
		_w4983_
	);
	LUT4 #(
		.INIT('h8000)
	) name1972 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 ,
		_w4984_
	);
	LUT4 #(
		.INIT('h8000)
	) name1973 (
		_w4960_,
		_w4973_,
		_w4974_,
		_w4984_,
		_w4985_
	);
	LUT3 #(
		.INIT('h8a)
	) name1974 (
		\wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131 ,
		_w3027_,
		_w3029_,
		_w4986_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1975 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4987_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w4986_,
		_w4987_,
		_w4988_
	);
	LUT4 #(
		.INIT('h00de)
	) name1977 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 ,
		_w3022_,
		_w4985_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131 ,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		_w4984_,
		_w4990_,
		_w4991_
	);
	LUT3 #(
		.INIT('h80)
	) name1980 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w4964_,
		_w4991_,
		_w4992_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1981 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131 ,
		_w4978_,
		_w4992_,
		_w4993_
	);
	LUT3 #(
		.INIT('h8a)
	) name1982 (
		\wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131 ,
		_w3027_,
		_w3029_,
		_w4994_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1983 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4995_
	);
	LUT2 #(
		.INIT('h4)
	) name1984 (
		_w4994_,
		_w4995_,
		_w4996_
	);
	LUT3 #(
		.INIT('h0e)
	) name1985 (
		_w3022_,
		_w4993_,
		_w4996_,
		_w4997_
	);
	LUT3 #(
		.INIT('h10)
	) name1986 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001 ,
		_w3027_,
		_w3029_,
		_w4998_
	);
	LUT4 #(
		.INIT('h8c88)
	) name1987 (
		\wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w4999_
	);
	LUT2 #(
		.INIT('h4)
	) name1988 (
		_w4998_,
		_w4999_,
		_w5000_
	);
	LUT4 #(
		.INIT('hff12)
	) name1989 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 ,
		_w3022_,
		_w4992_,
		_w5000_,
		_w5001_
	);
	LUT3 #(
		.INIT('h10)
	) name1990 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001 ,
		_w3027_,
		_w3029_,
		_w5002_
	);
	LUT4 #(
		.INIT('h8c88)
	) name1991 (
		\wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5003_
	);
	LUT2 #(
		.INIT('h4)
	) name1992 (
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT4 #(
		.INIT('h8000)
	) name1993 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 ,
		_w5005_
	);
	LUT4 #(
		.INIT('h8000)
	) name1994 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w4964_,
		_w4977_,
		_w5005_,
		_w5006_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name1995 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		_w3022_,
		_w5004_,
		_w5006_,
		_w5007_
	);
	LUT3 #(
		.INIT('h10)
	) name1996 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001 ,
		_w3027_,
		_w3029_,
		_w5008_
	);
	LUT4 #(
		.INIT('h8c88)
	) name1997 (
		\wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5009_
	);
	LUT2 #(
		.INIT('h4)
	) name1998 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		_w5011_
	);
	LUT3 #(
		.INIT('h80)
	) name2000 (
		_w4984_,
		_w4990_,
		_w5011_,
		_w5012_
	);
	LUT4 #(
		.INIT('h8000)
	) name2001 (
		_w4960_,
		_w4973_,
		_w4974_,
		_w5012_,
		_w5013_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name2002 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		_w3022_,
		_w5010_,
		_w5013_,
		_w5014_
	);
	LUT3 #(
		.INIT('h8a)
	) name2003 (
		\wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5015_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2004 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		_w5015_,
		_w5016_,
		_w5017_
	);
	LUT3 #(
		.INIT('h80)
	) name2006 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		_w5006_,
		_w5018_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name2007 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 ,
		_w3022_,
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT3 #(
		.INIT('h10)
	) name2008 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001 ,
		_w3027_,
		_w3029_,
		_w5020_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2009 (
		\wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5021_
	);
	LUT2 #(
		.INIT('h4)
	) name2010 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT4 #(
		.INIT('h8000)
	) name2011 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 ,
		_w5023_
	);
	LUT4 #(
		.INIT('h8000)
	) name2012 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w4964_,
		_w4991_,
		_w5023_,
		_w5024_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name2013 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 ,
		_w3022_,
		_w5022_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('h80)
	) name2014 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		_w5026_
	);
	LUT4 #(
		.INIT('h8000)
	) name2015 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		_w5006_,
		_w5026_,
		_w5027_
	);
	LUT4 #(
		.INIT('h8000)
	) name2016 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 ,
		_w5028_
	);
	LUT4 #(
		.INIT('h3222)
	) name2017 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		_w3022_,
		_w5006_,
		_w5028_,
		_w5029_
	);
	LUT3 #(
		.INIT('h10)
	) name2018 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001 ,
		_w3027_,
		_w3029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2019 (
		\wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name2020 (
		_w5030_,
		_w5031_,
		_w5032_
	);
	LUT3 #(
		.INIT('hf4)
	) name2021 (
		_w5027_,
		_w5029_,
		_w5032_,
		_w5033_
	);
	LUT3 #(
		.INIT('h80)
	) name2022 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]/NET0131 ,
		_w5013_,
		_w5026_,
		_w5034_
	);
	LUT3 #(
		.INIT('h10)
	) name2023 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001 ,
		_w3027_,
		_w3029_,
		_w5035_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2024 (
		\wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name2025 (
		_w5035_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('hff12)
	) name2026 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 ,
		_w3022_,
		_w5034_,
		_w5037_,
		_w5038_
	);
	LUT3 #(
		.INIT('h10)
	) name2027 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001 ,
		_w3027_,
		_w3029_,
		_w5039_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2028 (
		\wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w5039_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 ,
		_w5042_
	);
	LUT3 #(
		.INIT('h80)
	) name2031 (
		_w5006_,
		_w5028_,
		_w5042_,
		_w5043_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name2032 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131 ,
		_w3022_,
		_w5041_,
		_w5043_,
		_w5044_
	);
	LUT3 #(
		.INIT('h10)
	) name2033 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001 ,
		_w3027_,
		_w3029_,
		_w5045_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2034 (
		\wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name2035 (
		_w5045_,
		_w5046_,
		_w5047_
	);
	LUT3 #(
		.INIT('h80)
	) name2036 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131 ,
		_w5048_
	);
	LUT3 #(
		.INIT('h80)
	) name2037 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]/NET0131 ,
		_w5024_,
		_w5048_,
		_w5049_
	);
	LUT4 #(
		.INIT('hf1f2)
	) name2038 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131 ,
		_w3022_,
		_w5047_,
		_w5049_,
		_w5050_
	);
	LUT4 #(
		.INIT('h8000)
	) name2039 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]/NET0131 ,
		_w5051_
	);
	LUT3 #(
		.INIT('h80)
	) name2040 (
		_w5006_,
		_w5028_,
		_w5051_,
		_w5052_
	);
	LUT3 #(
		.INIT('h10)
	) name2041 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001 ,
		_w3027_,
		_w3029_,
		_w5053_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2042 (
		\wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5054_
	);
	LUT2 #(
		.INIT('h4)
	) name2043 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT4 #(
		.INIT('hff12)
	) name2044 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]/NET0131 ,
		_w3022_,
		_w5052_,
		_w5055_,
		_w5056_
	);
	LUT3 #(
		.INIT('h10)
	) name2045 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001 ,
		_w3027_,
		_w3029_,
		_w5057_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2046 (
		\wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5058_
	);
	LUT4 #(
		.INIT('h060c)
	) name2047 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]/NET0131 ,
		_w3022_,
		_w4957_,
		_w5059_
	);
	LUT3 #(
		.INIT('hf4)
	) name2048 (
		_w5057_,
		_w5058_,
		_w5059_,
		_w5060_
	);
	LUT4 #(
		.INIT('h2111)
	) name2049 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131 ,
		_w3022_,
		_w4957_,
		_w4958_,
		_w5061_
	);
	LUT3 #(
		.INIT('h8a)
	) name2050 (
		\wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5062_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2051 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5063_
	);
	LUT3 #(
		.INIT('h45)
	) name2052 (
		_w5061_,
		_w5062_,
		_w5063_,
		_w5064_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2053 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]/NET0131 ,
		_w4957_,
		_w4958_,
		_w5065_
	);
	LUT3 #(
		.INIT('h8a)
	) name2054 (
		\wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5066_
	);
	LUT3 #(
		.INIT('h20)
	) name2055 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001 ,
		_w3027_,
		_w3029_,
		_w5067_
	);
	LUT4 #(
		.INIT('heee4)
	) name2056 (
		_w3022_,
		_w5065_,
		_w5067_,
		_w5066_,
		_w5068_
	);
	LUT3 #(
		.INIT('h21)
	) name2057 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		_w3022_,
		_w4959_,
		_w5069_
	);
	LUT3 #(
		.INIT('h8a)
	) name2058 (
		\wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5070_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2059 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5071_
	);
	LUT2 #(
		.INIT('h4)
	) name2060 (
		_w5070_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w5069_,
		_w5072_,
		_w5073_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2062 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]/NET0131 ,
		_w4959_,
		_w5074_
	);
	LUT3 #(
		.INIT('h8a)
	) name2063 (
		\wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5075_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2064 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5076_
	);
	LUT2 #(
		.INIT('h4)
	) name2065 (
		_w5075_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h0e)
	) name2066 (
		_w3022_,
		_w5074_,
		_w5077_,
		_w5078_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2067 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w5079_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		_w3022_,
		_w5079_,
		_w5080_
	);
	LUT3 #(
		.INIT('h8a)
	) name2069 (
		\wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5081_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2070 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5082_
	);
	LUT3 #(
		.INIT('h45)
	) name2071 (
		_w5080_,
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT3 #(
		.INIT('h10)
	) name2072 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001 ,
		_w3027_,
		_w3029_,
		_w5084_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2073 (
		\wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5085_
	);
	LUT2 #(
		.INIT('h4)
	) name2074 (
		_w5084_,
		_w5085_,
		_w5086_
	);
	LUT3 #(
		.INIT('h80)
	) name2075 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		_w4964_,
		_w5087_
	);
	LUT4 #(
		.INIT('h8000)
	) name2076 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 ,
		_w4964_,
		_w5088_
	);
	LUT4 #(
		.INIT('h1333)
	) name2077 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w3022_,
		_w4964_,
		_w4977_,
		_w5089_
	);
	LUT4 #(
		.INIT('hfecc)
	) name2078 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]/NET0131 ,
		_w5086_,
		_w5088_,
		_w5089_,
		_w5090_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name2079 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]/NET0131 ,
		_w4960_,
		_w4963_,
		_w4973_,
		_w5091_
	);
	LUT3 #(
		.INIT('h8a)
	) name2080 (
		\wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5092_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2081 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5093_
	);
	LUT2 #(
		.INIT('h4)
	) name2082 (
		_w5092_,
		_w5093_,
		_w5094_
	);
	LUT3 #(
		.INIT('h0e)
	) name2083 (
		_w3022_,
		_w5091_,
		_w5094_,
		_w5095_
	);
	LUT4 #(
		.INIT('h2111)
	) name2084 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]/NET0131 ,
		_w3022_,
		_w4959_,
		_w4962_,
		_w5096_
	);
	LUT3 #(
		.INIT('h8a)
	) name2085 (
		\wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5097_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2086 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5098_
	);
	LUT2 #(
		.INIT('h4)
	) name2087 (
		_w5097_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w5096_,
		_w5099_,
		_w5100_
	);
	LUT3 #(
		.INIT('h8a)
	) name2089 (
		\wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5101_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2090 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5102_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		_w5101_,
		_w5102_,
		_w5103_
	);
	LUT4 #(
		.INIT('h00de)
	) name2092 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]/NET0131 ,
		_w3022_,
		_w4964_,
		_w5103_,
		_w5104_
	);
	LUT3 #(
		.INIT('h10)
	) name2093 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001 ,
		_w3027_,
		_w3029_,
		_w5105_
	);
	LUT4 #(
		.INIT('h8c88)
	) name2094 (
		\wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5106_
	);
	LUT2 #(
		.INIT('h4)
	) name2095 (
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT4 #(
		.INIT('hff12)
	) name2096 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]/NET0131 ,
		_w3022_,
		_w5087_,
		_w5107_,
		_w5108_
	);
	LUT3 #(
		.INIT('h21)
	) name2097 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]/NET0131 ,
		_w3022_,
		_w4957_,
		_w5109_
	);
	LUT3 #(
		.INIT('h8a)
	) name2098 (
		\wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5110_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2099 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5111_
	);
	LUT3 #(
		.INIT('h45)
	) name2100 (
		_w5109_,
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT4 #(
		.INIT('h0903)
	) name2101 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]/NET0131 ,
		_w3022_,
		_w4959_,
		_w5113_
	);
	LUT3 #(
		.INIT('h8a)
	) name2102 (
		\wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5114_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2103 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5115_
	);
	LUT2 #(
		.INIT('h4)
	) name2104 (
		_w5114_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w5113_,
		_w5116_,
		_w5117_
	);
	LUT3 #(
		.INIT('h8a)
	) name2106 (
		\wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5118_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2107 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5119_
	);
	LUT2 #(
		.INIT('h4)
	) name2108 (
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('h00de)
	) name2109 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131 ,
		_w3022_,
		_w4973_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('h0903)
	) name2110 (
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]/NET0131 ,
		_w3022_,
		_w4973_,
		_w5122_
	);
	LUT3 #(
		.INIT('h8a)
	) name2111 (
		\wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131 ,
		_w3027_,
		_w3029_,
		_w5123_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2112 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001 ,
		_w3022_,
		_w3027_,
		_w3029_,
		_w5124_
	);
	LUT2 #(
		.INIT('h4)
	) name2113 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w5122_,
		_w5125_,
		_w5126_
	);
	LUT4 #(
		.INIT('h333b)
	) name2115 (
		\pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131 ,
		\pci_target_unit_wishbone_master_wb_cyc_o_reg/NET0131 ,
		wbm_ack_i_pad,
		wbm_rty_i_pad,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name2116 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5128_
	);
	LUT3 #(
		.INIT('h20)
	) name2117 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]/P0001 ,
		_w3027_,
		_w3029_,
		_w5129_
	);
	LUT4 #(
		.INIT('hacaa)
	) name2118 (
		\wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]/P0001 ,
		_w3027_,
		_w3029_,
		_w5130_
	);
	LUT4 #(
		.INIT('hacaa)
	) name2119 (
		\wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]/P0001 ,
		_w3027_,
		_w3029_,
		_w5131_
	);
	LUT2 #(
		.INIT('h2)
	) name2120 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5132_
	);
	LUT4 #(
		.INIT('hacaa)
	) name2121 (
		\wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001 ,
		_w3027_,
		_w3029_,
		_w5133_
	);
	LUT4 #(
		.INIT('hacaa)
	) name2122 (
		\wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001 ,
		_w3027_,
		_w3029_,
		_w5134_
	);
	LUT2 #(
		.INIT('h2)
	) name2123 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5135_
	);
	LUT2 #(
		.INIT('h2)
	) name2124 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5136_
	);
	LUT2 #(
		.INIT('h2)
	) name2125 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5137_
	);
	LUT2 #(
		.INIT('h2)
	) name2126 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5138_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5139_
	);
	LUT2 #(
		.INIT('h2)
	) name2128 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5140_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5141_
	);
	LUT2 #(
		.INIT('h2)
	) name2130 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5142_
	);
	LUT2 #(
		.INIT('h2)
	) name2131 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5143_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5145_
	);
	LUT2 #(
		.INIT('h2)
	) name2134 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5146_
	);
	LUT2 #(
		.INIT('h2)
	) name2135 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5147_
	);
	LUT2 #(
		.INIT('h2)
	) name2136 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5148_
	);
	LUT2 #(
		.INIT('h2)
	) name2137 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5149_
	);
	LUT2 #(
		.INIT('h2)
	) name2138 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5150_
	);
	LUT2 #(
		.INIT('h2)
	) name2139 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5151_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5152_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name2142 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5154_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5155_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5156_
	);
	LUT2 #(
		.INIT('h2)
	) name2145 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5157_
	);
	LUT2 #(
		.INIT('h2)
	) name2146 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5159_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5160_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5161_
	);
	LUT2 #(
		.INIT('h2)
	) name2150 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5162_
	);
	LUT2 #(
		.INIT('h2)
	) name2151 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w5164_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		_w3081_,
		_w3097_,
		_w5165_
	);
	LUT4 #(
		.INIT('h2333)
	) name2154 (
		_w3165_,
		_w3168_,
		_w3149_,
		_w3147_,
		_w5166_
	);
	LUT3 #(
		.INIT('h35)
	) name2155 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131 ,
		_w5166_,
		_w5167_
	);
	LUT3 #(
		.INIT('h35)
	) name2156 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w5166_,
		_w5168_
	);
	LUT3 #(
		.INIT('h35)
	) name2157 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131 ,
		_w5166_,
		_w5169_
	);
	LUT3 #(
		.INIT('h35)
	) name2158 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w5166_,
		_w5170_
	);
	LUT4 #(
		.INIT('h0100)
	) name2159 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5171_
	);
	LUT4 #(
		.INIT('h0002)
	) name2160 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5172_
	);
	LUT4 #(
		.INIT('h135f)
	) name2161 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]/P0001 ,
		_w5171_,
		_w5172_,
		_w5173_
	);
	LUT4 #(
		.INIT('h0200)
	) name2162 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5174_
	);
	LUT4 #(
		.INIT('h0008)
	) name2163 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5175_
	);
	LUT4 #(
		.INIT('h135f)
	) name2164 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]/P0001 ,
		_w5174_,
		_w5175_,
		_w5176_
	);
	LUT4 #(
		.INIT('h0001)
	) name2165 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5177_
	);
	LUT4 #(
		.INIT('h0004)
	) name2166 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5178_
	);
	LUT4 #(
		.INIT('h153f)
	) name2167 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]/P0001 ,
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('h0080)
	) name2168 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5180_
	);
	LUT4 #(
		.INIT('h8000)
	) name2169 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5181_
	);
	LUT4 #(
		.INIT('h153f)
	) name2170 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]/P0001 ,
		_w5180_,
		_w5181_,
		_w5182_
	);
	LUT4 #(
		.INIT('h8000)
	) name2171 (
		_w5179_,
		_w5182_,
		_w5173_,
		_w5176_,
		_w5183_
	);
	LUT4 #(
		.INIT('h4000)
	) name2172 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5184_
	);
	LUT4 #(
		.INIT('h2000)
	) name2173 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5185_
	);
	LUT4 #(
		.INIT('h153f)
	) name2174 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]/P0001 ,
		_w5184_,
		_w5185_,
		_w5186_
	);
	LUT4 #(
		.INIT('h1000)
	) name2175 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5187_
	);
	LUT4 #(
		.INIT('h0400)
	) name2176 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5188_
	);
	LUT4 #(
		.INIT('h135f)
	) name2177 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]/P0001 ,
		_w5187_,
		_w5188_,
		_w5189_
	);
	LUT4 #(
		.INIT('h0040)
	) name2178 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5190_
	);
	LUT4 #(
		.INIT('h0010)
	) name2179 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5191_
	);
	LUT4 #(
		.INIT('h135f)
	) name2180 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]/P0001 ,
		_w5190_,
		_w5191_,
		_w5192_
	);
	LUT4 #(
		.INIT('h0800)
	) name2181 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5193_
	);
	LUT4 #(
		.INIT('h0020)
	) name2182 (
		_w5167_,
		_w5168_,
		_w5169_,
		_w5170_,
		_w5194_
	);
	LUT4 #(
		.INIT('h135f)
	) name2183 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]/P0001 ,
		_w5193_,
		_w5194_,
		_w5195_
	);
	LUT4 #(
		.INIT('h8000)
	) name2184 (
		_w5192_,
		_w5195_,
		_w5186_,
		_w5189_,
		_w5196_
	);
	LUT2 #(
		.INIT('h7)
	) name2185 (
		_w5183_,
		_w5196_,
		_w5197_
	);
	LUT4 #(
		.INIT('h135f)
	) name2186 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]/P0001 ,
		_w5178_,
		_w5184_,
		_w5198_
	);
	LUT4 #(
		.INIT('h135f)
	) name2187 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]/P0001 ,
		_w5174_,
		_w5175_,
		_w5199_
	);
	LUT4 #(
		.INIT('h135f)
	) name2188 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]/P0001 ,
		_w5187_,
		_w5188_,
		_w5200_
	);
	LUT4 #(
		.INIT('h153f)
	) name2189 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]/P0001 ,
		_w5180_,
		_w5181_,
		_w5201_
	);
	LUT4 #(
		.INIT('h8000)
	) name2190 (
		_w5200_,
		_w5201_,
		_w5198_,
		_w5199_,
		_w5202_
	);
	LUT4 #(
		.INIT('h135f)
	) name2191 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]/P0001 ,
		_w5171_,
		_w5191_,
		_w5203_
	);
	LUT4 #(
		.INIT('h153f)
	) name2192 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]/P0001 ,
		_w5172_,
		_w5194_,
		_w5204_
	);
	LUT4 #(
		.INIT('h135f)
	) name2193 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]/P0001 ,
		_w5193_,
		_w5185_,
		_w5205_
	);
	LUT4 #(
		.INIT('h153f)
	) name2194 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]/P0001 ,
		_w5177_,
		_w5190_,
		_w5206_
	);
	LUT4 #(
		.INIT('h8000)
	) name2195 (
		_w5205_,
		_w5206_,
		_w5203_,
		_w5204_,
		_w5207_
	);
	LUT2 #(
		.INIT('h7)
	) name2196 (
		_w5202_,
		_w5207_,
		_w5208_
	);
	LUT4 #(
		.INIT('h153f)
	) name2197 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]/P0001 ,
		_w5178_,
		_w5190_,
		_w5209_
	);
	LUT4 #(
		.INIT('h135f)
	) name2198 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]/P0001 ,
		_w5174_,
		_w5175_,
		_w5210_
	);
	LUT4 #(
		.INIT('h135f)
	) name2199 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]/P0001 ,
		_w5181_,
		_w5187_,
		_w5211_
	);
	LUT4 #(
		.INIT('h135f)
	) name2200 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]/P0001 ,
		_w5180_,
		_w5194_,
		_w5212_
	);
	LUT4 #(
		.INIT('h8000)
	) name2201 (
		_w5211_,
		_w5212_,
		_w5209_,
		_w5210_,
		_w5213_
	);
	LUT4 #(
		.INIT('h135f)
	) name2202 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]/P0001 ,
		_w5171_,
		_w5191_,
		_w5214_
	);
	LUT4 #(
		.INIT('h135f)
	) name2203 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]/P0001 ,
		_w5184_,
		_w5188_,
		_w5215_
	);
	LUT4 #(
		.INIT('h135f)
	) name2204 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]/P0001 ,
		_w5193_,
		_w5185_,
		_w5216_
	);
	LUT4 #(
		.INIT('h135f)
	) name2205 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]/P0001 ,
		_w5177_,
		_w5172_,
		_w5217_
	);
	LUT4 #(
		.INIT('h8000)
	) name2206 (
		_w5216_,
		_w5217_,
		_w5214_,
		_w5215_,
		_w5218_
	);
	LUT2 #(
		.INIT('h7)
	) name2207 (
		_w5213_,
		_w5218_,
		_w5219_
	);
	LUT4 #(
		.INIT('h135f)
	) name2208 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]/P0001 ,
		_w5171_,
		_w5185_,
		_w5220_
	);
	LUT4 #(
		.INIT('h135f)
	) name2209 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]/P0001 ,
		_w5190_,
		_w5191_,
		_w5221_
	);
	LUT4 #(
		.INIT('h153f)
	) name2210 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]/P0001 ,
		_w5172_,
		_w5194_,
		_w5222_
	);
	LUT4 #(
		.INIT('h153f)
	) name2211 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]/P0001 ,
		_w5177_,
		_w5178_,
		_w5223_
	);
	LUT4 #(
		.INIT('h8000)
	) name2212 (
		_w5222_,
		_w5223_,
		_w5220_,
		_w5221_,
		_w5224_
	);
	LUT4 #(
		.INIT('h153f)
	) name2213 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]/P0001 ,
		_w5180_,
		_w5193_,
		_w5225_
	);
	LUT4 #(
		.INIT('h135f)
	) name2214 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]/P0001 ,
		_w5187_,
		_w5188_,
		_w5226_
	);
	LUT4 #(
		.INIT('h135f)
	) name2215 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]/P0001 ,
		_w5174_,
		_w5175_,
		_w5227_
	);
	LUT4 #(
		.INIT('h135f)
	) name2216 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]/P0001 ,
		_w5181_,
		_w5184_,
		_w5228_
	);
	LUT4 #(
		.INIT('h8000)
	) name2217 (
		_w5227_,
		_w5228_,
		_w5225_,
		_w5226_,
		_w5229_
	);
	LUT2 #(
		.INIT('h7)
	) name2218 (
		_w5224_,
		_w5229_,
		_w5230_
	);
	LUT4 #(
		.INIT('h153f)
	) name2219 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]/P0001 ,
		_w5172_,
		_w5191_,
		_w5231_
	);
	LUT4 #(
		.INIT('h135f)
	) name2220 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]/P0001 ,
		_w5193_,
		_w5185_,
		_w5232_
	);
	LUT4 #(
		.INIT('h153f)
	) name2221 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]/P0001 ,
		_w5177_,
		_w5178_,
		_w5233_
	);
	LUT4 #(
		.INIT('h153f)
	) name2222 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]/P0001 ,
		_w5180_,
		_w5181_,
		_w5234_
	);
	LUT4 #(
		.INIT('h8000)
	) name2223 (
		_w5233_,
		_w5234_,
		_w5231_,
		_w5232_,
		_w5235_
	);
	LUT4 #(
		.INIT('h153f)
	) name2224 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]/P0001 ,
		_w5175_,
		_w5190_,
		_w5236_
	);
	LUT4 #(
		.INIT('h135f)
	) name2225 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]/P0001 ,
		_w5187_,
		_w5188_,
		_w5237_
	);
	LUT4 #(
		.INIT('h135f)
	) name2226 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]/P0001 ,
		_w5171_,
		_w5184_,
		_w5238_
	);
	LUT4 #(
		.INIT('h135f)
	) name2227 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]/P0001 ,
		_w5174_,
		_w5194_,
		_w5239_
	);
	LUT4 #(
		.INIT('h8000)
	) name2228 (
		_w5238_,
		_w5239_,
		_w5236_,
		_w5237_,
		_w5240_
	);
	LUT2 #(
		.INIT('h7)
	) name2229 (
		_w5235_,
		_w5240_,
		_w5241_
	);
	LUT4 #(
		.INIT('h153f)
	) name2230 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]/P0001 ,
		_w5174_,
		_w5185_,
		_w5242_
	);
	LUT4 #(
		.INIT('h135f)
	) name2231 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]/P0001 ,
		_w5171_,
		_w5184_,
		_w5243_
	);
	LUT4 #(
		.INIT('h153f)
	) name2232 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]/P0001 ,
		_w5172_,
		_w5194_,
		_w5244_
	);
	LUT4 #(
		.INIT('h135f)
	) name2233 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]/P0001 ,
		_w5187_,
		_w5188_,
		_w5245_
	);
	LUT4 #(
		.INIT('h8000)
	) name2234 (
		_w5244_,
		_w5245_,
		_w5242_,
		_w5243_,
		_w5246_
	);
	LUT4 #(
		.INIT('h135f)
	) name2235 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]/P0001 ,
		_w5180_,
		_w5175_,
		_w5247_
	);
	LUT4 #(
		.INIT('h153f)
	) name2236 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]/P0001 ,
		_w5177_,
		_w5178_,
		_w5248_
	);
	LUT4 #(
		.INIT('h135f)
	) name2237 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]/P0001 ,
		_w5190_,
		_w5191_,
		_w5249_
	);
	LUT4 #(
		.INIT('h135f)
	) name2238 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]/P0001 ,
		_w5181_,
		_w5193_,
		_w5250_
	);
	LUT4 #(
		.INIT('h8000)
	) name2239 (
		_w5249_,
		_w5250_,
		_w5247_,
		_w5248_,
		_w5251_
	);
	LUT2 #(
		.INIT('h7)
	) name2240 (
		_w5246_,
		_w5251_,
		_w5252_
	);
	LUT4 #(
		.INIT('h153f)
	) name2241 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]/P0001 ,
		_w5174_,
		_w5185_,
		_w5253_
	);
	LUT4 #(
		.INIT('h135f)
	) name2242 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]/P0001 ,
		_w5171_,
		_w5184_,
		_w5254_
	);
	LUT4 #(
		.INIT('h153f)
	) name2243 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]/P0001 ,
		_w5177_,
		_w5178_,
		_w5255_
	);
	LUT4 #(
		.INIT('h153f)
	) name2244 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]/P0001 ,
		_w5180_,
		_w5181_,
		_w5256_
	);
	LUT4 #(
		.INIT('h8000)
	) name2245 (
		_w5255_,
		_w5256_,
		_w5253_,
		_w5254_,
		_w5257_
	);
	LUT4 #(
		.INIT('h153f)
	) name2246 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]/P0001 ,
		_w5172_,
		_w5175_,
		_w5258_
	);
	LUT4 #(
		.INIT('h135f)
	) name2247 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]/P0001 ,
		_w5187_,
		_w5188_,
		_w5259_
	);
	LUT4 #(
		.INIT('h135f)
	) name2248 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]/P0001 ,
		_w5190_,
		_w5191_,
		_w5260_
	);
	LUT4 #(
		.INIT('h135f)
	) name2249 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]/P0001 ,
		_w5193_,
		_w5194_,
		_w5261_
	);
	LUT4 #(
		.INIT('h8000)
	) name2250 (
		_w5260_,
		_w5261_,
		_w5258_,
		_w5259_,
		_w5262_
	);
	LUT2 #(
		.INIT('h7)
	) name2251 (
		_w5257_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('h153f)
	) name2252 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]/P0001 ,
		_w5172_,
		_w5185_,
		_w5264_
	);
	LUT4 #(
		.INIT('h135f)
	) name2253 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]/P0001 ,
		_w5174_,
		_w5175_,
		_w5265_
	);
	LUT4 #(
		.INIT('h135f)
	) name2254 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]/P0001 ,
		_w5187_,
		_w5188_,
		_w5266_
	);
	LUT4 #(
		.INIT('h153f)
	) name2255 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]/P0001 ,
		_w5180_,
		_w5181_,
		_w5267_
	);
	LUT4 #(
		.INIT('h8000)
	) name2256 (
		_w5266_,
		_w5267_,
		_w5264_,
		_w5265_,
		_w5268_
	);
	LUT4 #(
		.INIT('h135f)
	) name2257 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]/P0001 ,
		_w5171_,
		_w5193_,
		_w5269_
	);
	LUT4 #(
		.INIT('h153f)
	) name2258 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]/P0001 ,
		_w5177_,
		_w5178_,
		_w5270_
	);
	LUT4 #(
		.INIT('h135f)
	) name2259 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]/P0001 ,
		_w5190_,
		_w5191_,
		_w5271_
	);
	LUT4 #(
		.INIT('h135f)
	) name2260 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]/P0001 ,
		_w5194_,
		_w5184_,
		_w5272_
	);
	LUT4 #(
		.INIT('h8000)
	) name2261 (
		_w5271_,
		_w5272_,
		_w5269_,
		_w5270_,
		_w5273_
	);
	LUT2 #(
		.INIT('h7)
	) name2262 (
		_w5268_,
		_w5273_,
		_w5274_
	);
	LUT4 #(
		.INIT('h153f)
	) name2263 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]/P0001 ,
		_w5180_,
		_w5171_,
		_w5275_
	);
	LUT4 #(
		.INIT('h135f)
	) name2264 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]/P0001 ,
		_w5193_,
		_w5185_,
		_w5276_
	);
	LUT4 #(
		.INIT('h153f)
	) name2265 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]/P0001 ,
		_w5172_,
		_w5194_,
		_w5277_
	);
	LUT4 #(
		.INIT('h153f)
	) name2266 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]/P0001 ,
		_w5177_,
		_w5178_,
		_w5278_
	);
	LUT4 #(
		.INIT('h8000)
	) name2267 (
		_w5277_,
		_w5278_,
		_w5275_,
		_w5276_,
		_w5279_
	);
	LUT4 #(
		.INIT('h135f)
	) name2268 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]/P0001 ,
		_w5175_,
		_w5184_,
		_w5280_
	);
	LUT4 #(
		.INIT('h135f)
	) name2269 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]/P0001 ,
		_w5187_,
		_w5188_,
		_w5281_
	);
	LUT4 #(
		.INIT('h135f)
	) name2270 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]/P0001 ,
		_w5190_,
		_w5191_,
		_w5282_
	);
	LUT4 #(
		.INIT('h135f)
	) name2271 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]/P0001 ,
		_w5181_,
		_w5174_,
		_w5283_
	);
	LUT4 #(
		.INIT('h8000)
	) name2272 (
		_w5282_,
		_w5283_,
		_w5280_,
		_w5281_,
		_w5284_
	);
	LUT2 #(
		.INIT('h7)
	) name2273 (
		_w5279_,
		_w5284_,
		_w5285_
	);
	LUT4 #(
		.INIT('h153f)
	) name2274 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]/P0001 ,
		_w5178_,
		_w5171_,
		_w5286_
	);
	LUT4 #(
		.INIT('h135f)
	) name2275 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]/P0001 ,
		_w5174_,
		_w5175_,
		_w5287_
	);
	LUT4 #(
		.INIT('h135f)
	) name2276 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]/P0001 ,
		_w5187_,
		_w5188_,
		_w5288_
	);
	LUT4 #(
		.INIT('h153f)
	) name2277 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]/P0001 ,
		_w5172_,
		_w5194_,
		_w5289_
	);
	LUT4 #(
		.INIT('h8000)
	) name2278 (
		_w5288_,
		_w5289_,
		_w5286_,
		_w5287_,
		_w5290_
	);
	LUT4 #(
		.INIT('h135f)
	) name2279 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]/P0001 ,
		_w5191_,
		_w5184_,
		_w5291_
	);
	LUT4 #(
		.INIT('h153f)
	) name2280 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]/P0001 ,
		_w5180_,
		_w5181_,
		_w5292_
	);
	LUT4 #(
		.INIT('h135f)
	) name2281 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]/P0001 ,
		_w5193_,
		_w5185_,
		_w5293_
	);
	LUT4 #(
		.INIT('h153f)
	) name2282 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]/P0001 ,
		_w5177_,
		_w5190_,
		_w5294_
	);
	LUT4 #(
		.INIT('h8000)
	) name2283 (
		_w5293_,
		_w5294_,
		_w5291_,
		_w5292_,
		_w5295_
	);
	LUT2 #(
		.INIT('h7)
	) name2284 (
		_w5290_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('h135f)
	) name2285 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]/P0001 ,
		_w5191_,
		_w5185_,
		_w5297_
	);
	LUT4 #(
		.INIT('h153f)
	) name2286 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]/P0001 ,
		_w5177_,
		_w5178_,
		_w5298_
	);
	LUT4 #(
		.INIT('h135f)
	) name2287 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]/P0001 ,
		_w5174_,
		_w5175_,
		_w5299_
	);
	LUT4 #(
		.INIT('h153f)
	) name2288 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]/P0001 ,
		_w5172_,
		_w5194_,
		_w5300_
	);
	LUT4 #(
		.INIT('h8000)
	) name2289 (
		_w5299_,
		_w5300_,
		_w5297_,
		_w5298_,
		_w5301_
	);
	LUT4 #(
		.INIT('h135f)
	) name2290 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]/P0001 ,
		_w5181_,
		_w5190_,
		_w5302_
	);
	LUT4 #(
		.INIT('h135f)
	) name2291 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]/P0001 ,
		_w5171_,
		_w5184_,
		_w5303_
	);
	LUT4 #(
		.INIT('h135f)
	) name2292 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]/P0001 ,
		_w5187_,
		_w5188_,
		_w5304_
	);
	LUT4 #(
		.INIT('h153f)
	) name2293 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]/P0001 ,
		_w5180_,
		_w5193_,
		_w5305_
	);
	LUT4 #(
		.INIT('h8000)
	) name2294 (
		_w5304_,
		_w5305_,
		_w5302_,
		_w5303_,
		_w5306_
	);
	LUT2 #(
		.INIT('h7)
	) name2295 (
		_w5301_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('h153f)
	) name2296 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]/P0001 ,
		_w5178_,
		_w5171_,
		_w5308_
	);
	LUT4 #(
		.INIT('h135f)
	) name2297 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]/P0001 ,
		_w5190_,
		_w5191_,
		_w5309_
	);
	LUT4 #(
		.INIT('h153f)
	) name2298 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]/P0001 ,
		_w5180_,
		_w5181_,
		_w5310_
	);
	LUT4 #(
		.INIT('h135f)
	) name2299 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]/P0001 ,
		_w5187_,
		_w5188_,
		_w5311_
	);
	LUT4 #(
		.INIT('h8000)
	) name2300 (
		_w5310_,
		_w5311_,
		_w5308_,
		_w5309_,
		_w5312_
	);
	LUT4 #(
		.INIT('h153f)
	) name2301 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]/P0001 ,
		_w5184_,
		_w5185_,
		_w5313_
	);
	LUT4 #(
		.INIT('h153f)
	) name2302 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]/P0001 ,
		_w5172_,
		_w5194_,
		_w5314_
	);
	LUT4 #(
		.INIT('h135f)
	) name2303 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]/P0001 ,
		_w5174_,
		_w5175_,
		_w5315_
	);
	LUT4 #(
		.INIT('h135f)
	) name2304 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]/P0001 ,
		_w5177_,
		_w5193_,
		_w5316_
	);
	LUT4 #(
		.INIT('h8000)
	) name2305 (
		_w5315_,
		_w5316_,
		_w5313_,
		_w5314_,
		_w5317_
	);
	LUT2 #(
		.INIT('h7)
	) name2306 (
		_w5312_,
		_w5317_,
		_w5318_
	);
	LUT4 #(
		.INIT('h153f)
	) name2307 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]/P0001 ,
		_w5180_,
		_w5185_,
		_w5319_
	);
	LUT4 #(
		.INIT('h135f)
	) name2308 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]/P0001 ,
		_w5171_,
		_w5184_,
		_w5320_
	);
	LUT4 #(
		.INIT('h135f)
	) name2309 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]/P0001 ,
		_w5187_,
		_w5188_,
		_w5321_
	);
	LUT4 #(
		.INIT('h153f)
	) name2310 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]/P0001 ,
		_w5177_,
		_w5178_,
		_w5322_
	);
	LUT4 #(
		.INIT('h8000)
	) name2311 (
		_w5321_,
		_w5322_,
		_w5319_,
		_w5320_,
		_w5323_
	);
	LUT4 #(
		.INIT('h153f)
	) name2312 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]/P0001 ,
		_w5175_,
		_w5193_,
		_w5324_
	);
	LUT4 #(
		.INIT('h153f)
	) name2313 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]/P0001 ,
		_w5172_,
		_w5194_,
		_w5325_
	);
	LUT4 #(
		.INIT('h135f)
	) name2314 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]/P0001 ,
		_w5190_,
		_w5191_,
		_w5326_
	);
	LUT4 #(
		.INIT('h135f)
	) name2315 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]/P0001 ,
		_w5181_,
		_w5174_,
		_w5327_
	);
	LUT4 #(
		.INIT('h8000)
	) name2316 (
		_w5326_,
		_w5327_,
		_w5324_,
		_w5325_,
		_w5328_
	);
	LUT2 #(
		.INIT('h7)
	) name2317 (
		_w5323_,
		_w5328_,
		_w5329_
	);
	LUT4 #(
		.INIT('h153f)
	) name2318 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]/P0001 ,
		_w5180_,
		_w5191_,
		_w5330_
	);
	LUT4 #(
		.INIT('h135f)
	) name2319 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]/P0001 ,
		_w5171_,
		_w5184_,
		_w5331_
	);
	LUT4 #(
		.INIT('h153f)
	) name2320 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]/P0001 ,
		_w5177_,
		_w5178_,
		_w5332_
	);
	LUT4 #(
		.INIT('h153f)
	) name2321 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]/P0001 ,
		_w5172_,
		_w5194_,
		_w5333_
	);
	LUT4 #(
		.INIT('h8000)
	) name2322 (
		_w5332_,
		_w5333_,
		_w5330_,
		_w5331_,
		_w5334_
	);
	LUT4 #(
		.INIT('h153f)
	) name2323 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]/P0001 ,
		_w5175_,
		_w5190_,
		_w5335_
	);
	LUT4 #(
		.INIT('h135f)
	) name2324 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]/P0001 ,
		_w5187_,
		_w5188_,
		_w5336_
	);
	LUT4 #(
		.INIT('h135f)
	) name2325 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]/P0001 ,
		_w5193_,
		_w5185_,
		_w5337_
	);
	LUT4 #(
		.INIT('h135f)
	) name2326 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]/P0001 ,
		_w5181_,
		_w5174_,
		_w5338_
	);
	LUT4 #(
		.INIT('h8000)
	) name2327 (
		_w5337_,
		_w5338_,
		_w5335_,
		_w5336_,
		_w5339_
	);
	LUT2 #(
		.INIT('h7)
	) name2328 (
		_w5334_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h153f)
	) name2329 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]/P0001 ,
		_w5184_,
		_w5185_,
		_w5341_
	);
	LUT4 #(
		.INIT('h135f)
	) name2330 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]/P0001 ,
		_w5174_,
		_w5175_,
		_w5342_
	);
	LUT4 #(
		.INIT('h153f)
	) name2331 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]/P0001 ,
		_w5172_,
		_w5194_,
		_w5343_
	);
	LUT4 #(
		.INIT('h135f)
	) name2332 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]/P0001 ,
		_w5187_,
		_w5188_,
		_w5344_
	);
	LUT4 #(
		.INIT('h8000)
	) name2333 (
		_w5343_,
		_w5344_,
		_w5341_,
		_w5342_,
		_w5345_
	);
	LUT4 #(
		.INIT('h153f)
	) name2334 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]/P0001 ,
		_w5178_,
		_w5171_,
		_w5346_
	);
	LUT4 #(
		.INIT('h153f)
	) name2335 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]/P0001 ,
		_w5180_,
		_w5181_,
		_w5347_
	);
	LUT4 #(
		.INIT('h135f)
	) name2336 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]/P0001 ,
		_w5190_,
		_w5191_,
		_w5348_
	);
	LUT4 #(
		.INIT('h135f)
	) name2337 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]/P0001 ,
		_w5177_,
		_w5193_,
		_w5349_
	);
	LUT4 #(
		.INIT('h8000)
	) name2338 (
		_w5348_,
		_w5349_,
		_w5346_,
		_w5347_,
		_w5350_
	);
	LUT2 #(
		.INIT('h7)
	) name2339 (
		_w5345_,
		_w5350_,
		_w5351_
	);
	LUT4 #(
		.INIT('h135f)
	) name2340 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]/P0001 ,
		_w5178_,
		_w5175_,
		_w5352_
	);
	LUT4 #(
		.INIT('h135f)
	) name2341 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]/P0001 ,
		_w5171_,
		_w5184_,
		_w5353_
	);
	LUT4 #(
		.INIT('h153f)
	) name2342 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]/P0001 ,
		_w5172_,
		_w5194_,
		_w5354_
	);
	LUT4 #(
		.INIT('h153f)
	) name2343 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]/P0001 ,
		_w5180_,
		_w5181_,
		_w5355_
	);
	LUT4 #(
		.INIT('h8000)
	) name2344 (
		_w5354_,
		_w5355_,
		_w5352_,
		_w5353_,
		_w5356_
	);
	LUT4 #(
		.INIT('h153f)
	) name2345 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]/P0001 ,
		_w5174_,
		_w5185_,
		_w5357_
	);
	LUT4 #(
		.INIT('h135f)
	) name2346 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]/P0001 ,
		_w5187_,
		_w5188_,
		_w5358_
	);
	LUT4 #(
		.INIT('h135f)
	) name2347 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]/P0001 ,
		_w5190_,
		_w5191_,
		_w5359_
	);
	LUT4 #(
		.INIT('h135f)
	) name2348 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]/P0001 ,
		_w5177_,
		_w5193_,
		_w5360_
	);
	LUT4 #(
		.INIT('h8000)
	) name2349 (
		_w5359_,
		_w5360_,
		_w5357_,
		_w5358_,
		_w5361_
	);
	LUT2 #(
		.INIT('h7)
	) name2350 (
		_w5356_,
		_w5361_,
		_w5362_
	);
	LUT4 #(
		.INIT('h135f)
	) name2351 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]/P0001 ,
		_w5171_,
		_w5175_,
		_w5363_
	);
	LUT4 #(
		.INIT('h153f)
	) name2352 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]/P0001 ,
		_w5172_,
		_w5194_,
		_w5364_
	);
	LUT4 #(
		.INIT('h135f)
	) name2353 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]/P0001 ,
		_w5193_,
		_w5185_,
		_w5365_
	);
	LUT4 #(
		.INIT('h153f)
	) name2354 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]/P0001 ,
		_w5177_,
		_w5178_,
		_w5366_
	);
	LUT4 #(
		.INIT('h8000)
	) name2355 (
		_w5365_,
		_w5366_,
		_w5363_,
		_w5364_,
		_w5367_
	);
	LUT4 #(
		.INIT('h135f)
	) name2356 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]/P0001 ,
		_w5181_,
		_w5174_,
		_w5368_
	);
	LUT4 #(
		.INIT('h135f)
	) name2357 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]/P0001 ,
		_w5190_,
		_w5191_,
		_w5369_
	);
	LUT4 #(
		.INIT('h135f)
	) name2358 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]/P0001 ,
		_w5187_,
		_w5188_,
		_w5370_
	);
	LUT4 #(
		.INIT('h135f)
	) name2359 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]/P0001 ,
		_w5180_,
		_w5184_,
		_w5371_
	);
	LUT4 #(
		.INIT('h8000)
	) name2360 (
		_w5370_,
		_w5371_,
		_w5368_,
		_w5369_,
		_w5372_
	);
	LUT2 #(
		.INIT('h7)
	) name2361 (
		_w5367_,
		_w5372_,
		_w5373_
	);
	LUT4 #(
		.INIT('h153f)
	) name2362 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001 ,
		_w5171_,
		_w5187_,
		_w5374_
	);
	LUT4 #(
		.INIT('h153f)
	) name2363 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001 ,
		_w5174_,
		_w5193_,
		_w5375_
	);
	LUT4 #(
		.INIT('h135f)
	) name2364 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001 ,
		_w5180_,
		_w5175_,
		_w5376_
	);
	LUT4 #(
		.INIT('h135f)
	) name2365 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001 ,
		_w5177_,
		_w5188_,
		_w5377_
	);
	LUT4 #(
		.INIT('h8000)
	) name2366 (
		_w5376_,
		_w5377_,
		_w5374_,
		_w5375_,
		_w5378_
	);
	LUT4 #(
		.INIT('h135f)
	) name2367 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001 ,
		_w5181_,
		_w5194_,
		_w5379_
	);
	LUT4 #(
		.INIT('h135f)
	) name2368 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001 ,
		_w5178_,
		_w5184_,
		_w5380_
	);
	LUT4 #(
		.INIT('h135f)
	) name2369 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001 ,
		_w5191_,
		_w5185_,
		_w5381_
	);
	LUT4 #(
		.INIT('h153f)
	) name2370 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001 ,
		_w5172_,
		_w5190_,
		_w5382_
	);
	LUT4 #(
		.INIT('h8000)
	) name2371 (
		_w5381_,
		_w5382_,
		_w5379_,
		_w5380_,
		_w5383_
	);
	LUT2 #(
		.INIT('h7)
	) name2372 (
		_w5378_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('h153f)
	) name2373 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]/P0001 ,
		_w5185_,
		_w5187_,
		_w5385_
	);
	LUT4 #(
		.INIT('h135f)
	) name2374 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]/P0001 ,
		_w5174_,
		_w5175_,
		_w5386_
	);
	LUT4 #(
		.INIT('h153f)
	) name2375 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]/P0001 ,
		_w5177_,
		_w5178_,
		_w5387_
	);
	LUT4 #(
		.INIT('h153f)
	) name2376 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]/P0001 ,
		_w5172_,
		_w5194_,
		_w5388_
	);
	LUT4 #(
		.INIT('h8000)
	) name2377 (
		_w5387_,
		_w5388_,
		_w5385_,
		_w5386_,
		_w5389_
	);
	LUT4 #(
		.INIT('h135f)
	) name2378 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]/P0001 ,
		_w5191_,
		_w5193_,
		_w5390_
	);
	LUT4 #(
		.INIT('h153f)
	) name2379 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]/P0001 ,
		_w5180_,
		_w5181_,
		_w5391_
	);
	LUT4 #(
		.INIT('h135f)
	) name2380 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]/P0001 ,
		_w5171_,
		_w5184_,
		_w5392_
	);
	LUT4 #(
		.INIT('h135f)
	) name2381 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]/P0001 ,
		_w5190_,
		_w5188_,
		_w5393_
	);
	LUT4 #(
		.INIT('h8000)
	) name2382 (
		_w5392_,
		_w5393_,
		_w5390_,
		_w5391_,
		_w5394_
	);
	LUT2 #(
		.INIT('h7)
	) name2383 (
		_w5389_,
		_w5394_,
		_w5395_
	);
	LUT4 #(
		.INIT('h153f)
	) name2384 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]/P0001 ,
		_w5171_,
		_w5187_,
		_w5396_
	);
	LUT4 #(
		.INIT('h135f)
	) name2385 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]/P0001 ,
		_w5190_,
		_w5191_,
		_w5397_
	);
	LUT4 #(
		.INIT('h153f)
	) name2386 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]/P0001 ,
		_w5180_,
		_w5181_,
		_w5398_
	);
	LUT4 #(
		.INIT('h153f)
	) name2387 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]/P0001 ,
		_w5172_,
		_w5194_,
		_w5399_
	);
	LUT4 #(
		.INIT('h8000)
	) name2388 (
		_w5398_,
		_w5399_,
		_w5396_,
		_w5397_,
		_w5400_
	);
	LUT4 #(
		.INIT('h153f)
	) name2389 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]/P0001 ,
		_w5184_,
		_w5185_,
		_w5401_
	);
	LUT4 #(
		.INIT('h153f)
	) name2390 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]/P0001 ,
		_w5177_,
		_w5178_,
		_w5402_
	);
	LUT4 #(
		.INIT('h135f)
	) name2391 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]/P0001 ,
		_w5174_,
		_w5175_,
		_w5403_
	);
	LUT4 #(
		.INIT('h135f)
	) name2392 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]/P0001 ,
		_w5193_,
		_w5188_,
		_w5404_
	);
	LUT4 #(
		.INIT('h8000)
	) name2393 (
		_w5403_,
		_w5404_,
		_w5401_,
		_w5402_,
		_w5405_
	);
	LUT2 #(
		.INIT('h7)
	) name2394 (
		_w5400_,
		_w5405_,
		_w5406_
	);
	LUT4 #(
		.INIT('h135f)
	) name2395 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]/P0001 ,
		_w5191_,
		_w5185_,
		_w5407_
	);
	LUT4 #(
		.INIT('h135f)
	) name2396 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]/P0001 ,
		_w5171_,
		_w5184_,
		_w5408_
	);
	LUT4 #(
		.INIT('h153f)
	) name2397 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]/P0001 ,
		_w5172_,
		_w5194_,
		_w5409_
	);
	LUT4 #(
		.INIT('h135f)
	) name2398 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]/P0001 ,
		_w5187_,
		_w5188_,
		_w5410_
	);
	LUT4 #(
		.INIT('h8000)
	) name2399 (
		_w5409_,
		_w5410_,
		_w5407_,
		_w5408_,
		_w5411_
	);
	LUT4 #(
		.INIT('h135f)
	) name2400 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]/P0001 ,
		_w5177_,
		_w5193_,
		_w5412_
	);
	LUT4 #(
		.INIT('h153f)
	) name2401 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]/P0001 ,
		_w5180_,
		_w5181_,
		_w5413_
	);
	LUT4 #(
		.INIT('h135f)
	) name2402 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]/P0001 ,
		_w5174_,
		_w5175_,
		_w5414_
	);
	LUT4 #(
		.INIT('h153f)
	) name2403 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]/P0001 ,
		_w5178_,
		_w5190_,
		_w5415_
	);
	LUT4 #(
		.INIT('h8000)
	) name2404 (
		_w5414_,
		_w5415_,
		_w5412_,
		_w5413_,
		_w5416_
	);
	LUT2 #(
		.INIT('h7)
	) name2405 (
		_w5411_,
		_w5416_,
		_w5417_
	);
	LUT4 #(
		.INIT('h153f)
	) name2406 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]/P0001 ,
		_w5175_,
		_w5185_,
		_w5418_
	);
	LUT4 #(
		.INIT('h135f)
	) name2407 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]/P0001 ,
		_w5171_,
		_w5184_,
		_w5419_
	);
	LUT4 #(
		.INIT('h153f)
	) name2408 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]/P0001 ,
		_w5172_,
		_w5194_,
		_w5420_
	);
	LUT4 #(
		.INIT('h153f)
	) name2409 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]/P0001 ,
		_w5180_,
		_w5181_,
		_w5421_
	);
	LUT4 #(
		.INIT('h8000)
	) name2410 (
		_w5420_,
		_w5421_,
		_w5418_,
		_w5419_,
		_w5422_
	);
	LUT4 #(
		.INIT('h135f)
	) name2411 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]/P0001 ,
		_w5178_,
		_w5193_,
		_w5423_
	);
	LUT4 #(
		.INIT('h135f)
	) name2412 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]/P0001 ,
		_w5187_,
		_w5188_,
		_w5424_
	);
	LUT4 #(
		.INIT('h135f)
	) name2413 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]/P0001 ,
		_w5190_,
		_w5191_,
		_w5425_
	);
	LUT4 #(
		.INIT('h135f)
	) name2414 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]/P0001 ,
		_w5177_,
		_w5174_,
		_w5426_
	);
	LUT4 #(
		.INIT('h8000)
	) name2415 (
		_w5425_,
		_w5426_,
		_w5423_,
		_w5424_,
		_w5427_
	);
	LUT2 #(
		.INIT('h7)
	) name2416 (
		_w5422_,
		_w5427_,
		_w5428_
	);
	LUT4 #(
		.INIT('h153f)
	) name2417 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]/P0001 ,
		_w5172_,
		_w5175_,
		_w5429_
	);
	LUT4 #(
		.INIT('h135f)
	) name2418 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]/P0001 ,
		_w5171_,
		_w5184_,
		_w5430_
	);
	LUT4 #(
		.INIT('h135f)
	) name2419 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]/P0001 ,
		_w5187_,
		_w5188_,
		_w5431_
	);
	LUT4 #(
		.INIT('h153f)
	) name2420 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]/P0001 ,
		_w5180_,
		_w5181_,
		_w5432_
	);
	LUT4 #(
		.INIT('h8000)
	) name2421 (
		_w5431_,
		_w5432_,
		_w5429_,
		_w5430_,
		_w5433_
	);
	LUT4 #(
		.INIT('h153f)
	) name2422 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]/P0001 ,
		_w5174_,
		_w5185_,
		_w5434_
	);
	LUT4 #(
		.INIT('h153f)
	) name2423 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]/P0001 ,
		_w5177_,
		_w5178_,
		_w5435_
	);
	LUT4 #(
		.INIT('h135f)
	) name2424 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]/P0001 ,
		_w5190_,
		_w5191_,
		_w5436_
	);
	LUT4 #(
		.INIT('h135f)
	) name2425 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]/P0001 ,
		_w5193_,
		_w5194_,
		_w5437_
	);
	LUT4 #(
		.INIT('h8000)
	) name2426 (
		_w5436_,
		_w5437_,
		_w5434_,
		_w5435_,
		_w5438_
	);
	LUT2 #(
		.INIT('h7)
	) name2427 (
		_w5433_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('h153f)
	) name2428 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]/P0001 ,
		_w5172_,
		_w5191_,
		_w5440_
	);
	LUT4 #(
		.INIT('h135f)
	) name2429 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]/P0001 ,
		_w5174_,
		_w5175_,
		_w5441_
	);
	LUT4 #(
		.INIT('h153f)
	) name2430 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]/P0001 ,
		_w5180_,
		_w5181_,
		_w5442_
	);
	LUT4 #(
		.INIT('h135f)
	) name2431 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]/P0001 ,
		_w5187_,
		_w5188_,
		_w5443_
	);
	LUT4 #(
		.INIT('h8000)
	) name2432 (
		_w5442_,
		_w5443_,
		_w5440_,
		_w5441_,
		_w5444_
	);
	LUT4 #(
		.INIT('h135f)
	) name2433 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]/P0001 ,
		_w5171_,
		_w5190_,
		_w5445_
	);
	LUT4 #(
		.INIT('h153f)
	) name2434 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]/P0001 ,
		_w5177_,
		_w5178_,
		_w5446_
	);
	LUT4 #(
		.INIT('h135f)
	) name2435 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]/P0001 ,
		_w5193_,
		_w5185_,
		_w5447_
	);
	LUT4 #(
		.INIT('h135f)
	) name2436 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]/P0001 ,
		_w5194_,
		_w5184_,
		_w5448_
	);
	LUT4 #(
		.INIT('h8000)
	) name2437 (
		_w5447_,
		_w5448_,
		_w5445_,
		_w5446_,
		_w5449_
	);
	LUT2 #(
		.INIT('h7)
	) name2438 (
		_w5444_,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('h153f)
	) name2439 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]/P0001 ,
		_w5180_,
		_w5191_,
		_w5451_
	);
	LUT4 #(
		.INIT('h135f)
	) name2440 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]/P0001 ,
		_w5193_,
		_w5185_,
		_w5452_
	);
	LUT4 #(
		.INIT('h135f)
	) name2441 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]/P0001 ,
		_w5187_,
		_w5188_,
		_w5453_
	);
	LUT4 #(
		.INIT('h153f)
	) name2442 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]/P0001 ,
		_w5172_,
		_w5194_,
		_w5454_
	);
	LUT4 #(
		.INIT('h8000)
	) name2443 (
		_w5453_,
		_w5454_,
		_w5451_,
		_w5452_,
		_w5455_
	);
	LUT4 #(
		.INIT('h153f)
	) name2444 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]/P0001 ,
		_w5175_,
		_w5190_,
		_w5456_
	);
	LUT4 #(
		.INIT('h153f)
	) name2445 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]/P0001 ,
		_w5177_,
		_w5178_,
		_w5457_
	);
	LUT4 #(
		.INIT('h135f)
	) name2446 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]/P0001 ,
		_w5171_,
		_w5184_,
		_w5458_
	);
	LUT4 #(
		.INIT('h135f)
	) name2447 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]/P0001 ,
		_w5181_,
		_w5174_,
		_w5459_
	);
	LUT4 #(
		.INIT('h8000)
	) name2448 (
		_w5458_,
		_w5459_,
		_w5456_,
		_w5457_,
		_w5460_
	);
	LUT2 #(
		.INIT('h7)
	) name2449 (
		_w5455_,
		_w5460_,
		_w5461_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 ,
		_w4478_,
		_w5462_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2451 (
		\pci_target_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 ,
		\pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131 ,
		_w4478_,
		_w5463_
	);
	LUT4 #(
		.INIT('h153f)
	) name2452 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]/P0001 ,
		_w5172_,
		_w5185_,
		_w5464_
	);
	LUT4 #(
		.INIT('h135f)
	) name2453 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]/P0001 ,
		_w5171_,
		_w5184_,
		_w5465_
	);
	LUT4 #(
		.INIT('h153f)
	) name2454 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]/P0001 ,
		_w5180_,
		_w5181_,
		_w5466_
	);
	LUT4 #(
		.INIT('h153f)
	) name2455 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]/P0001 ,
		_w5177_,
		_w5178_,
		_w5467_
	);
	LUT4 #(
		.INIT('h8000)
	) name2456 (
		_w5466_,
		_w5467_,
		_w5464_,
		_w5465_,
		_w5468_
	);
	LUT4 #(
		.INIT('h153f)
	) name2457 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]/P0001 ,
		_w5175_,
		_w5193_,
		_w5469_
	);
	LUT4 #(
		.INIT('h135f)
	) name2458 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]/P0001 ,
		_w5187_,
		_w5188_,
		_w5470_
	);
	LUT4 #(
		.INIT('h135f)
	) name2459 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]/P0001 ,
		_w5190_,
		_w5191_,
		_w5471_
	);
	LUT4 #(
		.INIT('h135f)
	) name2460 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]/P0001 ,
		_w5174_,
		_w5194_,
		_w5472_
	);
	LUT4 #(
		.INIT('h8000)
	) name2461 (
		_w5471_,
		_w5472_,
		_w5469_,
		_w5470_,
		_w5473_
	);
	LUT2 #(
		.INIT('h7)
	) name2462 (
		_w5468_,
		_w5473_,
		_w5474_
	);
	LUT4 #(
		.INIT('h135f)
	) name2463 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]/P0001 ,
		_w5191_,
		_w5185_,
		_w5475_
	);
	LUT4 #(
		.INIT('h135f)
	) name2464 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]/P0001 ,
		_w5171_,
		_w5184_,
		_w5476_
	);
	LUT4 #(
		.INIT('h153f)
	) name2465 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]/P0001 ,
		_w5172_,
		_w5194_,
		_w5477_
	);
	LUT4 #(
		.INIT('h153f)
	) name2466 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]/P0001 ,
		_w5180_,
		_w5181_,
		_w5478_
	);
	LUT4 #(
		.INIT('h8000)
	) name2467 (
		_w5477_,
		_w5478_,
		_w5475_,
		_w5476_,
		_w5479_
	);
	LUT4 #(
		.INIT('h135f)
	) name2468 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]/P0001 ,
		_w5177_,
		_w5193_,
		_w5480_
	);
	LUT4 #(
		.INIT('h135f)
	) name2469 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]/P0001 ,
		_w5187_,
		_w5188_,
		_w5481_
	);
	LUT4 #(
		.INIT('h135f)
	) name2470 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]/P0001 ,
		_w5174_,
		_w5175_,
		_w5482_
	);
	LUT4 #(
		.INIT('h153f)
	) name2471 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]/P0001 ,
		_w5178_,
		_w5190_,
		_w5483_
	);
	LUT4 #(
		.INIT('h8000)
	) name2472 (
		_w5482_,
		_w5483_,
		_w5480_,
		_w5481_,
		_w5484_
	);
	LUT2 #(
		.INIT('h7)
	) name2473 (
		_w5479_,
		_w5484_,
		_w5485_
	);
	LUT4 #(
		.INIT('h135f)
	) name2474 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]/P0001 ,
		_w5191_,
		_w5185_,
		_w5486_
	);
	LUT4 #(
		.INIT('h135f)
	) name2475 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]/P0001 ,
		_w5171_,
		_w5184_,
		_w5487_
	);
	LUT4 #(
		.INIT('h153f)
	) name2476 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]/P0001 ,
		_w5177_,
		_w5178_,
		_w5488_
	);
	LUT4 #(
		.INIT('h153f)
	) name2477 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]/P0001 ,
		_w5180_,
		_w5181_,
		_w5489_
	);
	LUT4 #(
		.INIT('h8000)
	) name2478 (
		_w5488_,
		_w5489_,
		_w5486_,
		_w5487_,
		_w5490_
	);
	LUT4 #(
		.INIT('h153f)
	) name2479 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]/P0001 ,
		_w5172_,
		_w5190_,
		_w5491_
	);
	LUT4 #(
		.INIT('h135f)
	) name2480 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]/P0001 ,
		_w5187_,
		_w5188_,
		_w5492_
	);
	LUT4 #(
		.INIT('h135f)
	) name2481 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]/P0001 ,
		_w5174_,
		_w5175_,
		_w5493_
	);
	LUT4 #(
		.INIT('h135f)
	) name2482 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]/P0001 ,
		_w5193_,
		_w5194_,
		_w5494_
	);
	LUT4 #(
		.INIT('h8000)
	) name2483 (
		_w5493_,
		_w5494_,
		_w5491_,
		_w5492_,
		_w5495_
	);
	LUT2 #(
		.INIT('h7)
	) name2484 (
		_w5490_,
		_w5495_,
		_w5496_
	);
	LUT4 #(
		.INIT('h135f)
	) name2485 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]/P0001 ,
		_w5178_,
		_w5191_,
		_w5497_
	);
	LUT4 #(
		.INIT('h135f)
	) name2486 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]/P0001 ,
		_w5174_,
		_w5175_,
		_w5498_
	);
	LUT4 #(
		.INIT('h153f)
	) name2487 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]/P0001 ,
		_w5180_,
		_w5181_,
		_w5499_
	);
	LUT4 #(
		.INIT('h135f)
	) name2488 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]/P0001 ,
		_w5187_,
		_w5188_,
		_w5500_
	);
	LUT4 #(
		.INIT('h8000)
	) name2489 (
		_w5499_,
		_w5500_,
		_w5497_,
		_w5498_,
		_w5501_
	);
	LUT4 #(
		.INIT('h135f)
	) name2490 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]/P0001 ,
		_w5171_,
		_w5190_,
		_w5502_
	);
	LUT4 #(
		.INIT('h153f)
	) name2491 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]/P0001 ,
		_w5172_,
		_w5194_,
		_w5503_
	);
	LUT4 #(
		.INIT('h135f)
	) name2492 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]/P0001 ,
		_w5193_,
		_w5185_,
		_w5504_
	);
	LUT4 #(
		.INIT('h135f)
	) name2493 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]/P0001 ,
		_w5177_,
		_w5184_,
		_w5505_
	);
	LUT4 #(
		.INIT('h8000)
	) name2494 (
		_w5504_,
		_w5505_,
		_w5502_,
		_w5503_,
		_w5506_
	);
	LUT2 #(
		.INIT('h7)
	) name2495 (
		_w5501_,
		_w5506_,
		_w5507_
	);
	LUT4 #(
		.INIT('h153f)
	) name2496 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]/P0001 ,
		_w5175_,
		_w5187_,
		_w5508_
	);
	LUT4 #(
		.INIT('h135f)
	) name2497 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]/P0001 ,
		_w5193_,
		_w5185_,
		_w5509_
	);
	LUT4 #(
		.INIT('h153f)
	) name2498 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]/P0001 ,
		_w5177_,
		_w5178_,
		_w5510_
	);
	LUT4 #(
		.INIT('h153f)
	) name2499 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]/P0001 ,
		_w5172_,
		_w5194_,
		_w5511_
	);
	LUT4 #(
		.INIT('h8000)
	) name2500 (
		_w5510_,
		_w5511_,
		_w5508_,
		_w5509_,
		_w5512_
	);
	LUT4 #(
		.INIT('h135f)
	) name2501 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]/P0001 ,
		_w5171_,
		_w5174_,
		_w5513_
	);
	LUT4 #(
		.INIT('h153f)
	) name2502 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]/P0001 ,
		_w5180_,
		_w5181_,
		_w5514_
	);
	LUT4 #(
		.INIT('h135f)
	) name2503 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]/P0001 ,
		_w5190_,
		_w5191_,
		_w5515_
	);
	LUT4 #(
		.INIT('h135f)
	) name2504 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]/P0001 ,
		_w5184_,
		_w5188_,
		_w5516_
	);
	LUT4 #(
		.INIT('h8000)
	) name2505 (
		_w5515_,
		_w5516_,
		_w5513_,
		_w5514_,
		_w5517_
	);
	LUT2 #(
		.INIT('h7)
	) name2506 (
		_w5512_,
		_w5517_,
		_w5518_
	);
	LUT4 #(
		.INIT('h153f)
	) name2507 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]/P0001 ,
		_w5180_,
		_w5191_,
		_w5519_
	);
	LUT4 #(
		.INIT('h135f)
	) name2508 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]/P0001 ,
		_w5174_,
		_w5175_,
		_w5520_
	);
	LUT4 #(
		.INIT('h153f)
	) name2509 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]/P0001 ,
		_w5172_,
		_w5194_,
		_w5521_
	);
	LUT4 #(
		.INIT('h135f)
	) name2510 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]/P0001 ,
		_w5187_,
		_w5188_,
		_w5522_
	);
	LUT4 #(
		.INIT('h8000)
	) name2511 (
		_w5521_,
		_w5522_,
		_w5519_,
		_w5520_,
		_w5523_
	);
	LUT4 #(
		.INIT('h135f)
	) name2512 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]/P0001 ,
		_w5190_,
		_w5185_,
		_w5524_
	);
	LUT4 #(
		.INIT('h153f)
	) name2513 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]/P0001 ,
		_w5177_,
		_w5178_,
		_w5525_
	);
	LUT4 #(
		.INIT('h135f)
	) name2514 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]/P0001 ,
		_w5171_,
		_w5184_,
		_w5526_
	);
	LUT4 #(
		.INIT('h135f)
	) name2515 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]/P0001 ,
		_w5181_,
		_w5193_,
		_w5527_
	);
	LUT4 #(
		.INIT('h8000)
	) name2516 (
		_w5526_,
		_w5527_,
		_w5524_,
		_w5525_,
		_w5528_
	);
	LUT2 #(
		.INIT('h7)
	) name2517 (
		_w5523_,
		_w5528_,
		_w5529_
	);
	LUT4 #(
		.INIT('h153f)
	) name2518 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]/P0001 ,
		_w5180_,
		_w5185_,
		_w5530_
	);
	LUT4 #(
		.INIT('h135f)
	) name2519 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]/P0001 ,
		_w5174_,
		_w5175_,
		_w5531_
	);
	LUT4 #(
		.INIT('h153f)
	) name2520 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]/P0001 ,
		_w5177_,
		_w5178_,
		_w5532_
	);
	LUT4 #(
		.INIT('h153f)
	) name2521 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]/P0001 ,
		_w5172_,
		_w5194_,
		_w5533_
	);
	LUT4 #(
		.INIT('h8000)
	) name2522 (
		_w5532_,
		_w5533_,
		_w5530_,
		_w5531_,
		_w5534_
	);
	LUT4 #(
		.INIT('h135f)
	) name2523 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]/P0001 ,
		_w5191_,
		_w5193_,
		_w5535_
	);
	LUT4 #(
		.INIT('h135f)
	) name2524 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]/P0001 ,
		_w5187_,
		_w5188_,
		_w5536_
	);
	LUT4 #(
		.INIT('h135f)
	) name2525 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]/P0001 ,
		_w5171_,
		_w5184_,
		_w5537_
	);
	LUT4 #(
		.INIT('h135f)
	) name2526 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]/P0001 ,
		_w5181_,
		_w5190_,
		_w5538_
	);
	LUT4 #(
		.INIT('h8000)
	) name2527 (
		_w5537_,
		_w5538_,
		_w5535_,
		_w5536_,
		_w5539_
	);
	LUT2 #(
		.INIT('h7)
	) name2528 (
		_w5534_,
		_w5539_,
		_w5540_
	);
	LUT4 #(
		.INIT('h153f)
	) name2529 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]/P0001 ,
		_w5172_,
		_w5190_,
		_w5541_
	);
	LUT4 #(
		.INIT('h135f)
	) name2530 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]/P0001 ,
		_w5171_,
		_w5184_,
		_w5542_
	);
	LUT4 #(
		.INIT('h135f)
	) name2531 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]/P0001 ,
		_w5180_,
		_w5175_,
		_w5543_
	);
	LUT4 #(
		.INIT('h153f)
	) name2532 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]/P0001 ,
		_w5177_,
		_w5178_,
		_w5544_
	);
	LUT4 #(
		.INIT('h8000)
	) name2533 (
		_w5543_,
		_w5544_,
		_w5541_,
		_w5542_,
		_w5545_
	);
	LUT4 #(
		.INIT('h153f)
	) name2534 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]/P0001 ,
		_w5191_,
		_w5187_,
		_w5546_
	);
	LUT4 #(
		.INIT('h135f)
	) name2535 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]/P0001 ,
		_w5181_,
		_w5174_,
		_w5547_
	);
	LUT4 #(
		.INIT('h135f)
	) name2536 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]/P0001 ,
		_w5193_,
		_w5185_,
		_w5548_
	);
	LUT4 #(
		.INIT('h135f)
	) name2537 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]/P0001 ,
		_w5194_,
		_w5188_,
		_w5549_
	);
	LUT4 #(
		.INIT('h8000)
	) name2538 (
		_w5548_,
		_w5549_,
		_w5546_,
		_w5547_,
		_w5550_
	);
	LUT2 #(
		.INIT('h7)
	) name2539 (
		_w5545_,
		_w5550_,
		_w5551_
	);
	LUT3 #(
		.INIT('h6c)
	) name2540 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]/NET0131 ,
		\pci_target_unit_fifos_pciw_outTransactionCount_reg[0]/NET0131 ,
		_w4478_,
		_w5552_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2541 (
		\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]/P0001 ,
		_w3252_,
		_w3253_,
		_w3254_,
		_w5553_
	);
	LUT3 #(
		.INIT('h40)
	) name2542 (
		_w3081_,
		_w3097_,
		_w3104_,
		_w5554_
	);
	LUT2 #(
		.INIT('h6)
	) name2543 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		_w4478_,
		_w5555_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2544 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5556_
	);
	LUT4 #(
		.INIT('h2022)
	) name2545 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5557_
	);
	LUT2 #(
		.INIT('he)
	) name2546 (
		_w5556_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('heee0)
	) name2547 (
		_w3032_,
		_w3033_,
		_w5556_,
		_w5557_,
		_w5559_
	);
	LUT4 #(
		.INIT('h1011)
	) name2548 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5560_
	);
	LUT4 #(
		.INIT('h4544)
	) name2549 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5561_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2550 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5562_
	);
	LUT4 #(
		.INIT('h2022)
	) name2551 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w5563_
	);
	LUT4 #(
		.INIT('heee0)
	) name2552 (
		_w5560_,
		_w5561_,
		_w5562_,
		_w5563_,
		_w5564_
	);
	LUT3 #(
		.INIT('h80)
	) name2553 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]/P0001 ,
		_w5559_,
		_w5564_,
		_w5565_
	);
	LUT4 #(
		.INIT('h1110)
	) name2554 (
		_w3032_,
		_w3033_,
		_w5556_,
		_w5557_,
		_w5566_
	);
	LUT4 #(
		.INIT('h1110)
	) name2555 (
		_w5560_,
		_w5561_,
		_w5562_,
		_w5563_,
		_w5567_
	);
	LUT3 #(
		.INIT('h80)
	) name2556 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]/P0001 ,
		_w5566_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('h0001)
	) name2557 (
		_w5560_,
		_w5561_,
		_w5562_,
		_w5563_,
		_w5569_
	);
	LUT4 #(
		.INIT('h000e)
	) name2558 (
		_w3032_,
		_w3033_,
		_w5556_,
		_w5557_,
		_w5570_
	);
	LUT3 #(
		.INIT('h80)
	) name2559 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]/P0001 ,
		_w5569_,
		_w5570_,
		_w5571_
	);
	LUT4 #(
		.INIT('h0001)
	) name2560 (
		_w3032_,
		_w3033_,
		_w5556_,
		_w5557_,
		_w5572_
	);
	LUT3 #(
		.INIT('h80)
	) name2561 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]/P0001 ,
		_w5567_,
		_w5572_,
		_w5573_
	);
	LUT4 #(
		.INIT('h0001)
	) name2562 (
		_w5565_,
		_w5568_,
		_w5571_,
		_w5573_,
		_w5574_
	);
	LUT3 #(
		.INIT('h80)
	) name2563 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]/P0001 ,
		_w5569_,
		_w5566_,
		_w5575_
	);
	LUT4 #(
		.INIT('h000e)
	) name2564 (
		_w5560_,
		_w5561_,
		_w5562_,
		_w5563_,
		_w5576_
	);
	LUT3 #(
		.INIT('h80)
	) name2565 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]/P0001 ,
		_w5576_,
		_w5559_,
		_w5577_
	);
	LUT3 #(
		.INIT('h80)
	) name2566 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]/P0001 ,
		_w5570_,
		_w5564_,
		_w5578_
	);
	LUT3 #(
		.INIT('h80)
	) name2567 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]/P0001 ,
		_w5570_,
		_w5567_,
		_w5579_
	);
	LUT4 #(
		.INIT('h0001)
	) name2568 (
		_w5575_,
		_w5577_,
		_w5578_,
		_w5579_,
		_w5580_
	);
	LUT3 #(
		.INIT('h80)
	) name2569 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]/P0001 ,
		_w5566_,
		_w5564_,
		_w5581_
	);
	LUT3 #(
		.INIT('h80)
	) name2570 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]/P0001 ,
		_w5576_,
		_w5570_,
		_w5582_
	);
	LUT3 #(
		.INIT('h80)
	) name2571 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]/P0001 ,
		_w5576_,
		_w5572_,
		_w5583_
	);
	LUT3 #(
		.INIT('h80)
	) name2572 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]/P0001 ,
		_w5564_,
		_w5572_,
		_w5584_
	);
	LUT4 #(
		.INIT('h0001)
	) name2573 (
		_w5581_,
		_w5582_,
		_w5583_,
		_w5584_,
		_w5585_
	);
	LUT3 #(
		.INIT('h80)
	) name2574 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]/P0001 ,
		_w5566_,
		_w5576_,
		_w5586_
	);
	LUT3 #(
		.INIT('h80)
	) name2575 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]/P0001 ,
		_w5569_,
		_w5559_,
		_w5587_
	);
	LUT3 #(
		.INIT('h80)
	) name2576 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]/P0001 ,
		_w5569_,
		_w5572_,
		_w5588_
	);
	LUT3 #(
		.INIT('h80)
	) name2577 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]/P0001 ,
		_w5559_,
		_w5567_,
		_w5589_
	);
	LUT4 #(
		.INIT('h0001)
	) name2578 (
		_w5586_,
		_w5587_,
		_w5588_,
		_w5589_,
		_w5590_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2579 (
		_w5585_,
		_w5590_,
		_w5574_,
		_w5580_,
		_w5591_
	);
	LUT3 #(
		.INIT('h80)
	) name2580 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]/P0001 ,
		_w5564_,
		_w5572_,
		_w5592_
	);
	LUT3 #(
		.INIT('h80)
	) name2581 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]/P0001 ,
		_w5559_,
		_w5564_,
		_w5593_
	);
	LUT3 #(
		.INIT('h80)
	) name2582 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]/P0001 ,
		_w5570_,
		_w5564_,
		_w5594_
	);
	LUT3 #(
		.INIT('h80)
	) name2583 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]/P0001 ,
		_w5570_,
		_w5567_,
		_w5595_
	);
	LUT4 #(
		.INIT('h0001)
	) name2584 (
		_w5592_,
		_w5593_,
		_w5594_,
		_w5595_,
		_w5596_
	);
	LUT3 #(
		.INIT('h80)
	) name2585 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]/P0001 ,
		_w5566_,
		_w5576_,
		_w5597_
	);
	LUT3 #(
		.INIT('h80)
	) name2586 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]/P0001 ,
		_w5569_,
		_w5559_,
		_w5598_
	);
	LUT3 #(
		.INIT('h80)
	) name2587 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]/P0001 ,
		_w5569_,
		_w5572_,
		_w5599_
	);
	LUT3 #(
		.INIT('h80)
	) name2588 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]/P0001 ,
		_w5576_,
		_w5570_,
		_w5600_
	);
	LUT4 #(
		.INIT('h0001)
	) name2589 (
		_w5597_,
		_w5598_,
		_w5599_,
		_w5600_,
		_w5601_
	);
	LUT3 #(
		.INIT('h80)
	) name2590 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]/P0001 ,
		_w5576_,
		_w5572_,
		_w5602_
	);
	LUT3 #(
		.INIT('h80)
	) name2591 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]/P0001 ,
		_w5566_,
		_w5567_,
		_w5603_
	);
	LUT3 #(
		.INIT('h80)
	) name2592 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]/P0001 ,
		_w5569_,
		_w5570_,
		_w5604_
	);
	LUT3 #(
		.INIT('h80)
	) name2593 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]/P0001 ,
		_w5567_,
		_w5572_,
		_w5605_
	);
	LUT4 #(
		.INIT('h0001)
	) name2594 (
		_w5602_,
		_w5603_,
		_w5604_,
		_w5605_,
		_w5606_
	);
	LUT3 #(
		.INIT('h80)
	) name2595 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]/P0001 ,
		_w5569_,
		_w5566_,
		_w5607_
	);
	LUT3 #(
		.INIT('h80)
	) name2596 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]/P0001 ,
		_w5576_,
		_w5559_,
		_w5608_
	);
	LUT3 #(
		.INIT('h80)
	) name2597 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]/P0001 ,
		_w5559_,
		_w5567_,
		_w5609_
	);
	LUT3 #(
		.INIT('h80)
	) name2598 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]/P0001 ,
		_w5566_,
		_w5564_,
		_w5610_
	);
	LUT4 #(
		.INIT('h0001)
	) name2599 (
		_w5607_,
		_w5608_,
		_w5609_,
		_w5610_,
		_w5611_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2600 (
		_w5606_,
		_w5611_,
		_w5596_,
		_w5601_,
		_w5612_
	);
	LUT3 #(
		.INIT('h80)
	) name2601 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]/P0001 ,
		_w5564_,
		_w5572_,
		_w5613_
	);
	LUT3 #(
		.INIT('h80)
	) name2602 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]/P0001 ,
		_w5569_,
		_w5559_,
		_w5614_
	);
	LUT3 #(
		.INIT('h80)
	) name2603 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]/P0001 ,
		_w5570_,
		_w5564_,
		_w5615_
	);
	LUT3 #(
		.INIT('h80)
	) name2604 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]/P0001 ,
		_w5570_,
		_w5567_,
		_w5616_
	);
	LUT4 #(
		.INIT('h0001)
	) name2605 (
		_w5613_,
		_w5614_,
		_w5615_,
		_w5616_,
		_w5617_
	);
	LUT3 #(
		.INIT('h80)
	) name2606 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]/P0001 ,
		_w5569_,
		_w5570_,
		_w5618_
	);
	LUT3 #(
		.INIT('h80)
	) name2607 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]/P0001 ,
		_w5567_,
		_w5572_,
		_w5619_
	);
	LUT3 #(
		.INIT('h80)
	) name2608 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]/P0001 ,
		_w5566_,
		_w5564_,
		_w5620_
	);
	LUT3 #(
		.INIT('h80)
	) name2609 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]/P0001 ,
		_w5559_,
		_w5564_,
		_w5621_
	);
	LUT4 #(
		.INIT('h0001)
	) name2610 (
		_w5618_,
		_w5619_,
		_w5620_,
		_w5621_,
		_w5622_
	);
	LUT3 #(
		.INIT('h80)
	) name2611 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]/P0001 ,
		_w5576_,
		_w5572_,
		_w5623_
	);
	LUT3 #(
		.INIT('h80)
	) name2612 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]/P0001 ,
		_w5566_,
		_w5567_,
		_w5624_
	);
	LUT3 #(
		.INIT('h80)
	) name2613 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]/P0001 ,
		_w5569_,
		_w5572_,
		_w5625_
	);
	LUT3 #(
		.INIT('h80)
	) name2614 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]/P0001 ,
		_w5576_,
		_w5570_,
		_w5626_
	);
	LUT4 #(
		.INIT('h0001)
	) name2615 (
		_w5623_,
		_w5624_,
		_w5625_,
		_w5626_,
		_w5627_
	);
	LUT3 #(
		.INIT('h80)
	) name2616 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]/P0001 ,
		_w5569_,
		_w5566_,
		_w5628_
	);
	LUT3 #(
		.INIT('h80)
	) name2617 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]/P0001 ,
		_w5576_,
		_w5559_,
		_w5629_
	);
	LUT3 #(
		.INIT('h80)
	) name2618 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]/P0001 ,
		_w5559_,
		_w5567_,
		_w5630_
	);
	LUT3 #(
		.INIT('h80)
	) name2619 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]/P0001 ,
		_w5566_,
		_w5576_,
		_w5631_
	);
	LUT4 #(
		.INIT('h0001)
	) name2620 (
		_w5628_,
		_w5629_,
		_w5630_,
		_w5631_,
		_w5632_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2621 (
		_w5627_,
		_w5632_,
		_w5617_,
		_w5622_,
		_w5633_
	);
	LUT3 #(
		.INIT('h80)
	) name2622 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]/P0001 ,
		_w5576_,
		_w5570_,
		_w5634_
	);
	LUT3 #(
		.INIT('h80)
	) name2623 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]/P0001 ,
		_w5566_,
		_w5567_,
		_w5635_
	);
	LUT3 #(
		.INIT('h80)
	) name2624 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]/P0001 ,
		_w5569_,
		_w5570_,
		_w5636_
	);
	LUT3 #(
		.INIT('h80)
	) name2625 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]/P0001 ,
		_w5567_,
		_w5572_,
		_w5637_
	);
	LUT4 #(
		.INIT('h0001)
	) name2626 (
		_w5634_,
		_w5635_,
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT3 #(
		.INIT('h80)
	) name2627 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]/P0001 ,
		_w5576_,
		_w5572_,
		_w5639_
	);
	LUT3 #(
		.INIT('h80)
	) name2628 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]/P0001 ,
		_w5564_,
		_w5572_,
		_w5640_
	);
	LUT3 #(
		.INIT('h80)
	) name2629 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]/P0001 ,
		_w5569_,
		_w5566_,
		_w5641_
	);
	LUT3 #(
		.INIT('h80)
	) name2630 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]/P0001 ,
		_w5576_,
		_w5559_,
		_w5642_
	);
	LUT4 #(
		.INIT('h0001)
	) name2631 (
		_w5639_,
		_w5640_,
		_w5641_,
		_w5642_,
		_w5643_
	);
	LUT3 #(
		.INIT('h80)
	) name2632 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]/P0001 ,
		_w5569_,
		_w5572_,
		_w5644_
	);
	LUT3 #(
		.INIT('h80)
	) name2633 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]/P0001 ,
		_w5559_,
		_w5564_,
		_w5645_
	);
	LUT3 #(
		.INIT('h80)
	) name2634 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]/P0001 ,
		_w5570_,
		_w5564_,
		_w5646_
	);
	LUT3 #(
		.INIT('h80)
	) name2635 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]/P0001 ,
		_w5570_,
		_w5567_,
		_w5647_
	);
	LUT4 #(
		.INIT('h0001)
	) name2636 (
		_w5644_,
		_w5645_,
		_w5646_,
		_w5647_,
		_w5648_
	);
	LUT3 #(
		.INIT('h80)
	) name2637 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]/P0001 ,
		_w5566_,
		_w5576_,
		_w5649_
	);
	LUT3 #(
		.INIT('h80)
	) name2638 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]/P0001 ,
		_w5569_,
		_w5559_,
		_w5650_
	);
	LUT3 #(
		.INIT('h80)
	) name2639 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]/P0001 ,
		_w5566_,
		_w5564_,
		_w5651_
	);
	LUT3 #(
		.INIT('h80)
	) name2640 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]/P0001 ,
		_w5559_,
		_w5567_,
		_w5652_
	);
	LUT4 #(
		.INIT('h0001)
	) name2641 (
		_w5649_,
		_w5650_,
		_w5651_,
		_w5652_,
		_w5653_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2642 (
		_w5648_,
		_w5653_,
		_w5638_,
		_w5643_,
		_w5654_
	);
	LUT3 #(
		.INIT('h80)
	) name2643 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]/P0001 ,
		_w5564_,
		_w5572_,
		_w5655_
	);
	LUT3 #(
		.INIT('h80)
	) name2644 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]/P0001 ,
		_w5559_,
		_w5564_,
		_w5656_
	);
	LUT3 #(
		.INIT('h80)
	) name2645 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]/P0001 ,
		_w5559_,
		_w5567_,
		_w5657_
	);
	LUT3 #(
		.INIT('h80)
	) name2646 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]/P0001 ,
		_w5566_,
		_w5567_,
		_w5658_
	);
	LUT4 #(
		.INIT('h0001)
	) name2647 (
		_w5655_,
		_w5656_,
		_w5657_,
		_w5658_,
		_w5659_
	);
	LUT3 #(
		.INIT('h80)
	) name2648 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]/P0001 ,
		_w5566_,
		_w5576_,
		_w5660_
	);
	LUT3 #(
		.INIT('h80)
	) name2649 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]/P0001 ,
		_w5569_,
		_w5559_,
		_w5661_
	);
	LUT3 #(
		.INIT('h80)
	) name2650 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]/P0001 ,
		_w5569_,
		_w5572_,
		_w5662_
	);
	LUT3 #(
		.INIT('h80)
	) name2651 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]/P0001 ,
		_w5576_,
		_w5570_,
		_w5663_
	);
	LUT4 #(
		.INIT('h0001)
	) name2652 (
		_w5660_,
		_w5661_,
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT3 #(
		.INIT('h80)
	) name2653 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]/P0001 ,
		_w5576_,
		_w5572_,
		_w5665_
	);
	LUT3 #(
		.INIT('h80)
	) name2654 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]/P0001 ,
		_w5570_,
		_w5567_,
		_w5666_
	);
	LUT3 #(
		.INIT('h80)
	) name2655 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]/P0001 ,
		_w5569_,
		_w5570_,
		_w5667_
	);
	LUT3 #(
		.INIT('h80)
	) name2656 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]/P0001 ,
		_w5567_,
		_w5572_,
		_w5668_
	);
	LUT4 #(
		.INIT('h0001)
	) name2657 (
		_w5665_,
		_w5666_,
		_w5667_,
		_w5668_,
		_w5669_
	);
	LUT3 #(
		.INIT('h80)
	) name2658 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]/P0001 ,
		_w5569_,
		_w5566_,
		_w5670_
	);
	LUT3 #(
		.INIT('h80)
	) name2659 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]/P0001 ,
		_w5576_,
		_w5559_,
		_w5671_
	);
	LUT3 #(
		.INIT('h80)
	) name2660 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]/P0001 ,
		_w5570_,
		_w5564_,
		_w5672_
	);
	LUT3 #(
		.INIT('h80)
	) name2661 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]/P0001 ,
		_w5566_,
		_w5564_,
		_w5673_
	);
	LUT4 #(
		.INIT('h0001)
	) name2662 (
		_w5670_,
		_w5671_,
		_w5672_,
		_w5673_,
		_w5674_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2663 (
		_w5669_,
		_w5674_,
		_w5659_,
		_w5664_,
		_w5675_
	);
	LUT3 #(
		.INIT('h80)
	) name2664 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]/P0001 ,
		_w5570_,
		_w5567_,
		_w5676_
	);
	LUT3 #(
		.INIT('h80)
	) name2665 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]/P0001 ,
		_w5576_,
		_w5570_,
		_w5677_
	);
	LUT3 #(
		.INIT('h80)
	) name2666 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]/P0001 ,
		_w5576_,
		_w5572_,
		_w5678_
	);
	LUT3 #(
		.INIT('h80)
	) name2667 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]/P0001 ,
		_w5564_,
		_w5572_,
		_w5679_
	);
	LUT4 #(
		.INIT('h0001)
	) name2668 (
		_w5676_,
		_w5677_,
		_w5678_,
		_w5679_,
		_w5680_
	);
	LUT3 #(
		.INIT('h80)
	) name2669 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]/P0001 ,
		_w5569_,
		_w5570_,
		_w5681_
	);
	LUT3 #(
		.INIT('h80)
	) name2670 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]/P0001 ,
		_w5567_,
		_w5572_,
		_w5682_
	);
	LUT3 #(
		.INIT('h80)
	) name2671 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]/P0001 ,
		_w5566_,
		_w5564_,
		_w5683_
	);
	LUT3 #(
		.INIT('h80)
	) name2672 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]/P0001 ,
		_w5559_,
		_w5564_,
		_w5684_
	);
	LUT4 #(
		.INIT('h0001)
	) name2673 (
		_w5681_,
		_w5682_,
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT3 #(
		.INIT('h80)
	) name2674 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]/P0001 ,
		_w5570_,
		_w5564_,
		_w5686_
	);
	LUT3 #(
		.INIT('h80)
	) name2675 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]/P0001 ,
		_w5566_,
		_w5567_,
		_w5687_
	);
	LUT3 #(
		.INIT('h80)
	) name2676 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]/P0001 ,
		_w5566_,
		_w5576_,
		_w5688_
	);
	LUT3 #(
		.INIT('h80)
	) name2677 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]/P0001 ,
		_w5569_,
		_w5559_,
		_w5689_
	);
	LUT4 #(
		.INIT('h0001)
	) name2678 (
		_w5686_,
		_w5687_,
		_w5688_,
		_w5689_,
		_w5690_
	);
	LUT3 #(
		.INIT('h80)
	) name2679 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]/P0001 ,
		_w5569_,
		_w5566_,
		_w5691_
	);
	LUT3 #(
		.INIT('h80)
	) name2680 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]/P0001 ,
		_w5576_,
		_w5559_,
		_w5692_
	);
	LUT3 #(
		.INIT('h80)
	) name2681 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]/P0001 ,
		_w5559_,
		_w5567_,
		_w5693_
	);
	LUT3 #(
		.INIT('h80)
	) name2682 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]/P0001 ,
		_w5569_,
		_w5572_,
		_w5694_
	);
	LUT4 #(
		.INIT('h0001)
	) name2683 (
		_w5691_,
		_w5692_,
		_w5693_,
		_w5694_,
		_w5695_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2684 (
		_w5690_,
		_w5695_,
		_w5680_,
		_w5685_,
		_w5696_
	);
	LUT3 #(
		.INIT('h80)
	) name2685 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]/P0001 ,
		_w5576_,
		_w5559_,
		_w5697_
	);
	LUT3 #(
		.INIT('h80)
	) name2686 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]/P0001 ,
		_w5567_,
		_w5572_,
		_w5698_
	);
	LUT3 #(
		.INIT('h80)
	) name2687 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]/P0001 ,
		_w5559_,
		_w5567_,
		_w5699_
	);
	LUT3 #(
		.INIT('h80)
	) name2688 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]/P0001 ,
		_w5566_,
		_w5567_,
		_w5700_
	);
	LUT4 #(
		.INIT('h0001)
	) name2689 (
		_w5697_,
		_w5698_,
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT3 #(
		.INIT('h80)
	) name2690 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]/P0001 ,
		_w5569_,
		_w5572_,
		_w5702_
	);
	LUT3 #(
		.INIT('h80)
	) name2691 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]/P0001 ,
		_w5576_,
		_w5570_,
		_w5703_
	);
	LUT3 #(
		.INIT('h80)
	) name2692 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]/P0001 ,
		_w5566_,
		_w5564_,
		_w5704_
	);
	LUT3 #(
		.INIT('h80)
	) name2693 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]/P0001 ,
		_w5559_,
		_w5564_,
		_w5705_
	);
	LUT4 #(
		.INIT('h0001)
	) name2694 (
		_w5702_,
		_w5703_,
		_w5704_,
		_w5705_,
		_w5706_
	);
	LUT3 #(
		.INIT('h80)
	) name2695 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]/P0001 ,
		_w5569_,
		_w5566_,
		_w5707_
	);
	LUT3 #(
		.INIT('h80)
	) name2696 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]/P0001 ,
		_w5570_,
		_w5567_,
		_w5708_
	);
	LUT3 #(
		.INIT('h80)
	) name2697 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]/P0001 ,
		_w5566_,
		_w5576_,
		_w5709_
	);
	LUT3 #(
		.INIT('h80)
	) name2698 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]/P0001 ,
		_w5569_,
		_w5559_,
		_w5710_
	);
	LUT4 #(
		.INIT('h0001)
	) name2699 (
		_w5707_,
		_w5708_,
		_w5709_,
		_w5710_,
		_w5711_
	);
	LUT3 #(
		.INIT('h80)
	) name2700 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]/P0001 ,
		_w5576_,
		_w5572_,
		_w5712_
	);
	LUT3 #(
		.INIT('h80)
	) name2701 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]/P0001 ,
		_w5564_,
		_w5572_,
		_w5713_
	);
	LUT3 #(
		.INIT('h80)
	) name2702 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]/P0001 ,
		_w5570_,
		_w5564_,
		_w5714_
	);
	LUT3 #(
		.INIT('h80)
	) name2703 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]/P0001 ,
		_w5569_,
		_w5570_,
		_w5715_
	);
	LUT4 #(
		.INIT('h0001)
	) name2704 (
		_w5712_,
		_w5713_,
		_w5714_,
		_w5715_,
		_w5716_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2705 (
		_w5711_,
		_w5716_,
		_w5701_,
		_w5706_,
		_w5717_
	);
	LUT3 #(
		.INIT('h80)
	) name2706 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]/P0001 ,
		_w5559_,
		_w5564_,
		_w5718_
	);
	LUT3 #(
		.INIT('h80)
	) name2707 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]/P0001 ,
		_w5566_,
		_w5567_,
		_w5719_
	);
	LUT3 #(
		.INIT('h80)
	) name2708 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]/P0001 ,
		_w5569_,
		_w5570_,
		_w5720_
	);
	LUT3 #(
		.INIT('h80)
	) name2709 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]/P0001 ,
		_w5567_,
		_w5572_,
		_w5721_
	);
	LUT4 #(
		.INIT('h0001)
	) name2710 (
		_w5718_,
		_w5719_,
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT3 #(
		.INIT('h80)
	) name2711 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]/P0001 ,
		_w5569_,
		_w5566_,
		_w5723_
	);
	LUT3 #(
		.INIT('h80)
	) name2712 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]/P0001 ,
		_w5576_,
		_w5559_,
		_w5724_
	);
	LUT3 #(
		.INIT('h80)
	) name2713 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]/P0001 ,
		_w5570_,
		_w5564_,
		_w5725_
	);
	LUT3 #(
		.INIT('h80)
	) name2714 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]/P0001 ,
		_w5570_,
		_w5567_,
		_w5726_
	);
	LUT4 #(
		.INIT('h0001)
	) name2715 (
		_w5723_,
		_w5724_,
		_w5725_,
		_w5726_,
		_w5727_
	);
	LUT3 #(
		.INIT('h80)
	) name2716 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]/P0001 ,
		_w5566_,
		_w5564_,
		_w5728_
	);
	LUT3 #(
		.INIT('h80)
	) name2717 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]/P0001 ,
		_w5576_,
		_w5570_,
		_w5729_
	);
	LUT3 #(
		.INIT('h80)
	) name2718 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]/P0001 ,
		_w5576_,
		_w5572_,
		_w5730_
	);
	LUT3 #(
		.INIT('h80)
	) name2719 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]/P0001 ,
		_w5564_,
		_w5572_,
		_w5731_
	);
	LUT4 #(
		.INIT('h0001)
	) name2720 (
		_w5728_,
		_w5729_,
		_w5730_,
		_w5731_,
		_w5732_
	);
	LUT3 #(
		.INIT('h80)
	) name2721 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]/P0001 ,
		_w5566_,
		_w5576_,
		_w5733_
	);
	LUT3 #(
		.INIT('h80)
	) name2722 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]/P0001 ,
		_w5569_,
		_w5559_,
		_w5734_
	);
	LUT3 #(
		.INIT('h80)
	) name2723 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]/P0001 ,
		_w5569_,
		_w5572_,
		_w5735_
	);
	LUT3 #(
		.INIT('h80)
	) name2724 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]/P0001 ,
		_w5559_,
		_w5567_,
		_w5736_
	);
	LUT4 #(
		.INIT('h0001)
	) name2725 (
		_w5733_,
		_w5734_,
		_w5735_,
		_w5736_,
		_w5737_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2726 (
		_w5732_,
		_w5737_,
		_w5722_,
		_w5727_,
		_w5738_
	);
	LUT3 #(
		.INIT('h80)
	) name2727 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]/P0001 ,
		_w5569_,
		_w5559_,
		_w5739_
	);
	LUT3 #(
		.INIT('h80)
	) name2728 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]/P0001 ,
		_w5564_,
		_w5572_,
		_w5740_
	);
	LUT3 #(
		.INIT('h80)
	) name2729 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]/P0001 ,
		_w5569_,
		_w5570_,
		_w5741_
	);
	LUT3 #(
		.INIT('h80)
	) name2730 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]/P0001 ,
		_w5567_,
		_w5572_,
		_w5742_
	);
	LUT4 #(
		.INIT('h0001)
	) name2731 (
		_w5739_,
		_w5740_,
		_w5741_,
		_w5742_,
		_w5743_
	);
	LUT3 #(
		.INIT('h80)
	) name2732 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]/P0001 ,
		_w5569_,
		_w5566_,
		_w5744_
	);
	LUT3 #(
		.INIT('h80)
	) name2733 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]/P0001 ,
		_w5576_,
		_w5559_,
		_w5745_
	);
	LUT3 #(
		.INIT('h80)
	) name2734 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]/P0001 ,
		_w5570_,
		_w5564_,
		_w5746_
	);
	LUT3 #(
		.INIT('h80)
	) name2735 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]/P0001 ,
		_w5570_,
		_w5567_,
		_w5747_
	);
	LUT4 #(
		.INIT('h0001)
	) name2736 (
		_w5744_,
		_w5745_,
		_w5746_,
		_w5747_,
		_w5748_
	);
	LUT3 #(
		.INIT('h80)
	) name2737 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]/P0001 ,
		_w5566_,
		_w5576_,
		_w5749_
	);
	LUT3 #(
		.INIT('h80)
	) name2738 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]/P0001 ,
		_w5559_,
		_w5564_,
		_w5750_
	);
	LUT3 #(
		.INIT('h80)
	) name2739 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]/P0001 ,
		_w5559_,
		_w5567_,
		_w5751_
	);
	LUT3 #(
		.INIT('h80)
	) name2740 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]/P0001 ,
		_w5566_,
		_w5567_,
		_w5752_
	);
	LUT4 #(
		.INIT('h0001)
	) name2741 (
		_w5749_,
		_w5750_,
		_w5751_,
		_w5752_,
		_w5753_
	);
	LUT3 #(
		.INIT('h80)
	) name2742 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]/P0001 ,
		_w5569_,
		_w5572_,
		_w5754_
	);
	LUT3 #(
		.INIT('h80)
	) name2743 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]/P0001 ,
		_w5576_,
		_w5570_,
		_w5755_
	);
	LUT3 #(
		.INIT('h80)
	) name2744 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]/P0001 ,
		_w5566_,
		_w5564_,
		_w5756_
	);
	LUT3 #(
		.INIT('h80)
	) name2745 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]/P0001 ,
		_w5576_,
		_w5572_,
		_w5757_
	);
	LUT4 #(
		.INIT('h0001)
	) name2746 (
		_w5754_,
		_w5755_,
		_w5756_,
		_w5757_,
		_w5758_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2747 (
		_w5753_,
		_w5758_,
		_w5743_,
		_w5748_,
		_w5759_
	);
	LUT3 #(
		.INIT('h80)
	) name2748 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]/P0001 ,
		_w5570_,
		_w5567_,
		_w5760_
	);
	LUT3 #(
		.INIT('h80)
	) name2749 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]/P0001 ,
		_w5569_,
		_w5559_,
		_w5761_
	);
	LUT3 #(
		.INIT('h80)
	) name2750 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]/P0001 ,
		_w5569_,
		_w5566_,
		_w5762_
	);
	LUT3 #(
		.INIT('h80)
	) name2751 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]/P0001 ,
		_w5576_,
		_w5559_,
		_w5763_
	);
	LUT4 #(
		.INIT('h0001)
	) name2752 (
		_w5760_,
		_w5761_,
		_w5762_,
		_w5763_,
		_w5764_
	);
	LUT3 #(
		.INIT('h80)
	) name2753 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]/P0001 ,
		_w5566_,
		_w5564_,
		_w5765_
	);
	LUT3 #(
		.INIT('h80)
	) name2754 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]/P0001 ,
		_w5559_,
		_w5564_,
		_w5766_
	);
	LUT3 #(
		.INIT('h80)
	) name2755 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]/P0001 ,
		_w5569_,
		_w5570_,
		_w5767_
	);
	LUT3 #(
		.INIT('h80)
	) name2756 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]/P0001 ,
		_w5567_,
		_w5572_,
		_w5768_
	);
	LUT4 #(
		.INIT('h0001)
	) name2757 (
		_w5765_,
		_w5766_,
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT3 #(
		.INIT('h80)
	) name2758 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]/P0001 ,
		_w5570_,
		_w5564_,
		_w5770_
	);
	LUT3 #(
		.INIT('h80)
	) name2759 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]/P0001 ,
		_w5566_,
		_w5567_,
		_w5771_
	);
	LUT3 #(
		.INIT('h80)
	) name2760 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]/P0001 ,
		_w5569_,
		_w5572_,
		_w5772_
	);
	LUT3 #(
		.INIT('h80)
	) name2761 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]/P0001 ,
		_w5576_,
		_w5570_,
		_w5773_
	);
	LUT4 #(
		.INIT('h0001)
	) name2762 (
		_w5770_,
		_w5771_,
		_w5772_,
		_w5773_,
		_w5774_
	);
	LUT3 #(
		.INIT('h80)
	) name2763 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]/P0001 ,
		_w5576_,
		_w5572_,
		_w5775_
	);
	LUT3 #(
		.INIT('h80)
	) name2764 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]/P0001 ,
		_w5564_,
		_w5572_,
		_w5776_
	);
	LUT3 #(
		.INIT('h80)
	) name2765 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]/P0001 ,
		_w5559_,
		_w5567_,
		_w5777_
	);
	LUT3 #(
		.INIT('h80)
	) name2766 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]/P0001 ,
		_w5566_,
		_w5576_,
		_w5778_
	);
	LUT4 #(
		.INIT('h0001)
	) name2767 (
		_w5775_,
		_w5776_,
		_w5777_,
		_w5778_,
		_w5779_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2768 (
		_w5774_,
		_w5779_,
		_w5764_,
		_w5769_,
		_w5780_
	);
	LUT3 #(
		.INIT('h80)
	) name2769 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]/P0001 ,
		_w5576_,
		_w5570_,
		_w5781_
	);
	LUT3 #(
		.INIT('h80)
	) name2770 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]/P0001 ,
		_w5576_,
		_w5559_,
		_w5782_
	);
	LUT3 #(
		.INIT('h80)
	) name2771 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]/P0001 ,
		_w5566_,
		_w5564_,
		_w5783_
	);
	LUT3 #(
		.INIT('h80)
	) name2772 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]/P0001 ,
		_w5559_,
		_w5564_,
		_w5784_
	);
	LUT4 #(
		.INIT('h0001)
	) name2773 (
		_w5781_,
		_w5782_,
		_w5783_,
		_w5784_,
		_w5785_
	);
	LUT3 #(
		.INIT('h80)
	) name2774 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]/P0001 ,
		_w5559_,
		_w5567_,
		_w5786_
	);
	LUT3 #(
		.INIT('h80)
	) name2775 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]/P0001 ,
		_w5566_,
		_w5567_,
		_w5787_
	);
	LUT3 #(
		.INIT('h80)
	) name2776 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]/P0001 ,
		_w5576_,
		_w5572_,
		_w5788_
	);
	LUT3 #(
		.INIT('h80)
	) name2777 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]/P0001 ,
		_w5564_,
		_w5572_,
		_w5789_
	);
	LUT4 #(
		.INIT('h0001)
	) name2778 (
		_w5786_,
		_w5787_,
		_w5788_,
		_w5789_,
		_w5790_
	);
	LUT3 #(
		.INIT('h80)
	) name2779 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]/P0001 ,
		_w5569_,
		_w5572_,
		_w5791_
	);
	LUT3 #(
		.INIT('h80)
	) name2780 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]/P0001 ,
		_w5567_,
		_w5572_,
		_w5792_
	);
	LUT3 #(
		.INIT('h80)
	) name2781 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]/P0001 ,
		_w5570_,
		_w5564_,
		_w5793_
	);
	LUT3 #(
		.INIT('h80)
	) name2782 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]/P0001 ,
		_w5570_,
		_w5567_,
		_w5794_
	);
	LUT4 #(
		.INIT('h0001)
	) name2783 (
		_w5791_,
		_w5792_,
		_w5793_,
		_w5794_,
		_w5795_
	);
	LUT3 #(
		.INIT('h80)
	) name2784 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]/P0001 ,
		_w5566_,
		_w5576_,
		_w5796_
	);
	LUT3 #(
		.INIT('h80)
	) name2785 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]/P0001 ,
		_w5569_,
		_w5559_,
		_w5797_
	);
	LUT3 #(
		.INIT('h80)
	) name2786 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]/P0001 ,
		_w5569_,
		_w5570_,
		_w5798_
	);
	LUT3 #(
		.INIT('h80)
	) name2787 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]/P0001 ,
		_w5569_,
		_w5566_,
		_w5799_
	);
	LUT4 #(
		.INIT('h0001)
	) name2788 (
		_w5796_,
		_w5797_,
		_w5798_,
		_w5799_,
		_w5800_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2789 (
		_w5795_,
		_w5800_,
		_w5785_,
		_w5790_,
		_w5801_
	);
	LUT3 #(
		.INIT('h80)
	) name2790 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]/P0001 ,
		_w5576_,
		_w5559_,
		_w5802_
	);
	LUT3 #(
		.INIT('h80)
	) name2791 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]/P0001 ,
		_w5559_,
		_w5564_,
		_w5803_
	);
	LUT3 #(
		.INIT('h80)
	) name2792 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]/P0001 ,
		_w5559_,
		_w5567_,
		_w5804_
	);
	LUT3 #(
		.INIT('h80)
	) name2793 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]/P0001 ,
		_w5566_,
		_w5567_,
		_w5805_
	);
	LUT4 #(
		.INIT('h0001)
	) name2794 (
		_w5802_,
		_w5803_,
		_w5804_,
		_w5805_,
		_w5806_
	);
	LUT3 #(
		.INIT('h80)
	) name2795 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]/P0001 ,
		_w5566_,
		_w5576_,
		_w5807_
	);
	LUT3 #(
		.INIT('h80)
	) name2796 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]/P0001 ,
		_w5569_,
		_w5559_,
		_w5808_
	);
	LUT3 #(
		.INIT('h80)
	) name2797 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]/P0001 ,
		_w5569_,
		_w5572_,
		_w5809_
	);
	LUT3 #(
		.INIT('h80)
	) name2798 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]/P0001 ,
		_w5576_,
		_w5570_,
		_w5810_
	);
	LUT4 #(
		.INIT('h0001)
	) name2799 (
		_w5807_,
		_w5808_,
		_w5809_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h80)
	) name2800 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]/P0001 ,
		_w5569_,
		_w5566_,
		_w5812_
	);
	LUT3 #(
		.INIT('h80)
	) name2801 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]/P0001 ,
		_w5570_,
		_w5567_,
		_w5813_
	);
	LUT3 #(
		.INIT('h80)
	) name2802 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]/P0001 ,
		_w5569_,
		_w5570_,
		_w5814_
	);
	LUT3 #(
		.INIT('h80)
	) name2803 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]/P0001 ,
		_w5567_,
		_w5572_,
		_w5815_
	);
	LUT4 #(
		.INIT('h0001)
	) name2804 (
		_w5812_,
		_w5813_,
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT3 #(
		.INIT('h80)
	) name2805 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]/P0001 ,
		_w5576_,
		_w5572_,
		_w5817_
	);
	LUT3 #(
		.INIT('h80)
	) name2806 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]/P0001 ,
		_w5564_,
		_w5572_,
		_w5818_
	);
	LUT3 #(
		.INIT('h80)
	) name2807 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]/P0001 ,
		_w5570_,
		_w5564_,
		_w5819_
	);
	LUT3 #(
		.INIT('h80)
	) name2808 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]/P0001 ,
		_w5566_,
		_w5564_,
		_w5820_
	);
	LUT4 #(
		.INIT('h0001)
	) name2809 (
		_w5817_,
		_w5818_,
		_w5819_,
		_w5820_,
		_w5821_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2810 (
		_w5816_,
		_w5821_,
		_w5806_,
		_w5811_,
		_w5822_
	);
	LUT3 #(
		.INIT('h80)
	) name2811 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]/P0001 ,
		_w5567_,
		_w5572_,
		_w5823_
	);
	LUT3 #(
		.INIT('h80)
	) name2812 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]/P0001 ,
		_w5576_,
		_w5559_,
		_w5824_
	);
	LUT3 #(
		.INIT('h80)
	) name2813 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]/P0001 ,
		_w5566_,
		_w5564_,
		_w5825_
	);
	LUT3 #(
		.INIT('h80)
	) name2814 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]/P0001 ,
		_w5559_,
		_w5564_,
		_w5826_
	);
	LUT4 #(
		.INIT('h0001)
	) name2815 (
		_w5823_,
		_w5824_,
		_w5825_,
		_w5826_,
		_w5827_
	);
	LUT3 #(
		.INIT('h80)
	) name2816 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]/P0001 ,
		_w5576_,
		_w5572_,
		_w5828_
	);
	LUT3 #(
		.INIT('h80)
	) name2817 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]/P0001 ,
		_w5564_,
		_w5572_,
		_w5829_
	);
	LUT3 #(
		.INIT('h80)
	) name2818 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]/P0001 ,
		_w5570_,
		_w5564_,
		_w5830_
	);
	LUT3 #(
		.INIT('h80)
	) name2819 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]/P0001 ,
		_w5570_,
		_w5567_,
		_w5831_
	);
	LUT4 #(
		.INIT('h0001)
	) name2820 (
		_w5828_,
		_w5829_,
		_w5830_,
		_w5831_,
		_w5832_
	);
	LUT3 #(
		.INIT('h80)
	) name2821 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]/P0001 ,
		_w5569_,
		_w5570_,
		_w5833_
	);
	LUT3 #(
		.INIT('h80)
	) name2822 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]/P0001 ,
		_w5569_,
		_w5559_,
		_w5834_
	);
	LUT3 #(
		.INIT('h80)
	) name2823 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]/P0001 ,
		_w5559_,
		_w5567_,
		_w5835_
	);
	LUT3 #(
		.INIT('h80)
	) name2824 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]/P0001 ,
		_w5566_,
		_w5567_,
		_w5836_
	);
	LUT4 #(
		.INIT('h0001)
	) name2825 (
		_w5833_,
		_w5834_,
		_w5835_,
		_w5836_,
		_w5837_
	);
	LUT3 #(
		.INIT('h80)
	) name2826 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]/P0001 ,
		_w5569_,
		_w5572_,
		_w5838_
	);
	LUT3 #(
		.INIT('h80)
	) name2827 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]/P0001 ,
		_w5576_,
		_w5570_,
		_w5839_
	);
	LUT3 #(
		.INIT('h80)
	) name2828 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]/P0001 ,
		_w5566_,
		_w5576_,
		_w5840_
	);
	LUT3 #(
		.INIT('h80)
	) name2829 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]/P0001 ,
		_w5569_,
		_w5566_,
		_w5841_
	);
	LUT4 #(
		.INIT('h0001)
	) name2830 (
		_w5838_,
		_w5839_,
		_w5840_,
		_w5841_,
		_w5842_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2831 (
		_w5837_,
		_w5842_,
		_w5827_,
		_w5832_,
		_w5843_
	);
	LUT3 #(
		.INIT('h80)
	) name2832 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]/P0001 ,
		_w5564_,
		_w5572_,
		_w5844_
	);
	LUT3 #(
		.INIT('h80)
	) name2833 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]/P0001 ,
		_w5559_,
		_w5564_,
		_w5845_
	);
	LUT3 #(
		.INIT('h80)
	) name2834 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]/P0001 ,
		_w5570_,
		_w5564_,
		_w5846_
	);
	LUT3 #(
		.INIT('h80)
	) name2835 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]/P0001 ,
		_w5570_,
		_w5567_,
		_w5847_
	);
	LUT4 #(
		.INIT('h0001)
	) name2836 (
		_w5844_,
		_w5845_,
		_w5846_,
		_w5847_,
		_w5848_
	);
	LUT3 #(
		.INIT('h80)
	) name2837 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]/P0001 ,
		_w5569_,
		_w5572_,
		_w5849_
	);
	LUT3 #(
		.INIT('h80)
	) name2838 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]/P0001 ,
		_w5576_,
		_w5570_,
		_w5850_
	);
	LUT3 #(
		.INIT('h80)
	) name2839 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]/P0001 ,
		_w5569_,
		_w5570_,
		_w5851_
	);
	LUT3 #(
		.INIT('h80)
	) name2840 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]/P0001 ,
		_w5567_,
		_w5572_,
		_w5852_
	);
	LUT4 #(
		.INIT('h0001)
	) name2841 (
		_w5849_,
		_w5850_,
		_w5851_,
		_w5852_,
		_w5853_
	);
	LUT3 #(
		.INIT('h80)
	) name2842 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]/P0001 ,
		_w5576_,
		_w5572_,
		_w5854_
	);
	LUT3 #(
		.INIT('h80)
	) name2843 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]/P0001 ,
		_w5566_,
		_w5567_,
		_w5855_
	);
	LUT3 #(
		.INIT('h80)
	) name2844 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]/P0001 ,
		_w5566_,
		_w5576_,
		_w5856_
	);
	LUT3 #(
		.INIT('h80)
	) name2845 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]/P0001 ,
		_w5569_,
		_w5559_,
		_w5857_
	);
	LUT4 #(
		.INIT('h0001)
	) name2846 (
		_w5854_,
		_w5855_,
		_w5856_,
		_w5857_,
		_w5858_
	);
	LUT3 #(
		.INIT('h80)
	) name2847 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]/P0001 ,
		_w5569_,
		_w5566_,
		_w5859_
	);
	LUT3 #(
		.INIT('h80)
	) name2848 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]/P0001 ,
		_w5576_,
		_w5559_,
		_w5860_
	);
	LUT3 #(
		.INIT('h80)
	) name2849 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]/P0001 ,
		_w5559_,
		_w5567_,
		_w5861_
	);
	LUT3 #(
		.INIT('h80)
	) name2850 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]/P0001 ,
		_w5566_,
		_w5564_,
		_w5862_
	);
	LUT4 #(
		.INIT('h0001)
	) name2851 (
		_w5859_,
		_w5860_,
		_w5861_,
		_w5862_,
		_w5863_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2852 (
		_w5858_,
		_w5863_,
		_w5848_,
		_w5853_,
		_w5864_
	);
	LUT3 #(
		.INIT('h80)
	) name2853 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]/P0001 ,
		_w5564_,
		_w5572_,
		_w5865_
	);
	LUT3 #(
		.INIT('h80)
	) name2854 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]/P0001 ,
		_w5576_,
		_w5559_,
		_w5866_
	);
	LUT3 #(
		.INIT('h80)
	) name2855 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]/P0001 ,
		_w5570_,
		_w5564_,
		_w5867_
	);
	LUT3 #(
		.INIT('h80)
	) name2856 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]/P0001 ,
		_w5570_,
		_w5567_,
		_w5868_
	);
	LUT4 #(
		.INIT('h0001)
	) name2857 (
		_w5865_,
		_w5866_,
		_w5867_,
		_w5868_,
		_w5869_
	);
	LUT3 #(
		.INIT('h80)
	) name2858 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]/P0001 ,
		_w5569_,
		_w5572_,
		_w5870_
	);
	LUT3 #(
		.INIT('h80)
	) name2859 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]/P0001 ,
		_w5576_,
		_w5570_,
		_w5871_
	);
	LUT3 #(
		.INIT('h80)
	) name2860 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]/P0001 ,
		_w5569_,
		_w5570_,
		_w5872_
	);
	LUT3 #(
		.INIT('h80)
	) name2861 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]/P0001 ,
		_w5567_,
		_w5572_,
		_w5873_
	);
	LUT4 #(
		.INIT('h0001)
	) name2862 (
		_w5870_,
		_w5871_,
		_w5872_,
		_w5873_,
		_w5874_
	);
	LUT3 #(
		.INIT('h80)
	) name2863 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]/P0001 ,
		_w5576_,
		_w5572_,
		_w5875_
	);
	LUT3 #(
		.INIT('h80)
	) name2864 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]/P0001 ,
		_w5569_,
		_w5559_,
		_w5876_
	);
	LUT3 #(
		.INIT('h80)
	) name2865 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]/P0001 ,
		_w5566_,
		_w5564_,
		_w5877_
	);
	LUT3 #(
		.INIT('h80)
	) name2866 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]/P0001 ,
		_w5559_,
		_w5564_,
		_w5878_
	);
	LUT4 #(
		.INIT('h0001)
	) name2867 (
		_w5875_,
		_w5876_,
		_w5877_,
		_w5878_,
		_w5879_
	);
	LUT3 #(
		.INIT('h80)
	) name2868 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]/P0001 ,
		_w5559_,
		_w5567_,
		_w5880_
	);
	LUT3 #(
		.INIT('h80)
	) name2869 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]/P0001 ,
		_w5566_,
		_w5567_,
		_w5881_
	);
	LUT3 #(
		.INIT('h80)
	) name2870 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]/P0001 ,
		_w5566_,
		_w5576_,
		_w5882_
	);
	LUT3 #(
		.INIT('h80)
	) name2871 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]/P0001 ,
		_w5569_,
		_w5566_,
		_w5883_
	);
	LUT4 #(
		.INIT('h0001)
	) name2872 (
		_w5880_,
		_w5881_,
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2873 (
		_w5879_,
		_w5884_,
		_w5869_,
		_w5874_,
		_w5885_
	);
	LUT3 #(
		.INIT('h80)
	) name2874 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]/P0001 ,
		_w5567_,
		_w5572_,
		_w5886_
	);
	LUT3 #(
		.INIT('h80)
	) name2875 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]/P0001 ,
		_w5576_,
		_w5559_,
		_w5887_
	);
	LUT3 #(
		.INIT('h80)
	) name2876 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]/P0001 ,
		_w5566_,
		_w5576_,
		_w5888_
	);
	LUT3 #(
		.INIT('h80)
	) name2877 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]/P0001 ,
		_w5569_,
		_w5559_,
		_w5889_
	);
	LUT4 #(
		.INIT('h0001)
	) name2878 (
		_w5886_,
		_w5887_,
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT3 #(
		.INIT('h80)
	) name2879 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]/P0001 ,
		_w5570_,
		_w5564_,
		_w5891_
	);
	LUT3 #(
		.INIT('h80)
	) name2880 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]/P0001 ,
		_w5570_,
		_w5567_,
		_w5892_
	);
	LUT3 #(
		.INIT('h80)
	) name2881 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]/P0001 ,
		_w5576_,
		_w5572_,
		_w5893_
	);
	LUT3 #(
		.INIT('h80)
	) name2882 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]/P0001 ,
		_w5564_,
		_w5572_,
		_w5894_
	);
	LUT4 #(
		.INIT('h0001)
	) name2883 (
		_w5891_,
		_w5892_,
		_w5893_,
		_w5894_,
		_w5895_
	);
	LUT3 #(
		.INIT('h80)
	) name2884 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]/P0001 ,
		_w5569_,
		_w5570_,
		_w5896_
	);
	LUT3 #(
		.INIT('h80)
	) name2885 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]/P0001 ,
		_w5559_,
		_w5564_,
		_w5897_
	);
	LUT3 #(
		.INIT('h80)
	) name2886 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]/P0001 ,
		_w5559_,
		_w5567_,
		_w5898_
	);
	LUT3 #(
		.INIT('h80)
	) name2887 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]/P0001 ,
		_w5566_,
		_w5567_,
		_w5899_
	);
	LUT4 #(
		.INIT('h0001)
	) name2888 (
		_w5896_,
		_w5897_,
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT3 #(
		.INIT('h80)
	) name2889 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]/P0001 ,
		_w5569_,
		_w5572_,
		_w5901_
	);
	LUT3 #(
		.INIT('h80)
	) name2890 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]/P0001 ,
		_w5576_,
		_w5570_,
		_w5902_
	);
	LUT3 #(
		.INIT('h80)
	) name2891 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]/P0001 ,
		_w5566_,
		_w5564_,
		_w5903_
	);
	LUT3 #(
		.INIT('h80)
	) name2892 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]/P0001 ,
		_w5569_,
		_w5566_,
		_w5904_
	);
	LUT4 #(
		.INIT('h0001)
	) name2893 (
		_w5901_,
		_w5902_,
		_w5903_,
		_w5904_,
		_w5905_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2894 (
		_w5900_,
		_w5905_,
		_w5890_,
		_w5895_,
		_w5906_
	);
	LUT3 #(
		.INIT('h80)
	) name2895 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]/P0001 ,
		_w5570_,
		_w5567_,
		_w5907_
	);
	LUT3 #(
		.INIT('h80)
	) name2896 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]/P0001 ,
		_w5576_,
		_w5570_,
		_w5908_
	);
	LUT3 #(
		.INIT('h80)
	) name2897 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]/P0001 ,
		_w5576_,
		_w5572_,
		_w5909_
	);
	LUT3 #(
		.INIT('h80)
	) name2898 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]/P0001 ,
		_w5564_,
		_w5572_,
		_w5910_
	);
	LUT4 #(
		.INIT('h0001)
	) name2899 (
		_w5907_,
		_w5908_,
		_w5909_,
		_w5910_,
		_w5911_
	);
	LUT3 #(
		.INIT('h80)
	) name2900 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]/P0001 ,
		_w5566_,
		_w5576_,
		_w5912_
	);
	LUT3 #(
		.INIT('h80)
	) name2901 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]/P0001 ,
		_w5569_,
		_w5559_,
		_w5913_
	);
	LUT3 #(
		.INIT('h80)
	) name2902 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]/P0001 ,
		_w5569_,
		_w5570_,
		_w5914_
	);
	LUT3 #(
		.INIT('h80)
	) name2903 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]/P0001 ,
		_w5567_,
		_w5572_,
		_w5915_
	);
	LUT4 #(
		.INIT('h0001)
	) name2904 (
		_w5912_,
		_w5913_,
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT3 #(
		.INIT('h80)
	) name2905 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]/P0001 ,
		_w5570_,
		_w5564_,
		_w5917_
	);
	LUT3 #(
		.INIT('h80)
	) name2906 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]/P0001 ,
		_w5576_,
		_w5559_,
		_w5918_
	);
	LUT3 #(
		.INIT('h80)
	) name2907 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]/P0001 ,
		_w5566_,
		_w5564_,
		_w5919_
	);
	LUT3 #(
		.INIT('h80)
	) name2908 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]/P0001 ,
		_w5559_,
		_w5564_,
		_w5920_
	);
	LUT4 #(
		.INIT('h0001)
	) name2909 (
		_w5917_,
		_w5918_,
		_w5919_,
		_w5920_,
		_w5921_
	);
	LUT3 #(
		.INIT('h80)
	) name2910 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]/P0001 ,
		_w5559_,
		_w5567_,
		_w5922_
	);
	LUT3 #(
		.INIT('h80)
	) name2911 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]/P0001 ,
		_w5566_,
		_w5567_,
		_w5923_
	);
	LUT3 #(
		.INIT('h80)
	) name2912 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]/P0001 ,
		_w5569_,
		_w5566_,
		_w5924_
	);
	LUT3 #(
		.INIT('h80)
	) name2913 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]/P0001 ,
		_w5569_,
		_w5572_,
		_w5925_
	);
	LUT4 #(
		.INIT('h0001)
	) name2914 (
		_w5922_,
		_w5923_,
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2915 (
		_w5921_,
		_w5926_,
		_w5911_,
		_w5916_,
		_w5927_
	);
	LUT3 #(
		.INIT('h80)
	) name2916 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]/P0001 ,
		_w5564_,
		_w5572_,
		_w5928_
	);
	LUT3 #(
		.INIT('h80)
	) name2917 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]/P0001 ,
		_w5569_,
		_w5559_,
		_w5929_
	);
	LUT3 #(
		.INIT('h80)
	) name2918 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]/P0001 ,
		_w5569_,
		_w5566_,
		_w5930_
	);
	LUT3 #(
		.INIT('h80)
	) name2919 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]/P0001 ,
		_w5576_,
		_w5559_,
		_w5931_
	);
	LUT4 #(
		.INIT('h0001)
	) name2920 (
		_w5928_,
		_w5929_,
		_w5930_,
		_w5931_,
		_w5932_
	);
	LUT3 #(
		.INIT('h80)
	) name2921 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]/P0001 ,
		_w5566_,
		_w5564_,
		_w5933_
	);
	LUT3 #(
		.INIT('h80)
	) name2922 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]/P0001 ,
		_w5559_,
		_w5564_,
		_w5934_
	);
	LUT3 #(
		.INIT('h80)
	) name2923 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]/P0001 ,
		_w5569_,
		_w5570_,
		_w5935_
	);
	LUT3 #(
		.INIT('h80)
	) name2924 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]/P0001 ,
		_w5567_,
		_w5572_,
		_w5936_
	);
	LUT4 #(
		.INIT('h0001)
	) name2925 (
		_w5933_,
		_w5934_,
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT3 #(
		.INIT('h80)
	) name2926 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]/P0001 ,
		_w5576_,
		_w5572_,
		_w5938_
	);
	LUT3 #(
		.INIT('h80)
	) name2927 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]/P0001 ,
		_w5566_,
		_w5567_,
		_w5939_
	);
	LUT3 #(
		.INIT('h80)
	) name2928 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]/P0001 ,
		_w5569_,
		_w5572_,
		_w5940_
	);
	LUT3 #(
		.INIT('h80)
	) name2929 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]/P0001 ,
		_w5576_,
		_w5570_,
		_w5941_
	);
	LUT4 #(
		.INIT('h0001)
	) name2930 (
		_w5938_,
		_w5939_,
		_w5940_,
		_w5941_,
		_w5942_
	);
	LUT3 #(
		.INIT('h80)
	) name2931 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]/P0001 ,
		_w5570_,
		_w5564_,
		_w5943_
	);
	LUT3 #(
		.INIT('h80)
	) name2932 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]/P0001 ,
		_w5570_,
		_w5567_,
		_w5944_
	);
	LUT3 #(
		.INIT('h80)
	) name2933 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]/P0001 ,
		_w5559_,
		_w5567_,
		_w5945_
	);
	LUT3 #(
		.INIT('h80)
	) name2934 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]/P0001 ,
		_w5566_,
		_w5576_,
		_w5946_
	);
	LUT4 #(
		.INIT('h0001)
	) name2935 (
		_w5943_,
		_w5944_,
		_w5945_,
		_w5946_,
		_w5947_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2936 (
		_w5942_,
		_w5947_,
		_w5932_,
		_w5937_,
		_w5948_
	);
	LUT3 #(
		.INIT('h80)
	) name2937 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]/P0001 ,
		_w5576_,
		_w5559_,
		_w5949_
	);
	LUT3 #(
		.INIT('h80)
	) name2938 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]/P0001 ,
		_w5576_,
		_w5570_,
		_w5950_
	);
	LUT3 #(
		.INIT('h80)
	) name2939 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]/P0001 ,
		_w5570_,
		_w5564_,
		_w5951_
	);
	LUT3 #(
		.INIT('h80)
	) name2940 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]/P0001 ,
		_w5570_,
		_w5567_,
		_w5952_
	);
	LUT4 #(
		.INIT('h0001)
	) name2941 (
		_w5949_,
		_w5950_,
		_w5951_,
		_w5952_,
		_w5953_
	);
	LUT3 #(
		.INIT('h80)
	) name2942 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]/P0001 ,
		_w5566_,
		_w5576_,
		_w5954_
	);
	LUT3 #(
		.INIT('h80)
	) name2943 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]/P0001 ,
		_w5569_,
		_w5559_,
		_w5955_
	);
	LUT3 #(
		.INIT('h80)
	) name2944 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]/P0001 ,
		_w5569_,
		_w5570_,
		_w5956_
	);
	LUT3 #(
		.INIT('h80)
	) name2945 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]/P0001 ,
		_w5567_,
		_w5572_,
		_w5957_
	);
	LUT4 #(
		.INIT('h0001)
	) name2946 (
		_w5954_,
		_w5955_,
		_w5956_,
		_w5957_,
		_w5958_
	);
	LUT3 #(
		.INIT('h80)
	) name2947 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]/P0001 ,
		_w5569_,
		_w5566_,
		_w5959_
	);
	LUT3 #(
		.INIT('h80)
	) name2948 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]/P0001 ,
		_w5564_,
		_w5572_,
		_w5960_
	);
	LUT3 #(
		.INIT('h80)
	) name2949 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]/P0001 ,
		_w5566_,
		_w5564_,
		_w5961_
	);
	LUT3 #(
		.INIT('h80)
	) name2950 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]/P0001 ,
		_w5559_,
		_w5564_,
		_w5962_
	);
	LUT4 #(
		.INIT('h0001)
	) name2951 (
		_w5959_,
		_w5960_,
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT3 #(
		.INIT('h80)
	) name2952 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]/P0001 ,
		_w5559_,
		_w5567_,
		_w5964_
	);
	LUT3 #(
		.INIT('h80)
	) name2953 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]/P0001 ,
		_w5566_,
		_w5567_,
		_w5965_
	);
	LUT3 #(
		.INIT('h80)
	) name2954 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]/P0001 ,
		_w5576_,
		_w5572_,
		_w5966_
	);
	LUT3 #(
		.INIT('h80)
	) name2955 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]/P0001 ,
		_w5569_,
		_w5572_,
		_w5967_
	);
	LUT4 #(
		.INIT('h0001)
	) name2956 (
		_w5964_,
		_w5965_,
		_w5966_,
		_w5967_,
		_w5968_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2957 (
		_w5963_,
		_w5968_,
		_w5953_,
		_w5958_,
		_w5969_
	);
	LUT3 #(
		.INIT('h80)
	) name2958 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]/P0001 ,
		_w5566_,
		_w5567_,
		_w5970_
	);
	LUT3 #(
		.INIT('h80)
	) name2959 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]/P0001 ,
		_w5569_,
		_w5559_,
		_w5971_
	);
	LUT3 #(
		.INIT('h80)
	) name2960 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]/P0001 ,
		_w5569_,
		_w5566_,
		_w5972_
	);
	LUT3 #(
		.INIT('h80)
	) name2961 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]/P0001 ,
		_w5576_,
		_w5559_,
		_w5973_
	);
	LUT4 #(
		.INIT('h0001)
	) name2962 (
		_w5970_,
		_w5971_,
		_w5972_,
		_w5973_,
		_w5974_
	);
	LUT3 #(
		.INIT('h80)
	) name2963 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]/P0001 ,
		_w5569_,
		_w5570_,
		_w5975_
	);
	LUT3 #(
		.INIT('h80)
	) name2964 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]/P0001 ,
		_w5567_,
		_w5572_,
		_w5976_
	);
	LUT3 #(
		.INIT('h80)
	) name2965 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]/P0001 ,
		_w5566_,
		_w5564_,
		_w5977_
	);
	LUT3 #(
		.INIT('h80)
	) name2966 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]/P0001 ,
		_w5559_,
		_w5564_,
		_w5978_
	);
	LUT4 #(
		.INIT('h0001)
	) name2967 (
		_w5975_,
		_w5976_,
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT3 #(
		.INIT('h80)
	) name2968 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]/P0001 ,
		_w5559_,
		_w5567_,
		_w5980_
	);
	LUT3 #(
		.INIT('h80)
	) name2969 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]/P0001 ,
		_w5564_,
		_w5572_,
		_w5981_
	);
	LUT3 #(
		.INIT('h80)
	) name2970 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]/P0001 ,
		_w5569_,
		_w5572_,
		_w5982_
	);
	LUT3 #(
		.INIT('h80)
	) name2971 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]/P0001 ,
		_w5576_,
		_w5570_,
		_w5983_
	);
	LUT4 #(
		.INIT('h0001)
	) name2972 (
		_w5980_,
		_w5981_,
		_w5982_,
		_w5983_,
		_w5984_
	);
	LUT3 #(
		.INIT('h80)
	) name2973 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]/P0001 ,
		_w5570_,
		_w5564_,
		_w5985_
	);
	LUT3 #(
		.INIT('h80)
	) name2974 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]/P0001 ,
		_w5570_,
		_w5567_,
		_w5986_
	);
	LUT3 #(
		.INIT('h80)
	) name2975 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]/P0001 ,
		_w5576_,
		_w5572_,
		_w5987_
	);
	LUT3 #(
		.INIT('h80)
	) name2976 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]/P0001 ,
		_w5566_,
		_w5576_,
		_w5988_
	);
	LUT4 #(
		.INIT('h0001)
	) name2977 (
		_w5985_,
		_w5986_,
		_w5987_,
		_w5988_,
		_w5989_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2978 (
		_w5984_,
		_w5989_,
		_w5974_,
		_w5979_,
		_w5990_
	);
	LUT3 #(
		.INIT('h80)
	) name2979 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]/P0001 ,
		_w5567_,
		_w5572_,
		_w5991_
	);
	LUT3 #(
		.INIT('h80)
	) name2980 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]/P0001 ,
		_w5566_,
		_w5567_,
		_w5992_
	);
	LUT3 #(
		.INIT('h80)
	) name2981 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]/P0001 ,
		_w5569_,
		_w5572_,
		_w5993_
	);
	LUT3 #(
		.INIT('h80)
	) name2982 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]/P0001 ,
		_w5576_,
		_w5570_,
		_w5994_
	);
	LUT4 #(
		.INIT('h0001)
	) name2983 (
		_w5991_,
		_w5992_,
		_w5993_,
		_w5994_,
		_w5995_
	);
	LUT3 #(
		.INIT('h80)
	) name2984 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]/P0001 ,
		_w5570_,
		_w5564_,
		_w5996_
	);
	LUT3 #(
		.INIT('h80)
	) name2985 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]/P0001 ,
		_w5570_,
		_w5567_,
		_w5997_
	);
	LUT3 #(
		.INIT('h80)
	) name2986 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]/P0001 ,
		_w5576_,
		_w5572_,
		_w5998_
	);
	LUT3 #(
		.INIT('h80)
	) name2987 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]/P0001 ,
		_w5564_,
		_w5572_,
		_w5999_
	);
	LUT4 #(
		.INIT('h0001)
	) name2988 (
		_w5996_,
		_w5997_,
		_w5998_,
		_w5999_,
		_w6000_
	);
	LUT3 #(
		.INIT('h80)
	) name2989 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]/P0001 ,
		_w5569_,
		_w5570_,
		_w6001_
	);
	LUT3 #(
		.INIT('h80)
	) name2990 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]/P0001 ,
		_w5559_,
		_w5564_,
		_w6002_
	);
	LUT3 #(
		.INIT('h80)
	) name2991 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]/P0001 ,
		_w5569_,
		_w5566_,
		_w6003_
	);
	LUT3 #(
		.INIT('h80)
	) name2992 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]/P0001 ,
		_w5576_,
		_w5559_,
		_w6004_
	);
	LUT4 #(
		.INIT('h0001)
	) name2993 (
		_w6001_,
		_w6002_,
		_w6003_,
		_w6004_,
		_w6005_
	);
	LUT3 #(
		.INIT('h80)
	) name2994 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]/P0001 ,
		_w5566_,
		_w5576_,
		_w6006_
	);
	LUT3 #(
		.INIT('h80)
	) name2995 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]/P0001 ,
		_w5569_,
		_w5559_,
		_w6007_
	);
	LUT3 #(
		.INIT('h80)
	) name2996 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]/P0001 ,
		_w5566_,
		_w5564_,
		_w6008_
	);
	LUT3 #(
		.INIT('h80)
	) name2997 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]/P0001 ,
		_w5559_,
		_w5567_,
		_w6009_
	);
	LUT4 #(
		.INIT('h0001)
	) name2998 (
		_w6006_,
		_w6007_,
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2999 (
		_w6005_,
		_w6010_,
		_w5995_,
		_w6000_,
		_w6011_
	);
	LUT3 #(
		.INIT('h80)
	) name3000 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]/P0001 ,
		_w5559_,
		_w5564_,
		_w6012_
	);
	LUT3 #(
		.INIT('h80)
	) name3001 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]/P0001 ,
		_w5576_,
		_w5559_,
		_w6013_
	);
	LUT3 #(
		.INIT('h80)
	) name3002 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]/P0001 ,
		_w5569_,
		_w5572_,
		_w6014_
	);
	LUT3 #(
		.INIT('h80)
	) name3003 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]/P0001 ,
		_w5576_,
		_w5570_,
		_w6015_
	);
	LUT4 #(
		.INIT('h0001)
	) name3004 (
		_w6012_,
		_w6013_,
		_w6014_,
		_w6015_,
		_w6016_
	);
	LUT3 #(
		.INIT('h80)
	) name3005 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]/P0001 ,
		_w5576_,
		_w5572_,
		_w6017_
	);
	LUT3 #(
		.INIT('h80)
	) name3006 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]/P0001 ,
		_w5564_,
		_w5572_,
		_w6018_
	);
	LUT3 #(
		.INIT('h80)
	) name3007 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]/P0001 ,
		_w5570_,
		_w5564_,
		_w6019_
	);
	LUT3 #(
		.INIT('h80)
	) name3008 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]/P0001 ,
		_w5570_,
		_w5567_,
		_w6020_
	);
	LUT4 #(
		.INIT('h0001)
	) name3009 (
		_w6017_,
		_w6018_,
		_w6019_,
		_w6020_,
		_w6021_
	);
	LUT3 #(
		.INIT('h80)
	) name3010 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]/P0001 ,
		_w5566_,
		_w5564_,
		_w6022_
	);
	LUT3 #(
		.INIT('h80)
	) name3011 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]/P0001 ,
		_w5567_,
		_w5572_,
		_w6023_
	);
	LUT3 #(
		.INIT('h80)
	) name3012 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]/P0001 ,
		_w5559_,
		_w5567_,
		_w6024_
	);
	LUT3 #(
		.INIT('h80)
	) name3013 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]/P0001 ,
		_w5566_,
		_w5567_,
		_w6025_
	);
	LUT4 #(
		.INIT('h0001)
	) name3014 (
		_w6022_,
		_w6023_,
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT3 #(
		.INIT('h80)
	) name3015 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]/P0001 ,
		_w5566_,
		_w5576_,
		_w6027_
	);
	LUT3 #(
		.INIT('h80)
	) name3016 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]/P0001 ,
		_w5569_,
		_w5559_,
		_w6028_
	);
	LUT3 #(
		.INIT('h80)
	) name3017 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]/P0001 ,
		_w5569_,
		_w5570_,
		_w6029_
	);
	LUT3 #(
		.INIT('h80)
	) name3018 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]/P0001 ,
		_w5569_,
		_w5566_,
		_w6030_
	);
	LUT4 #(
		.INIT('h0001)
	) name3019 (
		_w6027_,
		_w6028_,
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3020 (
		_w6026_,
		_w6031_,
		_w6016_,
		_w6021_,
		_w6032_
	);
	LUT3 #(
		.INIT('h80)
	) name3021 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]/P0001 ,
		_w5576_,
		_w5559_,
		_w6033_
	);
	LUT3 #(
		.INIT('h80)
	) name3022 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]/P0001 ,
		_w5567_,
		_w5572_,
		_w6034_
	);
	LUT3 #(
		.INIT('h80)
	) name3023 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]/P0001 ,
		_w5570_,
		_w5564_,
		_w6035_
	);
	LUT3 #(
		.INIT('h80)
	) name3024 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]/P0001 ,
		_w5570_,
		_w5567_,
		_w6036_
	);
	LUT4 #(
		.INIT('h0001)
	) name3025 (
		_w6033_,
		_w6034_,
		_w6035_,
		_w6036_,
		_w6037_
	);
	LUT3 #(
		.INIT('h80)
	) name3026 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]/P0001 ,
		_w5569_,
		_w5572_,
		_w6038_
	);
	LUT3 #(
		.INIT('h80)
	) name3027 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]/P0001 ,
		_w5576_,
		_w5570_,
		_w6039_
	);
	LUT3 #(
		.INIT('h80)
	) name3028 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]/P0001 ,
		_w5566_,
		_w5564_,
		_w6040_
	);
	LUT3 #(
		.INIT('h80)
	) name3029 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]/P0001 ,
		_w5559_,
		_w5564_,
		_w6041_
	);
	LUT4 #(
		.INIT('h0001)
	) name3030 (
		_w6038_,
		_w6039_,
		_w6040_,
		_w6041_,
		_w6042_
	);
	LUT3 #(
		.INIT('h80)
	) name3031 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]/P0001 ,
		_w5569_,
		_w5566_,
		_w6043_
	);
	LUT3 #(
		.INIT('h80)
	) name3032 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]/P0001 ,
		_w5564_,
		_w5572_,
		_w6044_
	);
	LUT3 #(
		.INIT('h80)
	) name3033 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]/P0001 ,
		_w5566_,
		_w5576_,
		_w6045_
	);
	LUT3 #(
		.INIT('h80)
	) name3034 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]/P0001 ,
		_w5569_,
		_w5559_,
		_w6046_
	);
	LUT4 #(
		.INIT('h0001)
	) name3035 (
		_w6043_,
		_w6044_,
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT3 #(
		.INIT('h80)
	) name3036 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]/P0001 ,
		_w5559_,
		_w5567_,
		_w6048_
	);
	LUT3 #(
		.INIT('h80)
	) name3037 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]/P0001 ,
		_w5566_,
		_w5567_,
		_w6049_
	);
	LUT3 #(
		.INIT('h80)
	) name3038 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]/P0001 ,
		_w5576_,
		_w5572_,
		_w6050_
	);
	LUT3 #(
		.INIT('h80)
	) name3039 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]/P0001 ,
		_w5569_,
		_w5570_,
		_w6051_
	);
	LUT4 #(
		.INIT('h0001)
	) name3040 (
		_w6048_,
		_w6049_,
		_w6050_,
		_w6051_,
		_w6052_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3041 (
		_w6047_,
		_w6052_,
		_w6037_,
		_w6042_,
		_w6053_
	);
	LUT3 #(
		.INIT('h80)
	) name3042 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]/P0001 ,
		_w5576_,
		_w5570_,
		_w6054_
	);
	LUT3 #(
		.INIT('h80)
	) name3043 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]/P0001 ,
		_w5564_,
		_w5572_,
		_w6055_
	);
	LUT3 #(
		.INIT('h80)
	) name3044 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]/P0001 ,
		_w5566_,
		_w5576_,
		_w6056_
	);
	LUT3 #(
		.INIT('h80)
	) name3045 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]/P0001 ,
		_w5569_,
		_w5559_,
		_w6057_
	);
	LUT4 #(
		.INIT('h0001)
	) name3046 (
		_w6054_,
		_w6055_,
		_w6056_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('h80)
	) name3047 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]/P0001 ,
		_w5559_,
		_w5567_,
		_w6059_
	);
	LUT3 #(
		.INIT('h80)
	) name3048 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]/P0001 ,
		_w5566_,
		_w5567_,
		_w6060_
	);
	LUT3 #(
		.INIT('h80)
	) name3049 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]/P0001 ,
		_w5570_,
		_w5564_,
		_w6061_
	);
	LUT3 #(
		.INIT('h80)
	) name3050 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]/P0001 ,
		_w5570_,
		_w5567_,
		_w6062_
	);
	LUT4 #(
		.INIT('h0001)
	) name3051 (
		_w6059_,
		_w6060_,
		_w6061_,
		_w6062_,
		_w6063_
	);
	LUT3 #(
		.INIT('h80)
	) name3052 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]/P0001 ,
		_w5569_,
		_w5572_,
		_w6064_
	);
	LUT3 #(
		.INIT('h80)
	) name3053 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]/P0001 ,
		_w5559_,
		_w5564_,
		_w6065_
	);
	LUT3 #(
		.INIT('h80)
	) name3054 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]/P0001 ,
		_w5569_,
		_w5566_,
		_w6066_
	);
	LUT3 #(
		.INIT('h80)
	) name3055 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]/P0001 ,
		_w5576_,
		_w5559_,
		_w6067_
	);
	LUT4 #(
		.INIT('h0001)
	) name3056 (
		_w6064_,
		_w6065_,
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT3 #(
		.INIT('h80)
	) name3057 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]/P0001 ,
		_w5569_,
		_w5570_,
		_w6069_
	);
	LUT3 #(
		.INIT('h80)
	) name3058 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]/P0001 ,
		_w5567_,
		_w5572_,
		_w6070_
	);
	LUT3 #(
		.INIT('h80)
	) name3059 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]/P0001 ,
		_w5566_,
		_w5564_,
		_w6071_
	);
	LUT3 #(
		.INIT('h80)
	) name3060 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]/P0001 ,
		_w5576_,
		_w5572_,
		_w6072_
	);
	LUT4 #(
		.INIT('h0001)
	) name3061 (
		_w6069_,
		_w6070_,
		_w6071_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3062 (
		_w6068_,
		_w6073_,
		_w6058_,
		_w6063_,
		_w6074_
	);
	LUT3 #(
		.INIT('h80)
	) name3063 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]/P0001 ,
		_w5566_,
		_w5567_,
		_w6075_
	);
	LUT3 #(
		.INIT('h80)
	) name3064 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]/P0001 ,
		_w5569_,
		_w5559_,
		_w6076_
	);
	LUT3 #(
		.INIT('h80)
	) name3065 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]/P0001 ,
		_w5569_,
		_w5566_,
		_w6077_
	);
	LUT3 #(
		.INIT('h80)
	) name3066 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]/P0001 ,
		_w5576_,
		_w5559_,
		_w6078_
	);
	LUT4 #(
		.INIT('h0001)
	) name3067 (
		_w6075_,
		_w6076_,
		_w6077_,
		_w6078_,
		_w6079_
	);
	LUT3 #(
		.INIT('h80)
	) name3068 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]/P0001 ,
		_w5569_,
		_w5570_,
		_w6080_
	);
	LUT3 #(
		.INIT('h80)
	) name3069 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]/P0001 ,
		_w5567_,
		_w5572_,
		_w6081_
	);
	LUT3 #(
		.INIT('h80)
	) name3070 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]/P0001 ,
		_w5566_,
		_w5564_,
		_w6082_
	);
	LUT3 #(
		.INIT('h80)
	) name3071 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]/P0001 ,
		_w5559_,
		_w5564_,
		_w6083_
	);
	LUT4 #(
		.INIT('h0001)
	) name3072 (
		_w6080_,
		_w6081_,
		_w6082_,
		_w6083_,
		_w6084_
	);
	LUT3 #(
		.INIT('h80)
	) name3073 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]/P0001 ,
		_w5559_,
		_w5567_,
		_w6085_
	);
	LUT3 #(
		.INIT('h80)
	) name3074 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]/P0001 ,
		_w5570_,
		_w5567_,
		_w6086_
	);
	LUT3 #(
		.INIT('h80)
	) name3075 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]/P0001 ,
		_w5569_,
		_w5572_,
		_w6087_
	);
	LUT3 #(
		.INIT('h80)
	) name3076 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]/P0001 ,
		_w5576_,
		_w5570_,
		_w6088_
	);
	LUT4 #(
		.INIT('h0001)
	) name3077 (
		_w6085_,
		_w6086_,
		_w6087_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h80)
	) name3078 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]/P0001 ,
		_w5576_,
		_w5572_,
		_w6090_
	);
	LUT3 #(
		.INIT('h80)
	) name3079 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]/P0001 ,
		_w5564_,
		_w5572_,
		_w6091_
	);
	LUT3 #(
		.INIT('h80)
	) name3080 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]/P0001 ,
		_w5570_,
		_w5564_,
		_w6092_
	);
	LUT3 #(
		.INIT('h80)
	) name3081 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]/P0001 ,
		_w5566_,
		_w5576_,
		_w6093_
	);
	LUT4 #(
		.INIT('h0001)
	) name3082 (
		_w6090_,
		_w6091_,
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3083 (
		_w6089_,
		_w6094_,
		_w6079_,
		_w6084_,
		_w6095_
	);
	LUT3 #(
		.INIT('h80)
	) name3084 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]/P0001 ,
		_w5559_,
		_w5564_,
		_w6096_
	);
	LUT3 #(
		.INIT('h80)
	) name3085 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]/P0001 ,
		_w5566_,
		_w5567_,
		_w6097_
	);
	LUT3 #(
		.INIT('h80)
	) name3086 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]/P0001 ,
		_w5569_,
		_w5570_,
		_w6098_
	);
	LUT3 #(
		.INIT('h80)
	) name3087 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]/P0001 ,
		_w5567_,
		_w5572_,
		_w6099_
	);
	LUT4 #(
		.INIT('h0001)
	) name3088 (
		_w6096_,
		_w6097_,
		_w6098_,
		_w6099_,
		_w6100_
	);
	LUT3 #(
		.INIT('h80)
	) name3089 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]/P0001 ,
		_w5576_,
		_w5572_,
		_w6101_
	);
	LUT3 #(
		.INIT('h80)
	) name3090 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]/P0001 ,
		_w5564_,
		_w5572_,
		_w6102_
	);
	LUT3 #(
		.INIT('h80)
	) name3091 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]/P0001 ,
		_w5569_,
		_w5566_,
		_w6103_
	);
	LUT3 #(
		.INIT('h80)
	) name3092 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]/P0001 ,
		_w5576_,
		_w5559_,
		_w6104_
	);
	LUT4 #(
		.INIT('h0001)
	) name3093 (
		_w6101_,
		_w6102_,
		_w6103_,
		_w6104_,
		_w6105_
	);
	LUT3 #(
		.INIT('h80)
	) name3094 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]/P0001 ,
		_w5566_,
		_w5564_,
		_w6106_
	);
	LUT3 #(
		.INIT('h80)
	) name3095 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]/P0001 ,
		_w5576_,
		_w5570_,
		_w6107_
	);
	LUT3 #(
		.INIT('h80)
	) name3096 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]/P0001 ,
		_w5570_,
		_w5564_,
		_w6108_
	);
	LUT3 #(
		.INIT('h80)
	) name3097 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]/P0001 ,
		_w5570_,
		_w5567_,
		_w6109_
	);
	LUT4 #(
		.INIT('h0001)
	) name3098 (
		_w6106_,
		_w6107_,
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT3 #(
		.INIT('h80)
	) name3099 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]/P0001 ,
		_w5566_,
		_w5576_,
		_w6111_
	);
	LUT3 #(
		.INIT('h80)
	) name3100 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]/P0001 ,
		_w5569_,
		_w5559_,
		_w6112_
	);
	LUT3 #(
		.INIT('h80)
	) name3101 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]/P0001 ,
		_w5569_,
		_w5572_,
		_w6113_
	);
	LUT3 #(
		.INIT('h80)
	) name3102 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]/P0001 ,
		_w5559_,
		_w5567_,
		_w6114_
	);
	LUT4 #(
		.INIT('h0001)
	) name3103 (
		_w6111_,
		_w6112_,
		_w6113_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3104 (
		_w6110_,
		_w6115_,
		_w6100_,
		_w6105_,
		_w6116_
	);
	LUT3 #(
		.INIT('h80)
	) name3105 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]/P0001 ,
		_w5559_,
		_w5567_,
		_w6117_
	);
	LUT3 #(
		.INIT('h80)
	) name3106 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]/P0001 ,
		_w5566_,
		_w5567_,
		_w6118_
	);
	LUT3 #(
		.INIT('h80)
	) name3107 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001 ,
		_w5567_,
		_w5572_,
		_w6119_
	);
	LUT3 #(
		.INIT('h80)
	) name3108 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001 ,
		_w5569_,
		_w5566_,
		_w6120_
	);
	LUT4 #(
		.INIT('h0001)
	) name3109 (
		_w6117_,
		_w6118_,
		_w6119_,
		_w6120_,
		_w6121_
	);
	LUT3 #(
		.INIT('h80)
	) name3110 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001 ,
		_w5570_,
		_w5564_,
		_w6122_
	);
	LUT3 #(
		.INIT('h80)
	) name3111 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001 ,
		_w5576_,
		_w5570_,
		_w6123_
	);
	LUT3 #(
		.INIT('h80)
	) name3112 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001 ,
		_w5564_,
		_w5572_,
		_w6124_
	);
	LUT3 #(
		.INIT('h80)
	) name3113 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001 ,
		_w5566_,
		_w5564_,
		_w6125_
	);
	LUT4 #(
		.INIT('h0001)
	) name3114 (
		_w6122_,
		_w6123_,
		_w6124_,
		_w6125_,
		_w6126_
	);
	LUT3 #(
		.INIT('h80)
	) name3115 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]/P0001 ,
		_w5569_,
		_w5559_,
		_w6127_
	);
	LUT3 #(
		.INIT('h80)
	) name3116 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]/P0001 ,
		_w5570_,
		_w5567_,
		_w6128_
	);
	LUT3 #(
		.INIT('h80)
	) name3117 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001 ,
		_w5569_,
		_w5570_,
		_w6129_
	);
	LUT3 #(
		.INIT('h80)
	) name3118 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]/P0001 ,
		_w5559_,
		_w5564_,
		_w6130_
	);
	LUT4 #(
		.INIT('h0001)
	) name3119 (
		_w6127_,
		_w6128_,
		_w6129_,
		_w6130_,
		_w6131_
	);
	LUT3 #(
		.INIT('h80)
	) name3120 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001 ,
		_w5566_,
		_w5576_,
		_w6132_
	);
	LUT3 #(
		.INIT('h80)
	) name3121 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001 ,
		_w5576_,
		_w5572_,
		_w6133_
	);
	LUT3 #(
		.INIT('h80)
	) name3122 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001 ,
		_w5576_,
		_w5559_,
		_w6134_
	);
	LUT3 #(
		.INIT('h80)
	) name3123 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001 ,
		_w5569_,
		_w5572_,
		_w6135_
	);
	LUT4 #(
		.INIT('h0001)
	) name3124 (
		_w6132_,
		_w6133_,
		_w6134_,
		_w6135_,
		_w6136_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3125 (
		_w6131_,
		_w6136_,
		_w6121_,
		_w6126_,
		_w6137_
	);
	LUT3 #(
		.INIT('h80)
	) name3126 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001 ,
		_w5566_,
		_w5576_,
		_w6138_
	);
	LUT3 #(
		.INIT('h80)
	) name3127 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001 ,
		_w5566_,
		_w5567_,
		_w6139_
	);
	LUT3 #(
		.INIT('h80)
	) name3128 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001 ,
		_w5569_,
		_w5570_,
		_w6140_
	);
	LUT3 #(
		.INIT('h80)
	) name3129 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001 ,
		_w5566_,
		_w5564_,
		_w6141_
	);
	LUT4 #(
		.INIT('h0001)
	) name3130 (
		_w6138_,
		_w6139_,
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT3 #(
		.INIT('h80)
	) name3131 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001 ,
		_w5570_,
		_w5567_,
		_w6143_
	);
	LUT3 #(
		.INIT('h80)
	) name3132 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001 ,
		_w5576_,
		_w5570_,
		_w6144_
	);
	LUT3 #(
		.INIT('h80)
	) name3133 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001 ,
		_w5576_,
		_w5572_,
		_w6145_
	);
	LUT3 #(
		.INIT('h80)
	) name3134 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001 ,
		_w5570_,
		_w5564_,
		_w6146_
	);
	LUT4 #(
		.INIT('h0001)
	) name3135 (
		_w6143_,
		_w6144_,
		_w6145_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h80)
	) name3136 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001 ,
		_w5569_,
		_w5566_,
		_w6148_
	);
	LUT3 #(
		.INIT('h80)
	) name3137 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001 ,
		_w5559_,
		_w5567_,
		_w6149_
	);
	LUT3 #(
		.INIT('h80)
	) name3138 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001 ,
		_w5576_,
		_w5559_,
		_w6150_
	);
	LUT3 #(
		.INIT('h80)
	) name3139 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001 ,
		_w5567_,
		_w5572_,
		_w6151_
	);
	LUT4 #(
		.INIT('h0001)
	) name3140 (
		_w6148_,
		_w6149_,
		_w6150_,
		_w6151_,
		_w6152_
	);
	LUT3 #(
		.INIT('h80)
	) name3141 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001 ,
		_w5569_,
		_w5572_,
		_w6153_
	);
	LUT3 #(
		.INIT('h80)
	) name3142 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001 ,
		_w5569_,
		_w5559_,
		_w6154_
	);
	LUT3 #(
		.INIT('h80)
	) name3143 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001 ,
		_w5564_,
		_w5572_,
		_w6155_
	);
	LUT3 #(
		.INIT('h80)
	) name3144 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001 ,
		_w5559_,
		_w5564_,
		_w6156_
	);
	LUT4 #(
		.INIT('h0001)
	) name3145 (
		_w6153_,
		_w6154_,
		_w6155_,
		_w6156_,
		_w6157_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3146 (
		_w6152_,
		_w6157_,
		_w6142_,
		_w6147_,
		_w6158_
	);
	LUT3 #(
		.INIT('h80)
	) name3147 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]/P0001 ,
		_w5569_,
		_w5559_,
		_w6159_
	);
	LUT3 #(
		.INIT('h80)
	) name3148 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]/P0001 ,
		_w5570_,
		_w5567_,
		_w6160_
	);
	LUT3 #(
		.INIT('h80)
	) name3149 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]/P0001 ,
		_w5569_,
		_w5572_,
		_w6161_
	);
	LUT3 #(
		.INIT('h80)
	) name3150 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]/P0001 ,
		_w5576_,
		_w5570_,
		_w6162_
	);
	LUT4 #(
		.INIT('h0001)
	) name3151 (
		_w6159_,
		_w6160_,
		_w6161_,
		_w6162_,
		_w6163_
	);
	LUT3 #(
		.INIT('h80)
	) name3152 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]/P0001 ,
		_w5569_,
		_w5566_,
		_w6164_
	);
	LUT3 #(
		.INIT('h80)
	) name3153 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]/P0001 ,
		_w5576_,
		_w5559_,
		_w6165_
	);
	LUT3 #(
		.INIT('h80)
	) name3154 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]/P0001 ,
		_w5576_,
		_w5572_,
		_w6166_
	);
	LUT3 #(
		.INIT('h80)
	) name3155 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]/P0001 ,
		_w5564_,
		_w5572_,
		_w6167_
	);
	LUT4 #(
		.INIT('h0001)
	) name3156 (
		_w6164_,
		_w6165_,
		_w6166_,
		_w6167_,
		_w6168_
	);
	LUT3 #(
		.INIT('h80)
	) name3157 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]/P0001 ,
		_w5566_,
		_w5576_,
		_w6169_
	);
	LUT3 #(
		.INIT('h80)
	) name3158 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]/P0001 ,
		_w5559_,
		_w5564_,
		_w6170_
	);
	LUT3 #(
		.INIT('h80)
	) name3159 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]/P0001 ,
		_w5559_,
		_w5567_,
		_w6171_
	);
	LUT3 #(
		.INIT('h80)
	) name3160 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]/P0001 ,
		_w5566_,
		_w5567_,
		_w6172_
	);
	LUT4 #(
		.INIT('h0001)
	) name3161 (
		_w6169_,
		_w6170_,
		_w6171_,
		_w6172_,
		_w6173_
	);
	LUT3 #(
		.INIT('h80)
	) name3162 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]/P0001 ,
		_w5569_,
		_w5570_,
		_w6174_
	);
	LUT3 #(
		.INIT('h80)
	) name3163 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]/P0001 ,
		_w5567_,
		_w5572_,
		_w6175_
	);
	LUT3 #(
		.INIT('h80)
	) name3164 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]/P0001 ,
		_w5566_,
		_w5564_,
		_w6176_
	);
	LUT3 #(
		.INIT('h80)
	) name3165 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]/P0001 ,
		_w5570_,
		_w5564_,
		_w6177_
	);
	LUT4 #(
		.INIT('h0001)
	) name3166 (
		_w6174_,
		_w6175_,
		_w6176_,
		_w6177_,
		_w6178_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3167 (
		_w6173_,
		_w6178_,
		_w6163_,
		_w6168_,
		_w6179_
	);
	LUT3 #(
		.INIT('h80)
	) name3168 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]/P0001 ,
		_w5569_,
		_w5559_,
		_w6180_
	);
	LUT3 #(
		.INIT('h80)
	) name3169 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]/P0001 ,
		_w5566_,
		_w5567_,
		_w6181_
	);
	LUT3 #(
		.INIT('h80)
	) name3170 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]/P0001 ,
		_w5566_,
		_w5564_,
		_w6182_
	);
	LUT3 #(
		.INIT('h80)
	) name3171 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]/P0001 ,
		_w5559_,
		_w5564_,
		_w6183_
	);
	LUT4 #(
		.INIT('h0001)
	) name3172 (
		_w6180_,
		_w6181_,
		_w6182_,
		_w6183_,
		_w6184_
	);
	LUT3 #(
		.INIT('h80)
	) name3173 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]/P0001 ,
		_w5576_,
		_w5572_,
		_w6185_
	);
	LUT3 #(
		.INIT('h80)
	) name3174 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]/P0001 ,
		_w5564_,
		_w5572_,
		_w6186_
	);
	LUT3 #(
		.INIT('h80)
	) name3175 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]/P0001 ,
		_w5570_,
		_w5564_,
		_w6187_
	);
	LUT3 #(
		.INIT('h80)
	) name3176 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]/P0001 ,
		_w5570_,
		_w5567_,
		_w6188_
	);
	LUT4 #(
		.INIT('h0001)
	) name3177 (
		_w6185_,
		_w6186_,
		_w6187_,
		_w6188_,
		_w6189_
	);
	LUT3 #(
		.INIT('h80)
	) name3178 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]/P0001 ,
		_w5566_,
		_w5576_,
		_w6190_
	);
	LUT3 #(
		.INIT('h80)
	) name3179 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]/P0001 ,
		_w5567_,
		_w5572_,
		_w6191_
	);
	LUT3 #(
		.INIT('h80)
	) name3180 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]/P0001 ,
		_w5569_,
		_w5566_,
		_w6192_
	);
	LUT3 #(
		.INIT('h80)
	) name3181 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]/P0001 ,
		_w5576_,
		_w5559_,
		_w6193_
	);
	LUT4 #(
		.INIT('h0001)
	) name3182 (
		_w6190_,
		_w6191_,
		_w6192_,
		_w6193_,
		_w6194_
	);
	LUT3 #(
		.INIT('h80)
	) name3183 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]/P0001 ,
		_w5569_,
		_w5572_,
		_w6195_
	);
	LUT3 #(
		.INIT('h80)
	) name3184 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]/P0001 ,
		_w5576_,
		_w5570_,
		_w6196_
	);
	LUT3 #(
		.INIT('h80)
	) name3185 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]/P0001 ,
		_w5569_,
		_w5570_,
		_w6197_
	);
	LUT3 #(
		.INIT('h80)
	) name3186 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]/P0001 ,
		_w5559_,
		_w5567_,
		_w6198_
	);
	LUT4 #(
		.INIT('h0001)
	) name3187 (
		_w6195_,
		_w6196_,
		_w6197_,
		_w6198_,
		_w6199_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3188 (
		_w6194_,
		_w6199_,
		_w6184_,
		_w6189_,
		_w6200_
	);
	LUT3 #(
		.INIT('h80)
	) name3189 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]/P0001 ,
		_w5576_,
		_w5559_,
		_w6201_
	);
	LUT3 #(
		.INIT('h80)
	) name3190 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]/P0001 ,
		_w5576_,
		_w5570_,
		_w6202_
	);
	LUT3 #(
		.INIT('h80)
	) name3191 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]/P0001 ,
		_w5559_,
		_w5567_,
		_w6203_
	);
	LUT3 #(
		.INIT('h80)
	) name3192 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]/P0001 ,
		_w5566_,
		_w5567_,
		_w6204_
	);
	LUT4 #(
		.INIT('h0001)
	) name3193 (
		_w6201_,
		_w6202_,
		_w6203_,
		_w6204_,
		_w6205_
	);
	LUT3 #(
		.INIT('h80)
	) name3194 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]/P0001 ,
		_w5566_,
		_w5576_,
		_w6206_
	);
	LUT3 #(
		.INIT('h80)
	) name3195 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]/P0001 ,
		_w5569_,
		_w5559_,
		_w6207_
	);
	LUT3 #(
		.INIT('h80)
	) name3196 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]/P0001 ,
		_w5569_,
		_w5570_,
		_w6208_
	);
	LUT3 #(
		.INIT('h80)
	) name3197 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]/P0001 ,
		_w5567_,
		_w5572_,
		_w6209_
	);
	LUT4 #(
		.INIT('h0001)
	) name3198 (
		_w6206_,
		_w6207_,
		_w6208_,
		_w6209_,
		_w6210_
	);
	LUT3 #(
		.INIT('h80)
	) name3199 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]/P0001 ,
		_w5569_,
		_w5566_,
		_w6211_
	);
	LUT3 #(
		.INIT('h80)
	) name3200 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]/P0001 ,
		_w5570_,
		_w5567_,
		_w6212_
	);
	LUT3 #(
		.INIT('h80)
	) name3201 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]/P0001 ,
		_w5566_,
		_w5564_,
		_w6213_
	);
	LUT3 #(
		.INIT('h80)
	) name3202 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]/P0001 ,
		_w5559_,
		_w5564_,
		_w6214_
	);
	LUT4 #(
		.INIT('h0001)
	) name3203 (
		_w6211_,
		_w6212_,
		_w6213_,
		_w6214_,
		_w6215_
	);
	LUT3 #(
		.INIT('h80)
	) name3204 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]/P0001 ,
		_w5576_,
		_w5572_,
		_w6216_
	);
	LUT3 #(
		.INIT('h80)
	) name3205 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]/P0001 ,
		_w5564_,
		_w5572_,
		_w6217_
	);
	LUT3 #(
		.INIT('h80)
	) name3206 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]/P0001 ,
		_w5570_,
		_w5564_,
		_w6218_
	);
	LUT3 #(
		.INIT('h80)
	) name3207 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]/P0001 ,
		_w5569_,
		_w5572_,
		_w6219_
	);
	LUT4 #(
		.INIT('h0001)
	) name3208 (
		_w6216_,
		_w6217_,
		_w6218_,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3209 (
		_w6215_,
		_w6220_,
		_w6205_,
		_w6210_,
		_w6221_
	);
	LUT3 #(
		.INIT('h80)
	) name3210 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]/P0001 ,
		_w5559_,
		_w5564_,
		_w6222_
	);
	LUT3 #(
		.INIT('h80)
	) name3211 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]/P0001 ,
		_w5566_,
		_w5567_,
		_w6223_
	);
	LUT3 #(
		.INIT('h80)
	) name3212 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]/P0001 ,
		_w5566_,
		_w5576_,
		_w6224_
	);
	LUT3 #(
		.INIT('h80)
	) name3213 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]/P0001 ,
		_w5569_,
		_w5559_,
		_w6225_
	);
	LUT4 #(
		.INIT('h0001)
	) name3214 (
		_w6222_,
		_w6223_,
		_w6224_,
		_w6225_,
		_w6226_
	);
	LUT3 #(
		.INIT('h80)
	) name3215 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]/P0001 ,
		_w5570_,
		_w5564_,
		_w6227_
	);
	LUT3 #(
		.INIT('h80)
	) name3216 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]/P0001 ,
		_w5570_,
		_w5567_,
		_w6228_
	);
	LUT3 #(
		.INIT('h80)
	) name3217 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]/P0001 ,
		_w5569_,
		_w5566_,
		_w6229_
	);
	LUT3 #(
		.INIT('h80)
	) name3218 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]/P0001 ,
		_w5576_,
		_w5559_,
		_w6230_
	);
	LUT4 #(
		.INIT('h0001)
	) name3219 (
		_w6227_,
		_w6228_,
		_w6229_,
		_w6230_,
		_w6231_
	);
	LUT3 #(
		.INIT('h80)
	) name3220 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]/P0001 ,
		_w5566_,
		_w5564_,
		_w6232_
	);
	LUT3 #(
		.INIT('h80)
	) name3221 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]/P0001 ,
		_w5567_,
		_w5572_,
		_w6233_
	);
	LUT3 #(
		.INIT('h80)
	) name3222 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]/P0001 ,
		_w5576_,
		_w5572_,
		_w6234_
	);
	LUT3 #(
		.INIT('h80)
	) name3223 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]/P0001 ,
		_w5564_,
		_w5572_,
		_w6235_
	);
	LUT4 #(
		.INIT('h0001)
	) name3224 (
		_w6232_,
		_w6233_,
		_w6234_,
		_w6235_,
		_w6236_
	);
	LUT3 #(
		.INIT('h80)
	) name3225 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]/P0001 ,
		_w5569_,
		_w5572_,
		_w6237_
	);
	LUT3 #(
		.INIT('h80)
	) name3226 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]/P0001 ,
		_w5576_,
		_w5570_,
		_w6238_
	);
	LUT3 #(
		.INIT('h80)
	) name3227 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]/P0001 ,
		_w5569_,
		_w5570_,
		_w6239_
	);
	LUT3 #(
		.INIT('h80)
	) name3228 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]/P0001 ,
		_w5559_,
		_w5567_,
		_w6240_
	);
	LUT4 #(
		.INIT('h0001)
	) name3229 (
		_w6237_,
		_w6238_,
		_w6239_,
		_w6240_,
		_w6241_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3230 (
		_w6236_,
		_w6241_,
		_w6226_,
		_w6231_,
		_w6242_
	);
	LUT3 #(
		.INIT('h80)
	) name3231 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]/P0001 ,
		_w5576_,
		_w5570_,
		_w6243_
	);
	LUT3 #(
		.INIT('h80)
	) name3232 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]/P0001 ,
		_w5566_,
		_w5567_,
		_w6244_
	);
	LUT3 #(
		.INIT('h80)
	) name3233 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]/P0001 ,
		_w5569_,
		_w5570_,
		_w6245_
	);
	LUT3 #(
		.INIT('h80)
	) name3234 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]/P0001 ,
		_w5567_,
		_w5572_,
		_w6246_
	);
	LUT4 #(
		.INIT('h0001)
	) name3235 (
		_w6243_,
		_w6244_,
		_w6245_,
		_w6246_,
		_w6247_
	);
	LUT3 #(
		.INIT('h80)
	) name3236 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]/P0001 ,
		_w5569_,
		_w5566_,
		_w6248_
	);
	LUT3 #(
		.INIT('h80)
	) name3237 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]/P0001 ,
		_w5576_,
		_w5559_,
		_w6249_
	);
	LUT3 #(
		.INIT('h80)
	) name3238 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]/P0001 ,
		_w5570_,
		_w5564_,
		_w6250_
	);
	LUT3 #(
		.INIT('h80)
	) name3239 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]/P0001 ,
		_w5570_,
		_w5567_,
		_w6251_
	);
	LUT4 #(
		.INIT('h0001)
	) name3240 (
		_w6248_,
		_w6249_,
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT3 #(
		.INIT('h80)
	) name3241 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]/P0001 ,
		_w5569_,
		_w5572_,
		_w6253_
	);
	LUT3 #(
		.INIT('h80)
	) name3242 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]/P0001 ,
		_w5559_,
		_w5564_,
		_w6254_
	);
	LUT3 #(
		.INIT('h80)
	) name3243 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]/P0001 ,
		_w5576_,
		_w5572_,
		_w6255_
	);
	LUT3 #(
		.INIT('h80)
	) name3244 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]/P0001 ,
		_w5564_,
		_w5572_,
		_w6256_
	);
	LUT4 #(
		.INIT('h0001)
	) name3245 (
		_w6253_,
		_w6254_,
		_w6255_,
		_w6256_,
		_w6257_
	);
	LUT3 #(
		.INIT('h80)
	) name3246 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]/P0001 ,
		_w5566_,
		_w5576_,
		_w6258_
	);
	LUT3 #(
		.INIT('h80)
	) name3247 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]/P0001 ,
		_w5569_,
		_w5559_,
		_w6259_
	);
	LUT3 #(
		.INIT('h80)
	) name3248 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]/P0001 ,
		_w5566_,
		_w5564_,
		_w6260_
	);
	LUT3 #(
		.INIT('h80)
	) name3249 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]/P0001 ,
		_w5559_,
		_w5567_,
		_w6261_
	);
	LUT4 #(
		.INIT('h0001)
	) name3250 (
		_w6258_,
		_w6259_,
		_w6260_,
		_w6261_,
		_w6262_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3251 (
		_w6257_,
		_w6262_,
		_w6247_,
		_w6252_,
		_w6263_
	);
	LUT3 #(
		.INIT('h80)
	) name3252 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]/P0001 ,
		_w5576_,
		_w5570_,
		_w6264_
	);
	LUT3 #(
		.INIT('h80)
	) name3253 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]/P0001 ,
		_w5566_,
		_w5567_,
		_w6265_
	);
	LUT3 #(
		.INIT('h80)
	) name3254 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]/P0001 ,
		_w5566_,
		_w5564_,
		_w6266_
	);
	LUT3 #(
		.INIT('h80)
	) name3255 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]/P0001 ,
		_w5559_,
		_w5564_,
		_w6267_
	);
	LUT4 #(
		.INIT('h0001)
	) name3256 (
		_w6264_,
		_w6265_,
		_w6266_,
		_w6267_,
		_w6268_
	);
	LUT3 #(
		.INIT('h80)
	) name3257 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]/P0001 ,
		_w5569_,
		_w5566_,
		_w6269_
	);
	LUT3 #(
		.INIT('h80)
	) name3258 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]/P0001 ,
		_w5576_,
		_w5559_,
		_w6270_
	);
	LUT3 #(
		.INIT('h80)
	) name3259 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]/P0001 ,
		_w5570_,
		_w5564_,
		_w6271_
	);
	LUT3 #(
		.INIT('h80)
	) name3260 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]/P0001 ,
		_w5570_,
		_w5567_,
		_w6272_
	);
	LUT4 #(
		.INIT('h0001)
	) name3261 (
		_w6269_,
		_w6270_,
		_w6271_,
		_w6272_,
		_w6273_
	);
	LUT3 #(
		.INIT('h80)
	) name3262 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]/P0001 ,
		_w5569_,
		_w5572_,
		_w6274_
	);
	LUT3 #(
		.INIT('h80)
	) name3263 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]/P0001 ,
		_w5567_,
		_w5572_,
		_w6275_
	);
	LUT3 #(
		.INIT('h80)
	) name3264 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]/P0001 ,
		_w5576_,
		_w5572_,
		_w6276_
	);
	LUT3 #(
		.INIT('h80)
	) name3265 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]/P0001 ,
		_w5564_,
		_w5572_,
		_w6277_
	);
	LUT4 #(
		.INIT('h0001)
	) name3266 (
		_w6274_,
		_w6275_,
		_w6276_,
		_w6277_,
		_w6278_
	);
	LUT3 #(
		.INIT('h80)
	) name3267 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]/P0001 ,
		_w5566_,
		_w5576_,
		_w6279_
	);
	LUT3 #(
		.INIT('h80)
	) name3268 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]/P0001 ,
		_w5569_,
		_w5559_,
		_w6280_
	);
	LUT3 #(
		.INIT('h80)
	) name3269 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]/P0001 ,
		_w5569_,
		_w5570_,
		_w6281_
	);
	LUT3 #(
		.INIT('h80)
	) name3270 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]/P0001 ,
		_w5559_,
		_w5567_,
		_w6282_
	);
	LUT4 #(
		.INIT('h0001)
	) name3271 (
		_w6279_,
		_w6280_,
		_w6281_,
		_w6282_,
		_w6283_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3272 (
		_w6278_,
		_w6283_,
		_w6268_,
		_w6273_,
		_w6284_
	);
	LUT3 #(
		.INIT('h80)
	) name3273 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]/P0001 ,
		_w5566_,
		_w5567_,
		_w6285_
	);
	LUT3 #(
		.INIT('h80)
	) name3274 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]/P0001 ,
		_w5567_,
		_w5572_,
		_w6286_
	);
	LUT3 #(
		.INIT('h80)
	) name3275 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]/P0001 ,
		_w5569_,
		_w5566_,
		_w6287_
	);
	LUT3 #(
		.INIT('h80)
	) name3276 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]/P0001 ,
		_w5576_,
		_w5559_,
		_w6288_
	);
	LUT4 #(
		.INIT('h0001)
	) name3277 (
		_w6285_,
		_w6286_,
		_w6287_,
		_w6288_,
		_w6289_
	);
	LUT3 #(
		.INIT('h80)
	) name3278 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]/P0001 ,
		_w5566_,
		_w5576_,
		_w6290_
	);
	LUT3 #(
		.INIT('h80)
	) name3279 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]/P0001 ,
		_w5569_,
		_w5559_,
		_w6291_
	);
	LUT3 #(
		.INIT('h80)
	) name3280 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]/P0001 ,
		_w5566_,
		_w5564_,
		_w6292_
	);
	LUT3 #(
		.INIT('h80)
	) name3281 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]/P0001 ,
		_w5559_,
		_w5564_,
		_w6293_
	);
	LUT4 #(
		.INIT('h0001)
	) name3282 (
		_w6290_,
		_w6291_,
		_w6292_,
		_w6293_,
		_w6294_
	);
	LUT3 #(
		.INIT('h80)
	) name3283 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]/P0001 ,
		_w5559_,
		_w5567_,
		_w6295_
	);
	LUT3 #(
		.INIT('h80)
	) name3284 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]/P0001 ,
		_w5570_,
		_w5567_,
		_w6296_
	);
	LUT3 #(
		.INIT('h80)
	) name3285 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]/P0001 ,
		_w5569_,
		_w5572_,
		_w6297_
	);
	LUT3 #(
		.INIT('h80)
	) name3286 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]/P0001 ,
		_w5576_,
		_w5570_,
		_w6298_
	);
	LUT4 #(
		.INIT('h0001)
	) name3287 (
		_w6295_,
		_w6296_,
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT3 #(
		.INIT('h80)
	) name3288 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]/P0001 ,
		_w5576_,
		_w5572_,
		_w6300_
	);
	LUT3 #(
		.INIT('h80)
	) name3289 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]/P0001 ,
		_w5564_,
		_w5572_,
		_w6301_
	);
	LUT3 #(
		.INIT('h80)
	) name3290 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]/P0001 ,
		_w5570_,
		_w5564_,
		_w6302_
	);
	LUT3 #(
		.INIT('h80)
	) name3291 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]/P0001 ,
		_w5569_,
		_w5570_,
		_w6303_
	);
	LUT4 #(
		.INIT('h0001)
	) name3292 (
		_w6300_,
		_w6301_,
		_w6302_,
		_w6303_,
		_w6304_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3293 (
		_w6299_,
		_w6304_,
		_w6289_,
		_w6294_,
		_w6305_
	);
	LUT4 #(
		.INIT('h2622)
	) name3294 (
		\pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg/NET0131 ,
		_w3229_,
		_w3251_,
		_w3259_,
		_w6306_
	);
	LUT3 #(
		.INIT('h47)
	) name3295 (
		\output_backup_stop_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		pci_stop_i_pad,
		_w6307_
	);
	LUT3 #(
		.INIT('hb8)
	) name3296 (
		\output_backup_stop_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		pci_stop_i_pad,
		_w6308_
	);
	LUT3 #(
		.INIT('h54)
	) name3297 (
		_w3206_,
		_w3789_,
		_w6307_,
		_w6309_
	);
	LUT4 #(
		.INIT('h0100)
	) name3298 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w6310_
	);
	LUT4 #(
		.INIT('haabf)
	) name3299 (
		pci_gnt_i_pad,
		_w3793_,
		_w3795_,
		_w6310_,
		_w6311_
	);
	LUT3 #(
		.INIT('h07)
	) name3300 (
		\output_backup_frame_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w6312_
	);
	LUT4 #(
		.INIT('hffeb)
	) name3301 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w6313_
	);
	LUT4 #(
		.INIT('h0014)
	) name3302 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w6314_
	);
	LUT4 #(
		.INIT('ha888)
	) name3303 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]/NET0131 ,
		_w3792_,
		_w3786_,
		_w6312_,
		_w6315_
	);
	LUT3 #(
		.INIT('h51)
	) name3304 (
		_w6309_,
		_w6311_,
		_w6315_,
		_w6316_
	);
	LUT4 #(
		.INIT('hfecf)
	) name3305 (
		\pci_target_unit_pci_target_sm_backoff_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w6317_
	);
	LUT4 #(
		.INIT('h1033)
	) name3306 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w3224_,
		_w6317_,
		_w6318_
	);
	LUT4 #(
		.INIT('h4044)
	) name3307 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3216_,
		_w3717_,
		_w3750_,
		_w6319_
	);
	LUT3 #(
		.INIT('h54)
	) name3308 (
		_w6309_,
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT4 #(
		.INIT('h0400)
	) name3309 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131 ,
		_w6321_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3310 (
		_w3212_,
		_w3215_,
		_w3221_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6323_
	);
	LUT3 #(
		.INIT('h02)
	) name3312 (
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_read_completed_reg_reg/NET0131 ,
		_w6324_
	);
	LUT3 #(
		.INIT('h01)
	) name3313 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\input_register_pci_trdy_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		_w6325_
	);
	LUT4 #(
		.INIT('h2000)
	) name3314 (
		\output_backup_trdy_en_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131 ,
		_w6326_
	);
	LUT3 #(
		.INIT('h15)
	) name3315 (
		_w6324_,
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('hb)
	) name3316 (
		_w6322_,
		_w6327_,
		_w6328_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3317 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6329_
	);
	LUT4 #(
		.INIT('h2022)
	) name3318 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6330_
	);
	LUT2 #(
		.INIT('h1)
	) name3319 (
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT4 #(
		.INIT('h2022)
	) name3320 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6332_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3321 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6333_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3322 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6334_
	);
	LUT4 #(
		.INIT('h2022)
	) name3323 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6335_
	);
	LUT4 #(
		.INIT('h000e)
	) name3324 (
		_w6332_,
		_w6333_,
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3325 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]/P0001 ,
		_w6331_,
		_w6336_,
		_w6337_
	);
	LUT4 #(
		.INIT('heee0)
	) name3326 (
		_w6332_,
		_w6333_,
		_w6334_,
		_w6335_,
		_w6338_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3327 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]/P0001 ,
		_w6331_,
		_w6338_,
		_w6339_
	);
	LUT4 #(
		.INIT('h0001)
	) name3328 (
		_w6332_,
		_w6333_,
		_w6334_,
		_w6335_,
		_w6340_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3329 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]/P0001 ,
		_w6331_,
		_w6340_,
		_w6341_
	);
	LUT4 #(
		.INIT('h1110)
	) name3330 (
		_w6332_,
		_w6333_,
		_w6334_,
		_w6335_,
		_w6342_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3331 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]/P0001 ,
		_w6331_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3332 (
		_w6341_,
		_w6343_,
		_w6337_,
		_w6339_,
		_w6344_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3333 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]/P0001 ,
		_w6331_,
		_w6342_,
		_w6345_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3334 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]/P0001 ,
		_w6331_,
		_w6338_,
		_w6346_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3335 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]/P0001 ,
		_w6331_,
		_w6336_,
		_w6347_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3336 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]/P0001 ,
		_w6331_,
		_w6340_,
		_w6348_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3337 (
		_w6347_,
		_w6348_,
		_w6345_,
		_w6346_,
		_w6349_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3338 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]/P0001 ,
		_w6331_,
		_w6342_,
		_w6350_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3339 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]/P0001 ,
		_w6331_,
		_w6340_,
		_w6351_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3340 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]/P0001 ,
		_w6331_,
		_w6336_,
		_w6352_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3341 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]/P0001 ,
		_w6331_,
		_w6338_,
		_w6353_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3342 (
		_w6352_,
		_w6353_,
		_w6350_,
		_w6351_,
		_w6354_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3343 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]/P0001 ,
		_w6331_,
		_w6340_,
		_w6355_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3344 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]/P0001 ,
		_w6331_,
		_w6342_,
		_w6356_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3345 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]/P0001 ,
		_w6331_,
		_w6336_,
		_w6357_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3346 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]/P0001 ,
		_w6331_,
		_w6338_,
		_w6358_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3347 (
		_w6357_,
		_w6358_,
		_w6355_,
		_w6356_,
		_w6359_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3348 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]/P0001 ,
		_w6331_,
		_w6340_,
		_w6360_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3349 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]/P0001 ,
		_w6331_,
		_w6342_,
		_w6361_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3350 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]/P0001 ,
		_w6331_,
		_w6336_,
		_w6362_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3351 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]/P0001 ,
		_w6331_,
		_w6338_,
		_w6363_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3352 (
		_w6362_,
		_w6363_,
		_w6360_,
		_w6361_,
		_w6364_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3353 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]/P0001 ,
		_w6331_,
		_w6340_,
		_w6365_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3354 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]/P0001 ,
		_w6331_,
		_w6338_,
		_w6366_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3355 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]/P0001 ,
		_w6331_,
		_w6336_,
		_w6367_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3356 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]/P0001 ,
		_w6331_,
		_w6342_,
		_w6368_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3357 (
		_w6367_,
		_w6368_,
		_w6365_,
		_w6366_,
		_w6369_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3358 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]/P0001 ,
		_w6331_,
		_w6338_,
		_w6370_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3359 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]/P0001 ,
		_w6331_,
		_w6336_,
		_w6371_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3360 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]/P0001 ,
		_w6331_,
		_w6342_,
		_w6372_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3361 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]/P0001 ,
		_w6331_,
		_w6340_,
		_w6373_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3362 (
		_w6372_,
		_w6373_,
		_w6370_,
		_w6371_,
		_w6374_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3363 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]/P0001 ,
		_w6331_,
		_w6340_,
		_w6375_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3364 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]/P0001 ,
		_w6331_,
		_w6342_,
		_w6376_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3365 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]/P0001 ,
		_w6331_,
		_w6336_,
		_w6377_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3366 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]/P0001 ,
		_w6331_,
		_w6338_,
		_w6378_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3367 (
		_w6377_,
		_w6378_,
		_w6375_,
		_w6376_,
		_w6379_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3368 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]/P0001 ,
		_w6331_,
		_w6338_,
		_w6380_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3369 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]/P0001 ,
		_w6331_,
		_w6342_,
		_w6381_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3370 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]/P0001 ,
		_w6331_,
		_w6340_,
		_w6382_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3371 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]/P0001 ,
		_w6331_,
		_w6336_,
		_w6383_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3372 (
		_w6382_,
		_w6383_,
		_w6380_,
		_w6381_,
		_w6384_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3373 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]/P0001 ,
		_w6331_,
		_w6342_,
		_w6385_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3374 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]/P0001 ,
		_w6331_,
		_w6338_,
		_w6386_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3375 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]/P0001 ,
		_w6331_,
		_w6340_,
		_w6387_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3376 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]/P0001 ,
		_w6331_,
		_w6336_,
		_w6388_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3377 (
		_w6387_,
		_w6388_,
		_w6385_,
		_w6386_,
		_w6389_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3378 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]/P0001 ,
		_w6331_,
		_w6340_,
		_w6390_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3379 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]/P0001 ,
		_w6331_,
		_w6338_,
		_w6391_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3380 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]/P0001 ,
		_w6331_,
		_w6336_,
		_w6392_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3381 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]/P0001 ,
		_w6331_,
		_w6342_,
		_w6393_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3382 (
		_w6392_,
		_w6393_,
		_w6390_,
		_w6391_,
		_w6394_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3383 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]/P0001 ,
		_w6331_,
		_w6340_,
		_w6395_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3384 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]/P0001 ,
		_w6331_,
		_w6342_,
		_w6396_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3385 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]/P0001 ,
		_w6331_,
		_w6338_,
		_w6397_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3386 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]/P0001 ,
		_w6331_,
		_w6336_,
		_w6398_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3387 (
		_w6397_,
		_w6398_,
		_w6395_,
		_w6396_,
		_w6399_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3388 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]/P0001 ,
		_w6331_,
		_w6336_,
		_w6400_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3389 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]/P0001 ,
		_w6331_,
		_w6342_,
		_w6401_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3390 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]/P0001 ,
		_w6331_,
		_w6340_,
		_w6402_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3391 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]/P0001 ,
		_w6331_,
		_w6338_,
		_w6403_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3392 (
		_w6402_,
		_w6403_,
		_w6400_,
		_w6401_,
		_w6404_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3393 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]/P0001 ,
		_w6331_,
		_w6340_,
		_w6405_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3394 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]/P0001 ,
		_w6331_,
		_w6336_,
		_w6406_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3395 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]/P0001 ,
		_w6331_,
		_w6342_,
		_w6407_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3396 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]/P0001 ,
		_w6331_,
		_w6338_,
		_w6408_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3397 (
		_w6407_,
		_w6408_,
		_w6405_,
		_w6406_,
		_w6409_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3398 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]/P0001 ,
		_w6331_,
		_w6336_,
		_w6410_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3399 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]/P0001 ,
		_w6331_,
		_w6340_,
		_w6411_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3400 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]/P0001 ,
		_w6331_,
		_w6338_,
		_w6412_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3401 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]/P0001 ,
		_w6331_,
		_w6342_,
		_w6413_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3402 (
		_w6412_,
		_w6413_,
		_w6410_,
		_w6411_,
		_w6414_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3403 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]/P0001 ,
		_w6331_,
		_w6342_,
		_w6415_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3404 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]/P0001 ,
		_w6331_,
		_w6338_,
		_w6416_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3405 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]/P0001 ,
		_w6331_,
		_w6340_,
		_w6417_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3406 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]/P0001 ,
		_w6331_,
		_w6336_,
		_w6418_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3407 (
		_w6417_,
		_w6418_,
		_w6415_,
		_w6416_,
		_w6419_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3408 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]/P0001 ,
		_w6331_,
		_w6338_,
		_w6420_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3409 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]/P0001 ,
		_w6331_,
		_w6340_,
		_w6421_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3410 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]/P0001 ,
		_w6331_,
		_w6336_,
		_w6422_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3411 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]/P0001 ,
		_w6331_,
		_w6342_,
		_w6423_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3412 (
		_w6422_,
		_w6423_,
		_w6420_,
		_w6421_,
		_w6424_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3413 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]/P0001 ,
		_w6331_,
		_w6338_,
		_w6425_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3414 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]/P0001 ,
		_w6331_,
		_w6342_,
		_w6426_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3415 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]/P0001 ,
		_w6331_,
		_w6340_,
		_w6427_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3416 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]/P0001 ,
		_w6331_,
		_w6336_,
		_w6428_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3417 (
		_w6427_,
		_w6428_,
		_w6425_,
		_w6426_,
		_w6429_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3418 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]/P0001 ,
		_w6331_,
		_w6336_,
		_w6430_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3419 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]/P0001 ,
		_w6331_,
		_w6342_,
		_w6431_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3420 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]/P0001 ,
		_w6331_,
		_w6340_,
		_w6432_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3421 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]/P0001 ,
		_w6331_,
		_w6338_,
		_w6433_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3422 (
		_w6432_,
		_w6433_,
		_w6430_,
		_w6431_,
		_w6434_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3423 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]/P0001 ,
		_w6331_,
		_w6340_,
		_w6435_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3424 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]/P0001 ,
		_w6331_,
		_w6342_,
		_w6436_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3425 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]/P0001 ,
		_w6331_,
		_w6336_,
		_w6437_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3426 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]/P0001 ,
		_w6331_,
		_w6338_,
		_w6438_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3427 (
		_w6437_,
		_w6438_,
		_w6435_,
		_w6436_,
		_w6439_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3428 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]/P0001 ,
		_w6331_,
		_w6342_,
		_w6440_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3429 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]/P0001 ,
		_w6331_,
		_w6340_,
		_w6441_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3430 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]/P0001 ,
		_w6331_,
		_w6338_,
		_w6442_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3431 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]/P0001 ,
		_w6331_,
		_w6336_,
		_w6443_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3432 (
		_w6442_,
		_w6443_,
		_w6440_,
		_w6441_,
		_w6444_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3433 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]/P0001 ,
		_w6331_,
		_w6342_,
		_w6445_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3434 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]/P0001 ,
		_w6331_,
		_w6336_,
		_w6446_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3435 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]/P0001 ,
		_w6331_,
		_w6338_,
		_w6447_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3436 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]/P0001 ,
		_w6331_,
		_w6340_,
		_w6448_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3437 (
		_w6447_,
		_w6448_,
		_w6445_,
		_w6446_,
		_w6449_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3438 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]/P0001 ,
		_w6331_,
		_w6336_,
		_w6450_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3439 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]/P0001 ,
		_w6331_,
		_w6340_,
		_w6451_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3440 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]/P0001 ,
		_w6331_,
		_w6338_,
		_w6452_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3441 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]/P0001 ,
		_w6331_,
		_w6342_,
		_w6453_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3442 (
		_w6452_,
		_w6453_,
		_w6450_,
		_w6451_,
		_w6454_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3443 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]/P0001 ,
		_w6331_,
		_w6338_,
		_w6455_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3444 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]/P0001 ,
		_w6331_,
		_w6342_,
		_w6456_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3445 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]/P0001 ,
		_w6331_,
		_w6340_,
		_w6457_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3446 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]/P0001 ,
		_w6331_,
		_w6336_,
		_w6458_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3447 (
		_w6457_,
		_w6458_,
		_w6455_,
		_w6456_,
		_w6459_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3448 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]/P0001 ,
		_w6331_,
		_w6342_,
		_w6460_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3449 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]/P0001 ,
		_w6331_,
		_w6336_,
		_w6461_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3450 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]/P0001 ,
		_w6331_,
		_w6338_,
		_w6462_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3451 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]/P0001 ,
		_w6331_,
		_w6340_,
		_w6463_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3452 (
		_w6462_,
		_w6463_,
		_w6460_,
		_w6461_,
		_w6464_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3453 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]/P0001 ,
		_w6331_,
		_w6342_,
		_w6465_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3454 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]/P0001 ,
		_w6331_,
		_w6340_,
		_w6466_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3455 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]/P0001 ,
		_w6331_,
		_w6336_,
		_w6467_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3456 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]/P0001 ,
		_w6331_,
		_w6338_,
		_w6468_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3457 (
		_w6467_,
		_w6468_,
		_w6465_,
		_w6466_,
		_w6469_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3458 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]/P0001 ,
		_w6331_,
		_w6336_,
		_w6470_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3459 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]/P0001 ,
		_w6331_,
		_w6338_,
		_w6471_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3460 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]/P0001 ,
		_w6331_,
		_w6340_,
		_w6472_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3461 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]/P0001 ,
		_w6331_,
		_w6342_,
		_w6473_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3462 (
		_w6472_,
		_w6473_,
		_w6470_,
		_w6471_,
		_w6474_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3463 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]/P0001 ,
		_w6331_,
		_w6340_,
		_w6475_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3464 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]/P0001 ,
		_w6331_,
		_w6336_,
		_w6476_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3465 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]/P0001 ,
		_w6331_,
		_w6338_,
		_w6477_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3466 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]/P0001 ,
		_w6331_,
		_w6342_,
		_w6478_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3467 (
		_w6477_,
		_w6478_,
		_w6475_,
		_w6476_,
		_w6479_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3468 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]/P0001 ,
		_w6331_,
		_w6336_,
		_w6480_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3469 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]/P0001 ,
		_w6331_,
		_w6338_,
		_w6481_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3470 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]/P0001 ,
		_w6331_,
		_w6342_,
		_w6482_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3471 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]/P0001 ,
		_w6331_,
		_w6340_,
		_w6483_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3472 (
		_w6482_,
		_w6483_,
		_w6480_,
		_w6481_,
		_w6484_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3473 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]/P0001 ,
		_w6331_,
		_w6336_,
		_w6485_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3474 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]/P0001 ,
		_w6331_,
		_w6342_,
		_w6486_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3475 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]/P0001 ,
		_w6331_,
		_w6340_,
		_w6487_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3476 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]/P0001 ,
		_w6331_,
		_w6338_,
		_w6488_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3477 (
		_w6487_,
		_w6488_,
		_w6485_,
		_w6486_,
		_w6489_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3478 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]/P0001 ,
		_w6331_,
		_w6338_,
		_w6490_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3479 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]/P0001 ,
		_w6331_,
		_w6340_,
		_w6491_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3480 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]/P0001 ,
		_w6331_,
		_w6342_,
		_w6492_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3481 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]/P0001 ,
		_w6331_,
		_w6336_,
		_w6493_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3482 (
		_w6492_,
		_w6493_,
		_w6490_,
		_w6491_,
		_w6494_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3483 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]/P0001 ,
		_w6331_,
		_w6336_,
		_w6495_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3484 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]/P0001 ,
		_w6331_,
		_w6338_,
		_w6496_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3485 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]/P0001 ,
		_w6331_,
		_w6340_,
		_w6497_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3486 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]/P0001 ,
		_w6331_,
		_w6342_,
		_w6498_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3487 (
		_w6497_,
		_w6498_,
		_w6495_,
		_w6496_,
		_w6499_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3488 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]/P0001 ,
		_w6331_,
		_w6340_,
		_w6500_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3489 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]/P0001 ,
		_w6331_,
		_w6336_,
		_w6501_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3490 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]/P0001 ,
		_w6331_,
		_w6342_,
		_w6502_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3491 (
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]/P0001 ,
		\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]/P0001 ,
		_w6331_,
		_w6338_,
		_w6503_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3492 (
		_w6502_,
		_w6503_,
		_w6500_,
		_w6501_,
		_w6504_
	);
	LUT3 #(
		.INIT('h80)
	) name3493 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		_w6505_
	);
	LUT4 #(
		.INIT('h8000)
	) name3494 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131 ,
		_w6506_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		_w6506_,
		_w6507_
	);
	LUT3 #(
		.INIT('h80)
	) name3496 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		_w6506_,
		_w6508_
	);
	LUT4 #(
		.INIT('h8000)
	) name3497 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131 ,
		_w6506_,
		_w6509_
	);
	LUT3 #(
		.INIT('h80)
	) name3498 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		_w6509_,
		_w6510_
	);
	LUT4 #(
		.INIT('h8000)
	) name3499 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131 ,
		_w6509_,
		_w6511_
	);
	LUT3 #(
		.INIT('h80)
	) name3500 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		_w6511_,
		_w6512_
	);
	LUT4 #(
		.INIT('h8000)
	) name3501 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131 ,
		_w6511_,
		_w6513_
	);
	LUT3 #(
		.INIT('h80)
	) name3502 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		_w6513_,
		_w6514_
	);
	LUT4 #(
		.INIT('h8000)
	) name3503 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131 ,
		_w6513_,
		_w6515_
	);
	LUT4 #(
		.INIT('h0004)
	) name3504 (
		\output_backup_trdy_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w6516_
	);
	LUT3 #(
		.INIT('h04)
	) name3505 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131 ,
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6517_
	);
	LUT2 #(
		.INIT('h4)
	) name3506 (
		_w6516_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		_w6515_,
		_w6518_,
		_w6519_
	);
	LUT4 #(
		.INIT('h8000)
	) name3508 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131 ,
		_w6520_
	);
	LUT4 #(
		.INIT('h8000)
	) name3509 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131 ,
		_w6520_,
		_w6521_
	);
	LUT4 #(
		.INIT('h8000)
	) name3510 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131 ,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		_w6522_,
		_w6523_
	);
	LUT3 #(
		.INIT('h80)
	) name3512 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		_w6522_,
		_w6524_
	);
	LUT4 #(
		.INIT('h8000)
	) name3513 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131 ,
		_w6522_,
		_w6525_
	);
	LUT3 #(
		.INIT('h80)
	) name3514 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		_w6525_,
		_w6526_
	);
	LUT4 #(
		.INIT('h8000)
	) name3515 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131 ,
		_w6525_,
		_w6527_
	);
	LUT3 #(
		.INIT('h04)
	) name3516 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]/NET0131 ,
		\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6528_
	);
	LUT2 #(
		.INIT('h4)
	) name3517 (
		_w3166_,
		_w6528_,
		_w6529_
	);
	LUT3 #(
		.INIT('h70)
	) name3518 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h8)
	) name3519 (
		_w6527_,
		_w6530_,
		_w6531_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3520 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6329_,
		_w6330_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name3521 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6533_
	);
	LUT3 #(
		.INIT('hc8)
	) name3522 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6534_
	);
	LUT4 #(
		.INIT('hca00)
	) name3523 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6535_
	);
	LUT2 #(
		.INIT('he)
	) name3524 (
		_w6534_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h2)
	) name3525 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		_w6537_
	);
	LUT4 #(
		.INIT('h0222)
	) name3526 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\input_register_pci_stop_reg_out_reg/NET0131 ,
		\input_register_pci_trdy_reg_out_reg/NET0131 ,
		_w6538_
	);
	LUT2 #(
		.INIT('h2)
	) name3527 (
		_w3205_,
		_w6538_,
		_w6539_
	);
	LUT4 #(
		.INIT('h1511)
	) name3528 (
		_w3212_,
		_w3216_,
		_w3717_,
		_w3750_,
		_w6540_
	);
	LUT2 #(
		.INIT('h4)
	) name3529 (
		_w6539_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('hb)
	) name3530 (
		_w6539_,
		_w6540_,
		_w6542_
	);
	LUT3 #(
		.INIT('h06)
	) name3531 (
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w6543_
	);
	LUT3 #(
		.INIT('hf9)
	) name3532 (
		\pci_target_unit_pci_target_sm_c_state_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_c_state_reg[2]/NET0131 ,
		_w6544_
	);
	LUT3 #(
		.INIT('h07)
	) name3533 (
		_w3205_,
		_w3206_,
		_w6543_,
		_w6545_
	);
	LUT2 #(
		.INIT('hd)
	) name3534 (
		_w6540_,
		_w6545_,
		_w6546_
	);
	LUT4 #(
		.INIT('h9a99)
	) name3535 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6547_
	);
	LUT3 #(
		.INIT('h74)
	) name3536 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6547_,
		_w6548_
	);
	LUT4 #(
		.INIT('ha533)
	) name3537 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6549_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3538 (
		_w3145_,
		_w3135_,
		_w3157_,
		_w3158_,
		_w6550_
	);
	LUT4 #(
		.INIT('haa08)
	) name3539 (
		_w3135_,
		_w3147_,
		_w3150_,
		_w3158_,
		_w6551_
	);
	LUT3 #(
		.INIT('h54)
	) name3540 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT4 #(
		.INIT('h0001)
	) name3541 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6553_
	);
	LUT4 #(
		.INIT('h5400)
	) name3542 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6555_
	);
	LUT3 #(
		.INIT('he2)
	) name3544 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]/P0001 ,
		_w6554_,
		_w6555_,
		_w6556_
	);
	LUT4 #(
		.INIT('h0400)
	) name3545 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6557_
	);
	LUT4 #(
		.INIT('h5400)
	) name3546 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6557_,
		_w6558_
	);
	LUT3 #(
		.INIT('hca)
	) name3547 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]/P0001 ,
		_w6555_,
		_w6558_,
		_w6559_
	);
	LUT4 #(
		.INIT('h1000)
	) name3548 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6560_
	);
	LUT4 #(
		.INIT('h5400)
	) name3549 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6560_,
		_w6561_
	);
	LUT3 #(
		.INIT('hca)
	) name3550 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]/P0001 ,
		_w6555_,
		_w6561_,
		_w6562_
	);
	LUT4 #(
		.INIT('h0002)
	) name3551 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6563_
	);
	LUT4 #(
		.INIT('h5400)
	) name3552 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6563_,
		_w6564_
	);
	LUT3 #(
		.INIT('hca)
	) name3553 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]/P0001 ,
		_w6555_,
		_w6564_,
		_w6565_
	);
	LUT4 #(
		.INIT('h0004)
	) name3554 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6566_
	);
	LUT4 #(
		.INIT('h5400)
	) name3555 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6566_,
		_w6567_
	);
	LUT3 #(
		.INIT('hca)
	) name3556 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]/P0001 ,
		_w6555_,
		_w6567_,
		_w6568_
	);
	LUT4 #(
		.INIT('h0008)
	) name3557 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6569_
	);
	LUT4 #(
		.INIT('h5400)
	) name3558 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6569_,
		_w6570_
	);
	LUT3 #(
		.INIT('hca)
	) name3559 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]/P0001 ,
		_w6555_,
		_w6570_,
		_w6571_
	);
	LUT4 #(
		.INIT('h0010)
	) name3560 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6572_
	);
	LUT4 #(
		.INIT('h5400)
	) name3561 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6572_,
		_w6573_
	);
	LUT3 #(
		.INIT('hca)
	) name3562 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]/P0001 ,
		_w6555_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h0020)
	) name3563 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6575_
	);
	LUT4 #(
		.INIT('h5400)
	) name3564 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6575_,
		_w6576_
	);
	LUT3 #(
		.INIT('hca)
	) name3565 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]/P0001 ,
		_w6555_,
		_w6576_,
		_w6577_
	);
	LUT4 #(
		.INIT('h0040)
	) name3566 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6578_
	);
	LUT4 #(
		.INIT('h5400)
	) name3567 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6578_,
		_w6579_
	);
	LUT3 #(
		.INIT('hca)
	) name3568 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]/P0001 ,
		_w6555_,
		_w6579_,
		_w6580_
	);
	LUT4 #(
		.INIT('h0100)
	) name3569 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6581_
	);
	LUT4 #(
		.INIT('h5400)
	) name3570 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6581_,
		_w6582_
	);
	LUT3 #(
		.INIT('hca)
	) name3571 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]/P0001 ,
		_w6555_,
		_w6582_,
		_w6583_
	);
	LUT4 #(
		.INIT('h0200)
	) name3572 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6584_
	);
	LUT4 #(
		.INIT('h5400)
	) name3573 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6584_,
		_w6585_
	);
	LUT3 #(
		.INIT('hca)
	) name3574 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]/P0001 ,
		_w6555_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name3575 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6587_
	);
	LUT4 #(
		.INIT('h2220)
	) name3576 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w3154_,
		_w6550_,
		_w6551_,
		_w6588_
	);
	LUT3 #(
		.INIT('h80)
	) name3577 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT4 #(
		.INIT('h0800)
	) name3578 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6590_
	);
	LUT4 #(
		.INIT('h5400)
	) name3579 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6590_,
		_w6591_
	);
	LUT4 #(
		.INIT('h2000)
	) name3580 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6592_
	);
	LUT4 #(
		.INIT('h5400)
	) name3581 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6592_,
		_w6593_
	);
	LUT4 #(
		.INIT('h4000)
	) name3582 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6594_
	);
	LUT4 #(
		.INIT('h5400)
	) name3583 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6594_,
		_w6595_
	);
	LUT4 #(
		.INIT('h8000)
	) name3584 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6596_
	);
	LUT4 #(
		.INIT('h5400)
	) name3585 (
		_w3154_,
		_w6550_,
		_w6551_,
		_w6596_,
		_w6597_
	);
	LUT3 #(
		.INIT('h60)
	) name3586 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[12]/NET0131 ,
		_w6512_,
		_w6518_,
		_w6598_
	);
	LUT3 #(
		.INIT('h60)
	) name3587 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]/NET0131 ,
		_w6524_,
		_w6530_,
		_w6599_
	);
	LUT3 #(
		.INIT('h08)
	) name3588 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w5166_,
		_w6600_
	);
	LUT4 #(
		.INIT('h0080)
	) name3589 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w5166_,
		_w6601_
	);
	LUT4 #(
		.INIT('h0080)
	) name3590 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6602_
	);
	LUT4 #(
		.INIT('h807f)
	) name3591 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6603_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3592 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6604_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		_w6533_,
		_w6603_,
		_w6605_
	);
	LUT4 #(
		.INIT('h007b)
	) name3594 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 ,
		_w6533_,
		_w6601_,
		_w6605_,
		_w6606_
	);
	LUT4 #(
		.INIT('h0903)
	) name3595 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6330_,
		_w6607_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w6608_
	);
	LUT3 #(
		.INIT('h78)
	) name3597 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w6609_
	);
	LUT4 #(
		.INIT('h8700)
	) name3598 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6610_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		_w6607_,
		_w6610_,
		_w6611_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w6612_
	);
	LUT3 #(
		.INIT('h60)
	) name3601 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6613_
	);
	LUT4 #(
		.INIT('hff12)
	) name3602 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6330_,
		_w6613_,
		_w6614_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3603 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6332_,
		_w6333_,
		_w6615_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3604 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6334_,
		_w6335_,
		_w6616_
	);
	LUT4 #(
		.INIT('h1011)
	) name3605 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6617_
	);
	LUT4 #(
		.INIT('h4544)
	) name3606 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6618_
	);
	LUT4 #(
		.INIT('h888b)
	) name3607 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6618_,
		_w6617_,
		_w6619_
	);
	LUT4 #(
		.INIT('h1011)
	) name3608 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6620_
	);
	LUT4 #(
		.INIT('h4544)
	) name3609 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6621_
	);
	LUT4 #(
		.INIT('h888b)
	) name3610 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6621_,
		_w6620_,
		_w6622_
	);
	LUT4 #(
		.INIT('h1011)
	) name3611 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6623_
	);
	LUT4 #(
		.INIT('h4544)
	) name3612 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6624_
	);
	LUT4 #(
		.INIT('h888b)
	) name3613 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6624_,
		_w6623_,
		_w6625_
	);
	LUT2 #(
		.INIT('h6)
	) name3614 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w6626_
	);
	LUT4 #(
		.INIT('h0045)
	) name3615 (
		_w3255_,
		_w6322_,
		_w6327_,
		_w6626_,
		_w6627_
	);
	LUT4 #(
		.INIT('h4544)
	) name3616 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6628_
	);
	LUT4 #(
		.INIT('h888b)
	) name3617 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6628_,
		_w6627_,
		_w6629_
	);
	LUT2 #(
		.INIT('h9)
	) name3618 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w6630_
	);
	LUT4 #(
		.INIT('h0045)
	) name3619 (
		_w3255_,
		_w6322_,
		_w6327_,
		_w6630_,
		_w6631_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3620 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6632_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3621 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6631_,
		_w6632_,
		_w6633_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3622 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6634_
	);
	LUT4 #(
		.INIT('h2022)
	) name3623 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w3255_,
		_w6322_,
		_w6327_,
		_w6635_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3624 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg/NET0131 ,
		_w6634_,
		_w6635_,
		_w6636_
	);
	LUT3 #(
		.INIT('h78)
	) name3625 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w6637_
	);
	LUT2 #(
		.INIT('h4)
	) name3626 (
		_w6533_,
		_w6637_,
		_w6638_
	);
	LUT4 #(
		.INIT('hff48)
	) name3627 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w6533_,
		_w6600_,
		_w6638_,
		_w6639_
	);
	LUT4 #(
		.INIT('h3c28)
	) name3628 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6640_
	);
	LUT4 #(
		.INIT('hc600)
	) name3629 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6641_
	);
	LUT2 #(
		.INIT('he)
	) name3630 (
		_w6640_,
		_w6641_,
		_w6642_
	);
	LUT3 #(
		.INIT('hc8)
	) name3631 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6643_
	);
	LUT4 #(
		.INIT('hca00)
	) name3632 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6644_
	);
	LUT2 #(
		.INIT('he)
	) name3633 (
		_w6643_,
		_w6644_,
		_w6645_
	);
	LUT4 #(
		.INIT('hca00)
	) name3634 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6646_
	);
	LUT3 #(
		.INIT('hc8)
	) name3635 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6647_
	);
	LUT2 #(
		.INIT('he)
	) name3636 (
		_w6646_,
		_w6647_,
		_w6648_
	);
	LUT4 #(
		.INIT('hca00)
	) name3637 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6649_
	);
	LUT3 #(
		.INIT('hc8)
	) name3638 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6650_
	);
	LUT2 #(
		.INIT('he)
	) name3639 (
		_w6649_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h6)
	) name3640 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w6652_
	);
	LUT4 #(
		.INIT('hb080)
	) name3641 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('he)
	) name3642 (
		_w6643_,
		_w6653_,
		_w6654_
	);
	LUT3 #(
		.INIT('hc8)
	) name3643 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6655_
	);
	LUT2 #(
		.INIT('h6)
	) name3644 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w6656_
	);
	LUT4 #(
		.INIT('hb080)
	) name3645 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6656_,
		_w6657_
	);
	LUT2 #(
		.INIT('he)
	) name3646 (
		_w6655_,
		_w6657_,
		_w6658_
	);
	LUT3 #(
		.INIT('hc8)
	) name3647 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6659_
	);
	LUT2 #(
		.INIT('h6)
	) name3648 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131 ,
		_w6660_
	);
	LUT4 #(
		.INIT('hb080)
	) name3649 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('he)
	) name3650 (
		_w6659_,
		_w6661_,
		_w6662_
	);
	LUT3 #(
		.INIT('hc8)
	) name3651 (
		\wishbone_slave_unit_del_sync_comp_flush_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg/NET0131 ,
		_w6663_
	);
	LUT4 #(
		.INIT('hca00)
	) name3652 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]/NET0131 ,
		_w5166_,
		_w6533_,
		_w6664_
	);
	LUT2 #(
		.INIT('he)
	) name3653 (
		_w6663_,
		_w6664_,
		_w6665_
	);
	LUT3 #(
		.INIT('h80)
	) name3654 (
		_w3216_,
		_w3728_,
		_w3747_,
		_w6666_
	);
	LUT4 #(
		.INIT('h0080)
	) name3655 (
		_w3216_,
		_w3728_,
		_w3747_,
		_w6323_,
		_w6667_
	);
	LUT4 #(
		.INIT('hef00)
	) name3656 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_progress_reg/NET0131 ,
		_w6668_
	);
	LUT3 #(
		.INIT('h02)
	) name3657 (
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w6669_
	);
	LUT4 #(
		.INIT('h8000)
	) name3658 (
		_w3015_,
		_w3016_,
		_w3216_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w6668_,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('hb)
	) name3660 (
		_w6667_,
		_w6671_,
		_w6672_
	);
	LUT3 #(
		.INIT('h14)
	) name3661 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 ,
		wbm_rty_i_pad,
		_w6673_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3662 (
		wbm_rty_i_pad,
		_w3053_,
		_w3055_,
		_w6673_,
		_w6674_
	);
	LUT2 #(
		.INIT('h4)
	) name3663 (
		_w3154_,
		_w6550_,
		_w6675_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name3664 (
		\wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131 ,
		_w3154_,
		_w6550_,
		_w6676_
	);
	LUT4 #(
		.INIT('hef00)
	) name3665 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_request_reg/NET0131 ,
		_w6677_
	);
	LUT2 #(
		.INIT('h1)
	) name3666 (
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6678_
	);
	LUT4 #(
		.INIT('h2a00)
	) name3667 (
		_w3216_,
		_w3728_,
		_w3747_,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('he)
	) name3668 (
		_w6677_,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6681_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		\wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131 ,
		_w3140_,
		_w6682_
	);
	LUT4 #(
		.INIT('h8000)
	) name3671 (
		_w3147_,
		_w3150_,
		_w6681_,
		_w6682_,
		_w6683_
	);
	LUT2 #(
		.INIT('h1)
	) name3672 (
		\wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131 ,
		_w6684_
	);
	LUT3 #(
		.INIT('h08)
	) name3673 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		_w6685_
	);
	LUT2 #(
		.INIT('h4)
	) name3674 (
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('he2)
	) name3675 (
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		_w6683_,
		_w6686_,
		_w6687_
	);
	LUT3 #(
		.INIT('h80)
	) name3676 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]/P0001 ,
		_w5566_,
		_w5567_,
		_w6688_
	);
	LUT3 #(
		.INIT('h80)
	) name3677 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]/P0001 ,
		_w5567_,
		_w5572_,
		_w6689_
	);
	LUT3 #(
		.INIT('h80)
	) name3678 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]/P0001 ,
		_w5570_,
		_w5567_,
		_w6690_
	);
	LUT3 #(
		.INIT('h80)
	) name3679 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]/P0001 ,
		_w5570_,
		_w5564_,
		_w6691_
	);
	LUT4 #(
		.INIT('h0001)
	) name3680 (
		_w6688_,
		_w6689_,
		_w6690_,
		_w6691_,
		_w6692_
	);
	LUT3 #(
		.INIT('h80)
	) name3681 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]/P0001 ,
		_w5566_,
		_w5576_,
		_w6693_
	);
	LUT3 #(
		.INIT('h80)
	) name3682 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]/P0001 ,
		_w5569_,
		_w5559_,
		_w6694_
	);
	LUT3 #(
		.INIT('h80)
	) name3683 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]/P0001 ,
		_w5566_,
		_w5564_,
		_w6695_
	);
	LUT3 #(
		.INIT('h80)
	) name3684 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]/P0001 ,
		_w5559_,
		_w5564_,
		_w6696_
	);
	LUT4 #(
		.INIT('h0001)
	) name3685 (
		_w6693_,
		_w6694_,
		_w6695_,
		_w6696_,
		_w6697_
	);
	LUT3 #(
		.INIT('h80)
	) name3686 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]/P0001 ,
		_w5559_,
		_w5567_,
		_w6698_
	);
	LUT3 #(
		.INIT('h80)
	) name3687 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]/P0001 ,
		_w5564_,
		_w5572_,
		_w6699_
	);
	LUT3 #(
		.INIT('h80)
	) name3688 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]/P0001 ,
		_w5569_,
		_w5572_,
		_w6700_
	);
	LUT3 #(
		.INIT('h80)
	) name3689 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]/P0001 ,
		_w5576_,
		_w5570_,
		_w6701_
	);
	LUT4 #(
		.INIT('h0001)
	) name3690 (
		_w6698_,
		_w6699_,
		_w6700_,
		_w6701_,
		_w6702_
	);
	LUT3 #(
		.INIT('h80)
	) name3691 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]/P0001 ,
		_w5576_,
		_w5559_,
		_w6703_
	);
	LUT3 #(
		.INIT('h80)
	) name3692 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]/P0001 ,
		_w5569_,
		_w5566_,
		_w6704_
	);
	LUT3 #(
		.INIT('h80)
	) name3693 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]/P0001 ,
		_w5576_,
		_w5572_,
		_w6705_
	);
	LUT3 #(
		.INIT('h80)
	) name3694 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]/P0001 ,
		_w5569_,
		_w5570_,
		_w6706_
	);
	LUT4 #(
		.INIT('h0001)
	) name3695 (
		_w6703_,
		_w6704_,
		_w6705_,
		_w6706_,
		_w6707_
	);
	LUT4 #(
		.INIT('h7fff)
	) name3696 (
		_w6702_,
		_w6707_,
		_w6692_,
		_w6697_,
		_w6708_
	);
	LUT3 #(
		.INIT('h9a)
	) name3697 (
		\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131 ,
		_w3154_,
		_w6550_,
		_w6709_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3698 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		_w6509_,
		_w6518_,
		_w6710_
	);
	LUT2 #(
		.INIT('h2)
	) name3699 (
		_w3050_,
		_w3062_,
		_w6711_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3700 (
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_c_state_reg[2]/NET0131 ,
		_w6712_
	);
	LUT4 #(
		.INIT('h0007)
	) name3701 (
		_w3060_,
		_w3068_,
		_w3101_,
		_w6712_,
		_w6713_
	);
	LUT3 #(
		.INIT('hb0)
	) name3702 (
		_w3067_,
		_w3070_,
		_w6713_,
		_w6714_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3703 (
		_w3084_,
		_w3087_,
		_w6711_,
		_w6714_,
		_w6715_
	);
	LUT3 #(
		.INIT('h6c)
	) name3704 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		_w6521_,
		_w6716_
	);
	LUT4 #(
		.INIT('h7000)
	) name3705 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h6)
	) name3706 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w6588_,
		_w6718_
	);
	LUT4 #(
		.INIT('hef00)
	) name3707 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_prf_en_reg/NET0131 ,
		_w6719_
	);
	LUT4 #(
		.INIT('h0888)
	) name3708 (
		\configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131 ,
		_w3216_,
		_w3728_,
		_w3747_,
		_w6720_
	);
	LUT2 #(
		.INIT('he)
	) name3709 (
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT4 #(
		.INIT('he222)
	) name3710 (
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w3216_,
		_w3728_,
		_w3747_,
		_w6722_
	);
	LUT4 #(
		.INIT('hef00)
	) name3711 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_wr_progress_reg/NET0131 ,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		_w6724_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		_w3216_,
		_w6724_,
		_w6725_
	);
	LUT3 #(
		.INIT('h10)
	) name3714 (
		_w3233_,
		_w3246_,
		_w6725_,
		_w6726_
	);
	LUT3 #(
		.INIT('h13)
	) name3715 (
		_w3242_,
		_w6723_,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('hb)
	) name3716 (
		_w6666_,
		_w6727_,
		_w6728_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131 ,
		_w6729_
	);
	LUT4 #(
		.INIT('h3a0a)
	) name3718 (
		\wishbone_slave_unit_del_sync_bc_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		_w6683_,
		_w6729_,
		_w6730_
	);
	LUT3 #(
		.INIT('hc8)
	) name3719 (
		_w3789_,
		_w3786_,
		_w6307_,
		_w6731_
	);
	LUT4 #(
		.INIT('h0006)
	) name3720 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w6732_
	);
	LUT2 #(
		.INIT('h1)
	) name3721 (
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		_w6732_,
		_w6733_
	);
	LUT3 #(
		.INIT('h20)
	) name3722 (
		\output_backup_frame_out_reg/NET0131 ,
		_w6731_,
		_w6733_,
		_w6734_
	);
	LUT3 #(
		.INIT('hc4)
	) name3723 (
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131 ,
		_w6735_
	);
	LUT3 #(
		.INIT('h40)
	) name3724 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		_w3018_,
		_w3019_,
		_w6736_
	);
	LUT4 #(
		.INIT('hc888)
	) name3725 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w6737_
	);
	LUT3 #(
		.INIT('hba)
	) name3726 (
		_w6735_,
		_w6736_,
		_w6737_,
		_w6738_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3727 (
		_w3786_,
		_w6735_,
		_w6736_,
		_w6737_,
		_w6739_
	);
	LUT3 #(
		.INIT('h01)
	) name3728 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131 ,
		_w6740_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131 ,
		_w6741_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131 ,
		_w6742_
	);
	LUT4 #(
		.INIT('h0001)
	) name3731 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131 ,
		_w6743_
	);
	LUT3 #(
		.INIT('h80)
	) name3732 (
		pci_gnt_i_pad,
		_w6740_,
		_w6743_,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		\wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		_w6745_
	);
	LUT2 #(
		.INIT('h4)
	) name3734 (
		_w6307_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h4)
	) name3735 (
		_w6744_,
		_w6746_,
		_w6747_
	);
	LUT3 #(
		.INIT('h45)
	) name3736 (
		_w3793_,
		_w6731_,
		_w6733_,
		_w6748_
	);
	LUT4 #(
		.INIT('hefaa)
	) name3737 (
		_w6734_,
		_w6739_,
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT3 #(
		.INIT('h20)
	) name3738 (
		pci_frame_o_pad,
		_w6731_,
		_w6733_,
		_w6750_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3739 (
		_w6739_,
		_w6747_,
		_w6748_,
		_w6750_,
		_w6751_
	);
	LUT4 #(
		.INIT('h999a)
	) name3740 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w3154_,
		_w6550_,
		_w6551_,
		_w6752_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		\configuration_latency_timer_reg[7]/NET0131 ,
		_w6313_,
		_w6753_
	);
	LUT4 #(
		.INIT('h0111)
	) name3742 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131 ,
		_w6313_,
		_w6740_,
		_w6743_,
		_w6754_
	);
	LUT3 #(
		.INIT('h40)
	) name3743 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131 ,
		_w6742_,
		_w6754_,
		_w6755_
	);
	LUT4 #(
		.INIT('h1000)
	) name3744 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131 ,
		_w6742_,
		_w6754_,
		_w6756_
	);
	LUT4 #(
		.INIT('h0222)
	) name3745 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]/NET0131 ,
		_w6313_,
		_w6741_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('he)
	) name3746 (
		_w6753_,
		_w6757_,
		_w6758_
	);
	LUT3 #(
		.INIT('h80)
	) name3747 (
		\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131 ,
		wbm_rty_i_pad,
		_w6759_
	);
	LUT4 #(
		.INIT('h8000)
	) name3748 (
		\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131 ,
		wbm_rty_i_pad,
		_w6760_
	);
	LUT3 #(
		.INIT('h80)
	) name3749 (
		\pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131 ,
		_w3054_,
		_w6760_,
		_w6761_
	);
	LUT4 #(
		.INIT('h1444)
	) name3750 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131 ,
		_w3054_,
		_w6760_,
		_w6762_
	);
	LUT4 #(
		.INIT('h8000)
	) name3751 (
		\pci_target_unit_wishbone_master_rty_counter_reg[5]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131 ,
		_w3054_,
		_w6760_,
		_w6763_
	);
	LUT3 #(
		.INIT('h14)
	) name3752 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[6]/NET0131 ,
		_w6761_,
		_w6764_
	);
	LUT3 #(
		.INIT('h14)
	) name3753 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[7]/NET0131 ,
		_w6763_,
		_w6765_
	);
	LUT2 #(
		.INIT('h6)
	) name3754 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		_w6766_
	);
	LUT4 #(
		.INIT('h7000)
	) name3755 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6766_,
		_w6767_
	);
	LUT3 #(
		.INIT('h60)
	) name3756 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		_w6522_,
		_w6530_,
		_w6768_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3757 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]/NET0131 ,
		_w6521_,
		_w6769_
	);
	LUT4 #(
		.INIT('h7000)
	) name3758 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('hd)
	) name3759 (
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6771_
	);
	LUT2 #(
		.INIT('hd)
	) name3760 (
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6772_
	);
	LUT4 #(
		.INIT('h1500)
	) name3761 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		_w3149_,
		_w3147_,
		_w6529_,
		_w6773_
	);
	LUT3 #(
		.INIT('h60)
	) name3762 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		_w6523_,
		_w6530_,
		_w6774_
	);
	LUT3 #(
		.INIT('h60)
	) name3763 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		_w6525_,
		_w6530_,
		_w6775_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3764 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		_w6525_,
		_w6530_,
		_w6776_
	);
	LUT3 #(
		.INIT('h60)
	) name3765 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]/NET0131 ,
		_w6526_,
		_w6530_,
		_w6777_
	);
	LUT3 #(
		.INIT('h78)
	) name3766 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		_w6778_
	);
	LUT4 #(
		.INIT('h7000)
	) name3767 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6778_,
		_w6779_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3768 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]/NET0131 ,
		_w6780_
	);
	LUT4 #(
		.INIT('h7000)
	) name3769 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6780_,
		_w6781_
	);
	LUT2 #(
		.INIT('h6)
	) name3770 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		_w6520_,
		_w6782_
	);
	LUT4 #(
		.INIT('h7000)
	) name3771 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6782_,
		_w6783_
	);
	LUT3 #(
		.INIT('h6c)
	) name3772 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		_w6520_,
		_w6784_
	);
	LUT4 #(
		.INIT('h7000)
	) name3773 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3774 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]/NET0131 ,
		_w6520_,
		_w6786_
	);
	LUT4 #(
		.INIT('h7000)
	) name3775 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h6)
	) name3776 (
		\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		_w6521_,
		_w6788_
	);
	LUT4 #(
		.INIT('h7000)
	) name3777 (
		_w3149_,
		_w3147_,
		_w6529_,
		_w6788_,
		_w6789_
	);
	LUT3 #(
		.INIT('h35)
	) name3778 (
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6790_
	);
	LUT3 #(
		.INIT('h14)
	) name3779 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[2]/NET0131 ,
		_w6759_,
		_w6791_
	);
	LUT3 #(
		.INIT('h14)
	) name3780 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131 ,
		_w6760_,
		_w6792_
	);
	LUT4 #(
		.INIT('h1450)
	) name3781 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[3]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[4]/NET0131 ,
		_w6760_,
		_w6793_
	);
	LUT3 #(
		.INIT('h3a)
	) name3782 (
		\wishbone_slave_unit_del_sync_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		_w6683_,
		_w6794_
	);
	LUT3 #(
		.INIT('h6c)
	) name3783 (
		\pci_target_unit_wishbone_master_rty_counter_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_rty_counter_reg[1]/NET0131 ,
		wbm_rty_i_pad,
		_w6795_
	);
	LUT4 #(
		.INIT('h007f)
	) name3784 (
		wbm_rty_i_pad,
		_w3053_,
		_w3055_,
		_w6795_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name3785 (
		\pci_target_unit_wishbone_master_reset_rty_cnt_reg/NET0131 ,
		_w6796_,
		_w6797_
	);
	LUT3 #(
		.INIT('hac)
	) name3786 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6798_
	);
	LUT3 #(
		.INIT('hac)
	) name3787 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6799_
	);
	LUT3 #(
		.INIT('hac)
	) name3788 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6800_
	);
	LUT3 #(
		.INIT('hac)
	) name3789 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6801_
	);
	LUT3 #(
		.INIT('hac)
	) name3790 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6802_
	);
	LUT3 #(
		.INIT('hac)
	) name3791 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6803_
	);
	LUT3 #(
		.INIT('hac)
	) name3792 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6804_
	);
	LUT3 #(
		.INIT('hac)
	) name3793 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6805_
	);
	LUT3 #(
		.INIT('hac)
	) name3794 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6806_
	);
	LUT3 #(
		.INIT('hac)
	) name3795 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6807_
	);
	LUT3 #(
		.INIT('hac)
	) name3796 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6808_
	);
	LUT3 #(
		.INIT('hac)
	) name3797 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6809_
	);
	LUT3 #(
		.INIT('hac)
	) name3798 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6810_
	);
	LUT3 #(
		.INIT('hac)
	) name3799 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6811_
	);
	LUT3 #(
		.INIT('hac)
	) name3800 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6812_
	);
	LUT3 #(
		.INIT('hac)
	) name3801 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6813_
	);
	LUT3 #(
		.INIT('hac)
	) name3802 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6814_
	);
	LUT3 #(
		.INIT('hac)
	) name3803 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6815_
	);
	LUT3 #(
		.INIT('hac)
	) name3804 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6816_
	);
	LUT3 #(
		.INIT('hac)
	) name3805 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6817_
	);
	LUT3 #(
		.INIT('hac)
	) name3806 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6818_
	);
	LUT3 #(
		.INIT('hac)
	) name3807 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6819_
	);
	LUT3 #(
		.INIT('hac)
	) name3808 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6820_
	);
	LUT3 #(
		.INIT('hac)
	) name3809 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6821_
	);
	LUT3 #(
		.INIT('hac)
	) name3810 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6822_
	);
	LUT3 #(
		.INIT('hac)
	) name3811 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6823_
	);
	LUT3 #(
		.INIT('hac)
	) name3812 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6824_
	);
	LUT3 #(
		.INIT('hac)
	) name3813 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6825_
	);
	LUT3 #(
		.INIT('hac)
	) name3814 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6826_
	);
	LUT3 #(
		.INIT('hac)
	) name3815 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6827_
	);
	LUT3 #(
		.INIT('hac)
	) name3816 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6828_
	);
	LUT3 #(
		.INIT('hac)
	) name3817 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg/NET0131 ,
		_w6829_
	);
	LUT2 #(
		.INIT('h8)
	) name3818 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w6830_
	);
	LUT2 #(
		.INIT('h2)
	) name3819 (
		\input_register_pci_devsel_reg_out_reg/NET0131 ,
		\input_register_pci_stop_reg_out_reg/NET0131 ,
		_w6831_
	);
	LUT2 #(
		.INIT('h2)
	) name3820 (
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w6832_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name3821 (
		\input_register_pci_devsel_reg_out_reg/NET0131 ,
		\input_register_pci_stop_reg_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w6833_
	);
	LUT2 #(
		.INIT('h4)
	) name3822 (
		\wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131 ,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('hd050)
	) name3823 (
		\input_register_pci_stop_reg_out_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131 ,
		_w6310_,
		_w6835_
	);
	LUT3 #(
		.INIT('ha2)
	) name3824 (
		_w6830_,
		_w6834_,
		_w6835_,
		_w6836_
	);
	LUT2 #(
		.INIT('h2)
	) name3825 (
		\wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 ,
		_w6837_
	);
	LUT3 #(
		.INIT('h80)
	) name3826 (
		_w3015_,
		_w3016_,
		_w6837_,
		_w6838_
	);
	LUT4 #(
		.INIT('h4000)
	) name3827 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3015_,
		_w3016_,
		_w6837_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w6836_,
		_w6840_,
		_w6841_
	);
	LUT3 #(
		.INIT('h60)
	) name3830 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[15]/NET0131 ,
		_w6514_,
		_w6518_,
		_w6842_
	);
	LUT2 #(
		.INIT('h4)
	) name3831 (
		\wishbone_slave_unit_del_sync_comp_done_reg_clr_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131 ,
		_w6843_
	);
	LUT4 #(
		.INIT('h8808)
	) name3832 (
		\wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131 ,
		_w6830_,
		_w6834_,
		_w6835_,
		_w6844_
	);
	LUT3 #(
		.INIT('h32)
	) name3833 (
		\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT4 #(
		.INIT('h1555)
	) name3834 (
		\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w3147_,
		_w3150_,
		_w6682_,
		_w6846_
	);
	LUT2 #(
		.INIT('h1)
	) name3835 (
		\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 ,
		_w6846_,
		_w6847_
	);
	LUT3 #(
		.INIT('h8a)
	) name3836 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		_w3021_,
		_w3030_,
		_w6848_
	);
	LUT4 #(
		.INIT('h8088)
	) name3837 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131 ,
		_w3021_,
		_w3030_,
		_w6849_
	);
	LUT2 #(
		.INIT('h6)
	) name3838 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		_w6849_,
		_w6850_
	);
	LUT3 #(
		.INIT('h0b)
	) name3839 (
		_w3064_,
		_w3065_,
		_w3632_,
		_w6851_
	);
	LUT4 #(
		.INIT('hff20)
	) name3840 (
		\pci_target_unit_wishbone_master_w_attempt_reg/NET0131 ,
		_w6711_,
		_w6714_,
		_w6851_,
		_w6852_
	);
	LUT4 #(
		.INIT('h9a99)
	) name3841 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		_w3017_,
		_w3021_,
		_w3030_,
		_w6853_
	);
	LUT4 #(
		.INIT('h6c66)
	) name3842 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131 ,
		_w3021_,
		_w3030_,
		_w6854_
	);
	LUT4 #(
		.INIT('h5540)
	) name3843 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131 ,
		_w3147_,
		_w3150_,
		_w3178_,
		_w6855_
	);
	LUT2 #(
		.INIT('h2)
	) name3844 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg/NET0131 ,
		wbs_stb_i_pad,
		_w6856_
	);
	LUT2 #(
		.INIT('he)
	) name3845 (
		_w6855_,
		_w6856_,
		_w6857_
	);
	LUT3 #(
		.INIT('hd8)
	) name3846 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[0]/NET0131 ,
		\pci_cbe_i[0]_pad ,
		_w6858_
	);
	LUT4 #(
		.INIT('h596a)
	) name3847 (
		\output_backup_ad_out_reg[19]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[0]/NET0131 ,
		\pci_cbe_i[0]_pad ,
		_w6859_
	);
	LUT3 #(
		.INIT('h27)
	) name3848 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[2]/NET0131 ,
		\pci_cbe_i[2]_pad ,
		_w6860_
	);
	LUT3 #(
		.INIT('hd8)
	) name3849 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[2]/NET0131 ,
		\pci_cbe_i[2]_pad ,
		_w6861_
	);
	LUT2 #(
		.INIT('h6)
	) name3850 (
		\output_backup_ad_out_reg[17]/NET0131 ,
		\output_backup_ad_out_reg[6]/NET0131 ,
		_w6862_
	);
	LUT4 #(
		.INIT('h6996)
	) name3851 (
		\output_backup_ad_out_reg[16]/NET0131 ,
		_w6859_,
		_w6860_,
		_w6862_,
		_w6863_
	);
	LUT4 #(
		.INIT('h9669)
	) name3852 (
		\output_backup_ad_out_reg[27]/NET0131 ,
		\output_backup_ad_out_reg[28]/NET0131 ,
		\output_backup_ad_out_reg[2]/NET0131 ,
		\output_backup_ad_out_reg[7]/NET0131 ,
		_w6864_
	);
	LUT4 #(
		.INIT('h6996)
	) name3853 (
		\output_backup_ad_out_reg[18]/NET0131 ,
		\output_backup_ad_out_reg[4]/NET0131 ,
		\output_backup_ad_out_reg[5]/NET0131 ,
		\output_backup_ad_out_reg[8]/NET0131 ,
		_w6865_
	);
	LUT2 #(
		.INIT('h9)
	) name3854 (
		\output_backup_ad_out_reg[12]/NET0131 ,
		\output_backup_ad_out_reg[9]/NET0131 ,
		_w6866_
	);
	LUT3 #(
		.INIT('h27)
	) name3855 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[3]/NET0131 ,
		\pci_cbe_i[3]_pad ,
		_w6867_
	);
	LUT3 #(
		.INIT('hd8)
	) name3856 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[3]/NET0131 ,
		\pci_cbe_i[3]_pad ,
		_w6868_
	);
	LUT2 #(
		.INIT('h9)
	) name3857 (
		\output_backup_ad_out_reg[24]/NET0131 ,
		\output_backup_ad_out_reg[26]/NET0131 ,
		_w6869_
	);
	LUT3 #(
		.INIT('hd8)
	) name3858 (
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[1]/NET0131 ,
		\pci_cbe_i[1]_pad ,
		_w6870_
	);
	LUT4 #(
		.INIT('h596a)
	) name3859 (
		\output_backup_ad_out_reg[0]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[1]/NET0131 ,
		\pci_cbe_i[1]_pad ,
		_w6871_
	);
	LUT4 #(
		.INIT('h6996)
	) name3860 (
		_w6866_,
		_w6867_,
		_w6869_,
		_w6871_,
		_w6872_
	);
	LUT4 #(
		.INIT('h9669)
	) name3861 (
		\output_backup_ad_out_reg[3]/NET0131 ,
		_w6864_,
		_w6865_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h9)
	) name3862 (
		\output_backup_ad_out_reg[30]/NET0131 ,
		\output_backup_ad_out_reg[31]/NET0131 ,
		_w6874_
	);
	LUT3 #(
		.INIT('h96)
	) name3863 (
		\output_backup_ad_out_reg[1]/NET0131 ,
		\output_backup_ad_out_reg[25]/NET0131 ,
		\output_backup_ad_out_reg[29]/NET0131 ,
		_w6875_
	);
	LUT2 #(
		.INIT('h6)
	) name3864 (
		\output_backup_ad_out_reg[11]/NET0131 ,
		\output_backup_ad_out_reg[13]/NET0131 ,
		_w6876_
	);
	LUT3 #(
		.INIT('h69)
	) name3865 (
		_w6874_,
		_w6875_,
		_w6876_,
		_w6877_
	);
	LUT2 #(
		.INIT('h9)
	) name3866 (
		\output_backup_ad_out_reg[14]/NET0131 ,
		\output_backup_ad_out_reg[15]/NET0131 ,
		_w6878_
	);
	LUT3 #(
		.INIT('h69)
	) name3867 (
		\output_backup_ad_out_reg[10]/NET0131 ,
		\output_backup_ad_out_reg[20]/NET0131 ,
		\output_backup_ad_out_reg[21]/NET0131 ,
		_w6879_
	);
	LUT2 #(
		.INIT('h6)
	) name3868 (
		\output_backup_ad_out_reg[22]/NET0131 ,
		\output_backup_ad_out_reg[23]/NET0131 ,
		_w6880_
	);
	LUT3 #(
		.INIT('h96)
	) name3869 (
		_w6878_,
		_w6879_,
		_w6880_,
		_w6881_
	);
	LUT2 #(
		.INIT('h9)
	) name3870 (
		_w6877_,
		_w6881_,
		_w6882_
	);
	LUT3 #(
		.INIT('h69)
	) name3871 (
		_w6863_,
		_w6873_,
		_w6882_,
		_w6883_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3872 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[14]/NET0131 ,
		_w6513_,
		_w6518_,
		_w6884_
	);
	LUT4 #(
		.INIT('h0600)
	) name3873 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[4]/NET0131 ,
		_w6506_,
		_w6516_,
		_w6517_,
		_w6885_
	);
	LUT3 #(
		.INIT('hdf)
	) name3874 (
		_w3051_,
		_w6711_,
		_w6714_,
		_w6886_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3875 (
		\wishbone_slave_unit_wishbone_slave_del_addr_hit_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6887_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3876 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131 ,
		_w6888_
	);
	LUT4 #(
		.INIT('hf531)
	) name3877 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131 ,
		_w6889_
	);
	LUT2 #(
		.INIT('h6)
	) name3878 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[2]/NET0131 ,
		_w6890_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3879 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[11]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131 ,
		_w6891_
	);
	LUT4 #(
		.INIT('h4000)
	) name3880 (
		_w6890_,
		_w6891_,
		_w6888_,
		_w6889_,
		_w6892_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3881 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131 ,
		_w6893_
	);
	LUT4 #(
		.INIT('hf531)
	) name3882 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131 ,
		_w6894_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3883 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[0]/NET0131 ,
		_w6895_
	);
	LUT4 #(
		.INIT('hf531)
	) name3884 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131 ,
		_w6896_
	);
	LUT4 #(
		.INIT('h8000)
	) name3885 (
		_w6895_,
		_w6896_,
		_w6893_,
		_w6894_,
		_w6897_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3886 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[15]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131 ,
		_w6898_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3887 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131 ,
		_w6899_
	);
	LUT4 #(
		.INIT('hf531)
	) name3888 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131 ,
		_w6900_
	);
	LUT4 #(
		.INIT('haf23)
	) name3889 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131 ,
		_w6901_
	);
	LUT4 #(
		.INIT('h8000)
	) name3890 (
		_w6900_,
		_w6901_,
		_w6898_,
		_w6899_,
		_w6902_
	);
	LUT3 #(
		.INIT('h80)
	) name3891 (
		_w6892_,
		_w6897_,
		_w6902_,
		_w6903_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3892 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[29]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131 ,
		_w6904_
	);
	LUT4 #(
		.INIT('hf531)
	) name3893 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[19]/NET0131 ,
		_w6905_
	);
	LUT4 #(
		.INIT('haf23)
	) name3894 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[14]/NET0131 ,
		_w6906_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3895 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131 ,
		_w6907_
	);
	LUT4 #(
		.INIT('h8000)
	) name3896 (
		_w6906_,
		_w6907_,
		_w6904_,
		_w6905_,
		_w6908_
	);
	LUT4 #(
		.INIT('haf23)
	) name3897 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[13]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131 ,
		_w6909_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3898 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131 ,
		_w6910_
	);
	LUT4 #(
		.INIT('haf23)
	) name3899 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[18]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[3]/NET0131 ,
		_w6911_
	);
	LUT4 #(
		.INIT('hf531)
	) name3900 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[12]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[26]/NET0131 ,
		_w6912_
	);
	LUT4 #(
		.INIT('h8000)
	) name3901 (
		_w6911_,
		_w6912_,
		_w6909_,
		_w6910_,
		_w6913_
	);
	LUT2 #(
		.INIT('h8)
	) name3902 (
		_w6908_,
		_w6913_,
		_w6914_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3903 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131 ,
		_w6915_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3904 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[25]/NET0131 ,
		_w6916_
	);
	LUT4 #(
		.INIT('hf531)
	) name3905 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[10]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[6]/NET0131 ,
		_w6917_
	);
	LUT4 #(
		.INIT('haf23)
	) name3906 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[21]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131 ,
		_w6918_
	);
	LUT4 #(
		.INIT('h8000)
	) name3907 (
		_w6917_,
		_w6918_,
		_w6915_,
		_w6916_,
		_w6919_
	);
	LUT4 #(
		.INIT('haf23)
	) name3908 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[16]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131 ,
		_w6920_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3909 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[20]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[30]/NET0131 ,
		_w6921_
	);
	LUT4 #(
		.INIT('hf531)
	) name3910 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[31]/NET0131 ,
		_w6922_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3911 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[24]/NET0131 ,
		_w6923_
	);
	LUT4 #(
		.INIT('h8000)
	) name3912 (
		_w6922_,
		_w6923_,
		_w6920_,
		_w6921_,
		_w6924_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3913 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[23]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[9]/NET0131 ,
		_w6925_
	);
	LUT4 #(
		.INIT('hf531)
	) name3914 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[22]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[8]/NET0131 ,
		_w6926_
	);
	LUT4 #(
		.INIT('haf23)
	) name3915 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131 ,
		_w6927_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3916 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[7]/NET0131 ,
		_w6928_
	);
	LUT4 #(
		.INIT('h8000)
	) name3917 (
		_w6927_,
		_w6928_,
		_w6925_,
		_w6926_,
		_w6929_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3918 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[17]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[2]/NET0131 ,
		_w6930_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3919 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[27]/NET0131 ,
		\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131 ,
		_w6931_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3920 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[5]/NET0131 ,
		_w6932_
	);
	LUT4 #(
		.INIT('hf531)
	) name3921 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[28]/NET0131 ,
		\wishbone_slave_unit_del_sync_addr_out_reg[4]/NET0131 ,
		_w6933_
	);
	LUT4 #(
		.INIT('h8000)
	) name3922 (
		_w6932_,
		_w6933_,
		_w6930_,
		_w6931_,
		_w6934_
	);
	LUT4 #(
		.INIT('h8000)
	) name3923 (
		_w6929_,
		_w6934_,
		_w6919_,
		_w6924_,
		_w6935_
	);
	LUT4 #(
		.INIT('h8000)
	) name3924 (
		_w3665_,
		_w6914_,
		_w6903_,
		_w6935_,
		_w6936_
	);
	LUT2 #(
		.INIT('he)
	) name3925 (
		_w6887_,
		_w6936_,
		_w6937_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3926 (
		\wishbone_slave_unit_wishbone_slave_do_del_request_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6938_
	);
	LUT4 #(
		.INIT('ha800)
	) name3927 (
		\configuration_sync_command_bit_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6939_
	);
	LUT3 #(
		.INIT('hec)
	) name3928 (
		_w6681_,
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3929 (
		\wishbone_slave_unit_wishbone_slave_img_wallow_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name3930 (
		\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w6942_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		_w3157_,
		_w6942_,
		_w6943_
	);
	LUT3 #(
		.INIT('hec)
	) name3932 (
		_w6939_,
		_w6941_,
		_w6943_,
		_w6944_
	);
	LUT3 #(
		.INIT('h82)
	) name3933 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6945_
	);
	LUT4 #(
		.INIT('h8020)
	) name3934 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		\configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6946_
	);
	LUT3 #(
		.INIT('h82)
	) name3935 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6947_
	);
	LUT4 #(
		.INIT('h8020)
	) name3936 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		\configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w6946_,
		_w6948_,
		_w6949_
	);
	LUT4 #(
		.INIT('ha800)
	) name3938 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6950_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3939 (
		\wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6951_
	);
	LUT3 #(
		.INIT('hf4)
	) name3940 (
		_w6949_,
		_w6950_,
		_w6951_,
		_w6952_
	);
	LUT4 #(
		.INIT('h8020)
	) name3941 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		\configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6953_
	);
	LUT4 #(
		.INIT('h8020)
	) name3942 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		\configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w6954_
	);
	LUT2 #(
		.INIT('h1)
	) name3943 (
		_w6953_,
		_w6954_,
		_w6955_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3944 (
		\wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w6956_
	);
	LUT3 #(
		.INIT('hf2)
	) name3945 (
		_w6950_,
		_w6955_,
		_w6956_,
		_w6957_
	);
	LUT4 #(
		.INIT('h2000)
	) name3946 (
		\output_backup_devsel_out_reg/NET0131 ,
		\output_backup_stop_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		_w6958_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w3224_,
		_w6958_,
		_w6959_
	);
	LUT4 #(
		.INIT('h0075)
	) name3948 (
		_w3212_,
		_w3215_,
		_w3221_,
		_w6959_,
		_w6960_
	);
	LUT4 #(
		.INIT('h0100)
	) name3949 (
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_request_reg/NET0131 ,
		_w6961_
	);
	LUT2 #(
		.INIT('h4)
	) name3950 (
		_w6960_,
		_w6961_,
		_w6962_
	);
	LUT3 #(
		.INIT('hca)
	) name3951 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]/P0001 ,
		_w6550_,
		_w6557_,
		_w6963_
	);
	LUT3 #(
		.INIT('hca)
	) name3952 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]/P0001 ,
		_w6550_,
		_w6553_,
		_w6964_
	);
	LUT3 #(
		.INIT('hca)
	) name3953 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]/P0001 ,
		_w6550_,
		_w6560_,
		_w6965_
	);
	LUT3 #(
		.INIT('hca)
	) name3954 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]/P0001 ,
		_w6550_,
		_w6563_,
		_w6966_
	);
	LUT3 #(
		.INIT('hca)
	) name3955 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]/P0001 ,
		_w6550_,
		_w6566_,
		_w6967_
	);
	LUT3 #(
		.INIT('hca)
	) name3956 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]/P0001 ,
		_w6550_,
		_w6569_,
		_w6968_
	);
	LUT3 #(
		.INIT('hca)
	) name3957 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]/P0001 ,
		_w6550_,
		_w6572_,
		_w6969_
	);
	LUT3 #(
		.INIT('hca)
	) name3958 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]/P0001 ,
		_w6550_,
		_w6575_,
		_w6970_
	);
	LUT3 #(
		.INIT('hca)
	) name3959 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]/P0001 ,
		_w6550_,
		_w6578_,
		_w6971_
	);
	LUT3 #(
		.INIT('hca)
	) name3960 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]/P0001 ,
		_w6550_,
		_w6581_,
		_w6972_
	);
	LUT3 #(
		.INIT('hca)
	) name3961 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]/P0001 ,
		_w6550_,
		_w6584_,
		_w6973_
	);
	LUT4 #(
		.INIT('h2111)
	) name3962 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]/NET0131 ,
		_w6313_,
		_w6742_,
		_w6754_,
		_w6974_
	);
	LUT2 #(
		.INIT('h4)
	) name3963 (
		\configuration_latency_timer_reg[3]/NET0131 ,
		_w6313_,
		_w6975_
	);
	LUT2 #(
		.INIT('h1)
	) name3964 (
		_w6974_,
		_w6975_,
		_w6976_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name3965 (
		\wishbone_slave_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_done_reg_main_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131 ,
		_w6977_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w6844_,
		_w6977_,
		_w6978_
	);
	LUT4 #(
		.INIT('h0080)
	) name3967 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w6979_
	);
	LUT3 #(
		.INIT('hca)
	) name3968 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]/P0001 ,
		_w6550_,
		_w6979_,
		_w6980_
	);
	LUT3 #(
		.INIT('hca)
	) name3969 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]/P0001 ,
		_w6550_,
		_w6590_,
		_w6981_
	);
	LUT3 #(
		.INIT('hca)
	) name3970 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]/P0001 ,
		_w6550_,
		_w6592_,
		_w6982_
	);
	LUT3 #(
		.INIT('hca)
	) name3971 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]/P0001 ,
		_w6550_,
		_w6594_,
		_w6983_
	);
	LUT3 #(
		.INIT('hca)
	) name3972 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]/P0001 ,
		_w6550_,
		_w6596_,
		_w6984_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3973 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[11]/NET0131 ,
		_w6511_,
		_w6518_,
		_w6985_
	);
	LUT4 #(
		.INIT('h8000)
	) name3974 (
		_w3053_,
		_w3055_,
		_w3050_,
		_w3093_,
		_w6986_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name3975 (
		\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131 ,
		_w6987_
	);
	LUT4 #(
		.INIT('h0001)
	) name3976 (
		\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131 ,
		\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]/NET0131 ,
		_w6988_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		_w6987_,
		_w6988_,
		_w6989_
	);
	LUT4 #(
		.INIT('h5700)
	) name3978 (
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131 ,
		_w6986_,
		_w6989_,
		_w6990_
	);
	LUT4 #(
		.INIT('hee0f)
	) name3979 (
		\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w6991_
	);
	LUT4 #(
		.INIT('h11f0)
	) name3980 (
		\wishbone_slave_unit_del_sync_be_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_data_source_reg/NET0131 ,
		_w6992_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w6991_,
		_w6993_
	);
	LUT3 #(
		.INIT('h40)
	) name3982 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001 ,
		_w3018_,
		_w3019_,
		_w6994_
	);
	LUT4 #(
		.INIT('h5444)
	) name3983 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131 ,
		_w3018_,
		_w3019_,
		_w6995_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3984 (
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w6993_,
		_w6994_,
		_w6995_,
		_w6996_
	);
	LUT4 #(
		.INIT('hff53)
	) name3985 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_be_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]/NET0131 ,
		_w6997_
	);
	LUT2 #(
		.INIT('hb)
	) name3986 (
		_w6996_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h4)
	) name3987 (
		\pci_target_unit_del_sync_comp_done_reg_clr_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_done_reg_main_reg/NET0131 ,
		_w6999_
	);
	LUT3 #(
		.INIT('h15)
	) name3988 (
		\pci_target_unit_del_sync_comp_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_wishbone_master_wb_read_done_out_reg/NET0131 ,
		_w7000_
	);
	LUT2 #(
		.INIT('h1)
	) name3989 (
		_w6999_,
		_w7000_,
		_w7001_
	);
	LUT4 #(
		.INIT('h2700)
	) name3990 (
		\output_backup_trdy_en_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		pci_trdy_i_pad,
		\wishbone_slave_unit_del_sync_burst_out_reg/NET0131 ,
		_w7002_
	);
	LUT3 #(
		.INIT('h2a)
	) name3991 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7003_
	);
	LUT3 #(
		.INIT('hd5)
	) name3992 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7004_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131 ,
		_w7005_
	);
	LUT3 #(
		.INIT('h01)
	) name3994 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131 ,
		_w7006_
	);
	LUT4 #(
		.INIT('hd555)
	) name3995 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7006_,
		_w7007_
	);
	LUT2 #(
		.INIT('h2)
	) name3996 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131 ,
		_w7007_,
		_w7008_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[3]/NET0131 ,
		_w7009_
	);
	LUT4 #(
		.INIT('h8000)
	) name3998 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7009_,
		_w7010_
	);
	LUT4 #(
		.INIT('h0001)
	) name3999 (
		\configuration_cache_line_size_reg_reg[4]/NET0131 ,
		\configuration_cache_line_size_reg_reg[5]/NET0131 ,
		\configuration_cache_line_size_reg_reg[6]/NET0131 ,
		\configuration_cache_line_size_reg_reg[7]/NET0131 ,
		_w7011_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name4000 (
		\configuration_cache_line_size_reg_reg[3]/NET0131 ,
		\wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w7011_,
		_w7012_
	);
	LUT3 #(
		.INIT('h07)
	) name4001 (
		_w7005_,
		_w7010_,
		_w7012_,
		_w7013_
	);
	LUT2 #(
		.INIT('hb)
	) name4002 (
		_w7008_,
		_w7013_,
		_w7014_
	);
	LUT4 #(
		.INIT('h001f)
	) name4003 (
		_w3140_,
		_w3135_,
		_w3143_,
		_w3158_,
		_w7015_
	);
	LUT4 #(
		.INIT('h8008)
	) name4004 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		\configuration_wb_ba2_bit0_reg/NET0131 ,
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w7016_
	);
	LUT4 #(
		.INIT('h8008)
	) name4005 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\configuration_wb_ba1_bit0_reg/NET0131 ,
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]/NET0131 ,
		_w7017_
	);
	LUT2 #(
		.INIT('h1)
	) name4006 (
		_w7016_,
		_w7017_,
		_w7018_
	);
	LUT4 #(
		.INIT('h00e0)
	) name4007 (
		_w3140_,
		_w3135_,
		_w3664_,
		_w7018_,
		_w7019_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4008 (
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		_w3140_,
		_w3135_,
		_w3664_,
		_w7020_
	);
	LUT2 #(
		.INIT('he)
	) name4009 (
		_w7019_,
		_w7020_,
		_w7021_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4010 (
		\pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg/NET0131 ,
		_w3234_,
		_w3235_,
		_w3236_,
		_w7022_
	);
	LUT3 #(
		.INIT('h40)
	) name4011 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7023_
	);
	LUT2 #(
		.INIT('h8)
	) name4012 (
		_w7022_,
		_w7023_,
		_w7024_
	);
	LUT3 #(
		.INIT('h10)
	) name4013 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7025_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		_w7022_,
		_w7025_,
		_w7026_
	);
	LUT3 #(
		.INIT('h20)
	) name4015 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7027_
	);
	LUT2 #(
		.INIT('h8)
	) name4016 (
		_w7022_,
		_w7027_,
		_w7028_
	);
	LUT3 #(
		.INIT('h80)
	) name4017 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7029_
	);
	LUT2 #(
		.INIT('h8)
	) name4018 (
		_w7022_,
		_w7029_,
		_w7030_
	);
	LUT3 #(
		.INIT('h04)
	) name4019 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7031_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		_w7022_,
		_w7031_,
		_w7032_
	);
	LUT3 #(
		.INIT('h01)
	) name4021 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7033_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		_w7022_,
		_w7033_,
		_w7034_
	);
	LUT3 #(
		.INIT('h02)
	) name4023 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7035_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		_w7022_,
		_w7035_,
		_w7036_
	);
	LUT3 #(
		.INIT('h08)
	) name4025 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7037_
	);
	LUT2 #(
		.INIT('h8)
	) name4026 (
		_w7022_,
		_w7037_,
		_w7038_
	);
	LUT3 #(
		.INIT('h1e)
	) name4027 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131 ,
		_w7039_
	);
	LUT4 #(
		.INIT('h0080)
	) name4028 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7039_,
		_w7040_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name4029 (
		\configuration_cache_line_size_reg_reg[2]/NET0131 ,
		\wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w7011_,
		_w7041_
	);
	LUT4 #(
		.INIT('hf8fb)
	) name4030 (
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]/NET0131 ,
		_w7003_,
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT3 #(
		.INIT('h60)
	) name4031 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[7]/NET0131 ,
		_w6509_,
		_w6518_,
		_w7043_
	);
	LUT3 #(
		.INIT('h10)
	) name4032 (
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		_w3044_,
		_w3046_,
		_w7044_
	);
	LUT3 #(
		.INIT('h80)
	) name4033 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w7045_
	);
	LUT2 #(
		.INIT('h8)
	) name4034 (
		_w3956_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4035 (
		\configuration_icr_bit31_reg/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7044_,
		_w7046_,
		_w7047_
	);
	LUT3 #(
		.INIT('h80)
	) name4036 (
		_w3782_,
		_w7044_,
		_w7046_,
		_w7048_
	);
	LUT2 #(
		.INIT('he)
	) name4037 (
		_w7047_,
		_w7048_,
		_w7049_
	);
	LUT4 #(
		.INIT('h2000)
	) name4038 (
		_w3040_,
		_w3044_,
		_w3046_,
		_w3806_,
		_w7050_
	);
	LUT2 #(
		.INIT('h2)
	) name4039 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7051_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4040 (
		\configuration_pci_ba1_bit31_8_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7052_
	);
	LUT2 #(
		.INIT('h2)
	) name4041 (
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7053_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4042 (
		\configuration_pci_ba1_bit31_8_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7054_
	);
	LUT2 #(
		.INIT('h2)
	) name4043 (
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7055_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4044 (
		\configuration_pci_ba1_bit31_8_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7056_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4045 (
		\configuration_icr_bit2_0_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7044_,
		_w7046_,
		_w7057_
	);
	LUT2 #(
		.INIT('h2)
	) name4046 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7058_
	);
	LUT3 #(
		.INIT('h80)
	) name4047 (
		_w7044_,
		_w7046_,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('he)
	) name4048 (
		_w7057_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('h2)
	) name4049 (
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7061_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4050 (
		\configuration_pci_ba1_bit31_8_reg[22]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7062_
	);
	LUT2 #(
		.INIT('h2)
	) name4051 (
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7063_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4052 (
		\configuration_pci_ba1_bit31_8_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7064_
	);
	LUT2 #(
		.INIT('h2)
	) name4053 (
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7065_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4054 (
		\configuration_pci_ba1_bit31_8_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7066_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4055 (
		\configuration_icr_bit2_0_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7044_,
		_w7046_,
		_w7067_
	);
	LUT2 #(
		.INIT('h2)
	) name4056 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7068_
	);
	LUT3 #(
		.INIT('h80)
	) name4057 (
		_w7044_,
		_w7046_,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('he)
	) name4058 (
		_w7067_,
		_w7069_,
		_w7070_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4059 (
		\configuration_pci_ba1_bit31_8_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7071_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4060 (
		\configuration_icr_bit2_0_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7044_,
		_w7046_,
		_w7072_
	);
	LUT2 #(
		.INIT('h2)
	) name4061 (
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7073_
	);
	LUT3 #(
		.INIT('h80)
	) name4062 (
		_w7044_,
		_w7046_,
		_w7073_,
		_w7074_
	);
	LUT2 #(
		.INIT('he)
	) name4063 (
		_w7072_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4064 (
		\configuration_pci_ba1_bit31_8_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7076_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4065 (
		\configuration_pci_ba1_bit31_8_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7077_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4066 (
		\configuration_pci_ba1_bit31_8_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7078_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4067 (
		\configuration_pci_ba1_bit31_8_reg[28]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7079_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4068 (
		\configuration_pci_ba1_bit31_8_reg[29]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7080_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4069 (
		\configuration_pci_ba1_bit31_8_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7081_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4070 (
		\configuration_pci_ba1_bit31_8_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7050_,
		_w7082_
	);
	LUT2 #(
		.INIT('h2)
	) name4071 (
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7083_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4072 (
		\configuration_pci_ba1_bit31_8_reg[9]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7084_
	);
	LUT2 #(
		.INIT('h2)
	) name4073 (
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7085_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4074 (
		\configuration_pci_ba1_bit31_8_reg[8]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7086_
	);
	LUT2 #(
		.INIT('h2)
	) name4075 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		_w7087_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w7088_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		_w3955_,
		_w7088_,
		_w7089_
	);
	LUT4 #(
		.INIT('h4000)
	) name4078 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7044_,
		_w7087_,
		_w7089_,
		_w7090_
	);
	LUT4 #(
		.INIT('h8000)
	) name4079 (
		_w7044_,
		_w7058_,
		_w7087_,
		_w7089_,
		_w7091_
	);
	LUT3 #(
		.INIT('hf2)
	) name4080 (
		\configuration_wb_img_ctrl1_bit2_0_reg[0]/NET0131 ,
		_w7090_,
		_w7091_,
		_w7092_
	);
	LUT4 #(
		.INIT('h8000)
	) name4081 (
		_w7044_,
		_w7073_,
		_w7087_,
		_w7089_,
		_w7093_
	);
	LUT3 #(
		.INIT('hf2)
	) name4082 (
		\configuration_wb_img_ctrl1_bit2_0_reg[2]/NET0131 ,
		_w7090_,
		_w7093_,
		_w7094_
	);
	LUT4 #(
		.INIT('h8000)
	) name4083 (
		_w7044_,
		_w7068_,
		_w7087_,
		_w7089_,
		_w7095_
	);
	LUT3 #(
		.INIT('hf2)
	) name4084 (
		\configuration_wb_img_ctrl1_bit2_0_reg[1]/NET0131 ,
		_w7090_,
		_w7095_,
		_w7096_
	);
	LUT3 #(
		.INIT('h40)
	) name4085 (
		_w3044_,
		_w3046_,
		_w3957_,
		_w7097_
	);
	LUT3 #(
		.INIT('h04)
	) name4086 (
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w7098_
	);
	LUT3 #(
		.INIT('h40)
	) name4087 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7088_,
		_w7098_,
		_w7099_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4088 (
		\configuration_pci_img_ctrl1_bit2_1_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7097_,
		_w7099_,
		_w7100_
	);
	LUT3 #(
		.INIT('h80)
	) name4089 (
		_w7068_,
		_w7097_,
		_w7099_,
		_w7101_
	);
	LUT2 #(
		.INIT('he)
	) name4090 (
		_w7100_,
		_w7101_,
		_w7102_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4091 (
		\configuration_pci_img_ctrl1_bit2_1_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7097_,
		_w7099_,
		_w7103_
	);
	LUT3 #(
		.INIT('h80)
	) name4092 (
		_w7073_,
		_w7097_,
		_w7099_,
		_w7104_
	);
	LUT2 #(
		.INIT('he)
	) name4093 (
		_w7103_,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h2)
	) name4094 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7106_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4095 (
		\configuration_pci_ba1_bit31_8_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7107_
	);
	LUT2 #(
		.INIT('h2)
	) name4096 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7108_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4097 (
		\configuration_pci_ba1_bit31_8_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7109_
	);
	LUT2 #(
		.INIT('h2)
	) name4098 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7110_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4099 (
		\configuration_pci_ba1_bit31_8_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7111_
	);
	LUT2 #(
		.INIT('h2)
	) name4100 (
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7112_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4101 (
		\configuration_pci_ba1_bit31_8_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7113_
	);
	LUT2 #(
		.INIT('h2)
	) name4102 (
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7114_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4103 (
		\configuration_pci_ba1_bit31_8_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7115_
	);
	LUT2 #(
		.INIT('h2)
	) name4104 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7116_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4105 (
		\configuration_pci_ba1_bit31_8_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7050_,
		_w7117_
	);
	LUT2 #(
		.INIT('h2)
	) name4106 (
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7118_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4107 (
		\configuration_pci_ba1_bit31_8_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7119_
	);
	LUT2 #(
		.INIT('h2)
	) name4108 (
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7120_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4109 (
		\configuration_pci_ba1_bit31_8_reg[17]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7050_,
		_w7121_
	);
	LUT4 #(
		.INIT('h8000)
	) name4110 (
		_w3052_,
		_w3053_,
		_w3055_,
		_w3068_,
		_w7122_
	);
	LUT2 #(
		.INIT('he)
	) name4111 (
		_w3069_,
		_w7122_,
		_w7123_
	);
	LUT4 #(
		.INIT('h8880)
	) name4112 (
		\configuration_icr_bit2_0_reg[2]/NET0131 ,
		\configuration_pci_err_cs_bit0_reg/NET0131 ,
		_w3069_,
		_w7122_,
		_w7124_
	);
	LUT3 #(
		.INIT('h8a)
	) name4113 (
		\configuration_set_isr_bit2_reg/NET0131 ,
		\configuration_sync_isr_2_delayed_del_bit_reg/NET0131 ,
		\configuration_sync_isr_2_sync_del_bit_reg/NET0131 ,
		_w7125_
	);
	LUT2 #(
		.INIT('he)
	) name4114 (
		_w7124_,
		_w7125_,
		_w7126_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4115 (
		\wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]/P0001 ,
		_w3027_,
		_w3029_,
		_w7127_
	);
	LUT4 #(
		.INIT('h0600)
	) name4116 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[3]/NET0131 ,
		_w6505_,
		_w6516_,
		_w6517_,
		_w7128_
	);
	LUT3 #(
		.INIT('h60)
	) name4117 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[10]/NET0131 ,
		_w6511_,
		_w6518_,
		_w7129_
	);
	LUT3 #(
		.INIT('h2a)
	) name4118 (
		\configuration_pci_err_cs_bit10_reg/NET0131 ,
		_w3060_,
		_w3068_,
		_w7130_
	);
	LUT2 #(
		.INIT('he)
	) name4119 (
		_w7122_,
		_w7130_,
		_w7131_
	);
	LUT4 #(
		.INIT('h0888)
	) name4120 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_bound_reg/NET0131 ,
		_w3019_,
		_w7002_,
		_w7132_
	);
	LUT2 #(
		.INIT('he)
	) name4121 (
		_w7010_,
		_w7132_,
		_w7133_
	);
	LUT3 #(
		.INIT('h2a)
	) name4122 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		_w3131_,
		_w3133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		\wbs_adr_i[2]_pad ,
		\wbs_adr_i[3]_pad ,
		_w7135_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4124 (
		\wbs_adr_i[2]_pad ,
		\wbs_adr_i[3]_pad ,
		\wbs_adr_i[4]_pad ,
		\wbs_bte_i[1]_pad ,
		_w7136_
	);
	LUT3 #(
		.INIT('he0)
	) name4125 (
		\wbs_adr_i[4]_pad ,
		\wbs_adr_i[5]_pad ,
		\wbs_bte_i[1]_pad ,
		_w7137_
	);
	LUT4 #(
		.INIT('hfa32)
	) name4126 (
		\wbs_bte_i[0]_pad ,
		_w7135_,
		_w7136_,
		_w7137_,
		_w7138_
	);
	LUT3 #(
		.INIT('h04)
	) name4127 (
		\wbs_cti_i[0]_pad ,
		\wbs_cti_i[1]_pad ,
		\wbs_cti_i[2]_pad ,
		_w7139_
	);
	LUT3 #(
		.INIT('h80)
	) name4128 (
		_w3131_,
		_w3133_,
		_w7139_,
		_w7140_
	);
	LUT3 #(
		.INIT('hba)
	) name4129 (
		_w7134_,
		_w7138_,
		_w7140_,
		_w7141_
	);
	LUT3 #(
		.INIT('h8a)
	) name4130 (
		\configuration_set_pci_err_cs_bit8_reg/NET0131 ,
		\configuration_sync_pci_err_cs_8_delayed_del_bit_reg/NET0131 ,
		\configuration_sync_pci_err_cs_8_sync_del_bit_reg/NET0131 ,
		_w7142_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4131 (
		\configuration_pci_err_cs_bit0_reg/NET0131 ,
		_w3069_,
		_w7122_,
		_w7142_,
		_w7143_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name4132 (
		\wishbone_slave_unit_pci_initiator_if_last_transfered_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6833_,
		_w7144_
	);
	LUT3 #(
		.INIT('hf4)
	) name4133 (
		_w3027_,
		_w3029_,
		_w7144_,
		_w7145_
	);
	LUT3 #(
		.INIT('h10)
	) name4134 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3044_,
		_w3046_,
		_w7146_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4135 (
		\configuration_wb_ta1_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w3819_,
		_w7146_,
		_w7147_
	);
	LUT3 #(
		.INIT('h10)
	) name4136 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3044_,
		_w3046_,
		_w7148_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4137 (
		\configuration_pci_err_cs_bit0_reg/NET0131 ,
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		_w3841_,
		_w7148_,
		_w7149_
	);
	LUT4 #(
		.INIT('h4000)
	) name4138 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		_w7044_,
		_w7089_,
		_w7150_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4139 (
		\configuration_wb_ba1_bit0_reg/NET0131 ,
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h4)
	) name4140 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7152_
	);
	LUT4 #(
		.INIT('h8000)
	) name4141 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		_w7044_,
		_w7089_,
		_w7152_,
		_w7153_
	);
	LUT3 #(
		.INIT('hca)
	) name4142 (
		\configuration_wb_am1_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h8)
	) name4143 (
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		_w7155_
	);
	LUT3 #(
		.INIT('h40)
	) name4144 (
		_w3044_,
		_w3046_,
		_w7155_,
		_w7156_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4145 (
		\configuration_wb_am2_reg[31]/NET0131 ,
		_w7089_,
		_w7152_,
		_w7156_,
		_w7157_
	);
	LUT4 #(
		.INIT('h8000)
	) name4146 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w7089_,
		_w7152_,
		_w7156_,
		_w7158_
	);
	LUT2 #(
		.INIT('he)
	) name4147 (
		_w7157_,
		_w7158_,
		_w7159_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4148 (
		\configuration_wb_ba1_bit31_12_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7150_,
		_w7160_
	);
	LUT4 #(
		.INIT('h1000)
	) name4149 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7089_,
		_w7156_,
		_w7161_
	);
	LUT4 #(
		.INIT('h4000)
	) name4150 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7058_,
		_w7089_,
		_w7156_,
		_w7162_
	);
	LUT3 #(
		.INIT('hf2)
	) name4151 (
		\configuration_wb_ba2_bit0_reg/NET0131 ,
		_w7161_,
		_w7162_,
		_w7163_
	);
	LUT4 #(
		.INIT('h1000)
	) name4152 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7089_,
		_w7156_,
		_w7164_
	);
	LUT4 #(
		.INIT('h4000)
	) name4153 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w3782_,
		_w7089_,
		_w7156_,
		_w7165_
	);
	LUT3 #(
		.INIT('hf2)
	) name4154 (
		\configuration_wb_ba2_bit31_12_reg[31]/NET0131 ,
		_w7164_,
		_w7165_,
		_w7166_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4155 (
		\configuration_command_bit8_reg/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7167_
	);
	LUT3 #(
		.INIT('h80)
	) name4156 (
		_w3043_,
		_w3047_,
		_w7085_,
		_w7168_
	);
	LUT2 #(
		.INIT('he)
	) name4157 (
		_w7167_,
		_w7168_,
		_w7169_
	);
	LUT3 #(
		.INIT('h20)
	) name4158 (
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w7170_
	);
	LUT3 #(
		.INIT('h80)
	) name4159 (
		_w3955_,
		_w7087_,
		_w7170_,
		_w7171_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4160 (
		\configuration_wb_err_cs_bit0_reg/NET0131 ,
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		_w7148_,
		_w7171_,
		_w7172_
	);
	LUT4 #(
		.INIT('h0001)
	) name4161 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w7173_
	);
	LUT2 #(
		.INIT('h8)
	) name4162 (
		_w3956_,
		_w7173_,
		_w7174_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4163 (
		\configuration_wb_ta2_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		_w7044_,
		_w7174_,
		_w7175_
	);
	LUT4 #(
		.INIT('h333a)
	) name4164 (
		\configuration_pci_err_cs_bit31_24_reg[28]/NET0131 ,
		\wbm_sel_o[0]_pad ,
		_w3069_,
		_w7122_,
		_w7176_
	);
	LUT4 #(
		.INIT('h333a)
	) name4165 (
		\configuration_pci_err_cs_bit31_24_reg[29]/NET0131 ,
		\wbm_sel_o[1]_pad ,
		_w3069_,
		_w7122_,
		_w7177_
	);
	LUT4 #(
		.INIT('h333a)
	) name4166 (
		\configuration_pci_err_cs_bit31_24_reg[30]/NET0131 ,
		\wbm_sel_o[2]_pad ,
		_w3069_,
		_w7122_,
		_w7178_
	);
	LUT4 #(
		.INIT('h333a)
	) name4167 (
		\configuration_pci_err_cs_bit31_24_reg[31]/NET0131 ,
		\wbm_sel_o[3]_pad ,
		_w3069_,
		_w7122_,
		_w7179_
	);
	LUT2 #(
		.INIT('h4)
	) name4168 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 ,
		_w7180_
	);
	LUT3 #(
		.INIT('h08)
	) name4169 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6833_,
		_w7181_
	);
	LUT3 #(
		.INIT('h01)
	) name4170 (
		\wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_err_recovery_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_intermediate_last_reg/NET0131 ,
		_w7182_
	);
	LUT4 #(
		.INIT('h0800)
	) name4171 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6833_,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('he)
	) name4172 (
		_w7180_,
		_w7183_,
		_w7184_
	);
	LUT3 #(
		.INIT('hca)
	) name4173 (
		\configuration_wb_err_addr_reg[0]/NET0131 ,
		_w4937_,
		_w7181_,
		_w7185_
	);
	LUT4 #(
		.INIT('h1000)
	) name4174 (
		\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_read_count_reg[1]/NET0131 ,
		_w3057_,
		_w3050_,
		_w7186_
	);
	LUT4 #(
		.INIT('h6333)
	) name4175 (
		\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_read_count_reg[1]/NET0131 ,
		_w3057_,
		_w3050_,
		_w7187_
	);
	LUT3 #(
		.INIT('h01)
	) name4176 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[5]/NET0131 ,
		\configuration_sync_cache_lsize_to_wb_bits_reg[6]/NET0131 ,
		\configuration_sync_cache_lsize_to_wb_bits_reg[7]/NET0131 ,
		_w7188_
	);
	LUT4 #(
		.INIT('h1110)
	) name4177 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[3]/NET0131 ,
		\configuration_sync_cache_lsize_to_wb_bits_reg[4]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[1]/NET0131 ,
		_w7189_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT4 #(
		.INIT('h038b)
	) name4179 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 ,
		_w3085_,
		_w7187_,
		_w7190_,
		_w7191_
	);
	LUT3 #(
		.INIT('h80)
	) name4180 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7088_,
		_w7098_,
		_w7192_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4181 (
		\configuration_pci_ta1_reg[19]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7193_
	);
	LUT3 #(
		.INIT('h80)
	) name4182 (
		_w7053_,
		_w7156_,
		_w7192_,
		_w7194_
	);
	LUT2 #(
		.INIT('he)
	) name4183 (
		_w7193_,
		_w7194_,
		_w7195_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4184 (
		\configuration_pci_ta1_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7196_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7197_
	);
	LUT3 #(
		.INIT('h80)
	) name4186 (
		_w7156_,
		_w7192_,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('he)
	) name4187 (
		_w7196_,
		_w7198_,
		_w7199_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4188 (
		\configuration_interrupt_line_reg[0]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7200_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4189 (
		\configuration_interrupt_line_reg[1]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7201_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4190 (
		\configuration_interrupt_line_reg[2]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7202_
	);
	LUT3 #(
		.INIT('h80)
	) name4191 (
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w3955_,
		_w7088_,
		_w7203_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4192 (
		\configuration_wb_img_ctrl2_bit2_0_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7097_,
		_w7203_,
		_w7204_
	);
	LUT3 #(
		.INIT('h80)
	) name4193 (
		_w7058_,
		_w7097_,
		_w7203_,
		_w7205_
	);
	LUT2 #(
		.INIT('he)
	) name4194 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4195 (
		\configuration_wb_img_ctrl2_bit2_0_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7097_,
		_w7203_,
		_w7207_
	);
	LUT3 #(
		.INIT('h80)
	) name4196 (
		_w7068_,
		_w7097_,
		_w7203_,
		_w7208_
	);
	LUT2 #(
		.INIT('he)
	) name4197 (
		_w7207_,
		_w7208_,
		_w7209_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4198 (
		\configuration_wb_img_ctrl2_bit2_0_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w7097_,
		_w7203_,
		_w7210_
	);
	LUT3 #(
		.INIT('h80)
	) name4199 (
		_w7073_,
		_w7097_,
		_w7203_,
		_w7211_
	);
	LUT2 #(
		.INIT('he)
	) name4200 (
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4201 (
		\configuration_interrupt_line_reg[6]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7213_
	);
	LUT4 #(
		.INIT('h4000)
	) name4202 (
		_w3044_,
		_w3046_,
		_w3824_,
		_w3807_,
		_w7214_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4203 (
		\configuration_pci_am1_reg[29]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7215_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4204 (
		\configuration_latency_timer_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7216_
	);
	LUT3 #(
		.INIT('h80)
	) name4205 (
		_w3047_,
		_w3948_,
		_w7085_,
		_w7217_
	);
	LUT2 #(
		.INIT('he)
	) name4206 (
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4207 (
		\configuration_latency_timer_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7219_
	);
	LUT3 #(
		.INIT('h80)
	) name4208 (
		_w3047_,
		_w3948_,
		_w7083_,
		_w7220_
	);
	LUT2 #(
		.INIT('he)
	) name4209 (
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4210 (
		\configuration_latency_timer_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7222_
	);
	LUT3 #(
		.INIT('h80)
	) name4211 (
		_w3047_,
		_w3948_,
		_w7106_,
		_w7223_
	);
	LUT2 #(
		.INIT('he)
	) name4212 (
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4213 (
		\configuration_pci_am1_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7225_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4214 (
		\configuration_latency_timer_reg[3]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7226_
	);
	LUT3 #(
		.INIT('h80)
	) name4215 (
		_w3047_,
		_w3948_,
		_w7108_,
		_w7227_
	);
	LUT2 #(
		.INIT('he)
	) name4216 (
		_w7226_,
		_w7227_,
		_w7228_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4217 (
		\configuration_pci_ba0_bit31_8_reg[16]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7229_
	);
	LUT3 #(
		.INIT('h20)
	) name4218 (
		_w3047_,
		_w3831_,
		_w7118_,
		_w7230_
	);
	LUT2 #(
		.INIT('he)
	) name4219 (
		_w7229_,
		_w7230_,
		_w7231_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4220 (
		\configuration_latency_timer_reg[4]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7232_
	);
	LUT3 #(
		.INIT('h80)
	) name4221 (
		_w3047_,
		_w3948_,
		_w7110_,
		_w7233_
	);
	LUT2 #(
		.INIT('he)
	) name4222 (
		_w7232_,
		_w7233_,
		_w7234_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4223 (
		\configuration_pci_am1_reg[8]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7235_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4224 (
		\configuration_latency_timer_reg[5]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7236_
	);
	LUT3 #(
		.INIT('h80)
	) name4225 (
		_w3047_,
		_w3948_,
		_w7112_,
		_w7237_
	);
	LUT2 #(
		.INIT('he)
	) name4226 (
		_w7236_,
		_w7237_,
		_w7238_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4227 (
		\configuration_pci_am1_reg[22]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7239_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4228 (
		\configuration_latency_timer_reg[6]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7240_
	);
	LUT3 #(
		.INIT('h80)
	) name4229 (
		_w3047_,
		_w3948_,
		_w7114_,
		_w7241_
	);
	LUT2 #(
		.INIT('he)
	) name4230 (
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4231 (
		\configuration_pci_am1_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7243_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4232 (
		\configuration_latency_timer_reg[7]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3948_,
		_w7244_
	);
	LUT3 #(
		.INIT('h80)
	) name4233 (
		_w3047_,
		_w3948_,
		_w7116_,
		_w7245_
	);
	LUT2 #(
		.INIT('he)
	) name4234 (
		_w7244_,
		_w7245_,
		_w7246_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4235 (
		\configuration_cache_line_size_reg_reg[0]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7247_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4236 (
		\configuration_pci_am1_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7248_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4237 (
		\configuration_pci_ta1_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7249_
	);
	LUT2 #(
		.INIT('h2)
	) name4238 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7250_
	);
	LUT3 #(
		.INIT('h80)
	) name4239 (
		_w7156_,
		_w7192_,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('he)
	) name4240 (
		_w7249_,
		_w7251_,
		_w7252_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4241 (
		\configuration_pci_am1_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7253_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4242 (
		\configuration_pci_am1_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7254_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4243 (
		\configuration_pci_am1_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7255_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4244 (
		\configuration_pci_am1_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7256_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4245 (
		\configuration_pci_am1_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7257_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4246 (
		\configuration_pci_am1_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7258_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4247 (
		\configuration_pci_ta1_reg[10]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7259_
	);
	LUT3 #(
		.INIT('h80)
	) name4248 (
		_w7106_,
		_w7156_,
		_w7192_,
		_w7260_
	);
	LUT2 #(
		.INIT('he)
	) name4249 (
		_w7259_,
		_w7260_,
		_w7261_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4250 (
		\configuration_pci_am1_reg[17]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7262_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4251 (
		\configuration_pci_am1_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7263_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4252 (
		\configuration_pci_am1_reg[20]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7264_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4253 (
		\configuration_pci_ta1_reg[11]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7265_
	);
	LUT3 #(
		.INIT('h80)
	) name4254 (
		_w7108_,
		_w7156_,
		_w7192_,
		_w7266_
	);
	LUT2 #(
		.INIT('he)
	) name4255 (
		_w7265_,
		_w7266_,
		_w7267_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4256 (
		\configuration_pci_ta1_reg[12]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7268_
	);
	LUT3 #(
		.INIT('h80)
	) name4257 (
		_w7110_,
		_w7156_,
		_w7192_,
		_w7269_
	);
	LUT2 #(
		.INIT('he)
	) name4258 (
		_w7268_,
		_w7269_,
		_w7270_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4259 (
		\configuration_pci_ta1_reg[13]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7271_
	);
	LUT3 #(
		.INIT('h80)
	) name4260 (
		_w7112_,
		_w7156_,
		_w7192_,
		_w7272_
	);
	LUT2 #(
		.INIT('he)
	) name4261 (
		_w7271_,
		_w7272_,
		_w7273_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4262 (
		\configuration_pci_ta1_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7274_
	);
	LUT3 #(
		.INIT('h80)
	) name4263 (
		_w7114_,
		_w7156_,
		_w7192_,
		_w7275_
	);
	LUT2 #(
		.INIT('he)
	) name4264 (
		_w7274_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4265 (
		\configuration_pci_am1_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7277_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4266 (
		\configuration_pci_ba0_bit31_8_reg[15]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7278_
	);
	LUT3 #(
		.INIT('h20)
	) name4267 (
		_w3047_,
		_w3831_,
		_w7116_,
		_w7279_
	);
	LUT2 #(
		.INIT('he)
	) name4268 (
		_w7278_,
		_w7279_,
		_w7280_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4269 (
		\configuration_pci_ta1_reg[16]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7281_
	);
	LUT3 #(
		.INIT('h80)
	) name4270 (
		_w7118_,
		_w7156_,
		_w7192_,
		_w7282_
	);
	LUT2 #(
		.INIT('he)
	) name4271 (
		_w7281_,
		_w7282_,
		_w7283_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4272 (
		\configuration_pci_ta1_reg[17]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7284_
	);
	LUT3 #(
		.INIT('h80)
	) name4273 (
		_w7120_,
		_w7156_,
		_w7192_,
		_w7285_
	);
	LUT2 #(
		.INIT('he)
	) name4274 (
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4275 (
		\configuration_pci_ta1_reg[18]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7287_
	);
	LUT3 #(
		.INIT('h80)
	) name4276 (
		_w7051_,
		_w7156_,
		_w7192_,
		_w7288_
	);
	LUT2 #(
		.INIT('he)
	) name4277 (
		_w7287_,
		_w7288_,
		_w7289_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4278 (
		\configuration_pci_am1_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7290_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4279 (
		\configuration_pci_ta1_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7291_
	);
	LUT3 #(
		.INIT('h80)
	) name4280 (
		_w7055_,
		_w7156_,
		_w7192_,
		_w7292_
	);
	LUT2 #(
		.INIT('he)
	) name4281 (
		_w7291_,
		_w7292_,
		_w7293_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4282 (
		\configuration_pci_ta1_reg[21]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7294_
	);
	LUT3 #(
		.INIT('h80)
	) name4283 (
		_w7063_,
		_w7156_,
		_w7192_,
		_w7295_
	);
	LUT2 #(
		.INIT('he)
	) name4284 (
		_w7294_,
		_w7295_,
		_w7296_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4285 (
		\configuration_pci_ta1_reg[22]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7297_
	);
	LUT3 #(
		.INIT('h80)
	) name4286 (
		_w7061_,
		_w7156_,
		_w7192_,
		_w7298_
	);
	LUT2 #(
		.INIT('he)
	) name4287 (
		_w7297_,
		_w7298_,
		_w7299_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4288 (
		\configuration_cache_line_size_reg_reg[1]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7300_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4289 (
		\configuration_pci_am1_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7301_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4290 (
		\configuration_pci_ta1_reg[23]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7302_
	);
	LUT3 #(
		.INIT('h80)
	) name4291 (
		_w7065_,
		_w7156_,
		_w7192_,
		_w7303_
	);
	LUT2 #(
		.INIT('he)
	) name4292 (
		_w7302_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4293 (
		\configuration_pci_ta1_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7305_
	);
	LUT3 #(
		.INIT('h80)
	) name4294 (
		_w3038_,
		_w7156_,
		_w7192_,
		_w7306_
	);
	LUT2 #(
		.INIT('he)
	) name4295 (
		_w7305_,
		_w7306_,
		_w7307_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4296 (
		\configuration_pci_ta1_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7308_
	);
	LUT4 #(
		.INIT('h2000)
	) name4297 (
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7309_
	);
	LUT2 #(
		.INIT('he)
	) name4298 (
		_w7308_,
		_w7309_,
		_w7310_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4299 (
		\configuration_pci_am1_reg[25]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7311_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4300 (
		\configuration_pci_ta1_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7312_
	);
	LUT4 #(
		.INIT('h2000)
	) name4301 (
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7313_
	);
	LUT2 #(
		.INIT('he)
	) name4302 (
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4303 (
		\configuration_cache_line_size_reg_reg[2]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7315_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4304 (
		\configuration_pci_am1_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w7214_,
		_w7316_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4305 (
		\configuration_pci_am1_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7317_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4306 (
		\configuration_pci_ta1_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7318_
	);
	LUT3 #(
		.INIT('h80)
	) name4307 (
		_w3782_,
		_w7156_,
		_w7192_,
		_w7319_
	);
	LUT2 #(
		.INIT('he)
	) name4308 (
		_w7318_,
		_w7319_,
		_w7320_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4309 (
		\configuration_pci_ta1_reg[8]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7321_
	);
	LUT3 #(
		.INIT('h80)
	) name4310 (
		_w7085_,
		_w7156_,
		_w7192_,
		_w7322_
	);
	LUT2 #(
		.INIT('he)
	) name4311 (
		_w7321_,
		_w7322_,
		_w7323_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4312 (
		\configuration_pci_ta1_reg[9]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7324_
	);
	LUT3 #(
		.INIT('h80)
	) name4313 (
		_w7083_,
		_w7156_,
		_w7192_,
		_w7325_
	);
	LUT2 #(
		.INIT('he)
	) name4314 (
		_w7324_,
		_w7325_,
		_w7326_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4315 (
		\configuration_pci_am1_reg[28]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7327_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4316 (
		\configuration_pci_am1_reg[31]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7214_,
		_w7328_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4317 (
		\configuration_pci_am1_reg[9]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7214_,
		_w7329_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4318 (
		\configuration_pci_ba0_bit31_8_reg[12]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7330_
	);
	LUT3 #(
		.INIT('h20)
	) name4319 (
		_w3047_,
		_w3831_,
		_w7110_,
		_w7331_
	);
	LUT2 #(
		.INIT('he)
	) name4320 (
		_w7330_,
		_w7331_,
		_w7332_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4321 (
		\configuration_pci_ba0_bit31_8_reg[13]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7333_
	);
	LUT3 #(
		.INIT('h20)
	) name4322 (
		_w3047_,
		_w3831_,
		_w7112_,
		_w7334_
	);
	LUT2 #(
		.INIT('he)
	) name4323 (
		_w7333_,
		_w7334_,
		_w7335_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4324 (
		\configuration_pci_ba0_bit31_8_reg[14]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7336_
	);
	LUT3 #(
		.INIT('h20)
	) name4325 (
		_w3047_,
		_w3831_,
		_w7114_,
		_w7337_
	);
	LUT2 #(
		.INIT('he)
	) name4326 (
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4327 (
		\configuration_pci_ba0_bit31_8_reg[18]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7339_
	);
	LUT3 #(
		.INIT('h20)
	) name4328 (
		_w3047_,
		_w3831_,
		_w7051_,
		_w7340_
	);
	LUT2 #(
		.INIT('he)
	) name4329 (
		_w7339_,
		_w7340_,
		_w7341_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4330 (
		\configuration_cache_line_size_reg_reg[6]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7342_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4331 (
		\configuration_pci_ba0_bit31_8_reg[17]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7343_
	);
	LUT3 #(
		.INIT('h20)
	) name4332 (
		_w3047_,
		_w3831_,
		_w7120_,
		_w7344_
	);
	LUT2 #(
		.INIT('he)
	) name4333 (
		_w7343_,
		_w7344_,
		_w7345_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4334 (
		\configuration_pci_ba0_bit31_8_reg[19]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7346_
	);
	LUT3 #(
		.INIT('h20)
	) name4335 (
		_w3047_,
		_w3831_,
		_w7053_,
		_w7347_
	);
	LUT2 #(
		.INIT('he)
	) name4336 (
		_w7346_,
		_w7347_,
		_w7348_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4337 (
		\configuration_pci_ba0_bit31_8_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7349_
	);
	LUT3 #(
		.INIT('h20)
	) name4338 (
		_w3047_,
		_w3831_,
		_w7055_,
		_w7350_
	);
	LUT2 #(
		.INIT('he)
	) name4339 (
		_w7349_,
		_w7350_,
		_w7351_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4340 (
		\configuration_pci_ba0_bit31_8_reg[21]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7352_
	);
	LUT3 #(
		.INIT('h20)
	) name4341 (
		_w3047_,
		_w3831_,
		_w7063_,
		_w7353_
	);
	LUT2 #(
		.INIT('he)
	) name4342 (
		_w7352_,
		_w7353_,
		_w7354_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4343 (
		\configuration_pci_ba0_bit31_8_reg[22]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7355_
	);
	LUT3 #(
		.INIT('h20)
	) name4344 (
		_w3047_,
		_w3831_,
		_w7061_,
		_w7356_
	);
	LUT2 #(
		.INIT('he)
	) name4345 (
		_w7355_,
		_w7356_,
		_w7357_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4346 (
		\configuration_pci_ba0_bit31_8_reg[23]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7358_
	);
	LUT3 #(
		.INIT('h20)
	) name4347 (
		_w3047_,
		_w3831_,
		_w7065_,
		_w7359_
	);
	LUT2 #(
		.INIT('he)
	) name4348 (
		_w7358_,
		_w7359_,
		_w7360_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4349 (
		\configuration_pci_ba0_bit31_8_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7361_
	);
	LUT4 #(
		.INIT('h0020)
	) name4350 (
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7362_
	);
	LUT2 #(
		.INIT('he)
	) name4351 (
		_w7361_,
		_w7362_,
		_w7363_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4352 (
		\configuration_pci_ba0_bit31_8_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7364_
	);
	LUT4 #(
		.INIT('h0020)
	) name4353 (
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7365_
	);
	LUT2 #(
		.INIT('he)
	) name4354 (
		_w7364_,
		_w7365_,
		_w7366_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4355 (
		\configuration_command_bit2_0_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7367_
	);
	LUT3 #(
		.INIT('h80)
	) name4356 (
		_w3043_,
		_w3047_,
		_w7058_,
		_w7368_
	);
	LUT2 #(
		.INIT('he)
	) name4357 (
		_w7367_,
		_w7368_,
		_w7369_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4358 (
		\configuration_pci_ba0_bit31_8_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7370_
	);
	LUT4 #(
		.INIT('h0020)
	) name4359 (
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7371_
	);
	LUT2 #(
		.INIT('he)
	) name4360 (
		_w7370_,
		_w7371_,
		_w7372_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4361 (
		\configuration_pci_ba0_bit31_8_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7373_
	);
	LUT4 #(
		.INIT('h0020)
	) name4362 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7374_
	);
	LUT2 #(
		.INIT('he)
	) name4363 (
		_w7373_,
		_w7374_,
		_w7375_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4364 (
		\configuration_pci_ba0_bit31_8_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7376_
	);
	LUT4 #(
		.INIT('h0020)
	) name4365 (
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7377_
	);
	LUT2 #(
		.INIT('he)
	) name4366 (
		_w7376_,
		_w7377_,
		_w7378_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4367 (
		\configuration_pci_ba0_bit31_8_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7379_
	);
	LUT4 #(
		.INIT('h0020)
	) name4368 (
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7380_
	);
	LUT2 #(
		.INIT('he)
	) name4369 (
		_w7379_,
		_w7380_,
		_w7381_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4370 (
		\configuration_pci_ba0_bit31_8_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7382_
	);
	LUT4 #(
		.INIT('h0020)
	) name4371 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7383_
	);
	LUT2 #(
		.INIT('he)
	) name4372 (
		_w7382_,
		_w7383_,
		_w7384_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4373 (
		\configuration_command_bit2_0_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7385_
	);
	LUT4 #(
		.INIT('h2000)
	) name4374 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7386_
	);
	LUT2 #(
		.INIT('he)
	) name4375 (
		_w7385_,
		_w7386_,
		_w7387_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4376 (
		\configuration_pci_ba0_bit31_8_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7388_
	);
	LUT4 #(
		.INIT('h0020)
	) name4377 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w3047_,
		_w3831_,
		_w7389_
	);
	LUT2 #(
		.INIT('he)
	) name4378 (
		_w7388_,
		_w7389_,
		_w7390_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4379 (
		\configuration_command_bit2_0_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7391_
	);
	LUT4 #(
		.INIT('h2000)
	) name4380 (
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7392_
	);
	LUT2 #(
		.INIT('he)
	) name4381 (
		_w7391_,
		_w7392_,
		_w7393_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4382 (
		\configuration_command_bit6_reg/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7394_
	);
	LUT4 #(
		.INIT('h2000)
	) name4383 (
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7395_
	);
	LUT2 #(
		.INIT('he)
	) name4384 (
		_w7394_,
		_w7395_,
		_w7396_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4385 (
		\configuration_pci_ta1_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7397_
	);
	LUT2 #(
		.INIT('h2)
	) name4386 (
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7398_
	);
	LUT3 #(
		.INIT('h80)
	) name4387 (
		_w7156_,
		_w7192_,
		_w7398_,
		_w7399_
	);
	LUT2 #(
		.INIT('he)
	) name4388 (
		_w7397_,
		_w7399_,
		_w7400_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4389 (
		\configuration_pci_ta1_reg[15]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7401_
	);
	LUT3 #(
		.INIT('h80)
	) name4390 (
		_w7116_,
		_w7156_,
		_w7192_,
		_w7402_
	);
	LUT2 #(
		.INIT('he)
	) name4391 (
		_w7401_,
		_w7402_,
		_w7403_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4392 (
		\configuration_pci_ta1_reg[30]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		_w7156_,
		_w7192_,
		_w7404_
	);
	LUT3 #(
		.INIT('h80)
	) name4393 (
		_w4475_,
		_w7156_,
		_w7192_,
		_w7405_
	);
	LUT2 #(
		.INIT('he)
	) name4394 (
		_w7404_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h4)
	) name4395 (
		\configuration_latency_timer_reg[6]/NET0131 ,
		_w6313_,
		_w7407_
	);
	LUT4 #(
		.INIT('h0603)
	) name4396 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]/NET0131 ,
		_w6313_,
		_w6756_,
		_w7408_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w7407_,
		_w7408_,
		_w7409_
	);
	LUT4 #(
		.INIT('h0603)
	) name4398 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]/NET0131 ,
		_w6313_,
		_w6754_,
		_w7410_
	);
	LUT2 #(
		.INIT('h4)
	) name4399 (
		\configuration_latency_timer_reg[2]/NET0131 ,
		_w6313_,
		_w7411_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w7410_,
		_w7411_,
		_w7412_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name4401 (
		\configuration_latency_timer_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]/NET0131 ,
		_w6313_,
		_w6756_,
		_w7413_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name4402 (
		\configuration_latency_timer_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]/NET0131 ,
		_w6313_,
		_w6754_,
		_w7414_
	);
	LUT3 #(
		.INIT('h40)
	) name4403 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[2]/NET0131 ,
		_w7188_,
		_w7189_,
		_w7415_
	);
	LUT2 #(
		.INIT('h2)
	) name4404 (
		_w3086_,
		_w7415_,
		_w7416_
	);
	LUT3 #(
		.INIT('h12)
	) name4405 (
		\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131 ,
		_w3085_,
		_w7186_,
		_w7417_
	);
	LUT2 #(
		.INIT('he)
	) name4406 (
		_w7416_,
		_w7417_,
		_w7418_
	);
	LUT4 #(
		.INIT('ha3ac)
	) name4407 (
		\configuration_latency_timer_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]/NET0131 ,
		_w6313_,
		_w6755_,
		_w7419_
	);
	LUT2 #(
		.INIT('h4)
	) name4408 (
		\configuration_latency_timer_reg[0]/NET0131 ,
		_w6313_,
		_w7420_
	);
	LUT4 #(
		.INIT('h1222)
	) name4409 (
		\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]/NET0131 ,
		_w6313_,
		_w6740_,
		_w6743_,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name4410 (
		_w7420_,
		_w7421_,
		_w7422_
	);
	LUT3 #(
		.INIT('h95)
	) name4411 (
		\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 ,
		_w3057_,
		_w3050_,
		_w7423_
	);
	LUT4 #(
		.INIT('h4c7f)
	) name4412 (
		\configuration_sync_cache_lsize_to_wb_bits_reg[8]/NET0131 ,
		_w3085_,
		_w7190_,
		_w7423_,
		_w7424_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4413 (
		\configuration_status_bit15_11_reg[11]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7250_,
		_w7425_
	);
	LUT2 #(
		.INIT('he)
	) name4414 (
		_w6958_,
		_w7425_,
		_w7426_
	);
	LUT3 #(
		.INIT('h2a)
	) name4415 (
		\pci_target_unit_wishbone_master_read_bound_reg/NET0131 ,
		_w3057_,
		_w3050_,
		_w7427_
	);
	LUT4 #(
		.INIT('h1000)
	) name4416 (
		\pci_target_unit_wishbone_master_read_count_reg[0]/NET0131 ,
		\pci_target_unit_wishbone_master_read_count_reg[2]/NET0131 ,
		_w3057_,
		_w3050_,
		_w7428_
	);
	LUT3 #(
		.INIT('h54)
	) name4417 (
		_w3085_,
		_w7427_,
		_w7428_,
		_w7429_
	);
	LUT4 #(
		.INIT('h0010)
	) name4418 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg/NET0131 ,
		\pci_target_unit_wishbone_master_w_attempt_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\wishbone_slave_unit_del_sync_req_req_pending_reg/NET0131 ,
		_w7430_
	);
	LUT3 #(
		.INIT('h70)
	) name4419 (
		_w3163_,
		_w3164_,
		_w7430_,
		_w7431_
	);
	LUT4 #(
		.INIT('h0080)
	) name4420 (
		\configuration_wb_err_cs_bit0_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6833_,
		_w7432_
	);
	LUT3 #(
		.INIT('h40)
	) name4421 (
		_w3044_,
		_w3046_,
		_w7085_,
		_w7433_
	);
	LUT4 #(
		.INIT('hf2fa)
	) name4422 (
		\configuration_wb_err_cs_bit8_reg/NET0131 ,
		_w7171_,
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4423 (
		\configuration_status_bit15_11_reg[12]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7398_,
		_w7435_
	);
	LUT2 #(
		.INIT('he)
	) name4424 (
		\wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg/NET0131 ,
		_w7435_,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name4425 (
		\configuration_icr_bit2_0_reg[1]/NET0131 ,
		_w7432_,
		_w7437_
	);
	LUT4 #(
		.INIT('h4000)
	) name4426 (
		_w3044_,
		_w3046_,
		_w3956_,
		_w3958_,
		_w7438_
	);
	LUT3 #(
		.INIT('h2a)
	) name4427 (
		\configuration_isr_bit2_0_reg[1]/NET0131 ,
		_w7068_,
		_w7438_,
		_w7439_
	);
	LUT2 #(
		.INIT('he)
	) name4428 (
		_w7437_,
		_w7439_,
		_w7440_
	);
	LUT4 #(
		.INIT('hef00)
	) name4429 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_wr_to_fifo_reg/NET0131 ,
		_w7441_
	);
	LUT3 #(
		.INIT('hf8)
	) name4430 (
		_w3242_,
		_w6726_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h4)
	) name4431 (
		\pci_target_unit_del_sync_comp_rty_exp_clr_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131 ,
		_w7443_
	);
	LUT2 #(
		.INIT('h2)
	) name4432 (
		\pci_target_unit_del_sync_comp_req_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_comp_rty_exp_reg_reg/NET0131 ,
		_w7444_
	);
	LUT3 #(
		.INIT('hec)
	) name4433 (
		_w6986_,
		_w7443_,
		_w7444_,
		_w7445_
	);
	LUT4 #(
		.INIT('hef00)
	) name4434 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_rd_from_fifo_reg/NET0131 ,
		_w7446_
	);
	LUT2 #(
		.INIT('he)
	) name4435 (
		_w6670_,
		_w7446_,
		_w7447_
	);
	LUT4 #(
		.INIT('hef00)
	) name4436 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		_w7448_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4437 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[12]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[1]/NET0131 ,
		_w7449_
	);
	LUT2 #(
		.INIT('h9)
	) name4438 (
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[17]/NET0131 ,
		_w7450_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4439 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[27]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[2]/NET0131 ,
		_w7451_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4440 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[15]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[19]/NET0131 ,
		_w7452_
	);
	LUT4 #(
		.INIT('h8000)
	) name4441 (
		_w7451_,
		_w7452_,
		_w7449_,
		_w7450_,
		_w7453_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4442 (
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[7]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[9]/NET0131 ,
		_w7454_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4443 (
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[14]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[20]/NET0131 ,
		_w7455_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4444 (
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[13]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[31]/NET0131 ,
		_w7456_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4445 (
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[28]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[0]/NET0131 ,
		_w7457_
	);
	LUT4 #(
		.INIT('h8000)
	) name4446 (
		_w7456_,
		_w7457_,
		_w7454_,
		_w7455_,
		_w7458_
	);
	LUT2 #(
		.INIT('h6)
	) name4447 (
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[29]/NET0131 ,
		_w7459_
	);
	LUT2 #(
		.INIT('h6)
	) name4448 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[1]/NET0131 ,
		_w7460_
	);
	LUT3 #(
		.INIT('h02)
	) name4449 (
		_w3216_,
		_w7460_,
		_w7459_,
		_w7461_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4450 (
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[19]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[30]/NET0131 ,
		_w7462_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4451 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[11]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[16]/NET0131 ,
		_w7463_
	);
	LUT4 #(
		.INIT('hf531)
	) name4452 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[18]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[4]/NET0131 ,
		_w7464_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4453 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[3]/NET0131 ,
		_w7465_
	);
	LUT4 #(
		.INIT('h8000)
	) name4454 (
		_w7464_,
		_w7465_,
		_w7462_,
		_w7463_,
		_w7466_
	);
	LUT4 #(
		.INIT('h8000)
	) name4455 (
		_w7461_,
		_w7466_,
		_w7453_,
		_w7458_,
		_w7467_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4456 (
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[13]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[24]/NET0131 ,
		_w7468_
	);
	LUT4 #(
		.INIT('haf23)
	) name4457 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[11]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[2]/NET0131 ,
		_w7469_
	);
	LUT2 #(
		.INIT('h8)
	) name4458 (
		_w7468_,
		_w7469_,
		_w7470_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4459 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[10]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[22]/NET0131 ,
		_w7471_
	);
	LUT4 #(
		.INIT('hf531)
	) name4460 (
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[26]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[5]/NET0131 ,
		_w7472_
	);
	LUT4 #(
		.INIT('haf23)
	) name4461 (
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[21]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[25]/NET0131 ,
		_w7473_
	);
	LUT4 #(
		.INIT('haf23)
	) name4462 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[12]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[14]/NET0131 ,
		_w7474_
	);
	LUT4 #(
		.INIT('h8000)
	) name4463 (
		_w7473_,
		_w7474_,
		_w7471_,
		_w7472_,
		_w7475_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		_w7470_,
		_w7475_,
		_w7476_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4465 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[31]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[2]/NET0131 ,
		_w7477_
	);
	LUT4 #(
		.INIT('hf531)
	) name4466 (
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[20]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[3]/NET0131 ,
		_w7478_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4467 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[30]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[6]/NET0131 ,
		_w7479_
	);
	LUT4 #(
		.INIT('haf23)
	) name4468 (
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[8]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[9]/NET0131 ,
		_w7480_
	);
	LUT4 #(
		.INIT('h8000)
	) name4469 (
		_w7479_,
		_w7480_,
		_w7477_,
		_w7478_,
		_w7481_
	);
	LUT4 #(
		.INIT('hf531)
	) name4470 (
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[16]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[3]/NET0131 ,
		_w7482_
	);
	LUT4 #(
		.INIT('haf23)
	) name4471 (
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[25]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[2]/NET0131 ,
		_w7483_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4472 (
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[23]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[7]/NET0131 ,
		_w7484_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4473 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[10]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[23]/NET0131 ,
		_w7485_
	);
	LUT4 #(
		.INIT('h8000)
	) name4474 (
		_w7484_,
		_w7485_,
		_w7482_,
		_w7483_,
		_w7486_
	);
	LUT4 #(
		.INIT('hf531)
	) name4475 (
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[24]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[8]/NET0131 ,
		_w7487_
	);
	LUT4 #(
		.INIT('haf23)
	) name4476 (
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[4]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[6]/NET0131 ,
		_w7488_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4477 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[18]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[3]/NET0131 ,
		_w7489_
	);
	LUT4 #(
		.INIT('hf531)
	) name4478 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_bc_out_reg[0]/NET0131 ,
		_w7490_
	);
	LUT4 #(
		.INIT('h8000)
	) name4479 (
		_w7489_,
		_w7490_,
		_w7487_,
		_w7488_,
		_w7491_
	);
	LUT4 #(
		.INIT('haf23)
	) name4480 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[15]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[22]/NET0131 ,
		_w7492_
	);
	LUT4 #(
		.INIT('haf23)
	) name4481 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[28]/NET0131 ,
		_w7493_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4482 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[27]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[5]/NET0131 ,
		_w7494_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4483 (
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[21]/NET0131 ,
		\pci_target_unit_del_sync_addr_out_reg[26]/NET0131 ,
		_w7495_
	);
	LUT4 #(
		.INIT('h8000)
	) name4484 (
		_w7494_,
		_w7495_,
		_w7492_,
		_w7493_,
		_w7496_
	);
	LUT4 #(
		.INIT('h8000)
	) name4485 (
		_w7491_,
		_w7496_,
		_w7481_,
		_w7486_,
		_w7497_
	);
	LUT4 #(
		.INIT('heaaa)
	) name4486 (
		_w7448_,
		_w7476_,
		_w7467_,
		_w7497_,
		_w7498_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4487 (
		\configuration_status_bit15_11_reg[13]/NET0131 ,
		_w3043_,
		_w3047_,
		_w7197_,
		_w7499_
	);
	LUT2 #(
		.INIT('he)
	) name4488 (
		_w6832_,
		_w7499_,
		_w7500_
	);
	LUT4 #(
		.INIT('haf23)
	) name4489 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131 ,
		_w7501_
	);
	LUT2 #(
		.INIT('h9)
	) name4490 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]/NET0131 ,
		_w7502_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4491 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]/NET0131 ,
		_w7503_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4492 (
		\pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg/NET0131 ,
		_w7501_,
		_w7502_,
		_w7503_,
		_w7504_
	);
	LUT3 #(
		.INIT('h6c)
	) name4493 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w7504_,
		_w7505_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name4494 (
		_w3789_,
		_w3786_,
		_w6307_,
		_w6312_,
		_w7506_
	);
	LUT2 #(
		.INIT('hb)
	) name4495 (
		_w3022_,
		_w3793_,
		_w7507_
	);
	LUT4 #(
		.INIT('h0800)
	) name4496 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		pci_gnt_i_pad,
		\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 ,
		_w7508_
	);
	LUT3 #(
		.INIT('h40)
	) name4497 (
		_w3022_,
		_w3793_,
		_w7508_,
		_w7509_
	);
	LUT4 #(
		.INIT('hfefb)
	) name4498 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w7510_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4499 (
		_w3022_,
		_w3793_,
		_w7508_,
		_w7510_,
		_w7511_
	);
	LUT2 #(
		.INIT('hb)
	) name4500 (
		_w7506_,
		_w7511_,
		_w7512_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4501 (
		\configuration_interrupt_line_reg[3]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7513_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4502 (
		\configuration_interrupt_line_reg[4]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7514_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4503 (
		\configuration_interrupt_line_reg[5]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7515_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4504 (
		\configuration_interrupt_line_reg[7]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		_w3933_,
		_w7148_,
		_w7516_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4505 (
		\configuration_cache_line_size_reg_reg[3]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7517_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4506 (
		\configuration_cache_line_size_reg_reg[4]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7518_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4507 (
		\configuration_cache_line_size_reg_reg[5]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7519_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7520_
	);
	LUT2 #(
		.INIT('h6)
	) name4509 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7521_
	);
	LUT3 #(
		.INIT('he2)
	) name4510 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		_w7504_,
		_w7521_,
		_w7522_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name4511 (
		\configuration_cache_line_size_reg_reg[7]/NET0131 ,
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		_w3948_,
		_w7148_,
		_w7523_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4512 (
		\configuration_wb_err_cs_bit9_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6833_,
		_w7524_
	);
	LUT3 #(
		.INIT('h80)
	) name4513 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w3019_,
		_w6832_,
		_w7525_
	);
	LUT2 #(
		.INIT('he)
	) name4514 (
		_w7524_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h4)
	) name4515 (
		\configuration_sync_isr_2_delayed_bckp_bit_reg/NET0131 ,
		\configuration_sync_isr_2_sync_bckp_bit_reg/NET0131 ,
		_w7527_
	);
	LUT4 #(
		.INIT('h00ea)
	) name4516 (
		\configuration_sync_isr_2_del_bit_reg/NET0131 ,
		_w7073_,
		_w7438_,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h4)
	) name4517 (
		\configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg/NET0131 ,
		\configuration_sync_pci_err_cs_8_sync_bckp_bit_reg/NET0131 ,
		_w7529_
	);
	LUT4 #(
		.INIT('h00ea)
	) name4518 (
		\configuration_sync_pci_err_cs_8_del_bit_reg/NET0131 ,
		_w3841_,
		_w7433_,
		_w7529_,
		_w7530_
	);
	LUT3 #(
		.INIT('h80)
	) name4519 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w6612_,
		_w7504_,
		_w7531_
	);
	LUT2 #(
		.INIT('h2)
	) name4520 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w7532_
	);
	LUT3 #(
		.INIT('h80)
	) name4521 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7504_,
		_w7532_,
		_w7533_
	);
	LUT2 #(
		.INIT('h4)
	) name4522 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w7534_
	);
	LUT3 #(
		.INIT('h80)
	) name4523 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7504_,
		_w7534_,
		_w7535_
	);
	LUT3 #(
		.INIT('h80)
	) name4524 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w7504_,
		_w7520_,
		_w7536_
	);
	LUT3 #(
		.INIT('h0d)
	) name4525 (
		\output_backup_frame_out_reg/NET0131 ,
		_w3792_,
		_w6313_,
		_w7537_
	);
	LUT2 #(
		.INIT('h8)
	) name4526 (
		\output_backup_frame_out_reg/NET0131 ,
		_w3786_,
		_w7538_
	);
	LUT2 #(
		.INIT('h1)
	) name4527 (
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7539_
	);
	LUT3 #(
		.INIT('h10)
	) name4528 (
		_w3789_,
		_w6307_,
		_w7539_,
		_w7540_
	);
	LUT4 #(
		.INIT('h0111)
	) name4529 (
		_w7509_,
		_w7537_,
		_w7538_,
		_w7540_,
		_w7541_
	);
	LUT4 #(
		.INIT('hfeee)
	) name4530 (
		_w7509_,
		_w7537_,
		_w7538_,
		_w7540_,
		_w7542_
	);
	LUT2 #(
		.INIT('h6)
	) name4531 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w7504_,
		_w7543_
	);
	LUT3 #(
		.INIT('h40)
	) name4532 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7504_,
		_w7532_,
		_w7544_
	);
	LUT3 #(
		.INIT('h40)
	) name4533 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7504_,
		_w7534_,
		_w7545_
	);
	LUT3 #(
		.INIT('h40)
	) name4534 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w6608_,
		_w7504_,
		_w7546_
	);
	LUT3 #(
		.INIT('h40)
	) name4535 (
		\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w6612_,
		_w7504_,
		_w7547_
	);
	LUT3 #(
		.INIT('h60)
	) name4536 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[13]/NET0131 ,
		_w6513_,
		_w6518_,
		_w7548_
	);
	LUT3 #(
		.INIT('h60)
	) name4537 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[6]/NET0131 ,
		_w6508_,
		_w6518_,
		_w7549_
	);
	LUT2 #(
		.INIT('h8)
	) name4538 (
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7022_,
		_w7550_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name4539 (
		\pci_target_unit_fifos_inGreyCount_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7022_,
		_w7551_
	);
	LUT4 #(
		.INIT('h4000)
	) name4540 (
		\output_backup_frame_out_reg/NET0131 ,
		pci_gnt_i_pad,
		_w6740_,
		_w6743_,
		_w7552_
	);
	LUT3 #(
		.INIT('hc8)
	) name4541 (
		\wishbone_slave_unit_pci_initiator_sm_timeout_reg/NET0131 ,
		_w3019_,
		_w7552_,
		_w7553_
	);
	LUT4 #(
		.INIT('h80a0)
	) name4542 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w6833_,
		_w7554_
	);
	LUT3 #(
		.INIT('h6c)
	) name4543 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w7554_,
		_w7555_
	);
	LUT4 #(
		.INIT('h0222)
	) name4544 (
		_w6311_,
		_w7537_,
		_w7538_,
		_w7540_,
		_w7556_
	);
	LUT4 #(
		.INIT('hfddd)
	) name4545 (
		_w6311_,
		_w7537_,
		_w7538_,
		_w7540_,
		_w7557_
	);
	LUT4 #(
		.INIT('h0400)
	) name4546 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7558_
	);
	LUT2 #(
		.INIT('h8)
	) name4547 (
		_w7554_,
		_w7558_,
		_w7559_
	);
	LUT4 #(
		.INIT('h1000)
	) name4548 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7560_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		_w7554_,
		_w7560_,
		_w7561_
	);
	LUT4 #(
		.INIT('h0001)
	) name4550 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name4551 (
		_w7554_,
		_w7562_,
		_w7563_
	);
	LUT4 #(
		.INIT('h0002)
	) name4552 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7564_
	);
	LUT2 #(
		.INIT('h8)
	) name4553 (
		_w7554_,
		_w7564_,
		_w7565_
	);
	LUT4 #(
		.INIT('h0004)
	) name4554 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7566_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		_w7554_,
		_w7566_,
		_w7567_
	);
	LUT4 #(
		.INIT('h0008)
	) name4556 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7568_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		_w7554_,
		_w7568_,
		_w7569_
	);
	LUT4 #(
		.INIT('h0010)
	) name4558 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7570_
	);
	LUT2 #(
		.INIT('h8)
	) name4559 (
		_w7554_,
		_w7570_,
		_w7571_
	);
	LUT4 #(
		.INIT('h0020)
	) name4560 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name4561 (
		_w7554_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('h0040)
	) name4562 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7574_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		_w7554_,
		_w7574_,
		_w7575_
	);
	LUT4 #(
		.INIT('h0100)
	) name4564 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7576_
	);
	LUT2 #(
		.INIT('h8)
	) name4565 (
		_w7554_,
		_w7576_,
		_w7577_
	);
	LUT4 #(
		.INIT('h0200)
	) name4566 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7578_
	);
	LUT2 #(
		.INIT('h8)
	) name4567 (
		_w7554_,
		_w7578_,
		_w7579_
	);
	LUT3 #(
		.INIT('h02)
	) name4568 (
		\pci_target_unit_pci_target_if_target_rd_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg/NET0131 ,
		_w7580_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		_w6537_,
		_w7580_,
		_w7581_
	);
	LUT3 #(
		.INIT('hba)
	) name4570 (
		\pci_target_unit_del_sync_comp_flush_out_reg/NET0131 ,
		_w3255_,
		_w7581_,
		_w7582_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4571 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]/NET0131 ,
		_w7583_
	);
	LUT2 #(
		.INIT('h6)
	) name4572 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w7554_,
		_w7584_
	);
	LUT4 #(
		.INIT('h0800)
	) name4573 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7585_
	);
	LUT2 #(
		.INIT('h8)
	) name4574 (
		_w7554_,
		_w7585_,
		_w7586_
	);
	LUT4 #(
		.INIT('h4000)
	) name4575 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7587_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		_w7554_,
		_w7587_,
		_w7588_
	);
	LUT4 #(
		.INIT('h2000)
	) name4577 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7589_
	);
	LUT2 #(
		.INIT('h8)
	) name4578 (
		_w7554_,
		_w7589_,
		_w7590_
	);
	LUT4 #(
		.INIT('h8000)
	) name4579 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7591_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		_w7554_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('h8)
	) name4581 (
		_w6602_,
		_w7554_,
		_w7593_
	);
	LUT3 #(
		.INIT('h6a)
	) name4582 (
		\pci_target_unit_fifos_pciw_inTransactionCount_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7022_,
		_w7594_
	);
	LUT3 #(
		.INIT('h78)
	) name4583 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[2]/NET0131 ,
		_w7595_
	);
	LUT3 #(
		.INIT('h40)
	) name4584 (
		_w6516_,
		_w6517_,
		_w7595_,
		_w7596_
	);
	LUT3 #(
		.INIT('h60)
	) name4585 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[9]/NET0131 ,
		_w6510_,
		_w6518_,
		_w7597_
	);
	LUT4 #(
		.INIT('h3111)
	) name4586 (
		\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 ,
		_w3022_,
		_w3019_,
		_w3789_,
		_w7598_
	);
	LUT4 #(
		.INIT('ha222)
	) name4587 (
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_rdy_out_reg/NET0131 ,
		_w3018_,
		_w3019_,
		_w7599_
	);
	LUT4 #(
		.INIT('ha695)
	) name4588 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[1]/NET0131 ,
		\pci_cbe_i[1]_pad ,
		_w7600_
	);
	LUT4 #(
		.INIT('ha695)
	) name4589 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[0]/NET0131 ,
		\pci_cbe_i[0]_pad ,
		_w7601_
	);
	LUT4 #(
		.INIT('h596a)
	) name4590 (
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[2]/NET0131 ,
		\pci_cbe_i[2]_pad ,
		_w7602_
	);
	LUT4 #(
		.INIT('ha695)
	) name4591 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\output_backup_cbe_en_out_reg/NET0131 ,
		\output_backup_cbe_out_reg[3]/NET0131 ,
		\pci_cbe_i[3]_pad ,
		_w7603_
	);
	LUT4 #(
		.INIT('h4000)
	) name4592 (
		_w7602_,
		_w7603_,
		_w7600_,
		_w7601_,
		_w7604_
	);
	LUT2 #(
		.INIT('h1)
	) name4593 (
		\output_backup_trdy_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7605_
	);
	LUT2 #(
		.INIT('h4)
	) name4594 (
		_w7604_,
		_w7605_,
		_w7606_
	);
	LUT3 #(
		.INIT('h6c)
	) name4595 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 ,
		_w7022_,
		_w7607_
	);
	LUT3 #(
		.INIT('h6c)
	) name4596 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		_w7022_,
		_w7608_
	);
	LUT4 #(
		.INIT('he222)
	) name4597 (
		\pci_target_unit_pci_target_sm_cnf_progress_reg/NET0131 ,
		_w3216_,
		_w3698_,
		_w3748_,
		_w7609_
	);
	LUT2 #(
		.INIT('h9)
	) name4598 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7610_
	);
	LUT3 #(
		.INIT('h2e)
	) name4599 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]/NET0131 ,
		_w7022_,
		_w7610_,
		_w7611_
	);
	LUT2 #(
		.INIT('h6)
	) name4600 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131 ,
		_w7022_,
		_w7612_
	);
	LUT2 #(
		.INIT('h6)
	) name4601 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		_w7022_,
		_w7613_
	);
	LUT3 #(
		.INIT('h47)
	) name4602 (
		\output_backup_devsel_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		pci_devsel_i_pad,
		_w7614_
	);
	LUT3 #(
		.INIT('hb8)
	) name4603 (
		\output_backup_devsel_out_reg/NET0131 ,
		\output_backup_trdy_en_out_reg/NET0131 ,
		pci_devsel_i_pad,
		_w7615_
	);
	LUT4 #(
		.INIT('h0004)
	) name4604 (
		_w3789_,
		_w3786_,
		_w6307_,
		_w7614_,
		_w7616_
	);
	LUT3 #(
		.INIT('h1e)
	) name4605 (
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131 ,
		_w7617_
	);
	LUT2 #(
		.INIT('h7)
	) name4606 (
		_w7616_,
		_w7617_,
		_w7618_
	);
	LUT3 #(
		.INIT('h23)
	) name4607 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131 ,
		_w7619_
	);
	LUT3 #(
		.INIT('h45)
	) name4608 (
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131 ,
		\pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131 ,
		_w7620_
	);
	LUT2 #(
		.INIT('h4)
	) name4609 (
		_w7619_,
		_w7620_,
		_w7621_
	);
	LUT2 #(
		.INIT('h6)
	) name4610 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_comp_cycle_count_reg[1]/NET0131 ,
		_w7622_
	);
	LUT3 #(
		.INIT('h40)
	) name4611 (
		_w6516_,
		_w6517_,
		_w7622_,
		_w7623_
	);
	LUT3 #(
		.INIT('h60)
	) name4612 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[5]/NET0131 ,
		_w6507_,
		_w6518_,
		_w7624_
	);
	LUT3 #(
		.INIT('h78)
	) name4613 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7625_
	);
	LUT2 #(
		.INIT('h4)
	) name4614 (
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131 ,
		_w7616_,
		_w7626_
	);
	LUT2 #(
		.INIT('h6)
	) name4615 (
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131 ,
		_w7627_
	);
	LUT2 #(
		.INIT('h2)
	) name4616 (
		_w7616_,
		_w7627_,
		_w7628_
	);
	LUT3 #(
		.INIT('h10)
	) name4617 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[0]/NET0131 ,
		_w6516_,
		_w6517_,
		_w7629_
	);
	LUT4 #(
		.INIT('h0111)
	) name4618 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131 ,
		\pci_target_unit_del_sync_req_done_reg_reg/NET0131 ,
		_w6537_,
		_w7580_,
		_w7630_
	);
	LUT2 #(
		.INIT('h2)
	) name4619 (
		\pci_target_unit_del_sync_req_comp_pending_sample_reg/NET0131 ,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]/P0001 ,
		_w7558_,
		_w7632_
	);
	LUT3 #(
		.INIT('h20)
	) name4621 (
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]/NET0131 ,
		_w7633_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4622 (
		_w6831_,
		_w6832_,
		_w7558_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('he)
	) name4623 (
		_w7632_,
		_w7634_,
		_w7635_
	);
	LUT2 #(
		.INIT('h2)
	) name4624 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]/P0001 ,
		_w7560_,
		_w7636_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4625 (
		_w6831_,
		_w6832_,
		_w7560_,
		_w7633_,
		_w7637_
	);
	LUT2 #(
		.INIT('he)
	) name4626 (
		_w7636_,
		_w7637_,
		_w7638_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]/P0001 ,
		_w7587_,
		_w7639_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4628 (
		_w6831_,
		_w6832_,
		_w7587_,
		_w7633_,
		_w7640_
	);
	LUT2 #(
		.INIT('he)
	) name4629 (
		_w7639_,
		_w7640_,
		_w7641_
	);
	LUT2 #(
		.INIT('h2)
	) name4630 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]/P0001 ,
		_w7566_,
		_w7642_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4631 (
		_w6831_,
		_w6832_,
		_w7566_,
		_w7633_,
		_w7643_
	);
	LUT2 #(
		.INIT('he)
	) name4632 (
		_w7642_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h2)
	) name4633 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]/P0001 ,
		_w7570_,
		_w7645_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4634 (
		_w6831_,
		_w6832_,
		_w7570_,
		_w7633_,
		_w7646_
	);
	LUT2 #(
		.INIT('he)
	) name4635 (
		_w7645_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h2)
	) name4636 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]/P0001 ,
		_w7574_,
		_w7648_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4637 (
		_w6831_,
		_w6832_,
		_w7574_,
		_w7633_,
		_w7649_
	);
	LUT2 #(
		.INIT('he)
	) name4638 (
		_w7648_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]/P0001 ,
		_w7576_,
		_w7651_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4640 (
		_w6831_,
		_w6832_,
		_w7576_,
		_w7633_,
		_w7652_
	);
	LUT2 #(
		.INIT('he)
	) name4641 (
		_w7651_,
		_w7652_,
		_w7653_
	);
	LUT2 #(
		.INIT('h2)
	) name4642 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]/P0001 ,
		_w7585_,
		_w7654_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4643 (
		_w6831_,
		_w6832_,
		_w7585_,
		_w7633_,
		_w7655_
	);
	LUT2 #(
		.INIT('he)
	) name4644 (
		_w7654_,
		_w7655_,
		_w7656_
	);
	LUT2 #(
		.INIT('h2)
	) name4645 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]/P0001 ,
		_w7578_,
		_w7657_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4646 (
		_w6831_,
		_w6832_,
		_w7578_,
		_w7633_,
		_w7658_
	);
	LUT2 #(
		.INIT('he)
	) name4647 (
		_w7657_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h2)
	) name4648 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]/P0001 ,
		_w6602_,
		_w7660_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4649 (
		_w6602_,
		_w6831_,
		_w6832_,
		_w7633_,
		_w7661_
	);
	LUT2 #(
		.INIT('he)
	) name4650 (
		_w7660_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h2)
	) name4651 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]/P0001 ,
		_w7572_,
		_w7663_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4652 (
		_w6831_,
		_w6832_,
		_w7572_,
		_w7633_,
		_w7664_
	);
	LUT2 #(
		.INIT('he)
	) name4653 (
		_w7663_,
		_w7664_,
		_w7665_
	);
	LUT2 #(
		.INIT('h2)
	) name4654 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]/P0001 ,
		_w7568_,
		_w7666_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4655 (
		_w6831_,
		_w6832_,
		_w7568_,
		_w7633_,
		_w7667_
	);
	LUT2 #(
		.INIT('he)
	) name4656 (
		_w7666_,
		_w7667_,
		_w7668_
	);
	LUT2 #(
		.INIT('h2)
	) name4657 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]/P0001 ,
		_w7591_,
		_w7669_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4658 (
		_w6831_,
		_w6832_,
		_w7591_,
		_w7633_,
		_w7670_
	);
	LUT2 #(
		.INIT('he)
	) name4659 (
		_w7669_,
		_w7670_,
		_w7671_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]/P0001 ,
		_w7589_,
		_w7672_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4661 (
		_w6831_,
		_w6832_,
		_w7589_,
		_w7633_,
		_w7673_
	);
	LUT2 #(
		.INIT('he)
	) name4662 (
		_w7672_,
		_w7673_,
		_w7674_
	);
	LUT2 #(
		.INIT('h2)
	) name4663 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]/P0001 ,
		_w7564_,
		_w7675_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4664 (
		_w6831_,
		_w6832_,
		_w7564_,
		_w7633_,
		_w7676_
	);
	LUT2 #(
		.INIT('he)
	) name4665 (
		_w7675_,
		_w7676_,
		_w7677_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]/P0001 ,
		_w7562_,
		_w7678_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name4667 (
		_w6831_,
		_w6832_,
		_w7562_,
		_w7633_,
		_w7679_
	);
	LUT2 #(
		.INIT('he)
	) name4668 (
		_w7678_,
		_w7679_,
		_w7680_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4669 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001 ,
		_w7681_
	);
	LUT4 #(
		.INIT('h4000)
	) name4670 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7682_
	);
	LUT2 #(
		.INIT('he)
	) name4671 (
		_w7681_,
		_w7682_,
		_w7683_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4672 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001 ,
		_w7684_
	);
	LUT4 #(
		.INIT('h2000)
	) name4673 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7685_
	);
	LUT2 #(
		.INIT('he)
	) name4674 (
		_w7684_,
		_w7685_,
		_w7686_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4675 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001 ,
		_w7687_
	);
	LUT4 #(
		.INIT('h8000)
	) name4676 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7688_
	);
	LUT2 #(
		.INIT('he)
	) name4677 (
		_w7687_,
		_w7688_,
		_w7689_
	);
	LUT4 #(
		.INIT('hef00)
	) name4678 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001 ,
		_w7690_
	);
	LUT4 #(
		.INIT('h1000)
	) name4679 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7691_
	);
	LUT2 #(
		.INIT('he)
	) name4680 (
		_w7690_,
		_w7691_,
		_w7692_
	);
	LUT4 #(
		.INIT('hfb00)
	) name4681 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001 ,
		_w7693_
	);
	LUT4 #(
		.INIT('h0400)
	) name4682 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7694_
	);
	LUT2 #(
		.INIT('he)
	) name4683 (
		_w7693_,
		_w7694_,
		_w7695_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4684 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001 ,
		_w7696_
	);
	LUT4 #(
		.INIT('h0200)
	) name4685 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7697_
	);
	LUT2 #(
		.INIT('he)
	) name4686 (
		_w7696_,
		_w7697_,
		_w7698_
	);
	LUT4 #(
		.INIT('hf700)
	) name4687 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001 ,
		_w7699_
	);
	LUT4 #(
		.INIT('h0800)
	) name4688 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7700_
	);
	LUT2 #(
		.INIT('he)
	) name4689 (
		_w7699_,
		_w7700_,
		_w7701_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4690 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001 ,
		_w7702_
	);
	LUT4 #(
		.INIT('h0100)
	) name4691 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]/NET0131 ,
		_w7703_
	);
	LUT2 #(
		.INIT('he)
	) name4692 (
		_w7702_,
		_w7703_,
		_w7704_
	);
	LUT4 #(
		.INIT('he0a0)
	) name4693 (
		\wishbone_slave_unit_pci_initiator_sm_transfer_reg/NET0131 ,
		_w3789_,
		_w3786_,
		_w7614_,
		_w7705_
	);
	LUT3 #(
		.INIT('h78)
	) name4694 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7706_
	);
	LUT2 #(
		.INIT('h8)
	) name4695 (
		_w3019_,
		_w6831_,
		_w7707_
	);
	LUT3 #(
		.INIT('h82)
	) name4696 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]/NET0131 ,
		_w7708_
	);
	LUT4 #(
		.INIT('hff13)
	) name4697 (
		\wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		_w7011_,
		_w7708_,
		_w7709_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name4698 (
		\pci_target_unit_wishbone_master_first_wb_data_access_reg/NET0131 ,
		_w3052_,
		_w3068_,
		_w3050_,
		_w7710_
	);
	LUT3 #(
		.INIT('hca)
	) name4699 (
		\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]/NET0131 ,
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_done_reg_reg/NET0131 ,
		_w7711_
	);
	LUT4 #(
		.INIT('h1500)
	) name4700 (
		\pci_target_unit_del_sync_comp_cycle_count_reg[16]/NET0131 ,
		_w6537_,
		_w7580_,
		_w7711_,
		_w7712_
	);
	LUT3 #(
		.INIT('hd0)
	) name4701 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_if_target_rd_reg/NET0131 ,
		_w7713_
	);
	LUT3 #(
		.INIT('hd0)
	) name4702 (
		\output_backup_devsel_out_reg/NET0131 ,
		\output_backup_stop_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		_w7714_
	);
	LUT3 #(
		.INIT('h8a)
	) name4703 (
		\pci_target_unit_pci_target_if_same_read_reg_reg/NET0131 ,
		_w7713_,
		_w7714_,
		_w7715_
	);
	LUT3 #(
		.INIT('h80)
	) name4704 (
		\wishbone_slave_unit_pci_initiator_if_current_last_reg/NET0131 ,
		_w3019_,
		_w3789_,
		_w7716_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4705 (
		\output_backup_frame_out_reg/NET0131 ,
		_w3789_,
		_w6307_,
		_w6312_,
		_w7717_
	);
	LUT2 #(
		.INIT('h1)
	) name4706 (
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]/NET0131 ,
		_w7718_
	);
	LUT4 #(
		.INIT('h0100)
	) name4707 (
		_w3789_,
		_w6307_,
		_w7614_,
		_w7718_,
		_w7719_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name4708 (
		\wishbone_slave_unit_del_sync_bc_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]/NET0131 ,
		_w7011_,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		_w3216_,
		_w3739_,
		_w7721_
	);
	LUT3 #(
		.INIT('h78)
	) name4710 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w7722_
	);
	LUT3 #(
		.INIT('h78)
	) name4711 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]/NET0131 ,
		_w7723_
	);
	LUT3 #(
		.INIT('h8b)
	) name4712 (
		\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w6991_,
		_w7724_
	);
	LUT2 #(
		.INIT('h2)
	) name4713 (
		_w3050_,
		_w3075_,
		_w7725_
	);
	LUT3 #(
		.INIT('h78)
	) name4714 (
		\wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131 ,
		_w7726_
	);
	LUT3 #(
		.INIT('h78)
	) name4715 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131 ,
		_w7727_
	);
	LUT3 #(
		.INIT('hea)
	) name4716 (
		\wishbone_slave_unit_pci_initiator_if_del_read_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_if_write_req_int_reg/NET0131 ,
		_w7728_
	);
	LUT3 #(
		.INIT('h78)
	) name4717 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131 ,
		_w7729_
	);
	LUT4 #(
		.INIT('hef00)
	) name4718 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		_w7730_
	);
	LUT4 #(
		.INIT('h0200)
	) name4719 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7731_
	);
	LUT2 #(
		.INIT('he)
	) name4720 (
		_w7730_,
		_w7731_,
		_w7732_
	);
	LUT4 #(
		.INIT('h0200)
	) name4721 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7733_
	);
	LUT2 #(
		.INIT('he)
	) name4722 (
		_w3217_,
		_w7733_,
		_w7734_
	);
	LUT4 #(
		.INIT('hef00)
	) name4723 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		_w7735_
	);
	LUT4 #(
		.INIT('h0200)
	) name4724 (
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7736_
	);
	LUT2 #(
		.INIT('he)
	) name4725 (
		_w7735_,
		_w7736_,
		_w7737_
	);
	LUT4 #(
		.INIT('hef00)
	) name4726 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		_w7738_
	);
	LUT4 #(
		.INIT('h0200)
	) name4727 (
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7739_
	);
	LUT2 #(
		.INIT('he)
	) name4728 (
		_w7738_,
		_w7739_,
		_w7740_
	);
	LUT4 #(
		.INIT('hef00)
	) name4729 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		_w7741_
	);
	LUT4 #(
		.INIT('h0200)
	) name4730 (
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7742_
	);
	LUT2 #(
		.INIT('he)
	) name4731 (
		_w7741_,
		_w7742_,
		_w7743_
	);
	LUT4 #(
		.INIT('hef00)
	) name4732 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		_w7744_
	);
	LUT4 #(
		.INIT('h0200)
	) name4733 (
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7745_
	);
	LUT2 #(
		.INIT('he)
	) name4734 (
		_w7744_,
		_w7745_,
		_w7746_
	);
	LUT4 #(
		.INIT('hef00)
	) name4735 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		_w7747_
	);
	LUT4 #(
		.INIT('h0200)
	) name4736 (
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7748_
	);
	LUT2 #(
		.INIT('he)
	) name4737 (
		_w7747_,
		_w7748_,
		_w7749_
	);
	LUT4 #(
		.INIT('hef00)
	) name4738 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		_w7750_
	);
	LUT4 #(
		.INIT('h0200)
	) name4739 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7751_
	);
	LUT2 #(
		.INIT('he)
	) name4740 (
		_w7750_,
		_w7751_,
		_w7752_
	);
	LUT4 #(
		.INIT('hef00)
	) name4741 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		_w7753_
	);
	LUT4 #(
		.INIT('h0200)
	) name4742 (
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7754_
	);
	LUT2 #(
		.INIT('he)
	) name4743 (
		_w7753_,
		_w7754_,
		_w7755_
	);
	LUT4 #(
		.INIT('hef00)
	) name4744 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		_w7756_
	);
	LUT4 #(
		.INIT('h0200)
	) name4745 (
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7757_
	);
	LUT2 #(
		.INIT('he)
	) name4746 (
		_w7756_,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h8)
	) name4747 (
		\pci_target_unit_del_sync_req_rty_exp_clr_reg/NET0131 ,
		\pci_target_unit_del_sync_req_rty_exp_reg_reg/NET0131 ,
		_w7759_
	);
	LUT4 #(
		.INIT('hffe9)
	) name4748 (
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]/NET0131 ,
		_w7760_
	);
	LUT4 #(
		.INIT('hef00)
	) name4749 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		_w7761_
	);
	LUT4 #(
		.INIT('h0200)
	) name4750 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7762_
	);
	LUT2 #(
		.INIT('he)
	) name4751 (
		_w7761_,
		_w7762_,
		_w7763_
	);
	LUT4 #(
		.INIT('hef00)
	) name4752 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		_w7764_
	);
	LUT4 #(
		.INIT('h0200)
	) name4753 (
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_frame_en_out_reg/NET0131 ,
		\parity_checker_frame_dec2_reg/NET0131 ,
		_w7765_
	);
	LUT2 #(
		.INIT('he)
	) name4754 (
		_w7764_,
		_w7765_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		\configuration_cache_line_size_reg_reg[2]/NET0131 ,
		\configuration_cache_line_size_reg_reg[3]/NET0131 ,
		_w7767_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		\configuration_cache_line_size_reg_reg[0]/NET0131 ,
		\configuration_cache_line_size_reg_reg[1]/NET0131 ,
		_w7768_
	);
	LUT3 #(
		.INIT('h70)
	) name4757 (
		_w7011_,
		_w7767_,
		_w7768_,
		_w7769_
	);
	LUT2 #(
		.INIT('h2)
	) name4758 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7770_
	);
	LUT4 #(
		.INIT('h0200)
	) name4759 (
		\pci_target_unit_pci_target_if_norm_address_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7771_
	);
	LUT2 #(
		.INIT('he)
	) name4760 (
		_w7770_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h2)
	) name4761 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7773_
	);
	LUT4 #(
		.INIT('h0200)
	) name4762 (
		\pci_target_unit_pci_target_if_norm_address_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7774_
	);
	LUT2 #(
		.INIT('he)
	) name4763 (
		_w7773_,
		_w7774_,
		_w7775_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4764 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7776_
	);
	LUT3 #(
		.INIT('hae)
	) name4765 (
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7777_
	);
	LUT3 #(
		.INIT('hae)
	) name4766 (
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7778_
	);
	LUT3 #(
		.INIT('hae)
	) name4767 (
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7779_
	);
	LUT3 #(
		.INIT('hae)
	) name4768 (
		\input_register_pci_ad_reg_out_reg[0]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7780_
	);
	LUT3 #(
		.INIT('hae)
	) name4769 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7781_
	);
	LUT3 #(
		.INIT('hae)
	) name4770 (
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7782_
	);
	LUT3 #(
		.INIT('hae)
	) name4771 (
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7783_
	);
	LUT3 #(
		.INIT('hae)
	) name4772 (
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7784_
	);
	LUT3 #(
		.INIT('hae)
	) name4773 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7785_
	);
	LUT3 #(
		.INIT('hae)
	) name4774 (
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7786_
	);
	LUT3 #(
		.INIT('hae)
	) name4775 (
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7787_
	);
	LUT3 #(
		.INIT('hae)
	) name4776 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7788_
	);
	LUT3 #(
		.INIT('hae)
	) name4777 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7789_
	);
	LUT3 #(
		.INIT('hae)
	) name4778 (
		\input_register_pci_ad_reg_out_reg[1]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7790_
	);
	LUT3 #(
		.INIT('hae)
	) name4779 (
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7791_
	);
	LUT3 #(
		.INIT('hae)
	) name4780 (
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7792_
	);
	LUT3 #(
		.INIT('hae)
	) name4781 (
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7793_
	);
	LUT3 #(
		.INIT('hae)
	) name4782 (
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7794_
	);
	LUT3 #(
		.INIT('hae)
	) name4783 (
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7795_
	);
	LUT3 #(
		.INIT('hae)
	) name4784 (
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7796_
	);
	LUT3 #(
		.INIT('hae)
	) name4785 (
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7797_
	);
	LUT3 #(
		.INIT('hae)
	) name4786 (
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7798_
	);
	LUT3 #(
		.INIT('hae)
	) name4787 (
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7799_
	);
	LUT3 #(
		.INIT('hae)
	) name4788 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7800_
	);
	LUT3 #(
		.INIT('hae)
	) name4789 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7801_
	);
	LUT3 #(
		.INIT('hae)
	) name4790 (
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7802_
	);
	LUT3 #(
		.INIT('hae)
	) name4791 (
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7803_
	);
	LUT3 #(
		.INIT('hae)
	) name4792 (
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7804_
	);
	LUT3 #(
		.INIT('hae)
	) name4793 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7805_
	);
	LUT3 #(
		.INIT('hae)
	) name4794 (
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7806_
	);
	LUT3 #(
		.INIT('hae)
	) name4795 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7807_
	);
	LUT3 #(
		.INIT('hae)
	) name4796 (
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort1_reg/NET0131 ,
		\wishbone_slave_unit_pci_initiator_sm_mabort2_reg/NET0131 ,
		_w7808_
	);
	LUT4 #(
		.INIT('h0100)
	) name4797 (
		\input_register_pci_irdy_reg_out_reg/NET0131 ,
		\pci_target_unit_del_sync_req_comp_pending_reg/NET0131 ,
		\pci_target_unit_del_sync_req_req_pending_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_master_will_request_read_reg/NET0131 ,
		_w7809_
	);
	LUT2 #(
		.INIT('he)
	) name4798 (
		\configuration_init_complete_reg/NET0131 ,
		\configuration_rst_inactive_reg/NET0131 ,
		_w7810_
	);
	LUT2 #(
		.INIT('h2)
	) name4799 (
		\configuration_set_isr_bit2_reg/NET0131 ,
		\configuration_sync_isr_2_del_bit_reg/NET0131 ,
		_w7811_
	);
	LUT2 #(
		.INIT('h8)
	) name4800 (
		\configuration_icr_bit2_0_reg[0]/NET0131 ,
		wb_int_i_pad,
		_w7812_
	);
	LUT3 #(
		.INIT('h13)
	) name4801 (
		\configuration_icr_bit2_0_reg[0]/NET0131 ,
		\configuration_isr_bit2_0_reg[1]/NET0131 ,
		wb_int_i_pad,
		_w7813_
	);
	LUT2 #(
		.INIT('hb)
	) name4802 (
		_w7811_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		_w3060_,
		_w3050_,
		_w7815_
	);
	LUT4 #(
		.INIT('h00ba)
	) name4804 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\output_backup_stop_out_reg/NET0131 ,
		\output_backup_trdy_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7816_
	);
	LUT3 #(
		.INIT('hca)
	) name4805 (
		\input_register_pci_ad_reg_out_reg[12]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[12]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7817_
	);
	LUT3 #(
		.INIT('hca)
	) name4806 (
		\input_register_pci_ad_reg_out_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[5]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7818_
	);
	LUT3 #(
		.INIT('hca)
	) name4807 (
		\input_register_pci_ad_reg_out_reg[27]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[27]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7819_
	);
	LUT3 #(
		.INIT('hca)
	) name4808 (
		\input_register_pci_ad_reg_out_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[7]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7820_
	);
	LUT3 #(
		.INIT('hca)
	) name4809 (
		\input_register_pci_ad_reg_out_reg[20]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[20]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7821_
	);
	LUT3 #(
		.INIT('hca)
	) name4810 (
		\input_register_pci_ad_reg_out_reg[23]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[23]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7822_
	);
	LUT3 #(
		.INIT('hca)
	) name4811 (
		\input_register_pci_ad_reg_out_reg[16]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[16]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7823_
	);
	LUT3 #(
		.INIT('hca)
	) name4812 (
		\input_register_pci_ad_reg_out_reg[17]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[17]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7824_
	);
	LUT3 #(
		.INIT('hca)
	) name4813 (
		\input_register_pci_ad_reg_out_reg[13]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[13]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7825_
	);
	LUT3 #(
		.INIT('hca)
	) name4814 (
		\input_register_pci_ad_reg_out_reg[26]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[26]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7826_
	);
	LUT3 #(
		.INIT('hca)
	) name4815 (
		\input_register_pci_ad_reg_out_reg[21]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[21]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7827_
	);
	LUT3 #(
		.INIT('hca)
	) name4816 (
		\input_register_pci_ad_reg_out_reg[18]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[18]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7828_
	);
	LUT3 #(
		.INIT('hca)
	) name4817 (
		\input_register_pci_ad_reg_out_reg[19]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[19]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7829_
	);
	LUT3 #(
		.INIT('hca)
	) name4818 (
		\input_register_pci_ad_reg_out_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[4]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7830_
	);
	LUT3 #(
		.INIT('hca)
	) name4819 (
		\input_register_pci_cbe_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7831_
	);
	LUT3 #(
		.INIT('hca)
	) name4820 (
		\input_register_pci_ad_reg_out_reg[25]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[25]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7832_
	);
	LUT3 #(
		.INIT('hca)
	) name4821 (
		\input_register_pci_cbe_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7833_
	);
	LUT3 #(
		.INIT('hca)
	) name4822 (
		\input_register_pci_ad_reg_out_reg[10]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[10]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7834_
	);
	LUT3 #(
		.INIT('hca)
	) name4823 (
		\input_register_pci_ad_reg_out_reg[28]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[28]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7835_
	);
	LUT3 #(
		.INIT('hca)
	) name4824 (
		\input_register_pci_ad_reg_out_reg[11]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[11]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7836_
	);
	LUT3 #(
		.INIT('hca)
	) name4825 (
		\input_register_pci_ad_reg_out_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[2]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7837_
	);
	LUT3 #(
		.INIT('hca)
	) name4826 (
		\input_register_pci_ad_reg_out_reg[22]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[22]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7838_
	);
	LUT3 #(
		.INIT('hca)
	) name4827 (
		\input_register_pci_ad_reg_out_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[6]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7839_
	);
	LUT3 #(
		.INIT('hca)
	) name4828 (
		\input_register_pci_ad_reg_out_reg[30]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[30]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7840_
	);
	LUT3 #(
		.INIT('hca)
	) name4829 (
		\input_register_pci_ad_reg_out_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[8]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7841_
	);
	LUT3 #(
		.INIT('hca)
	) name4830 (
		\input_register_pci_ad_reg_out_reg[29]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[29]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7842_
	);
	LUT3 #(
		.INIT('hca)
	) name4831 (
		\input_register_pci_ad_reg_out_reg[9]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[9]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7843_
	);
	LUT3 #(
		.INIT('hca)
	) name4832 (
		\input_register_pci_ad_reg_out_reg[24]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[24]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7844_
	);
	LUT3 #(
		.INIT('hca)
	) name4833 (
		\input_register_pci_cbe_reg_out_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[1]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7845_
	);
	LUT3 #(
		.INIT('hca)
	) name4834 (
		\input_register_pci_ad_reg_out_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[3]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7846_
	);
	LUT3 #(
		.INIT('hca)
	) name4835 (
		\input_register_pci_cbe_reg_out_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_bc_reg[0]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7847_
	);
	LUT3 #(
		.INIT('hca)
	) name4836 (
		\input_register_pci_ad_reg_out_reg[15]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[15]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7848_
	);
	LUT3 #(
		.INIT('hca)
	) name4837 (
		\input_register_pci_ad_reg_out_reg[31]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[31]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7849_
	);
	LUT3 #(
		.INIT('hca)
	) name4838 (
		\input_register_pci_ad_reg_out_reg[14]/NET0131 ,
		\pci_target_unit_pci_target_if_norm_address_reg[14]/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7850_
	);
	LUT2 #(
		.INIT('h6)
	) name4839 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w7851_
	);
	LUT2 #(
		.INIT('h6)
	) name4840 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]/NET0131 ,
		_w7852_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		\input_register_pci_frame_reg_out_reg/NET0131 ,
		\pci_target_unit_pci_target_sm_bckp_trdy_reg_reg/NET0131 ,
		_w7853_
	);
	LUT2 #(
		.INIT('h6)
	) name4842 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7854_
	);
	LUT2 #(
		.INIT('h6)
	) name4843 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		_w7855_
	);
	LUT2 #(
		.INIT('h8)
	) name4844 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]/P0001 ,
		\wishbone_slave_unit_pci_initiator_if_posted_write_req_reg/NET0131 ,
		_w7856_
	);
	LUT2 #(
		.INIT('h6)
	) name4845 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]/NET0131 ,
		_w7857_
	);
	LUT2 #(
		.INIT('h6)
	) name4846 (
		\wishbone_slave_unit_fifos_outGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]/NET0131 ,
		_w7858_
	);
	LUT2 #(
		.INIT('h6)
	) name4847 (
		\wishbone_slave_unit_fifos_inGreyCount_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]/NET0131 ,
		_w7859_
	);
	LUT4 #(
		.INIT('hdfff)
	) name4848 (
		\i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_map_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_mrl_en_reg/NET0131 ,
		\wishbone_slave_unit_wishbone_slave_pref_en_reg/NET0131 ,
		_w7860_
	);
	LUT2 #(
		.INIT('h6)
	) name4849 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w7861_
	);
	LUT2 #(
		.INIT('h6)
	) name4850 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]/NET0131 ,
		_w7862_
	);
	LUT2 #(
		.INIT('h6)
	) name4851 (
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7863_
	);
	LUT2 #(
		.INIT('h6)
	) name4852 (
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]/NET0131 ,
		\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w7864_
	);
	LUT2 #(
		.INIT('h6)
	) name4853 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]/NET0131 ,
		_w7865_
	);
	LUT2 #(
		.INIT('h6)
	) name4854 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]/NET0131 ,
		_w7866_
	);
	LUT2 #(
		.INIT('h6)
	) name4855 (
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]/NET0131 ,
		\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]/NET0131 ,
		_w7867_
	);
	LUT2 #(
		.INIT('h2)
	) name4856 (
		\configuration_set_pci_err_cs_bit8_reg/NET0131 ,
		\configuration_sync_pci_err_cs_8_del_bit_reg/NET0131 ,
		_w7868_
	);
	LUT2 #(
		.INIT('h8)
	) name4857 (
		\output_backup_frame_en_out_reg/NET0131 ,
		\output_backup_irdy_en_out_reg/NET0131 ,
		_w7869_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4858 (
		\wbm_dat_o[10]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w7870_
	);
	LUT4 #(
		.INIT('h0080)
	) name4859 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w7871_
	);
	LUT2 #(
		.INIT('he)
	) name4860 (
		_w7870_,
		_w7871_,
		_w7872_
	);
	LUT3 #(
		.INIT('h80)
	) name4861 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]/P0001 ,
		_w5559_,
		_w5564_,
		_w7873_
	);
	LUT3 #(
		.INIT('h80)
	) name4862 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]/P0001 ,
		_w5566_,
		_w5567_,
		_w7874_
	);
	LUT3 #(
		.INIT('h80)
	) name4863 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]/P0001 ,
		_w5566_,
		_w5576_,
		_w7875_
	);
	LUT3 #(
		.INIT('h80)
	) name4864 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]/P0001 ,
		_w5569_,
		_w5559_,
		_w7876_
	);
	LUT4 #(
		.INIT('h0001)
	) name4865 (
		_w7873_,
		_w7874_,
		_w7875_,
		_w7876_,
		_w7877_
	);
	LUT3 #(
		.INIT('h80)
	) name4866 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]/P0001 ,
		_w5576_,
		_w5570_,
		_w7878_
	);
	LUT3 #(
		.INIT('h80)
	) name4867 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]/P0001 ,
		_w5570_,
		_w5567_,
		_w7879_
	);
	LUT3 #(
		.INIT('h80)
	) name4868 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]/P0001 ,
		_w5570_,
		_w5564_,
		_w7880_
	);
	LUT3 #(
		.INIT('h80)
	) name4869 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]/P0001 ,
		_w5576_,
		_w5559_,
		_w7881_
	);
	LUT4 #(
		.INIT('h0001)
	) name4870 (
		_w7878_,
		_w7879_,
		_w7880_,
		_w7881_,
		_w7882_
	);
	LUT3 #(
		.INIT('h80)
	) name4871 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]/P0001 ,
		_w5566_,
		_w5564_,
		_w7883_
	);
	LUT3 #(
		.INIT('h80)
	) name4872 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]/P0001 ,
		_w5569_,
		_w5570_,
		_w7884_
	);
	LUT3 #(
		.INIT('h80)
	) name4873 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]/P0001 ,
		_w5569_,
		_w5566_,
		_w7885_
	);
	LUT3 #(
		.INIT('h80)
	) name4874 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]/P0001 ,
		_w5569_,
		_w5572_,
		_w7886_
	);
	LUT4 #(
		.INIT('h0001)
	) name4875 (
		_w7883_,
		_w7884_,
		_w7885_,
		_w7886_,
		_w7887_
	);
	LUT3 #(
		.INIT('h80)
	) name4876 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]/P0001 ,
		_w5567_,
		_w5572_,
		_w7888_
	);
	LUT3 #(
		.INIT('h80)
	) name4877 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]/P0001 ,
		_w5576_,
		_w5572_,
		_w7889_
	);
	LUT3 #(
		.INIT('h80)
	) name4878 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]/P0001 ,
		_w5564_,
		_w5572_,
		_w7890_
	);
	LUT3 #(
		.INIT('h80)
	) name4879 (
		\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]/P0001 ,
		_w5559_,
		_w5567_,
		_w7891_
	);
	LUT4 #(
		.INIT('h0001)
	) name4880 (
		_w7888_,
		_w7889_,
		_w7890_,
		_w7891_,
		_w7892_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4881 (
		_w7887_,
		_w7892_,
		_w7877_,
		_w7882_,
		_w7893_
	);
	LUT4 #(
		.INIT('h2223)
	) name4882 (
		_w6309_,
		_w6316_,
		_w6318_,
		_w6319_,
		_w7894_
	);
	LUT4 #(
		.INIT('h153f)
	) name4883 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]/P0001 ,
		_w5184_,
		_w5185_,
		_w7895_
	);
	LUT4 #(
		.INIT('h135f)
	) name4884 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]/P0001 ,
		_w5172_,
		_w5188_,
		_w7896_
	);
	LUT4 #(
		.INIT('h153f)
	) name4885 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]/P0001 ,
		_w5177_,
		_w5178_,
		_w7897_
	);
	LUT4 #(
		.INIT('h153f)
	) name4886 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]/P0001 ,
		_w5174_,
		_w5190_,
		_w7898_
	);
	LUT4 #(
		.INIT('h8000)
	) name4887 (
		_w7897_,
		_w7898_,
		_w7895_,
		_w7896_,
		_w7899_
	);
	LUT4 #(
		.INIT('h135f)
	) name4888 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]/P0001 ,
		_w5181_,
		_w5193_,
		_w7900_
	);
	LUT4 #(
		.INIT('h153f)
	) name4889 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]/P0001 ,
		_w5191_,
		_w5187_,
		_w7901_
	);
	LUT4 #(
		.INIT('h135f)
	) name4890 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]/P0001 ,
		_w5180_,
		_w5194_,
		_w7902_
	);
	LUT4 #(
		.INIT('h135f)
	) name4891 (
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]/P0001 ,
		\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]/P0001 ,
		_w5171_,
		_w5175_,
		_w7903_
	);
	LUT4 #(
		.INIT('h8000)
	) name4892 (
		_w7902_,
		_w7903_,
		_w7900_,
		_w7901_,
		_w7904_
	);
	LUT2 #(
		.INIT('h7)
	) name4893 (
		_w7899_,
		_w7904_,
		_w7905_
	);
	LUT4 #(
		.INIT('h2000)
	) name4894 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7906_
	);
	LUT4 #(
		.INIT('h8000)
	) name4895 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7907_
	);
	LUT4 #(
		.INIT('h0200)
	) name4896 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7908_
	);
	LUT4 #(
		.INIT('h0800)
	) name4897 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7909_
	);
	LUT4 #(
		.INIT('h0001)
	) name4898 (
		_w7906_,
		_w7907_,
		_w7908_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('h0080)
	) name4899 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7911_
	);
	LUT4 #(
		.INIT('h0020)
	) name4900 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7912_
	);
	LUT4 #(
		.INIT('h0002)
	) name4901 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7913_
	);
	LUT4 #(
		.INIT('h0008)
	) name4902 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7914_
	);
	LUT4 #(
		.INIT('h0001)
	) name4903 (
		_w7911_,
		_w7912_,
		_w7913_,
		_w7914_,
		_w7915_
	);
	LUT2 #(
		.INIT('h7)
	) name4904 (
		_w7910_,
		_w7915_,
		_w7916_
	);
	LUT4 #(
		.INIT('h8000)
	) name4905 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7917_
	);
	LUT4 #(
		.INIT('h2000)
	) name4906 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7918_
	);
	LUT4 #(
		.INIT('h0002)
	) name4907 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7919_
	);
	LUT4 #(
		.INIT('h0008)
	) name4908 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7920_
	);
	LUT4 #(
		.INIT('h0001)
	) name4909 (
		_w7917_,
		_w7918_,
		_w7919_,
		_w7920_,
		_w7921_
	);
	LUT4 #(
		.INIT('h0020)
	) name4910 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7922_
	);
	LUT4 #(
		.INIT('h0080)
	) name4911 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7923_
	);
	LUT4 #(
		.INIT('h0200)
	) name4912 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7924_
	);
	LUT4 #(
		.INIT('h0800)
	) name4913 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7925_
	);
	LUT4 #(
		.INIT('h0001)
	) name4914 (
		_w7922_,
		_w7923_,
		_w7924_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h7)
	) name4915 (
		_w7921_,
		_w7926_,
		_w7927_
	);
	LUT4 #(
		.INIT('h2000)
	) name4916 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7928_
	);
	LUT4 #(
		.INIT('h0002)
	) name4917 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7929_
	);
	LUT4 #(
		.INIT('h0008)
	) name4918 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7930_
	);
	LUT4 #(
		.INIT('h8000)
	) name4919 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7931_
	);
	LUT4 #(
		.INIT('h0001)
	) name4920 (
		_w7928_,
		_w7929_,
		_w7930_,
		_w7931_,
		_w7932_
	);
	LUT4 #(
		.INIT('h0020)
	) name4921 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7933_
	);
	LUT4 #(
		.INIT('h0080)
	) name4922 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7934_
	);
	LUT4 #(
		.INIT('h0200)
	) name4923 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7935_
	);
	LUT4 #(
		.INIT('h0800)
	) name4924 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7936_
	);
	LUT4 #(
		.INIT('h0001)
	) name4925 (
		_w7933_,
		_w7934_,
		_w7935_,
		_w7936_,
		_w7937_
	);
	LUT2 #(
		.INIT('h7)
	) name4926 (
		_w7932_,
		_w7937_,
		_w7938_
	);
	LUT4 #(
		.INIT('h0020)
	) name4927 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7939_
	);
	LUT4 #(
		.INIT('h0080)
	) name4928 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7940_
	);
	LUT4 #(
		.INIT('h0002)
	) name4929 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7941_
	);
	LUT4 #(
		.INIT('h0008)
	) name4930 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7942_
	);
	LUT4 #(
		.INIT('h0001)
	) name4931 (
		_w7939_,
		_w7940_,
		_w7941_,
		_w7942_,
		_w7943_
	);
	LUT4 #(
		.INIT('h0200)
	) name4932 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7944_
	);
	LUT4 #(
		.INIT('h0800)
	) name4933 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7945_
	);
	LUT4 #(
		.INIT('h2000)
	) name4934 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7946_
	);
	LUT4 #(
		.INIT('h8000)
	) name4935 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7947_
	);
	LUT4 #(
		.INIT('h0001)
	) name4936 (
		_w7944_,
		_w7945_,
		_w7946_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('h7)
	) name4937 (
		_w7943_,
		_w7948_,
		_w7949_
	);
	LUT4 #(
		.INIT('h0020)
	) name4938 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7950_
	);
	LUT4 #(
		.INIT('h0080)
	) name4939 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7951_
	);
	LUT4 #(
		.INIT('h0002)
	) name4940 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7952_
	);
	LUT4 #(
		.INIT('h0008)
	) name4941 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7953_
	);
	LUT4 #(
		.INIT('h0001)
	) name4942 (
		_w7950_,
		_w7951_,
		_w7952_,
		_w7953_,
		_w7954_
	);
	LUT4 #(
		.INIT('h0200)
	) name4943 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7955_
	);
	LUT4 #(
		.INIT('h0800)
	) name4944 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7956_
	);
	LUT4 #(
		.INIT('h2000)
	) name4945 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7957_
	);
	LUT4 #(
		.INIT('h8000)
	) name4946 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7958_
	);
	LUT4 #(
		.INIT('h0001)
	) name4947 (
		_w7955_,
		_w7956_,
		_w7957_,
		_w7958_,
		_w7959_
	);
	LUT2 #(
		.INIT('h7)
	) name4948 (
		_w7954_,
		_w7959_,
		_w7960_
	);
	LUT4 #(
		.INIT('h0008)
	) name4949 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7961_
	);
	LUT4 #(
		.INIT('h0002)
	) name4950 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7962_
	);
	LUT4 #(
		.INIT('h0080)
	) name4951 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7963_
	);
	LUT4 #(
		.INIT('h0020)
	) name4952 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7964_
	);
	LUT4 #(
		.INIT('h0001)
	) name4953 (
		_w7961_,
		_w7962_,
		_w7963_,
		_w7964_,
		_w7965_
	);
	LUT4 #(
		.INIT('h0800)
	) name4954 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7966_
	);
	LUT4 #(
		.INIT('h0200)
	) name4955 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7967_
	);
	LUT4 #(
		.INIT('h2000)
	) name4956 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7968_
	);
	LUT4 #(
		.INIT('h8000)
	) name4957 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7969_
	);
	LUT4 #(
		.INIT('h0001)
	) name4958 (
		_w7966_,
		_w7967_,
		_w7968_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h7)
	) name4959 (
		_w7965_,
		_w7970_,
		_w7971_
	);
	LUT4 #(
		.INIT('h0008)
	) name4960 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7972_
	);
	LUT4 #(
		.INIT('h0002)
	) name4961 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7973_
	);
	LUT4 #(
		.INIT('h0080)
	) name4962 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7974_
	);
	LUT4 #(
		.INIT('h0020)
	) name4963 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7975_
	);
	LUT4 #(
		.INIT('h0001)
	) name4964 (
		_w7972_,
		_w7973_,
		_w7974_,
		_w7975_,
		_w7976_
	);
	LUT4 #(
		.INIT('h0800)
	) name4965 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7977_
	);
	LUT4 #(
		.INIT('h0200)
	) name4966 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7978_
	);
	LUT4 #(
		.INIT('h2000)
	) name4967 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7979_
	);
	LUT4 #(
		.INIT('h8000)
	) name4968 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7980_
	);
	LUT4 #(
		.INIT('h0001)
	) name4969 (
		_w7977_,
		_w7978_,
		_w7979_,
		_w7980_,
		_w7981_
	);
	LUT2 #(
		.INIT('h7)
	) name4970 (
		_w7976_,
		_w7981_,
		_w7982_
	);
	LUT4 #(
		.INIT('h0008)
	) name4971 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7983_
	);
	LUT4 #(
		.INIT('h0002)
	) name4972 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7984_
	);
	LUT4 #(
		.INIT('h0080)
	) name4973 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7985_
	);
	LUT4 #(
		.INIT('h0020)
	) name4974 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7986_
	);
	LUT4 #(
		.INIT('h0001)
	) name4975 (
		_w7983_,
		_w7984_,
		_w7985_,
		_w7986_,
		_w7987_
	);
	LUT4 #(
		.INIT('h0800)
	) name4976 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7988_
	);
	LUT4 #(
		.INIT('h0200)
	) name4977 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7989_
	);
	LUT4 #(
		.INIT('h2000)
	) name4978 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7990_
	);
	LUT4 #(
		.INIT('h8000)
	) name4979 (
		\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]/P0001 ,
		_w4480_,
		_w4479_,
		_w4481_,
		_w7991_
	);
	LUT4 #(
		.INIT('h0001)
	) name4980 (
		_w7988_,
		_w7989_,
		_w7990_,
		_w7991_,
		_w7992_
	);
	LUT2 #(
		.INIT('h7)
	) name4981 (
		_w7987_,
		_w7992_,
		_w7993_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4982 (
		\wbm_dat_o[22]_pad ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w7994_
	);
	LUT4 #(
		.INIT('h0080)
	) name4983 (
		\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]/P0001 ,
		_w3097_,
		_w3104_,
		_w3183_,
		_w7995_
	);
	LUT2 #(
		.INIT('he)
	) name4984 (
		_w7994_,
		_w7995_,
		_w7996_
	);
	LUT4 #(
		.INIT('haa08)
	) name4985 (
		_w3135_,
		_w3147_,
		_w3150_,
		_w3160_,
		_w7997_
	);
	LUT2 #(
		.INIT('hb)
	) name4986 (
		\configuration_icr_bit31_reg/NET0131 ,
		pci_rst_i_pad,
		_w7998_
	);
	assign \configuration_init_complete_reg/P0001  = _w20_ ;
	assign \configuration_interrupt_out_reg/P0001  = _w30_ ;
	assign \g21/_0_  = _w3034_ ;
	assign \g52241/_0_  = _w3049_ ;
	assign \g52244/_0_  = _w3129_ ;
	assign \g52348/_0_  = _w3181_ ;
	assign \g52349/_0_  = _w3188_ ;
	assign \g52350/_0_  = _w3193_ ;
	assign \g52351/_0_  = _w3198_ ;
	assign \g52352/_0_  = _w3203_ ;
	assign \g52390/_0_  = _w3274_ ;
	assign \g52391/_0_  = _w3275_ ;
	assign \g52393/_3_  = _w3287_ ;
	assign \g52394/_3_  = _w3293_ ;
	assign \g52395/_3_  = _w3298_ ;
	assign \g52396/_3_  = _w3301_ ;
	assign \g52397/_3_  = _w3308_ ;
	assign \g52398/_3_  = _w3313_ ;
	assign \g52399/_3_  = _w3317_ ;
	assign \g52400/_3_  = _w3323_ ;
	assign \g52401/_3_  = _w3327_ ;
	assign \g52402/_3_  = _w3331_ ;
	assign \g52403/_3_  = _w3337_ ;
	assign \g52404/_3_  = _w3340_ ;
	assign \g52405/_3_  = _w3344_ ;
	assign \g52406/_0_  = _w3347_ ;
	assign \g52408/_0_  = _w3350_ ;
	assign \g52409/_0_  = _w3353_ ;
	assign \g52410/_0_  = _w3356_ ;
	assign \g52411/_0_  = _w3359_ ;
	assign \g52412/_0_  = _w3362_ ;
	assign \g52413/_0_  = _w3365_ ;
	assign \g52414/_0_  = _w3368_ ;
	assign \g52415/_0_  = _w3371_ ;
	assign \g52416/_0_  = _w3374_ ;
	assign \g52417/_0_  = _w3377_ ;
	assign \g52418/_0_  = _w3380_ ;
	assign \g52419/_0_  = _w3383_ ;
	assign \g52421/_0_  = _w3386_ ;
	assign \g52422/_0_  = _w3389_ ;
	assign \g52423/_0_  = _w3392_ ;
	assign \g52424/_0_  = _w3395_ ;
	assign \g52425/_0_  = _w3398_ ;
	assign \g52426/_0_  = _w3401_ ;
	assign \g52427/_0_  = _w3404_ ;
	assign \g52428/_0_  = _w3407_ ;
	assign \g52429/_0_  = _w3410_ ;
	assign \g52430/_0_  = _w3413_ ;
	assign \g52431/_0_  = _w3416_ ;
	assign \g52432/_0_  = _w3419_ ;
	assign \g52433/_0_  = _w3422_ ;
	assign \g52434/_0_  = _w3425_ ;
	assign \g52435/_0_  = _w3428_ ;
	assign \g52436/_0_  = _w3431_ ;
	assign \g52437/_0_  = _w3434_ ;
	assign \g52439/_3_  = _w3438_ ;
	assign \g52440/_3_  = _w3443_ ;
	assign \g52441/_3_  = _w3447_ ;
	assign \g52442/_3_  = _w3450_ ;
	assign \g52443/_3_  = _w3454_ ;
	assign \g52444/_3_  = _w3457_ ;
	assign \g52445/_3_  = _w3461_ ;
	assign \g52446/_3_  = _w3464_ ;
	assign \g52447/_3_  = _w3468_ ;
	assign \g52448/_3_  = _w3472_ ;
	assign \g52449/_3_  = _w3474_ ;
	assign \g52450/_3_  = _w3478_ ;
	assign \g52451/_3_  = _w3483_ ;
	assign \g52452/_3_  = _w3487_ ;
	assign \g52453/_3_  = _w3490_ ;
	assign \g52454/_3_  = _w3494_ ;
	assign \g52455/_3_  = _w3499_ ;
	assign \g52456/_3_  = _w3507_ ;
	assign \g52457/_3_  = _w3513_ ;
	assign \g52458/_3_  = _w3515_ ;
	assign \g52459/_3_  = _w3521_ ;
	assign \g52460/_3_  = _w3525_ ;
	assign \g52461/_3_  = _w3528_ ;
	assign \g52462/_3_  = _w3530_ ;
	assign \g52463/_3_  = _w3535_ ;
	assign \g52464/_3_  = _w3536_ ;
	assign \g52465/_3_  = _w3540_ ;
	assign \g52466/_3_  = _w3543_ ;
	assign \g52467/_3_  = _w3547_ ;
	assign \g52468/_3_  = _w3551_ ;
	assign \g52469/_3_  = _w3556_ ;
	assign \g52470/_3_  = _w3563_ ;
	assign \g52471/_3_  = _w3567_ ;
	assign \g52472/_3_  = _w3571_ ;
	assign \g52473/_3_  = _w3577_ ;
	assign \g52474/_3_  = _w3581_ ;
	assign \g52475/_3_  = _w3585_ ;
	assign \g52476/_3_  = _w3591_ ;
	assign \g52477/_3_  = _w3597_ ;
	assign \g52478/_3_  = _w3601_ ;
	assign \g52479/_3_  = _w3602_ ;
	assign \g52480/_3_  = _w3606_ ;
	assign \g52481/_3_  = _w3607_ ;
	assign \g52482/_3_  = _w3610_ ;
	assign \g52483/_3_  = _w3614_ ;
	assign \g52484/_3_  = _w3615_ ;
	assign \g52485/_3_  = _w3616_ ;
	assign \g52499/_0_  = _w3621_ ;
	assign \g52500/_0_  = _w3627_ ;
	assign \g52501/_0_  = _w3631_ ;
	assign \g52547/_0_  = _w3634_ ;
	assign \g52550/_0_  = _w3641_ ;
	assign \g52553/_0_  = _w3655_ ;
	assign \g52675/_0__syn_2  = _w3656_ ;
	assign \g52714/_0_  = _w3658_ ;
	assign \g52715/_0_  = _w3660_ ;
	assign \g52716/_0_  = _w3667_ ;
	assign \g52717/_0_  = _w3670_ ;
	assign \g52718/_0_  = _w3675_ ;
	assign \g52720/_0_  = _w3676_ ;
	assign \g52865/_0_  = _w3752_ ;
	assign \g52867/_0_  = _w3780_ ;
	assign \g52867/_1_  = _w3781_ ;
	assign \g52868/_0_  = _w3785_ ;
	assign \g52871/_2_  = _w3855_ ;
	assign \g52897/_0_  = _w3880_ ;
	assign \g52898/_0_  = _w3902_ ;
	assign \g52899/_0_  = _w3924_ ;
	assign \g52900/_0_  = _w3945_ ;
	assign \g52901/_0_  = _w3980_ ;
	assign \g52902/_0_  = _w4002_ ;
	assign \g52903/_0_  = _w4022_ ;
	assign \g52904/_0_  = _w4042_ ;
	assign \g52905/_0_  = _w4062_ ;
	assign \g52906/_0_  = _w4085_ ;
	assign \g52907/_0_  = _w4110_ ;
	assign \g52908/_0_  = _w4135_ ;
	assign \g52909/_0_  = _w4161_ ;
	assign \g52910/_0_  = _w4189_ ;
	assign \g52911/_0_  = _w4212_ ;
	assign \g52912/_0_  = _w4229_ ;
	assign \g52913/_0_  = _w4248_ ;
	assign \g52914/_0_  = _w4265_ ;
	assign \g52915/_0_  = _w4283_ ;
	assign \g52916/_0_  = _w4302_ ;
	assign \g52917/_0_  = _w4327_ ;
	assign \g52918/_0_  = _w4349_ ;
	assign \g52920/_0_  = _w4370_ ;
	assign \g52921/_0_  = _w4390_ ;
	assign \g52922/_0_  = _w4414_ ;
	assign \g52923/_0_  = _w4434_ ;
	assign \g52924/_0_  = _w4454_ ;
	assign \g52925/_0_  = _w4474_ ;
	assign \g52948/_0_  = _w4477_ ;
	assign \g52958/_0_  = _w4492_ ;
	assign \g52959/_0_  = _w4503_ ;
	assign \g52960/_0_  = _w4514_ ;
	assign \g52961/_0_  = _w4525_ ;
	assign \g52962/_0_  = _w4536_ ;
	assign \g52963/_0_  = _w4547_ ;
	assign \g52965/_0_  = _w4558_ ;
	assign \g52966/_0_  = _w4569_ ;
	assign \g52969/_0_  = _w4580_ ;
	assign \g52970/_0_  = _w4591_ ;
	assign \g52971/_0_  = _w4602_ ;
	assign \g52972/_0_  = _w4613_ ;
	assign \g52973/_0_  = _w4624_ ;
	assign \g52975/_0_  = _w4635_ ;
	assign \g52976/_0_  = _w4646_ ;
	assign \g52977/_0_  = _w4657_ ;
	assign \g52978/_0_  = _w4668_ ;
	assign \g52979/_0_  = _w4679_ ;
	assign \g52980/_0_  = _w4690_ ;
	assign \g52981/_0_  = _w4701_ ;
	assign \g52982/_0_  = _w4712_ ;
	assign \g52983/_0_  = _w4723_ ;
	assign \g52984/_0_  = _w4734_ ;
	assign \g52985/_0_  = _w4745_ ;
	assign \g52986/_0_  = _w4756_ ;
	assign \g52988/_0_  = _w4767_ ;
	assign \g52990/_0_  = _w4778_ ;
	assign \g52991/_0_  = _w4789_ ;
	assign \g52993/_0_  = _w4800_ ;
	assign \g52994/_0_  = _w4811_ ;
	assign \g52996/_0_  = _w4822_ ;
	assign \g52997/_0_  = _w4833_ ;
	assign \g53068/_0_  = _w3779_ ;
	assign \g53085/_0_  = _w4858_ ;
	assign \g53086/_0_  = _w4882_ ;
	assign \g53088/_0_  = _w4890_ ;
	assign \g53089/_0_  = _w4898_ ;
	assign \g53090/_0_  = _w4906_ ;
	assign \g53091/_0_  = _w4941_ ;
	assign \g53096/_0_  = _w4942_ ;
	assign \g53123/_0_  = _w3778_ ;
	assign \g53124/_0_  = _w4944_ ;
	assign \g53137/_0_  = _w4946_ ;
	assign \g53137/_1_  = _w4947_ ;
	assign \g53145/_0_  = _w4952_ ;
	assign \g53146/_0_  = _w4954_ ;
	assign \g53147/_0_  = _w4956_ ;
	assign \g53870/_0_  = _w4969_ ;
	assign \g53871/_0_  = _w4976_ ;
	assign \g53872/_0_  = _w4983_ ;
	assign \g53873/_0_  = _w4989_ ;
	assign \g53874/_0_  = _w4997_ ;
	assign \g53875/_0_  = _w5001_ ;
	assign \g53876/_0_  = _w5007_ ;
	assign \g53877/_0_  = _w5014_ ;
	assign \g53878/_0_  = _w5019_ ;
	assign \g53879/_0_  = _w5025_ ;
	assign \g53880/_0_  = _w5033_ ;
	assign \g53881/_0_  = _w5038_ ;
	assign \g53882/_0_  = _w5044_ ;
	assign \g53883/_0_  = _w5050_ ;
	assign \g53884/_0_  = _w5056_ ;
	assign \g53885/_0_  = _w5060_ ;
	assign \g53886/_0_  = _w5064_ ;
	assign \g53887/_0_  = _w5068_ ;
	assign \g53888/_0_  = _w5073_ ;
	assign \g53889/_0_  = _w5078_ ;
	assign \g53890/_3_  = _w5083_ ;
	assign \g53897/_3_  = _w5090_ ;
	assign \g53935/_3_  = _w5095_ ;
	assign \g53936/_3_  = _w5100_ ;
	assign \g53937/_3_  = _w5104_ ;
	assign \g53938/_3_  = _w5108_ ;
	assign \g53939/_3_  = _w5112_ ;
	assign \g53940/_3_  = _w5117_ ;
	assign \g53941/_3_  = _w5121_ ;
	assign \g53942/_3_  = _w5126_ ;
	assign \g54022/_0_  = _w5127_ ;
	assign \g54160/_3_  = _w4884_ ;
	assign \g54163/_3_  = _w4892_ ;
	assign \g54166/_3_  = _w4900_ ;
	assign \g54167/_2_  = _w5128_ ;
	assign \g54168/_3_  = _w5129_ ;
	assign \g54169/_3_  = _w5130_ ;
	assign \g54170/_3_  = _w5131_ ;
	assign \g54171/_2_  = _w5132_ ;
	assign \g54172/_3_  = _w5133_ ;
	assign \g54173/_3_  = _w5134_ ;
	assign \g54204/_2_  = _w5135_ ;
	assign \g54205/_2_  = _w5136_ ;
	assign \g54206/_2_  = _w5137_ ;
	assign \g54207/_2_  = _w5138_ ;
	assign \g54208/_2_  = _w5139_ ;
	assign \g54209/_2_  = _w5140_ ;
	assign \g54210/_2_  = _w5141_ ;
	assign \g54211/_2_  = _w5142_ ;
	assign \g54212/_2_  = _w5143_ ;
	assign \g54213/_2_  = _w5144_ ;
	assign \g54214/_2_  = _w5145_ ;
	assign \g54215/_2_  = _w5146_ ;
	assign \g54216/_2_  = _w5147_ ;
	assign \g54217/_2_  = _w5148_ ;
	assign \g54218/_2_  = _w5149_ ;
	assign \g54219/_2_  = _w5150_ ;
	assign \g54220/_2_  = _w5151_ ;
	assign \g54221/_2_  = _w5152_ ;
	assign \g54222/_2_  = _w5153_ ;
	assign \g54223/_2_  = _w5154_ ;
	assign \g54224/_2_  = _w5155_ ;
	assign \g54225/_2_  = _w5156_ ;
	assign \g54226/_2_  = _w5157_ ;
	assign \g54227/_2_  = _w5158_ ;
	assign \g54228/_2_  = _w5159_ ;
	assign \g54229/_2_  = _w5160_ ;
	assign \g54230/_2_  = _w5161_ ;
	assign \g54231/_2_  = _w5162_ ;
	assign \g54232/_2_  = _w5163_ ;
	assign \g54233/_2_  = _w5164_ ;
	assign \g54267/_0_  = _w5165_ ;
	assign \g54268/_0_  = _w5197_ ;
	assign \g54269/_0_  = _w5208_ ;
	assign \g54270/_0_  = _w5219_ ;
	assign \g54271/_0_  = _w5230_ ;
	assign \g54272/_0_  = _w5241_ ;
	assign \g54273/_0_  = _w5252_ ;
	assign \g54274/_0_  = _w5263_ ;
	assign \g54275/_0_  = _w5274_ ;
	assign \g54276/_0_  = _w5285_ ;
	assign \g54278/_0_  = _w5296_ ;
	assign \g54279/_0_  = _w5307_ ;
	assign \g54280/_0_  = _w5318_ ;
	assign \g54281/_0_  = _w5329_ ;
	assign \g54282/_0_  = _w5340_ ;
	assign \g54283/_0_  = _w5351_ ;
	assign \g54284/_0_  = _w5362_ ;
	assign \g54285/_0_  = _w5373_ ;
	assign \g54286/_0_  = _w5384_ ;
	assign \g54287/_0_  = _w5395_ ;
	assign \g54288/_0_  = _w5406_ ;
	assign \g54289/_0_  = _w5417_ ;
	assign \g54290/_0_  = _w5428_ ;
	assign \g54291/_0_  = _w5439_ ;
	assign \g54292/_0_  = _w5450_ ;
	assign \g54293/_0_  = _w5461_ ;
	assign \g54294/_0_  = _w5463_ ;
	assign \g54296/_0_  = _w5474_ ;
	assign \g54297/_0_  = _w5485_ ;
	assign \g54298/_0_  = _w5496_ ;
	assign \g54299/_0_  = _w5507_ ;
	assign \g54300/_0_  = _w5518_ ;
	assign \g54301/_0_  = _w5529_ ;
	assign \g54302/_0_  = _w5540_ ;
	assign \g54303/_0_  = _w5551_ ;
	assign \g54329/_0_  = _w5552_ ;
	assign \g54453/_0_  = _w5553_ ;
	assign \g54466/_0_  = _w5554_ ;
	assign \g54470/_0_  = _w3774_ ;
	assign \g54470/_1_  = _w3775_ ;
	assign \g54496/_0_  = _w5555_ ;
	assign \g54597/_0_  = _w5462_ ;
	assign \g54628/_0_  = _w5591_ ;
	assign \g54629/_0_  = _w5612_ ;
	assign \g54630/_0_  = _w5633_ ;
	assign \g54631/_0_  = _w5654_ ;
	assign \g54632/_0_  = _w5675_ ;
	assign \g54633/_0_  = _w5696_ ;
	assign \g54634/_0_  = _w5717_ ;
	assign \g54635/_0_  = _w5738_ ;
	assign \g54636/_0_  = _w5759_ ;
	assign \g54638/_0_  = _w5780_ ;
	assign \g54639/_0_  = _w5801_ ;
	assign \g54640/_0_  = _w5822_ ;
	assign \g54641/_0_  = _w5843_ ;
	assign \g54642/_0_  = _w5864_ ;
	assign \g54643/_0_  = _w5885_ ;
	assign \g54645/_0_  = _w5906_ ;
	assign \g54646/_0_  = _w5927_ ;
	assign \g54647/_0_  = _w5948_ ;
	assign \g54648/_0_  = _w5969_ ;
	assign \g54649/_0_  = _w5990_ ;
	assign \g54650/_0_  = _w6011_ ;
	assign \g54651/_0_  = _w6032_ ;
	assign \g54652/_0_  = _w6053_ ;
	assign \g54653/_0_  = _w6074_ ;
	assign \g54654/_0_  = _w6095_ ;
	assign \g54655/_0_  = _w6116_ ;
	assign \g54656/_0_  = _w6137_ ;
	assign \g54657/_0_  = _w6158_ ;
	assign \g54658/_0_  = _w6179_ ;
	assign \g54659/_0_  = _w6200_ ;
	assign \g54660/_0_  = _w6221_ ;
	assign \g54661/_0_  = _w6242_ ;
	assign \g54662/_0_  = _w6263_ ;
	assign \g54663/_0_  = _w6284_ ;
	assign \g54664/_0_  = _w6305_ ;
	assign \g54669/_0_  = _w6306_ ;
	assign \g54832/_0_  = _w6316_ ;
	assign \g54833/_0_  = _w6320_ ;
	assign \g54867/_0_  = _w6344_ ;
	assign \g54868/_0_  = _w6349_ ;
	assign \g54869/_0_  = _w6354_ ;
	assign \g54870/_0_  = _w6359_ ;
	assign \g54871/_0_  = _w6364_ ;
	assign \g54872/_0_  = _w6369_ ;
	assign \g54873/_0_  = _w6374_ ;
	assign \g54874/_0_  = _w6379_ ;
	assign \g54875/_0_  = _w6384_ ;
	assign \g54876/_0_  = _w6389_ ;
	assign \g54877/_0_  = _w6394_ ;
	assign \g54878/_0_  = _w6399_ ;
	assign \g54879/_0_  = _w6404_ ;
	assign \g54880/_0_  = _w6409_ ;
	assign \g54881/_0_  = _w6414_ ;
	assign \g54882/_0_  = _w6419_ ;
	assign \g54883/_0_  = _w6424_ ;
	assign \g54884/_0_  = _w6429_ ;
	assign \g54885/_0_  = _w6434_ ;
	assign \g54886/_0_  = _w6439_ ;
	assign \g54887/_0_  = _w6444_ ;
	assign \g54888/_0_  = _w6449_ ;
	assign \g54889/_0_  = _w6454_ ;
	assign \g54890/_0_  = _w6459_ ;
	assign \g54891/_0_  = _w6464_ ;
	assign \g54892/_0_  = _w6469_ ;
	assign \g54893/_0_  = _w6474_ ;
	assign \g54894/_0_  = _w6479_ ;
	assign \g54895/_0_  = _w6484_ ;
	assign \g54896/_0_  = _w6489_ ;
	assign \g54897/_0_  = _w6494_ ;
	assign \g54898/_0_  = _w6499_ ;
	assign \g54899/_0_  = _w6504_ ;
	assign \g56438/_0_  = _w6519_ ;
	assign \g56439/_0_  = _w6531_ ;
	assign \g56933/_3_  = _w6532_ ;
	assign \g56934/_3_  = _w6536_ ;
	assign \g56960/_0_  = _w6541_ ;
	assign \g56960/_1_  = _w6542_ ;
	assign \g56961/_3__syn_2  = _w6546_ ;
	assign \g57019/_0_  = _w6548_ ;
	assign \g57020/_0_  = _w6549_ ;
	assign \g57021/_0_  = _w6556_ ;
	assign \g57022/_0_  = _w6559_ ;
	assign \g57023/_0_  = _w6562_ ;
	assign \g57024/_0_  = _w6565_ ;
	assign \g57025/_0_  = _w6568_ ;
	assign \g57026/_0_  = _w6571_ ;
	assign \g57027/_0_  = _w6574_ ;
	assign \g57028/_0_  = _w6577_ ;
	assign \g57029/_0_  = _w6580_ ;
	assign \g57031/_0_  = _w6583_ ;
	assign \g57032/_0_  = _w6586_ ;
	assign \g57034/u3_syn_4  = _w6558_ ;
	assign \g57069/u3_syn_4  = _w6561_ ;
	assign \g57104/u3_syn_4  = _w6570_ ;
	assign \g57139/u3_syn_4  = _w6576_ ;
	assign \g57174/u3_syn_4  = _w6579_ ;
	assign \g57209/u3_syn_4  = _w6585_ ;
	assign \g57244/u3_syn_4  = _w6554_ ;
	assign \g57276/u3_syn_4  = _w6564_ ;
	assign \g57308/u3_syn_4  = _w6567_ ;
	assign \g57340/u3_syn_4  = _w6573_ ;
	assign \g57372/u3_syn_4  = _w6582_ ;
	assign \g57404/u3_syn_4  = _w6589_ ;
	assign \g57408/u3_syn_4  = _w6591_ ;
	assign \g57444/u3_syn_4  = _w6593_ ;
	assign \g57480/u3_syn_4  = _w6595_ ;
	assign \g57516/u3_syn_4  = _w6597_ ;
	assign \g57646/_0_  = _w6598_ ;
	assign \g57649/_0_  = _w6599_ ;
	assign \g57779/_3_  = _w6606_ ;
	assign \g57780/_3_  = _w6611_ ;
	assign \g57781/_3_  = _w6614_ ;
	assign \g57782/_3_  = _w6615_ ;
	assign \g57783/_3_  = _w6616_ ;
	assign \g57784/_3_  = _w6619_ ;
	assign \g57785/_3_  = _w6622_ ;
	assign \g57786/_3_  = _w6625_ ;
	assign \g57787/_3_  = _w6629_ ;
	assign \g57788/_3_  = _w6633_ ;
	assign \g57789/_3_  = _w6636_ ;
	assign \g57791/_3_  = _w6639_ ;
	assign \g57795/_3_  = _w6642_ ;
	assign \g57796/_3_  = _w6645_ ;
	assign \g57797/_3_  = _w6648_ ;
	assign \g57798/_3_  = _w6651_ ;
	assign \g57799/_3_  = _w6654_ ;
	assign \g57800/_3_  = _w6658_ ;
	assign \g57801/_3_  = _w6662_ ;
	assign \g57802/_3_  = _w6665_ ;
	assign \g57850/_0_  = _w6672_ ;
	assign \g57852/_0_  = _w6674_ ;
	assign \g57871/_0_  = _w6676_ ;
	assign \g57872/_0_  = _w6680_ ;
	assign \g57873/_0_  = _w6687_ ;
	assign \g58/_0_  = _w6708_ ;
	assign \g58490/_0_  = _w6709_ ;
	assign \g58564/_0_  = _w6710_ ;
	assign \g58569/_0_  = _w6715_ ;
	assign \g58571/_0_  = _w6717_ ;
	assign \g58573/_0_  = _w6718_ ;
	assign \g58577/_0_  = _w6721_ ;
	assign \g58578/_0_  = _w6722_ ;
	assign \g58579/_0_  = _w6728_ ;
	assign \g58580/_0_  = _w6730_ ;
	assign \g58583/_0_  = _w6749_ ;
	assign \g58584/_0_  = _w6751_ ;
	assign \g58603/_0_  = _w6752_ ;
	assign \g58611/_3_  = _w6758_ ;
	assign \g58637/_0_  = _w6762_ ;
	assign \g58638/_0_  = _w6764_ ;
	assign \g58639/_0_  = _w6765_ ;
	assign \g58691/_0_  = _w6767_ ;
	assign \g58693/_0_  = _w6768_ ;
	assign \g58696/_0_  = _w6770_ ;
	assign \g58700/_0_  = _w6771_ ;
	assign \g58701/_0_  = _w6772_ ;
	assign \g58708/_1_  = _w6555_ ;
	assign \g58730/_0_  = _w6773_ ;
	assign \g58731/_0_  = _w6774_ ;
	assign \g58732/_0_  = _w6775_ ;
	assign \g58733/_0_  = _w6776_ ;
	assign \g58734/_0_  = _w6777_ ;
	assign \g58735/_0_  = _w6779_ ;
	assign \g58736/_0_  = _w6781_ ;
	assign \g58737/_0_  = _w6783_ ;
	assign \g58738/_0_  = _w6785_ ;
	assign \g58739/_0_  = _w6787_ ;
	assign \g58740/_0_  = _w6789_ ;
	assign \g58741/_1__syn_2  = _w6675_ ;
	assign \g58748/_0_  = _w6790_ ;
	assign \g58751/_0_  = _w6791_ ;
	assign \g58752/_0_  = _w6792_ ;
	assign \g58753/_0_  = _w6793_ ;
	assign \g58754/_0_  = _w6794_ ;
	assign \g58756/_0_  = _w6797_ ;
	assign \g58767/_3_  = _w6798_ ;
	assign \g58768/_3_  = _w6799_ ;
	assign \g58769/_3_  = _w6800_ ;
	assign \g58770/_3_  = _w6801_ ;
	assign \g58771/_3_  = _w6802_ ;
	assign \g58772/_3_  = _w6803_ ;
	assign \g58773/_3_  = _w6804_ ;
	assign \g58774/_3_  = _w6805_ ;
	assign \g58775/_3_  = _w6806_ ;
	assign \g58776/_3_  = _w6807_ ;
	assign \g58777/_3_  = _w6808_ ;
	assign \g58778/_3_  = _w6809_ ;
	assign \g58779/_3_  = _w6810_ ;
	assign \g58780/_3_  = _w6811_ ;
	assign \g58781/_3_  = _w6812_ ;
	assign \g58782/_3_  = _w6813_ ;
	assign \g58783/_3_  = _w6814_ ;
	assign \g58784/_3_  = _w6815_ ;
	assign \g58785/_3_  = _w6816_ ;
	assign \g58786/_3_  = _w6817_ ;
	assign \g58787/_3_  = _w6818_ ;
	assign \g58788/_3_  = _w6819_ ;
	assign \g58789/_3_  = _w6820_ ;
	assign \g58790/_3_  = _w6821_ ;
	assign \g58791/_3_  = _w6822_ ;
	assign \g58792/_3_  = _w6823_ ;
	assign \g58793/_3_  = _w6824_ ;
	assign \g58794/_3_  = _w6825_ ;
	assign \g58795/_3_  = _w6826_ ;
	assign \g58796/_3_  = _w6827_ ;
	assign \g58797/_3_  = _w6828_ ;
	assign \g58798/_3_  = _w6829_ ;
	assign \g58874/_0_  = _w6841_ ;
	assign \g59064/_1_  = _w6552_ ;
	assign \g59072/_0_  = _w6842_ ;
	assign \g59080/_0_  = _w3229_ ;
	assign \g59083/_0_  = _w6845_ ;
	assign \g59084/_0_  = _w6847_ ;
	assign \g59085/_0_  = _w6850_ ;
	assign \g59088/_0_  = _w6852_ ;
	assign \g59094/_0_  = _w6853_ ;
	assign \g59095/_0_  = _w6854_ ;
	assign \g59126/_3_  = _w6857_ ;
	assign \g59128/_0_  = _w6883_ ;
	assign \g59174/_2_  = _w6683_ ;
	assign \g59180/_0_  = _w6884_ ;
	assign \g59181/_0_  = _w6885_ ;
	assign \g59182/_0_  = _w6886_ ;
	assign \g59190/_0_  = _w6937_ ;
	assign \g59191/_0_  = _w6940_ ;
	assign \g59192/_0_  = _w6944_ ;
	assign \g59204/_0_  = _w6952_ ;
	assign \g59205/_0_  = _w6957_ ;
	assign \g59210/_3_  = _w6962_ ;
	assign \g59213/_0_  = _w6963_ ;
	assign \g59214/_0_  = _w6964_ ;
	assign \g59215/_0_  = _w6965_ ;
	assign \g59216/_0_  = _w6966_ ;
	assign \g59217/_0_  = _w6967_ ;
	assign \g59218/_0_  = _w6968_ ;
	assign \g59219/_0_  = _w6969_ ;
	assign \g59220/_0_  = _w6970_ ;
	assign \g59221/_0_  = _w6971_ ;
	assign \g59222/_0_  = _w6972_ ;
	assign \g59223/_0_  = _w6973_ ;
	assign \g59226/_3_  = _w6976_ ;
	assign \g59232/_00_  = _w6978_ ;
	assign \g59233/_0_  = _w6980_ ;
	assign \g59235/_0_  = _w6981_ ;
	assign \g59236/_0_  = _w6982_ ;
	assign \g59237/_0_  = _w6983_ ;
	assign \g59238/_0_  = _w6984_ ;
	assign \g59318/_0_  = _w6985_ ;
	assign \g59331/_0_  = _w6848_ ;
	assign \g59336/_0_  = _w6990_ ;
	assign \g59351/_0_  = _w6998_ ;
	assign \g59354/_0_  = _w7001_ ;
	assign \g59358/_0_  = _w7014_ ;
	assign \g59363/_0_  = _w7015_ ;
	assign \g59366/_0_  = _w7021_ ;
	assign \g59370/u3_syn_4  = _w7024_ ;
	assign \g59371/u3_syn_4  = _w7026_ ;
	assign \g59372/u3_syn_4  = _w7028_ ;
	assign \g59373/u3_syn_4  = _w7030_ ;
	assign \g59378/u3_syn_4  = _w7032_ ;
	assign \g59379/u3_syn_4  = _w7034_ ;
	assign \g59380/u3_syn_4  = _w7036_ ;
	assign \g59381/u3_syn_4  = _w7038_ ;
	assign \g59589/_0_  = _w7042_ ;
	assign \g59655/_0_  = _w7043_ ;
	assign \g59662/_0_  = _w3105_ ;
	assign \g59735/_0_  = _w7049_ ;
	assign \g59739/_0_  = _w7052_ ;
	assign \g59740/_0_  = _w7054_ ;
	assign \g59741/_0_  = _w7056_ ;
	assign \g59742/_0_  = _w7060_ ;
	assign \g59743/_0_  = _w7062_ ;
	assign \g59744/_0_  = _w7064_ ;
	assign \g59745/_0_  = _w7066_ ;
	assign \g59746/_0_  = _w7070_ ;
	assign \g59747/_0_  = _w7071_ ;
	assign \g59748/_0_  = _w7075_ ;
	assign \g59749/_0_  = _w7076_ ;
	assign \g59750/_0_  = _w7077_ ;
	assign \g59751/_0_  = _w7078_ ;
	assign \g59752/_0_  = _w7079_ ;
	assign \g59753/_0_  = _w7080_ ;
	assign \g59754/_0_  = _w7081_ ;
	assign \g59755/_0_  = _w7082_ ;
	assign \g59756/_0_  = _w7084_ ;
	assign \g59757/_0_  = _w7086_ ;
	assign \g59758/_0_  = _w7092_ ;
	assign \g59759/_0_  = _w7094_ ;
	assign \g59760/_0_  = _w7096_ ;
	assign \g59764/_0_  = _w7102_ ;
	assign \g59766/_0_  = _w7105_ ;
	assign \g59774/_0_  = _w7107_ ;
	assign \g59775/_0_  = _w7109_ ;
	assign \g59776/_0_  = _w7111_ ;
	assign \g59777/_0_  = _w7113_ ;
	assign \g59778/_0_  = _w7115_ ;
	assign \g59779/_0_  = _w7117_ ;
	assign \g59780/_0_  = _w7119_ ;
	assign \g59781/_0_  = _w7121_ ;
	assign \g59789/_3_  = _w7126_ ;
	assign \g59799/_3_  = _w7127_ ;
	assign \g60311/_0_  = _w6738_ ;
	assign \g60326/_0_  = _w7128_ ;
	assign \g60333/_0_  = _w7129_ ;
	assign \g60336/_3_  = _w3665_ ;
	assign \g60341/_0_  = _w7131_ ;
	assign \g60343/_0_  = _w7133_ ;
	assign \g60344/_0_  = _w7141_ ;
	assign \g60345/_0_  = _w7143_ ;
	assign \g60354/_0_  = _w7145_ ;
	assign \g60355/_0_  = _w7147_ ;
	assign \g60356/_0_  = _w7149_ ;
	assign \g60357/_0_  = _w7151_ ;
	assign \g60358/_0_  = _w7154_ ;
	assign \g60359/_0_  = _w7159_ ;
	assign \g60360/_0_  = _w7160_ ;
	assign \g60361/_0_  = _w7163_ ;
	assign \g60362/_0_  = _w7166_ ;
	assign \g60363/_0_  = _w7169_ ;
	assign \g60364/_0_  = _w7172_ ;
	assign \g60398/_2_  = _w3800_ ;
	assign \g60399/_0_  = _w7175_ ;
	assign \g60400/_0_  = _w7176_ ;
	assign \g60401/_0_  = _w7177_ ;
	assign \g60402/_0_  = _w7178_ ;
	assign \g60403/_0_  = _w7179_ ;
	assign \g60406/_0_  = _w7184_ ;
	assign \g60410/_0_  = _w7185_ ;
	assign \g60411/_0_  = _w7191_ ;
	assign \g60417/_3_  = _w7195_ ;
	assign \g60419/_3_  = _w7199_ ;
	assign \g60421/_3_  = _w7200_ ;
	assign \g60423/_3_  = _w7201_ ;
	assign \g60425/_3_  = _w7202_ ;
	assign \g60427/_3_  = _w7206_ ;
	assign \g60429/_3_  = _w7209_ ;
	assign \g60431/_3_  = _w7212_ ;
	assign \g60433/_3_  = _w7213_ ;
	assign \g60435/_3_  = _w7215_ ;
	assign \g60437/_3_  = _w7218_ ;
	assign \g60439/_3_  = _w7221_ ;
	assign \g60441/_3_  = _w7224_ ;
	assign \g60443/_3_  = _w7225_ ;
	assign \g60445/_3_  = _w7228_ ;
	assign \g60447/_3_  = _w7231_ ;
	assign \g60449/_3_  = _w7234_ ;
	assign \g60451/_3_  = _w7235_ ;
	assign \g60453/_3_  = _w7238_ ;
	assign \g60455/_3_  = _w7239_ ;
	assign \g60457/_3_  = _w7242_ ;
	assign \g60459/_3_  = _w7243_ ;
	assign \g60461/_3_  = _w7246_ ;
	assign \g60463/_3_  = _w7247_ ;
	assign \g60465/_3_  = _w7248_ ;
	assign \g60467/_3_  = _w7252_ ;
	assign \g60469/_3_  = _w7253_ ;
	assign \g60471/_3_  = _w7254_ ;
	assign \g60473/_3_  = _w7255_ ;
	assign \g60475/_3_  = _w7256_ ;
	assign \g60477/_3_  = _w7257_ ;
	assign \g60479/_3_  = _w7258_ ;
	assign \g60481/_3_  = _w7261_ ;
	assign \g60483/_3_  = _w7262_ ;
	assign \g60485/_3_  = _w7263_ ;
	assign \g60487/_3_  = _w7264_ ;
	assign \g60489/_3_  = _w7267_ ;
	assign \g60491/_3_  = _w7270_ ;
	assign \g60493/_3_  = _w7273_ ;
	assign \g60495/_3_  = _w7276_ ;
	assign \g60497/_3_  = _w7277_ ;
	assign \g60499/_3_  = _w7280_ ;
	assign \g60501/_3_  = _w7283_ ;
	assign \g60503/_3_  = _w7286_ ;
	assign \g60505/_3_  = _w7289_ ;
	assign \g60507/_3_  = _w7290_ ;
	assign \g60509/_3_  = _w7293_ ;
	assign \g60511/_3_  = _w7296_ ;
	assign \g60513/_3_  = _w7299_ ;
	assign \g60515/_3_  = _w7300_ ;
	assign \g60517/_3_  = _w7301_ ;
	assign \g60519/_3_  = _w7304_ ;
	assign \g60521/_3_  = _w7307_ ;
	assign \g60523/_3_  = _w7310_ ;
	assign \g60525/_3_  = _w7311_ ;
	assign \g60527/_3_  = _w7314_ ;
	assign \g60529/_3_  = _w7315_ ;
	assign \g60531/_3_  = _w7316_ ;
	assign \g60533/_3_  = _w7317_ ;
	assign \g60535/_3_  = _w7320_ ;
	assign \g60537/_3_  = _w7323_ ;
	assign \g60539/_3_  = _w7326_ ;
	assign \g60541/_3_  = _w7327_ ;
	assign \g60544/_3_  = _w7328_ ;
	assign \g60546/_3_  = _w7329_ ;
	assign \g60548/_3_  = _w7332_ ;
	assign \g60550/_3_  = _w7335_ ;
	assign \g60552/_3_  = _w7338_ ;
	assign \g60554/_3_  = _w7341_ ;
	assign \g60556/_3_  = _w7342_ ;
	assign \g60559/_3_  = _w7345_ ;
	assign \g60561/_3_  = _w7348_ ;
	assign \g60563/_3_  = _w7351_ ;
	assign \g60565/_3_  = _w7354_ ;
	assign \g60567/_3_  = _w7357_ ;
	assign \g60569/_3_  = _w7360_ ;
	assign \g60571/_3_  = _w7363_ ;
	assign \g60573/_3_  = _w7366_ ;
	assign \g60575/_3_  = _w7369_ ;
	assign \g60577/_3_  = _w7372_ ;
	assign \g60579/_3_  = _w7375_ ;
	assign \g60581/_3_  = _w7378_ ;
	assign \g60583/_3_  = _w7381_ ;
	assign \g60585/_3_  = _w7384_ ;
	assign \g60588/_3_  = _w7387_ ;
	assign \g60590/_3_  = _w7390_ ;
	assign \g60593/_3_  = _w7393_ ;
	assign \g60596/_3_  = _w7396_ ;
	assign \g60598/_3_  = _w7400_ ;
	assign \g60600/_3_  = _w7403_ ;
	assign \g60602/_3_  = _w7406_ ;
	assign \g60603/_3_  = _w7409_ ;
	assign \g60671/_3_  = _w7412_ ;
	assign \g60672/_3_  = _w7413_ ;
	assign \g60674/_3_  = _w7414_ ;
	assign \g60680/_0_  = _w7418_ ;
	assign \g60682/_3_  = _w7419_ ;
	assign \g60690/_3_  = _w7422_ ;
	assign \g60692/_3_  = _w7424_ ;
	assign \g61594/_0_  = _w7426_ ;
	assign \g61614/_0_  = _w7429_ ;
	assign \g61618/_00_  = _w7431_ ;
	assign \g61649/_0_  = _w7434_ ;
	assign \g61651/_0_  = _w7436_ ;
	assign \g61656/_0_  = _w7440_ ;
	assign \g61657/_0_  = _w7442_ ;
	assign \g61659/_0_  = _w7445_ ;
	assign \g61662/_0_  = _w7447_ ;
	assign \g61663/_0_  = _w7498_ ;
	assign \g61664/_0_  = _w7500_ ;
	assign \g61665/_0_  = _w7505_ ;
	assign \g61667/_2_  = _w6838_ ;
	assign \g61669/_3__syn_2  = _w7512_ ;
	assign \g61678/_0_  = _w7513_ ;
	assign \g61679/_0_  = _w7514_ ;
	assign \g61680/_0_  = _w7515_ ;
	assign \g61681/_0_  = _w7516_ ;
	assign \g61684/_0_  = _w7517_ ;
	assign \g61685/_0_  = _w7518_ ;
	assign \g61686/_0_  = _w7519_ ;
	assign \g61690/_0_  = _w7522_ ;
	assign \g61692/_0_  = _w7523_ ;
	assign \g61694/_0_  = _w7526_ ;
	assign \g61695/_0_  = _w7528_ ;
	assign \g61696/_0_  = _w7530_ ;
	assign \g61699/u3_syn_4  = _w7531_ ;
	assign \g61732/u3_syn_4  = _w7533_ ;
	assign \g61765/u3_syn_4  = _w7535_ ;
	assign \g61798/u3_syn_4  = _w7536_ ;
	assign \g61848/_0_  = _w7542_ ;
	assign \g61848/_3_  = _w7541_ ;
	assign \g61853/_0_  = _w7543_ ;
	assign \g61854/_1__syn_2  = _w3021_ ;
	assign \g61858/u3_syn_4  = _w7544_ ;
	assign \g61880/u3_syn_4  = _w3618_ ;
	assign \g61887/u3_syn_4  = _w7545_ ;
	assign \g61920/u3_syn_4  = _w7546_ ;
	assign \g61990/u3_syn_4  = _w7547_ ;
	assign \g62254/_0__syn_2  = _w7123_ ;
	assign \g62260/_0_  = _w7548_ ;
	assign \g62262/_1__syn_2  = _w7004_ ;
	assign \g62290/_0_  = _w7549_ ;
	assign \g62317/_0_  = _w7551_ ;
	assign \g62319/_0_  = _w7553_ ;
	assign \g62324/_0_  = _w7555_ ;
	assign \g62329/_0_  = _w6711_ ;
	assign \g62331/_0_  = _w7556_ ;
	assign \g62331/_1_  = _w7557_ ;
	assign \g62333/u3_syn_4  = _w7559_ ;
	assign \g62335/u3_syn_4  = _w7561_ ;
	assign \g62336/u3_syn_4  = _w7563_ ;
	assign \g62428/u3_syn_4  = _w7565_ ;
	assign \g62454/u3_syn_4  = _w7567_ ;
	assign \g62487/u3_syn_4  = _w7569_ ;
	assign \g62520/u3_syn_4  = _w7571_ ;
	assign \g62552/u3_syn_4  = _w7573_ ;
	assign \g62584/u3_syn_4  = _w7575_ ;
	assign \g62619/u3_syn_4  = _w7577_ ;
	assign \g62651/u3_syn_4  = _w7579_ ;
	assign \g62692/_0_  = _w7582_ ;
	assign \g62873/_0_  = _w7583_ ;
	assign \g62882/_0_  = _w7584_ ;
	assign \g62883/u3_syn_4  = _w7586_ ;
	assign \g62886/u3_syn_4  = _w7588_ ;
	assign \g62908/u3_syn_4  = _w7590_ ;
	assign \g62952/u3_syn_4  = _w7592_ ;
	assign \g62974/u3_syn_4  = _w7593_ ;
	assign \g63207/_0_  = _w7594_ ;
	assign \g63214/_3_  = _w3209_ ;
	assign \g63227/_0_  = _w3975_ ;
	assign \g63250/_1__syn_2  = _w7181_ ;
	assign \g63315/_0__syn_2  = _w4950_ ;
	assign \g63320/_0_  = _w7596_ ;
	assign \g63322/_0_  = _w7597_ ;
	assign \g63324/_2_  = _w7598_ ;
	assign \g63338/_0__syn_2  = _w7599_ ;
	assign \g63340/_0_  = _w7606_ ;
	assign \g63376/_0_  = _w7607_ ;
	assign \g63395/_2_  = _w7608_ ;
	assign \g63398/_0_  = _w7609_ ;
	assign \g63419/_0_  = _w7611_ ;
	assign \g63524/_3_  = _w7504_ ;
	assign \g63540/_0_  = _w7612_ ;
	assign \g63541/_0_  = _w7613_ ;
	assign \g63682/_0_  = _w7618_ ;
	assign \g63890/_1_  = _w7554_ ;
	assign \g63892/_0_  = _w7621_ ;
	assign \g63894/_0_  = _w7623_ ;
	assign \g63897/_1_  = _w3797_ ;
	assign \g63908/_0_  = _w7624_ ;
	assign \g63913/_0_  = _w7625_ ;
	assign \g63914/_0_  = _w7626_ ;
	assign \g63927/_1__syn_2  = _w7550_ ;
	assign \g63934/_0_  = _w7628_ ;
	assign \g63942/_0_  = _w7629_ ;
	assign \g63952/_0_  = _w6637_ ;
	assign \g63965/_0_  = _w7631_ ;
	assign \g63969/_0_  = _w7537_ ;
	assign \g63985/_0_  = _w7635_ ;
	assign \g63986/_0_  = _w7638_ ;
	assign \g63987/_0_  = _w7641_ ;
	assign \g63988/_0_  = _w7644_ ;
	assign \g63990/_0_  = _w7647_ ;
	assign \g63991/_0_  = _w7650_ ;
	assign \g63992/_0_  = _w7653_ ;
	assign \g63993/_0_  = _w7656_ ;
	assign \g64016/_0_  = _w7659_ ;
	assign \g64017/_0_  = _w7662_ ;
	assign \g64018/_0_  = _w7665_ ;
	assign \g64019/_0_  = _w7668_ ;
	assign \g64020/_0_  = _w7671_ ;
	assign \g64021/_0_  = _w7674_ ;
	assign \g64023/_0_  = _w7677_ ;
	assign \g64024/_0_  = _w7680_ ;
	assign \g64101/_0_  = _w7683_ ;
	assign \g64104/_0_  = _w7686_ ;
	assign \g64121/_0_  = _w7689_ ;
	assign \g64174/_0_  = _w7692_ ;
	assign \g64249/_0_  = _w7695_ ;
	assign \g64299/_0_  = _w7698_ ;
	assign \g64338/_0_  = _w7701_ ;
	assign \g64364/_0_  = _w7704_ ;
	assign \g64459/_0_  = _w7705_ ;
	assign \g64461/_0_  = _w6609_ ;
	assign \g64466/_0_  = _w7706_ ;
	assign \g64577/_0_  = _w7022_ ;
	assign \g64583/_0_  = _w6314_ ;
	assign \g64589/_1_  = _w7507_ ;
	assign \g64595/_0_  = _w7707_ ;
	assign \g64598/_0_  = _w7709_ ;
	assign \g64649/_0_  = _w7710_ ;
	assign \g64678/_0_  = _w7712_ ;
	assign \g64688/_3_  = _w3134_ ;
	assign \g64689/_0_  = _w7715_ ;
	assign \g64694/_0_  = _w7716_ ;
	assign \g64695/_0_  = _w7717_ ;
	assign \g64700/_0_  = _w7719_ ;
	assign \g64714/_0_  = _w7720_ ;
	assign \g64744/_2_  = _w7721_ ;
	assign \g65255/_0_  = _w7722_ ;
	assign \g65258/_0_  = _w7723_ ;
	assign \g65269/_3_  = _w7724_ ;
	assign \g65489/_0_  = _w6947_ ;
	assign \g65513/_0_  = _w6945_ ;
	assign \g65530/_0_  = _w7725_ ;
	assign \g65561/_0_  = _w7538_ ;
	assign \g65563/_0_  = _w7726_ ;
	assign \g65564/_0_  = _w7727_ ;
	assign \g65573/_0_  = _w7728_ ;
	assign \g65578/_2_  = _w3793_ ;
	assign \g65597/_0_  = _w7729_ ;
	assign \g65605/_0_  = _w7732_ ;
	assign \g65606/_0_  = _w7734_ ;
	assign \g65609/_0_  = _w7737_ ;
	assign \g65611/_0_  = _w7740_ ;
	assign \g65612/_0_  = _w7743_ ;
	assign \g65613/_0_  = _w7746_ ;
	assign \g65615/_0_  = _w7749_ ;
	assign \g65618/_0_  = _w7752_ ;
	assign \g65631/_0_  = _w7755_ ;
	assign \g65634/_0_  = _w7758_ ;
	assign \g65635/_0_  = _w7759_ ;
	assign \g65639/_0_  = _w7760_ ;
	assign \g65644/_0_  = _w7763_ ;
	assign \g65648/_0_  = _w7766_ ;
	assign \g65650/_0_  = _w7769_ ;
	assign \g65662/_3_  = _w7772_ ;
	assign \g65665/_3_  = _w7775_ ;
	assign \g65729/_0_  = _w7776_ ;
	assign \g65801/_0_  = _w6604_ ;
	assign \g66072/_0_  = _w7777_ ;
	assign \g66074/_0_  = _w7778_ ;
	assign \g66075/_0_  = _w7779_ ;
	assign \g66076/_0_  = _w7780_ ;
	assign \g66077/_0_  = _w7781_ ;
	assign \g66078/_0_  = _w7782_ ;
	assign \g66079/_0_  = _w7783_ ;
	assign \g66080/_0_  = _w7784_ ;
	assign \g66081/_0_  = _w7785_ ;
	assign \g66082/_0_  = _w7786_ ;
	assign \g66085/_0_  = _w7787_ ;
	assign \g66086/_0_  = _w7788_ ;
	assign \g66087/_0_  = _w7789_ ;
	assign \g66089/_0_  = _w7790_ ;
	assign \g66090/_0_  = _w7791_ ;
	assign \g66093/_0_  = _w7792_ ;
	assign \g66094/_0_  = _w7793_ ;
	assign \g66095/_0_  = _w7794_ ;
	assign \g66098/_0_  = _w7795_ ;
	assign \g66100/_0_  = _w7796_ ;
	assign \g66106/_1_  = _w3224_ ;
	assign \g66107/_0_  = _w7797_ ;
	assign \g66108/_0_  = _w7798_ ;
	assign \g66110/_0_  = _w7799_ ;
	assign \g66114/_0_  = _w3257_ ;
	assign \g66124/_0_  = _w7800_ ;
	assign \g66125/_0_  = _w7801_ ;
	assign \g66127/_0_  = _w7802_ ;
	assign \g66128/_0_  = _w7803_ ;
	assign \g66129/_0_  = _w7804_ ;
	assign \g66130/_0_  = _w7805_ ;
	assign \g66133/_0_  = _w7806_ ;
	assign \g66134/_0_  = _w7807_ ;
	assign \g66136/_0_  = _w7808_ ;
	assign \g66141/_1_  = _w7809_ ;
	assign \g66153/_0_  = _w7810_ ;
	assign \g66182/_0_  = _w3645_ ;
	assign \g66187/_0_  = _w6544_ ;
	assign \g66240/_0_  = _w7814_ ;
	assign \g66268/_0_  = _w7815_ ;
	assign \g66354/_0_  = _w7816_ ;
	assign \g66397/_3_  = _w7817_ ;
	assign \g66398/_3_  = _w7818_ ;
	assign \g66399/_3_  = _w7819_ ;
	assign \g66400/_3_  = _w7820_ ;
	assign \g66401/_3_  = _w7821_ ;
	assign \g66402/_3_  = _w7822_ ;
	assign \g66403/_3_  = _w7823_ ;
	assign \g66404/_3_  = _w7824_ ;
	assign \g66405/_3_  = _w7825_ ;
	assign \g66406/_3_  = _w7826_ ;
	assign \g66407/_3_  = _w7827_ ;
	assign \g66408/_3_  = _w7828_ ;
	assign \g66409/_3_  = _w7829_ ;
	assign \g66410/_3_  = _w7830_ ;
	assign \g66411/_3_  = _w7831_ ;
	assign \g66412/_3_  = _w7832_ ;
	assign \g66413/_3_  = _w7833_ ;
	assign \g66414/_3_  = _w7834_ ;
	assign \g66415/_3_  = _w7835_ ;
	assign \g66416/_3_  = _w7836_ ;
	assign \g66417/_3_  = _w7837_ ;
	assign \g66418/_3_  = _w7838_ ;
	assign \g66419/_3_  = _w7839_ ;
	assign \g66420/_3_  = _w7840_ ;
	assign \g66421/_3_  = _w7841_ ;
	assign \g66422/_3_  = _w7842_ ;
	assign \g66423/_3_  = _w7843_ ;
	assign \g66424/_3_  = _w7844_ ;
	assign \g66425/_3_  = _w7845_ ;
	assign \g66426/_3_  = _w7846_ ;
	assign \g66427/_3_  = _w7847_ ;
	assign \g66428/_3_  = _w7848_ ;
	assign \g66429/_3_  = _w7849_ ;
	assign \g66430/_3_  = _w7850_ ;
	assign \g66464/_0_  = _w7851_ ;
	assign \g66465/_0_  = _w7852_ ;
	assign \g66477/_3_  = _w6992_ ;
	assign \g66643/_0_  = _w3794_ ;
	assign \g66733/_2_  = _w3212_ ;
	assign \g66735/_1_  = _w3204_ ;
	assign \g66801/_0_  = _w7853_ ;
	assign \g66866/_0_  = _w7854_ ;
	assign \g66875/_0_  = _w7855_ ;
	assign \g66885/_1_  = _w7856_ ;
	assign \g66890/_0_  = _w7857_ ;
	assign \g66939/_0_  = _w7615_ ;
	assign \g66950/_0_  = _w7858_ ;
	assign \g67035/_0_  = _w7859_ ;
	assign \g67038/_0_  = _w7860_ ;
	assign \g67044/_3_  = _w6858_ ;
	assign \g67045/_3_  = _w6870_ ;
	assign \g67046/_3_  = _w6868_ ;
	assign \g67070/_3_  = _w6861_ ;
	assign \g67082/_3_  = _w3790_ ;
	assign \g67090/_3_  = _w6308_ ;
	assign \g67106/_0_  = _w7861_ ;
	assign \g67107/_0_  = _w7862_ ;
	assign \g67108/_0_  = _w7863_ ;
	assign \g67109/_0_  = _w7864_ ;
	assign \g67117/_0_  = _w7865_ ;
	assign \g67131/_0_  = _w7866_ ;
	assign \g67142/_0_  = _w7867_ ;
	assign \g67421/_0_  = _w6323_ ;
	assign \g67456/_0_  = _w7811_ ;
	assign \g67464/_0_  = _w7868_ ;
	assign \g67617/_1_  = _w7812_ ;
	assign \g67772/_0_  = _w7869_ ;
	assign \g68523/_0_  = _w452_ ;
	assign \g73970/_0_  = _w7872_ ;
	assign \g73976/_0_  = _w3074_ ;
	assign \g74120/_1_  = _w3216_ ;
	assign \g74148/_2_  = _w6328_ ;
	assign \g74245/_0_  = _w7893_ ;
	assign \g74426/_0_  = _w7894_ ;
	assign \g74434/_3_  = _w3207_ ;
	assign \g74589/_0_  = _w7905_ ;
	assign \g74626/_1__syn_2  = _w3022_ ;
	assign \g74790/_0_  = _w3096_ ;
	assign \g74801/_0_  = _w7916_ ;
	assign \g74838/_0_  = _w7927_ ;
	assign \g74850/_0_  = _w7938_ ;
	assign \g74855/_0_  = _w7949_ ;
	assign \g74862/_0_  = _w7960_ ;
	assign \g74871/_0_  = _w7971_ ;
	assign \g74878/_0_  = _w7982_ ;
	assign \g74885/_0_  = _w7993_ ;
	assign \g74922/_0_  = _w7996_ ;
	assign \g75066/_1__syn_2  = _w7997_ ;
	assign \g75100/_1_  = _w3081_ ;
	assign \g75201/_1_  = _w5558_ ;
	assign \g75205/_1_  = _w3031_ ;
	assign \g75420/_1_  = _w4478_ ;
	assign pci_rst_oe_o_pad = 1'b1;
	assign wb_int_o_pad = 1'b0;
	assign wb_rst_o_pad = _w7998_ ;
endmodule;